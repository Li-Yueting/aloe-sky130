magic
tech sky130A
magscale 1 2
timestamp 1654748007
<< pwell >>
rect -2706 -970 2608 526
<< psubdiff >>
rect -2668 -840 -2628 -800
rect -2668 -920 -2628 -880
rect -1610 -872 -1490 -870
rect -1610 -908 -1570 -872
rect -1526 -908 -1490 -872
rect -1610 -920 -1490 -908
rect -310 -872 -190 -870
rect -310 -908 -270 -872
rect -226 -908 -190 -872
rect -310 -920 -190 -908
rect 990 -872 1110 -870
rect 990 -908 1030 -872
rect 1074 -908 1110 -872
rect 990 -920 1110 -908
<< psubdiffcont >>
rect -2668 -880 -2628 -840
rect -1570 -908 -1526 -872
rect -270 -908 -226 -872
rect 1030 -908 1074 -872
<< poly >>
rect -2488 -716 -2368 -466
rect -2232 -716 -2112 -466
rect -1976 -716 -1856 -466
rect -1720 -716 -1600 -466
rect -1464 -716 -1344 -466
rect -1208 -716 -1088 -466
rect -952 -716 -832 -466
rect -696 -716 -576 -466
rect -440 -716 -320 -466
rect -184 -716 -64 -466
rect 72 -716 192 -466
rect 328 -716 448 -466
rect 584 -716 704 -466
rect 840 -716 960 -466
rect 1096 -716 1216 -466
rect 1352 -716 1472 -466
rect 1608 -716 1728 -466
rect 1864 -716 1984 -466
rect 2120 -716 2240 -466
rect 2376 -716 2496 -466
rect -2528 -736 2608 -716
rect -2528 -796 -2438 -736
rect -2378 -796 -2238 -736
rect -2178 -796 -2038 -736
rect -1978 -796 -1838 -736
rect -1778 -796 -1638 -736
rect -1578 -796 -1438 -736
rect -1378 -796 -1238 -736
rect -1178 -796 -1038 -736
rect -978 -796 -838 -736
rect -778 -796 -638 -736
rect -578 -796 -438 -736
rect -378 -796 -238 -736
rect -178 -796 -38 -736
rect 22 -796 162 -736
rect 222 -796 362 -736
rect 422 -796 562 -736
rect 622 -796 762 -736
rect 822 -796 962 -736
rect 1022 -796 1162 -736
rect 1222 -796 1362 -736
rect 1422 -796 1562 -736
rect 1622 -796 1762 -736
rect 1822 -796 1962 -736
rect 2022 -796 2162 -736
rect 2222 -796 2362 -736
rect 2422 -796 2608 -736
rect -2528 -816 2608 -796
<< polycont >>
rect -2438 -796 -2378 -736
rect -2238 -796 -2178 -736
rect -2038 -796 -1978 -736
rect -1838 -796 -1778 -736
rect -1638 -796 -1578 -736
rect -1438 -796 -1378 -736
rect -1238 -796 -1178 -736
rect -1038 -796 -978 -736
rect -838 -796 -778 -736
rect -638 -796 -578 -736
rect -438 -796 -378 -736
rect -238 -796 -178 -736
rect -38 -796 22 -736
rect 162 -796 222 -736
rect 362 -796 422 -736
rect 562 -796 622 -736
rect 762 -796 822 -736
rect 962 -796 1022 -736
rect 1162 -796 1222 -736
rect 1362 -796 1422 -736
rect 1562 -796 1622 -736
rect 1762 -796 1822 -736
rect 1962 -796 2022 -736
rect 2162 -796 2222 -736
rect 2362 -796 2422 -736
<< locali >>
rect -2706 850 -2438 910
rect -2378 850 -2238 910
rect -2178 850 -2038 910
rect -1978 850 -1838 910
rect -1778 850 -1638 910
rect -1578 850 -1438 910
rect -1378 850 -1238 910
rect -1178 850 -1038 910
rect -978 850 -838 910
rect -778 850 -638 910
rect -578 850 -438 910
rect -378 850 -238 910
rect -178 850 -38 910
rect 22 850 162 910
rect 222 850 362 910
rect 422 850 562 910
rect 622 850 762 910
rect 822 850 962 910
rect 1022 850 1162 910
rect 1222 850 1362 910
rect 1422 850 1562 910
rect 1622 850 1762 910
rect 1822 850 1962 910
rect 2022 850 2162 910
rect 2222 850 2362 910
rect 2422 850 2608 910
rect -2608 690 2608 750
rect -2339 486 -2305 690
rect -1823 486 -1789 690
rect -1307 486 -1273 690
rect -791 486 -757 690
rect -275 486 -241 690
rect 241 486 275 690
rect 757 486 791 690
rect 1273 486 1307 690
rect 1789 486 1823 690
rect 2305 486 2339 690
rect -2597 -470 -2563 -446
rect -2081 -470 -2047 -446
rect -1565 -470 -1531 -446
rect -1049 -470 -1015 -446
rect -533 -470 -499 -446
rect -17 -470 17 -446
rect 499 -470 533 -446
rect 1015 -470 1049 -446
rect 1531 -470 1565 -446
rect 2047 -470 2081 -446
rect -2608 -530 2608 -470
rect -2678 -840 -2618 -760
rect -2528 -796 -2438 -736
rect -2378 -796 -2238 -736
rect -2178 -796 -2038 -736
rect -1978 -796 -1838 -736
rect -1778 -796 -1638 -736
rect -1578 -796 -1438 -736
rect -1378 -796 -1238 -736
rect -1178 -796 -1038 -736
rect -978 -796 -838 -736
rect -778 -796 -638 -736
rect -578 -796 -438 -736
rect -378 -796 -238 -736
rect -178 -796 -38 -736
rect 22 -796 162 -736
rect 222 -796 362 -736
rect 422 -796 562 -736
rect 622 -796 762 -736
rect 822 -796 962 -736
rect 1022 -796 1162 -736
rect 1222 -796 1362 -736
rect 1422 -796 1562 -736
rect 1622 -796 1762 -736
rect 1822 -796 1962 -736
rect 2022 -796 2162 -736
rect 2222 -796 2362 -736
rect 2422 -796 2608 -736
rect -2678 -880 -2668 -840
rect -2628 -880 -2618 -840
rect -2678 -970 -2618 -880
rect -1630 -872 -1470 -850
rect -1630 -908 -1570 -872
rect -1526 -908 -1470 -872
rect -1630 -970 -1470 -908
rect -330 -872 -170 -850
rect -330 -908 -270 -872
rect -226 -908 -170 -872
rect -330 -970 -170 -908
rect 970 -872 1130 -850
rect 970 -908 1030 -872
rect 1074 -908 1130 -872
rect 970 -970 1130 -908
rect -2706 -1030 -2438 -970
rect -2378 -1030 -2238 -970
rect -2178 -1030 -2038 -970
rect -1978 -1030 -1838 -970
rect -1778 -1030 -1638 -970
rect -1578 -1030 -1438 -970
rect -1378 -1030 -1238 -970
rect -1178 -1030 -1038 -970
rect -978 -1030 -838 -970
rect -778 -1030 -638 -970
rect -578 -1030 -438 -970
rect -378 -1030 -238 -970
rect -178 -1030 -38 -970
rect 22 -1030 162 -970
rect 222 -1030 362 -970
rect 422 -1030 562 -970
rect 622 -1030 762 -970
rect 822 -1030 962 -970
rect 1022 -1030 1162 -970
rect 1222 -1030 1362 -970
rect 1422 -1030 1562 -970
rect 1622 -1030 1762 -970
rect 1822 -1030 1962 -970
rect 2022 -1030 2162 -970
rect 2222 -1030 2362 -970
rect 2422 -1030 2608 -970
<< viali >>
rect -2438 850 -2378 910
rect -2238 850 -2178 910
rect -2038 850 -1978 910
rect -1838 850 -1778 910
rect -1638 850 -1578 910
rect -1438 850 -1378 910
rect -1238 850 -1178 910
rect -1038 850 -978 910
rect -838 850 -778 910
rect -638 850 -578 910
rect -438 850 -378 910
rect -238 850 -178 910
rect -38 850 22 910
rect 162 850 222 910
rect 362 850 422 910
rect 562 850 622 910
rect 762 850 822 910
rect 962 850 1022 910
rect 1162 850 1222 910
rect 1362 850 1422 910
rect 1562 850 1622 910
rect 1762 850 1822 910
rect 1962 850 2022 910
rect 2162 850 2222 910
rect 2362 850 2422 910
rect -2438 -1030 -2378 -970
rect -2238 -1030 -2178 -970
rect -2038 -1030 -1978 -970
rect -1838 -1030 -1778 -970
rect -1638 -1030 -1578 -970
rect -1438 -1030 -1378 -970
rect -1238 -1030 -1178 -970
rect -1038 -1030 -978 -970
rect -838 -1030 -778 -970
rect -638 -1030 -578 -970
rect -438 -1030 -378 -970
rect -238 -1030 -178 -970
rect -38 -1030 22 -970
rect 162 -1030 222 -970
rect 362 -1030 422 -970
rect 562 -1030 622 -970
rect 762 -1030 822 -970
rect 962 -1030 1022 -970
rect 1162 -1030 1222 -970
rect 1362 -1030 1422 -970
rect 1562 -1030 1622 -970
rect 1762 -1030 1822 -970
rect 1962 -1030 2022 -970
rect 2162 -1030 2222 -970
rect 2362 -1030 2422 -970
<< metal1 >>
rect -2706 910 2608 940
rect -2706 850 -2438 910
rect -2378 850 -2238 910
rect -2178 850 -2038 910
rect -1978 850 -1838 910
rect -1778 850 -1638 910
rect -1578 850 -1438 910
rect -1378 850 -1238 910
rect -1178 850 -1038 910
rect -978 850 -838 910
rect -778 850 -638 910
rect -578 850 -438 910
rect -378 850 -238 910
rect -178 850 -38 910
rect 22 850 162 910
rect 222 850 362 910
rect 422 850 562 910
rect 622 850 762 910
rect 822 850 962 910
rect 1022 850 1162 910
rect 1222 850 1362 910
rect 1422 850 1562 910
rect 1622 850 1762 910
rect 1822 850 1962 910
rect 2022 850 2162 910
rect 2222 850 2362 910
rect 2422 850 2608 910
rect -2706 820 2608 850
rect -2706 -970 2608 -940
rect -2706 -1030 -2438 -970
rect -2378 -1030 -2238 -970
rect -2178 -1030 -2038 -970
rect -1978 -1030 -1838 -970
rect -1778 -1030 -1638 -970
rect -1578 -1030 -1438 -970
rect -1378 -1030 -1238 -970
rect -1178 -1030 -1038 -970
rect -978 -1030 -838 -970
rect -778 -1030 -638 -970
rect -578 -1030 -438 -970
rect -378 -1030 -238 -970
rect -178 -1030 -38 -970
rect 22 -1030 162 -970
rect 222 -1030 362 -970
rect 422 -1030 562 -970
rect 622 -1030 762 -970
rect 822 -1030 962 -970
rect 1022 -1030 1162 -970
rect 1222 -1030 1362 -970
rect 1422 -1030 1562 -970
rect 1622 -1030 1762 -970
rect 1822 -1030 1962 -970
rect 2022 -1030 2162 -970
rect 2222 -1030 2362 -970
rect 2422 -1030 2608 -970
rect -2706 -1060 2608 -1030
use sky130_fd_pr__nfet_01v8_lvt_W76TCA  xm0
timestamp 0
transform 1 0 0 0 1 0
box 0 0 1 1
<< labels >>
flabel metal1 -2608 850 -2548 910 1 FreeSans 800 0 0 0 VPWR
flabel metal1 -2608 -1030 -2548 -970 1 FreeSans 800 0 0 0 VGND
flabel locali 2548 690 2608 750 1 FreeSans 800 0 0 0 SOURCE
flabel locali 2548 -530 2608 -470 1 FreeSans 800 0 0 0 DRAIN
flabel locali 2548 -796 2608 -736 1 FreeSans 800 0 0 0 GATE
<< end >>
