magic
tech sky130A
magscale 1 2
timestamp 1652936931
<< nwell >>
rect 90 294 4440 1940
rect 188 293 4440 294
<< pmoslvt >>
rect 282 355 682 1645
rect 740 355 1140 1645
rect 1198 355 1598 1645
rect 1656 355 2056 1645
rect 2114 355 2514 1645
rect 2572 355 2972 1645
rect 3030 355 3430 1645
rect 3488 355 3888 1645
rect 3946 355 4346 1645
<< pdiff >>
rect 224 1633 282 1645
rect 224 367 236 1633
rect 270 367 282 1633
rect 224 355 282 367
rect 682 1633 740 1645
rect 682 367 694 1633
rect 728 367 740 1633
rect 682 355 740 367
rect 1140 1633 1198 1645
rect 1140 367 1152 1633
rect 1186 367 1198 1633
rect 1140 355 1198 367
rect 1598 1633 1656 1645
rect 1598 367 1610 1633
rect 1644 367 1656 1633
rect 1598 355 1656 367
rect 2056 1633 2114 1645
rect 2056 367 2068 1633
rect 2102 367 2114 1633
rect 2056 355 2114 367
rect 2514 1633 2572 1645
rect 2514 367 2526 1633
rect 2560 367 2572 1633
rect 2514 355 2572 367
rect 2972 1633 3030 1645
rect 2972 367 2984 1633
rect 3018 367 3030 1633
rect 2972 355 3030 367
rect 3430 1633 3488 1645
rect 3430 367 3442 1633
rect 3476 367 3488 1633
rect 3430 355 3488 367
rect 3888 1633 3946 1645
rect 3888 367 3900 1633
rect 3934 367 3946 1633
rect 3888 355 3946 367
rect 4346 1633 4404 1645
rect 4346 367 4358 1633
rect 4392 367 4404 1633
rect 4346 355 4404 367
<< pdiffc >>
rect 236 367 270 1633
rect 694 367 728 1633
rect 1152 367 1186 1633
rect 1610 367 1644 1633
rect 2068 367 2102 1633
rect 2526 367 2560 1633
rect 2984 367 3018 1633
rect 3442 367 3476 1633
rect 3900 367 3934 1633
rect 4358 367 4392 1633
<< nsubdiff >>
rect 1188 1808 1308 1810
rect 128 1760 168 1800
rect 1188 1772 1228 1808
rect 1272 1772 1308 1808
rect 1188 1770 1308 1772
rect 2488 1808 2608 1810
rect 2488 1772 2528 1808
rect 2572 1772 2608 1808
rect 2488 1770 2608 1772
rect 128 1680 168 1720
<< nsubdiffcont >>
rect 1228 1772 1272 1808
rect 2528 1772 2572 1808
rect 128 1720 168 1760
<< poly >>
rect 282 1645 682 1671
rect 740 1645 1140 1671
rect 1198 1645 1598 1671
rect 1656 1645 2056 1671
rect 2114 1645 2514 1671
rect 2572 1645 2972 1671
rect 3030 1645 3430 1671
rect 3488 1645 3888 1671
rect 3946 1645 4346 1671
rect 282 329 682 355
rect 740 329 1140 355
rect 1198 329 1598 355
rect 1656 329 2056 355
rect 2114 329 2514 355
rect 2572 329 2972 355
rect 3030 329 3430 355
rect 3488 329 3888 355
rect 3946 329 4346 355
rect 428 184 548 329
rect 884 184 1004 329
rect 1340 184 1460 329
rect 1796 184 1916 329
rect 2252 184 2372 329
rect 2708 184 2828 329
rect 3164 184 3284 329
rect 3620 184 3740 329
rect 4076 184 4196 329
rect 188 164 4440 184
rect 188 104 358 164
rect 418 104 758 164
rect 818 104 1158 164
rect 1218 104 1558 164
rect 1618 104 1958 164
rect 2018 104 2358 164
rect 2418 104 2758 164
rect 2818 104 3158 164
rect 3218 104 3558 164
rect 3618 104 3958 164
rect 4018 104 4440 164
rect 188 84 4440 104
<< polycont >>
rect 358 104 418 164
rect 758 104 818 164
rect 1158 104 1218 164
rect 1558 104 1618 164
rect 1958 104 2018 164
rect 2358 104 2418 164
rect 2758 104 2818 164
rect 3158 104 3218 164
rect 3558 104 3618 164
rect 3958 104 4018 164
<< locali >>
rect 90 1850 358 1910
rect 418 1850 758 1910
rect 818 1850 1158 1910
rect 1218 1850 1558 1910
rect 1618 1850 1958 1910
rect 2018 1850 2358 1910
rect 2418 1850 2758 1910
rect 2818 1850 3158 1910
rect 3218 1850 3558 1910
rect 3618 1850 3958 1910
rect 4018 1850 4440 1910
rect 118 1760 178 1850
rect 1168 1808 1328 1850
rect 1168 1772 1228 1808
rect 1272 1772 1328 1808
rect 1168 1770 1328 1772
rect 2468 1808 2628 1850
rect 2468 1772 2528 1808
rect 2572 1772 2628 1808
rect 2468 1770 2628 1772
rect 118 1720 128 1760
rect 168 1720 178 1760
rect 118 1640 178 1720
rect 248 1690 4440 1730
rect 693 1649 727 1690
rect 1609 1649 1643 1690
rect 2525 1649 2559 1690
rect 3441 1649 3475 1690
rect 4357 1649 4391 1690
rect 236 1633 270 1649
rect 235 367 236 374
rect 693 1633 728 1649
rect 693 1626 694 1633
rect 235 351 270 367
rect 1152 1633 1186 1649
rect 694 351 728 367
rect 1151 367 1152 374
rect 1609 1633 1644 1649
rect 1609 1626 1610 1633
rect 1151 351 1186 367
rect 2068 1633 2102 1649
rect 1610 351 1644 367
rect 2067 367 2068 374
rect 2525 1633 2560 1649
rect 2525 1626 2526 1633
rect 2067 351 2102 367
rect 2984 1633 3018 1649
rect 2526 351 2560 367
rect 2983 367 2984 374
rect 3441 1633 3476 1649
rect 3441 1626 3442 1633
rect 2983 351 3018 367
rect 3900 1633 3934 1649
rect 3442 351 3476 367
rect 3899 367 3900 374
rect 4357 1633 4392 1649
rect 4357 1626 4358 1633
rect 3899 351 3934 367
rect 4358 351 4392 367
rect 235 270 269 351
rect 1151 270 1185 351
rect 2067 270 2101 351
rect 2983 270 3017 351
rect 3899 270 3933 351
rect 188 210 4440 270
rect 188 104 358 164
rect 418 104 758 164
rect 818 104 1158 164
rect 1218 104 1558 164
rect 1618 104 1958 164
rect 2018 104 2358 164
rect 2418 104 2758 164
rect 2818 104 3158 164
rect 3218 104 3558 164
rect 3618 104 3958 164
rect 4018 104 4440 164
rect 90 -30 358 30
rect 418 -30 758 30
rect 818 -30 1158 30
rect 1218 -30 1558 30
rect 1618 -30 1958 30
rect 2018 -30 2358 30
rect 2418 -30 2758 30
rect 2818 -30 3158 30
rect 3218 -30 3558 30
rect 3618 -30 3958 30
rect 4018 -30 4440 30
<< viali >>
rect 358 1850 418 1910
rect 758 1850 818 1910
rect 1158 1850 1218 1910
rect 1558 1850 1618 1910
rect 1958 1850 2018 1910
rect 2358 1850 2418 1910
rect 2758 1850 2818 1910
rect 3158 1850 3218 1910
rect 3558 1850 3618 1910
rect 3958 1850 4018 1910
rect 236 367 270 1633
rect 694 367 728 1633
rect 1152 367 1186 1633
rect 1610 367 1644 1633
rect 2068 367 2102 1633
rect 2526 367 2560 1633
rect 2984 367 3018 1633
rect 3442 367 3476 1633
rect 3900 367 3934 1633
rect 4358 367 4392 1633
rect 358 -30 418 30
rect 758 -30 818 30
rect 1158 -30 1218 30
rect 1558 -30 1618 30
rect 1958 -30 2018 30
rect 2358 -30 2418 30
rect 2758 -30 2818 30
rect 3158 -30 3218 30
rect 3558 -30 3618 30
rect 3958 -30 4018 30
<< metal1 >>
rect 90 1910 4440 1940
rect 90 1850 358 1910
rect 418 1850 758 1910
rect 818 1850 1158 1910
rect 1218 1850 1558 1910
rect 1618 1850 1958 1910
rect 2018 1850 2358 1910
rect 2418 1850 2758 1910
rect 2818 1850 3158 1910
rect 3218 1850 3558 1910
rect 3618 1850 3958 1910
rect 4018 1850 4440 1910
rect 90 1820 4440 1850
rect 230 1633 276 1645
rect 230 367 236 1633
rect 270 367 276 1633
rect 230 355 276 367
rect 688 1633 734 1645
rect 688 367 694 1633
rect 728 367 734 1633
rect 688 355 734 367
rect 1146 1633 1192 1645
rect 1146 367 1152 1633
rect 1186 367 1192 1633
rect 1146 355 1192 367
rect 1604 1633 1650 1645
rect 1604 367 1610 1633
rect 1644 367 1650 1633
rect 1604 355 1650 367
rect 2062 1633 2108 1645
rect 2062 367 2068 1633
rect 2102 367 2108 1633
rect 2062 355 2108 367
rect 2520 1633 2566 1645
rect 2520 367 2526 1633
rect 2560 367 2566 1633
rect 2520 355 2566 367
rect 2978 1633 3024 1645
rect 2978 367 2984 1633
rect 3018 367 3024 1633
rect 2978 355 3024 367
rect 3436 1633 3482 1645
rect 3436 367 3442 1633
rect 3476 367 3482 1633
rect 3436 355 3482 367
rect 3894 1633 3940 1645
rect 3894 367 3900 1633
rect 3934 367 3940 1633
rect 3894 355 3940 367
rect 4352 1633 4398 1645
rect 4352 367 4358 1633
rect 4392 367 4398 1633
rect 4352 355 4398 367
rect 90 30 4440 60
rect 90 -30 358 30
rect 418 -30 758 30
rect 818 -30 1158 30
rect 1218 -30 1558 30
rect 1618 -30 1958 30
rect 2018 -30 2358 30
rect 2418 -30 2758 30
rect 2818 -30 3158 30
rect 3218 -30 3558 30
rect 3618 -30 3958 30
rect 4018 -30 4440 30
rect 90 -60 4440 -30
<< labels >>
flabel nwell 90 1850 150 1910 1 FreeSans 800 0 0 0 VPWR
port 4 n power bidirectional
flabel metal1 90 -30 248 30 1 FreeSans 800 0 0 0 VGND
port 5 n ground bidirectional
flabel locali 4380 1690 4440 1730 1 FreeSans 800 0 0 0 SOURCE
port 2 n signal bidirectional
flabel locali 4380 210 4440 270 1 FreeSans 800 0 0 0 DRAIN
port 3 n signal bidirectional
flabel locali 4380 104 4440 164 1 FreeSans 800 0 0 0 GATE
port 1 n signal bidirectional
<< properties >>
string FIXED_BBOX 0 0 4530 1880
string LEFclass CORE
string LEFsite unitasc
<< end >>
