magic
tech sky130A
magscale 1 2
timestamp 1652142384
<< nwell >>
rect 0 1707 5722 1940
rect 0 294 5723 1707
rect 97 293 5723 294
<< pmoslvt >>
rect 191 355 591 1645
rect 649 355 1049 1645
rect 1107 355 1507 1645
rect 1565 355 1965 1645
rect 2023 355 2423 1645
rect 2481 355 2881 1645
rect 2939 355 3339 1645
rect 3397 355 3797 1645
rect 3855 355 4255 1645
rect 4313 355 4713 1645
rect 4771 355 5171 1645
rect 5229 355 5629 1645
<< pdiff >>
rect 133 1633 191 1645
rect 133 367 145 1633
rect 179 367 191 1633
rect 133 355 191 367
rect 591 1633 649 1645
rect 591 367 603 1633
rect 637 367 649 1633
rect 591 355 649 367
rect 1049 1633 1107 1645
rect 1049 367 1061 1633
rect 1095 367 1107 1633
rect 1049 355 1107 367
rect 1507 1633 1565 1645
rect 1507 367 1519 1633
rect 1553 367 1565 1633
rect 1507 355 1565 367
rect 1965 1633 2023 1645
rect 1965 367 1977 1633
rect 2011 367 2023 1633
rect 1965 355 2023 367
rect 2423 1633 2481 1645
rect 2423 367 2435 1633
rect 2469 367 2481 1633
rect 2423 355 2481 367
rect 2881 1633 2939 1645
rect 2881 367 2893 1633
rect 2927 367 2939 1633
rect 2881 355 2939 367
rect 3339 1633 3397 1645
rect 3339 367 3351 1633
rect 3385 367 3397 1633
rect 3339 355 3397 367
rect 3797 1633 3855 1645
rect 3797 367 3809 1633
rect 3843 367 3855 1633
rect 3797 355 3855 367
rect 4255 1633 4313 1645
rect 4255 367 4267 1633
rect 4301 367 4313 1633
rect 4255 355 4313 367
rect 4713 1633 4771 1645
rect 4713 367 4725 1633
rect 4759 367 4771 1633
rect 4713 355 4771 367
rect 5171 1633 5229 1645
rect 5171 367 5183 1633
rect 5217 367 5229 1633
rect 5171 355 5229 367
rect 5629 1633 5687 1645
rect 5629 367 5641 1633
rect 5675 367 5687 1633
rect 5629 355 5687 367
<< pdiffc >>
rect 145 367 179 1633
rect 603 367 637 1633
rect 1061 367 1095 1633
rect 1519 367 1553 1633
rect 1977 367 2011 1633
rect 2435 367 2469 1633
rect 2893 367 2927 1633
rect 3351 367 3385 1633
rect 3809 367 3843 1633
rect 4267 367 4301 1633
rect 4725 367 4759 1633
rect 5183 367 5217 1633
rect 5641 367 5675 1633
<< nsubdiff >>
rect 38 1760 78 1800
rect 38 1680 78 1720
<< nsubdiffcont >>
rect 38 1720 78 1760
<< poly >>
rect 191 1645 591 1671
rect 649 1645 1049 1671
rect 1107 1645 1507 1671
rect 1565 1645 1965 1671
rect 2023 1645 2423 1671
rect 2481 1645 2881 1671
rect 2939 1645 3339 1671
rect 3397 1645 3797 1671
rect 3855 1645 4255 1671
rect 4313 1645 4713 1671
rect 4771 1645 5171 1671
rect 5229 1645 5629 1671
rect 191 329 591 355
rect 649 329 1049 355
rect 1107 329 1507 355
rect 1565 329 1965 355
rect 2023 329 2423 355
rect 2481 329 2881 355
rect 2939 329 3339 355
rect 3397 329 3797 355
rect 3855 329 4255 355
rect 4313 329 4713 355
rect 4771 329 5171 355
rect 5229 329 5629 355
rect 338 184 458 329
rect 794 184 914 329
rect 1250 184 1370 329
rect 1706 184 1826 329
rect 2162 184 2282 329
rect 2618 184 2738 329
rect 3074 184 3194 329
rect 3530 184 3650 329
rect 3986 184 4106 329
rect 4442 184 4562 329
rect 4898 184 5018 329
rect 5354 184 5474 329
rect 98 164 5722 184
rect 98 104 268 164
rect 328 104 668 164
rect 728 104 1068 164
rect 1128 104 1468 164
rect 1528 104 1868 164
rect 1928 104 2268 164
rect 2328 104 2668 164
rect 2728 104 3068 164
rect 3128 104 3468 164
rect 3528 104 3868 164
rect 3928 104 4268 164
rect 4328 104 4668 164
rect 4728 104 5068 164
rect 5128 104 5468 164
rect 5528 104 5722 164
rect 98 84 5722 104
<< polycont >>
rect 268 104 328 164
rect 668 104 728 164
rect 1068 104 1128 164
rect 1468 104 1528 164
rect 1868 104 1928 164
rect 2268 104 2328 164
rect 2668 104 2728 164
rect 3068 104 3128 164
rect 3468 104 3528 164
rect 3868 104 3928 164
rect 4268 104 4328 164
rect 4668 104 4728 164
rect 5068 104 5128 164
rect 5468 104 5528 164
<< locali >>
rect 0 1850 268 1910
rect 328 1850 668 1910
rect 728 1850 1068 1910
rect 1128 1850 1468 1910
rect 1528 1850 1868 1910
rect 1928 1850 2268 1910
rect 2328 1850 2668 1910
rect 2728 1850 3068 1910
rect 3128 1850 3468 1910
rect 3528 1850 3868 1910
rect 3928 1850 4268 1910
rect 4328 1850 4668 1910
rect 4728 1850 5068 1910
rect 5128 1850 5468 1910
rect 5528 1850 5722 1910
rect 28 1760 88 1850
rect 28 1720 38 1760
rect 78 1720 88 1760
rect 158 1730 5722 1790
rect 28 1640 88 1720
rect 145 1633 179 1649
rect 145 270 179 367
rect 603 1633 637 1730
rect 603 351 637 367
rect 1061 1633 1095 1649
rect 1061 270 1095 367
rect 1519 1633 1553 1730
rect 1519 351 1553 367
rect 1977 1633 2011 1649
rect 1977 270 2011 367
rect 2435 1633 2469 1730
rect 2435 351 2469 367
rect 2893 1633 2927 1649
rect 2893 270 2927 367
rect 3351 1633 3385 1730
rect 3351 351 3385 367
rect 3809 1633 3843 1649
rect 3809 270 3843 367
rect 4267 1633 4301 1730
rect 4267 351 4301 367
rect 4725 1633 4759 1649
rect 4725 270 4759 367
rect 5183 1633 5217 1730
rect 5183 351 5217 367
rect 5641 1633 5675 1649
rect 5641 270 5675 367
rect 98 210 5722 270
rect 98 104 268 164
rect 328 104 668 164
rect 728 104 1068 164
rect 1128 104 1468 164
rect 1528 104 1868 164
rect 1928 104 2268 164
rect 2328 104 2668 164
rect 2728 104 3068 164
rect 3128 104 3468 164
rect 3528 104 3868 164
rect 3928 104 4268 164
rect 4328 104 4668 164
rect 4728 104 5068 164
rect 5128 104 5468 164
rect 5528 104 5722 164
rect 0 -30 268 30
rect 328 -30 668 30
rect 728 -30 1068 30
rect 1128 -30 1468 30
rect 1528 -30 1868 30
rect 1928 -30 2268 30
rect 2328 -30 2668 30
rect 2728 -30 3068 30
rect 3128 -30 3468 30
rect 3528 -30 3868 30
rect 3928 -30 4268 30
rect 4328 -30 4668 30
rect 4728 -30 5068 30
rect 5128 -30 5468 30
rect 5528 -30 5722 30
<< viali >>
rect 268 1850 328 1910
rect 668 1850 728 1910
rect 1068 1850 1128 1910
rect 1468 1850 1528 1910
rect 1868 1850 1928 1910
rect 2268 1850 2328 1910
rect 2668 1850 2728 1910
rect 3068 1850 3128 1910
rect 3468 1850 3528 1910
rect 3868 1850 3928 1910
rect 4268 1850 4328 1910
rect 4668 1850 4728 1910
rect 5068 1850 5128 1910
rect 5468 1850 5528 1910
rect 145 367 179 1633
rect 603 367 637 1633
rect 1061 367 1095 1633
rect 1519 367 1553 1633
rect 1977 367 2011 1633
rect 2435 367 2469 1633
rect 2893 367 2927 1633
rect 3351 367 3385 1633
rect 3809 367 3843 1633
rect 4267 367 4301 1633
rect 4725 367 4759 1633
rect 5183 367 5217 1633
rect 5641 367 5675 1633
rect 268 -30 328 30
rect 668 -30 728 30
rect 1068 -30 1128 30
rect 1468 -30 1528 30
rect 1868 -30 1928 30
rect 2268 -30 2328 30
rect 2668 -30 2728 30
rect 3068 -30 3128 30
rect 3468 -30 3528 30
rect 3868 -30 3928 30
rect 4268 -30 4328 30
rect 4668 -30 4728 30
rect 5068 -30 5128 30
rect 5468 -30 5528 30
<< metal1 >>
rect 0 1910 5722 1940
rect 0 1850 268 1910
rect 328 1850 668 1910
rect 728 1850 1068 1910
rect 1128 1850 1468 1910
rect 1528 1850 1868 1910
rect 1928 1850 2268 1910
rect 2328 1850 2668 1910
rect 2728 1850 3068 1910
rect 3128 1850 3468 1910
rect 3528 1850 3868 1910
rect 3928 1850 4268 1910
rect 4328 1850 4668 1910
rect 4728 1850 5068 1910
rect 5128 1850 5468 1910
rect 5528 1850 5722 1910
rect 0 1820 5722 1850
rect 139 1633 185 1645
rect 139 367 145 1633
rect 179 367 185 1633
rect 139 355 185 367
rect 597 1633 643 1645
rect 597 367 603 1633
rect 637 367 643 1633
rect 597 355 643 367
rect 1055 1633 1101 1645
rect 1055 367 1061 1633
rect 1095 367 1101 1633
rect 1055 355 1101 367
rect 1513 1633 1559 1645
rect 1513 367 1519 1633
rect 1553 367 1559 1633
rect 1513 355 1559 367
rect 1971 1633 2017 1645
rect 1971 367 1977 1633
rect 2011 367 2017 1633
rect 1971 355 2017 367
rect 2429 1633 2475 1645
rect 2429 367 2435 1633
rect 2469 367 2475 1633
rect 2429 355 2475 367
rect 2887 1633 2933 1645
rect 2887 367 2893 1633
rect 2927 367 2933 1633
rect 2887 355 2933 367
rect 3345 1633 3391 1645
rect 3345 367 3351 1633
rect 3385 367 3391 1633
rect 3345 355 3391 367
rect 3803 1633 3849 1645
rect 3803 367 3809 1633
rect 3843 367 3849 1633
rect 3803 355 3849 367
rect 4261 1633 4307 1645
rect 4261 367 4267 1633
rect 4301 367 4307 1633
rect 4261 355 4307 367
rect 4719 1633 4765 1645
rect 4719 367 4725 1633
rect 4759 367 4765 1633
rect 4719 355 4765 367
rect 5177 1633 5223 1645
rect 5177 367 5183 1633
rect 5217 367 5223 1633
rect 5177 355 5223 367
rect 5635 1633 5681 1645
rect 5635 367 5641 1633
rect 5675 367 5681 1633
rect 5635 355 5681 367
rect 0 30 5722 60
rect 0 -30 268 30
rect 328 -30 668 30
rect 728 -30 1068 30
rect 1128 -30 1468 30
rect 1528 -30 1868 30
rect 1928 -30 2268 30
rect 2328 -30 2668 30
rect 2728 -30 3068 30
rect 3128 -30 3468 30
rect 3528 -30 3868 30
rect 3928 -30 4268 30
rect 4328 -30 4668 30
rect 4728 -30 5068 30
rect 5128 -30 5468 30
rect 5528 -30 5722 30
rect 0 -60 5722 -30
<< labels >>
flabel nwell 0 1850 60 1910 1 FreeSans 800 0 0 0 VPWR
port 4 n power bidirectional
flabel metal1 0 -30 158 30 1 FreeSans 800 0 0 0 VGND
port 5 n ground bidirectional
flabel locali 5662 1730 5722 1790 1 FreeSans 800 0 0 0 SOURCE
port 2 n signal bidirectional
flabel locali 5662 210 5722 270 1 FreeSans 800 0 0 0 DRAIN
port 3 n signal bidirectional
flabel locali 5662 104 5722 164 1 FreeSans 800 0 0 0 GATE
port 1 n signal bidirectional
<< properties >>
string FIXED_BBOX 0 0 5723 1880
string LEFclass CORE
string LEFsite unitasc
<< end >>
