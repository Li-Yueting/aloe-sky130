VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO sky130_asc_pfet_01v8_lvt_60
  CLASS CORE ;
  FOREIGN sky130_asc_pfet_01v8_lvt_60 ;
  ORIGIN 0.000 0.000 ;
  SIZE 139.435 BY 9.400 ;
  SITE unitasc ;
  PIN GATE
    DIRECTION INOUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 774.000000 ;
    PORT
      LAYER li1 ;
        RECT 0.940 0.520 138.980 0.820 ;
    END
  END GATE
  PIN SOURCE
    DIRECTION INOUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 56.114998 ;
    PORT
      LAYER li1 ;
        RECT 1.240 8.650 138.980 8.950 ;
        RECT 3.465 1.755 3.635 8.650 ;
        RECT 8.045 1.755 8.215 8.650 ;
        RECT 12.625 1.755 12.795 8.650 ;
        RECT 17.205 1.755 17.375 8.650 ;
        RECT 21.785 1.755 21.955 8.650 ;
        RECT 26.365 1.755 26.535 8.650 ;
        RECT 30.945 1.755 31.115 8.650 ;
        RECT 35.525 1.755 35.695 8.650 ;
        RECT 40.105 1.755 40.275 8.650 ;
        RECT 44.685 1.755 44.855 8.650 ;
        RECT 49.265 1.755 49.435 8.650 ;
        RECT 53.845 1.755 54.015 8.650 ;
        RECT 58.425 1.755 58.595 8.650 ;
        RECT 63.005 1.755 63.175 8.650 ;
        RECT 67.585 1.755 67.755 8.650 ;
        RECT 72.165 1.755 72.335 8.650 ;
        RECT 76.745 1.755 76.915 8.650 ;
        RECT 81.325 1.755 81.495 8.650 ;
        RECT 85.905 1.755 86.075 8.650 ;
        RECT 90.485 1.755 90.655 8.650 ;
        RECT 95.065 1.755 95.235 8.650 ;
        RECT 99.645 1.755 99.815 8.650 ;
        RECT 104.225 1.755 104.395 8.650 ;
        RECT 108.805 1.755 108.975 8.650 ;
        RECT 113.385 1.755 113.555 8.650 ;
        RECT 117.965 1.755 118.135 8.650 ;
        RECT 122.545 1.755 122.715 8.650 ;
        RECT 127.125 1.755 127.295 8.650 ;
        RECT 131.705 1.755 131.875 8.650 ;
        RECT 136.285 1.755 136.455 8.650 ;
      LAYER mcon ;
        RECT 3.465 1.835 3.635 8.165 ;
        RECT 8.045 1.835 8.215 8.165 ;
        RECT 12.625 1.835 12.795 8.165 ;
        RECT 17.205 1.835 17.375 8.165 ;
        RECT 21.785 1.835 21.955 8.165 ;
        RECT 26.365 1.835 26.535 8.165 ;
        RECT 30.945 1.835 31.115 8.165 ;
        RECT 35.525 1.835 35.695 8.165 ;
        RECT 40.105 1.835 40.275 8.165 ;
        RECT 44.685 1.835 44.855 8.165 ;
        RECT 49.265 1.835 49.435 8.165 ;
        RECT 53.845 1.835 54.015 8.165 ;
        RECT 58.425 1.835 58.595 8.165 ;
        RECT 63.005 1.835 63.175 8.165 ;
        RECT 67.585 1.835 67.755 8.165 ;
        RECT 72.165 1.835 72.335 8.165 ;
        RECT 76.745 1.835 76.915 8.165 ;
        RECT 81.325 1.835 81.495 8.165 ;
        RECT 85.905 1.835 86.075 8.165 ;
        RECT 90.485 1.835 90.655 8.165 ;
        RECT 95.065 1.835 95.235 8.165 ;
        RECT 99.645 1.835 99.815 8.165 ;
        RECT 104.225 1.835 104.395 8.165 ;
        RECT 108.805 1.835 108.975 8.165 ;
        RECT 113.385 1.835 113.555 8.165 ;
        RECT 117.965 1.835 118.135 8.165 ;
        RECT 122.545 1.835 122.715 8.165 ;
        RECT 127.125 1.835 127.295 8.165 ;
        RECT 131.705 1.835 131.875 8.165 ;
        RECT 136.285 1.835 136.455 8.165 ;
      LAYER met1 ;
        RECT 3.435 1.775 3.665 8.225 ;
        RECT 8.015 1.775 8.245 8.225 ;
        RECT 12.595 1.775 12.825 8.225 ;
        RECT 17.175 1.775 17.405 8.225 ;
        RECT 21.755 1.775 21.985 8.225 ;
        RECT 26.335 1.775 26.565 8.225 ;
        RECT 30.915 1.775 31.145 8.225 ;
        RECT 35.495 1.775 35.725 8.225 ;
        RECT 40.075 1.775 40.305 8.225 ;
        RECT 44.655 1.775 44.885 8.225 ;
        RECT 49.235 1.775 49.465 8.225 ;
        RECT 53.815 1.775 54.045 8.225 ;
        RECT 58.395 1.775 58.625 8.225 ;
        RECT 62.975 1.775 63.205 8.225 ;
        RECT 67.555 1.775 67.785 8.225 ;
        RECT 72.135 1.775 72.365 8.225 ;
        RECT 76.715 1.775 76.945 8.225 ;
        RECT 81.295 1.775 81.525 8.225 ;
        RECT 85.875 1.775 86.105 8.225 ;
        RECT 90.455 1.775 90.685 8.225 ;
        RECT 95.035 1.775 95.265 8.225 ;
        RECT 99.615 1.775 99.845 8.225 ;
        RECT 104.195 1.775 104.425 8.225 ;
        RECT 108.775 1.775 109.005 8.225 ;
        RECT 113.355 1.775 113.585 8.225 ;
        RECT 117.935 1.775 118.165 8.225 ;
        RECT 122.515 1.775 122.745 8.225 ;
        RECT 127.095 1.775 127.325 8.225 ;
        RECT 131.675 1.775 131.905 8.225 ;
        RECT 136.255 1.775 136.485 8.225 ;
    END
  END SOURCE
  PIN DRAIN
    DIRECTION INOUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 57.985500 ;
    PORT
      LAYER li1 ;
        RECT 1.175 1.350 1.345 8.245 ;
        RECT 5.755 1.350 5.925 8.245 ;
        RECT 10.335 1.350 10.505 8.245 ;
        RECT 14.915 1.350 15.085 8.245 ;
        RECT 19.495 1.350 19.665 8.245 ;
        RECT 24.075 1.350 24.245 8.245 ;
        RECT 28.655 1.350 28.825 8.245 ;
        RECT 33.235 1.350 33.405 8.245 ;
        RECT 37.815 1.350 37.985 8.245 ;
        RECT 42.395 1.350 42.565 8.245 ;
        RECT 46.975 1.350 47.145 8.245 ;
        RECT 51.555 1.350 51.725 8.245 ;
        RECT 56.135 1.350 56.305 8.245 ;
        RECT 60.715 1.350 60.885 8.245 ;
        RECT 65.295 1.350 65.465 8.245 ;
        RECT 69.875 1.350 70.045 8.245 ;
        RECT 74.455 1.350 74.625 8.245 ;
        RECT 79.035 1.350 79.205 8.245 ;
        RECT 83.615 1.350 83.785 8.245 ;
        RECT 88.195 1.350 88.365 8.245 ;
        RECT 92.775 1.350 92.945 8.245 ;
        RECT 97.355 1.350 97.525 8.245 ;
        RECT 101.935 1.350 102.105 8.245 ;
        RECT 106.515 1.350 106.685 8.245 ;
        RECT 111.095 1.350 111.265 8.245 ;
        RECT 115.675 1.350 115.845 8.245 ;
        RECT 120.255 1.350 120.425 8.245 ;
        RECT 124.835 1.350 125.005 8.245 ;
        RECT 129.415 1.350 129.585 8.245 ;
        RECT 133.995 1.350 134.165 8.245 ;
        RECT 138.575 1.350 138.745 8.245 ;
        RECT 0.940 1.050 138.980 1.350 ;
      LAYER mcon ;
        RECT 1.175 1.835 1.345 8.165 ;
        RECT 5.755 1.835 5.925 8.165 ;
        RECT 10.335 1.835 10.505 8.165 ;
        RECT 14.915 1.835 15.085 8.165 ;
        RECT 19.495 1.835 19.665 8.165 ;
        RECT 24.075 1.835 24.245 8.165 ;
        RECT 28.655 1.835 28.825 8.165 ;
        RECT 33.235 1.835 33.405 8.165 ;
        RECT 37.815 1.835 37.985 8.165 ;
        RECT 42.395 1.835 42.565 8.165 ;
        RECT 46.975 1.835 47.145 8.165 ;
        RECT 51.555 1.835 51.725 8.165 ;
        RECT 56.135 1.835 56.305 8.165 ;
        RECT 60.715 1.835 60.885 8.165 ;
        RECT 65.295 1.835 65.465 8.165 ;
        RECT 69.875 1.835 70.045 8.165 ;
        RECT 74.455 1.835 74.625 8.165 ;
        RECT 79.035 1.835 79.205 8.165 ;
        RECT 83.615 1.835 83.785 8.165 ;
        RECT 88.195 1.835 88.365 8.165 ;
        RECT 92.775 1.835 92.945 8.165 ;
        RECT 97.355 1.835 97.525 8.165 ;
        RECT 101.935 1.835 102.105 8.165 ;
        RECT 106.515 1.835 106.685 8.165 ;
        RECT 111.095 1.835 111.265 8.165 ;
        RECT 115.675 1.835 115.845 8.165 ;
        RECT 120.255 1.835 120.425 8.165 ;
        RECT 124.835 1.835 125.005 8.165 ;
        RECT 129.415 1.835 129.585 8.165 ;
        RECT 133.995 1.835 134.165 8.165 ;
        RECT 138.575 1.835 138.745 8.165 ;
      LAYER met1 ;
        RECT 1.145 1.775 1.375 8.225 ;
        RECT 5.725 1.775 5.955 8.225 ;
        RECT 10.305 1.775 10.535 8.225 ;
        RECT 14.885 1.775 15.115 8.225 ;
        RECT 19.465 1.775 19.695 8.225 ;
        RECT 24.045 1.775 24.275 8.225 ;
        RECT 28.625 1.775 28.855 8.225 ;
        RECT 33.205 1.775 33.435 8.225 ;
        RECT 37.785 1.775 38.015 8.225 ;
        RECT 42.365 1.775 42.595 8.225 ;
        RECT 46.945 1.775 47.175 8.225 ;
        RECT 51.525 1.775 51.755 8.225 ;
        RECT 56.105 1.775 56.335 8.225 ;
        RECT 60.685 1.775 60.915 8.225 ;
        RECT 65.265 1.775 65.495 8.225 ;
        RECT 69.845 1.775 70.075 8.225 ;
        RECT 74.425 1.775 74.655 8.225 ;
        RECT 79.005 1.775 79.235 8.225 ;
        RECT 83.585 1.775 83.815 8.225 ;
        RECT 88.165 1.775 88.395 8.225 ;
        RECT 92.745 1.775 92.975 8.225 ;
        RECT 97.325 1.775 97.555 8.225 ;
        RECT 101.905 1.775 102.135 8.225 ;
        RECT 106.485 1.775 106.715 8.225 ;
        RECT 111.065 1.775 111.295 8.225 ;
        RECT 115.645 1.775 115.875 8.225 ;
        RECT 120.225 1.775 120.455 8.225 ;
        RECT 124.805 1.775 125.035 8.225 ;
        RECT 129.385 1.775 129.615 8.225 ;
        RECT 133.965 1.775 134.195 8.225 ;
        RECT 138.545 1.775 138.775 8.225 ;
    END
  END DRAIN
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT 0.450 8.535 138.980 9.700 ;
        RECT 0.450 1.470 138.985 8.535 ;
        RECT 0.935 1.465 138.985 1.470 ;
      LAYER li1 ;
        RECT 0.450 9.250 138.980 9.550 ;
        RECT 0.590 8.200 0.890 9.250 ;
      LAYER mcon ;
        RECT 1.790 9.250 2.090 9.550 ;
        RECT 3.790 9.250 4.090 9.550 ;
        RECT 5.790 9.250 6.090 9.550 ;
        RECT 7.790 9.250 8.090 9.550 ;
        RECT 9.790 9.250 10.090 9.550 ;
        RECT 11.790 9.250 12.090 9.550 ;
        RECT 13.790 9.250 14.090 9.550 ;
        RECT 15.790 9.250 16.090 9.550 ;
        RECT 17.790 9.250 18.090 9.550 ;
        RECT 19.790 9.250 20.090 9.550 ;
        RECT 21.790 9.250 22.090 9.550 ;
        RECT 23.790 9.250 24.090 9.550 ;
        RECT 25.790 9.250 26.090 9.550 ;
        RECT 27.790 9.250 28.090 9.550 ;
        RECT 29.790 9.250 30.090 9.550 ;
        RECT 31.790 9.250 32.090 9.550 ;
        RECT 33.790 9.250 34.090 9.550 ;
        RECT 35.790 9.250 36.090 9.550 ;
        RECT 37.790 9.250 38.090 9.550 ;
        RECT 39.790 9.250 40.090 9.550 ;
        RECT 41.790 9.250 42.090 9.550 ;
        RECT 43.790 9.250 44.090 9.550 ;
        RECT 45.790 9.250 46.090 9.550 ;
        RECT 47.790 9.250 48.090 9.550 ;
        RECT 49.790 9.250 50.090 9.550 ;
        RECT 51.790 9.250 52.090 9.550 ;
        RECT 53.790 9.250 54.090 9.550 ;
        RECT 55.790 9.250 56.090 9.550 ;
        RECT 57.790 9.250 58.090 9.550 ;
        RECT 59.790 9.250 60.090 9.550 ;
        RECT 61.790 9.250 62.090 9.550 ;
        RECT 63.790 9.250 64.090 9.550 ;
        RECT 65.790 9.250 66.090 9.550 ;
        RECT 67.790 9.250 68.090 9.550 ;
        RECT 69.790 9.250 70.090 9.550 ;
        RECT 71.790 9.250 72.090 9.550 ;
        RECT 73.790 9.250 74.090 9.550 ;
        RECT 75.790 9.250 76.090 9.550 ;
        RECT 77.790 9.250 78.090 9.550 ;
        RECT 79.790 9.250 80.090 9.550 ;
        RECT 81.790 9.250 82.090 9.550 ;
        RECT 83.790 9.250 84.090 9.550 ;
        RECT 85.790 9.250 86.090 9.550 ;
        RECT 87.790 9.250 88.090 9.550 ;
        RECT 89.790 9.250 90.090 9.550 ;
        RECT 91.790 9.250 92.090 9.550 ;
        RECT 93.790 9.250 94.090 9.550 ;
        RECT 95.790 9.250 96.090 9.550 ;
        RECT 97.790 9.250 98.090 9.550 ;
        RECT 99.790 9.250 100.090 9.550 ;
        RECT 101.790 9.250 102.090 9.550 ;
        RECT 103.790 9.250 104.090 9.550 ;
        RECT 105.790 9.250 106.090 9.550 ;
        RECT 107.790 9.250 108.090 9.550 ;
        RECT 109.790 9.250 110.090 9.550 ;
        RECT 111.790 9.250 112.090 9.550 ;
        RECT 113.790 9.250 114.090 9.550 ;
        RECT 115.790 9.250 116.090 9.550 ;
        RECT 117.790 9.250 118.090 9.550 ;
        RECT 119.790 9.250 120.090 9.550 ;
        RECT 121.790 9.250 122.090 9.550 ;
        RECT 123.790 9.250 124.090 9.550 ;
        RECT 125.790 9.250 126.090 9.550 ;
        RECT 127.790 9.250 128.090 9.550 ;
        RECT 129.790 9.250 130.090 9.550 ;
        RECT 131.790 9.250 132.090 9.550 ;
        RECT 133.790 9.250 134.090 9.550 ;
        RECT 135.790 9.250 136.090 9.550 ;
        RECT 137.790 9.250 138.090 9.550 ;
      LAYER met1 ;
        RECT 0.450 9.100 138.980 9.700 ;
    END
  END VPWR
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER li1 ;
        RECT 0.450 -0.150 138.980 0.150 ;
      LAYER mcon ;
        RECT 1.790 -0.150 2.090 0.150 ;
        RECT 3.790 -0.150 4.090 0.150 ;
        RECT 5.790 -0.150 6.090 0.150 ;
        RECT 7.790 -0.150 8.090 0.150 ;
        RECT 9.790 -0.150 10.090 0.150 ;
        RECT 11.790 -0.150 12.090 0.150 ;
        RECT 13.790 -0.150 14.090 0.150 ;
        RECT 15.790 -0.150 16.090 0.150 ;
        RECT 17.790 -0.150 18.090 0.150 ;
        RECT 19.790 -0.150 20.090 0.150 ;
        RECT 21.790 -0.150 22.090 0.150 ;
        RECT 23.790 -0.150 24.090 0.150 ;
        RECT 25.790 -0.150 26.090 0.150 ;
        RECT 27.790 -0.150 28.090 0.150 ;
        RECT 29.790 -0.150 30.090 0.150 ;
        RECT 31.790 -0.150 32.090 0.150 ;
        RECT 33.790 -0.150 34.090 0.150 ;
        RECT 35.790 -0.150 36.090 0.150 ;
        RECT 37.790 -0.150 38.090 0.150 ;
        RECT 39.790 -0.150 40.090 0.150 ;
        RECT 41.790 -0.150 42.090 0.150 ;
        RECT 43.790 -0.150 44.090 0.150 ;
        RECT 45.790 -0.150 46.090 0.150 ;
        RECT 47.790 -0.150 48.090 0.150 ;
        RECT 49.790 -0.150 50.090 0.150 ;
        RECT 51.790 -0.150 52.090 0.150 ;
        RECT 53.790 -0.150 54.090 0.150 ;
        RECT 55.790 -0.150 56.090 0.150 ;
        RECT 57.790 -0.150 58.090 0.150 ;
        RECT 59.790 -0.150 60.090 0.150 ;
        RECT 61.790 -0.150 62.090 0.150 ;
        RECT 63.790 -0.150 64.090 0.150 ;
        RECT 65.790 -0.150 66.090 0.150 ;
        RECT 67.790 -0.150 68.090 0.150 ;
        RECT 69.790 -0.150 70.090 0.150 ;
        RECT 71.790 -0.150 72.090 0.150 ;
        RECT 73.790 -0.150 74.090 0.150 ;
        RECT 75.790 -0.150 76.090 0.150 ;
        RECT 77.790 -0.150 78.090 0.150 ;
        RECT 79.790 -0.150 80.090 0.150 ;
        RECT 81.790 -0.150 82.090 0.150 ;
        RECT 83.790 -0.150 84.090 0.150 ;
        RECT 85.790 -0.150 86.090 0.150 ;
        RECT 87.790 -0.150 88.090 0.150 ;
        RECT 89.790 -0.150 90.090 0.150 ;
        RECT 91.790 -0.150 92.090 0.150 ;
        RECT 93.790 -0.150 94.090 0.150 ;
        RECT 95.790 -0.150 96.090 0.150 ;
        RECT 97.790 -0.150 98.090 0.150 ;
        RECT 99.790 -0.150 100.090 0.150 ;
        RECT 101.790 -0.150 102.090 0.150 ;
        RECT 103.790 -0.150 104.090 0.150 ;
        RECT 105.790 -0.150 106.090 0.150 ;
        RECT 107.790 -0.150 108.090 0.150 ;
        RECT 109.790 -0.150 110.090 0.150 ;
        RECT 111.790 -0.150 112.090 0.150 ;
        RECT 113.790 -0.150 114.090 0.150 ;
        RECT 115.790 -0.150 116.090 0.150 ;
        RECT 117.790 -0.150 118.090 0.150 ;
        RECT 119.790 -0.150 120.090 0.150 ;
        RECT 121.790 -0.150 122.090 0.150 ;
        RECT 123.790 -0.150 124.090 0.150 ;
        RECT 125.790 -0.150 126.090 0.150 ;
        RECT 127.790 -0.150 128.090 0.150 ;
        RECT 129.790 -0.150 130.090 0.150 ;
        RECT 131.790 -0.150 132.090 0.150 ;
        RECT 133.790 -0.150 134.090 0.150 ;
        RECT 135.790 -0.150 136.090 0.150 ;
        RECT 137.790 -0.150 138.090 0.150 ;
      LAYER met1 ;
        RECT 0.450 -0.300 138.980 0.300 ;
    END
  END VGND
END sky130_asc_pfet_01v8_lvt_60
END LIBRARY

