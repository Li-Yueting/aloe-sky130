magic
tech sky130A
magscale 1 2
timestamp 1653341788
<< nwell >>
rect 120 294 4470 1940
rect 218 293 4470 294
<< pmoslvt >>
rect 312 355 712 1645
rect 770 355 1170 1645
rect 1228 355 1628 1645
rect 1686 355 2086 1645
rect 2144 355 2544 1645
rect 2602 355 3002 1645
rect 3060 355 3460 1645
rect 3518 355 3918 1645
rect 3976 355 4376 1645
<< pdiff >>
rect 254 1633 312 1645
rect 254 367 266 1633
rect 300 367 312 1633
rect 254 355 312 367
rect 712 1633 770 1645
rect 712 367 724 1633
rect 758 367 770 1633
rect 712 355 770 367
rect 1170 1633 1228 1645
rect 1170 367 1182 1633
rect 1216 367 1228 1633
rect 1170 355 1228 367
rect 1628 1633 1686 1645
rect 1628 367 1640 1633
rect 1674 367 1686 1633
rect 1628 355 1686 367
rect 2086 1633 2144 1645
rect 2086 367 2098 1633
rect 2132 367 2144 1633
rect 2086 355 2144 367
rect 2544 1633 2602 1645
rect 2544 367 2556 1633
rect 2590 367 2602 1633
rect 2544 355 2602 367
rect 3002 1633 3060 1645
rect 3002 367 3014 1633
rect 3048 367 3060 1633
rect 3002 355 3060 367
rect 3460 1633 3518 1645
rect 3460 367 3472 1633
rect 3506 367 3518 1633
rect 3460 355 3518 367
rect 3918 1633 3976 1645
rect 3918 367 3930 1633
rect 3964 367 3976 1633
rect 3918 355 3976 367
rect 4376 1633 4434 1645
rect 4376 367 4388 1633
rect 4422 367 4434 1633
rect 4376 355 4434 367
<< pdiffc >>
rect 266 367 300 1633
rect 724 367 758 1633
rect 1182 367 1216 1633
rect 1640 367 1674 1633
rect 2098 367 2132 1633
rect 2556 367 2590 1633
rect 3014 367 3048 1633
rect 3472 367 3506 1633
rect 3930 367 3964 1633
rect 4388 367 4422 1633
<< nsubdiff >>
rect 1218 1808 1338 1810
rect 158 1760 198 1800
rect 1218 1772 1258 1808
rect 1302 1772 1338 1808
rect 1218 1770 1338 1772
rect 2518 1808 2638 1810
rect 2518 1772 2558 1808
rect 2602 1772 2638 1808
rect 2518 1770 2638 1772
rect 158 1680 198 1720
<< nsubdiffcont >>
rect 1258 1772 1302 1808
rect 2558 1772 2602 1808
rect 158 1720 198 1760
<< poly >>
rect 312 1645 712 1671
rect 770 1645 1170 1671
rect 1228 1645 1628 1671
rect 1686 1645 2086 1671
rect 2144 1645 2544 1671
rect 2602 1645 3002 1671
rect 3060 1645 3460 1671
rect 3518 1645 3918 1671
rect 3976 1645 4376 1671
rect 312 329 712 355
rect 770 329 1170 355
rect 1228 329 1628 355
rect 1686 329 2086 355
rect 2144 329 2544 355
rect 2602 329 3002 355
rect 3060 329 3460 355
rect 3518 329 3918 355
rect 3976 329 4376 355
rect 458 184 578 329
rect 914 184 1034 329
rect 1370 184 1490 329
rect 1826 184 1946 329
rect 2282 184 2402 329
rect 2738 184 2858 329
rect 3194 184 3314 329
rect 3650 184 3770 329
rect 4106 184 4226 329
rect 218 164 4470 184
rect 218 104 388 164
rect 448 104 788 164
rect 848 104 1188 164
rect 1248 104 1588 164
rect 1648 104 1988 164
rect 2048 104 2388 164
rect 2448 104 2788 164
rect 2848 104 3188 164
rect 3248 104 3588 164
rect 3648 104 3988 164
rect 4048 104 4470 164
rect 218 84 4470 104
<< polycont >>
rect 388 104 448 164
rect 788 104 848 164
rect 1188 104 1248 164
rect 1588 104 1648 164
rect 1988 104 2048 164
rect 2388 104 2448 164
rect 2788 104 2848 164
rect 3188 104 3248 164
rect 3588 104 3648 164
rect 3988 104 4048 164
<< locali >>
rect 120 1850 388 1910
rect 448 1850 788 1910
rect 848 1850 1188 1910
rect 1248 1850 1588 1910
rect 1648 1850 1988 1910
rect 2048 1850 2388 1910
rect 2448 1850 2788 1910
rect 2848 1850 3188 1910
rect 3248 1850 3588 1910
rect 3648 1850 3988 1910
rect 4048 1850 4470 1910
rect 148 1760 208 1850
rect 1198 1808 1358 1850
rect 1198 1772 1258 1808
rect 1302 1772 1358 1808
rect 1198 1770 1358 1772
rect 2498 1808 2658 1850
rect 2498 1772 2558 1808
rect 2602 1772 2658 1808
rect 2498 1770 2658 1772
rect 148 1720 158 1760
rect 198 1720 208 1760
rect 148 1640 208 1720
rect 278 1690 4470 1730
rect 723 1649 757 1690
rect 1639 1649 1673 1690
rect 2555 1649 2589 1690
rect 3471 1649 3505 1690
rect 4387 1649 4421 1690
rect 266 1633 300 1649
rect 265 367 266 374
rect 723 1633 758 1649
rect 723 1626 724 1633
rect 265 351 300 367
rect 1182 1633 1216 1649
rect 724 351 758 367
rect 1181 367 1182 374
rect 1639 1633 1674 1649
rect 1639 1626 1640 1633
rect 1181 351 1216 367
rect 2098 1633 2132 1649
rect 1640 351 1674 367
rect 2097 367 2098 374
rect 2555 1633 2590 1649
rect 2555 1626 2556 1633
rect 2097 351 2132 367
rect 3014 1633 3048 1649
rect 2556 351 2590 367
rect 3013 367 3014 374
rect 3471 1633 3506 1649
rect 3471 1626 3472 1633
rect 3013 351 3048 367
rect 3930 1633 3964 1649
rect 3472 351 3506 367
rect 3929 367 3930 374
rect 4387 1633 4422 1649
rect 4387 1626 4388 1633
rect 3929 351 3964 367
rect 4388 351 4422 367
rect 265 270 299 351
rect 1181 270 1215 351
rect 2097 270 2131 351
rect 3013 270 3047 351
rect 3929 270 3963 351
rect 218 210 4470 270
rect 218 104 388 164
rect 448 104 788 164
rect 848 104 1188 164
rect 1248 104 1588 164
rect 1648 104 1988 164
rect 2048 104 2388 164
rect 2448 104 2788 164
rect 2848 104 3188 164
rect 3248 104 3588 164
rect 3648 104 3988 164
rect 4048 104 4470 164
rect 120 -30 388 30
rect 448 -30 788 30
rect 848 -30 1188 30
rect 1248 -30 1588 30
rect 1648 -30 1988 30
rect 2048 -30 2388 30
rect 2448 -30 2788 30
rect 2848 -30 3188 30
rect 3248 -30 3588 30
rect 3648 -30 3988 30
rect 4048 -30 4470 30
<< viali >>
rect 388 1850 448 1910
rect 788 1850 848 1910
rect 1188 1850 1248 1910
rect 1588 1850 1648 1910
rect 1988 1850 2048 1910
rect 2388 1850 2448 1910
rect 2788 1850 2848 1910
rect 3188 1850 3248 1910
rect 3588 1850 3648 1910
rect 3988 1850 4048 1910
rect 266 367 300 1633
rect 724 367 758 1633
rect 1182 367 1216 1633
rect 1640 367 1674 1633
rect 2098 367 2132 1633
rect 2556 367 2590 1633
rect 3014 367 3048 1633
rect 3472 367 3506 1633
rect 3930 367 3964 1633
rect 4388 367 4422 1633
rect 388 -30 448 30
rect 788 -30 848 30
rect 1188 -30 1248 30
rect 1588 -30 1648 30
rect 1988 -30 2048 30
rect 2388 -30 2448 30
rect 2788 -30 2848 30
rect 3188 -30 3248 30
rect 3588 -30 3648 30
rect 3988 -30 4048 30
<< metal1 >>
rect 120 1910 4470 1940
rect 120 1850 388 1910
rect 448 1850 788 1910
rect 848 1850 1188 1910
rect 1248 1850 1588 1910
rect 1648 1850 1988 1910
rect 2048 1850 2388 1910
rect 2448 1850 2788 1910
rect 2848 1850 3188 1910
rect 3248 1850 3588 1910
rect 3648 1850 3988 1910
rect 4048 1850 4470 1910
rect 120 1820 4470 1850
rect 260 1633 306 1645
rect 260 367 266 1633
rect 300 367 306 1633
rect 260 355 306 367
rect 718 1633 764 1645
rect 718 367 724 1633
rect 758 367 764 1633
rect 718 355 764 367
rect 1176 1633 1222 1645
rect 1176 367 1182 1633
rect 1216 367 1222 1633
rect 1176 355 1222 367
rect 1634 1633 1680 1645
rect 1634 367 1640 1633
rect 1674 367 1680 1633
rect 1634 355 1680 367
rect 2092 1633 2138 1645
rect 2092 367 2098 1633
rect 2132 367 2138 1633
rect 2092 355 2138 367
rect 2550 1633 2596 1645
rect 2550 367 2556 1633
rect 2590 367 2596 1633
rect 2550 355 2596 367
rect 3008 1633 3054 1645
rect 3008 367 3014 1633
rect 3048 367 3054 1633
rect 3008 355 3054 367
rect 3466 1633 3512 1645
rect 3466 367 3472 1633
rect 3506 367 3512 1633
rect 3466 355 3512 367
rect 3924 1633 3970 1645
rect 3924 367 3930 1633
rect 3964 367 3970 1633
rect 3924 355 3970 367
rect 4382 1633 4428 1645
rect 4382 367 4388 1633
rect 4422 367 4428 1633
rect 4382 355 4428 367
rect 120 30 4470 60
rect 120 -30 388 30
rect 448 -30 788 30
rect 848 -30 1188 30
rect 1248 -30 1588 30
rect 1648 -30 1988 30
rect 2048 -30 2388 30
rect 2448 -30 2788 30
rect 2848 -30 3188 30
rect 3248 -30 3588 30
rect 3648 -30 3988 30
rect 4048 -30 4470 30
rect 120 -60 4470 -30
<< labels >>
flabel nwell 120 1850 180 1910 1 FreeSans 800 0 0 0 VPWR
port 4 n power bidirectional
flabel metal1 120 -30 278 30 1 FreeSans 800 0 0 0 VGND
port 5 n ground bidirectional
flabel locali 4410 1690 4470 1730 1 FreeSans 800 0 0 0 SOURCE
port 2 n signal bidirectional
flabel locali 4410 210 4470 270 1 FreeSans 800 0 0 0 DRAIN
port 3 n signal bidirectional
flabel locali 4410 104 4470 164 1 FreeSans 800 0 0 0 GATE
port 1 n signal bidirectional
<< properties >>
string FIXED_BBOX 0 0 4770 1880
string LEFclass CORE
string LEFsite unitasc
<< end >>
