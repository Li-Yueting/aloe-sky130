VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO sky130_asc_pfet_01v8_lvt_9
  CLASS CORE ;
  FOREIGN sky130_asc_pfet_01v8_lvt_9 ;
  ORIGIN 0.000 0.000 ;
  SIZE 23.850 BY 9.400 ;
  SITE unitasc ;
  PIN GATE
    DIRECTION INOUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 116.099998 ;
    PORT
      LAYER li1 ;
        RECT 0.650 0.510 21.910 0.810 ;
    END
  END GATE
  PIN SOURCE
    DIRECTION INOUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 9.352500 ;
    PORT
      LAYER li1 ;
        RECT 0.650 8.650 21.910 8.950 ;
        RECT 3.175 8.245 3.345 8.650 ;
        RECT 7.755 8.245 7.925 8.650 ;
        RECT 12.335 8.245 12.505 8.650 ;
        RECT 16.915 8.245 17.085 8.650 ;
        RECT 21.495 8.245 21.665 8.650 ;
        RECT 3.175 8.130 3.350 8.245 ;
        RECT 7.755 8.130 7.930 8.245 ;
        RECT 12.335 8.130 12.510 8.245 ;
        RECT 16.915 8.130 17.090 8.245 ;
        RECT 21.495 8.130 21.670 8.245 ;
        RECT 3.180 1.755 3.350 8.130 ;
        RECT 7.760 1.755 7.930 8.130 ;
        RECT 12.340 1.755 12.510 8.130 ;
        RECT 16.920 1.755 17.090 8.130 ;
        RECT 21.500 1.755 21.670 8.130 ;
      LAYER mcon ;
        RECT 3.180 1.835 3.350 8.165 ;
        RECT 7.760 1.835 7.930 8.165 ;
        RECT 12.340 1.835 12.510 8.165 ;
        RECT 16.920 1.835 17.090 8.165 ;
        RECT 21.500 1.835 21.670 8.165 ;
      LAYER met1 ;
        RECT 3.150 1.775 3.380 8.225 ;
        RECT 7.730 1.775 7.960 8.225 ;
        RECT 12.310 1.775 12.540 8.225 ;
        RECT 16.890 1.775 17.120 8.225 ;
        RECT 21.470 1.775 21.700 8.225 ;
    END
  END SOURCE
  PIN DRAIN
    DIRECTION INOUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 9.352500 ;
    PORT
      LAYER li1 ;
        RECT 0.890 1.860 1.060 8.245 ;
        RECT 5.470 1.860 5.640 8.245 ;
        RECT 10.050 1.860 10.220 8.245 ;
        RECT 14.630 1.860 14.800 8.245 ;
        RECT 19.210 1.860 19.380 8.245 ;
        RECT 0.885 1.755 1.060 1.860 ;
        RECT 5.465 1.755 5.640 1.860 ;
        RECT 10.045 1.755 10.220 1.860 ;
        RECT 14.625 1.755 14.800 1.860 ;
        RECT 19.205 1.755 19.380 1.860 ;
        RECT 0.885 1.350 1.055 1.755 ;
        RECT 5.465 1.350 5.635 1.755 ;
        RECT 10.045 1.350 10.215 1.755 ;
        RECT 14.625 1.350 14.795 1.755 ;
        RECT 19.205 1.350 19.375 1.755 ;
        RECT 0.650 1.050 21.910 1.350 ;
      LAYER mcon ;
        RECT 0.890 1.835 1.060 8.165 ;
        RECT 5.470 1.835 5.640 8.165 ;
        RECT 10.050 1.835 10.220 8.165 ;
        RECT 14.630 1.835 14.800 8.165 ;
        RECT 19.210 1.835 19.380 8.165 ;
      LAYER met1 ;
        RECT 0.860 1.775 1.090 8.225 ;
        RECT 5.440 1.775 5.670 8.225 ;
        RECT 10.020 1.775 10.250 8.225 ;
        RECT 14.600 1.775 14.830 8.225 ;
        RECT 19.180 1.775 19.410 8.225 ;
    END
  END DRAIN
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER li1 ;
        RECT 0.650 9.250 21.910 9.550 ;
      LAYER mcon ;
        RECT 1.500 9.250 1.800 9.550 ;
        RECT 3.500 9.250 3.800 9.550 ;
        RECT 5.500 9.250 5.800 9.550 ;
        RECT 7.500 9.250 7.800 9.550 ;
        RECT 9.500 9.250 9.800 9.550 ;
        RECT 11.500 9.250 11.800 9.550 ;
        RECT 13.500 9.250 13.800 9.550 ;
        RECT 15.500 9.250 15.800 9.550 ;
        RECT 17.500 9.250 17.800 9.550 ;
        RECT 19.500 9.250 19.800 9.550 ;
      LAYER met1 ;
        RECT 0.650 9.100 21.910 9.700 ;
    END
  END VPWR
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER li1 ;
        RECT 0.650 -0.150 21.910 0.150 ;
      LAYER mcon ;
        RECT 1.500 -0.150 1.800 0.150 ;
        RECT 3.500 -0.150 3.800 0.150 ;
        RECT 5.500 -0.150 5.800 0.150 ;
        RECT 7.500 -0.150 7.800 0.150 ;
        RECT 9.500 -0.150 9.800 0.150 ;
        RECT 11.500 -0.150 11.800 0.150 ;
        RECT 13.500 -0.150 13.800 0.150 ;
        RECT 15.500 -0.150 15.800 0.150 ;
        RECT 17.500 -0.150 17.800 0.150 ;
        RECT 19.500 -0.150 19.800 0.150 ;
      LAYER met1 ;
        RECT 0.650 -0.300 21.910 0.300 ;
    END
  END VGND
  OBS
      LAYER nwell ;
        RECT 0.650 1.465 21.910 9.700 ;
  END
END sky130_asc_pfet_01v8_lvt_9
END LIBRARY

