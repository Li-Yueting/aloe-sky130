VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO ls
  CLASS CORE ;
  FOREIGN ls ;
  ORIGIN 0.000 0.000 ;
  SIZE 4.270 BY 9.400 ;
  SITE unitasc ;
  PIN GATE
    DIRECTION INOUT ;
    ANTENNAGATEAREA 10.000000 ;
    PORT
      LAYER li1 ;
        RECT 1.490 1.020 3.670 1.320 ;
    END
  END GATE
  PIN SOURCE
    DIRECTION INOUT ;
    ANTENNADIFFAREA 1.450000 ;
    PORT
      LAYER li1 ;
        RECT 1.090 8.450 3.670 8.750 ;
        RECT 3.435 7.520 3.605 8.450 ;
        RECT 3.435 7.430 3.610 7.520 ;
        RECT 3.440 2.480 3.610 7.430 ;
      LAYER mcon ;
        RECT 3.440 2.560 3.610 7.440 ;
      LAYER met1 ;
        RECT 3.410 2.500 3.640 7.500 ;
    END
  END SOURCE
  PIN DRAIN
    DIRECTION INOUT ;
    ANTENNADIFFAREA 1.450000 ;
    PORT
      LAYER li1 ;
        RECT 1.150 2.770 1.320 7.520 ;
        RECT 1.145 2.480 1.320 2.770 ;
        RECT 1.145 2.150 1.315 2.480 ;
        RECT 1.090 1.850 3.670 2.150 ;
      LAYER mcon ;
        RECT 1.150 2.560 1.320 7.440 ;
      LAYER met1 ;
        RECT 1.120 2.500 1.350 7.500 ;
    END
  END DRAIN
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER li1 ;
        RECT 0.600 9.250 3.670 9.550 ;
      LAYER mcon ;
        RECT 1.940 9.250 2.240 9.550 ;
      LAYER met1 ;
        RECT 0.600 9.100 3.670 9.700 ;
    END
  END VPWR
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.600 0.150 3.670 7.630 ;
      LAYER li1 ;
        RECT 0.740 0.150 1.040 1.200 ;
        RECT 0.600 -0.150 3.670 0.150 ;
      LAYER mcon ;
        RECT 1.940 -0.150 2.240 0.150 ;
      LAYER met1 ;
        RECT 0.600 -0.300 3.670 0.300 ;
    END
  END VGND
END ls
END LIBRARY

