VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO sky130_asc_pnp_05v5_W3p40L3p40_1
  CLASS CORE ;
  FOREIGN sky130_asc_pnp_05v5_W3p40L3p40_1 ;
  ORIGIN 0.000 0.000 ;
  SIZE 7.600 BY 9.400 ;
  SITE unitasc ;
  PIN Emitter
    DIRECTION INOUT ;
    ANTENNADIFFAREA 11.559999 ;
    PORT
      LAYER li1 ;
        RECT 2.065 2.965 5.535 6.435 ;
      LAYER mcon ;
        RECT 2.430 5.830 2.600 6.000 ;
        RECT 2.930 5.830 3.100 6.000 ;
        RECT 3.430 5.830 3.600 6.000 ;
        RECT 3.930 5.830 4.100 6.000 ;
        RECT 4.430 5.830 4.600 6.000 ;
        RECT 4.930 5.830 5.100 6.000 ;
        RECT 2.430 5.330 2.600 5.500 ;
        RECT 2.930 5.330 3.100 5.500 ;
        RECT 3.430 5.330 3.600 5.500 ;
        RECT 3.930 5.330 4.100 5.500 ;
        RECT 4.430 5.330 4.600 5.500 ;
        RECT 4.930 5.330 5.100 5.500 ;
        RECT 2.430 4.830 2.600 5.000 ;
        RECT 2.930 4.830 3.100 5.000 ;
        RECT 3.430 4.830 3.600 5.000 ;
        RECT 3.930 4.830 4.100 5.000 ;
        RECT 4.430 4.830 4.600 5.000 ;
        RECT 4.930 4.830 5.100 5.000 ;
        RECT 2.430 4.330 2.600 4.500 ;
        RECT 2.930 4.330 3.100 4.500 ;
        RECT 3.430 4.330 3.600 4.500 ;
        RECT 3.930 4.330 4.100 4.500 ;
        RECT 4.430 4.330 4.600 4.500 ;
        RECT 4.930 4.330 5.100 4.500 ;
        RECT 2.430 3.830 2.600 4.000 ;
        RECT 2.930 3.830 3.100 4.000 ;
        RECT 3.430 3.830 3.600 4.000 ;
        RECT 3.930 3.830 4.100 4.000 ;
        RECT 4.430 3.830 4.600 4.000 ;
        RECT 4.930 3.830 5.100 4.000 ;
        RECT 2.430 3.330 2.600 3.500 ;
        RECT 2.930 3.330 3.100 3.500 ;
        RECT 3.430 3.330 3.600 3.500 ;
        RECT 3.930 3.330 4.100 3.500 ;
        RECT 4.430 3.330 4.600 3.500 ;
        RECT 4.930 3.330 5.100 3.500 ;
      LAYER met1 ;
        RECT 2.275 3.175 5.325 6.225 ;
    END
  END Emitter
  PIN Base
    DIRECTION INOUT ;
    ANTENNAGATEAREA 26.728899 ;
    ANTENNADIFFAREA 6.408000 ;
    PORT
      LAYER li1 ;
        RECT 1.395 6.745 6.205 7.105 ;
        RECT 1.395 2.655 1.755 6.745 ;
        RECT 5.845 2.655 6.205 6.745 ;
        RECT 1.395 2.295 6.205 2.655 ;
    END
  END Base
  PIN Collector
    DIRECTION INOUT ;
    ANTENNADIFFAREA 11.988700 ;
    PORT
      LAYER pwell ;
        RECT 0.450 7.285 7.150 8.050 ;
        RECT 0.450 2.115 1.215 7.285 ;
        RECT 6.385 2.115 7.150 7.285 ;
        RECT 0.450 1.350 7.150 2.115 ;
      LAYER li1 ;
        RECT 0.580 7.425 7.020 7.920 ;
        RECT 0.580 1.975 1.075 7.425 ;
        RECT 6.525 1.975 7.020 7.425 ;
        RECT 0.580 1.480 7.020 1.975 ;
    END
  END Collector
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER li1 ;
        RECT 0.450 9.250 7.150 9.550 ;
      LAYER mcon ;
        RECT 1.300 9.250 1.600 9.550 ;
        RECT 2.300 9.250 2.600 9.550 ;
        RECT 3.300 9.250 3.600 9.550 ;
        RECT 4.300 9.250 4.600 9.550 ;
        RECT 5.300 9.250 5.600 9.550 ;
        RECT 6.300 9.250 6.600 9.550 ;
      LAYER met1 ;
        RECT 0.450 9.100 7.150 9.700 ;
    END
  END VPWR
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER li1 ;
        RECT 0.450 -0.150 7.150 0.150 ;
      LAYER mcon ;
        RECT 1.300 -0.150 1.600 0.150 ;
        RECT 2.300 -0.150 2.600 0.150 ;
        RECT 3.300 -0.150 3.600 0.150 ;
        RECT 4.300 -0.150 4.600 0.150 ;
        RECT 5.300 -0.150 5.600 0.150 ;
        RECT 6.300 -0.150 6.600 0.150 ;
      LAYER met1 ;
        RECT 0.450 -0.300 7.150 0.300 ;
    END
  END VGND
END sky130_asc_pnp_05v5_W3p40L3p40_1
END LIBRARY

