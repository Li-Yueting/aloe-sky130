magic
tech sky130A
magscale 1 2
timestamp 1652221573
<< nwell >>
rect 0 1707 2974 1940
rect 0 294 2975 1707
rect 97 293 2975 294
<< pmoslvt >>
rect 191 355 591 1645
rect 649 355 1049 1645
rect 1107 355 1507 1645
rect 1565 355 1965 1645
rect 2023 355 2423 1645
rect 2481 355 2881 1645
<< pdiff >>
rect 133 1633 191 1645
rect 133 367 145 1633
rect 179 367 191 1633
rect 133 355 191 367
rect 591 1633 649 1645
rect 591 367 603 1633
rect 637 367 649 1633
rect 591 355 649 367
rect 1049 1633 1107 1645
rect 1049 367 1061 1633
rect 1095 367 1107 1633
rect 1049 355 1107 367
rect 1507 1633 1565 1645
rect 1507 367 1519 1633
rect 1553 367 1565 1633
rect 1507 355 1565 367
rect 1965 1633 2023 1645
rect 1965 367 1977 1633
rect 2011 367 2023 1633
rect 1965 355 2023 367
rect 2423 1633 2481 1645
rect 2423 367 2435 1633
rect 2469 367 2481 1633
rect 2423 355 2481 367
rect 2881 1633 2939 1645
rect 2881 367 2893 1633
rect 2927 367 2939 1633
rect 2881 355 2939 367
<< pdiffc >>
rect 145 367 179 1633
rect 603 367 637 1633
rect 1061 367 1095 1633
rect 1519 367 1553 1633
rect 1977 367 2011 1633
rect 2435 367 2469 1633
rect 2893 367 2927 1633
<< nsubdiff >>
rect 38 1760 78 1800
rect 38 1680 78 1720
<< nsubdiffcont >>
rect 38 1720 78 1760
<< poly >>
rect 191 1645 591 1671
rect 649 1645 1049 1671
rect 1107 1645 1507 1671
rect 1565 1645 1965 1671
rect 2023 1645 2423 1671
rect 2481 1645 2881 1671
rect 191 329 591 355
rect 649 329 1049 355
rect 1107 329 1507 355
rect 1565 329 1965 355
rect 2023 329 2423 355
rect 2481 329 2881 355
rect 338 184 458 329
rect 794 184 914 329
rect 1250 184 1370 329
rect 1706 184 1826 329
rect 2162 184 2282 329
rect 2618 184 2738 329
rect 98 164 2974 184
rect 98 104 268 164
rect 328 104 668 164
rect 728 104 1068 164
rect 1128 104 1468 164
rect 1528 104 1868 164
rect 1928 104 2268 164
rect 2328 104 2668 164
rect 2728 104 2974 164
rect 98 84 2974 104
<< polycont >>
rect 268 104 328 164
rect 668 104 728 164
rect 1068 104 1128 164
rect 1468 104 1528 164
rect 1868 104 1928 164
rect 2268 104 2328 164
rect 2668 104 2728 164
<< locali >>
rect 0 1850 268 1910
rect 328 1850 668 1910
rect 728 1850 1068 1910
rect 1128 1850 1468 1910
rect 1528 1850 1868 1910
rect 1928 1850 2268 1910
rect 2328 1850 2668 1910
rect 2728 1850 2974 1910
rect 28 1760 88 1850
rect 28 1720 38 1760
rect 78 1720 88 1760
rect 158 1730 2974 1790
rect 28 1640 88 1720
rect 145 1633 179 1649
rect 145 270 179 367
rect 603 1633 637 1730
rect 603 351 637 367
rect 1061 1633 1095 1649
rect 1061 270 1095 367
rect 1519 1633 1553 1730
rect 1519 351 1553 367
rect 1977 1633 2011 1649
rect 1977 270 2011 367
rect 2435 1633 2469 1730
rect 2435 351 2469 367
rect 2893 1633 2927 1649
rect 2893 270 2927 367
rect 98 210 2974 270
rect 98 104 268 164
rect 328 104 668 164
rect 728 104 1068 164
rect 1128 104 1468 164
rect 1528 104 1868 164
rect 1928 104 2268 164
rect 2328 104 2668 164
rect 2728 104 2974 164
rect 0 -30 268 30
rect 328 -30 668 30
rect 728 -30 1068 30
rect 1128 -30 1468 30
rect 1528 -30 1868 30
rect 1928 -30 2268 30
rect 2328 -30 2668 30
rect 2728 -30 2974 30
<< viali >>
rect 268 1850 328 1910
rect 668 1850 728 1910
rect 1068 1850 1128 1910
rect 1468 1850 1528 1910
rect 1868 1850 1928 1910
rect 2268 1850 2328 1910
rect 2668 1850 2728 1910
rect 145 367 179 1633
rect 603 367 637 1633
rect 1061 367 1095 1633
rect 1519 367 1553 1633
rect 1977 367 2011 1633
rect 2435 367 2469 1633
rect 2893 367 2927 1633
rect 268 -30 328 30
rect 668 -30 728 30
rect 1068 -30 1128 30
rect 1468 -30 1528 30
rect 1868 -30 1928 30
rect 2268 -30 2328 30
rect 2668 -30 2728 30
<< metal1 >>
rect 0 1910 2974 1940
rect 0 1850 268 1910
rect 328 1850 668 1910
rect 728 1850 1068 1910
rect 1128 1850 1468 1910
rect 1528 1850 1868 1910
rect 1928 1850 2268 1910
rect 2328 1850 2668 1910
rect 2728 1850 2974 1910
rect 0 1820 2974 1850
rect 139 1633 185 1645
rect 139 367 145 1633
rect 179 367 185 1633
rect 139 355 185 367
rect 597 1633 643 1645
rect 597 367 603 1633
rect 637 367 643 1633
rect 597 355 643 367
rect 1055 1633 1101 1645
rect 1055 367 1061 1633
rect 1095 367 1101 1633
rect 1055 355 1101 367
rect 1513 1633 1559 1645
rect 1513 367 1519 1633
rect 1553 367 1559 1633
rect 1513 355 1559 367
rect 1971 1633 2017 1645
rect 1971 367 1977 1633
rect 2011 367 2017 1633
rect 1971 355 2017 367
rect 2429 1633 2475 1645
rect 2429 367 2435 1633
rect 2469 367 2475 1633
rect 2429 355 2475 367
rect 2887 1633 2933 1645
rect 2887 367 2893 1633
rect 2927 367 2933 1633
rect 2887 355 2933 367
rect 0 30 2974 60
rect 0 -30 268 30
rect 328 -30 668 30
rect 728 -30 1068 30
rect 1128 -30 1468 30
rect 1528 -30 1868 30
rect 1928 -30 2268 30
rect 2328 -30 2668 30
rect 2728 -30 2974 30
rect 0 -60 2974 -30
<< labels >>
flabel nwell 0 1850 60 1910 1 FreeSans 800 0 0 0 VPWR
port 4 n power bidirectional
flabel metal1 0 -30 158 30 1 FreeSans 800 0 0 0 VGND
port 5 n ground bidirectional
flabel locali 2914 1730 2974 1790 1 FreeSans 800 0 0 0 SOURCE
port 2 n signal bidirectional
flabel locali 2914 210 2974 270 1 FreeSans 800 0 0 0 DRAIN
port 3 n signal bidirectional
flabel locali 2914 104 2974 164 1 FreeSans 800 0 0 0 GATE
port 1 n signal bidirectional
<< properties >>
string FIXED_BBOX 0 0 2975 1880
string LEFclass CORE
string LEFsite unitasc
<< end >>
