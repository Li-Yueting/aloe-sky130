magic
tech sky130A
magscale 1 2
timestamp 1654749236
<< pwell >>
rect -284 -426 284 426
rect -344 -946 -252 -774
<< nmoslvt >>
rect -200 -400 200 400
<< ndiff >>
rect -258 357 -200 400
rect -258 323 -246 357
rect -212 323 -200 357
rect -258 289 -200 323
rect -258 255 -246 289
rect -212 255 -200 289
rect -258 221 -200 255
rect -258 187 -246 221
rect -212 187 -200 221
rect -258 153 -200 187
rect -258 119 -246 153
rect -212 119 -200 153
rect -258 85 -200 119
rect -258 51 -246 85
rect -212 51 -200 85
rect -258 17 -200 51
rect -258 -17 -246 17
rect -212 -17 -200 17
rect -258 -51 -200 -17
rect -258 -85 -246 -51
rect -212 -85 -200 -51
rect -258 -119 -200 -85
rect -258 -153 -246 -119
rect -212 -153 -200 -119
rect -258 -187 -200 -153
rect -258 -221 -246 -187
rect -212 -221 -200 -187
rect -258 -255 -200 -221
rect -258 -289 -246 -255
rect -212 -289 -200 -255
rect -258 -323 -200 -289
rect -258 -357 -246 -323
rect -212 -357 -200 -323
rect -258 -400 -200 -357
rect 200 357 258 400
rect 200 323 212 357
rect 246 323 258 357
rect 200 289 258 323
rect 200 255 212 289
rect 246 255 258 289
rect 200 221 258 255
rect 200 187 212 221
rect 246 187 258 221
rect 200 153 258 187
rect 200 119 212 153
rect 246 119 258 153
rect 200 85 258 119
rect 200 51 212 85
rect 246 51 258 85
rect 200 17 258 51
rect 200 -17 212 17
rect 246 -17 258 17
rect 200 -51 258 -17
rect 200 -85 212 -51
rect 246 -85 258 -51
rect 200 -119 258 -85
rect 200 -153 212 -119
rect 246 -153 258 -119
rect 200 -187 258 -153
rect 200 -221 212 -187
rect 246 -221 258 -187
rect 200 -255 258 -221
rect 200 -289 212 -255
rect 246 -289 258 -255
rect 200 -323 258 -289
rect 200 -357 212 -323
rect 246 -357 258 -323
rect 200 -400 258 -357
<< ndiffc >>
rect -246 323 -212 357
rect -246 255 -212 289
rect -246 187 -212 221
rect -246 119 -212 153
rect -246 51 -212 85
rect -246 -17 -212 17
rect -246 -85 -212 -51
rect -246 -153 -212 -119
rect -246 -221 -212 -187
rect -246 -289 -212 -255
rect -246 -357 -212 -323
rect 212 323 246 357
rect 212 255 246 289
rect 212 187 246 221
rect 212 119 246 153
rect 212 51 246 85
rect 212 -17 246 17
rect 212 -85 246 -51
rect 212 -153 246 -119
rect 212 -221 246 -187
rect 212 -289 246 -255
rect 212 -357 246 -323
<< psubdiff >>
rect -318 -843 -278 -800
rect -318 -877 -315 -843
rect -281 -877 -278 -843
rect -318 -920 -278 -877
<< psubdiffcont >>
rect -315 -877 -281 -843
<< poly >>
rect -200 400 200 426
rect -200 -426 200 -400
rect -52 -616 68 -426
rect -178 -649 258 -616
rect -178 -683 -75 -649
rect -41 -683 258 -649
rect -178 -716 258 -683
<< polycont >>
rect -75 -683 -41 -649
<< locali >>
rect -356 897 258 910
rect -356 863 -75 897
rect -41 863 258 897
rect -356 850 258 863
rect -258 690 258 750
rect 211 404 245 690
rect -246 377 -212 404
rect 211 386 246 404
rect -246 305 -212 323
rect -246 233 -212 255
rect -246 161 -212 187
rect -246 89 -212 119
rect -246 17 -212 51
rect -246 -51 -212 -17
rect -246 -119 -212 -89
rect -246 -187 -212 -161
rect -246 -255 -212 -233
rect -246 -323 -212 -305
rect -247 -377 -246 -346
rect -247 -404 -212 -377
rect 212 377 246 386
rect 212 305 246 323
rect 212 233 246 255
rect 212 161 246 187
rect 212 89 246 119
rect 212 17 246 51
rect 212 -51 246 -17
rect 212 -119 246 -89
rect 212 -187 246 -161
rect 212 -255 246 -233
rect 212 -323 246 -305
rect 212 -404 246 -377
rect -247 -470 -213 -404
rect -258 -530 258 -470
rect -178 -649 258 -636
rect -178 -683 -75 -649
rect -41 -683 258 -649
rect -178 -696 258 -683
rect -328 -843 -268 -760
rect -328 -877 -315 -843
rect -281 -877 -268 -843
rect -328 -970 -268 -877
rect -356 -983 258 -970
rect -356 -1017 -75 -983
rect -41 -1017 258 -983
rect -356 -1030 258 -1017
<< viali >>
rect -75 863 -41 897
rect -246 357 -212 377
rect -246 343 -212 357
rect -246 289 -212 305
rect -246 271 -212 289
rect -246 221 -212 233
rect -246 199 -212 221
rect -246 153 -212 161
rect -246 127 -212 153
rect -246 85 -212 89
rect -246 55 -212 85
rect -246 -17 -212 17
rect -246 -85 -212 -55
rect -246 -89 -212 -85
rect -246 -153 -212 -127
rect -246 -161 -212 -153
rect -246 -221 -212 -199
rect -246 -233 -212 -221
rect -246 -289 -212 -271
rect -246 -305 -212 -289
rect -246 -357 -212 -343
rect -246 -377 -212 -357
rect 212 357 246 377
rect 212 343 246 357
rect 212 289 246 305
rect 212 271 246 289
rect 212 221 246 233
rect 212 199 246 221
rect 212 153 246 161
rect 212 127 246 153
rect 212 85 246 89
rect 212 55 246 85
rect 212 -17 246 17
rect 212 -85 246 -55
rect 212 -89 246 -85
rect 212 -153 246 -127
rect 212 -161 246 -153
rect 212 -221 246 -199
rect 212 -233 246 -221
rect 212 -289 246 -271
rect 212 -305 246 -289
rect 212 -357 246 -343
rect 212 -377 246 -357
rect -75 -1017 -41 -983
<< metal1 >>
rect -356 897 258 940
rect -356 863 -75 897
rect -41 863 258 897
rect -356 820 258 863
rect -252 377 -206 400
rect -252 343 -246 377
rect -212 343 -206 377
rect -252 305 -206 343
rect -252 271 -246 305
rect -212 271 -206 305
rect -252 233 -206 271
rect -252 199 -246 233
rect -212 199 -206 233
rect -252 161 -206 199
rect -252 127 -246 161
rect -212 127 -206 161
rect -252 89 -206 127
rect -252 55 -246 89
rect -212 55 -206 89
rect -252 17 -206 55
rect -252 -17 -246 17
rect -212 -17 -206 17
rect -252 -55 -206 -17
rect -252 -89 -246 -55
rect -212 -89 -206 -55
rect -252 -127 -206 -89
rect -252 -161 -246 -127
rect -212 -161 -206 -127
rect -252 -199 -206 -161
rect -252 -233 -246 -199
rect -212 -233 -206 -199
rect -252 -271 -206 -233
rect -252 -305 -246 -271
rect -212 -305 -206 -271
rect -252 -343 -206 -305
rect -252 -377 -246 -343
rect -212 -377 -206 -343
rect -252 -400 -206 -377
rect 206 377 252 400
rect 206 343 212 377
rect 246 343 252 377
rect 206 305 252 343
rect 206 271 212 305
rect 246 271 252 305
rect 206 233 252 271
rect 206 199 212 233
rect 246 199 252 233
rect 206 161 252 199
rect 206 127 212 161
rect 246 127 252 161
rect 206 89 252 127
rect 206 55 212 89
rect 246 55 252 89
rect 206 17 252 55
rect 206 -17 212 17
rect 246 -17 252 17
rect 206 -55 252 -17
rect 206 -89 212 -55
rect 246 -89 252 -55
rect 206 -127 252 -89
rect 206 -161 212 -127
rect 246 -161 252 -127
rect 206 -199 252 -161
rect 206 -233 212 -199
rect 246 -233 252 -199
rect 206 -271 252 -233
rect 206 -305 212 -271
rect 246 -305 252 -271
rect 206 -343 252 -305
rect 206 -377 212 -343
rect 246 -377 252 -343
rect 206 -400 252 -377
rect -356 -983 258 -940
rect -356 -1017 -75 -983
rect -41 -1017 258 -983
rect -356 -1060 258 -1017
<< labels >>
flabel metal1 s -258 850 -198 910 1 FreeSans 1000 0 0 0 VPWR
port 1 nsew
flabel metal1 s -258 -1030 -198 -970 1 FreeSans 1000 0 0 0 VGND
port 2 nsew
flabel locali s 198 690 258 750 1 FreeSans 1000 0 0 0 SOURCE
port 3 nsew
flabel locali s 198 -530 258 -470 1 FreeSans 1000 0 0 0 DRAIN
port 4 nsew
flabel locali s 198 -696 258 -636 1 FreeSans 1000 0 0 0 GATE
port 5 nsew
<< end >>
