magic
tech sky130A
magscale 1 2
timestamp 1653360443
<< pwell >>
rect 90 30 4368 1426
<< nmoslvt >>
rect 246 600 646 1400
rect 704 600 1104 1400
rect 1162 600 1562 1400
rect 1620 600 2020 1400
rect 2078 600 2478 1400
rect 2536 600 2936 1400
rect 2994 600 3394 1400
rect 3452 600 3852 1400
rect 3910 600 4310 1400
<< ndiff >>
rect 188 1388 246 1400
rect 188 612 200 1388
rect 234 612 246 1388
rect 188 600 246 612
rect 646 1388 704 1400
rect 646 612 658 1388
rect 692 612 704 1388
rect 646 600 704 612
rect 1104 1388 1162 1400
rect 1104 612 1116 1388
rect 1150 612 1162 1388
rect 1104 600 1162 612
rect 1562 1388 1620 1400
rect 1562 612 1574 1388
rect 1608 612 1620 1388
rect 1562 600 1620 612
rect 2020 1388 2078 1400
rect 2020 612 2032 1388
rect 2066 612 2078 1388
rect 2020 600 2078 612
rect 2478 1388 2536 1400
rect 2478 612 2490 1388
rect 2524 612 2536 1388
rect 2478 600 2536 612
rect 2936 1388 2994 1400
rect 2936 612 2948 1388
rect 2982 612 2994 1388
rect 2936 600 2994 612
rect 3394 1388 3452 1400
rect 3394 612 3406 1388
rect 3440 612 3452 1388
rect 3394 600 3452 612
rect 3852 1388 3910 1400
rect 3852 612 3864 1388
rect 3898 612 3910 1388
rect 3852 600 3910 612
rect 4310 1388 4368 1400
rect 4310 612 4322 1388
rect 4356 612 4368 1388
rect 4310 600 4368 612
<< ndiffc >>
rect 200 612 234 1388
rect 658 612 692 1388
rect 1116 612 1150 1388
rect 1574 612 1608 1388
rect 2032 612 2066 1388
rect 2490 612 2524 1388
rect 2948 612 2982 1388
rect 3406 612 3440 1388
rect 3864 612 3898 1388
rect 4322 612 4356 1388
<< psubdiff >>
rect 128 160 168 200
rect 128 80 168 120
<< psubdiffcont >>
rect 128 120 168 160
<< poly >>
rect 246 1400 646 1426
rect 704 1400 1104 1426
rect 1162 1400 1562 1426
rect 1620 1400 2020 1426
rect 2078 1400 2478 1426
rect 2536 1400 2936 1426
rect 2994 1400 3394 1426
rect 3452 1400 3852 1426
rect 3910 1400 4310 1426
rect 246 574 646 600
rect 704 574 1104 600
rect 1162 574 1562 600
rect 1620 574 2020 600
rect 2078 574 2478 600
rect 2536 574 2936 600
rect 2994 574 3394 600
rect 3452 574 3852 600
rect 3910 574 4310 600
rect 394 224 514 574
rect 850 224 970 574
rect 1306 224 1426 574
rect 1762 224 1882 574
rect 2218 224 2338 574
rect 2674 224 2794 574
rect 3130 224 3250 574
rect 3586 224 3706 574
rect 4042 224 4162 574
rect 268 204 4368 224
rect 268 144 358 204
rect 418 144 758 204
rect 818 144 1158 204
rect 1218 144 1558 204
rect 1618 144 1958 204
rect 2018 144 2358 204
rect 2418 144 2758 204
rect 2818 144 3158 204
rect 3218 144 3558 204
rect 3618 144 3958 204
rect 4018 144 4368 204
rect 268 124 4368 144
<< polycont >>
rect 358 144 418 204
rect 758 144 818 204
rect 1158 144 1218 204
rect 1558 144 1618 204
rect 1958 144 2018 204
rect 2358 144 2418 204
rect 2758 144 2818 204
rect 3158 144 3218 204
rect 3558 144 3618 204
rect 3958 144 4018 204
<< locali >>
rect 90 1850 358 1910
rect 418 1850 758 1910
rect 818 1850 1158 1910
rect 1218 1850 1558 1910
rect 1618 1850 1958 1910
rect 2018 1850 2358 1910
rect 2418 1850 2758 1910
rect 2818 1850 3158 1910
rect 3218 1850 3558 1910
rect 3618 1850 3958 1910
rect 4018 1850 4368 1910
rect 188 1690 4368 1750
rect 657 1404 691 1690
rect 1573 1404 1607 1690
rect 2489 1404 2523 1690
rect 3405 1404 3439 1690
rect 4321 1404 4355 1690
rect 200 1388 234 1404
rect 199 612 200 654
rect 657 1388 692 1404
rect 657 1386 658 1388
rect 199 596 234 612
rect 1116 1388 1150 1404
rect 658 596 692 612
rect 1115 612 1116 654
rect 1573 1388 1608 1404
rect 1573 1386 1574 1388
rect 1115 596 1150 612
rect 2032 1388 2066 1404
rect 1574 596 1608 612
rect 2031 612 2032 654
rect 2489 1388 2524 1404
rect 2489 1386 2490 1388
rect 2031 596 2066 612
rect 2948 1388 2982 1404
rect 2490 596 2524 612
rect 2947 612 2948 654
rect 3405 1388 3440 1404
rect 3405 1386 3406 1388
rect 2947 596 2982 612
rect 3864 1388 3898 1404
rect 3406 596 3440 612
rect 3863 612 3864 654
rect 4321 1388 4356 1404
rect 4321 1386 4322 1388
rect 3863 596 3898 612
rect 4322 596 4356 612
rect 199 430 233 596
rect 1115 430 1149 596
rect 2031 430 2065 596
rect 2947 430 2981 596
rect 3863 430 3897 596
rect 188 370 4368 430
rect 118 160 178 240
rect 118 120 128 160
rect 168 120 178 160
rect 268 144 358 204
rect 418 144 758 204
rect 818 144 1158 204
rect 1218 144 1558 204
rect 1618 144 1958 204
rect 2018 144 2358 204
rect 2418 144 2758 204
rect 2818 144 3158 204
rect 3218 144 3558 204
rect 3618 144 3958 204
rect 4018 144 4368 204
rect 118 30 178 120
rect 90 -30 358 30
rect 418 -30 758 30
rect 818 -30 1158 30
rect 1218 -30 1558 30
rect 1618 -30 1958 30
rect 2018 -30 2358 30
rect 2418 -30 2758 30
rect 2818 -30 3158 30
rect 3218 -30 3558 30
rect 3618 -30 3958 30
rect 4018 -30 4368 30
<< viali >>
rect 358 1850 418 1910
rect 758 1850 818 1910
rect 1158 1850 1218 1910
rect 1558 1850 1618 1910
rect 1958 1850 2018 1910
rect 2358 1850 2418 1910
rect 2758 1850 2818 1910
rect 3158 1850 3218 1910
rect 3558 1850 3618 1910
rect 3958 1850 4018 1910
rect 200 612 234 1388
rect 658 612 692 1388
rect 1116 612 1150 1388
rect 1574 612 1608 1388
rect 2032 612 2066 1388
rect 2490 612 2524 1388
rect 2948 612 2982 1388
rect 3406 612 3440 1388
rect 3864 612 3898 1388
rect 4322 612 4356 1388
rect 358 -30 418 30
rect 758 -30 818 30
rect 1158 -30 1218 30
rect 1558 -30 1618 30
rect 1958 -30 2018 30
rect 2358 -30 2418 30
rect 2758 -30 2818 30
rect 3158 -30 3218 30
rect 3558 -30 3618 30
rect 3958 -30 4018 30
<< metal1 >>
rect 90 1910 4368 1940
rect 90 1850 358 1910
rect 418 1850 758 1910
rect 818 1850 1158 1910
rect 1218 1850 1558 1910
rect 1618 1850 1958 1910
rect 2018 1850 2358 1910
rect 2418 1850 2758 1910
rect 2818 1850 3158 1910
rect 3218 1850 3558 1910
rect 3618 1850 3958 1910
rect 4018 1850 4368 1910
rect 90 1820 4368 1850
rect 194 1388 240 1400
rect 194 612 200 1388
rect 234 612 240 1388
rect 194 600 240 612
rect 652 1388 698 1400
rect 652 612 658 1388
rect 692 612 698 1388
rect 652 600 698 612
rect 1110 1388 1156 1400
rect 1110 612 1116 1388
rect 1150 612 1156 1388
rect 1110 600 1156 612
rect 1568 1388 1614 1400
rect 1568 612 1574 1388
rect 1608 612 1614 1388
rect 1568 600 1614 612
rect 2026 1388 2072 1400
rect 2026 612 2032 1388
rect 2066 612 2072 1388
rect 2026 600 2072 612
rect 2484 1388 2530 1400
rect 2484 612 2490 1388
rect 2524 612 2530 1388
rect 2484 600 2530 612
rect 2942 1388 2988 1400
rect 2942 612 2948 1388
rect 2982 612 2988 1388
rect 2942 600 2988 612
rect 3400 1388 3446 1400
rect 3400 612 3406 1388
rect 3440 612 3446 1388
rect 3400 600 3446 612
rect 3858 1388 3904 1400
rect 3858 612 3864 1388
rect 3898 612 3904 1388
rect 3858 600 3904 612
rect 4316 1388 4362 1400
rect 4316 612 4322 1388
rect 4356 612 4362 1388
rect 4316 600 4362 612
rect 90 30 4368 60
rect 90 -30 358 30
rect 418 -30 758 30
rect 818 -30 1158 30
rect 1218 -30 1558 30
rect 1618 -30 1958 30
rect 2018 -30 2358 30
rect 2418 -30 2758 30
rect 2818 -30 3158 30
rect 3218 -30 3558 30
rect 3618 -30 3958 30
rect 4018 -30 4368 30
rect 90 -60 4368 -30
<< labels >>
flabel metal1 188 1850 248 1910 1 FreeSans 800 0 0 0 VPWR
port 4 n power bidirectional
flabel metal1 188 -30 248 30 1 FreeSans 800 0 0 0 VGND
port 5 n ground bidirectional
flabel locali 4308 1690 4368 1750 1 FreeSans 800 0 0 0 SOURCE
port 2 n default bidirectional
flabel locali 4308 370 4368 430 1 FreeSans 800 0 0 0 DRAIN
port 3 n default bidirectional
flabel locali 4308 144 4368 204 1 FreeSans 800 0 0 0 GATE
port 1 n default bidirectional
<< properties >>
string FIXED_BBOX 0 0 4500 1880
string LEFclass CORE
string LEFsite unitasc
<< end >>
