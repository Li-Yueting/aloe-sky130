.subckt sky130_asc_pfet_01v8_lvt_1 GATE SOURCE DRAIN VGND VPWR
X0 SOURCE GATE DRAIN VPWR sky130_fd_pr__pfet_01v8_lvt ad=1.8705e+12p pd=1.348e+07u as=1.8705e+12p ps=1.348e+07u w=6.45e+06u l=2e+06u
.ends


.subckt sky130_fd_pr__cap_mim_m3_1 c0 c1 VPWR VGND
X0 c1 c0 sky130_fd_pr__cap_mim_m3_1 l=2e+06u w=2e+06u
X1 c1 c0 sky130_fd_pr__cap_mim_m3_1 l=2e+06u w=2e+06u
X2 c1 c0 sky130_fd_pr__cap_mim_m3_1 l=2e+06u w=2e+06u
X3 c1 c0 sky130_fd_pr__cap_mim_m3_1 l=2e+06u w=2e+06u
X4 c1 c0 sky130_fd_pr__cap_mim_m3_1 l=2e+06u w=2e+06u
X5 c1 c0 sky130_fd_pr__cap_mim_m3_1 l=2e+06u w=2e+06u
X6 c1 c0 sky130_fd_pr__cap_mim_m3_1 l=2e+06u w=2e+06u
X7 c1 c0 sky130_fd_pr__cap_mim_m3_1 l=2e+06u w=2e+06u
X8 c1 c0 sky130_fd_pr__cap_mim_m3_1 l=2e+06u w=2e+06u
X9 c1 c0 sky130_fd_pr__cap_mim_m3_1 l=2e+06u w=2e+06u
X10 c1 c0 sky130_fd_pr__cap_mim_m3_1 l=2e+06u w=2e+06u
X11 c1 c0 sky130_fd_pr__cap_mim_m3_1 l=2e+06u w=2e+06u
X12 c1 c0 sky130_fd_pr__cap_mim_m3_1 l=2e+06u w=2e+06u
X13 c1 c0 sky130_fd_pr__cap_mim_m3_1 l=2e+06u w=2e+06u
X14 c1 c0 sky130_fd_pr__cap_mim_m3_1 l=2e+06u w=2e+06u
X15 c1 c0 sky130_fd_pr__cap_mim_m3_1 l=2e+06u w=2e+06u
X16 c1 c0 sky130_fd_pr__cap_mim_m3_1 l=2e+06u w=2e+06u
X17 c1 c0 sky130_fd_pr__cap_mim_m3_1 l=2e+06u w=2e+06u
X18 c1 c0 sky130_fd_pr__cap_mim_m3_1 l=2e+06u w=2e+06u
X19 c1 c0 sky130_fd_pr__cap_mim_m3_1 l=2e+06u w=2e+06u
.ends


.subckt sky130_asc_nfet_01v8_lvt_1 GATE SOURCE DRAIN VPWR VGND
X0 SOURCE GATE DRAIN VGND sky130_fd_pr__nfet_01v8_lvt ad=1.16e+12p pd=8.58e+06u as=1.16e+12p ps=8.58e+06u w=4e+06u l=2e+06u
.ends


