VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO bgr_0
  CLASS BLOCK ;
  FOREIGN bgr_0 ;
  ORIGIN 0.000 0.000 ;
  SIZE 292.560 BY 282.880 ;
  PIN porst
    ANTENNAGATEAREA 72.000000 ;
    PORT
      LAYER li1 ;
        RECT 127.490 124.080 147.990 124.380 ;
      LAYER mcon ;
        RECT 137.685 124.185 137.855 124.355 ;
      LAYER met1 ;
        RECT 137.610 124.340 137.930 124.400 ;
        RECT 137.335 124.200 137.930 124.340 ;
        RECT 137.610 124.140 137.930 124.200 ;
        RECT 127.490 22.680 127.810 22.740 ;
        RECT 137.610 22.680 137.930 22.740 ;
        RECT 127.490 22.540 137.930 22.680 ;
        RECT 127.490 22.480 127.810 22.540 ;
        RECT 137.610 22.480 137.930 22.540 ;
      LAYER via ;
        RECT 137.640 124.140 137.900 124.400 ;
        RECT 127.520 22.480 127.780 22.740 ;
        RECT 137.640 22.480 137.900 22.740 ;
      LAYER met2 ;
        RECT 137.640 124.110 137.900 124.430 ;
        RECT 137.700 22.770 137.840 124.110 ;
        RECT 127.520 22.450 127.780 22.770 ;
        RECT 137.640 22.450 137.900 22.770 ;
        RECT 127.580 0.000 127.720 22.450 ;
    END
  END porst
  PIN va
    ANTENNAGATEAREA 72.000000 ;
    ANTENNADIFFAREA 82.639000 ;
    PORT
      LAYER li1 ;
        RECT 75.385 217.910 75.555 224.805 ;
        RECT 79.965 217.910 80.135 224.805 ;
        RECT 84.545 217.910 84.715 224.805 ;
        RECT 89.125 217.910 89.295 224.805 ;
        RECT 93.705 217.910 93.875 224.805 ;
        RECT 98.285 217.910 98.455 224.805 ;
        RECT 102.865 217.910 103.035 224.805 ;
        RECT 107.445 217.910 107.615 224.805 ;
        RECT 112.025 217.910 112.195 224.805 ;
        RECT 116.605 217.910 116.775 224.805 ;
        RECT 121.185 217.910 121.355 224.805 ;
        RECT 125.765 217.910 125.935 224.805 ;
        RECT 130.345 217.910 130.515 224.805 ;
        RECT 134.925 217.910 135.095 224.805 ;
        RECT 139.505 217.910 139.675 224.805 ;
        RECT 144.085 217.910 144.255 224.805 ;
        RECT 148.665 217.910 148.835 224.805 ;
        RECT 153.245 217.910 153.415 224.805 ;
        RECT 157.825 217.910 157.995 224.805 ;
        RECT 162.405 217.910 162.575 224.805 ;
        RECT 166.985 217.910 167.155 224.805 ;
        RECT 171.565 217.910 171.735 224.805 ;
        RECT 176.145 217.910 176.315 224.805 ;
        RECT 180.725 217.910 180.895 224.805 ;
        RECT 185.305 217.910 185.475 224.805 ;
        RECT 189.885 217.910 190.055 224.805 ;
        RECT 194.465 217.910 194.635 224.805 ;
        RECT 199.045 217.910 199.215 224.805 ;
        RECT 203.625 217.910 203.795 224.805 ;
        RECT 208.205 217.910 208.375 224.805 ;
        RECT 212.785 217.910 212.955 224.805 ;
        RECT 75.150 217.855 213.190 217.910 ;
        RECT 75.125 217.685 213.190 217.855 ;
        RECT 75.150 217.610 213.190 217.685 ;
        RECT 113.605 199.155 113.775 206.005 ;
        RECT 113.605 199.110 113.935 199.155 ;
        RECT 118.185 199.110 118.355 206.005 ;
        RECT 122.765 199.110 122.935 206.005 ;
        RECT 127.345 199.110 127.515 206.005 ;
        RECT 131.925 199.110 132.095 206.005 ;
        RECT 136.505 199.110 136.675 206.005 ;
        RECT 140.445 199.110 140.615 199.155 ;
        RECT 141.085 199.110 141.255 206.005 ;
        RECT 113.370 198.810 141.490 199.110 ;
        RECT 61.575 181.925 65.045 185.395 ;
        RECT 140.445 180.780 140.615 180.795 ;
        RECT 127.490 180.480 147.990 180.780 ;
        RECT 110.040 146.735 112.200 149.585 ;
      LAYER mcon ;
        RECT 75.385 224.535 75.555 224.705 ;
        RECT 75.385 224.175 75.555 224.345 ;
        RECT 75.385 223.815 75.555 223.985 ;
        RECT 75.385 223.455 75.555 223.625 ;
        RECT 75.385 223.095 75.555 223.265 ;
        RECT 75.385 222.735 75.555 222.905 ;
        RECT 75.385 222.375 75.555 222.545 ;
        RECT 75.385 222.015 75.555 222.185 ;
        RECT 75.385 221.655 75.555 221.825 ;
        RECT 75.385 221.295 75.555 221.465 ;
        RECT 75.385 220.935 75.555 221.105 ;
        RECT 75.385 220.575 75.555 220.745 ;
        RECT 75.385 220.215 75.555 220.385 ;
        RECT 75.385 219.855 75.555 220.025 ;
        RECT 75.385 219.495 75.555 219.665 ;
        RECT 75.385 219.135 75.555 219.305 ;
        RECT 75.385 218.775 75.555 218.945 ;
        RECT 75.385 218.415 75.555 218.585 ;
        RECT 79.965 224.535 80.135 224.705 ;
        RECT 79.965 224.175 80.135 224.345 ;
        RECT 79.965 223.815 80.135 223.985 ;
        RECT 79.965 223.455 80.135 223.625 ;
        RECT 79.965 223.095 80.135 223.265 ;
        RECT 79.965 222.735 80.135 222.905 ;
        RECT 79.965 222.375 80.135 222.545 ;
        RECT 79.965 222.015 80.135 222.185 ;
        RECT 79.965 221.655 80.135 221.825 ;
        RECT 79.965 221.295 80.135 221.465 ;
        RECT 79.965 220.935 80.135 221.105 ;
        RECT 79.965 220.575 80.135 220.745 ;
        RECT 79.965 220.215 80.135 220.385 ;
        RECT 79.965 219.855 80.135 220.025 ;
        RECT 79.965 219.495 80.135 219.665 ;
        RECT 79.965 219.135 80.135 219.305 ;
        RECT 79.965 218.775 80.135 218.945 ;
        RECT 79.965 218.415 80.135 218.585 ;
        RECT 84.545 224.535 84.715 224.705 ;
        RECT 84.545 224.175 84.715 224.345 ;
        RECT 84.545 223.815 84.715 223.985 ;
        RECT 84.545 223.455 84.715 223.625 ;
        RECT 84.545 223.095 84.715 223.265 ;
        RECT 84.545 222.735 84.715 222.905 ;
        RECT 84.545 222.375 84.715 222.545 ;
        RECT 84.545 222.015 84.715 222.185 ;
        RECT 84.545 221.655 84.715 221.825 ;
        RECT 84.545 221.295 84.715 221.465 ;
        RECT 84.545 220.935 84.715 221.105 ;
        RECT 84.545 220.575 84.715 220.745 ;
        RECT 84.545 220.215 84.715 220.385 ;
        RECT 84.545 219.855 84.715 220.025 ;
        RECT 84.545 219.495 84.715 219.665 ;
        RECT 84.545 219.135 84.715 219.305 ;
        RECT 84.545 218.775 84.715 218.945 ;
        RECT 84.545 218.415 84.715 218.585 ;
        RECT 89.125 224.535 89.295 224.705 ;
        RECT 89.125 224.175 89.295 224.345 ;
        RECT 89.125 223.815 89.295 223.985 ;
        RECT 89.125 223.455 89.295 223.625 ;
        RECT 89.125 223.095 89.295 223.265 ;
        RECT 89.125 222.735 89.295 222.905 ;
        RECT 89.125 222.375 89.295 222.545 ;
        RECT 89.125 222.015 89.295 222.185 ;
        RECT 89.125 221.655 89.295 221.825 ;
        RECT 89.125 221.295 89.295 221.465 ;
        RECT 89.125 220.935 89.295 221.105 ;
        RECT 89.125 220.575 89.295 220.745 ;
        RECT 89.125 220.215 89.295 220.385 ;
        RECT 89.125 219.855 89.295 220.025 ;
        RECT 89.125 219.495 89.295 219.665 ;
        RECT 89.125 219.135 89.295 219.305 ;
        RECT 89.125 218.775 89.295 218.945 ;
        RECT 89.125 218.415 89.295 218.585 ;
        RECT 93.705 224.535 93.875 224.705 ;
        RECT 93.705 224.175 93.875 224.345 ;
        RECT 93.705 223.815 93.875 223.985 ;
        RECT 93.705 223.455 93.875 223.625 ;
        RECT 93.705 223.095 93.875 223.265 ;
        RECT 93.705 222.735 93.875 222.905 ;
        RECT 93.705 222.375 93.875 222.545 ;
        RECT 93.705 222.015 93.875 222.185 ;
        RECT 93.705 221.655 93.875 221.825 ;
        RECT 93.705 221.295 93.875 221.465 ;
        RECT 93.705 220.935 93.875 221.105 ;
        RECT 93.705 220.575 93.875 220.745 ;
        RECT 93.705 220.215 93.875 220.385 ;
        RECT 93.705 219.855 93.875 220.025 ;
        RECT 93.705 219.495 93.875 219.665 ;
        RECT 93.705 219.135 93.875 219.305 ;
        RECT 93.705 218.775 93.875 218.945 ;
        RECT 93.705 218.415 93.875 218.585 ;
        RECT 98.285 224.535 98.455 224.705 ;
        RECT 98.285 224.175 98.455 224.345 ;
        RECT 98.285 223.815 98.455 223.985 ;
        RECT 98.285 223.455 98.455 223.625 ;
        RECT 98.285 223.095 98.455 223.265 ;
        RECT 98.285 222.735 98.455 222.905 ;
        RECT 98.285 222.375 98.455 222.545 ;
        RECT 98.285 222.015 98.455 222.185 ;
        RECT 98.285 221.655 98.455 221.825 ;
        RECT 98.285 221.295 98.455 221.465 ;
        RECT 98.285 220.935 98.455 221.105 ;
        RECT 98.285 220.575 98.455 220.745 ;
        RECT 98.285 220.215 98.455 220.385 ;
        RECT 98.285 219.855 98.455 220.025 ;
        RECT 98.285 219.495 98.455 219.665 ;
        RECT 98.285 219.135 98.455 219.305 ;
        RECT 98.285 218.775 98.455 218.945 ;
        RECT 98.285 218.415 98.455 218.585 ;
        RECT 102.865 224.535 103.035 224.705 ;
        RECT 102.865 224.175 103.035 224.345 ;
        RECT 102.865 223.815 103.035 223.985 ;
        RECT 102.865 223.455 103.035 223.625 ;
        RECT 102.865 223.095 103.035 223.265 ;
        RECT 102.865 222.735 103.035 222.905 ;
        RECT 102.865 222.375 103.035 222.545 ;
        RECT 102.865 222.015 103.035 222.185 ;
        RECT 102.865 221.655 103.035 221.825 ;
        RECT 102.865 221.295 103.035 221.465 ;
        RECT 102.865 220.935 103.035 221.105 ;
        RECT 102.865 220.575 103.035 220.745 ;
        RECT 102.865 220.215 103.035 220.385 ;
        RECT 102.865 219.855 103.035 220.025 ;
        RECT 102.865 219.495 103.035 219.665 ;
        RECT 102.865 219.135 103.035 219.305 ;
        RECT 102.865 218.775 103.035 218.945 ;
        RECT 102.865 218.415 103.035 218.585 ;
        RECT 107.445 224.535 107.615 224.705 ;
        RECT 107.445 224.175 107.615 224.345 ;
        RECT 107.445 223.815 107.615 223.985 ;
        RECT 107.445 223.455 107.615 223.625 ;
        RECT 107.445 223.095 107.615 223.265 ;
        RECT 107.445 222.735 107.615 222.905 ;
        RECT 107.445 222.375 107.615 222.545 ;
        RECT 107.445 222.015 107.615 222.185 ;
        RECT 107.445 221.655 107.615 221.825 ;
        RECT 107.445 221.295 107.615 221.465 ;
        RECT 107.445 220.935 107.615 221.105 ;
        RECT 107.445 220.575 107.615 220.745 ;
        RECT 107.445 220.215 107.615 220.385 ;
        RECT 107.445 219.855 107.615 220.025 ;
        RECT 107.445 219.495 107.615 219.665 ;
        RECT 107.445 219.135 107.615 219.305 ;
        RECT 107.445 218.775 107.615 218.945 ;
        RECT 107.445 218.415 107.615 218.585 ;
        RECT 112.025 224.535 112.195 224.705 ;
        RECT 112.025 224.175 112.195 224.345 ;
        RECT 112.025 223.815 112.195 223.985 ;
        RECT 112.025 223.455 112.195 223.625 ;
        RECT 112.025 223.095 112.195 223.265 ;
        RECT 112.025 222.735 112.195 222.905 ;
        RECT 112.025 222.375 112.195 222.545 ;
        RECT 112.025 222.015 112.195 222.185 ;
        RECT 112.025 221.655 112.195 221.825 ;
        RECT 112.025 221.295 112.195 221.465 ;
        RECT 112.025 220.935 112.195 221.105 ;
        RECT 112.025 220.575 112.195 220.745 ;
        RECT 112.025 220.215 112.195 220.385 ;
        RECT 112.025 219.855 112.195 220.025 ;
        RECT 112.025 219.495 112.195 219.665 ;
        RECT 112.025 219.135 112.195 219.305 ;
        RECT 112.025 218.775 112.195 218.945 ;
        RECT 112.025 218.415 112.195 218.585 ;
        RECT 116.605 224.535 116.775 224.705 ;
        RECT 116.605 224.175 116.775 224.345 ;
        RECT 116.605 223.815 116.775 223.985 ;
        RECT 116.605 223.455 116.775 223.625 ;
        RECT 116.605 223.095 116.775 223.265 ;
        RECT 116.605 222.735 116.775 222.905 ;
        RECT 116.605 222.375 116.775 222.545 ;
        RECT 116.605 222.015 116.775 222.185 ;
        RECT 116.605 221.655 116.775 221.825 ;
        RECT 116.605 221.295 116.775 221.465 ;
        RECT 116.605 220.935 116.775 221.105 ;
        RECT 116.605 220.575 116.775 220.745 ;
        RECT 116.605 220.215 116.775 220.385 ;
        RECT 116.605 219.855 116.775 220.025 ;
        RECT 116.605 219.495 116.775 219.665 ;
        RECT 116.605 219.135 116.775 219.305 ;
        RECT 116.605 218.775 116.775 218.945 ;
        RECT 116.605 218.415 116.775 218.585 ;
        RECT 121.185 224.535 121.355 224.705 ;
        RECT 121.185 224.175 121.355 224.345 ;
        RECT 121.185 223.815 121.355 223.985 ;
        RECT 121.185 223.455 121.355 223.625 ;
        RECT 121.185 223.095 121.355 223.265 ;
        RECT 121.185 222.735 121.355 222.905 ;
        RECT 121.185 222.375 121.355 222.545 ;
        RECT 121.185 222.015 121.355 222.185 ;
        RECT 121.185 221.655 121.355 221.825 ;
        RECT 121.185 221.295 121.355 221.465 ;
        RECT 121.185 220.935 121.355 221.105 ;
        RECT 121.185 220.575 121.355 220.745 ;
        RECT 121.185 220.215 121.355 220.385 ;
        RECT 121.185 219.855 121.355 220.025 ;
        RECT 121.185 219.495 121.355 219.665 ;
        RECT 121.185 219.135 121.355 219.305 ;
        RECT 121.185 218.775 121.355 218.945 ;
        RECT 121.185 218.415 121.355 218.585 ;
        RECT 125.765 224.535 125.935 224.705 ;
        RECT 125.765 224.175 125.935 224.345 ;
        RECT 125.765 223.815 125.935 223.985 ;
        RECT 125.765 223.455 125.935 223.625 ;
        RECT 125.765 223.095 125.935 223.265 ;
        RECT 125.765 222.735 125.935 222.905 ;
        RECT 125.765 222.375 125.935 222.545 ;
        RECT 125.765 222.015 125.935 222.185 ;
        RECT 125.765 221.655 125.935 221.825 ;
        RECT 125.765 221.295 125.935 221.465 ;
        RECT 125.765 220.935 125.935 221.105 ;
        RECT 125.765 220.575 125.935 220.745 ;
        RECT 125.765 220.215 125.935 220.385 ;
        RECT 125.765 219.855 125.935 220.025 ;
        RECT 125.765 219.495 125.935 219.665 ;
        RECT 125.765 219.135 125.935 219.305 ;
        RECT 125.765 218.775 125.935 218.945 ;
        RECT 125.765 218.415 125.935 218.585 ;
        RECT 130.345 224.535 130.515 224.705 ;
        RECT 130.345 224.175 130.515 224.345 ;
        RECT 130.345 223.815 130.515 223.985 ;
        RECT 130.345 223.455 130.515 223.625 ;
        RECT 130.345 223.095 130.515 223.265 ;
        RECT 130.345 222.735 130.515 222.905 ;
        RECT 130.345 222.375 130.515 222.545 ;
        RECT 130.345 222.015 130.515 222.185 ;
        RECT 130.345 221.655 130.515 221.825 ;
        RECT 130.345 221.295 130.515 221.465 ;
        RECT 130.345 220.935 130.515 221.105 ;
        RECT 130.345 220.575 130.515 220.745 ;
        RECT 130.345 220.215 130.515 220.385 ;
        RECT 130.345 219.855 130.515 220.025 ;
        RECT 130.345 219.495 130.515 219.665 ;
        RECT 130.345 219.135 130.515 219.305 ;
        RECT 130.345 218.775 130.515 218.945 ;
        RECT 130.345 218.415 130.515 218.585 ;
        RECT 134.925 224.535 135.095 224.705 ;
        RECT 134.925 224.175 135.095 224.345 ;
        RECT 134.925 223.815 135.095 223.985 ;
        RECT 134.925 223.455 135.095 223.625 ;
        RECT 134.925 223.095 135.095 223.265 ;
        RECT 134.925 222.735 135.095 222.905 ;
        RECT 134.925 222.375 135.095 222.545 ;
        RECT 134.925 222.015 135.095 222.185 ;
        RECT 134.925 221.655 135.095 221.825 ;
        RECT 134.925 221.295 135.095 221.465 ;
        RECT 134.925 220.935 135.095 221.105 ;
        RECT 134.925 220.575 135.095 220.745 ;
        RECT 134.925 220.215 135.095 220.385 ;
        RECT 134.925 219.855 135.095 220.025 ;
        RECT 134.925 219.495 135.095 219.665 ;
        RECT 134.925 219.135 135.095 219.305 ;
        RECT 134.925 218.775 135.095 218.945 ;
        RECT 134.925 218.415 135.095 218.585 ;
        RECT 139.505 224.535 139.675 224.705 ;
        RECT 139.505 224.175 139.675 224.345 ;
        RECT 139.505 223.815 139.675 223.985 ;
        RECT 139.505 223.455 139.675 223.625 ;
        RECT 139.505 223.095 139.675 223.265 ;
        RECT 139.505 222.735 139.675 222.905 ;
        RECT 139.505 222.375 139.675 222.545 ;
        RECT 139.505 222.015 139.675 222.185 ;
        RECT 139.505 221.655 139.675 221.825 ;
        RECT 139.505 221.295 139.675 221.465 ;
        RECT 139.505 220.935 139.675 221.105 ;
        RECT 139.505 220.575 139.675 220.745 ;
        RECT 139.505 220.215 139.675 220.385 ;
        RECT 139.505 219.855 139.675 220.025 ;
        RECT 139.505 219.495 139.675 219.665 ;
        RECT 139.505 219.135 139.675 219.305 ;
        RECT 139.505 218.775 139.675 218.945 ;
        RECT 139.505 218.415 139.675 218.585 ;
        RECT 144.085 224.535 144.255 224.705 ;
        RECT 144.085 224.175 144.255 224.345 ;
        RECT 144.085 223.815 144.255 223.985 ;
        RECT 144.085 223.455 144.255 223.625 ;
        RECT 144.085 223.095 144.255 223.265 ;
        RECT 144.085 222.735 144.255 222.905 ;
        RECT 144.085 222.375 144.255 222.545 ;
        RECT 144.085 222.015 144.255 222.185 ;
        RECT 144.085 221.655 144.255 221.825 ;
        RECT 144.085 221.295 144.255 221.465 ;
        RECT 144.085 220.935 144.255 221.105 ;
        RECT 144.085 220.575 144.255 220.745 ;
        RECT 144.085 220.215 144.255 220.385 ;
        RECT 144.085 219.855 144.255 220.025 ;
        RECT 144.085 219.495 144.255 219.665 ;
        RECT 144.085 219.135 144.255 219.305 ;
        RECT 144.085 218.775 144.255 218.945 ;
        RECT 144.085 218.415 144.255 218.585 ;
        RECT 148.665 224.535 148.835 224.705 ;
        RECT 148.665 224.175 148.835 224.345 ;
        RECT 148.665 223.815 148.835 223.985 ;
        RECT 148.665 223.455 148.835 223.625 ;
        RECT 148.665 223.095 148.835 223.265 ;
        RECT 148.665 222.735 148.835 222.905 ;
        RECT 148.665 222.375 148.835 222.545 ;
        RECT 148.665 222.015 148.835 222.185 ;
        RECT 148.665 221.655 148.835 221.825 ;
        RECT 148.665 221.295 148.835 221.465 ;
        RECT 148.665 220.935 148.835 221.105 ;
        RECT 148.665 220.575 148.835 220.745 ;
        RECT 148.665 220.215 148.835 220.385 ;
        RECT 148.665 219.855 148.835 220.025 ;
        RECT 148.665 219.495 148.835 219.665 ;
        RECT 148.665 219.135 148.835 219.305 ;
        RECT 148.665 218.775 148.835 218.945 ;
        RECT 148.665 218.415 148.835 218.585 ;
        RECT 153.245 224.535 153.415 224.705 ;
        RECT 153.245 224.175 153.415 224.345 ;
        RECT 153.245 223.815 153.415 223.985 ;
        RECT 153.245 223.455 153.415 223.625 ;
        RECT 153.245 223.095 153.415 223.265 ;
        RECT 153.245 222.735 153.415 222.905 ;
        RECT 153.245 222.375 153.415 222.545 ;
        RECT 153.245 222.015 153.415 222.185 ;
        RECT 153.245 221.655 153.415 221.825 ;
        RECT 153.245 221.295 153.415 221.465 ;
        RECT 153.245 220.935 153.415 221.105 ;
        RECT 153.245 220.575 153.415 220.745 ;
        RECT 153.245 220.215 153.415 220.385 ;
        RECT 153.245 219.855 153.415 220.025 ;
        RECT 153.245 219.495 153.415 219.665 ;
        RECT 153.245 219.135 153.415 219.305 ;
        RECT 153.245 218.775 153.415 218.945 ;
        RECT 153.245 218.415 153.415 218.585 ;
        RECT 157.825 224.535 157.995 224.705 ;
        RECT 157.825 224.175 157.995 224.345 ;
        RECT 157.825 223.815 157.995 223.985 ;
        RECT 157.825 223.455 157.995 223.625 ;
        RECT 157.825 223.095 157.995 223.265 ;
        RECT 157.825 222.735 157.995 222.905 ;
        RECT 157.825 222.375 157.995 222.545 ;
        RECT 157.825 222.015 157.995 222.185 ;
        RECT 157.825 221.655 157.995 221.825 ;
        RECT 157.825 221.295 157.995 221.465 ;
        RECT 157.825 220.935 157.995 221.105 ;
        RECT 157.825 220.575 157.995 220.745 ;
        RECT 157.825 220.215 157.995 220.385 ;
        RECT 157.825 219.855 157.995 220.025 ;
        RECT 157.825 219.495 157.995 219.665 ;
        RECT 157.825 219.135 157.995 219.305 ;
        RECT 157.825 218.775 157.995 218.945 ;
        RECT 157.825 218.415 157.995 218.585 ;
        RECT 162.405 224.535 162.575 224.705 ;
        RECT 162.405 224.175 162.575 224.345 ;
        RECT 162.405 223.815 162.575 223.985 ;
        RECT 162.405 223.455 162.575 223.625 ;
        RECT 162.405 223.095 162.575 223.265 ;
        RECT 162.405 222.735 162.575 222.905 ;
        RECT 162.405 222.375 162.575 222.545 ;
        RECT 162.405 222.015 162.575 222.185 ;
        RECT 162.405 221.655 162.575 221.825 ;
        RECT 162.405 221.295 162.575 221.465 ;
        RECT 162.405 220.935 162.575 221.105 ;
        RECT 162.405 220.575 162.575 220.745 ;
        RECT 162.405 220.215 162.575 220.385 ;
        RECT 162.405 219.855 162.575 220.025 ;
        RECT 162.405 219.495 162.575 219.665 ;
        RECT 162.405 219.135 162.575 219.305 ;
        RECT 162.405 218.775 162.575 218.945 ;
        RECT 162.405 218.415 162.575 218.585 ;
        RECT 166.985 224.535 167.155 224.705 ;
        RECT 166.985 224.175 167.155 224.345 ;
        RECT 166.985 223.815 167.155 223.985 ;
        RECT 166.985 223.455 167.155 223.625 ;
        RECT 166.985 223.095 167.155 223.265 ;
        RECT 166.985 222.735 167.155 222.905 ;
        RECT 166.985 222.375 167.155 222.545 ;
        RECT 166.985 222.015 167.155 222.185 ;
        RECT 166.985 221.655 167.155 221.825 ;
        RECT 166.985 221.295 167.155 221.465 ;
        RECT 166.985 220.935 167.155 221.105 ;
        RECT 166.985 220.575 167.155 220.745 ;
        RECT 166.985 220.215 167.155 220.385 ;
        RECT 166.985 219.855 167.155 220.025 ;
        RECT 166.985 219.495 167.155 219.665 ;
        RECT 166.985 219.135 167.155 219.305 ;
        RECT 166.985 218.775 167.155 218.945 ;
        RECT 166.985 218.415 167.155 218.585 ;
        RECT 171.565 224.535 171.735 224.705 ;
        RECT 171.565 224.175 171.735 224.345 ;
        RECT 171.565 223.815 171.735 223.985 ;
        RECT 171.565 223.455 171.735 223.625 ;
        RECT 171.565 223.095 171.735 223.265 ;
        RECT 171.565 222.735 171.735 222.905 ;
        RECT 171.565 222.375 171.735 222.545 ;
        RECT 171.565 222.015 171.735 222.185 ;
        RECT 171.565 221.655 171.735 221.825 ;
        RECT 171.565 221.295 171.735 221.465 ;
        RECT 171.565 220.935 171.735 221.105 ;
        RECT 171.565 220.575 171.735 220.745 ;
        RECT 171.565 220.215 171.735 220.385 ;
        RECT 171.565 219.855 171.735 220.025 ;
        RECT 171.565 219.495 171.735 219.665 ;
        RECT 171.565 219.135 171.735 219.305 ;
        RECT 171.565 218.775 171.735 218.945 ;
        RECT 171.565 218.415 171.735 218.585 ;
        RECT 176.145 224.535 176.315 224.705 ;
        RECT 176.145 224.175 176.315 224.345 ;
        RECT 176.145 223.815 176.315 223.985 ;
        RECT 176.145 223.455 176.315 223.625 ;
        RECT 176.145 223.095 176.315 223.265 ;
        RECT 176.145 222.735 176.315 222.905 ;
        RECT 176.145 222.375 176.315 222.545 ;
        RECT 176.145 222.015 176.315 222.185 ;
        RECT 176.145 221.655 176.315 221.825 ;
        RECT 176.145 221.295 176.315 221.465 ;
        RECT 176.145 220.935 176.315 221.105 ;
        RECT 176.145 220.575 176.315 220.745 ;
        RECT 176.145 220.215 176.315 220.385 ;
        RECT 176.145 219.855 176.315 220.025 ;
        RECT 176.145 219.495 176.315 219.665 ;
        RECT 176.145 219.135 176.315 219.305 ;
        RECT 176.145 218.775 176.315 218.945 ;
        RECT 176.145 218.415 176.315 218.585 ;
        RECT 180.725 224.535 180.895 224.705 ;
        RECT 180.725 224.175 180.895 224.345 ;
        RECT 180.725 223.815 180.895 223.985 ;
        RECT 180.725 223.455 180.895 223.625 ;
        RECT 180.725 223.095 180.895 223.265 ;
        RECT 180.725 222.735 180.895 222.905 ;
        RECT 180.725 222.375 180.895 222.545 ;
        RECT 180.725 222.015 180.895 222.185 ;
        RECT 180.725 221.655 180.895 221.825 ;
        RECT 180.725 221.295 180.895 221.465 ;
        RECT 180.725 220.935 180.895 221.105 ;
        RECT 180.725 220.575 180.895 220.745 ;
        RECT 180.725 220.215 180.895 220.385 ;
        RECT 180.725 219.855 180.895 220.025 ;
        RECT 180.725 219.495 180.895 219.665 ;
        RECT 180.725 219.135 180.895 219.305 ;
        RECT 180.725 218.775 180.895 218.945 ;
        RECT 180.725 218.415 180.895 218.585 ;
        RECT 185.305 224.535 185.475 224.705 ;
        RECT 185.305 224.175 185.475 224.345 ;
        RECT 185.305 223.815 185.475 223.985 ;
        RECT 185.305 223.455 185.475 223.625 ;
        RECT 185.305 223.095 185.475 223.265 ;
        RECT 185.305 222.735 185.475 222.905 ;
        RECT 185.305 222.375 185.475 222.545 ;
        RECT 185.305 222.015 185.475 222.185 ;
        RECT 185.305 221.655 185.475 221.825 ;
        RECT 185.305 221.295 185.475 221.465 ;
        RECT 185.305 220.935 185.475 221.105 ;
        RECT 185.305 220.575 185.475 220.745 ;
        RECT 185.305 220.215 185.475 220.385 ;
        RECT 185.305 219.855 185.475 220.025 ;
        RECT 185.305 219.495 185.475 219.665 ;
        RECT 185.305 219.135 185.475 219.305 ;
        RECT 185.305 218.775 185.475 218.945 ;
        RECT 185.305 218.415 185.475 218.585 ;
        RECT 189.885 224.535 190.055 224.705 ;
        RECT 189.885 224.175 190.055 224.345 ;
        RECT 189.885 223.815 190.055 223.985 ;
        RECT 189.885 223.455 190.055 223.625 ;
        RECT 189.885 223.095 190.055 223.265 ;
        RECT 189.885 222.735 190.055 222.905 ;
        RECT 189.885 222.375 190.055 222.545 ;
        RECT 189.885 222.015 190.055 222.185 ;
        RECT 189.885 221.655 190.055 221.825 ;
        RECT 189.885 221.295 190.055 221.465 ;
        RECT 189.885 220.935 190.055 221.105 ;
        RECT 189.885 220.575 190.055 220.745 ;
        RECT 189.885 220.215 190.055 220.385 ;
        RECT 189.885 219.855 190.055 220.025 ;
        RECT 189.885 219.495 190.055 219.665 ;
        RECT 189.885 219.135 190.055 219.305 ;
        RECT 189.885 218.775 190.055 218.945 ;
        RECT 189.885 218.415 190.055 218.585 ;
        RECT 194.465 224.535 194.635 224.705 ;
        RECT 194.465 224.175 194.635 224.345 ;
        RECT 194.465 223.815 194.635 223.985 ;
        RECT 194.465 223.455 194.635 223.625 ;
        RECT 194.465 223.095 194.635 223.265 ;
        RECT 194.465 222.735 194.635 222.905 ;
        RECT 194.465 222.375 194.635 222.545 ;
        RECT 194.465 222.015 194.635 222.185 ;
        RECT 194.465 221.655 194.635 221.825 ;
        RECT 194.465 221.295 194.635 221.465 ;
        RECT 194.465 220.935 194.635 221.105 ;
        RECT 194.465 220.575 194.635 220.745 ;
        RECT 194.465 220.215 194.635 220.385 ;
        RECT 194.465 219.855 194.635 220.025 ;
        RECT 194.465 219.495 194.635 219.665 ;
        RECT 194.465 219.135 194.635 219.305 ;
        RECT 194.465 218.775 194.635 218.945 ;
        RECT 194.465 218.415 194.635 218.585 ;
        RECT 199.045 224.535 199.215 224.705 ;
        RECT 199.045 224.175 199.215 224.345 ;
        RECT 199.045 223.815 199.215 223.985 ;
        RECT 199.045 223.455 199.215 223.625 ;
        RECT 199.045 223.095 199.215 223.265 ;
        RECT 199.045 222.735 199.215 222.905 ;
        RECT 199.045 222.375 199.215 222.545 ;
        RECT 199.045 222.015 199.215 222.185 ;
        RECT 199.045 221.655 199.215 221.825 ;
        RECT 199.045 221.295 199.215 221.465 ;
        RECT 199.045 220.935 199.215 221.105 ;
        RECT 199.045 220.575 199.215 220.745 ;
        RECT 199.045 220.215 199.215 220.385 ;
        RECT 199.045 219.855 199.215 220.025 ;
        RECT 199.045 219.495 199.215 219.665 ;
        RECT 199.045 219.135 199.215 219.305 ;
        RECT 199.045 218.775 199.215 218.945 ;
        RECT 199.045 218.415 199.215 218.585 ;
        RECT 203.625 224.535 203.795 224.705 ;
        RECT 203.625 224.175 203.795 224.345 ;
        RECT 203.625 223.815 203.795 223.985 ;
        RECT 203.625 223.455 203.795 223.625 ;
        RECT 203.625 223.095 203.795 223.265 ;
        RECT 203.625 222.735 203.795 222.905 ;
        RECT 203.625 222.375 203.795 222.545 ;
        RECT 203.625 222.015 203.795 222.185 ;
        RECT 203.625 221.655 203.795 221.825 ;
        RECT 203.625 221.295 203.795 221.465 ;
        RECT 203.625 220.935 203.795 221.105 ;
        RECT 203.625 220.575 203.795 220.745 ;
        RECT 203.625 220.215 203.795 220.385 ;
        RECT 203.625 219.855 203.795 220.025 ;
        RECT 203.625 219.495 203.795 219.665 ;
        RECT 203.625 219.135 203.795 219.305 ;
        RECT 203.625 218.775 203.795 218.945 ;
        RECT 203.625 218.415 203.795 218.585 ;
        RECT 208.205 224.535 208.375 224.705 ;
        RECT 208.205 224.175 208.375 224.345 ;
        RECT 208.205 223.815 208.375 223.985 ;
        RECT 208.205 223.455 208.375 223.625 ;
        RECT 208.205 223.095 208.375 223.265 ;
        RECT 208.205 222.735 208.375 222.905 ;
        RECT 208.205 222.375 208.375 222.545 ;
        RECT 208.205 222.015 208.375 222.185 ;
        RECT 208.205 221.655 208.375 221.825 ;
        RECT 208.205 221.295 208.375 221.465 ;
        RECT 208.205 220.935 208.375 221.105 ;
        RECT 208.205 220.575 208.375 220.745 ;
        RECT 208.205 220.215 208.375 220.385 ;
        RECT 208.205 219.855 208.375 220.025 ;
        RECT 208.205 219.495 208.375 219.665 ;
        RECT 208.205 219.135 208.375 219.305 ;
        RECT 208.205 218.775 208.375 218.945 ;
        RECT 208.205 218.415 208.375 218.585 ;
        RECT 212.785 224.535 212.955 224.705 ;
        RECT 212.785 224.175 212.955 224.345 ;
        RECT 212.785 223.815 212.955 223.985 ;
        RECT 212.785 223.455 212.955 223.625 ;
        RECT 212.785 223.095 212.955 223.265 ;
        RECT 212.785 222.735 212.955 222.905 ;
        RECT 212.785 222.375 212.955 222.545 ;
        RECT 212.785 222.015 212.955 222.185 ;
        RECT 212.785 221.655 212.955 221.825 ;
        RECT 212.785 221.295 212.955 221.465 ;
        RECT 212.785 220.935 212.955 221.105 ;
        RECT 212.785 220.575 212.955 220.745 ;
        RECT 212.785 220.215 212.955 220.385 ;
        RECT 212.785 219.855 212.955 220.025 ;
        RECT 212.785 219.495 212.955 219.665 ;
        RECT 212.785 219.135 212.955 219.305 ;
        RECT 212.785 218.775 212.955 218.945 ;
        RECT 212.785 218.415 212.955 218.585 ;
        RECT 113.605 205.735 113.775 205.905 ;
        RECT 113.605 205.375 113.775 205.545 ;
        RECT 113.605 205.015 113.775 205.185 ;
        RECT 113.605 204.655 113.775 204.825 ;
        RECT 113.605 204.295 113.775 204.465 ;
        RECT 113.605 203.935 113.775 204.105 ;
        RECT 113.605 203.575 113.775 203.745 ;
        RECT 113.605 203.215 113.775 203.385 ;
        RECT 113.605 202.855 113.775 203.025 ;
        RECT 113.605 202.495 113.775 202.665 ;
        RECT 113.605 202.135 113.775 202.305 ;
        RECT 113.605 201.775 113.775 201.945 ;
        RECT 113.605 201.415 113.775 201.585 ;
        RECT 113.605 201.055 113.775 201.225 ;
        RECT 113.605 200.695 113.775 200.865 ;
        RECT 113.605 200.335 113.775 200.505 ;
        RECT 113.605 199.975 113.775 200.145 ;
        RECT 113.605 199.615 113.775 199.785 ;
        RECT 118.185 205.735 118.355 205.905 ;
        RECT 118.185 205.375 118.355 205.545 ;
        RECT 118.185 205.015 118.355 205.185 ;
        RECT 118.185 204.655 118.355 204.825 ;
        RECT 118.185 204.295 118.355 204.465 ;
        RECT 118.185 203.935 118.355 204.105 ;
        RECT 118.185 203.575 118.355 203.745 ;
        RECT 118.185 203.215 118.355 203.385 ;
        RECT 118.185 202.855 118.355 203.025 ;
        RECT 118.185 202.495 118.355 202.665 ;
        RECT 118.185 202.135 118.355 202.305 ;
        RECT 118.185 201.775 118.355 201.945 ;
        RECT 118.185 201.415 118.355 201.585 ;
        RECT 118.185 201.055 118.355 201.225 ;
        RECT 118.185 200.695 118.355 200.865 ;
        RECT 118.185 200.335 118.355 200.505 ;
        RECT 118.185 199.975 118.355 200.145 ;
        RECT 118.185 199.615 118.355 199.785 ;
        RECT 113.765 198.985 113.935 199.155 ;
        RECT 122.765 205.735 122.935 205.905 ;
        RECT 122.765 205.375 122.935 205.545 ;
        RECT 122.765 205.015 122.935 205.185 ;
        RECT 122.765 204.655 122.935 204.825 ;
        RECT 122.765 204.295 122.935 204.465 ;
        RECT 122.765 203.935 122.935 204.105 ;
        RECT 122.765 203.575 122.935 203.745 ;
        RECT 122.765 203.215 122.935 203.385 ;
        RECT 122.765 202.855 122.935 203.025 ;
        RECT 122.765 202.495 122.935 202.665 ;
        RECT 122.765 202.135 122.935 202.305 ;
        RECT 122.765 201.775 122.935 201.945 ;
        RECT 122.765 201.415 122.935 201.585 ;
        RECT 122.765 201.055 122.935 201.225 ;
        RECT 122.765 200.695 122.935 200.865 ;
        RECT 122.765 200.335 122.935 200.505 ;
        RECT 122.765 199.975 122.935 200.145 ;
        RECT 122.765 199.615 122.935 199.785 ;
        RECT 127.345 205.735 127.515 205.905 ;
        RECT 127.345 205.375 127.515 205.545 ;
        RECT 127.345 205.015 127.515 205.185 ;
        RECT 127.345 204.655 127.515 204.825 ;
        RECT 127.345 204.295 127.515 204.465 ;
        RECT 127.345 203.935 127.515 204.105 ;
        RECT 127.345 203.575 127.515 203.745 ;
        RECT 127.345 203.215 127.515 203.385 ;
        RECT 127.345 202.855 127.515 203.025 ;
        RECT 127.345 202.495 127.515 202.665 ;
        RECT 127.345 202.135 127.515 202.305 ;
        RECT 127.345 201.775 127.515 201.945 ;
        RECT 127.345 201.415 127.515 201.585 ;
        RECT 127.345 201.055 127.515 201.225 ;
        RECT 127.345 200.695 127.515 200.865 ;
        RECT 127.345 200.335 127.515 200.505 ;
        RECT 127.345 199.975 127.515 200.145 ;
        RECT 127.345 199.615 127.515 199.785 ;
        RECT 131.925 205.735 132.095 205.905 ;
        RECT 131.925 205.375 132.095 205.545 ;
        RECT 131.925 205.015 132.095 205.185 ;
        RECT 131.925 204.655 132.095 204.825 ;
        RECT 131.925 204.295 132.095 204.465 ;
        RECT 131.925 203.935 132.095 204.105 ;
        RECT 131.925 203.575 132.095 203.745 ;
        RECT 131.925 203.215 132.095 203.385 ;
        RECT 131.925 202.855 132.095 203.025 ;
        RECT 131.925 202.495 132.095 202.665 ;
        RECT 131.925 202.135 132.095 202.305 ;
        RECT 131.925 201.775 132.095 201.945 ;
        RECT 131.925 201.415 132.095 201.585 ;
        RECT 131.925 201.055 132.095 201.225 ;
        RECT 131.925 200.695 132.095 200.865 ;
        RECT 131.925 200.335 132.095 200.505 ;
        RECT 131.925 199.975 132.095 200.145 ;
        RECT 131.925 199.615 132.095 199.785 ;
        RECT 136.505 205.735 136.675 205.905 ;
        RECT 136.505 205.375 136.675 205.545 ;
        RECT 136.505 205.015 136.675 205.185 ;
        RECT 136.505 204.655 136.675 204.825 ;
        RECT 136.505 204.295 136.675 204.465 ;
        RECT 136.505 203.935 136.675 204.105 ;
        RECT 136.505 203.575 136.675 203.745 ;
        RECT 136.505 203.215 136.675 203.385 ;
        RECT 136.505 202.855 136.675 203.025 ;
        RECT 136.505 202.495 136.675 202.665 ;
        RECT 136.505 202.135 136.675 202.305 ;
        RECT 136.505 201.775 136.675 201.945 ;
        RECT 136.505 201.415 136.675 201.585 ;
        RECT 136.505 201.055 136.675 201.225 ;
        RECT 136.505 200.695 136.675 200.865 ;
        RECT 136.505 200.335 136.675 200.505 ;
        RECT 136.505 199.975 136.675 200.145 ;
        RECT 136.505 199.615 136.675 199.785 ;
        RECT 141.085 205.735 141.255 205.905 ;
        RECT 141.085 205.375 141.255 205.545 ;
        RECT 141.085 205.015 141.255 205.185 ;
        RECT 141.085 204.655 141.255 204.825 ;
        RECT 141.085 204.295 141.255 204.465 ;
        RECT 141.085 203.935 141.255 204.105 ;
        RECT 141.085 203.575 141.255 203.745 ;
        RECT 141.085 203.215 141.255 203.385 ;
        RECT 141.085 202.855 141.255 203.025 ;
        RECT 141.085 202.495 141.255 202.665 ;
        RECT 141.085 202.135 141.255 202.305 ;
        RECT 141.085 201.775 141.255 201.945 ;
        RECT 141.085 201.415 141.255 201.585 ;
        RECT 141.085 201.055 141.255 201.225 ;
        RECT 141.085 200.695 141.255 200.865 ;
        RECT 141.085 200.335 141.255 200.505 ;
        RECT 141.085 199.975 141.255 200.145 ;
        RECT 141.085 199.615 141.255 199.785 ;
        RECT 140.445 198.985 140.615 199.155 ;
        RECT 61.940 184.790 62.110 184.960 ;
        RECT 62.440 184.790 62.610 184.960 ;
        RECT 62.940 184.790 63.110 184.960 ;
        RECT 63.440 184.790 63.610 184.960 ;
        RECT 63.940 184.790 64.110 184.960 ;
        RECT 64.440 184.790 64.610 184.960 ;
        RECT 61.940 184.290 62.110 184.460 ;
        RECT 62.440 184.290 62.610 184.460 ;
        RECT 62.940 184.290 63.110 184.460 ;
        RECT 63.440 184.290 63.610 184.460 ;
        RECT 63.940 184.290 64.110 184.460 ;
        RECT 64.440 184.290 64.610 184.460 ;
        RECT 61.940 183.790 62.110 183.960 ;
        RECT 62.440 183.790 62.610 183.960 ;
        RECT 62.940 183.790 63.110 183.960 ;
        RECT 63.440 183.790 63.610 183.960 ;
        RECT 63.940 183.790 64.110 183.960 ;
        RECT 64.440 183.790 64.610 183.960 ;
        RECT 61.940 183.290 62.110 183.460 ;
        RECT 62.440 183.290 62.610 183.460 ;
        RECT 62.940 183.290 63.110 183.460 ;
        RECT 63.440 183.290 63.610 183.460 ;
        RECT 63.940 183.290 64.110 183.460 ;
        RECT 64.440 183.290 64.610 183.460 ;
        RECT 61.940 182.790 62.110 182.960 ;
        RECT 62.440 182.790 62.610 182.960 ;
        RECT 62.940 182.790 63.110 182.960 ;
        RECT 63.440 182.790 63.610 182.960 ;
        RECT 63.940 182.790 64.110 182.960 ;
        RECT 64.440 182.790 64.610 182.960 ;
        RECT 61.940 182.290 62.110 182.460 ;
        RECT 62.440 182.290 62.610 182.460 ;
        RECT 62.940 182.290 63.110 182.460 ;
        RECT 63.440 182.290 63.610 182.460 ;
        RECT 63.940 182.290 64.110 182.460 ;
        RECT 64.440 182.290 64.610 182.460 ;
        RECT 140.445 180.625 140.615 180.795 ;
        RECT 110.135 146.815 112.105 149.505 ;
      LAYER met1 ;
        RECT 75.355 218.335 75.585 224.785 ;
        RECT 79.935 218.335 80.165 224.785 ;
        RECT 84.515 218.335 84.745 224.785 ;
        RECT 89.095 218.335 89.325 224.785 ;
        RECT 93.675 218.335 93.905 224.785 ;
        RECT 98.255 218.335 98.485 224.785 ;
        RECT 102.835 218.335 103.065 224.785 ;
        RECT 107.415 218.335 107.645 224.785 ;
        RECT 110.930 218.520 111.250 218.580 ;
        RECT 111.995 218.520 112.225 224.785 ;
        RECT 110.930 218.380 112.225 218.520 ;
        RECT 110.930 218.320 111.250 218.380 ;
        RECT 111.995 218.335 112.225 218.380 ;
        RECT 116.575 218.335 116.805 224.785 ;
        RECT 121.155 218.335 121.385 224.785 ;
        RECT 125.735 218.335 125.965 224.785 ;
        RECT 130.315 218.335 130.545 224.785 ;
        RECT 134.895 218.335 135.125 224.785 ;
        RECT 139.475 218.335 139.705 224.785 ;
        RECT 144.055 218.335 144.285 224.785 ;
        RECT 148.635 218.335 148.865 224.785 ;
        RECT 153.215 218.335 153.445 224.785 ;
        RECT 157.795 218.335 158.025 224.785 ;
        RECT 162.375 218.335 162.605 224.785 ;
        RECT 166.955 218.335 167.185 224.785 ;
        RECT 171.535 218.335 171.765 224.785 ;
        RECT 176.115 218.335 176.345 224.785 ;
        RECT 180.695 218.335 180.925 224.785 ;
        RECT 185.275 218.335 185.505 224.785 ;
        RECT 189.855 218.335 190.085 224.785 ;
        RECT 194.435 218.335 194.665 224.785 ;
        RECT 199.015 218.335 199.245 224.785 ;
        RECT 203.595 218.335 203.825 224.785 ;
        RECT 208.175 218.335 208.405 224.785 ;
        RECT 212.755 218.335 212.985 224.785 ;
        RECT 75.050 217.840 75.370 217.900 ;
        RECT 74.775 217.700 75.370 217.840 ;
        RECT 75.050 217.640 75.370 217.700 ;
        RECT 113.575 199.535 113.805 205.985 ;
        RECT 118.155 199.535 118.385 205.985 ;
        RECT 122.735 199.535 122.965 205.985 ;
        RECT 127.315 199.535 127.545 205.985 ;
        RECT 131.895 199.535 132.125 205.985 ;
        RECT 136.475 199.535 136.705 205.985 ;
        RECT 141.055 199.535 141.285 205.985 ;
        RECT 110.930 199.140 111.250 199.200 ;
        RECT 113.705 199.140 113.995 199.185 ;
        RECT 140.370 199.140 140.690 199.200 ;
        RECT 110.930 199.000 113.995 199.140 ;
        RECT 140.095 199.000 140.690 199.140 ;
        RECT 110.930 198.940 111.250 199.000 ;
        RECT 113.705 198.955 113.995 199.000 ;
        RECT 140.370 198.940 140.690 199.000 ;
        RECT 64.470 185.680 64.790 185.940 ;
        RECT 64.560 185.185 64.700 185.680 ;
        RECT 61.785 182.135 64.835 185.185 ;
        RECT 140.370 180.780 140.690 180.840 ;
        RECT 140.095 180.640 140.690 180.780 ;
        RECT 140.370 180.580 140.690 180.640 ;
        RECT 110.095 146.755 112.145 149.565 ;
      LAYER via ;
        RECT 110.960 218.320 111.220 218.580 ;
        RECT 75.080 217.640 75.340 217.900 ;
        RECT 110.960 198.940 111.220 199.200 ;
        RECT 140.400 198.940 140.660 199.200 ;
        RECT 64.500 185.680 64.760 185.940 ;
        RECT 140.400 180.580 140.660 180.840 ;
        RECT 110.960 149.300 111.220 149.560 ;
      LAYER met2 ;
        RECT 29.580 243.210 30.580 243.610 ;
        RECT 66.820 243.210 67.820 243.610 ;
        RECT 29.580 224.410 30.580 224.810 ;
        RECT 75.070 218.865 75.350 219.235 ;
        RECT 75.140 217.930 75.280 218.865 ;
        RECT 110.960 218.290 111.220 218.610 ;
        RECT 75.080 217.610 75.340 217.930 ;
        RECT 111.020 207.035 111.160 218.290 ;
        RECT 110.950 206.665 111.230 207.035 ;
        RECT 31.540 205.610 32.540 206.010 ;
        RECT 75.640 205.610 76.640 206.010 ;
        RECT 111.020 199.230 111.160 206.665 ;
        RECT 110.960 198.910 111.220 199.230 ;
        RECT 140.400 198.910 140.660 199.230 ;
        RECT 64.490 185.925 64.770 186.295 ;
        RECT 64.500 185.650 64.760 185.925 ;
        RECT 111.020 149.590 111.160 198.910 ;
        RECT 140.460 180.870 140.600 198.910 ;
        RECT 140.400 180.550 140.660 180.870 ;
        RECT 110.960 149.270 111.220 149.590 ;
      LAYER via2 ;
        RECT 29.740 243.270 30.020 243.550 ;
        RECT 30.140 243.270 30.420 243.550 ;
        RECT 66.980 243.270 67.260 243.550 ;
        RECT 67.380 243.270 67.660 243.550 ;
        RECT 29.740 224.470 30.020 224.750 ;
        RECT 30.140 224.470 30.420 224.750 ;
        RECT 75.070 218.910 75.350 219.190 ;
        RECT 110.950 206.710 111.230 206.990 ;
        RECT 31.700 205.670 31.980 205.950 ;
        RECT 32.100 205.670 32.380 205.950 ;
        RECT 75.800 205.670 76.080 205.950 ;
        RECT 76.200 205.670 76.480 205.950 ;
        RECT 64.490 185.970 64.770 186.250 ;
      LAYER met3 ;
        RECT 29.580 237.110 65.440 243.610 ;
        RECT 66.820 237.110 102.680 243.610 ;
        RECT 29.580 218.310 65.440 224.810 ;
        RECT 66.970 219.200 67.350 219.210 ;
        RECT 75.045 219.200 75.375 219.215 ;
        RECT 66.970 218.900 75.375 219.200 ;
        RECT 66.970 218.890 67.350 218.900 ;
        RECT 75.045 218.885 75.375 218.900 ;
        RECT 110.925 207.010 111.255 207.015 ;
        RECT 34.540 207.000 34.920 207.010 ;
        RECT 110.925 207.000 111.510 207.010 ;
        RECT 25.840 206.700 34.920 207.000 ;
        RECT 110.710 206.700 111.510 207.000 ;
        RECT 25.840 205.170 26.140 206.700 ;
        RECT 34.540 206.690 34.920 206.700 ;
        RECT 110.925 206.690 111.510 206.700 ;
        RECT 110.925 206.685 111.255 206.690 ;
        RECT 0.000 204.870 26.140 205.170 ;
        RECT 31.540 199.510 67.400 206.010 ;
        RECT 75.640 199.510 111.500 206.010 ;
        RECT 64.465 186.260 64.795 186.275 ;
        RECT 67.660 186.260 68.040 186.270 ;
        RECT 64.465 185.960 68.040 186.260 ;
        RECT 64.465 185.945 64.795 185.960 ;
        RECT 67.660 185.950 68.040 185.960 ;
      LAYER via3 ;
        RECT 32.660 243.150 32.980 243.470 ;
        RECT 36.255 243.150 36.575 243.470 ;
        RECT 39.850 243.150 40.170 243.470 ;
        RECT 43.445 243.150 43.765 243.470 ;
        RECT 47.040 243.150 47.360 243.470 ;
        RECT 50.635 243.150 50.955 243.470 ;
        RECT 54.230 243.150 54.550 243.470 ;
        RECT 57.825 243.150 58.145 243.470 ;
        RECT 61.420 243.150 61.740 243.470 ;
        RECT 65.015 243.150 65.335 243.470 ;
        RECT 32.660 242.750 32.980 243.070 ;
        RECT 36.255 242.750 36.575 243.070 ;
        RECT 39.850 242.750 40.170 243.070 ;
        RECT 43.445 242.750 43.765 243.070 ;
        RECT 47.040 242.750 47.360 243.070 ;
        RECT 50.635 242.750 50.955 243.070 ;
        RECT 54.230 242.750 54.550 243.070 ;
        RECT 57.825 242.750 58.145 243.070 ;
        RECT 61.420 242.750 61.740 243.070 ;
        RECT 65.015 242.750 65.335 243.070 ;
        RECT 32.660 242.350 32.980 242.670 ;
        RECT 36.255 242.350 36.575 242.670 ;
        RECT 39.850 242.350 40.170 242.670 ;
        RECT 43.445 242.350 43.765 242.670 ;
        RECT 47.040 242.350 47.360 242.670 ;
        RECT 50.635 242.350 50.955 242.670 ;
        RECT 54.230 242.350 54.550 242.670 ;
        RECT 57.825 242.350 58.145 242.670 ;
        RECT 61.420 242.350 61.740 242.670 ;
        RECT 65.015 242.350 65.335 242.670 ;
        RECT 32.660 241.950 32.980 242.270 ;
        RECT 36.255 241.950 36.575 242.270 ;
        RECT 39.850 241.950 40.170 242.270 ;
        RECT 43.445 241.950 43.765 242.270 ;
        RECT 47.040 241.950 47.360 242.270 ;
        RECT 50.635 241.950 50.955 242.270 ;
        RECT 54.230 241.950 54.550 242.270 ;
        RECT 57.825 241.950 58.145 242.270 ;
        RECT 61.420 241.950 61.740 242.270 ;
        RECT 65.015 241.950 65.335 242.270 ;
        RECT 32.660 241.550 32.980 241.870 ;
        RECT 36.255 241.550 36.575 241.870 ;
        RECT 39.850 241.550 40.170 241.870 ;
        RECT 43.445 241.550 43.765 241.870 ;
        RECT 47.040 241.550 47.360 241.870 ;
        RECT 50.635 241.550 50.955 241.870 ;
        RECT 54.230 241.550 54.550 241.870 ;
        RECT 57.825 241.550 58.145 241.870 ;
        RECT 61.420 241.550 61.740 241.870 ;
        RECT 65.015 241.550 65.335 241.870 ;
        RECT 32.660 241.150 32.980 241.470 ;
        RECT 36.255 241.150 36.575 241.470 ;
        RECT 39.850 241.150 40.170 241.470 ;
        RECT 43.445 241.150 43.765 241.470 ;
        RECT 47.040 241.150 47.360 241.470 ;
        RECT 50.635 241.150 50.955 241.470 ;
        RECT 54.230 241.150 54.550 241.470 ;
        RECT 57.825 241.150 58.145 241.470 ;
        RECT 61.420 241.150 61.740 241.470 ;
        RECT 65.015 241.150 65.335 241.470 ;
        RECT 32.660 240.750 32.980 241.070 ;
        RECT 36.255 240.750 36.575 241.070 ;
        RECT 39.850 240.750 40.170 241.070 ;
        RECT 43.445 240.750 43.765 241.070 ;
        RECT 47.040 240.750 47.360 241.070 ;
        RECT 50.635 240.750 50.955 241.070 ;
        RECT 54.230 240.750 54.550 241.070 ;
        RECT 57.825 240.750 58.145 241.070 ;
        RECT 61.420 240.750 61.740 241.070 ;
        RECT 65.015 240.750 65.335 241.070 ;
        RECT 32.660 239.650 32.980 239.970 ;
        RECT 36.255 239.650 36.575 239.970 ;
        RECT 39.850 239.650 40.170 239.970 ;
        RECT 43.445 239.650 43.765 239.970 ;
        RECT 47.040 239.650 47.360 239.970 ;
        RECT 50.635 239.650 50.955 239.970 ;
        RECT 54.230 239.650 54.550 239.970 ;
        RECT 57.825 239.650 58.145 239.970 ;
        RECT 61.420 239.650 61.740 239.970 ;
        RECT 65.015 239.650 65.335 239.970 ;
        RECT 32.660 239.250 32.980 239.570 ;
        RECT 36.255 239.250 36.575 239.570 ;
        RECT 39.850 239.250 40.170 239.570 ;
        RECT 43.445 239.250 43.765 239.570 ;
        RECT 47.040 239.250 47.360 239.570 ;
        RECT 50.635 239.250 50.955 239.570 ;
        RECT 54.230 239.250 54.550 239.570 ;
        RECT 57.825 239.250 58.145 239.570 ;
        RECT 61.420 239.250 61.740 239.570 ;
        RECT 65.015 239.250 65.335 239.570 ;
        RECT 32.660 238.850 32.980 239.170 ;
        RECT 36.255 238.850 36.575 239.170 ;
        RECT 39.850 238.850 40.170 239.170 ;
        RECT 43.445 238.850 43.765 239.170 ;
        RECT 47.040 238.850 47.360 239.170 ;
        RECT 50.635 238.850 50.955 239.170 ;
        RECT 54.230 238.850 54.550 239.170 ;
        RECT 57.825 238.850 58.145 239.170 ;
        RECT 61.420 238.850 61.740 239.170 ;
        RECT 65.015 238.850 65.335 239.170 ;
        RECT 32.660 238.450 32.980 238.770 ;
        RECT 36.255 238.450 36.575 238.770 ;
        RECT 39.850 238.450 40.170 238.770 ;
        RECT 43.445 238.450 43.765 238.770 ;
        RECT 47.040 238.450 47.360 238.770 ;
        RECT 50.635 238.450 50.955 238.770 ;
        RECT 54.230 238.450 54.550 238.770 ;
        RECT 57.825 238.450 58.145 238.770 ;
        RECT 61.420 238.450 61.740 238.770 ;
        RECT 65.015 238.450 65.335 238.770 ;
        RECT 32.660 238.050 32.980 238.370 ;
        RECT 36.255 238.050 36.575 238.370 ;
        RECT 39.850 238.050 40.170 238.370 ;
        RECT 43.445 238.050 43.765 238.370 ;
        RECT 47.040 238.050 47.360 238.370 ;
        RECT 50.635 238.050 50.955 238.370 ;
        RECT 54.230 238.050 54.550 238.370 ;
        RECT 57.825 238.050 58.145 238.370 ;
        RECT 61.420 238.050 61.740 238.370 ;
        RECT 65.015 238.050 65.335 238.370 ;
        RECT 32.660 237.650 32.980 237.970 ;
        RECT 36.255 237.650 36.575 237.970 ;
        RECT 39.850 237.650 40.170 237.970 ;
        RECT 43.445 237.650 43.765 237.970 ;
        RECT 47.040 237.650 47.360 237.970 ;
        RECT 50.635 237.650 50.955 237.970 ;
        RECT 54.230 237.650 54.550 237.970 ;
        RECT 57.825 237.650 58.145 237.970 ;
        RECT 61.420 237.650 61.740 237.970 ;
        RECT 65.015 237.650 65.335 237.970 ;
        RECT 32.660 237.250 32.980 237.570 ;
        RECT 36.255 237.250 36.575 237.570 ;
        RECT 39.850 237.250 40.170 237.570 ;
        RECT 43.445 237.250 43.765 237.570 ;
        RECT 47.040 237.250 47.360 237.570 ;
        RECT 50.635 237.250 50.955 237.570 ;
        RECT 54.230 237.250 54.550 237.570 ;
        RECT 57.825 237.250 58.145 237.570 ;
        RECT 61.420 237.250 61.740 237.570 ;
        RECT 65.015 237.250 65.335 237.570 ;
        RECT 69.900 243.150 70.220 243.470 ;
        RECT 73.495 243.150 73.815 243.470 ;
        RECT 77.090 243.150 77.410 243.470 ;
        RECT 80.685 243.150 81.005 243.470 ;
        RECT 84.280 243.150 84.600 243.470 ;
        RECT 87.875 243.150 88.195 243.470 ;
        RECT 91.470 243.150 91.790 243.470 ;
        RECT 95.065 243.150 95.385 243.470 ;
        RECT 98.660 243.150 98.980 243.470 ;
        RECT 102.255 243.150 102.575 243.470 ;
        RECT 69.900 242.750 70.220 243.070 ;
        RECT 73.495 242.750 73.815 243.070 ;
        RECT 77.090 242.750 77.410 243.070 ;
        RECT 80.685 242.750 81.005 243.070 ;
        RECT 84.280 242.750 84.600 243.070 ;
        RECT 87.875 242.750 88.195 243.070 ;
        RECT 91.470 242.750 91.790 243.070 ;
        RECT 95.065 242.750 95.385 243.070 ;
        RECT 98.660 242.750 98.980 243.070 ;
        RECT 102.255 242.750 102.575 243.070 ;
        RECT 69.900 242.350 70.220 242.670 ;
        RECT 73.495 242.350 73.815 242.670 ;
        RECT 77.090 242.350 77.410 242.670 ;
        RECT 80.685 242.350 81.005 242.670 ;
        RECT 84.280 242.350 84.600 242.670 ;
        RECT 87.875 242.350 88.195 242.670 ;
        RECT 91.470 242.350 91.790 242.670 ;
        RECT 95.065 242.350 95.385 242.670 ;
        RECT 98.660 242.350 98.980 242.670 ;
        RECT 102.255 242.350 102.575 242.670 ;
        RECT 69.900 241.950 70.220 242.270 ;
        RECT 73.495 241.950 73.815 242.270 ;
        RECT 77.090 241.950 77.410 242.270 ;
        RECT 80.685 241.950 81.005 242.270 ;
        RECT 84.280 241.950 84.600 242.270 ;
        RECT 87.875 241.950 88.195 242.270 ;
        RECT 91.470 241.950 91.790 242.270 ;
        RECT 95.065 241.950 95.385 242.270 ;
        RECT 98.660 241.950 98.980 242.270 ;
        RECT 102.255 241.950 102.575 242.270 ;
        RECT 69.900 241.550 70.220 241.870 ;
        RECT 73.495 241.550 73.815 241.870 ;
        RECT 77.090 241.550 77.410 241.870 ;
        RECT 80.685 241.550 81.005 241.870 ;
        RECT 84.280 241.550 84.600 241.870 ;
        RECT 87.875 241.550 88.195 241.870 ;
        RECT 91.470 241.550 91.790 241.870 ;
        RECT 95.065 241.550 95.385 241.870 ;
        RECT 98.660 241.550 98.980 241.870 ;
        RECT 102.255 241.550 102.575 241.870 ;
        RECT 69.900 241.150 70.220 241.470 ;
        RECT 73.495 241.150 73.815 241.470 ;
        RECT 77.090 241.150 77.410 241.470 ;
        RECT 80.685 241.150 81.005 241.470 ;
        RECT 84.280 241.150 84.600 241.470 ;
        RECT 87.875 241.150 88.195 241.470 ;
        RECT 91.470 241.150 91.790 241.470 ;
        RECT 95.065 241.150 95.385 241.470 ;
        RECT 98.660 241.150 98.980 241.470 ;
        RECT 102.255 241.150 102.575 241.470 ;
        RECT 69.900 240.750 70.220 241.070 ;
        RECT 73.495 240.750 73.815 241.070 ;
        RECT 77.090 240.750 77.410 241.070 ;
        RECT 80.685 240.750 81.005 241.070 ;
        RECT 84.280 240.750 84.600 241.070 ;
        RECT 87.875 240.750 88.195 241.070 ;
        RECT 91.470 240.750 91.790 241.070 ;
        RECT 95.065 240.750 95.385 241.070 ;
        RECT 98.660 240.750 98.980 241.070 ;
        RECT 102.255 240.750 102.575 241.070 ;
        RECT 69.900 239.650 70.220 239.970 ;
        RECT 73.495 239.650 73.815 239.970 ;
        RECT 77.090 239.650 77.410 239.970 ;
        RECT 80.685 239.650 81.005 239.970 ;
        RECT 84.280 239.650 84.600 239.970 ;
        RECT 87.875 239.650 88.195 239.970 ;
        RECT 91.470 239.650 91.790 239.970 ;
        RECT 95.065 239.650 95.385 239.970 ;
        RECT 98.660 239.650 98.980 239.970 ;
        RECT 102.255 239.650 102.575 239.970 ;
        RECT 69.900 239.250 70.220 239.570 ;
        RECT 73.495 239.250 73.815 239.570 ;
        RECT 77.090 239.250 77.410 239.570 ;
        RECT 80.685 239.250 81.005 239.570 ;
        RECT 84.280 239.250 84.600 239.570 ;
        RECT 87.875 239.250 88.195 239.570 ;
        RECT 91.470 239.250 91.790 239.570 ;
        RECT 95.065 239.250 95.385 239.570 ;
        RECT 98.660 239.250 98.980 239.570 ;
        RECT 102.255 239.250 102.575 239.570 ;
        RECT 69.900 238.850 70.220 239.170 ;
        RECT 73.495 238.850 73.815 239.170 ;
        RECT 77.090 238.850 77.410 239.170 ;
        RECT 80.685 238.850 81.005 239.170 ;
        RECT 84.280 238.850 84.600 239.170 ;
        RECT 87.875 238.850 88.195 239.170 ;
        RECT 91.470 238.850 91.790 239.170 ;
        RECT 95.065 238.850 95.385 239.170 ;
        RECT 98.660 238.850 98.980 239.170 ;
        RECT 102.255 238.850 102.575 239.170 ;
        RECT 69.900 238.450 70.220 238.770 ;
        RECT 73.495 238.450 73.815 238.770 ;
        RECT 77.090 238.450 77.410 238.770 ;
        RECT 80.685 238.450 81.005 238.770 ;
        RECT 84.280 238.450 84.600 238.770 ;
        RECT 87.875 238.450 88.195 238.770 ;
        RECT 91.470 238.450 91.790 238.770 ;
        RECT 95.065 238.450 95.385 238.770 ;
        RECT 98.660 238.450 98.980 238.770 ;
        RECT 102.255 238.450 102.575 238.770 ;
        RECT 69.900 238.050 70.220 238.370 ;
        RECT 73.495 238.050 73.815 238.370 ;
        RECT 77.090 238.050 77.410 238.370 ;
        RECT 80.685 238.050 81.005 238.370 ;
        RECT 84.280 238.050 84.600 238.370 ;
        RECT 87.875 238.050 88.195 238.370 ;
        RECT 91.470 238.050 91.790 238.370 ;
        RECT 95.065 238.050 95.385 238.370 ;
        RECT 98.660 238.050 98.980 238.370 ;
        RECT 102.255 238.050 102.575 238.370 ;
        RECT 69.900 237.650 70.220 237.970 ;
        RECT 73.495 237.650 73.815 237.970 ;
        RECT 77.090 237.650 77.410 237.970 ;
        RECT 80.685 237.650 81.005 237.970 ;
        RECT 84.280 237.650 84.600 237.970 ;
        RECT 87.875 237.650 88.195 237.970 ;
        RECT 91.470 237.650 91.790 237.970 ;
        RECT 95.065 237.650 95.385 237.970 ;
        RECT 98.660 237.650 98.980 237.970 ;
        RECT 102.255 237.650 102.575 237.970 ;
        RECT 69.900 237.250 70.220 237.570 ;
        RECT 73.495 237.250 73.815 237.570 ;
        RECT 77.090 237.250 77.410 237.570 ;
        RECT 80.685 237.250 81.005 237.570 ;
        RECT 84.280 237.250 84.600 237.570 ;
        RECT 87.875 237.250 88.195 237.570 ;
        RECT 91.470 237.250 91.790 237.570 ;
        RECT 95.065 237.250 95.385 237.570 ;
        RECT 98.660 237.250 98.980 237.570 ;
        RECT 102.255 237.250 102.575 237.570 ;
        RECT 32.660 224.350 32.980 224.670 ;
        RECT 36.255 224.350 36.575 224.670 ;
        RECT 39.850 224.350 40.170 224.670 ;
        RECT 43.445 224.350 43.765 224.670 ;
        RECT 47.040 224.350 47.360 224.670 ;
        RECT 50.635 224.350 50.955 224.670 ;
        RECT 54.230 224.350 54.550 224.670 ;
        RECT 57.825 224.350 58.145 224.670 ;
        RECT 61.420 224.350 61.740 224.670 ;
        RECT 65.015 224.350 65.335 224.670 ;
        RECT 32.660 223.950 32.980 224.270 ;
        RECT 36.255 223.950 36.575 224.270 ;
        RECT 39.850 223.950 40.170 224.270 ;
        RECT 43.445 223.950 43.765 224.270 ;
        RECT 47.040 223.950 47.360 224.270 ;
        RECT 50.635 223.950 50.955 224.270 ;
        RECT 54.230 223.950 54.550 224.270 ;
        RECT 57.825 223.950 58.145 224.270 ;
        RECT 61.420 223.950 61.740 224.270 ;
        RECT 65.015 223.950 65.335 224.270 ;
        RECT 32.660 223.550 32.980 223.870 ;
        RECT 36.255 223.550 36.575 223.870 ;
        RECT 39.850 223.550 40.170 223.870 ;
        RECT 43.445 223.550 43.765 223.870 ;
        RECT 47.040 223.550 47.360 223.870 ;
        RECT 50.635 223.550 50.955 223.870 ;
        RECT 54.230 223.550 54.550 223.870 ;
        RECT 57.825 223.550 58.145 223.870 ;
        RECT 61.420 223.550 61.740 223.870 ;
        RECT 65.015 223.550 65.335 223.870 ;
        RECT 32.660 223.150 32.980 223.470 ;
        RECT 36.255 223.150 36.575 223.470 ;
        RECT 39.850 223.150 40.170 223.470 ;
        RECT 43.445 223.150 43.765 223.470 ;
        RECT 47.040 223.150 47.360 223.470 ;
        RECT 50.635 223.150 50.955 223.470 ;
        RECT 54.230 223.150 54.550 223.470 ;
        RECT 57.825 223.150 58.145 223.470 ;
        RECT 61.420 223.150 61.740 223.470 ;
        RECT 65.015 223.150 65.335 223.470 ;
        RECT 32.660 222.750 32.980 223.070 ;
        RECT 36.255 222.750 36.575 223.070 ;
        RECT 39.850 222.750 40.170 223.070 ;
        RECT 43.445 222.750 43.765 223.070 ;
        RECT 47.040 222.750 47.360 223.070 ;
        RECT 50.635 222.750 50.955 223.070 ;
        RECT 54.230 222.750 54.550 223.070 ;
        RECT 57.825 222.750 58.145 223.070 ;
        RECT 61.420 222.750 61.740 223.070 ;
        RECT 65.015 222.750 65.335 223.070 ;
        RECT 32.660 222.350 32.980 222.670 ;
        RECT 36.255 222.350 36.575 222.670 ;
        RECT 39.850 222.350 40.170 222.670 ;
        RECT 43.445 222.350 43.765 222.670 ;
        RECT 47.040 222.350 47.360 222.670 ;
        RECT 50.635 222.350 50.955 222.670 ;
        RECT 54.230 222.350 54.550 222.670 ;
        RECT 57.825 222.350 58.145 222.670 ;
        RECT 61.420 222.350 61.740 222.670 ;
        RECT 65.015 222.350 65.335 222.670 ;
        RECT 32.660 221.950 32.980 222.270 ;
        RECT 36.255 221.950 36.575 222.270 ;
        RECT 39.850 221.950 40.170 222.270 ;
        RECT 43.445 221.950 43.765 222.270 ;
        RECT 47.040 221.950 47.360 222.270 ;
        RECT 50.635 221.950 50.955 222.270 ;
        RECT 54.230 221.950 54.550 222.270 ;
        RECT 57.825 221.950 58.145 222.270 ;
        RECT 61.420 221.950 61.740 222.270 ;
        RECT 65.015 221.950 65.335 222.270 ;
        RECT 32.660 220.850 32.980 221.170 ;
        RECT 36.255 220.850 36.575 221.170 ;
        RECT 39.850 220.850 40.170 221.170 ;
        RECT 43.445 220.850 43.765 221.170 ;
        RECT 47.040 220.850 47.360 221.170 ;
        RECT 50.635 220.850 50.955 221.170 ;
        RECT 54.230 220.850 54.550 221.170 ;
        RECT 57.825 220.850 58.145 221.170 ;
        RECT 61.420 220.850 61.740 221.170 ;
        RECT 65.015 220.850 65.335 221.170 ;
        RECT 32.660 220.450 32.980 220.770 ;
        RECT 36.255 220.450 36.575 220.770 ;
        RECT 39.850 220.450 40.170 220.770 ;
        RECT 43.445 220.450 43.765 220.770 ;
        RECT 47.040 220.450 47.360 220.770 ;
        RECT 50.635 220.450 50.955 220.770 ;
        RECT 54.230 220.450 54.550 220.770 ;
        RECT 57.825 220.450 58.145 220.770 ;
        RECT 61.420 220.450 61.740 220.770 ;
        RECT 65.015 220.450 65.335 220.770 ;
        RECT 32.660 220.050 32.980 220.370 ;
        RECT 36.255 220.050 36.575 220.370 ;
        RECT 39.850 220.050 40.170 220.370 ;
        RECT 43.445 220.050 43.765 220.370 ;
        RECT 47.040 220.050 47.360 220.370 ;
        RECT 50.635 220.050 50.955 220.370 ;
        RECT 54.230 220.050 54.550 220.370 ;
        RECT 57.825 220.050 58.145 220.370 ;
        RECT 61.420 220.050 61.740 220.370 ;
        RECT 65.015 220.050 65.335 220.370 ;
        RECT 32.660 219.650 32.980 219.970 ;
        RECT 36.255 219.650 36.575 219.970 ;
        RECT 39.850 219.650 40.170 219.970 ;
        RECT 43.445 219.650 43.765 219.970 ;
        RECT 47.040 219.650 47.360 219.970 ;
        RECT 50.635 219.650 50.955 219.970 ;
        RECT 54.230 219.650 54.550 219.970 ;
        RECT 57.825 219.650 58.145 219.970 ;
        RECT 61.420 219.650 61.740 219.970 ;
        RECT 65.015 219.650 65.335 219.970 ;
        RECT 32.660 219.250 32.980 219.570 ;
        RECT 36.255 219.250 36.575 219.570 ;
        RECT 39.850 219.250 40.170 219.570 ;
        RECT 43.445 219.250 43.765 219.570 ;
        RECT 47.040 219.250 47.360 219.570 ;
        RECT 50.635 219.250 50.955 219.570 ;
        RECT 54.230 219.250 54.550 219.570 ;
        RECT 57.825 219.250 58.145 219.570 ;
        RECT 61.420 219.250 61.740 219.570 ;
        RECT 65.015 219.250 65.335 219.570 ;
        RECT 32.660 218.850 32.980 219.170 ;
        RECT 36.255 218.850 36.575 219.170 ;
        RECT 39.850 218.850 40.170 219.170 ;
        RECT 43.445 218.850 43.765 219.170 ;
        RECT 47.040 218.850 47.360 219.170 ;
        RECT 50.635 218.850 50.955 219.170 ;
        RECT 54.230 218.850 54.550 219.170 ;
        RECT 57.825 218.850 58.145 219.170 ;
        RECT 61.420 218.850 61.740 219.170 ;
        RECT 65.015 218.850 65.335 219.170 ;
        RECT 67.000 218.890 67.320 219.210 ;
        RECT 32.660 218.450 32.980 218.770 ;
        RECT 36.255 218.450 36.575 218.770 ;
        RECT 39.850 218.450 40.170 218.770 ;
        RECT 43.445 218.450 43.765 218.770 ;
        RECT 47.040 218.450 47.360 218.770 ;
        RECT 50.635 218.450 50.955 218.770 ;
        RECT 54.230 218.450 54.550 218.770 ;
        RECT 57.825 218.450 58.145 218.770 ;
        RECT 61.420 218.450 61.740 218.770 ;
        RECT 65.015 218.450 65.335 218.770 ;
        RECT 34.570 206.690 34.890 207.010 ;
        RECT 111.160 206.690 111.480 207.010 ;
        RECT 34.620 205.550 34.940 205.870 ;
        RECT 38.215 205.550 38.535 205.870 ;
        RECT 41.810 205.550 42.130 205.870 ;
        RECT 45.405 205.550 45.725 205.870 ;
        RECT 49.000 205.550 49.320 205.870 ;
        RECT 52.595 205.550 52.915 205.870 ;
        RECT 56.190 205.550 56.510 205.870 ;
        RECT 59.785 205.550 60.105 205.870 ;
        RECT 63.380 205.550 63.700 205.870 ;
        RECT 66.975 205.550 67.295 205.870 ;
        RECT 34.620 205.150 34.940 205.470 ;
        RECT 38.215 205.150 38.535 205.470 ;
        RECT 41.810 205.150 42.130 205.470 ;
        RECT 45.405 205.150 45.725 205.470 ;
        RECT 49.000 205.150 49.320 205.470 ;
        RECT 52.595 205.150 52.915 205.470 ;
        RECT 56.190 205.150 56.510 205.470 ;
        RECT 59.785 205.150 60.105 205.470 ;
        RECT 63.380 205.150 63.700 205.470 ;
        RECT 66.975 205.150 67.295 205.470 ;
        RECT 34.620 204.750 34.940 205.070 ;
        RECT 38.215 204.750 38.535 205.070 ;
        RECT 41.810 204.750 42.130 205.070 ;
        RECT 45.405 204.750 45.725 205.070 ;
        RECT 49.000 204.750 49.320 205.070 ;
        RECT 52.595 204.750 52.915 205.070 ;
        RECT 56.190 204.750 56.510 205.070 ;
        RECT 59.785 204.750 60.105 205.070 ;
        RECT 63.380 204.750 63.700 205.070 ;
        RECT 66.975 204.750 67.295 205.070 ;
        RECT 34.620 204.350 34.940 204.670 ;
        RECT 38.215 204.350 38.535 204.670 ;
        RECT 41.810 204.350 42.130 204.670 ;
        RECT 45.405 204.350 45.725 204.670 ;
        RECT 49.000 204.350 49.320 204.670 ;
        RECT 52.595 204.350 52.915 204.670 ;
        RECT 56.190 204.350 56.510 204.670 ;
        RECT 59.785 204.350 60.105 204.670 ;
        RECT 63.380 204.350 63.700 204.670 ;
        RECT 66.975 204.350 67.295 204.670 ;
        RECT 34.620 203.950 34.940 204.270 ;
        RECT 38.215 203.950 38.535 204.270 ;
        RECT 41.810 203.950 42.130 204.270 ;
        RECT 45.405 203.950 45.725 204.270 ;
        RECT 49.000 203.950 49.320 204.270 ;
        RECT 52.595 203.950 52.915 204.270 ;
        RECT 56.190 203.950 56.510 204.270 ;
        RECT 59.785 203.950 60.105 204.270 ;
        RECT 63.380 203.950 63.700 204.270 ;
        RECT 66.975 203.950 67.295 204.270 ;
        RECT 34.620 203.550 34.940 203.870 ;
        RECT 38.215 203.550 38.535 203.870 ;
        RECT 41.810 203.550 42.130 203.870 ;
        RECT 45.405 203.550 45.725 203.870 ;
        RECT 49.000 203.550 49.320 203.870 ;
        RECT 52.595 203.550 52.915 203.870 ;
        RECT 56.190 203.550 56.510 203.870 ;
        RECT 59.785 203.550 60.105 203.870 ;
        RECT 63.380 203.550 63.700 203.870 ;
        RECT 66.975 203.550 67.295 203.870 ;
        RECT 34.620 203.150 34.940 203.470 ;
        RECT 38.215 203.150 38.535 203.470 ;
        RECT 41.810 203.150 42.130 203.470 ;
        RECT 45.405 203.150 45.725 203.470 ;
        RECT 49.000 203.150 49.320 203.470 ;
        RECT 52.595 203.150 52.915 203.470 ;
        RECT 56.190 203.150 56.510 203.470 ;
        RECT 59.785 203.150 60.105 203.470 ;
        RECT 63.380 203.150 63.700 203.470 ;
        RECT 66.975 203.150 67.295 203.470 ;
        RECT 34.620 202.050 34.940 202.370 ;
        RECT 38.215 202.050 38.535 202.370 ;
        RECT 41.810 202.050 42.130 202.370 ;
        RECT 45.405 202.050 45.725 202.370 ;
        RECT 49.000 202.050 49.320 202.370 ;
        RECT 52.595 202.050 52.915 202.370 ;
        RECT 56.190 202.050 56.510 202.370 ;
        RECT 59.785 202.050 60.105 202.370 ;
        RECT 63.380 202.050 63.700 202.370 ;
        RECT 66.975 202.050 67.295 202.370 ;
        RECT 34.620 201.650 34.940 201.970 ;
        RECT 38.215 201.650 38.535 201.970 ;
        RECT 41.810 201.650 42.130 201.970 ;
        RECT 45.405 201.650 45.725 201.970 ;
        RECT 49.000 201.650 49.320 201.970 ;
        RECT 52.595 201.650 52.915 201.970 ;
        RECT 56.190 201.650 56.510 201.970 ;
        RECT 59.785 201.650 60.105 201.970 ;
        RECT 63.380 201.650 63.700 201.970 ;
        RECT 66.975 201.650 67.295 201.970 ;
        RECT 34.620 201.250 34.940 201.570 ;
        RECT 38.215 201.250 38.535 201.570 ;
        RECT 41.810 201.250 42.130 201.570 ;
        RECT 45.405 201.250 45.725 201.570 ;
        RECT 49.000 201.250 49.320 201.570 ;
        RECT 52.595 201.250 52.915 201.570 ;
        RECT 56.190 201.250 56.510 201.570 ;
        RECT 59.785 201.250 60.105 201.570 ;
        RECT 63.380 201.250 63.700 201.570 ;
        RECT 66.975 201.250 67.295 201.570 ;
        RECT 34.620 200.850 34.940 201.170 ;
        RECT 38.215 200.850 38.535 201.170 ;
        RECT 41.810 200.850 42.130 201.170 ;
        RECT 45.405 200.850 45.725 201.170 ;
        RECT 49.000 200.850 49.320 201.170 ;
        RECT 52.595 200.850 52.915 201.170 ;
        RECT 56.190 200.850 56.510 201.170 ;
        RECT 59.785 200.850 60.105 201.170 ;
        RECT 63.380 200.850 63.700 201.170 ;
        RECT 66.975 200.850 67.295 201.170 ;
        RECT 34.620 200.450 34.940 200.770 ;
        RECT 38.215 200.450 38.535 200.770 ;
        RECT 41.810 200.450 42.130 200.770 ;
        RECT 45.405 200.450 45.725 200.770 ;
        RECT 49.000 200.450 49.320 200.770 ;
        RECT 52.595 200.450 52.915 200.770 ;
        RECT 56.190 200.450 56.510 200.770 ;
        RECT 59.785 200.450 60.105 200.770 ;
        RECT 63.380 200.450 63.700 200.770 ;
        RECT 66.975 200.450 67.295 200.770 ;
        RECT 34.620 200.050 34.940 200.370 ;
        RECT 38.215 200.050 38.535 200.370 ;
        RECT 41.810 200.050 42.130 200.370 ;
        RECT 45.405 200.050 45.725 200.370 ;
        RECT 49.000 200.050 49.320 200.370 ;
        RECT 52.595 200.050 52.915 200.370 ;
        RECT 56.190 200.050 56.510 200.370 ;
        RECT 59.785 200.050 60.105 200.370 ;
        RECT 63.380 200.050 63.700 200.370 ;
        RECT 66.975 200.050 67.295 200.370 ;
        RECT 34.620 199.650 34.940 199.970 ;
        RECT 38.215 199.650 38.535 199.970 ;
        RECT 41.810 199.650 42.130 199.970 ;
        RECT 45.405 199.650 45.725 199.970 ;
        RECT 49.000 199.650 49.320 199.970 ;
        RECT 52.595 199.650 52.915 199.970 ;
        RECT 56.190 199.650 56.510 199.970 ;
        RECT 59.785 199.650 60.105 199.970 ;
        RECT 63.380 199.650 63.700 199.970 ;
        RECT 66.975 199.650 67.295 199.970 ;
        RECT 78.720 205.550 79.040 205.870 ;
        RECT 82.315 205.550 82.635 205.870 ;
        RECT 85.910 205.550 86.230 205.870 ;
        RECT 89.505 205.550 89.825 205.870 ;
        RECT 93.100 205.550 93.420 205.870 ;
        RECT 96.695 205.550 97.015 205.870 ;
        RECT 100.290 205.550 100.610 205.870 ;
        RECT 103.885 205.550 104.205 205.870 ;
        RECT 107.480 205.550 107.800 205.870 ;
        RECT 111.075 205.550 111.395 205.870 ;
        RECT 78.720 205.150 79.040 205.470 ;
        RECT 82.315 205.150 82.635 205.470 ;
        RECT 85.910 205.150 86.230 205.470 ;
        RECT 89.505 205.150 89.825 205.470 ;
        RECT 93.100 205.150 93.420 205.470 ;
        RECT 96.695 205.150 97.015 205.470 ;
        RECT 100.290 205.150 100.610 205.470 ;
        RECT 103.885 205.150 104.205 205.470 ;
        RECT 107.480 205.150 107.800 205.470 ;
        RECT 111.075 205.150 111.395 205.470 ;
        RECT 78.720 204.750 79.040 205.070 ;
        RECT 82.315 204.750 82.635 205.070 ;
        RECT 85.910 204.750 86.230 205.070 ;
        RECT 89.505 204.750 89.825 205.070 ;
        RECT 93.100 204.750 93.420 205.070 ;
        RECT 96.695 204.750 97.015 205.070 ;
        RECT 100.290 204.750 100.610 205.070 ;
        RECT 103.885 204.750 104.205 205.070 ;
        RECT 107.480 204.750 107.800 205.070 ;
        RECT 111.075 204.750 111.395 205.070 ;
        RECT 78.720 204.350 79.040 204.670 ;
        RECT 82.315 204.350 82.635 204.670 ;
        RECT 85.910 204.350 86.230 204.670 ;
        RECT 89.505 204.350 89.825 204.670 ;
        RECT 93.100 204.350 93.420 204.670 ;
        RECT 96.695 204.350 97.015 204.670 ;
        RECT 100.290 204.350 100.610 204.670 ;
        RECT 103.885 204.350 104.205 204.670 ;
        RECT 107.480 204.350 107.800 204.670 ;
        RECT 111.075 204.350 111.395 204.670 ;
        RECT 78.720 203.950 79.040 204.270 ;
        RECT 82.315 203.950 82.635 204.270 ;
        RECT 85.910 203.950 86.230 204.270 ;
        RECT 89.505 203.950 89.825 204.270 ;
        RECT 93.100 203.950 93.420 204.270 ;
        RECT 96.695 203.950 97.015 204.270 ;
        RECT 100.290 203.950 100.610 204.270 ;
        RECT 103.885 203.950 104.205 204.270 ;
        RECT 107.480 203.950 107.800 204.270 ;
        RECT 111.075 203.950 111.395 204.270 ;
        RECT 78.720 203.550 79.040 203.870 ;
        RECT 82.315 203.550 82.635 203.870 ;
        RECT 85.910 203.550 86.230 203.870 ;
        RECT 89.505 203.550 89.825 203.870 ;
        RECT 93.100 203.550 93.420 203.870 ;
        RECT 96.695 203.550 97.015 203.870 ;
        RECT 100.290 203.550 100.610 203.870 ;
        RECT 103.885 203.550 104.205 203.870 ;
        RECT 107.480 203.550 107.800 203.870 ;
        RECT 111.075 203.550 111.395 203.870 ;
        RECT 78.720 203.150 79.040 203.470 ;
        RECT 82.315 203.150 82.635 203.470 ;
        RECT 85.910 203.150 86.230 203.470 ;
        RECT 89.505 203.150 89.825 203.470 ;
        RECT 93.100 203.150 93.420 203.470 ;
        RECT 96.695 203.150 97.015 203.470 ;
        RECT 100.290 203.150 100.610 203.470 ;
        RECT 103.885 203.150 104.205 203.470 ;
        RECT 107.480 203.150 107.800 203.470 ;
        RECT 111.075 203.150 111.395 203.470 ;
        RECT 78.720 202.050 79.040 202.370 ;
        RECT 82.315 202.050 82.635 202.370 ;
        RECT 85.910 202.050 86.230 202.370 ;
        RECT 89.505 202.050 89.825 202.370 ;
        RECT 93.100 202.050 93.420 202.370 ;
        RECT 96.695 202.050 97.015 202.370 ;
        RECT 100.290 202.050 100.610 202.370 ;
        RECT 103.885 202.050 104.205 202.370 ;
        RECT 107.480 202.050 107.800 202.370 ;
        RECT 111.075 202.050 111.395 202.370 ;
        RECT 78.720 201.650 79.040 201.970 ;
        RECT 82.315 201.650 82.635 201.970 ;
        RECT 85.910 201.650 86.230 201.970 ;
        RECT 89.505 201.650 89.825 201.970 ;
        RECT 93.100 201.650 93.420 201.970 ;
        RECT 96.695 201.650 97.015 201.970 ;
        RECT 100.290 201.650 100.610 201.970 ;
        RECT 103.885 201.650 104.205 201.970 ;
        RECT 107.480 201.650 107.800 201.970 ;
        RECT 111.075 201.650 111.395 201.970 ;
        RECT 78.720 201.250 79.040 201.570 ;
        RECT 82.315 201.250 82.635 201.570 ;
        RECT 85.910 201.250 86.230 201.570 ;
        RECT 89.505 201.250 89.825 201.570 ;
        RECT 93.100 201.250 93.420 201.570 ;
        RECT 96.695 201.250 97.015 201.570 ;
        RECT 100.290 201.250 100.610 201.570 ;
        RECT 103.885 201.250 104.205 201.570 ;
        RECT 107.480 201.250 107.800 201.570 ;
        RECT 111.075 201.250 111.395 201.570 ;
        RECT 78.720 200.850 79.040 201.170 ;
        RECT 82.315 200.850 82.635 201.170 ;
        RECT 85.910 200.850 86.230 201.170 ;
        RECT 89.505 200.850 89.825 201.170 ;
        RECT 93.100 200.850 93.420 201.170 ;
        RECT 96.695 200.850 97.015 201.170 ;
        RECT 100.290 200.850 100.610 201.170 ;
        RECT 103.885 200.850 104.205 201.170 ;
        RECT 107.480 200.850 107.800 201.170 ;
        RECT 111.075 200.850 111.395 201.170 ;
        RECT 78.720 200.450 79.040 200.770 ;
        RECT 82.315 200.450 82.635 200.770 ;
        RECT 85.910 200.450 86.230 200.770 ;
        RECT 89.505 200.450 89.825 200.770 ;
        RECT 93.100 200.450 93.420 200.770 ;
        RECT 96.695 200.450 97.015 200.770 ;
        RECT 100.290 200.450 100.610 200.770 ;
        RECT 103.885 200.450 104.205 200.770 ;
        RECT 107.480 200.450 107.800 200.770 ;
        RECT 111.075 200.450 111.395 200.770 ;
        RECT 78.720 200.050 79.040 200.370 ;
        RECT 82.315 200.050 82.635 200.370 ;
        RECT 85.910 200.050 86.230 200.370 ;
        RECT 89.505 200.050 89.825 200.370 ;
        RECT 93.100 200.050 93.420 200.370 ;
        RECT 96.695 200.050 97.015 200.370 ;
        RECT 100.290 200.050 100.610 200.370 ;
        RECT 103.885 200.050 104.205 200.370 ;
        RECT 107.480 200.050 107.800 200.370 ;
        RECT 111.075 200.050 111.395 200.370 ;
        RECT 78.720 199.650 79.040 199.970 ;
        RECT 82.315 199.650 82.635 199.970 ;
        RECT 85.910 199.650 86.230 199.970 ;
        RECT 89.505 199.650 89.825 199.970 ;
        RECT 93.100 199.650 93.420 199.970 ;
        RECT 96.695 199.650 97.015 199.970 ;
        RECT 100.290 199.650 100.610 199.970 ;
        RECT 103.885 199.650 104.205 199.970 ;
        RECT 107.480 199.650 107.800 199.970 ;
        RECT 111.075 199.650 111.395 199.970 ;
        RECT 67.690 185.950 68.010 186.270 ;
      LAYER met4 ;
        RECT 28.370 244.520 32.980 244.820 ;
        RECT 28.370 226.520 28.670 244.520 ;
        RECT 32.680 243.550 32.980 244.520 ;
        RECT 64.940 244.520 70.240 244.820 ;
        RECT 64.940 243.550 65.240 244.520 ;
        RECT 69.940 243.550 70.240 244.520 ;
        RECT 32.580 240.670 33.060 243.550 ;
        RECT 36.175 240.670 36.655 243.550 ;
        RECT 39.770 240.670 40.250 243.550 ;
        RECT 43.365 240.670 43.845 243.550 ;
        RECT 46.960 240.670 47.440 243.550 ;
        RECT 50.555 240.670 51.035 243.550 ;
        RECT 54.150 240.670 54.630 243.550 ;
        RECT 57.745 240.670 58.225 243.550 ;
        RECT 61.340 240.670 61.820 243.550 ;
        RECT 64.935 240.670 65.415 243.550 ;
        RECT 69.820 240.670 70.300 243.550 ;
        RECT 73.415 240.670 73.895 243.550 ;
        RECT 77.010 240.670 77.490 243.550 ;
        RECT 80.605 240.670 81.085 243.550 ;
        RECT 84.200 240.670 84.680 243.550 ;
        RECT 87.795 240.670 88.275 243.550 ;
        RECT 91.390 240.670 91.870 243.550 ;
        RECT 94.985 240.670 95.465 243.550 ;
        RECT 98.580 240.670 99.060 243.550 ;
        RECT 102.175 240.670 102.655 243.550 ;
        RECT 32.580 237.170 33.060 240.050 ;
        RECT 36.175 237.170 36.655 240.050 ;
        RECT 39.770 237.170 40.250 240.050 ;
        RECT 43.365 237.170 43.845 240.050 ;
        RECT 46.960 237.170 47.440 240.050 ;
        RECT 50.555 237.170 51.035 240.050 ;
        RECT 54.150 237.170 54.630 240.050 ;
        RECT 57.745 237.170 58.225 240.050 ;
        RECT 61.340 237.170 61.820 240.050 ;
        RECT 64.935 237.170 65.415 240.050 ;
        RECT 69.820 237.170 70.300 240.050 ;
        RECT 73.415 237.170 73.895 240.050 ;
        RECT 77.010 237.170 77.490 240.050 ;
        RECT 80.605 237.170 81.085 240.050 ;
        RECT 84.200 237.170 84.680 240.050 ;
        RECT 87.795 237.170 88.275 240.050 ;
        RECT 91.390 237.170 91.870 240.050 ;
        RECT 94.985 237.170 95.465 240.050 ;
        RECT 98.580 237.170 99.060 240.050 ;
        RECT 102.175 237.170 102.655 240.050 ;
        RECT 28.370 226.220 32.980 226.520 ;
        RECT 32.680 224.750 32.980 226.220 ;
        RECT 32.580 221.870 33.060 224.750 ;
        RECT 36.175 221.870 36.655 224.750 ;
        RECT 39.770 221.870 40.250 224.750 ;
        RECT 43.365 221.870 43.845 224.750 ;
        RECT 46.960 221.870 47.440 224.750 ;
        RECT 50.555 221.870 51.035 224.750 ;
        RECT 54.150 221.870 54.630 224.750 ;
        RECT 57.745 221.870 58.225 224.750 ;
        RECT 61.340 221.870 61.820 224.750 ;
        RECT 64.935 221.870 65.415 224.750 ;
        RECT 32.580 218.370 33.060 221.250 ;
        RECT 36.175 218.370 36.655 221.250 ;
        RECT 39.770 218.370 40.250 221.250 ;
        RECT 43.365 218.370 43.845 221.250 ;
        RECT 46.960 218.370 47.440 221.250 ;
        RECT 50.555 218.370 51.035 221.250 ;
        RECT 54.150 218.370 54.630 221.250 ;
        RECT 57.745 218.370 58.225 221.250 ;
        RECT 61.340 218.370 61.820 221.250 ;
        RECT 64.935 219.200 65.415 221.250 ;
        RECT 66.995 219.200 67.325 219.215 ;
        RECT 64.935 218.900 67.325 219.200 ;
        RECT 64.935 218.370 65.415 218.900 ;
        RECT 66.995 218.885 67.325 218.900 ;
        RECT 34.565 206.685 34.895 207.015 ;
        RECT 34.580 205.950 34.880 206.685 ;
        RECT 67.010 205.950 67.310 218.885 ;
        RECT 111.155 206.685 111.485 207.015 ;
        RECT 111.170 205.950 111.470 206.685 ;
        RECT 34.540 203.070 35.020 205.950 ;
        RECT 38.135 203.070 38.615 205.950 ;
        RECT 41.730 203.070 42.210 205.950 ;
        RECT 45.325 203.070 45.805 205.950 ;
        RECT 48.920 203.070 49.400 205.950 ;
        RECT 52.515 203.070 52.995 205.950 ;
        RECT 56.110 203.070 56.590 205.950 ;
        RECT 59.705 203.070 60.185 205.950 ;
        RECT 63.300 203.070 63.780 205.950 ;
        RECT 66.895 203.070 67.375 205.950 ;
        RECT 78.640 203.070 79.120 205.950 ;
        RECT 82.235 203.070 82.715 205.950 ;
        RECT 85.830 203.070 86.310 205.950 ;
        RECT 89.425 203.070 89.905 205.950 ;
        RECT 93.020 203.070 93.500 205.950 ;
        RECT 96.615 203.070 97.095 205.950 ;
        RECT 100.210 203.070 100.690 205.950 ;
        RECT 103.805 203.070 104.285 205.950 ;
        RECT 107.400 203.070 107.880 205.950 ;
        RECT 110.995 203.070 111.475 205.950 ;
        RECT 34.540 199.570 35.020 202.450 ;
        RECT 38.135 199.570 38.615 202.450 ;
        RECT 41.730 199.570 42.210 202.450 ;
        RECT 45.325 199.570 45.805 202.450 ;
        RECT 48.920 199.570 49.400 202.450 ;
        RECT 52.515 199.570 52.995 202.450 ;
        RECT 56.110 199.570 56.590 202.450 ;
        RECT 59.705 199.570 60.185 202.450 ;
        RECT 63.300 199.570 63.780 202.450 ;
        RECT 66.895 199.680 67.375 202.450 ;
        RECT 66.895 199.570 68.000 199.680 ;
        RECT 78.640 199.570 79.120 202.450 ;
        RECT 82.235 199.570 82.715 202.450 ;
        RECT 85.830 199.570 86.310 202.450 ;
        RECT 89.425 199.570 89.905 202.450 ;
        RECT 93.020 199.570 93.500 202.450 ;
        RECT 96.615 199.570 97.095 202.450 ;
        RECT 100.210 199.570 100.690 202.450 ;
        RECT 103.805 199.570 104.285 202.450 ;
        RECT 107.400 199.570 107.880 202.450 ;
        RECT 110.995 199.570 111.475 202.450 ;
        RECT 67.010 199.380 68.000 199.570 ;
        RECT 67.700 186.275 68.000 199.380 ;
        RECT 67.685 185.945 68.015 186.275 ;
    END
  END va
  PIN vb
    ANTENNAGATEAREA 72.000000 ;
    ANTENNADIFFAREA 57.985500 ;
    PORT
      LAYER li1 ;
        RECT 124.385 236.710 124.555 243.605 ;
        RECT 128.965 236.710 129.135 243.605 ;
        RECT 133.545 236.710 133.715 243.605 ;
        RECT 138.125 236.710 138.295 243.605 ;
        RECT 142.705 236.710 142.875 243.605 ;
        RECT 147.285 236.710 147.455 243.605 ;
        RECT 151.865 236.710 152.035 243.605 ;
        RECT 156.445 236.710 156.615 243.605 ;
        RECT 161.025 236.710 161.195 243.605 ;
        RECT 165.605 236.710 165.775 243.605 ;
        RECT 170.185 236.710 170.355 243.605 ;
        RECT 174.765 236.710 174.935 243.605 ;
        RECT 179.345 236.710 179.515 243.605 ;
        RECT 183.925 236.710 184.095 243.605 ;
        RECT 188.505 236.710 188.675 243.605 ;
        RECT 193.085 236.710 193.255 243.605 ;
        RECT 197.665 236.710 197.835 243.605 ;
        RECT 202.245 236.710 202.415 243.605 ;
        RECT 206.825 236.710 206.995 243.605 ;
        RECT 211.405 236.710 211.575 243.605 ;
        RECT 215.985 236.710 216.155 243.605 ;
        RECT 220.565 236.710 220.735 243.605 ;
        RECT 225.145 236.710 225.315 243.605 ;
        RECT 229.725 236.710 229.895 243.605 ;
        RECT 234.305 236.710 234.475 243.605 ;
        RECT 238.885 236.710 239.055 243.605 ;
        RECT 243.465 236.710 243.635 243.605 ;
        RECT 248.045 236.710 248.215 243.605 ;
        RECT 252.625 236.710 252.795 243.605 ;
        RECT 257.205 236.710 257.375 243.605 ;
        RECT 261.785 236.710 261.955 243.605 ;
        RECT 124.150 236.410 262.190 236.710 ;
        RECT 186.780 199.495 207.280 199.580 ;
        RECT 186.780 199.325 207.315 199.495 ;
        RECT 186.780 199.280 207.280 199.325 ;
        RECT 228.130 123.135 230.290 125.985 ;
        RECT 241.850 109.135 244.010 111.985 ;
      LAYER mcon ;
        RECT 124.385 243.335 124.555 243.505 ;
        RECT 124.385 242.975 124.555 243.145 ;
        RECT 124.385 242.615 124.555 242.785 ;
        RECT 124.385 242.255 124.555 242.425 ;
        RECT 124.385 241.895 124.555 242.065 ;
        RECT 124.385 241.535 124.555 241.705 ;
        RECT 124.385 241.175 124.555 241.345 ;
        RECT 124.385 240.815 124.555 240.985 ;
        RECT 124.385 240.455 124.555 240.625 ;
        RECT 124.385 240.095 124.555 240.265 ;
        RECT 124.385 239.735 124.555 239.905 ;
        RECT 124.385 239.375 124.555 239.545 ;
        RECT 124.385 239.015 124.555 239.185 ;
        RECT 124.385 238.655 124.555 238.825 ;
        RECT 124.385 238.295 124.555 238.465 ;
        RECT 124.385 237.935 124.555 238.105 ;
        RECT 124.385 237.575 124.555 237.745 ;
        RECT 124.385 237.215 124.555 237.385 ;
        RECT 128.965 243.335 129.135 243.505 ;
        RECT 128.965 242.975 129.135 243.145 ;
        RECT 128.965 242.615 129.135 242.785 ;
        RECT 128.965 242.255 129.135 242.425 ;
        RECT 128.965 241.895 129.135 242.065 ;
        RECT 128.965 241.535 129.135 241.705 ;
        RECT 128.965 241.175 129.135 241.345 ;
        RECT 128.965 240.815 129.135 240.985 ;
        RECT 128.965 240.455 129.135 240.625 ;
        RECT 128.965 240.095 129.135 240.265 ;
        RECT 128.965 239.735 129.135 239.905 ;
        RECT 128.965 239.375 129.135 239.545 ;
        RECT 128.965 239.015 129.135 239.185 ;
        RECT 128.965 238.655 129.135 238.825 ;
        RECT 128.965 238.295 129.135 238.465 ;
        RECT 128.965 237.935 129.135 238.105 ;
        RECT 128.965 237.575 129.135 237.745 ;
        RECT 128.965 237.215 129.135 237.385 ;
        RECT 133.545 243.335 133.715 243.505 ;
        RECT 133.545 242.975 133.715 243.145 ;
        RECT 133.545 242.615 133.715 242.785 ;
        RECT 133.545 242.255 133.715 242.425 ;
        RECT 133.545 241.895 133.715 242.065 ;
        RECT 133.545 241.535 133.715 241.705 ;
        RECT 133.545 241.175 133.715 241.345 ;
        RECT 133.545 240.815 133.715 240.985 ;
        RECT 133.545 240.455 133.715 240.625 ;
        RECT 133.545 240.095 133.715 240.265 ;
        RECT 133.545 239.735 133.715 239.905 ;
        RECT 133.545 239.375 133.715 239.545 ;
        RECT 133.545 239.015 133.715 239.185 ;
        RECT 133.545 238.655 133.715 238.825 ;
        RECT 133.545 238.295 133.715 238.465 ;
        RECT 133.545 237.935 133.715 238.105 ;
        RECT 133.545 237.575 133.715 237.745 ;
        RECT 133.545 237.215 133.715 237.385 ;
        RECT 138.125 243.335 138.295 243.505 ;
        RECT 138.125 242.975 138.295 243.145 ;
        RECT 138.125 242.615 138.295 242.785 ;
        RECT 138.125 242.255 138.295 242.425 ;
        RECT 138.125 241.895 138.295 242.065 ;
        RECT 138.125 241.535 138.295 241.705 ;
        RECT 138.125 241.175 138.295 241.345 ;
        RECT 138.125 240.815 138.295 240.985 ;
        RECT 138.125 240.455 138.295 240.625 ;
        RECT 138.125 240.095 138.295 240.265 ;
        RECT 138.125 239.735 138.295 239.905 ;
        RECT 138.125 239.375 138.295 239.545 ;
        RECT 138.125 239.015 138.295 239.185 ;
        RECT 138.125 238.655 138.295 238.825 ;
        RECT 138.125 238.295 138.295 238.465 ;
        RECT 138.125 237.935 138.295 238.105 ;
        RECT 138.125 237.575 138.295 237.745 ;
        RECT 138.125 237.215 138.295 237.385 ;
        RECT 142.705 243.335 142.875 243.505 ;
        RECT 142.705 242.975 142.875 243.145 ;
        RECT 142.705 242.615 142.875 242.785 ;
        RECT 142.705 242.255 142.875 242.425 ;
        RECT 142.705 241.895 142.875 242.065 ;
        RECT 142.705 241.535 142.875 241.705 ;
        RECT 142.705 241.175 142.875 241.345 ;
        RECT 142.705 240.815 142.875 240.985 ;
        RECT 142.705 240.455 142.875 240.625 ;
        RECT 142.705 240.095 142.875 240.265 ;
        RECT 142.705 239.735 142.875 239.905 ;
        RECT 142.705 239.375 142.875 239.545 ;
        RECT 142.705 239.015 142.875 239.185 ;
        RECT 142.705 238.655 142.875 238.825 ;
        RECT 142.705 238.295 142.875 238.465 ;
        RECT 142.705 237.935 142.875 238.105 ;
        RECT 142.705 237.575 142.875 237.745 ;
        RECT 142.705 237.215 142.875 237.385 ;
        RECT 147.285 243.335 147.455 243.505 ;
        RECT 147.285 242.975 147.455 243.145 ;
        RECT 147.285 242.615 147.455 242.785 ;
        RECT 147.285 242.255 147.455 242.425 ;
        RECT 147.285 241.895 147.455 242.065 ;
        RECT 147.285 241.535 147.455 241.705 ;
        RECT 147.285 241.175 147.455 241.345 ;
        RECT 147.285 240.815 147.455 240.985 ;
        RECT 147.285 240.455 147.455 240.625 ;
        RECT 147.285 240.095 147.455 240.265 ;
        RECT 147.285 239.735 147.455 239.905 ;
        RECT 147.285 239.375 147.455 239.545 ;
        RECT 147.285 239.015 147.455 239.185 ;
        RECT 147.285 238.655 147.455 238.825 ;
        RECT 147.285 238.295 147.455 238.465 ;
        RECT 147.285 237.935 147.455 238.105 ;
        RECT 147.285 237.575 147.455 237.745 ;
        RECT 147.285 237.215 147.455 237.385 ;
        RECT 151.865 243.335 152.035 243.505 ;
        RECT 151.865 242.975 152.035 243.145 ;
        RECT 151.865 242.615 152.035 242.785 ;
        RECT 151.865 242.255 152.035 242.425 ;
        RECT 151.865 241.895 152.035 242.065 ;
        RECT 151.865 241.535 152.035 241.705 ;
        RECT 151.865 241.175 152.035 241.345 ;
        RECT 151.865 240.815 152.035 240.985 ;
        RECT 151.865 240.455 152.035 240.625 ;
        RECT 151.865 240.095 152.035 240.265 ;
        RECT 151.865 239.735 152.035 239.905 ;
        RECT 151.865 239.375 152.035 239.545 ;
        RECT 151.865 239.015 152.035 239.185 ;
        RECT 151.865 238.655 152.035 238.825 ;
        RECT 151.865 238.295 152.035 238.465 ;
        RECT 151.865 237.935 152.035 238.105 ;
        RECT 151.865 237.575 152.035 237.745 ;
        RECT 151.865 237.215 152.035 237.385 ;
        RECT 156.445 243.335 156.615 243.505 ;
        RECT 156.445 242.975 156.615 243.145 ;
        RECT 156.445 242.615 156.615 242.785 ;
        RECT 156.445 242.255 156.615 242.425 ;
        RECT 156.445 241.895 156.615 242.065 ;
        RECT 156.445 241.535 156.615 241.705 ;
        RECT 156.445 241.175 156.615 241.345 ;
        RECT 156.445 240.815 156.615 240.985 ;
        RECT 156.445 240.455 156.615 240.625 ;
        RECT 156.445 240.095 156.615 240.265 ;
        RECT 156.445 239.735 156.615 239.905 ;
        RECT 156.445 239.375 156.615 239.545 ;
        RECT 156.445 239.015 156.615 239.185 ;
        RECT 156.445 238.655 156.615 238.825 ;
        RECT 156.445 238.295 156.615 238.465 ;
        RECT 156.445 237.935 156.615 238.105 ;
        RECT 156.445 237.575 156.615 237.745 ;
        RECT 156.445 237.215 156.615 237.385 ;
        RECT 161.025 243.335 161.195 243.505 ;
        RECT 161.025 242.975 161.195 243.145 ;
        RECT 161.025 242.615 161.195 242.785 ;
        RECT 161.025 242.255 161.195 242.425 ;
        RECT 161.025 241.895 161.195 242.065 ;
        RECT 161.025 241.535 161.195 241.705 ;
        RECT 161.025 241.175 161.195 241.345 ;
        RECT 161.025 240.815 161.195 240.985 ;
        RECT 161.025 240.455 161.195 240.625 ;
        RECT 161.025 240.095 161.195 240.265 ;
        RECT 161.025 239.735 161.195 239.905 ;
        RECT 161.025 239.375 161.195 239.545 ;
        RECT 161.025 239.015 161.195 239.185 ;
        RECT 161.025 238.655 161.195 238.825 ;
        RECT 161.025 238.295 161.195 238.465 ;
        RECT 161.025 237.935 161.195 238.105 ;
        RECT 161.025 237.575 161.195 237.745 ;
        RECT 161.025 237.215 161.195 237.385 ;
        RECT 165.605 243.335 165.775 243.505 ;
        RECT 165.605 242.975 165.775 243.145 ;
        RECT 165.605 242.615 165.775 242.785 ;
        RECT 165.605 242.255 165.775 242.425 ;
        RECT 165.605 241.895 165.775 242.065 ;
        RECT 165.605 241.535 165.775 241.705 ;
        RECT 165.605 241.175 165.775 241.345 ;
        RECT 165.605 240.815 165.775 240.985 ;
        RECT 165.605 240.455 165.775 240.625 ;
        RECT 165.605 240.095 165.775 240.265 ;
        RECT 165.605 239.735 165.775 239.905 ;
        RECT 165.605 239.375 165.775 239.545 ;
        RECT 165.605 239.015 165.775 239.185 ;
        RECT 165.605 238.655 165.775 238.825 ;
        RECT 165.605 238.295 165.775 238.465 ;
        RECT 165.605 237.935 165.775 238.105 ;
        RECT 165.605 237.575 165.775 237.745 ;
        RECT 165.605 237.215 165.775 237.385 ;
        RECT 170.185 243.335 170.355 243.505 ;
        RECT 170.185 242.975 170.355 243.145 ;
        RECT 170.185 242.615 170.355 242.785 ;
        RECT 170.185 242.255 170.355 242.425 ;
        RECT 170.185 241.895 170.355 242.065 ;
        RECT 170.185 241.535 170.355 241.705 ;
        RECT 170.185 241.175 170.355 241.345 ;
        RECT 170.185 240.815 170.355 240.985 ;
        RECT 170.185 240.455 170.355 240.625 ;
        RECT 170.185 240.095 170.355 240.265 ;
        RECT 170.185 239.735 170.355 239.905 ;
        RECT 170.185 239.375 170.355 239.545 ;
        RECT 170.185 239.015 170.355 239.185 ;
        RECT 170.185 238.655 170.355 238.825 ;
        RECT 170.185 238.295 170.355 238.465 ;
        RECT 170.185 237.935 170.355 238.105 ;
        RECT 170.185 237.575 170.355 237.745 ;
        RECT 170.185 237.215 170.355 237.385 ;
        RECT 174.765 243.335 174.935 243.505 ;
        RECT 174.765 242.975 174.935 243.145 ;
        RECT 174.765 242.615 174.935 242.785 ;
        RECT 174.765 242.255 174.935 242.425 ;
        RECT 174.765 241.895 174.935 242.065 ;
        RECT 174.765 241.535 174.935 241.705 ;
        RECT 174.765 241.175 174.935 241.345 ;
        RECT 174.765 240.815 174.935 240.985 ;
        RECT 174.765 240.455 174.935 240.625 ;
        RECT 174.765 240.095 174.935 240.265 ;
        RECT 174.765 239.735 174.935 239.905 ;
        RECT 174.765 239.375 174.935 239.545 ;
        RECT 174.765 239.015 174.935 239.185 ;
        RECT 174.765 238.655 174.935 238.825 ;
        RECT 174.765 238.295 174.935 238.465 ;
        RECT 174.765 237.935 174.935 238.105 ;
        RECT 174.765 237.575 174.935 237.745 ;
        RECT 174.765 237.215 174.935 237.385 ;
        RECT 179.345 243.335 179.515 243.505 ;
        RECT 179.345 242.975 179.515 243.145 ;
        RECT 179.345 242.615 179.515 242.785 ;
        RECT 179.345 242.255 179.515 242.425 ;
        RECT 179.345 241.895 179.515 242.065 ;
        RECT 179.345 241.535 179.515 241.705 ;
        RECT 179.345 241.175 179.515 241.345 ;
        RECT 179.345 240.815 179.515 240.985 ;
        RECT 179.345 240.455 179.515 240.625 ;
        RECT 179.345 240.095 179.515 240.265 ;
        RECT 179.345 239.735 179.515 239.905 ;
        RECT 179.345 239.375 179.515 239.545 ;
        RECT 179.345 239.015 179.515 239.185 ;
        RECT 179.345 238.655 179.515 238.825 ;
        RECT 179.345 238.295 179.515 238.465 ;
        RECT 179.345 237.935 179.515 238.105 ;
        RECT 179.345 237.575 179.515 237.745 ;
        RECT 179.345 237.215 179.515 237.385 ;
        RECT 183.925 243.335 184.095 243.505 ;
        RECT 183.925 242.975 184.095 243.145 ;
        RECT 183.925 242.615 184.095 242.785 ;
        RECT 183.925 242.255 184.095 242.425 ;
        RECT 183.925 241.895 184.095 242.065 ;
        RECT 183.925 241.535 184.095 241.705 ;
        RECT 183.925 241.175 184.095 241.345 ;
        RECT 183.925 240.815 184.095 240.985 ;
        RECT 183.925 240.455 184.095 240.625 ;
        RECT 183.925 240.095 184.095 240.265 ;
        RECT 183.925 239.735 184.095 239.905 ;
        RECT 183.925 239.375 184.095 239.545 ;
        RECT 183.925 239.015 184.095 239.185 ;
        RECT 183.925 238.655 184.095 238.825 ;
        RECT 183.925 238.295 184.095 238.465 ;
        RECT 183.925 237.935 184.095 238.105 ;
        RECT 183.925 237.575 184.095 237.745 ;
        RECT 183.925 237.215 184.095 237.385 ;
        RECT 188.505 243.335 188.675 243.505 ;
        RECT 188.505 242.975 188.675 243.145 ;
        RECT 188.505 242.615 188.675 242.785 ;
        RECT 188.505 242.255 188.675 242.425 ;
        RECT 188.505 241.895 188.675 242.065 ;
        RECT 188.505 241.535 188.675 241.705 ;
        RECT 188.505 241.175 188.675 241.345 ;
        RECT 188.505 240.815 188.675 240.985 ;
        RECT 188.505 240.455 188.675 240.625 ;
        RECT 188.505 240.095 188.675 240.265 ;
        RECT 188.505 239.735 188.675 239.905 ;
        RECT 188.505 239.375 188.675 239.545 ;
        RECT 188.505 239.015 188.675 239.185 ;
        RECT 188.505 238.655 188.675 238.825 ;
        RECT 188.505 238.295 188.675 238.465 ;
        RECT 188.505 237.935 188.675 238.105 ;
        RECT 188.505 237.575 188.675 237.745 ;
        RECT 188.505 237.215 188.675 237.385 ;
        RECT 193.085 243.335 193.255 243.505 ;
        RECT 193.085 242.975 193.255 243.145 ;
        RECT 193.085 242.615 193.255 242.785 ;
        RECT 193.085 242.255 193.255 242.425 ;
        RECT 193.085 241.895 193.255 242.065 ;
        RECT 193.085 241.535 193.255 241.705 ;
        RECT 193.085 241.175 193.255 241.345 ;
        RECT 193.085 240.815 193.255 240.985 ;
        RECT 193.085 240.455 193.255 240.625 ;
        RECT 193.085 240.095 193.255 240.265 ;
        RECT 193.085 239.735 193.255 239.905 ;
        RECT 193.085 239.375 193.255 239.545 ;
        RECT 193.085 239.015 193.255 239.185 ;
        RECT 193.085 238.655 193.255 238.825 ;
        RECT 193.085 238.295 193.255 238.465 ;
        RECT 193.085 237.935 193.255 238.105 ;
        RECT 193.085 237.575 193.255 237.745 ;
        RECT 193.085 237.215 193.255 237.385 ;
        RECT 197.665 243.335 197.835 243.505 ;
        RECT 197.665 242.975 197.835 243.145 ;
        RECT 197.665 242.615 197.835 242.785 ;
        RECT 197.665 242.255 197.835 242.425 ;
        RECT 197.665 241.895 197.835 242.065 ;
        RECT 197.665 241.535 197.835 241.705 ;
        RECT 197.665 241.175 197.835 241.345 ;
        RECT 197.665 240.815 197.835 240.985 ;
        RECT 197.665 240.455 197.835 240.625 ;
        RECT 197.665 240.095 197.835 240.265 ;
        RECT 197.665 239.735 197.835 239.905 ;
        RECT 197.665 239.375 197.835 239.545 ;
        RECT 197.665 239.015 197.835 239.185 ;
        RECT 197.665 238.655 197.835 238.825 ;
        RECT 197.665 238.295 197.835 238.465 ;
        RECT 197.665 237.935 197.835 238.105 ;
        RECT 197.665 237.575 197.835 237.745 ;
        RECT 197.665 237.215 197.835 237.385 ;
        RECT 202.245 243.335 202.415 243.505 ;
        RECT 202.245 242.975 202.415 243.145 ;
        RECT 202.245 242.615 202.415 242.785 ;
        RECT 202.245 242.255 202.415 242.425 ;
        RECT 202.245 241.895 202.415 242.065 ;
        RECT 202.245 241.535 202.415 241.705 ;
        RECT 202.245 241.175 202.415 241.345 ;
        RECT 202.245 240.815 202.415 240.985 ;
        RECT 202.245 240.455 202.415 240.625 ;
        RECT 202.245 240.095 202.415 240.265 ;
        RECT 202.245 239.735 202.415 239.905 ;
        RECT 202.245 239.375 202.415 239.545 ;
        RECT 202.245 239.015 202.415 239.185 ;
        RECT 202.245 238.655 202.415 238.825 ;
        RECT 202.245 238.295 202.415 238.465 ;
        RECT 202.245 237.935 202.415 238.105 ;
        RECT 202.245 237.575 202.415 237.745 ;
        RECT 202.245 237.215 202.415 237.385 ;
        RECT 206.825 243.335 206.995 243.505 ;
        RECT 206.825 242.975 206.995 243.145 ;
        RECT 206.825 242.615 206.995 242.785 ;
        RECT 206.825 242.255 206.995 242.425 ;
        RECT 206.825 241.895 206.995 242.065 ;
        RECT 206.825 241.535 206.995 241.705 ;
        RECT 206.825 241.175 206.995 241.345 ;
        RECT 206.825 240.815 206.995 240.985 ;
        RECT 206.825 240.455 206.995 240.625 ;
        RECT 206.825 240.095 206.995 240.265 ;
        RECT 206.825 239.735 206.995 239.905 ;
        RECT 206.825 239.375 206.995 239.545 ;
        RECT 206.825 239.015 206.995 239.185 ;
        RECT 206.825 238.655 206.995 238.825 ;
        RECT 206.825 238.295 206.995 238.465 ;
        RECT 206.825 237.935 206.995 238.105 ;
        RECT 206.825 237.575 206.995 237.745 ;
        RECT 206.825 237.215 206.995 237.385 ;
        RECT 211.405 243.335 211.575 243.505 ;
        RECT 211.405 242.975 211.575 243.145 ;
        RECT 211.405 242.615 211.575 242.785 ;
        RECT 211.405 242.255 211.575 242.425 ;
        RECT 211.405 241.895 211.575 242.065 ;
        RECT 211.405 241.535 211.575 241.705 ;
        RECT 211.405 241.175 211.575 241.345 ;
        RECT 211.405 240.815 211.575 240.985 ;
        RECT 211.405 240.455 211.575 240.625 ;
        RECT 211.405 240.095 211.575 240.265 ;
        RECT 211.405 239.735 211.575 239.905 ;
        RECT 211.405 239.375 211.575 239.545 ;
        RECT 211.405 239.015 211.575 239.185 ;
        RECT 211.405 238.655 211.575 238.825 ;
        RECT 211.405 238.295 211.575 238.465 ;
        RECT 211.405 237.935 211.575 238.105 ;
        RECT 211.405 237.575 211.575 237.745 ;
        RECT 211.405 237.215 211.575 237.385 ;
        RECT 215.985 243.335 216.155 243.505 ;
        RECT 215.985 242.975 216.155 243.145 ;
        RECT 215.985 242.615 216.155 242.785 ;
        RECT 215.985 242.255 216.155 242.425 ;
        RECT 215.985 241.895 216.155 242.065 ;
        RECT 215.985 241.535 216.155 241.705 ;
        RECT 215.985 241.175 216.155 241.345 ;
        RECT 215.985 240.815 216.155 240.985 ;
        RECT 215.985 240.455 216.155 240.625 ;
        RECT 215.985 240.095 216.155 240.265 ;
        RECT 215.985 239.735 216.155 239.905 ;
        RECT 215.985 239.375 216.155 239.545 ;
        RECT 215.985 239.015 216.155 239.185 ;
        RECT 215.985 238.655 216.155 238.825 ;
        RECT 215.985 238.295 216.155 238.465 ;
        RECT 215.985 237.935 216.155 238.105 ;
        RECT 215.985 237.575 216.155 237.745 ;
        RECT 215.985 237.215 216.155 237.385 ;
        RECT 220.565 243.335 220.735 243.505 ;
        RECT 220.565 242.975 220.735 243.145 ;
        RECT 220.565 242.615 220.735 242.785 ;
        RECT 220.565 242.255 220.735 242.425 ;
        RECT 220.565 241.895 220.735 242.065 ;
        RECT 220.565 241.535 220.735 241.705 ;
        RECT 220.565 241.175 220.735 241.345 ;
        RECT 220.565 240.815 220.735 240.985 ;
        RECT 220.565 240.455 220.735 240.625 ;
        RECT 220.565 240.095 220.735 240.265 ;
        RECT 220.565 239.735 220.735 239.905 ;
        RECT 220.565 239.375 220.735 239.545 ;
        RECT 220.565 239.015 220.735 239.185 ;
        RECT 220.565 238.655 220.735 238.825 ;
        RECT 220.565 238.295 220.735 238.465 ;
        RECT 220.565 237.935 220.735 238.105 ;
        RECT 220.565 237.575 220.735 237.745 ;
        RECT 220.565 237.215 220.735 237.385 ;
        RECT 225.145 243.335 225.315 243.505 ;
        RECT 225.145 242.975 225.315 243.145 ;
        RECT 225.145 242.615 225.315 242.785 ;
        RECT 225.145 242.255 225.315 242.425 ;
        RECT 225.145 241.895 225.315 242.065 ;
        RECT 225.145 241.535 225.315 241.705 ;
        RECT 225.145 241.175 225.315 241.345 ;
        RECT 225.145 240.815 225.315 240.985 ;
        RECT 225.145 240.455 225.315 240.625 ;
        RECT 225.145 240.095 225.315 240.265 ;
        RECT 225.145 239.735 225.315 239.905 ;
        RECT 225.145 239.375 225.315 239.545 ;
        RECT 225.145 239.015 225.315 239.185 ;
        RECT 225.145 238.655 225.315 238.825 ;
        RECT 225.145 238.295 225.315 238.465 ;
        RECT 225.145 237.935 225.315 238.105 ;
        RECT 225.145 237.575 225.315 237.745 ;
        RECT 225.145 237.215 225.315 237.385 ;
        RECT 229.725 243.335 229.895 243.505 ;
        RECT 229.725 242.975 229.895 243.145 ;
        RECT 229.725 242.615 229.895 242.785 ;
        RECT 229.725 242.255 229.895 242.425 ;
        RECT 229.725 241.895 229.895 242.065 ;
        RECT 229.725 241.535 229.895 241.705 ;
        RECT 229.725 241.175 229.895 241.345 ;
        RECT 229.725 240.815 229.895 240.985 ;
        RECT 229.725 240.455 229.895 240.625 ;
        RECT 229.725 240.095 229.895 240.265 ;
        RECT 229.725 239.735 229.895 239.905 ;
        RECT 229.725 239.375 229.895 239.545 ;
        RECT 229.725 239.015 229.895 239.185 ;
        RECT 229.725 238.655 229.895 238.825 ;
        RECT 229.725 238.295 229.895 238.465 ;
        RECT 229.725 237.935 229.895 238.105 ;
        RECT 229.725 237.575 229.895 237.745 ;
        RECT 229.725 237.215 229.895 237.385 ;
        RECT 234.305 243.335 234.475 243.505 ;
        RECT 234.305 242.975 234.475 243.145 ;
        RECT 234.305 242.615 234.475 242.785 ;
        RECT 234.305 242.255 234.475 242.425 ;
        RECT 234.305 241.895 234.475 242.065 ;
        RECT 234.305 241.535 234.475 241.705 ;
        RECT 234.305 241.175 234.475 241.345 ;
        RECT 234.305 240.815 234.475 240.985 ;
        RECT 234.305 240.455 234.475 240.625 ;
        RECT 234.305 240.095 234.475 240.265 ;
        RECT 234.305 239.735 234.475 239.905 ;
        RECT 234.305 239.375 234.475 239.545 ;
        RECT 234.305 239.015 234.475 239.185 ;
        RECT 234.305 238.655 234.475 238.825 ;
        RECT 234.305 238.295 234.475 238.465 ;
        RECT 234.305 237.935 234.475 238.105 ;
        RECT 234.305 237.575 234.475 237.745 ;
        RECT 234.305 237.215 234.475 237.385 ;
        RECT 238.885 243.335 239.055 243.505 ;
        RECT 238.885 242.975 239.055 243.145 ;
        RECT 238.885 242.615 239.055 242.785 ;
        RECT 238.885 242.255 239.055 242.425 ;
        RECT 238.885 241.895 239.055 242.065 ;
        RECT 238.885 241.535 239.055 241.705 ;
        RECT 238.885 241.175 239.055 241.345 ;
        RECT 238.885 240.815 239.055 240.985 ;
        RECT 238.885 240.455 239.055 240.625 ;
        RECT 238.885 240.095 239.055 240.265 ;
        RECT 238.885 239.735 239.055 239.905 ;
        RECT 238.885 239.375 239.055 239.545 ;
        RECT 238.885 239.015 239.055 239.185 ;
        RECT 238.885 238.655 239.055 238.825 ;
        RECT 238.885 238.295 239.055 238.465 ;
        RECT 238.885 237.935 239.055 238.105 ;
        RECT 238.885 237.575 239.055 237.745 ;
        RECT 238.885 237.215 239.055 237.385 ;
        RECT 243.465 243.335 243.635 243.505 ;
        RECT 243.465 242.975 243.635 243.145 ;
        RECT 243.465 242.615 243.635 242.785 ;
        RECT 243.465 242.255 243.635 242.425 ;
        RECT 243.465 241.895 243.635 242.065 ;
        RECT 243.465 241.535 243.635 241.705 ;
        RECT 243.465 241.175 243.635 241.345 ;
        RECT 243.465 240.815 243.635 240.985 ;
        RECT 243.465 240.455 243.635 240.625 ;
        RECT 243.465 240.095 243.635 240.265 ;
        RECT 243.465 239.735 243.635 239.905 ;
        RECT 243.465 239.375 243.635 239.545 ;
        RECT 243.465 239.015 243.635 239.185 ;
        RECT 243.465 238.655 243.635 238.825 ;
        RECT 243.465 238.295 243.635 238.465 ;
        RECT 243.465 237.935 243.635 238.105 ;
        RECT 243.465 237.575 243.635 237.745 ;
        RECT 243.465 237.215 243.635 237.385 ;
        RECT 248.045 243.335 248.215 243.505 ;
        RECT 248.045 242.975 248.215 243.145 ;
        RECT 248.045 242.615 248.215 242.785 ;
        RECT 248.045 242.255 248.215 242.425 ;
        RECT 248.045 241.895 248.215 242.065 ;
        RECT 248.045 241.535 248.215 241.705 ;
        RECT 248.045 241.175 248.215 241.345 ;
        RECT 248.045 240.815 248.215 240.985 ;
        RECT 248.045 240.455 248.215 240.625 ;
        RECT 248.045 240.095 248.215 240.265 ;
        RECT 248.045 239.735 248.215 239.905 ;
        RECT 248.045 239.375 248.215 239.545 ;
        RECT 248.045 239.015 248.215 239.185 ;
        RECT 248.045 238.655 248.215 238.825 ;
        RECT 248.045 238.295 248.215 238.465 ;
        RECT 248.045 237.935 248.215 238.105 ;
        RECT 248.045 237.575 248.215 237.745 ;
        RECT 248.045 237.215 248.215 237.385 ;
        RECT 252.625 243.335 252.795 243.505 ;
        RECT 252.625 242.975 252.795 243.145 ;
        RECT 252.625 242.615 252.795 242.785 ;
        RECT 252.625 242.255 252.795 242.425 ;
        RECT 252.625 241.895 252.795 242.065 ;
        RECT 252.625 241.535 252.795 241.705 ;
        RECT 252.625 241.175 252.795 241.345 ;
        RECT 252.625 240.815 252.795 240.985 ;
        RECT 252.625 240.455 252.795 240.625 ;
        RECT 252.625 240.095 252.795 240.265 ;
        RECT 252.625 239.735 252.795 239.905 ;
        RECT 252.625 239.375 252.795 239.545 ;
        RECT 252.625 239.015 252.795 239.185 ;
        RECT 252.625 238.655 252.795 238.825 ;
        RECT 252.625 238.295 252.795 238.465 ;
        RECT 252.625 237.935 252.795 238.105 ;
        RECT 252.625 237.575 252.795 237.745 ;
        RECT 252.625 237.215 252.795 237.385 ;
        RECT 257.205 243.335 257.375 243.505 ;
        RECT 257.205 242.975 257.375 243.145 ;
        RECT 257.205 242.615 257.375 242.785 ;
        RECT 257.205 242.255 257.375 242.425 ;
        RECT 257.205 241.895 257.375 242.065 ;
        RECT 257.205 241.535 257.375 241.705 ;
        RECT 257.205 241.175 257.375 241.345 ;
        RECT 257.205 240.815 257.375 240.985 ;
        RECT 257.205 240.455 257.375 240.625 ;
        RECT 257.205 240.095 257.375 240.265 ;
        RECT 257.205 239.735 257.375 239.905 ;
        RECT 257.205 239.375 257.375 239.545 ;
        RECT 257.205 239.015 257.375 239.185 ;
        RECT 257.205 238.655 257.375 238.825 ;
        RECT 257.205 238.295 257.375 238.465 ;
        RECT 257.205 237.935 257.375 238.105 ;
        RECT 257.205 237.575 257.375 237.745 ;
        RECT 257.205 237.215 257.375 237.385 ;
        RECT 261.785 243.335 261.955 243.505 ;
        RECT 261.785 242.975 261.955 243.145 ;
        RECT 261.785 242.615 261.955 242.785 ;
        RECT 261.785 242.255 261.955 242.425 ;
        RECT 261.785 241.895 261.955 242.065 ;
        RECT 261.785 241.535 261.955 241.705 ;
        RECT 261.785 241.175 261.955 241.345 ;
        RECT 261.785 240.815 261.955 240.985 ;
        RECT 261.785 240.455 261.955 240.625 ;
        RECT 261.785 240.095 261.955 240.265 ;
        RECT 261.785 239.735 261.955 239.905 ;
        RECT 261.785 239.375 261.955 239.545 ;
        RECT 261.785 239.015 261.955 239.185 ;
        RECT 261.785 238.655 261.955 238.825 ;
        RECT 261.785 238.295 261.955 238.465 ;
        RECT 261.785 237.935 261.955 238.105 ;
        RECT 261.785 237.575 261.955 237.745 ;
        RECT 261.785 237.215 261.955 237.385 ;
        RECT 207.145 199.325 207.315 199.495 ;
        RECT 228.225 123.215 230.195 125.905 ;
        RECT 241.945 109.215 243.915 111.905 ;
      LAYER met1 ;
        RECT 124.355 237.135 124.585 243.585 ;
        RECT 128.935 237.135 129.165 243.585 ;
        RECT 133.515 237.135 133.745 243.585 ;
        RECT 138.095 237.135 138.325 243.585 ;
        RECT 142.675 237.135 142.905 243.585 ;
        RECT 147.255 237.135 147.485 243.585 ;
        RECT 151.835 237.135 152.065 243.585 ;
        RECT 156.415 237.135 156.645 243.585 ;
        RECT 160.995 237.135 161.225 243.585 ;
        RECT 165.575 237.135 165.805 243.585 ;
        RECT 170.155 237.135 170.385 243.585 ;
        RECT 174.735 237.135 174.965 243.585 ;
        RECT 179.315 237.135 179.545 243.585 ;
        RECT 183.895 237.135 184.125 243.585 ;
        RECT 188.475 237.135 188.705 243.585 ;
        RECT 193.055 237.135 193.285 243.585 ;
        RECT 197.635 237.135 197.865 243.585 ;
        RECT 202.215 237.135 202.445 243.585 ;
        RECT 206.795 237.135 207.025 243.585 ;
        RECT 211.375 237.135 211.605 243.585 ;
        RECT 215.955 237.135 216.185 243.585 ;
        RECT 220.535 237.135 220.765 243.585 ;
        RECT 225.115 237.135 225.345 243.585 ;
        RECT 229.695 237.135 229.925 243.585 ;
        RECT 234.275 237.135 234.505 243.585 ;
        RECT 238.855 237.135 239.085 243.585 ;
        RECT 241.570 237.560 241.890 237.620 ;
        RECT 243.435 237.560 243.665 243.585 ;
        RECT 241.570 237.420 243.665 237.560 ;
        RECT 241.570 237.360 241.890 237.420 ;
        RECT 243.435 237.135 243.665 237.420 ;
        RECT 248.015 237.135 248.245 243.585 ;
        RECT 252.595 237.135 252.825 243.585 ;
        RECT 257.175 237.135 257.405 243.585 ;
        RECT 261.755 237.135 261.985 243.585 ;
        RECT 207.085 199.480 207.375 199.525 ;
        RECT 241.570 199.480 241.890 199.540 ;
        RECT 207.085 199.340 241.890 199.480 ;
        RECT 207.085 199.295 207.375 199.340 ;
        RECT 241.570 199.280 241.890 199.340 ;
        RECT 243.410 168.680 243.730 168.940 ;
        RECT 243.500 168.540 243.640 168.680 ;
        RECT 243.500 168.400 292.330 168.540 ;
        RECT 292.190 167.180 292.330 168.400 ;
        RECT 291.965 167.040 292.560 167.180 ;
        RECT 230.070 131.140 230.390 131.200 ;
        RECT 242.490 131.140 242.810 131.200 ;
        RECT 230.070 131.000 242.810 131.140 ;
        RECT 230.070 130.940 230.390 131.000 ;
        RECT 242.490 130.940 242.810 131.000 ;
        RECT 228.185 125.760 230.235 125.965 ;
        RECT 228.185 125.500 230.390 125.760 ;
        RECT 228.185 123.155 230.235 125.500 ;
        RECT 242.490 112.240 242.810 112.500 ;
        RECT 242.580 111.965 242.720 112.240 ;
        RECT 241.905 109.155 243.955 111.965 ;
      LAYER via ;
        RECT 241.600 237.360 241.860 237.620 ;
        RECT 241.600 199.280 241.860 199.540 ;
        RECT 243.440 168.680 243.700 168.940 ;
        RECT 230.100 130.940 230.360 131.200 ;
        RECT 242.520 130.940 242.780 131.200 ;
        RECT 230.100 125.500 230.360 125.760 ;
        RECT 242.520 112.240 242.780 112.500 ;
      LAYER met2 ;
        RECT 241.600 237.330 241.860 237.650 ;
        RECT 241.660 199.570 241.800 237.330 ;
        RECT 241.600 199.250 241.860 199.570 ;
        RECT 241.660 185.880 241.800 199.250 ;
        RECT 241.660 185.740 242.720 185.880 ;
        RECT 242.580 168.880 242.720 185.740 ;
        RECT 243.440 168.880 243.700 168.970 ;
        RECT 242.580 168.740 243.700 168.880 ;
        RECT 242.580 131.230 242.720 168.740 ;
        RECT 243.440 168.650 243.700 168.740 ;
        RECT 230.100 130.910 230.360 131.230 ;
        RECT 242.520 130.910 242.780 131.230 ;
        RECT 230.160 125.790 230.300 130.910 ;
        RECT 230.100 125.470 230.360 125.790 ;
        RECT 242.580 112.530 242.720 130.910 ;
        RECT 242.520 112.210 242.780 112.530 ;
    END
  END vb
  PIN vbg
    ANTENNADIFFAREA 57.985500 ;
    PORT
      LAYER li1 ;
        RECT 124.385 86.310 124.555 93.205 ;
        RECT 128.965 86.310 129.135 93.205 ;
        RECT 133.545 86.310 133.715 93.205 ;
        RECT 138.125 86.310 138.295 93.205 ;
        RECT 142.705 86.310 142.875 93.205 ;
        RECT 147.285 86.310 147.455 93.205 ;
        RECT 151.865 86.310 152.035 93.205 ;
        RECT 156.445 86.310 156.615 93.205 ;
        RECT 161.025 86.310 161.195 93.205 ;
        RECT 165.605 86.310 165.775 93.205 ;
        RECT 170.185 86.310 170.355 93.205 ;
        RECT 174.765 86.310 174.935 93.205 ;
        RECT 179.345 86.310 179.515 93.205 ;
        RECT 183.925 86.310 184.095 93.205 ;
        RECT 188.505 86.310 188.675 93.205 ;
        RECT 193.085 86.310 193.255 93.205 ;
        RECT 197.665 86.310 197.835 93.205 ;
        RECT 202.245 86.310 202.415 93.205 ;
        RECT 206.825 86.310 206.995 93.205 ;
        RECT 211.405 86.310 211.575 93.205 ;
        RECT 215.985 86.310 216.155 93.205 ;
        RECT 220.565 86.310 220.735 93.205 ;
        RECT 225.145 86.310 225.315 93.205 ;
        RECT 229.725 86.310 229.895 93.205 ;
        RECT 234.305 86.310 234.475 93.205 ;
        RECT 238.885 86.310 239.055 93.205 ;
        RECT 243.465 86.310 243.635 93.205 ;
        RECT 248.045 86.310 248.215 93.205 ;
        RECT 252.625 86.310 252.795 93.205 ;
        RECT 257.205 86.310 257.375 93.205 ;
        RECT 261.785 86.310 261.955 93.205 ;
        RECT 124.150 86.010 262.190 86.310 ;
        RECT 218.820 52.735 220.980 55.585 ;
      LAYER mcon ;
        RECT 124.385 92.935 124.555 93.105 ;
        RECT 124.385 92.575 124.555 92.745 ;
        RECT 124.385 92.215 124.555 92.385 ;
        RECT 124.385 91.855 124.555 92.025 ;
        RECT 124.385 91.495 124.555 91.665 ;
        RECT 124.385 91.135 124.555 91.305 ;
        RECT 124.385 90.775 124.555 90.945 ;
        RECT 124.385 90.415 124.555 90.585 ;
        RECT 124.385 90.055 124.555 90.225 ;
        RECT 124.385 89.695 124.555 89.865 ;
        RECT 124.385 89.335 124.555 89.505 ;
        RECT 124.385 88.975 124.555 89.145 ;
        RECT 124.385 88.615 124.555 88.785 ;
        RECT 124.385 88.255 124.555 88.425 ;
        RECT 124.385 87.895 124.555 88.065 ;
        RECT 124.385 87.535 124.555 87.705 ;
        RECT 124.385 87.175 124.555 87.345 ;
        RECT 124.385 86.815 124.555 86.985 ;
        RECT 128.965 92.935 129.135 93.105 ;
        RECT 128.965 92.575 129.135 92.745 ;
        RECT 128.965 92.215 129.135 92.385 ;
        RECT 128.965 91.855 129.135 92.025 ;
        RECT 128.965 91.495 129.135 91.665 ;
        RECT 128.965 91.135 129.135 91.305 ;
        RECT 128.965 90.775 129.135 90.945 ;
        RECT 128.965 90.415 129.135 90.585 ;
        RECT 128.965 90.055 129.135 90.225 ;
        RECT 128.965 89.695 129.135 89.865 ;
        RECT 128.965 89.335 129.135 89.505 ;
        RECT 128.965 88.975 129.135 89.145 ;
        RECT 128.965 88.615 129.135 88.785 ;
        RECT 128.965 88.255 129.135 88.425 ;
        RECT 128.965 87.895 129.135 88.065 ;
        RECT 128.965 87.535 129.135 87.705 ;
        RECT 128.965 87.175 129.135 87.345 ;
        RECT 128.965 86.815 129.135 86.985 ;
        RECT 133.545 92.935 133.715 93.105 ;
        RECT 133.545 92.575 133.715 92.745 ;
        RECT 133.545 92.215 133.715 92.385 ;
        RECT 133.545 91.855 133.715 92.025 ;
        RECT 133.545 91.495 133.715 91.665 ;
        RECT 133.545 91.135 133.715 91.305 ;
        RECT 133.545 90.775 133.715 90.945 ;
        RECT 133.545 90.415 133.715 90.585 ;
        RECT 133.545 90.055 133.715 90.225 ;
        RECT 133.545 89.695 133.715 89.865 ;
        RECT 133.545 89.335 133.715 89.505 ;
        RECT 133.545 88.975 133.715 89.145 ;
        RECT 133.545 88.615 133.715 88.785 ;
        RECT 133.545 88.255 133.715 88.425 ;
        RECT 133.545 87.895 133.715 88.065 ;
        RECT 133.545 87.535 133.715 87.705 ;
        RECT 133.545 87.175 133.715 87.345 ;
        RECT 133.545 86.815 133.715 86.985 ;
        RECT 138.125 92.935 138.295 93.105 ;
        RECT 138.125 92.575 138.295 92.745 ;
        RECT 138.125 92.215 138.295 92.385 ;
        RECT 138.125 91.855 138.295 92.025 ;
        RECT 138.125 91.495 138.295 91.665 ;
        RECT 138.125 91.135 138.295 91.305 ;
        RECT 138.125 90.775 138.295 90.945 ;
        RECT 138.125 90.415 138.295 90.585 ;
        RECT 138.125 90.055 138.295 90.225 ;
        RECT 138.125 89.695 138.295 89.865 ;
        RECT 138.125 89.335 138.295 89.505 ;
        RECT 138.125 88.975 138.295 89.145 ;
        RECT 138.125 88.615 138.295 88.785 ;
        RECT 138.125 88.255 138.295 88.425 ;
        RECT 138.125 87.895 138.295 88.065 ;
        RECT 138.125 87.535 138.295 87.705 ;
        RECT 138.125 87.175 138.295 87.345 ;
        RECT 138.125 86.815 138.295 86.985 ;
        RECT 142.705 92.935 142.875 93.105 ;
        RECT 142.705 92.575 142.875 92.745 ;
        RECT 142.705 92.215 142.875 92.385 ;
        RECT 142.705 91.855 142.875 92.025 ;
        RECT 142.705 91.495 142.875 91.665 ;
        RECT 142.705 91.135 142.875 91.305 ;
        RECT 142.705 90.775 142.875 90.945 ;
        RECT 142.705 90.415 142.875 90.585 ;
        RECT 142.705 90.055 142.875 90.225 ;
        RECT 142.705 89.695 142.875 89.865 ;
        RECT 142.705 89.335 142.875 89.505 ;
        RECT 142.705 88.975 142.875 89.145 ;
        RECT 142.705 88.615 142.875 88.785 ;
        RECT 142.705 88.255 142.875 88.425 ;
        RECT 142.705 87.895 142.875 88.065 ;
        RECT 142.705 87.535 142.875 87.705 ;
        RECT 142.705 87.175 142.875 87.345 ;
        RECT 142.705 86.815 142.875 86.985 ;
        RECT 147.285 92.935 147.455 93.105 ;
        RECT 147.285 92.575 147.455 92.745 ;
        RECT 147.285 92.215 147.455 92.385 ;
        RECT 147.285 91.855 147.455 92.025 ;
        RECT 147.285 91.495 147.455 91.665 ;
        RECT 147.285 91.135 147.455 91.305 ;
        RECT 147.285 90.775 147.455 90.945 ;
        RECT 147.285 90.415 147.455 90.585 ;
        RECT 147.285 90.055 147.455 90.225 ;
        RECT 147.285 89.695 147.455 89.865 ;
        RECT 147.285 89.335 147.455 89.505 ;
        RECT 147.285 88.975 147.455 89.145 ;
        RECT 147.285 88.615 147.455 88.785 ;
        RECT 147.285 88.255 147.455 88.425 ;
        RECT 147.285 87.895 147.455 88.065 ;
        RECT 147.285 87.535 147.455 87.705 ;
        RECT 147.285 87.175 147.455 87.345 ;
        RECT 147.285 86.815 147.455 86.985 ;
        RECT 151.865 92.935 152.035 93.105 ;
        RECT 151.865 92.575 152.035 92.745 ;
        RECT 151.865 92.215 152.035 92.385 ;
        RECT 151.865 91.855 152.035 92.025 ;
        RECT 151.865 91.495 152.035 91.665 ;
        RECT 151.865 91.135 152.035 91.305 ;
        RECT 151.865 90.775 152.035 90.945 ;
        RECT 151.865 90.415 152.035 90.585 ;
        RECT 151.865 90.055 152.035 90.225 ;
        RECT 151.865 89.695 152.035 89.865 ;
        RECT 151.865 89.335 152.035 89.505 ;
        RECT 151.865 88.975 152.035 89.145 ;
        RECT 151.865 88.615 152.035 88.785 ;
        RECT 151.865 88.255 152.035 88.425 ;
        RECT 151.865 87.895 152.035 88.065 ;
        RECT 151.865 87.535 152.035 87.705 ;
        RECT 151.865 87.175 152.035 87.345 ;
        RECT 151.865 86.815 152.035 86.985 ;
        RECT 156.445 92.935 156.615 93.105 ;
        RECT 156.445 92.575 156.615 92.745 ;
        RECT 156.445 92.215 156.615 92.385 ;
        RECT 156.445 91.855 156.615 92.025 ;
        RECT 156.445 91.495 156.615 91.665 ;
        RECT 156.445 91.135 156.615 91.305 ;
        RECT 156.445 90.775 156.615 90.945 ;
        RECT 156.445 90.415 156.615 90.585 ;
        RECT 156.445 90.055 156.615 90.225 ;
        RECT 156.445 89.695 156.615 89.865 ;
        RECT 156.445 89.335 156.615 89.505 ;
        RECT 156.445 88.975 156.615 89.145 ;
        RECT 156.445 88.615 156.615 88.785 ;
        RECT 156.445 88.255 156.615 88.425 ;
        RECT 156.445 87.895 156.615 88.065 ;
        RECT 156.445 87.535 156.615 87.705 ;
        RECT 156.445 87.175 156.615 87.345 ;
        RECT 156.445 86.815 156.615 86.985 ;
        RECT 161.025 92.935 161.195 93.105 ;
        RECT 161.025 92.575 161.195 92.745 ;
        RECT 161.025 92.215 161.195 92.385 ;
        RECT 161.025 91.855 161.195 92.025 ;
        RECT 161.025 91.495 161.195 91.665 ;
        RECT 161.025 91.135 161.195 91.305 ;
        RECT 161.025 90.775 161.195 90.945 ;
        RECT 161.025 90.415 161.195 90.585 ;
        RECT 161.025 90.055 161.195 90.225 ;
        RECT 161.025 89.695 161.195 89.865 ;
        RECT 161.025 89.335 161.195 89.505 ;
        RECT 161.025 88.975 161.195 89.145 ;
        RECT 161.025 88.615 161.195 88.785 ;
        RECT 161.025 88.255 161.195 88.425 ;
        RECT 161.025 87.895 161.195 88.065 ;
        RECT 161.025 87.535 161.195 87.705 ;
        RECT 161.025 87.175 161.195 87.345 ;
        RECT 161.025 86.815 161.195 86.985 ;
        RECT 165.605 92.935 165.775 93.105 ;
        RECT 165.605 92.575 165.775 92.745 ;
        RECT 165.605 92.215 165.775 92.385 ;
        RECT 165.605 91.855 165.775 92.025 ;
        RECT 165.605 91.495 165.775 91.665 ;
        RECT 165.605 91.135 165.775 91.305 ;
        RECT 165.605 90.775 165.775 90.945 ;
        RECT 165.605 90.415 165.775 90.585 ;
        RECT 165.605 90.055 165.775 90.225 ;
        RECT 165.605 89.695 165.775 89.865 ;
        RECT 165.605 89.335 165.775 89.505 ;
        RECT 165.605 88.975 165.775 89.145 ;
        RECT 165.605 88.615 165.775 88.785 ;
        RECT 165.605 88.255 165.775 88.425 ;
        RECT 165.605 87.895 165.775 88.065 ;
        RECT 165.605 87.535 165.775 87.705 ;
        RECT 165.605 87.175 165.775 87.345 ;
        RECT 165.605 86.815 165.775 86.985 ;
        RECT 170.185 92.935 170.355 93.105 ;
        RECT 170.185 92.575 170.355 92.745 ;
        RECT 170.185 92.215 170.355 92.385 ;
        RECT 170.185 91.855 170.355 92.025 ;
        RECT 170.185 91.495 170.355 91.665 ;
        RECT 170.185 91.135 170.355 91.305 ;
        RECT 170.185 90.775 170.355 90.945 ;
        RECT 170.185 90.415 170.355 90.585 ;
        RECT 170.185 90.055 170.355 90.225 ;
        RECT 170.185 89.695 170.355 89.865 ;
        RECT 170.185 89.335 170.355 89.505 ;
        RECT 170.185 88.975 170.355 89.145 ;
        RECT 170.185 88.615 170.355 88.785 ;
        RECT 170.185 88.255 170.355 88.425 ;
        RECT 170.185 87.895 170.355 88.065 ;
        RECT 170.185 87.535 170.355 87.705 ;
        RECT 170.185 87.175 170.355 87.345 ;
        RECT 170.185 86.815 170.355 86.985 ;
        RECT 174.765 92.935 174.935 93.105 ;
        RECT 174.765 92.575 174.935 92.745 ;
        RECT 174.765 92.215 174.935 92.385 ;
        RECT 174.765 91.855 174.935 92.025 ;
        RECT 174.765 91.495 174.935 91.665 ;
        RECT 174.765 91.135 174.935 91.305 ;
        RECT 174.765 90.775 174.935 90.945 ;
        RECT 174.765 90.415 174.935 90.585 ;
        RECT 174.765 90.055 174.935 90.225 ;
        RECT 174.765 89.695 174.935 89.865 ;
        RECT 174.765 89.335 174.935 89.505 ;
        RECT 174.765 88.975 174.935 89.145 ;
        RECT 174.765 88.615 174.935 88.785 ;
        RECT 174.765 88.255 174.935 88.425 ;
        RECT 174.765 87.895 174.935 88.065 ;
        RECT 174.765 87.535 174.935 87.705 ;
        RECT 174.765 87.175 174.935 87.345 ;
        RECT 174.765 86.815 174.935 86.985 ;
        RECT 179.345 92.935 179.515 93.105 ;
        RECT 179.345 92.575 179.515 92.745 ;
        RECT 179.345 92.215 179.515 92.385 ;
        RECT 179.345 91.855 179.515 92.025 ;
        RECT 179.345 91.495 179.515 91.665 ;
        RECT 179.345 91.135 179.515 91.305 ;
        RECT 179.345 90.775 179.515 90.945 ;
        RECT 179.345 90.415 179.515 90.585 ;
        RECT 179.345 90.055 179.515 90.225 ;
        RECT 179.345 89.695 179.515 89.865 ;
        RECT 179.345 89.335 179.515 89.505 ;
        RECT 179.345 88.975 179.515 89.145 ;
        RECT 179.345 88.615 179.515 88.785 ;
        RECT 179.345 88.255 179.515 88.425 ;
        RECT 179.345 87.895 179.515 88.065 ;
        RECT 179.345 87.535 179.515 87.705 ;
        RECT 179.345 87.175 179.515 87.345 ;
        RECT 179.345 86.815 179.515 86.985 ;
        RECT 183.925 92.935 184.095 93.105 ;
        RECT 183.925 92.575 184.095 92.745 ;
        RECT 183.925 92.215 184.095 92.385 ;
        RECT 183.925 91.855 184.095 92.025 ;
        RECT 183.925 91.495 184.095 91.665 ;
        RECT 183.925 91.135 184.095 91.305 ;
        RECT 183.925 90.775 184.095 90.945 ;
        RECT 183.925 90.415 184.095 90.585 ;
        RECT 183.925 90.055 184.095 90.225 ;
        RECT 183.925 89.695 184.095 89.865 ;
        RECT 183.925 89.335 184.095 89.505 ;
        RECT 183.925 88.975 184.095 89.145 ;
        RECT 183.925 88.615 184.095 88.785 ;
        RECT 183.925 88.255 184.095 88.425 ;
        RECT 183.925 87.895 184.095 88.065 ;
        RECT 183.925 87.535 184.095 87.705 ;
        RECT 183.925 87.175 184.095 87.345 ;
        RECT 183.925 86.815 184.095 86.985 ;
        RECT 188.505 92.935 188.675 93.105 ;
        RECT 188.505 92.575 188.675 92.745 ;
        RECT 188.505 92.215 188.675 92.385 ;
        RECT 188.505 91.855 188.675 92.025 ;
        RECT 188.505 91.495 188.675 91.665 ;
        RECT 188.505 91.135 188.675 91.305 ;
        RECT 188.505 90.775 188.675 90.945 ;
        RECT 188.505 90.415 188.675 90.585 ;
        RECT 188.505 90.055 188.675 90.225 ;
        RECT 188.505 89.695 188.675 89.865 ;
        RECT 188.505 89.335 188.675 89.505 ;
        RECT 188.505 88.975 188.675 89.145 ;
        RECT 188.505 88.615 188.675 88.785 ;
        RECT 188.505 88.255 188.675 88.425 ;
        RECT 188.505 87.895 188.675 88.065 ;
        RECT 188.505 87.535 188.675 87.705 ;
        RECT 188.505 87.175 188.675 87.345 ;
        RECT 188.505 86.815 188.675 86.985 ;
        RECT 193.085 92.935 193.255 93.105 ;
        RECT 193.085 92.575 193.255 92.745 ;
        RECT 193.085 92.215 193.255 92.385 ;
        RECT 193.085 91.855 193.255 92.025 ;
        RECT 193.085 91.495 193.255 91.665 ;
        RECT 193.085 91.135 193.255 91.305 ;
        RECT 193.085 90.775 193.255 90.945 ;
        RECT 193.085 90.415 193.255 90.585 ;
        RECT 193.085 90.055 193.255 90.225 ;
        RECT 193.085 89.695 193.255 89.865 ;
        RECT 193.085 89.335 193.255 89.505 ;
        RECT 193.085 88.975 193.255 89.145 ;
        RECT 193.085 88.615 193.255 88.785 ;
        RECT 193.085 88.255 193.255 88.425 ;
        RECT 193.085 87.895 193.255 88.065 ;
        RECT 193.085 87.535 193.255 87.705 ;
        RECT 193.085 87.175 193.255 87.345 ;
        RECT 193.085 86.815 193.255 86.985 ;
        RECT 197.665 92.935 197.835 93.105 ;
        RECT 197.665 92.575 197.835 92.745 ;
        RECT 197.665 92.215 197.835 92.385 ;
        RECT 197.665 91.855 197.835 92.025 ;
        RECT 197.665 91.495 197.835 91.665 ;
        RECT 197.665 91.135 197.835 91.305 ;
        RECT 197.665 90.775 197.835 90.945 ;
        RECT 197.665 90.415 197.835 90.585 ;
        RECT 197.665 90.055 197.835 90.225 ;
        RECT 197.665 89.695 197.835 89.865 ;
        RECT 197.665 89.335 197.835 89.505 ;
        RECT 197.665 88.975 197.835 89.145 ;
        RECT 197.665 88.615 197.835 88.785 ;
        RECT 197.665 88.255 197.835 88.425 ;
        RECT 197.665 87.895 197.835 88.065 ;
        RECT 197.665 87.535 197.835 87.705 ;
        RECT 197.665 87.175 197.835 87.345 ;
        RECT 197.665 86.815 197.835 86.985 ;
        RECT 202.245 92.935 202.415 93.105 ;
        RECT 202.245 92.575 202.415 92.745 ;
        RECT 202.245 92.215 202.415 92.385 ;
        RECT 202.245 91.855 202.415 92.025 ;
        RECT 202.245 91.495 202.415 91.665 ;
        RECT 202.245 91.135 202.415 91.305 ;
        RECT 202.245 90.775 202.415 90.945 ;
        RECT 202.245 90.415 202.415 90.585 ;
        RECT 202.245 90.055 202.415 90.225 ;
        RECT 202.245 89.695 202.415 89.865 ;
        RECT 202.245 89.335 202.415 89.505 ;
        RECT 202.245 88.975 202.415 89.145 ;
        RECT 202.245 88.615 202.415 88.785 ;
        RECT 202.245 88.255 202.415 88.425 ;
        RECT 202.245 87.895 202.415 88.065 ;
        RECT 202.245 87.535 202.415 87.705 ;
        RECT 202.245 87.175 202.415 87.345 ;
        RECT 202.245 86.815 202.415 86.985 ;
        RECT 206.825 92.935 206.995 93.105 ;
        RECT 206.825 92.575 206.995 92.745 ;
        RECT 206.825 92.215 206.995 92.385 ;
        RECT 206.825 91.855 206.995 92.025 ;
        RECT 206.825 91.495 206.995 91.665 ;
        RECT 206.825 91.135 206.995 91.305 ;
        RECT 206.825 90.775 206.995 90.945 ;
        RECT 206.825 90.415 206.995 90.585 ;
        RECT 206.825 90.055 206.995 90.225 ;
        RECT 206.825 89.695 206.995 89.865 ;
        RECT 206.825 89.335 206.995 89.505 ;
        RECT 206.825 88.975 206.995 89.145 ;
        RECT 206.825 88.615 206.995 88.785 ;
        RECT 206.825 88.255 206.995 88.425 ;
        RECT 206.825 87.895 206.995 88.065 ;
        RECT 206.825 87.535 206.995 87.705 ;
        RECT 206.825 87.175 206.995 87.345 ;
        RECT 206.825 86.815 206.995 86.985 ;
        RECT 211.405 92.935 211.575 93.105 ;
        RECT 211.405 92.575 211.575 92.745 ;
        RECT 211.405 92.215 211.575 92.385 ;
        RECT 211.405 91.855 211.575 92.025 ;
        RECT 211.405 91.495 211.575 91.665 ;
        RECT 211.405 91.135 211.575 91.305 ;
        RECT 211.405 90.775 211.575 90.945 ;
        RECT 211.405 90.415 211.575 90.585 ;
        RECT 211.405 90.055 211.575 90.225 ;
        RECT 211.405 89.695 211.575 89.865 ;
        RECT 211.405 89.335 211.575 89.505 ;
        RECT 211.405 88.975 211.575 89.145 ;
        RECT 211.405 88.615 211.575 88.785 ;
        RECT 211.405 88.255 211.575 88.425 ;
        RECT 211.405 87.895 211.575 88.065 ;
        RECT 211.405 87.535 211.575 87.705 ;
        RECT 211.405 87.175 211.575 87.345 ;
        RECT 211.405 86.815 211.575 86.985 ;
        RECT 215.985 92.935 216.155 93.105 ;
        RECT 215.985 92.575 216.155 92.745 ;
        RECT 215.985 92.215 216.155 92.385 ;
        RECT 215.985 91.855 216.155 92.025 ;
        RECT 215.985 91.495 216.155 91.665 ;
        RECT 215.985 91.135 216.155 91.305 ;
        RECT 215.985 90.775 216.155 90.945 ;
        RECT 215.985 90.415 216.155 90.585 ;
        RECT 215.985 90.055 216.155 90.225 ;
        RECT 215.985 89.695 216.155 89.865 ;
        RECT 215.985 89.335 216.155 89.505 ;
        RECT 215.985 88.975 216.155 89.145 ;
        RECT 215.985 88.615 216.155 88.785 ;
        RECT 215.985 88.255 216.155 88.425 ;
        RECT 215.985 87.895 216.155 88.065 ;
        RECT 215.985 87.535 216.155 87.705 ;
        RECT 215.985 87.175 216.155 87.345 ;
        RECT 215.985 86.815 216.155 86.985 ;
        RECT 220.565 92.935 220.735 93.105 ;
        RECT 220.565 92.575 220.735 92.745 ;
        RECT 220.565 92.215 220.735 92.385 ;
        RECT 220.565 91.855 220.735 92.025 ;
        RECT 220.565 91.495 220.735 91.665 ;
        RECT 220.565 91.135 220.735 91.305 ;
        RECT 220.565 90.775 220.735 90.945 ;
        RECT 220.565 90.415 220.735 90.585 ;
        RECT 220.565 90.055 220.735 90.225 ;
        RECT 220.565 89.695 220.735 89.865 ;
        RECT 220.565 89.335 220.735 89.505 ;
        RECT 220.565 88.975 220.735 89.145 ;
        RECT 220.565 88.615 220.735 88.785 ;
        RECT 220.565 88.255 220.735 88.425 ;
        RECT 220.565 87.895 220.735 88.065 ;
        RECT 220.565 87.535 220.735 87.705 ;
        RECT 220.565 87.175 220.735 87.345 ;
        RECT 220.565 86.815 220.735 86.985 ;
        RECT 225.145 92.935 225.315 93.105 ;
        RECT 225.145 92.575 225.315 92.745 ;
        RECT 225.145 92.215 225.315 92.385 ;
        RECT 225.145 91.855 225.315 92.025 ;
        RECT 225.145 91.495 225.315 91.665 ;
        RECT 225.145 91.135 225.315 91.305 ;
        RECT 225.145 90.775 225.315 90.945 ;
        RECT 225.145 90.415 225.315 90.585 ;
        RECT 225.145 90.055 225.315 90.225 ;
        RECT 225.145 89.695 225.315 89.865 ;
        RECT 225.145 89.335 225.315 89.505 ;
        RECT 225.145 88.975 225.315 89.145 ;
        RECT 225.145 88.615 225.315 88.785 ;
        RECT 225.145 88.255 225.315 88.425 ;
        RECT 225.145 87.895 225.315 88.065 ;
        RECT 225.145 87.535 225.315 87.705 ;
        RECT 225.145 87.175 225.315 87.345 ;
        RECT 225.145 86.815 225.315 86.985 ;
        RECT 229.725 92.935 229.895 93.105 ;
        RECT 229.725 92.575 229.895 92.745 ;
        RECT 229.725 92.215 229.895 92.385 ;
        RECT 229.725 91.855 229.895 92.025 ;
        RECT 229.725 91.495 229.895 91.665 ;
        RECT 229.725 91.135 229.895 91.305 ;
        RECT 229.725 90.775 229.895 90.945 ;
        RECT 229.725 90.415 229.895 90.585 ;
        RECT 229.725 90.055 229.895 90.225 ;
        RECT 229.725 89.695 229.895 89.865 ;
        RECT 229.725 89.335 229.895 89.505 ;
        RECT 229.725 88.975 229.895 89.145 ;
        RECT 229.725 88.615 229.895 88.785 ;
        RECT 229.725 88.255 229.895 88.425 ;
        RECT 229.725 87.895 229.895 88.065 ;
        RECT 229.725 87.535 229.895 87.705 ;
        RECT 229.725 87.175 229.895 87.345 ;
        RECT 229.725 86.815 229.895 86.985 ;
        RECT 234.305 92.935 234.475 93.105 ;
        RECT 234.305 92.575 234.475 92.745 ;
        RECT 234.305 92.215 234.475 92.385 ;
        RECT 234.305 91.855 234.475 92.025 ;
        RECT 234.305 91.495 234.475 91.665 ;
        RECT 234.305 91.135 234.475 91.305 ;
        RECT 234.305 90.775 234.475 90.945 ;
        RECT 234.305 90.415 234.475 90.585 ;
        RECT 234.305 90.055 234.475 90.225 ;
        RECT 234.305 89.695 234.475 89.865 ;
        RECT 234.305 89.335 234.475 89.505 ;
        RECT 234.305 88.975 234.475 89.145 ;
        RECT 234.305 88.615 234.475 88.785 ;
        RECT 234.305 88.255 234.475 88.425 ;
        RECT 234.305 87.895 234.475 88.065 ;
        RECT 234.305 87.535 234.475 87.705 ;
        RECT 234.305 87.175 234.475 87.345 ;
        RECT 234.305 86.815 234.475 86.985 ;
        RECT 238.885 92.935 239.055 93.105 ;
        RECT 238.885 92.575 239.055 92.745 ;
        RECT 238.885 92.215 239.055 92.385 ;
        RECT 238.885 91.855 239.055 92.025 ;
        RECT 238.885 91.495 239.055 91.665 ;
        RECT 238.885 91.135 239.055 91.305 ;
        RECT 238.885 90.775 239.055 90.945 ;
        RECT 238.885 90.415 239.055 90.585 ;
        RECT 238.885 90.055 239.055 90.225 ;
        RECT 238.885 89.695 239.055 89.865 ;
        RECT 238.885 89.335 239.055 89.505 ;
        RECT 238.885 88.975 239.055 89.145 ;
        RECT 238.885 88.615 239.055 88.785 ;
        RECT 238.885 88.255 239.055 88.425 ;
        RECT 238.885 87.895 239.055 88.065 ;
        RECT 238.885 87.535 239.055 87.705 ;
        RECT 238.885 87.175 239.055 87.345 ;
        RECT 238.885 86.815 239.055 86.985 ;
        RECT 243.465 92.935 243.635 93.105 ;
        RECT 243.465 92.575 243.635 92.745 ;
        RECT 243.465 92.215 243.635 92.385 ;
        RECT 243.465 91.855 243.635 92.025 ;
        RECT 243.465 91.495 243.635 91.665 ;
        RECT 243.465 91.135 243.635 91.305 ;
        RECT 243.465 90.775 243.635 90.945 ;
        RECT 243.465 90.415 243.635 90.585 ;
        RECT 243.465 90.055 243.635 90.225 ;
        RECT 243.465 89.695 243.635 89.865 ;
        RECT 243.465 89.335 243.635 89.505 ;
        RECT 243.465 88.975 243.635 89.145 ;
        RECT 243.465 88.615 243.635 88.785 ;
        RECT 243.465 88.255 243.635 88.425 ;
        RECT 243.465 87.895 243.635 88.065 ;
        RECT 243.465 87.535 243.635 87.705 ;
        RECT 243.465 87.175 243.635 87.345 ;
        RECT 243.465 86.815 243.635 86.985 ;
        RECT 248.045 92.935 248.215 93.105 ;
        RECT 248.045 92.575 248.215 92.745 ;
        RECT 248.045 92.215 248.215 92.385 ;
        RECT 248.045 91.855 248.215 92.025 ;
        RECT 248.045 91.495 248.215 91.665 ;
        RECT 248.045 91.135 248.215 91.305 ;
        RECT 248.045 90.775 248.215 90.945 ;
        RECT 248.045 90.415 248.215 90.585 ;
        RECT 248.045 90.055 248.215 90.225 ;
        RECT 248.045 89.695 248.215 89.865 ;
        RECT 248.045 89.335 248.215 89.505 ;
        RECT 248.045 88.975 248.215 89.145 ;
        RECT 248.045 88.615 248.215 88.785 ;
        RECT 248.045 88.255 248.215 88.425 ;
        RECT 248.045 87.895 248.215 88.065 ;
        RECT 248.045 87.535 248.215 87.705 ;
        RECT 248.045 87.175 248.215 87.345 ;
        RECT 248.045 86.815 248.215 86.985 ;
        RECT 252.625 92.935 252.795 93.105 ;
        RECT 252.625 92.575 252.795 92.745 ;
        RECT 252.625 92.215 252.795 92.385 ;
        RECT 252.625 91.855 252.795 92.025 ;
        RECT 252.625 91.495 252.795 91.665 ;
        RECT 252.625 91.135 252.795 91.305 ;
        RECT 252.625 90.775 252.795 90.945 ;
        RECT 252.625 90.415 252.795 90.585 ;
        RECT 252.625 90.055 252.795 90.225 ;
        RECT 252.625 89.695 252.795 89.865 ;
        RECT 252.625 89.335 252.795 89.505 ;
        RECT 252.625 88.975 252.795 89.145 ;
        RECT 252.625 88.615 252.795 88.785 ;
        RECT 252.625 88.255 252.795 88.425 ;
        RECT 252.625 87.895 252.795 88.065 ;
        RECT 252.625 87.535 252.795 87.705 ;
        RECT 252.625 87.175 252.795 87.345 ;
        RECT 252.625 86.815 252.795 86.985 ;
        RECT 257.205 92.935 257.375 93.105 ;
        RECT 257.205 92.575 257.375 92.745 ;
        RECT 257.205 92.215 257.375 92.385 ;
        RECT 257.205 91.855 257.375 92.025 ;
        RECT 257.205 91.495 257.375 91.665 ;
        RECT 257.205 91.135 257.375 91.305 ;
        RECT 257.205 90.775 257.375 90.945 ;
        RECT 257.205 90.415 257.375 90.585 ;
        RECT 257.205 90.055 257.375 90.225 ;
        RECT 257.205 89.695 257.375 89.865 ;
        RECT 257.205 89.335 257.375 89.505 ;
        RECT 257.205 88.975 257.375 89.145 ;
        RECT 257.205 88.615 257.375 88.785 ;
        RECT 257.205 88.255 257.375 88.425 ;
        RECT 257.205 87.895 257.375 88.065 ;
        RECT 257.205 87.535 257.375 87.705 ;
        RECT 257.205 87.175 257.375 87.345 ;
        RECT 257.205 86.815 257.375 86.985 ;
        RECT 261.785 92.935 261.955 93.105 ;
        RECT 261.785 92.575 261.955 92.745 ;
        RECT 261.785 92.215 261.955 92.385 ;
        RECT 261.785 91.855 261.955 92.025 ;
        RECT 261.785 91.495 261.955 91.665 ;
        RECT 261.785 91.135 261.955 91.305 ;
        RECT 261.785 90.775 261.955 90.945 ;
        RECT 261.785 90.415 261.955 90.585 ;
        RECT 261.785 90.055 261.955 90.225 ;
        RECT 261.785 89.695 261.955 89.865 ;
        RECT 261.785 89.335 261.955 89.505 ;
        RECT 261.785 88.975 261.955 89.145 ;
        RECT 261.785 88.615 261.955 88.785 ;
        RECT 261.785 88.255 261.955 88.425 ;
        RECT 261.785 87.895 261.955 88.065 ;
        RECT 261.785 87.535 261.955 87.705 ;
        RECT 261.785 87.175 261.955 87.345 ;
        RECT 261.785 86.815 261.955 86.985 ;
        RECT 171.725 86.105 171.895 86.275 ;
        RECT 218.915 52.815 220.885 55.505 ;
      LAYER met1 ;
        RECT 124.355 86.735 124.585 93.185 ;
        RECT 128.935 86.735 129.165 93.185 ;
        RECT 133.515 86.735 133.745 93.185 ;
        RECT 138.095 86.735 138.325 93.185 ;
        RECT 142.675 86.735 142.905 93.185 ;
        RECT 147.255 86.735 147.485 93.185 ;
        RECT 151.835 86.735 152.065 93.185 ;
        RECT 156.415 86.735 156.645 93.185 ;
        RECT 160.995 86.735 161.225 93.185 ;
        RECT 165.575 86.735 165.805 93.185 ;
        RECT 170.155 86.735 170.385 93.185 ;
        RECT 174.735 86.735 174.965 93.185 ;
        RECT 179.315 86.735 179.545 93.185 ;
        RECT 183.895 86.735 184.125 93.185 ;
        RECT 188.475 86.735 188.705 93.185 ;
        RECT 193.055 86.735 193.285 93.185 ;
        RECT 197.635 86.735 197.865 93.185 ;
        RECT 202.215 86.735 202.445 93.185 ;
        RECT 206.795 86.735 207.025 93.185 ;
        RECT 211.375 86.735 211.605 93.185 ;
        RECT 215.955 86.735 216.185 93.185 ;
        RECT 219.950 86.940 220.270 87.000 ;
        RECT 220.535 86.940 220.765 93.185 ;
        RECT 219.950 86.800 220.765 86.940 ;
        RECT 219.950 86.740 220.270 86.800 ;
        RECT 220.535 86.735 220.765 86.800 ;
        RECT 225.115 86.735 225.345 93.185 ;
        RECT 229.695 86.735 229.925 93.185 ;
        RECT 234.275 86.735 234.505 93.185 ;
        RECT 238.855 86.735 239.085 93.185 ;
        RECT 243.435 86.735 243.665 93.185 ;
        RECT 248.015 86.735 248.245 93.185 ;
        RECT 252.595 86.735 252.825 93.185 ;
        RECT 257.175 86.735 257.405 93.185 ;
        RECT 261.755 86.735 261.985 93.185 ;
        RECT 171.650 86.260 171.970 86.320 ;
        RECT 171.375 86.120 171.970 86.260 ;
        RECT 171.650 86.060 171.970 86.120 ;
        RECT 218.875 52.755 220.925 55.565 ;
      LAYER via ;
        RECT 219.980 86.740 220.240 87.000 ;
        RECT 171.680 86.060 171.940 86.320 ;
        RECT 219.980 55.120 220.240 55.380 ;
      LAYER met2 ;
        RECT 219.980 86.710 220.240 87.030 ;
        RECT 171.680 86.030 171.940 86.350 ;
        RECT 171.740 0.000 171.880 86.030 ;
        RECT 220.040 55.410 220.180 86.710 ;
        RECT 219.980 55.090 220.240 55.410 ;
    END
  END vbg
  PIN VSS
    ANTENNAGATEAREA 1069.156006 ;
    ANTENNADIFFAREA 893.893555 ;
    PORT
      LAYER pwell ;
        RECT 108.590 239.180 111.930 240.340 ;
        RECT 119.160 235.630 119.620 236.490 ;
        RECT 214.800 223.845 261.700 224.610 ;
        RECT 214.800 218.675 215.565 223.845 ;
        RECT 220.735 218.675 222.265 223.845 ;
        RECT 227.435 218.675 228.965 223.845 ;
        RECT 234.135 218.675 235.665 223.845 ;
        RECT 240.835 218.675 242.365 223.845 ;
        RECT 247.535 218.675 249.065 223.845 ;
        RECT 254.235 218.675 255.765 223.845 ;
        RECT 260.935 218.675 261.700 223.845 ;
        RECT 214.800 217.910 261.700 218.675 ;
        RECT 70.160 216.830 70.620 217.690 ;
        RECT 208.920 205.045 262.520 205.810 ;
        RECT 208.920 199.875 209.685 205.045 ;
        RECT 214.855 199.875 216.385 205.045 ;
        RECT 221.555 199.875 223.085 205.045 ;
        RECT 228.255 199.875 229.785 205.045 ;
        RECT 234.955 199.875 236.485 205.045 ;
        RECT 241.655 199.875 243.185 205.045 ;
        RECT 248.355 199.875 249.885 205.045 ;
        RECT 255.055 199.875 256.585 205.045 ;
        RECT 261.755 199.875 262.520 205.045 ;
        RECT 208.920 199.110 262.520 199.875 ;
        RECT 185.950 198.030 186.410 198.890 ;
        RECT 191.250 198.030 192.110 198.540 ;
        RECT 197.750 198.030 198.610 198.540 ;
        RECT 59.960 186.245 66.660 187.010 ;
        RECT 59.960 181.075 60.725 186.245 ;
        RECT 65.895 181.075 66.660 186.245 ;
        RECT 208.920 186.245 262.520 187.010 ;
        RECT 72.820 182.780 76.160 183.940 ;
        RECT 86.540 182.780 89.880 183.940 ;
        RECT 101.700 182.780 105.040 183.940 ;
        RECT 116.920 182.780 120.260 183.940 ;
        RECT 59.960 180.310 66.660 181.075 ;
        RECT 208.920 181.075 209.685 186.245 ;
        RECT 214.855 181.075 216.385 186.245 ;
        RECT 221.555 181.075 223.085 186.245 ;
        RECT 228.255 181.075 229.785 186.245 ;
        RECT 234.955 181.075 236.485 186.245 ;
        RECT 241.655 181.075 243.185 186.245 ;
        RECT 248.355 181.075 249.885 186.245 ;
        RECT 255.055 181.075 256.585 186.245 ;
        RECT 261.755 181.075 262.520 186.245 ;
        RECT 208.920 180.310 262.520 181.075 ;
        RECT 126.660 179.230 127.120 180.090 ;
        RECT 131.960 179.230 132.820 179.740 ;
        RECT 138.460 179.230 139.320 179.740 ;
        RECT 208.920 167.445 262.520 168.210 ;
        RECT 100.750 163.980 104.090 165.140 ;
        RECT 115.910 163.980 119.250 165.140 ;
        RECT 208.920 162.275 209.685 167.445 ;
        RECT 214.855 162.275 216.385 167.445 ;
        RECT 221.555 162.275 223.085 167.445 ;
        RECT 228.255 162.275 229.785 167.445 ;
        RECT 234.955 162.275 236.485 167.445 ;
        RECT 241.655 162.275 243.185 167.445 ;
        RECT 248.355 162.275 249.885 167.445 ;
        RECT 255.055 162.275 256.585 167.445 ;
        RECT 261.755 162.275 262.520 167.445 ;
        RECT 208.920 161.510 262.520 162.275 ;
        RECT 208.920 148.645 262.520 149.410 ;
        RECT 87.030 145.180 90.370 146.340 ;
        RECT 100.750 145.180 104.090 146.340 ;
        RECT 114.470 145.180 117.810 146.340 ;
        RECT 140.440 145.180 143.780 146.340 ;
        RECT 208.920 143.475 209.685 148.645 ;
        RECT 214.855 143.475 216.385 148.645 ;
        RECT 221.555 143.475 223.085 148.645 ;
        RECT 228.255 143.475 229.785 148.645 ;
        RECT 234.955 143.475 236.485 148.645 ;
        RECT 241.655 143.475 243.185 148.645 ;
        RECT 248.355 143.475 249.885 148.645 ;
        RECT 255.055 143.475 256.585 148.645 ;
        RECT 261.755 143.475 262.520 148.645 ;
        RECT 208.920 142.710 262.520 143.475 ;
        RECT 116.430 126.380 119.770 127.540 ;
        RECT 191.400 126.380 194.740 127.540 ;
        RECT 205.120 126.380 208.460 127.540 ;
        RECT 218.840 126.380 222.180 127.540 ;
        RECT 232.560 126.380 235.900 127.540 ;
        RECT 246.280 126.380 249.620 127.540 ;
        RECT 126.660 122.830 127.120 123.690 ;
        RECT 131.960 122.830 132.820 123.340 ;
        RECT 138.460 122.830 139.320 123.340 ;
        RECT 123.780 107.580 127.120 108.740 ;
        RECT 140.440 107.580 143.780 108.740 ;
        RECT 154.160 107.580 157.500 108.740 ;
        RECT 170.330 107.580 173.670 108.740 ;
        RECT 191.400 107.580 194.740 108.740 ;
        RECT 205.120 107.580 208.460 108.740 ;
        RECT 246.280 107.580 249.620 108.740 ;
        RECT 223.740 69.980 227.080 71.140 ;
        RECT 237.460 69.980 240.800 71.140 ;
        RECT 251.180 69.980 254.520 71.140 ;
        RECT 223.250 51.180 226.590 52.340 ;
        RECT 236.970 51.180 240.310 52.340 ;
        RECT 250.690 51.180 254.030 52.340 ;
        RECT 227.170 32.380 230.510 33.540 ;
        RECT 240.890 32.380 244.230 33.540 ;
        RECT 254.610 32.380 257.950 33.540 ;
      LAYER li1 ;
        RECT 119.590 243.810 122.170 244.110 ;
        RECT 121.935 242.380 122.105 243.810 ;
        RECT 121.935 242.290 122.110 242.380 ;
        RECT 108.720 235.510 111.800 240.210 ;
        RECT 121.940 238.340 122.110 242.290 ;
        RECT 119.240 235.510 119.540 236.560 ;
        RECT 29.590 235.210 65.430 235.510 ;
        RECT 66.830 235.210 102.670 235.510 ;
        RECT 104.160 235.210 116.360 235.510 ;
        RECT 119.100 235.210 122.170 235.510 ;
        RECT 123.660 235.210 262.190 235.510 ;
        RECT 70.590 225.010 73.170 225.310 ;
        RECT 72.935 223.580 73.105 225.010 ;
        RECT 214.930 223.985 261.570 224.480 ;
        RECT 72.935 223.490 73.110 223.580 ;
        RECT 72.940 219.540 73.110 223.490 ;
        RECT 214.930 218.535 215.425 223.985 ;
        RECT 215.745 223.305 220.555 223.665 ;
        RECT 215.745 219.215 216.105 223.305 ;
        RECT 220.195 219.215 220.555 223.305 ;
        RECT 215.745 218.855 220.555 219.215 ;
        RECT 220.875 218.535 222.125 223.985 ;
        RECT 222.445 223.305 227.255 223.665 ;
        RECT 222.445 219.215 222.805 223.305 ;
        RECT 226.895 219.215 227.255 223.305 ;
        RECT 222.445 218.855 227.255 219.215 ;
        RECT 227.575 218.535 228.825 223.985 ;
        RECT 229.145 223.305 233.955 223.665 ;
        RECT 229.145 219.215 229.505 223.305 ;
        RECT 233.595 219.215 233.955 223.305 ;
        RECT 229.145 218.855 233.955 219.215 ;
        RECT 234.275 218.535 235.525 223.985 ;
        RECT 235.845 223.305 240.655 223.665 ;
        RECT 235.845 219.215 236.205 223.305 ;
        RECT 240.295 219.215 240.655 223.305 ;
        RECT 235.845 218.855 240.655 219.215 ;
        RECT 240.975 218.535 242.225 223.985 ;
        RECT 242.545 223.305 247.355 223.665 ;
        RECT 242.545 219.215 242.905 223.305 ;
        RECT 246.995 219.215 247.355 223.305 ;
        RECT 242.545 218.855 247.355 219.215 ;
        RECT 247.675 218.535 248.925 223.985 ;
        RECT 249.245 223.305 254.055 223.665 ;
        RECT 249.245 219.215 249.605 223.305 ;
        RECT 253.695 219.215 254.055 223.305 ;
        RECT 249.245 218.855 254.055 219.215 ;
        RECT 254.375 218.535 255.625 223.985 ;
        RECT 255.945 223.305 260.755 223.665 ;
        RECT 255.945 219.215 256.305 223.305 ;
        RECT 260.395 219.215 260.755 223.305 ;
        RECT 255.945 218.855 260.755 219.215 ;
        RECT 261.075 218.535 261.570 223.985 ;
        RECT 214.930 218.040 261.570 218.535 ;
        RECT 70.240 216.710 70.540 217.760 ;
        RECT 29.590 216.410 65.430 216.710 ;
        RECT 70.100 216.410 73.170 216.710 ;
        RECT 74.660 216.410 213.190 216.710 ;
        RECT 214.800 216.410 261.700 216.710 ;
        RECT 209.050 205.185 262.390 205.680 ;
        RECT 209.050 199.735 209.545 205.185 ;
        RECT 209.865 204.505 214.675 204.865 ;
        RECT 209.865 200.415 210.225 204.505 ;
        RECT 214.315 200.415 214.675 204.505 ;
        RECT 209.865 200.055 214.675 200.415 ;
        RECT 214.995 199.735 216.245 205.185 ;
        RECT 216.565 204.505 221.375 204.865 ;
        RECT 216.565 200.415 216.925 204.505 ;
        RECT 221.015 200.415 221.375 204.505 ;
        RECT 216.565 200.055 221.375 200.415 ;
        RECT 221.695 199.735 222.945 205.185 ;
        RECT 223.265 204.505 228.075 204.865 ;
        RECT 223.265 200.415 223.625 204.505 ;
        RECT 227.715 200.415 228.075 204.505 ;
        RECT 223.265 200.055 228.075 200.415 ;
        RECT 228.395 199.735 229.645 205.185 ;
        RECT 229.965 204.505 234.775 204.865 ;
        RECT 229.965 200.415 230.325 204.505 ;
        RECT 234.415 200.415 234.775 204.505 ;
        RECT 229.965 200.055 234.775 200.415 ;
        RECT 235.095 199.735 236.345 205.185 ;
        RECT 236.665 204.505 241.475 204.865 ;
        RECT 236.665 200.415 237.025 204.505 ;
        RECT 241.115 200.415 241.475 204.505 ;
        RECT 236.665 200.055 241.475 200.415 ;
        RECT 241.795 199.735 243.045 205.185 ;
        RECT 243.365 204.505 248.175 204.865 ;
        RECT 243.365 200.415 243.725 204.505 ;
        RECT 247.815 200.415 248.175 204.505 ;
        RECT 243.365 200.055 248.175 200.415 ;
        RECT 248.495 199.735 249.745 205.185 ;
        RECT 250.065 204.505 254.875 204.865 ;
        RECT 250.065 200.415 250.425 204.505 ;
        RECT 254.515 200.415 254.875 204.505 ;
        RECT 250.065 200.055 254.875 200.415 ;
        RECT 255.195 199.735 256.445 205.185 ;
        RECT 256.765 204.505 261.575 204.865 ;
        RECT 256.765 200.415 257.125 204.505 ;
        RECT 261.215 200.415 261.575 204.505 ;
        RECT 256.765 200.055 261.575 200.415 ;
        RECT 261.895 199.735 262.390 205.185 ;
        RECT 209.050 199.240 262.390 199.735 ;
        RECT 186.030 197.910 186.330 198.960 ;
        RECT 191.280 197.910 192.080 198.510 ;
        RECT 197.780 197.910 198.580 198.510 ;
        RECT 31.550 197.610 67.390 197.910 ;
        RECT 75.650 197.610 111.490 197.910 ;
        RECT 112.880 197.610 141.490 197.910 ;
        RECT 146.200 197.610 174.810 197.910 ;
        RECT 185.890 197.610 207.280 197.910 ;
        RECT 208.920 197.610 262.520 197.910 ;
        RECT 60.090 186.385 66.530 186.880 ;
        RECT 60.090 180.935 60.585 186.385 ;
        RECT 60.905 185.705 65.715 186.065 ;
        RECT 60.905 181.615 61.265 185.705 ;
        RECT 65.355 181.615 65.715 185.705 ;
        RECT 60.905 181.255 65.715 181.615 ;
        RECT 66.035 180.935 66.530 186.385 ;
        RECT 209.050 186.385 262.390 186.880 ;
        RECT 60.090 180.795 66.530 180.935 ;
        RECT 60.090 180.625 66.555 180.795 ;
        RECT 60.090 180.440 66.530 180.625 ;
        RECT 72.950 179.110 76.030 183.810 ;
        RECT 86.670 179.110 89.750 183.810 ;
        RECT 95.835 179.535 97.995 182.385 ;
        RECT 101.830 179.110 104.910 183.810 ;
        RECT 117.050 179.110 120.130 183.810 ;
        RECT 209.050 180.935 209.545 186.385 ;
        RECT 209.865 185.705 214.675 186.065 ;
        RECT 209.865 181.615 210.225 185.705 ;
        RECT 214.315 181.615 214.675 185.705 ;
        RECT 209.865 181.255 214.675 181.615 ;
        RECT 214.995 180.935 216.245 186.385 ;
        RECT 216.565 185.705 221.375 186.065 ;
        RECT 216.565 181.615 216.925 185.705 ;
        RECT 221.015 181.615 221.375 185.705 ;
        RECT 216.565 181.255 221.375 181.615 ;
        RECT 221.695 180.935 222.945 186.385 ;
        RECT 223.265 185.705 228.075 186.065 ;
        RECT 223.265 181.615 223.625 185.705 ;
        RECT 227.715 181.615 228.075 185.705 ;
        RECT 223.265 181.255 228.075 181.615 ;
        RECT 228.395 180.935 229.645 186.385 ;
        RECT 229.965 185.705 234.775 186.065 ;
        RECT 229.965 181.615 230.325 185.705 ;
        RECT 234.415 181.615 234.775 185.705 ;
        RECT 229.965 181.255 234.775 181.615 ;
        RECT 235.095 180.935 236.345 186.385 ;
        RECT 236.665 185.705 241.475 186.065 ;
        RECT 236.665 181.615 237.025 185.705 ;
        RECT 241.115 181.615 241.475 185.705 ;
        RECT 236.665 181.255 241.475 181.615 ;
        RECT 241.795 180.935 243.045 186.385 ;
        RECT 243.365 185.705 248.175 186.065 ;
        RECT 243.365 181.615 243.725 185.705 ;
        RECT 247.815 181.615 248.175 185.705 ;
        RECT 243.365 181.255 248.175 181.615 ;
        RECT 248.495 180.935 249.745 186.385 ;
        RECT 250.065 185.705 254.875 186.065 ;
        RECT 250.065 181.615 250.425 185.705 ;
        RECT 254.515 181.615 254.875 185.705 ;
        RECT 250.065 181.255 254.875 181.615 ;
        RECT 255.195 180.935 256.445 186.385 ;
        RECT 256.765 185.705 261.575 186.065 ;
        RECT 256.765 181.615 257.125 185.705 ;
        RECT 261.215 181.615 261.575 185.705 ;
        RECT 256.765 181.255 261.575 181.615 ;
        RECT 261.895 180.935 262.390 186.385 ;
        RECT 209.050 180.440 262.390 180.935 ;
        RECT 126.740 179.110 127.040 180.160 ;
        RECT 131.990 179.110 132.790 179.710 ;
        RECT 138.490 179.110 139.290 179.710 ;
        RECT 59.960 178.810 66.660 179.110 ;
        RECT 68.390 178.810 80.590 179.110 ;
        RECT 82.110 178.810 94.310 179.110 ;
        RECT 95.840 178.810 110.900 179.110 ;
        RECT 112.490 178.810 124.690 179.110 ;
        RECT 126.600 178.810 147.990 179.110 ;
        RECT 149.640 178.810 185.480 179.110 ;
        RECT 186.870 178.810 201.740 179.110 ;
        RECT 208.920 178.810 262.520 179.110 ;
        RECT 209.050 167.585 262.390 168.080 ;
        RECT 100.880 160.310 103.960 165.010 ;
        RECT 110.045 160.735 112.205 163.585 ;
        RECT 116.040 160.310 119.120 165.010 ;
        RECT 209.050 162.135 209.545 167.585 ;
        RECT 209.865 166.905 214.675 167.265 ;
        RECT 209.865 162.815 210.225 166.905 ;
        RECT 214.315 162.815 214.675 166.905 ;
        RECT 209.865 162.455 214.675 162.815 ;
        RECT 214.995 162.135 216.245 167.585 ;
        RECT 216.565 166.905 221.375 167.265 ;
        RECT 216.565 162.815 216.925 166.905 ;
        RECT 221.015 162.815 221.375 166.905 ;
        RECT 216.565 162.455 221.375 162.815 ;
        RECT 221.695 162.135 222.945 167.585 ;
        RECT 223.265 166.905 228.075 167.265 ;
        RECT 223.265 162.815 223.625 166.905 ;
        RECT 227.715 162.815 228.075 166.905 ;
        RECT 223.265 162.455 228.075 162.815 ;
        RECT 228.395 162.135 229.645 167.585 ;
        RECT 229.965 166.905 234.775 167.265 ;
        RECT 229.965 162.815 230.325 166.905 ;
        RECT 234.415 162.815 234.775 166.905 ;
        RECT 229.965 162.455 234.775 162.815 ;
        RECT 235.095 162.135 236.345 167.585 ;
        RECT 236.665 166.905 241.475 167.265 ;
        RECT 236.665 162.815 237.025 166.905 ;
        RECT 241.115 162.815 241.475 166.905 ;
        RECT 236.665 162.455 241.475 162.815 ;
        RECT 241.795 162.135 243.045 167.585 ;
        RECT 243.365 166.905 248.175 167.265 ;
        RECT 243.365 162.815 243.725 166.905 ;
        RECT 247.815 162.815 248.175 166.905 ;
        RECT 243.365 162.455 248.175 162.815 ;
        RECT 248.495 162.135 249.745 167.585 ;
        RECT 250.065 166.905 254.875 167.265 ;
        RECT 250.065 162.815 250.425 166.905 ;
        RECT 254.515 162.815 254.875 166.905 ;
        RECT 250.065 162.455 254.875 162.815 ;
        RECT 255.195 162.135 256.445 167.585 ;
        RECT 256.765 166.905 261.575 167.265 ;
        RECT 256.765 162.815 257.125 166.905 ;
        RECT 261.215 162.815 261.575 166.905 ;
        RECT 256.765 162.455 261.575 162.815 ;
        RECT 261.895 162.135 262.390 167.585 ;
        RECT 209.050 161.640 262.390 162.135 ;
        RECT 96.320 160.010 108.520 160.310 ;
        RECT 110.050 160.010 125.110 160.310 ;
        RECT 131.020 160.010 166.860 160.310 ;
        RECT 168.260 160.010 204.100 160.310 ;
        RECT 208.920 160.010 262.520 160.310 ;
        RECT 209.050 148.785 262.390 149.280 ;
        RECT 87.160 141.510 90.240 146.210 ;
        RECT 100.880 141.510 103.960 146.210 ;
        RECT 114.600 141.510 117.680 146.210 ;
        RECT 140.570 141.510 143.650 146.210 ;
        RECT 209.050 143.335 209.545 148.785 ;
        RECT 209.865 148.105 214.675 148.465 ;
        RECT 209.865 144.015 210.225 148.105 ;
        RECT 214.315 144.015 214.675 148.105 ;
        RECT 209.865 143.655 214.675 144.015 ;
        RECT 214.995 143.335 216.245 148.785 ;
        RECT 216.565 148.105 221.375 148.465 ;
        RECT 216.565 144.015 216.925 148.105 ;
        RECT 221.015 144.015 221.375 148.105 ;
        RECT 216.565 143.655 221.375 144.015 ;
        RECT 221.695 143.335 222.945 148.785 ;
        RECT 223.265 148.105 228.075 148.465 ;
        RECT 223.265 144.015 223.625 148.105 ;
        RECT 227.715 144.015 228.075 148.105 ;
        RECT 223.265 143.655 228.075 144.015 ;
        RECT 228.395 143.335 229.645 148.785 ;
        RECT 229.965 148.105 234.775 148.465 ;
        RECT 229.965 144.015 230.325 148.105 ;
        RECT 234.415 144.015 234.775 148.105 ;
        RECT 229.965 143.655 234.775 144.015 ;
        RECT 235.095 143.335 236.345 148.785 ;
        RECT 236.665 148.105 241.475 148.465 ;
        RECT 236.665 144.015 237.025 148.105 ;
        RECT 241.115 144.015 241.475 148.105 ;
        RECT 236.665 143.655 241.475 144.015 ;
        RECT 241.795 143.335 243.045 148.785 ;
        RECT 243.365 148.105 248.175 148.465 ;
        RECT 243.365 144.015 243.725 148.105 ;
        RECT 247.815 144.015 248.175 148.105 ;
        RECT 243.365 143.655 248.175 144.015 ;
        RECT 248.495 143.335 249.745 148.785 ;
        RECT 250.065 148.105 254.875 148.465 ;
        RECT 250.065 144.015 250.425 148.105 ;
        RECT 254.515 144.015 254.875 148.105 ;
        RECT 250.065 143.655 254.875 144.015 ;
        RECT 255.195 143.335 256.445 148.785 ;
        RECT 256.765 148.105 261.575 148.465 ;
        RECT 256.765 144.015 257.125 148.105 ;
        RECT 261.215 144.015 261.575 148.105 ;
        RECT 256.765 143.655 261.575 144.015 ;
        RECT 261.895 143.335 262.390 148.785 ;
        RECT 209.050 142.840 262.390 143.335 ;
        RECT 82.600 141.210 94.800 141.510 ;
        RECT 96.320 141.210 108.520 141.510 ;
        RECT 110.040 141.210 122.240 141.510 ;
        RECT 136.010 141.210 148.210 141.510 ;
        RECT 149.640 141.210 185.480 141.510 ;
        RECT 186.870 141.210 201.740 141.510 ;
        RECT 208.920 141.210 262.520 141.510 ;
        RECT 127.090 131.010 147.990 131.310 ;
        RECT 129.435 129.580 129.605 131.010 ;
        RECT 134.015 129.580 134.185 131.010 ;
        RECT 138.595 129.580 138.765 131.010 ;
        RECT 143.175 129.580 143.345 131.010 ;
        RECT 147.755 129.580 147.925 131.010 ;
        RECT 129.435 129.490 129.610 129.580 ;
        RECT 134.015 129.490 134.190 129.580 ;
        RECT 138.595 129.490 138.770 129.580 ;
        RECT 143.175 129.490 143.350 129.580 ;
        RECT 147.755 129.490 147.930 129.580 ;
        RECT 116.560 122.710 119.640 127.410 ;
        RECT 129.440 125.540 129.610 129.490 ;
        RECT 134.020 125.540 134.190 129.490 ;
        RECT 138.600 125.540 138.770 129.490 ;
        RECT 143.180 125.540 143.350 129.490 ;
        RECT 147.760 125.540 147.930 129.490 ;
        RECT 126.740 122.710 127.040 123.760 ;
        RECT 131.990 122.710 132.790 123.310 ;
        RECT 138.490 122.710 139.290 123.310 ;
        RECT 191.530 122.710 194.610 127.410 ;
        RECT 205.250 122.710 208.330 127.410 ;
        RECT 218.970 122.710 222.050 127.410 ;
        RECT 232.690 122.710 235.770 127.410 ;
        RECT 246.410 122.710 249.490 127.410 ;
        RECT 112.000 122.410 124.200 122.710 ;
        RECT 126.600 122.410 147.990 122.710 ;
        RECT 149.640 122.410 185.480 122.710 ;
        RECT 186.970 122.410 199.170 122.710 ;
        RECT 200.690 122.410 212.890 122.710 ;
        RECT 214.410 122.410 226.610 122.710 ;
        RECT 228.130 122.410 240.330 122.710 ;
        RECT 241.850 122.410 254.050 122.710 ;
        RECT 123.910 103.910 126.990 108.610 ;
        RECT 140.570 103.910 143.650 108.610 ;
        RECT 154.290 103.910 157.370 108.610 ;
        RECT 170.460 103.910 173.540 108.610 ;
        RECT 191.530 103.910 194.610 108.610 ;
        RECT 205.250 103.910 208.330 108.610 ;
        RECT 246.410 103.910 249.490 108.610 ;
        RECT 119.350 103.610 131.550 103.910 ;
        RECT 136.010 103.610 148.210 103.910 ;
        RECT 149.730 103.610 161.930 103.910 ;
        RECT 165.900 103.610 178.100 103.910 ;
        RECT 186.970 103.610 199.170 103.910 ;
        RECT 200.690 103.610 212.890 103.910 ;
        RECT 241.850 103.610 254.050 103.910 ;
        RECT 123.660 84.810 262.190 85.110 ;
        RECT 223.870 66.310 226.950 71.010 ;
        RECT 237.590 66.310 240.670 71.010 ;
        RECT 251.310 66.310 254.390 71.010 ;
        RECT 219.310 66.010 231.510 66.310 ;
        RECT 233.030 66.010 245.230 66.310 ;
        RECT 246.750 66.010 258.950 66.310 ;
        RECT 223.380 47.510 226.460 52.210 ;
        RECT 237.100 47.510 240.180 52.210 ;
        RECT 250.820 47.510 253.900 52.210 ;
        RECT 218.820 47.210 231.020 47.510 ;
        RECT 232.540 47.210 244.740 47.510 ;
        RECT 246.260 47.210 258.460 47.510 ;
        RECT 227.300 28.710 230.380 33.410 ;
        RECT 236.460 29.135 238.620 31.985 ;
        RECT 241.020 28.710 244.100 33.410 ;
        RECT 254.740 28.710 257.820 33.410 ;
        RECT 222.740 28.410 234.940 28.710 ;
        RECT 236.460 28.410 248.660 28.710 ;
        RECT 250.180 28.410 262.380 28.710 ;
      LAYER mcon ;
        RECT 121.940 242.075 122.110 242.245 ;
        RECT 121.940 241.715 122.110 241.885 ;
        RECT 121.940 241.355 122.110 241.525 ;
        RECT 121.940 240.995 122.110 241.165 ;
        RECT 121.940 240.635 122.110 240.805 ;
        RECT 121.940 240.275 122.110 240.445 ;
        RECT 121.940 239.915 122.110 240.085 ;
        RECT 121.940 239.555 122.110 239.725 ;
        RECT 121.940 239.195 122.110 239.365 ;
        RECT 121.940 238.835 122.110 239.005 ;
        RECT 121.940 238.475 122.110 238.645 ;
        RECT 30.505 235.275 30.675 235.445 ;
        RECT 32.505 235.275 32.675 235.445 ;
        RECT 34.505 235.275 34.675 235.445 ;
        RECT 36.505 235.275 36.675 235.445 ;
        RECT 38.505 235.275 38.675 235.445 ;
        RECT 40.505 235.275 40.675 235.445 ;
        RECT 42.505 235.275 42.675 235.445 ;
        RECT 44.505 235.275 44.675 235.445 ;
        RECT 46.505 235.275 46.675 235.445 ;
        RECT 48.505 235.275 48.675 235.445 ;
        RECT 50.505 235.275 50.675 235.445 ;
        RECT 52.505 235.275 52.675 235.445 ;
        RECT 54.505 235.275 54.675 235.445 ;
        RECT 56.505 235.275 56.675 235.445 ;
        RECT 58.505 235.275 58.675 235.445 ;
        RECT 60.505 235.275 60.675 235.445 ;
        RECT 62.505 235.275 62.675 235.445 ;
        RECT 64.505 235.275 64.675 235.445 ;
        RECT 67.745 235.275 67.915 235.445 ;
        RECT 69.745 235.275 69.915 235.445 ;
        RECT 71.745 235.275 71.915 235.445 ;
        RECT 73.745 235.275 73.915 235.445 ;
        RECT 75.745 235.275 75.915 235.445 ;
        RECT 77.745 235.275 77.915 235.445 ;
        RECT 79.745 235.275 79.915 235.445 ;
        RECT 81.745 235.275 81.915 235.445 ;
        RECT 83.745 235.275 83.915 235.445 ;
        RECT 85.745 235.275 85.915 235.445 ;
        RECT 87.745 235.275 87.915 235.445 ;
        RECT 89.745 235.275 89.915 235.445 ;
        RECT 91.745 235.275 91.915 235.445 ;
        RECT 93.745 235.275 93.915 235.445 ;
        RECT 95.745 235.275 95.915 235.445 ;
        RECT 97.745 235.275 97.915 235.445 ;
        RECT 99.745 235.275 99.915 235.445 ;
        RECT 101.745 235.275 101.915 235.445 ;
        RECT 105.075 235.275 105.245 235.445 ;
        RECT 106.075 235.275 106.245 235.445 ;
        RECT 107.075 235.275 107.245 235.445 ;
        RECT 108.075 235.275 108.245 235.445 ;
        RECT 109.075 235.275 109.245 235.445 ;
        RECT 110.075 235.275 110.245 235.445 ;
        RECT 111.075 235.275 111.245 235.445 ;
        RECT 112.075 235.275 112.245 235.445 ;
        RECT 113.075 235.275 113.245 235.445 ;
        RECT 114.075 235.275 114.245 235.445 ;
        RECT 115.075 235.275 115.245 235.445 ;
        RECT 120.505 235.275 120.675 235.445 ;
        RECT 125.065 235.275 125.235 235.445 ;
        RECT 127.065 235.275 127.235 235.445 ;
        RECT 129.065 235.275 129.235 235.445 ;
        RECT 131.065 235.275 131.235 235.445 ;
        RECT 133.065 235.275 133.235 235.445 ;
        RECT 135.065 235.275 135.235 235.445 ;
        RECT 137.065 235.275 137.235 235.445 ;
        RECT 139.065 235.275 139.235 235.445 ;
        RECT 141.065 235.275 141.235 235.445 ;
        RECT 143.065 235.275 143.235 235.445 ;
        RECT 145.065 235.275 145.235 235.445 ;
        RECT 147.065 235.275 147.235 235.445 ;
        RECT 149.065 235.275 149.235 235.445 ;
        RECT 151.065 235.275 151.235 235.445 ;
        RECT 153.065 235.275 153.235 235.445 ;
        RECT 155.065 235.275 155.235 235.445 ;
        RECT 157.065 235.275 157.235 235.445 ;
        RECT 159.065 235.275 159.235 235.445 ;
        RECT 161.065 235.275 161.235 235.445 ;
        RECT 163.065 235.275 163.235 235.445 ;
        RECT 165.065 235.275 165.235 235.445 ;
        RECT 167.065 235.275 167.235 235.445 ;
        RECT 169.065 235.275 169.235 235.445 ;
        RECT 171.065 235.275 171.235 235.445 ;
        RECT 173.065 235.275 173.235 235.445 ;
        RECT 175.065 235.275 175.235 235.445 ;
        RECT 177.065 235.275 177.235 235.445 ;
        RECT 179.065 235.275 179.235 235.445 ;
        RECT 181.065 235.275 181.235 235.445 ;
        RECT 183.065 235.275 183.235 235.445 ;
        RECT 185.065 235.275 185.235 235.445 ;
        RECT 187.065 235.275 187.235 235.445 ;
        RECT 189.065 235.275 189.235 235.445 ;
        RECT 191.065 235.275 191.235 235.445 ;
        RECT 193.065 235.275 193.235 235.445 ;
        RECT 195.065 235.275 195.235 235.445 ;
        RECT 197.065 235.275 197.235 235.445 ;
        RECT 199.065 235.275 199.235 235.445 ;
        RECT 201.065 235.275 201.235 235.445 ;
        RECT 203.065 235.275 203.235 235.445 ;
        RECT 205.065 235.275 205.235 235.445 ;
        RECT 207.065 235.275 207.235 235.445 ;
        RECT 209.065 235.275 209.235 235.445 ;
        RECT 211.065 235.275 211.235 235.445 ;
        RECT 213.065 235.275 213.235 235.445 ;
        RECT 215.065 235.275 215.235 235.445 ;
        RECT 217.065 235.275 217.235 235.445 ;
        RECT 219.065 235.275 219.235 235.445 ;
        RECT 221.065 235.275 221.235 235.445 ;
        RECT 223.065 235.275 223.235 235.445 ;
        RECT 225.065 235.275 225.235 235.445 ;
        RECT 227.065 235.275 227.235 235.445 ;
        RECT 229.065 235.275 229.235 235.445 ;
        RECT 231.065 235.275 231.235 235.445 ;
        RECT 233.065 235.275 233.235 235.445 ;
        RECT 235.065 235.275 235.235 235.445 ;
        RECT 237.065 235.275 237.235 235.445 ;
        RECT 239.065 235.275 239.235 235.445 ;
        RECT 241.065 235.275 241.235 235.445 ;
        RECT 243.065 235.275 243.235 235.445 ;
        RECT 245.065 235.275 245.235 235.445 ;
        RECT 247.065 235.275 247.235 235.445 ;
        RECT 249.065 235.275 249.235 235.445 ;
        RECT 251.065 235.275 251.235 235.445 ;
        RECT 253.065 235.275 253.235 235.445 ;
        RECT 255.065 235.275 255.235 235.445 ;
        RECT 257.065 235.275 257.235 235.445 ;
        RECT 259.065 235.275 259.235 235.445 ;
        RECT 261.065 235.275 261.235 235.445 ;
        RECT 215.030 224.210 215.200 224.380 ;
        RECT 215.480 224.210 215.650 224.380 ;
        RECT 215.930 224.210 216.100 224.380 ;
        RECT 216.380 224.210 216.550 224.380 ;
        RECT 216.830 224.210 217.000 224.380 ;
        RECT 217.280 224.210 217.450 224.380 ;
        RECT 217.730 224.210 217.900 224.380 ;
        RECT 218.180 224.210 218.350 224.380 ;
        RECT 218.630 224.210 218.800 224.380 ;
        RECT 219.080 224.210 219.250 224.380 ;
        RECT 219.530 224.210 219.700 224.380 ;
        RECT 219.980 224.210 220.150 224.380 ;
        RECT 220.430 224.210 220.600 224.380 ;
        RECT 220.880 224.210 221.050 224.380 ;
        RECT 221.730 224.210 221.900 224.380 ;
        RECT 222.180 224.210 222.350 224.380 ;
        RECT 222.630 224.210 222.800 224.380 ;
        RECT 223.080 224.210 223.250 224.380 ;
        RECT 223.530 224.210 223.700 224.380 ;
        RECT 223.980 224.210 224.150 224.380 ;
        RECT 224.430 224.210 224.600 224.380 ;
        RECT 224.880 224.210 225.050 224.380 ;
        RECT 225.330 224.210 225.500 224.380 ;
        RECT 225.780 224.210 225.950 224.380 ;
        RECT 226.230 224.210 226.400 224.380 ;
        RECT 226.680 224.210 226.850 224.380 ;
        RECT 227.130 224.210 227.300 224.380 ;
        RECT 227.580 224.210 227.750 224.380 ;
        RECT 228.430 224.210 228.600 224.380 ;
        RECT 228.880 224.210 229.050 224.380 ;
        RECT 229.330 224.210 229.500 224.380 ;
        RECT 229.780 224.210 229.950 224.380 ;
        RECT 230.230 224.210 230.400 224.380 ;
        RECT 230.680 224.210 230.850 224.380 ;
        RECT 231.130 224.210 231.300 224.380 ;
        RECT 231.580 224.210 231.750 224.380 ;
        RECT 232.030 224.210 232.200 224.380 ;
        RECT 232.480 224.210 232.650 224.380 ;
        RECT 232.930 224.210 233.100 224.380 ;
        RECT 233.380 224.210 233.550 224.380 ;
        RECT 233.830 224.210 234.000 224.380 ;
        RECT 234.280 224.210 234.450 224.380 ;
        RECT 235.130 224.210 235.300 224.380 ;
        RECT 235.580 224.210 235.750 224.380 ;
        RECT 236.030 224.210 236.200 224.380 ;
        RECT 236.480 224.210 236.650 224.380 ;
        RECT 236.930 224.210 237.100 224.380 ;
        RECT 237.380 224.210 237.550 224.380 ;
        RECT 237.830 224.210 238.000 224.380 ;
        RECT 238.280 224.210 238.450 224.380 ;
        RECT 238.730 224.210 238.900 224.380 ;
        RECT 239.180 224.210 239.350 224.380 ;
        RECT 239.630 224.210 239.800 224.380 ;
        RECT 240.080 224.210 240.250 224.380 ;
        RECT 240.530 224.210 240.700 224.380 ;
        RECT 240.980 224.210 241.150 224.380 ;
        RECT 241.830 224.210 242.000 224.380 ;
        RECT 242.280 224.210 242.450 224.380 ;
        RECT 242.730 224.210 242.900 224.380 ;
        RECT 243.180 224.210 243.350 224.380 ;
        RECT 243.630 224.210 243.800 224.380 ;
        RECT 244.080 224.210 244.250 224.380 ;
        RECT 244.530 224.210 244.700 224.380 ;
        RECT 244.980 224.210 245.150 224.380 ;
        RECT 245.430 224.210 245.600 224.380 ;
        RECT 245.880 224.210 246.050 224.380 ;
        RECT 246.330 224.210 246.500 224.380 ;
        RECT 246.780 224.210 246.950 224.380 ;
        RECT 247.230 224.210 247.400 224.380 ;
        RECT 247.680 224.210 247.850 224.380 ;
        RECT 248.530 224.210 248.700 224.380 ;
        RECT 248.980 224.210 249.150 224.380 ;
        RECT 249.430 224.210 249.600 224.380 ;
        RECT 249.880 224.210 250.050 224.380 ;
        RECT 250.330 224.210 250.500 224.380 ;
        RECT 250.780 224.210 250.950 224.380 ;
        RECT 251.230 224.210 251.400 224.380 ;
        RECT 251.680 224.210 251.850 224.380 ;
        RECT 252.130 224.210 252.300 224.380 ;
        RECT 252.580 224.210 252.750 224.380 ;
        RECT 253.030 224.210 253.200 224.380 ;
        RECT 253.480 224.210 253.650 224.380 ;
        RECT 253.930 224.210 254.100 224.380 ;
        RECT 254.380 224.210 254.550 224.380 ;
        RECT 255.230 224.210 255.400 224.380 ;
        RECT 255.680 224.210 255.850 224.380 ;
        RECT 256.130 224.210 256.300 224.380 ;
        RECT 256.580 224.210 256.750 224.380 ;
        RECT 257.030 224.210 257.200 224.380 ;
        RECT 257.480 224.210 257.650 224.380 ;
        RECT 257.930 224.210 258.100 224.380 ;
        RECT 258.380 224.210 258.550 224.380 ;
        RECT 258.830 224.210 259.000 224.380 ;
        RECT 259.280 224.210 259.450 224.380 ;
        RECT 259.730 224.210 259.900 224.380 ;
        RECT 260.180 224.210 260.350 224.380 ;
        RECT 260.630 224.210 260.800 224.380 ;
        RECT 261.080 224.210 261.250 224.380 ;
        RECT 72.940 223.275 73.110 223.445 ;
        RECT 72.940 222.915 73.110 223.085 ;
        RECT 72.940 222.555 73.110 222.725 ;
        RECT 72.940 222.195 73.110 222.365 ;
        RECT 72.940 221.835 73.110 222.005 ;
        RECT 72.940 221.475 73.110 221.645 ;
        RECT 72.940 221.115 73.110 221.285 ;
        RECT 72.940 220.755 73.110 220.925 ;
        RECT 72.940 220.395 73.110 220.565 ;
        RECT 72.940 220.035 73.110 220.205 ;
        RECT 72.940 219.675 73.110 219.845 ;
        RECT 215.850 223.410 216.020 223.580 ;
        RECT 216.300 223.410 216.470 223.580 ;
        RECT 216.750 223.410 216.920 223.580 ;
        RECT 217.200 223.410 217.370 223.580 ;
        RECT 217.650 223.410 217.820 223.580 ;
        RECT 218.100 223.410 218.270 223.580 ;
        RECT 218.550 223.410 218.720 223.580 ;
        RECT 219.000 223.410 219.170 223.580 ;
        RECT 219.450 223.410 219.620 223.580 ;
        RECT 219.900 223.410 220.070 223.580 ;
        RECT 220.350 223.410 220.520 223.580 ;
        RECT 222.550 223.410 222.720 223.580 ;
        RECT 223.000 223.410 223.170 223.580 ;
        RECT 223.450 223.410 223.620 223.580 ;
        RECT 223.900 223.410 224.070 223.580 ;
        RECT 224.350 223.410 224.520 223.580 ;
        RECT 224.800 223.410 224.970 223.580 ;
        RECT 225.250 223.410 225.420 223.580 ;
        RECT 225.700 223.410 225.870 223.580 ;
        RECT 226.150 223.410 226.320 223.580 ;
        RECT 226.600 223.410 226.770 223.580 ;
        RECT 227.050 223.410 227.220 223.580 ;
        RECT 229.250 223.410 229.420 223.580 ;
        RECT 229.700 223.410 229.870 223.580 ;
        RECT 230.150 223.410 230.320 223.580 ;
        RECT 230.600 223.410 230.770 223.580 ;
        RECT 231.050 223.410 231.220 223.580 ;
        RECT 231.500 223.410 231.670 223.580 ;
        RECT 231.950 223.410 232.120 223.580 ;
        RECT 232.400 223.410 232.570 223.580 ;
        RECT 232.850 223.410 233.020 223.580 ;
        RECT 233.300 223.410 233.470 223.580 ;
        RECT 233.750 223.410 233.920 223.580 ;
        RECT 235.950 223.410 236.120 223.580 ;
        RECT 236.400 223.410 236.570 223.580 ;
        RECT 236.850 223.410 237.020 223.580 ;
        RECT 237.300 223.410 237.470 223.580 ;
        RECT 237.750 223.410 237.920 223.580 ;
        RECT 238.200 223.410 238.370 223.580 ;
        RECT 238.650 223.410 238.820 223.580 ;
        RECT 239.100 223.410 239.270 223.580 ;
        RECT 239.550 223.410 239.720 223.580 ;
        RECT 240.000 223.410 240.170 223.580 ;
        RECT 240.450 223.410 240.620 223.580 ;
        RECT 242.650 223.410 242.820 223.580 ;
        RECT 243.100 223.410 243.270 223.580 ;
        RECT 243.550 223.410 243.720 223.580 ;
        RECT 244.000 223.410 244.170 223.580 ;
        RECT 244.450 223.410 244.620 223.580 ;
        RECT 244.900 223.410 245.070 223.580 ;
        RECT 245.350 223.410 245.520 223.580 ;
        RECT 245.800 223.410 245.970 223.580 ;
        RECT 246.250 223.410 246.420 223.580 ;
        RECT 246.700 223.410 246.870 223.580 ;
        RECT 247.150 223.410 247.320 223.580 ;
        RECT 249.350 223.410 249.520 223.580 ;
        RECT 249.800 223.410 249.970 223.580 ;
        RECT 250.250 223.410 250.420 223.580 ;
        RECT 250.700 223.410 250.870 223.580 ;
        RECT 251.150 223.410 251.320 223.580 ;
        RECT 251.600 223.410 251.770 223.580 ;
        RECT 252.050 223.410 252.220 223.580 ;
        RECT 252.500 223.410 252.670 223.580 ;
        RECT 252.950 223.410 253.120 223.580 ;
        RECT 253.400 223.410 253.570 223.580 ;
        RECT 253.850 223.410 254.020 223.580 ;
        RECT 256.050 223.410 256.220 223.580 ;
        RECT 256.500 223.410 256.670 223.580 ;
        RECT 256.950 223.410 257.120 223.580 ;
        RECT 257.400 223.410 257.570 223.580 ;
        RECT 257.850 223.410 258.020 223.580 ;
        RECT 258.300 223.410 258.470 223.580 ;
        RECT 258.750 223.410 258.920 223.580 ;
        RECT 259.200 223.410 259.370 223.580 ;
        RECT 259.650 223.410 259.820 223.580 ;
        RECT 260.100 223.410 260.270 223.580 ;
        RECT 260.550 223.410 260.720 223.580 ;
        RECT 30.505 216.475 30.675 216.645 ;
        RECT 32.505 216.475 32.675 216.645 ;
        RECT 34.505 216.475 34.675 216.645 ;
        RECT 36.505 216.475 36.675 216.645 ;
        RECT 38.505 216.475 38.675 216.645 ;
        RECT 40.505 216.475 40.675 216.645 ;
        RECT 42.505 216.475 42.675 216.645 ;
        RECT 44.505 216.475 44.675 216.645 ;
        RECT 46.505 216.475 46.675 216.645 ;
        RECT 48.505 216.475 48.675 216.645 ;
        RECT 50.505 216.475 50.675 216.645 ;
        RECT 52.505 216.475 52.675 216.645 ;
        RECT 54.505 216.475 54.675 216.645 ;
        RECT 56.505 216.475 56.675 216.645 ;
        RECT 58.505 216.475 58.675 216.645 ;
        RECT 60.505 216.475 60.675 216.645 ;
        RECT 62.505 216.475 62.675 216.645 ;
        RECT 64.505 216.475 64.675 216.645 ;
        RECT 71.505 216.475 71.675 216.645 ;
        RECT 76.065 216.475 76.235 216.645 ;
        RECT 78.065 216.475 78.235 216.645 ;
        RECT 80.065 216.475 80.235 216.645 ;
        RECT 82.065 216.475 82.235 216.645 ;
        RECT 84.065 216.475 84.235 216.645 ;
        RECT 86.065 216.475 86.235 216.645 ;
        RECT 88.065 216.475 88.235 216.645 ;
        RECT 90.065 216.475 90.235 216.645 ;
        RECT 92.065 216.475 92.235 216.645 ;
        RECT 94.065 216.475 94.235 216.645 ;
        RECT 96.065 216.475 96.235 216.645 ;
        RECT 98.065 216.475 98.235 216.645 ;
        RECT 100.065 216.475 100.235 216.645 ;
        RECT 102.065 216.475 102.235 216.645 ;
        RECT 104.065 216.475 104.235 216.645 ;
        RECT 106.065 216.475 106.235 216.645 ;
        RECT 108.065 216.475 108.235 216.645 ;
        RECT 110.065 216.475 110.235 216.645 ;
        RECT 112.065 216.475 112.235 216.645 ;
        RECT 114.065 216.475 114.235 216.645 ;
        RECT 116.065 216.475 116.235 216.645 ;
        RECT 118.065 216.475 118.235 216.645 ;
        RECT 120.065 216.475 120.235 216.645 ;
        RECT 122.065 216.475 122.235 216.645 ;
        RECT 124.065 216.475 124.235 216.645 ;
        RECT 126.065 216.475 126.235 216.645 ;
        RECT 128.065 216.475 128.235 216.645 ;
        RECT 130.065 216.475 130.235 216.645 ;
        RECT 132.065 216.475 132.235 216.645 ;
        RECT 134.065 216.475 134.235 216.645 ;
        RECT 136.065 216.475 136.235 216.645 ;
        RECT 138.065 216.475 138.235 216.645 ;
        RECT 140.065 216.475 140.235 216.645 ;
        RECT 142.065 216.475 142.235 216.645 ;
        RECT 144.065 216.475 144.235 216.645 ;
        RECT 146.065 216.475 146.235 216.645 ;
        RECT 148.065 216.475 148.235 216.645 ;
        RECT 150.065 216.475 150.235 216.645 ;
        RECT 152.065 216.475 152.235 216.645 ;
        RECT 154.065 216.475 154.235 216.645 ;
        RECT 156.065 216.475 156.235 216.645 ;
        RECT 158.065 216.475 158.235 216.645 ;
        RECT 160.065 216.475 160.235 216.645 ;
        RECT 162.065 216.475 162.235 216.645 ;
        RECT 164.065 216.475 164.235 216.645 ;
        RECT 166.065 216.475 166.235 216.645 ;
        RECT 168.065 216.475 168.235 216.645 ;
        RECT 170.065 216.475 170.235 216.645 ;
        RECT 172.065 216.475 172.235 216.645 ;
        RECT 174.065 216.475 174.235 216.645 ;
        RECT 176.065 216.475 176.235 216.645 ;
        RECT 178.065 216.475 178.235 216.645 ;
        RECT 180.065 216.475 180.235 216.645 ;
        RECT 182.065 216.475 182.235 216.645 ;
        RECT 184.065 216.475 184.235 216.645 ;
        RECT 186.065 216.475 186.235 216.645 ;
        RECT 188.065 216.475 188.235 216.645 ;
        RECT 190.065 216.475 190.235 216.645 ;
        RECT 192.065 216.475 192.235 216.645 ;
        RECT 194.065 216.475 194.235 216.645 ;
        RECT 196.065 216.475 196.235 216.645 ;
        RECT 198.065 216.475 198.235 216.645 ;
        RECT 200.065 216.475 200.235 216.645 ;
        RECT 202.065 216.475 202.235 216.645 ;
        RECT 204.065 216.475 204.235 216.645 ;
        RECT 206.065 216.475 206.235 216.645 ;
        RECT 208.065 216.475 208.235 216.645 ;
        RECT 210.065 216.475 210.235 216.645 ;
        RECT 212.065 216.475 212.235 216.645 ;
        RECT 215.715 216.475 215.885 216.645 ;
        RECT 216.715 216.475 216.885 216.645 ;
        RECT 217.715 216.475 217.885 216.645 ;
        RECT 218.715 216.475 218.885 216.645 ;
        RECT 219.715 216.475 219.885 216.645 ;
        RECT 220.715 216.475 220.885 216.645 ;
        RECT 221.715 216.475 221.885 216.645 ;
        RECT 222.715 216.475 222.885 216.645 ;
        RECT 223.715 216.475 223.885 216.645 ;
        RECT 224.715 216.475 224.885 216.645 ;
        RECT 225.715 216.475 225.885 216.645 ;
        RECT 226.715 216.475 226.885 216.645 ;
        RECT 227.715 216.475 227.885 216.645 ;
        RECT 228.715 216.475 228.885 216.645 ;
        RECT 229.715 216.475 229.885 216.645 ;
        RECT 230.715 216.475 230.885 216.645 ;
        RECT 231.715 216.475 231.885 216.645 ;
        RECT 232.715 216.475 232.885 216.645 ;
        RECT 233.715 216.475 233.885 216.645 ;
        RECT 234.715 216.475 234.885 216.645 ;
        RECT 235.715 216.475 235.885 216.645 ;
        RECT 236.715 216.475 236.885 216.645 ;
        RECT 237.715 216.475 237.885 216.645 ;
        RECT 238.715 216.475 238.885 216.645 ;
        RECT 239.715 216.475 239.885 216.645 ;
        RECT 240.715 216.475 240.885 216.645 ;
        RECT 241.715 216.475 241.885 216.645 ;
        RECT 242.715 216.475 242.885 216.645 ;
        RECT 243.715 216.475 243.885 216.645 ;
        RECT 244.715 216.475 244.885 216.645 ;
        RECT 245.715 216.475 245.885 216.645 ;
        RECT 246.715 216.475 246.885 216.645 ;
        RECT 247.715 216.475 247.885 216.645 ;
        RECT 248.715 216.475 248.885 216.645 ;
        RECT 249.715 216.475 249.885 216.645 ;
        RECT 250.715 216.475 250.885 216.645 ;
        RECT 251.715 216.475 251.885 216.645 ;
        RECT 252.715 216.475 252.885 216.645 ;
        RECT 253.715 216.475 253.885 216.645 ;
        RECT 254.715 216.475 254.885 216.645 ;
        RECT 255.715 216.475 255.885 216.645 ;
        RECT 256.715 216.475 256.885 216.645 ;
        RECT 257.715 216.475 257.885 216.645 ;
        RECT 258.715 216.475 258.885 216.645 ;
        RECT 259.715 216.475 259.885 216.645 ;
        RECT 260.715 216.475 260.885 216.645 ;
        RECT 209.150 205.410 209.320 205.580 ;
        RECT 209.600 205.410 209.770 205.580 ;
        RECT 210.050 205.410 210.220 205.580 ;
        RECT 210.500 205.410 210.670 205.580 ;
        RECT 210.950 205.410 211.120 205.580 ;
        RECT 211.400 205.410 211.570 205.580 ;
        RECT 211.850 205.410 212.020 205.580 ;
        RECT 212.300 205.410 212.470 205.580 ;
        RECT 212.750 205.410 212.920 205.580 ;
        RECT 213.200 205.410 213.370 205.580 ;
        RECT 213.650 205.410 213.820 205.580 ;
        RECT 214.100 205.410 214.270 205.580 ;
        RECT 214.550 205.410 214.720 205.580 ;
        RECT 215.000 205.410 215.170 205.580 ;
        RECT 215.850 205.410 216.020 205.580 ;
        RECT 216.300 205.410 216.470 205.580 ;
        RECT 216.750 205.410 216.920 205.580 ;
        RECT 217.200 205.410 217.370 205.580 ;
        RECT 217.650 205.410 217.820 205.580 ;
        RECT 218.100 205.410 218.270 205.580 ;
        RECT 218.550 205.410 218.720 205.580 ;
        RECT 219.000 205.410 219.170 205.580 ;
        RECT 219.450 205.410 219.620 205.580 ;
        RECT 219.900 205.410 220.070 205.580 ;
        RECT 220.350 205.410 220.520 205.580 ;
        RECT 220.800 205.410 220.970 205.580 ;
        RECT 221.250 205.410 221.420 205.580 ;
        RECT 221.700 205.410 221.870 205.580 ;
        RECT 222.550 205.410 222.720 205.580 ;
        RECT 223.000 205.410 223.170 205.580 ;
        RECT 223.450 205.410 223.620 205.580 ;
        RECT 223.900 205.410 224.070 205.580 ;
        RECT 224.350 205.410 224.520 205.580 ;
        RECT 224.800 205.410 224.970 205.580 ;
        RECT 225.250 205.410 225.420 205.580 ;
        RECT 225.700 205.410 225.870 205.580 ;
        RECT 226.150 205.410 226.320 205.580 ;
        RECT 226.600 205.410 226.770 205.580 ;
        RECT 227.050 205.410 227.220 205.580 ;
        RECT 227.500 205.410 227.670 205.580 ;
        RECT 227.950 205.410 228.120 205.580 ;
        RECT 228.400 205.410 228.570 205.580 ;
        RECT 229.250 205.410 229.420 205.580 ;
        RECT 229.700 205.410 229.870 205.580 ;
        RECT 230.150 205.410 230.320 205.580 ;
        RECT 230.600 205.410 230.770 205.580 ;
        RECT 231.050 205.410 231.220 205.580 ;
        RECT 231.500 205.410 231.670 205.580 ;
        RECT 231.950 205.410 232.120 205.580 ;
        RECT 232.400 205.410 232.570 205.580 ;
        RECT 232.850 205.410 233.020 205.580 ;
        RECT 233.300 205.410 233.470 205.580 ;
        RECT 233.750 205.410 233.920 205.580 ;
        RECT 234.200 205.410 234.370 205.580 ;
        RECT 234.650 205.410 234.820 205.580 ;
        RECT 235.100 205.410 235.270 205.580 ;
        RECT 235.950 205.410 236.120 205.580 ;
        RECT 236.400 205.410 236.570 205.580 ;
        RECT 236.850 205.410 237.020 205.580 ;
        RECT 237.300 205.410 237.470 205.580 ;
        RECT 237.750 205.410 237.920 205.580 ;
        RECT 238.200 205.410 238.370 205.580 ;
        RECT 238.650 205.410 238.820 205.580 ;
        RECT 239.100 205.410 239.270 205.580 ;
        RECT 239.550 205.410 239.720 205.580 ;
        RECT 240.000 205.410 240.170 205.580 ;
        RECT 240.450 205.410 240.620 205.580 ;
        RECT 240.900 205.410 241.070 205.580 ;
        RECT 241.350 205.410 241.520 205.580 ;
        RECT 241.800 205.410 241.970 205.580 ;
        RECT 242.650 205.410 242.820 205.580 ;
        RECT 243.100 205.410 243.270 205.580 ;
        RECT 243.550 205.410 243.720 205.580 ;
        RECT 244.000 205.410 244.170 205.580 ;
        RECT 244.450 205.410 244.620 205.580 ;
        RECT 244.900 205.410 245.070 205.580 ;
        RECT 245.350 205.410 245.520 205.580 ;
        RECT 245.800 205.410 245.970 205.580 ;
        RECT 246.250 205.410 246.420 205.580 ;
        RECT 246.700 205.410 246.870 205.580 ;
        RECT 247.150 205.410 247.320 205.580 ;
        RECT 247.600 205.410 247.770 205.580 ;
        RECT 248.050 205.410 248.220 205.580 ;
        RECT 248.500 205.410 248.670 205.580 ;
        RECT 249.350 205.410 249.520 205.580 ;
        RECT 249.800 205.410 249.970 205.580 ;
        RECT 250.250 205.410 250.420 205.580 ;
        RECT 250.700 205.410 250.870 205.580 ;
        RECT 251.150 205.410 251.320 205.580 ;
        RECT 251.600 205.410 251.770 205.580 ;
        RECT 252.050 205.410 252.220 205.580 ;
        RECT 252.500 205.410 252.670 205.580 ;
        RECT 252.950 205.410 253.120 205.580 ;
        RECT 253.400 205.410 253.570 205.580 ;
        RECT 253.850 205.410 254.020 205.580 ;
        RECT 254.300 205.410 254.470 205.580 ;
        RECT 254.750 205.410 254.920 205.580 ;
        RECT 255.200 205.410 255.370 205.580 ;
        RECT 256.050 205.410 256.220 205.580 ;
        RECT 256.500 205.410 256.670 205.580 ;
        RECT 256.950 205.410 257.120 205.580 ;
        RECT 257.400 205.410 257.570 205.580 ;
        RECT 257.850 205.410 258.020 205.580 ;
        RECT 258.300 205.410 258.470 205.580 ;
        RECT 258.750 205.410 258.920 205.580 ;
        RECT 259.200 205.410 259.370 205.580 ;
        RECT 259.650 205.410 259.820 205.580 ;
        RECT 260.100 205.410 260.270 205.580 ;
        RECT 260.550 205.410 260.720 205.580 ;
        RECT 261.000 205.410 261.170 205.580 ;
        RECT 261.450 205.410 261.620 205.580 ;
        RECT 261.900 205.410 262.070 205.580 ;
        RECT 209.970 204.610 210.140 204.780 ;
        RECT 210.420 204.610 210.590 204.780 ;
        RECT 210.870 204.610 211.040 204.780 ;
        RECT 211.320 204.610 211.490 204.780 ;
        RECT 211.770 204.610 211.940 204.780 ;
        RECT 212.220 204.610 212.390 204.780 ;
        RECT 212.670 204.610 212.840 204.780 ;
        RECT 213.120 204.610 213.290 204.780 ;
        RECT 213.570 204.610 213.740 204.780 ;
        RECT 214.020 204.610 214.190 204.780 ;
        RECT 214.470 204.610 214.640 204.780 ;
        RECT 216.670 204.610 216.840 204.780 ;
        RECT 217.120 204.610 217.290 204.780 ;
        RECT 217.570 204.610 217.740 204.780 ;
        RECT 218.020 204.610 218.190 204.780 ;
        RECT 218.470 204.610 218.640 204.780 ;
        RECT 218.920 204.610 219.090 204.780 ;
        RECT 219.370 204.610 219.540 204.780 ;
        RECT 219.820 204.610 219.990 204.780 ;
        RECT 220.270 204.610 220.440 204.780 ;
        RECT 220.720 204.610 220.890 204.780 ;
        RECT 221.170 204.610 221.340 204.780 ;
        RECT 223.370 204.610 223.540 204.780 ;
        RECT 223.820 204.610 223.990 204.780 ;
        RECT 224.270 204.610 224.440 204.780 ;
        RECT 224.720 204.610 224.890 204.780 ;
        RECT 225.170 204.610 225.340 204.780 ;
        RECT 225.620 204.610 225.790 204.780 ;
        RECT 226.070 204.610 226.240 204.780 ;
        RECT 226.520 204.610 226.690 204.780 ;
        RECT 226.970 204.610 227.140 204.780 ;
        RECT 227.420 204.610 227.590 204.780 ;
        RECT 227.870 204.610 228.040 204.780 ;
        RECT 230.070 204.610 230.240 204.780 ;
        RECT 230.520 204.610 230.690 204.780 ;
        RECT 230.970 204.610 231.140 204.780 ;
        RECT 231.420 204.610 231.590 204.780 ;
        RECT 231.870 204.610 232.040 204.780 ;
        RECT 232.320 204.610 232.490 204.780 ;
        RECT 232.770 204.610 232.940 204.780 ;
        RECT 233.220 204.610 233.390 204.780 ;
        RECT 233.670 204.610 233.840 204.780 ;
        RECT 234.120 204.610 234.290 204.780 ;
        RECT 234.570 204.610 234.740 204.780 ;
        RECT 236.770 204.610 236.940 204.780 ;
        RECT 237.220 204.610 237.390 204.780 ;
        RECT 237.670 204.610 237.840 204.780 ;
        RECT 238.120 204.610 238.290 204.780 ;
        RECT 238.570 204.610 238.740 204.780 ;
        RECT 239.020 204.610 239.190 204.780 ;
        RECT 239.470 204.610 239.640 204.780 ;
        RECT 239.920 204.610 240.090 204.780 ;
        RECT 240.370 204.610 240.540 204.780 ;
        RECT 240.820 204.610 240.990 204.780 ;
        RECT 241.270 204.610 241.440 204.780 ;
        RECT 243.470 204.610 243.640 204.780 ;
        RECT 243.920 204.610 244.090 204.780 ;
        RECT 244.370 204.610 244.540 204.780 ;
        RECT 244.820 204.610 244.990 204.780 ;
        RECT 245.270 204.610 245.440 204.780 ;
        RECT 245.720 204.610 245.890 204.780 ;
        RECT 246.170 204.610 246.340 204.780 ;
        RECT 246.620 204.610 246.790 204.780 ;
        RECT 247.070 204.610 247.240 204.780 ;
        RECT 247.520 204.610 247.690 204.780 ;
        RECT 247.970 204.610 248.140 204.780 ;
        RECT 250.170 204.610 250.340 204.780 ;
        RECT 250.620 204.610 250.790 204.780 ;
        RECT 251.070 204.610 251.240 204.780 ;
        RECT 251.520 204.610 251.690 204.780 ;
        RECT 251.970 204.610 252.140 204.780 ;
        RECT 252.420 204.610 252.590 204.780 ;
        RECT 252.870 204.610 253.040 204.780 ;
        RECT 253.320 204.610 253.490 204.780 ;
        RECT 253.770 204.610 253.940 204.780 ;
        RECT 254.220 204.610 254.390 204.780 ;
        RECT 254.670 204.610 254.840 204.780 ;
        RECT 256.870 204.610 257.040 204.780 ;
        RECT 257.320 204.610 257.490 204.780 ;
        RECT 257.770 204.610 257.940 204.780 ;
        RECT 258.220 204.610 258.390 204.780 ;
        RECT 258.670 204.610 258.840 204.780 ;
        RECT 259.120 204.610 259.290 204.780 ;
        RECT 259.570 204.610 259.740 204.780 ;
        RECT 260.020 204.610 260.190 204.780 ;
        RECT 260.470 204.610 260.640 204.780 ;
        RECT 260.920 204.610 261.090 204.780 ;
        RECT 261.370 204.610 261.540 204.780 ;
        RECT 32.465 197.675 32.635 197.845 ;
        RECT 34.465 197.675 34.635 197.845 ;
        RECT 36.465 197.675 36.635 197.845 ;
        RECT 38.465 197.675 38.635 197.845 ;
        RECT 40.465 197.675 40.635 197.845 ;
        RECT 42.465 197.675 42.635 197.845 ;
        RECT 44.465 197.675 44.635 197.845 ;
        RECT 46.465 197.675 46.635 197.845 ;
        RECT 48.465 197.675 48.635 197.845 ;
        RECT 50.465 197.675 50.635 197.845 ;
        RECT 52.465 197.675 52.635 197.845 ;
        RECT 54.465 197.675 54.635 197.845 ;
        RECT 56.465 197.675 56.635 197.845 ;
        RECT 58.465 197.675 58.635 197.845 ;
        RECT 60.465 197.675 60.635 197.845 ;
        RECT 62.465 197.675 62.635 197.845 ;
        RECT 64.465 197.675 64.635 197.845 ;
        RECT 66.465 197.675 66.635 197.845 ;
        RECT 76.565 197.675 76.735 197.845 ;
        RECT 78.565 197.675 78.735 197.845 ;
        RECT 80.565 197.675 80.735 197.845 ;
        RECT 82.565 197.675 82.735 197.845 ;
        RECT 84.565 197.675 84.735 197.845 ;
        RECT 86.565 197.675 86.735 197.845 ;
        RECT 88.565 197.675 88.735 197.845 ;
        RECT 90.565 197.675 90.735 197.845 ;
        RECT 92.565 197.675 92.735 197.845 ;
        RECT 94.565 197.675 94.735 197.845 ;
        RECT 96.565 197.675 96.735 197.845 ;
        RECT 98.565 197.675 98.735 197.845 ;
        RECT 100.565 197.675 100.735 197.845 ;
        RECT 102.565 197.675 102.735 197.845 ;
        RECT 104.565 197.675 104.735 197.845 ;
        RECT 106.565 197.675 106.735 197.845 ;
        RECT 108.565 197.675 108.735 197.845 ;
        RECT 110.565 197.675 110.735 197.845 ;
        RECT 114.285 197.675 114.455 197.845 ;
        RECT 116.285 197.675 116.455 197.845 ;
        RECT 118.285 197.675 118.455 197.845 ;
        RECT 120.285 197.675 120.455 197.845 ;
        RECT 122.285 197.675 122.455 197.845 ;
        RECT 124.285 197.675 124.455 197.845 ;
        RECT 126.285 197.675 126.455 197.845 ;
        RECT 128.285 197.675 128.455 197.845 ;
        RECT 130.285 197.675 130.455 197.845 ;
        RECT 132.285 197.675 132.455 197.845 ;
        RECT 134.285 197.675 134.455 197.845 ;
        RECT 136.285 197.675 136.455 197.845 ;
        RECT 138.285 197.675 138.455 197.845 ;
        RECT 140.285 197.675 140.455 197.845 ;
        RECT 147.605 197.675 147.775 197.845 ;
        RECT 149.605 197.675 149.775 197.845 ;
        RECT 151.605 197.675 151.775 197.845 ;
        RECT 153.605 197.675 153.775 197.845 ;
        RECT 155.605 197.675 155.775 197.845 ;
        RECT 157.605 197.675 157.775 197.845 ;
        RECT 159.605 197.675 159.775 197.845 ;
        RECT 161.605 197.675 161.775 197.845 ;
        RECT 163.605 197.675 163.775 197.845 ;
        RECT 165.605 197.675 165.775 197.845 ;
        RECT 167.605 197.675 167.775 197.845 ;
        RECT 169.605 197.675 169.775 197.845 ;
        RECT 171.605 197.675 171.775 197.845 ;
        RECT 173.605 197.675 173.775 197.845 ;
        RECT 187.295 197.675 187.465 197.845 ;
        RECT 189.295 197.675 189.465 197.845 ;
        RECT 191.295 197.675 191.465 197.845 ;
        RECT 193.295 197.675 193.465 197.845 ;
        RECT 195.295 197.675 195.465 197.845 ;
        RECT 197.295 197.675 197.465 197.845 ;
        RECT 199.295 197.675 199.465 197.845 ;
        RECT 201.295 197.675 201.465 197.845 ;
        RECT 203.295 197.675 203.465 197.845 ;
        RECT 205.295 197.675 205.465 197.845 ;
        RECT 209.835 197.675 210.005 197.845 ;
        RECT 210.835 197.675 211.005 197.845 ;
        RECT 211.835 197.675 212.005 197.845 ;
        RECT 212.835 197.675 213.005 197.845 ;
        RECT 213.835 197.675 214.005 197.845 ;
        RECT 214.835 197.675 215.005 197.845 ;
        RECT 215.835 197.675 216.005 197.845 ;
        RECT 216.835 197.675 217.005 197.845 ;
        RECT 217.835 197.675 218.005 197.845 ;
        RECT 218.835 197.675 219.005 197.845 ;
        RECT 219.835 197.675 220.005 197.845 ;
        RECT 220.835 197.675 221.005 197.845 ;
        RECT 221.835 197.675 222.005 197.845 ;
        RECT 222.835 197.675 223.005 197.845 ;
        RECT 223.835 197.675 224.005 197.845 ;
        RECT 224.835 197.675 225.005 197.845 ;
        RECT 225.835 197.675 226.005 197.845 ;
        RECT 226.835 197.675 227.005 197.845 ;
        RECT 227.835 197.675 228.005 197.845 ;
        RECT 228.835 197.675 229.005 197.845 ;
        RECT 229.835 197.675 230.005 197.845 ;
        RECT 230.835 197.675 231.005 197.845 ;
        RECT 231.835 197.675 232.005 197.845 ;
        RECT 232.835 197.675 233.005 197.845 ;
        RECT 233.835 197.675 234.005 197.845 ;
        RECT 234.835 197.675 235.005 197.845 ;
        RECT 235.835 197.675 236.005 197.845 ;
        RECT 236.835 197.675 237.005 197.845 ;
        RECT 237.835 197.675 238.005 197.845 ;
        RECT 238.835 197.675 239.005 197.845 ;
        RECT 239.835 197.675 240.005 197.845 ;
        RECT 240.835 197.675 241.005 197.845 ;
        RECT 241.835 197.675 242.005 197.845 ;
        RECT 242.835 197.675 243.005 197.845 ;
        RECT 243.835 197.675 244.005 197.845 ;
        RECT 244.835 197.675 245.005 197.845 ;
        RECT 245.835 197.675 246.005 197.845 ;
        RECT 246.835 197.675 247.005 197.845 ;
        RECT 247.835 197.675 248.005 197.845 ;
        RECT 248.835 197.675 249.005 197.845 ;
        RECT 249.835 197.675 250.005 197.845 ;
        RECT 250.835 197.675 251.005 197.845 ;
        RECT 251.835 197.675 252.005 197.845 ;
        RECT 252.835 197.675 253.005 197.845 ;
        RECT 253.835 197.675 254.005 197.845 ;
        RECT 254.835 197.675 255.005 197.845 ;
        RECT 255.835 197.675 256.005 197.845 ;
        RECT 256.835 197.675 257.005 197.845 ;
        RECT 257.835 197.675 258.005 197.845 ;
        RECT 258.835 197.675 259.005 197.845 ;
        RECT 259.835 197.675 260.005 197.845 ;
        RECT 260.835 197.675 261.005 197.845 ;
        RECT 261.835 197.675 262.005 197.845 ;
        RECT 65.465 181.305 65.635 181.475 ;
        RECT 209.150 186.610 209.320 186.780 ;
        RECT 209.600 186.610 209.770 186.780 ;
        RECT 210.050 186.610 210.220 186.780 ;
        RECT 210.500 186.610 210.670 186.780 ;
        RECT 210.950 186.610 211.120 186.780 ;
        RECT 211.400 186.610 211.570 186.780 ;
        RECT 211.850 186.610 212.020 186.780 ;
        RECT 212.300 186.610 212.470 186.780 ;
        RECT 212.750 186.610 212.920 186.780 ;
        RECT 213.200 186.610 213.370 186.780 ;
        RECT 213.650 186.610 213.820 186.780 ;
        RECT 214.100 186.610 214.270 186.780 ;
        RECT 214.550 186.610 214.720 186.780 ;
        RECT 215.000 186.610 215.170 186.780 ;
        RECT 215.850 186.610 216.020 186.780 ;
        RECT 216.300 186.610 216.470 186.780 ;
        RECT 216.750 186.610 216.920 186.780 ;
        RECT 217.200 186.610 217.370 186.780 ;
        RECT 217.650 186.610 217.820 186.780 ;
        RECT 218.100 186.610 218.270 186.780 ;
        RECT 218.550 186.610 218.720 186.780 ;
        RECT 219.000 186.610 219.170 186.780 ;
        RECT 219.450 186.610 219.620 186.780 ;
        RECT 219.900 186.610 220.070 186.780 ;
        RECT 220.350 186.610 220.520 186.780 ;
        RECT 220.800 186.610 220.970 186.780 ;
        RECT 221.250 186.610 221.420 186.780 ;
        RECT 221.700 186.610 221.870 186.780 ;
        RECT 222.550 186.610 222.720 186.780 ;
        RECT 223.000 186.610 223.170 186.780 ;
        RECT 223.450 186.610 223.620 186.780 ;
        RECT 223.900 186.610 224.070 186.780 ;
        RECT 224.350 186.610 224.520 186.780 ;
        RECT 224.800 186.610 224.970 186.780 ;
        RECT 225.250 186.610 225.420 186.780 ;
        RECT 225.700 186.610 225.870 186.780 ;
        RECT 226.150 186.610 226.320 186.780 ;
        RECT 226.600 186.610 226.770 186.780 ;
        RECT 227.050 186.610 227.220 186.780 ;
        RECT 227.500 186.610 227.670 186.780 ;
        RECT 227.950 186.610 228.120 186.780 ;
        RECT 228.400 186.610 228.570 186.780 ;
        RECT 229.250 186.610 229.420 186.780 ;
        RECT 229.700 186.610 229.870 186.780 ;
        RECT 230.150 186.610 230.320 186.780 ;
        RECT 230.600 186.610 230.770 186.780 ;
        RECT 231.050 186.610 231.220 186.780 ;
        RECT 231.500 186.610 231.670 186.780 ;
        RECT 231.950 186.610 232.120 186.780 ;
        RECT 232.400 186.610 232.570 186.780 ;
        RECT 232.850 186.610 233.020 186.780 ;
        RECT 233.300 186.610 233.470 186.780 ;
        RECT 233.750 186.610 233.920 186.780 ;
        RECT 234.200 186.610 234.370 186.780 ;
        RECT 234.650 186.610 234.820 186.780 ;
        RECT 235.100 186.610 235.270 186.780 ;
        RECT 235.950 186.610 236.120 186.780 ;
        RECT 236.400 186.610 236.570 186.780 ;
        RECT 236.850 186.610 237.020 186.780 ;
        RECT 237.300 186.610 237.470 186.780 ;
        RECT 237.750 186.610 237.920 186.780 ;
        RECT 238.200 186.610 238.370 186.780 ;
        RECT 238.650 186.610 238.820 186.780 ;
        RECT 239.100 186.610 239.270 186.780 ;
        RECT 239.550 186.610 239.720 186.780 ;
        RECT 240.000 186.610 240.170 186.780 ;
        RECT 240.450 186.610 240.620 186.780 ;
        RECT 240.900 186.610 241.070 186.780 ;
        RECT 241.350 186.610 241.520 186.780 ;
        RECT 241.800 186.610 241.970 186.780 ;
        RECT 242.650 186.610 242.820 186.780 ;
        RECT 243.100 186.610 243.270 186.780 ;
        RECT 243.550 186.610 243.720 186.780 ;
        RECT 244.000 186.610 244.170 186.780 ;
        RECT 244.450 186.610 244.620 186.780 ;
        RECT 244.900 186.610 245.070 186.780 ;
        RECT 245.350 186.610 245.520 186.780 ;
        RECT 245.800 186.610 245.970 186.780 ;
        RECT 246.250 186.610 246.420 186.780 ;
        RECT 246.700 186.610 246.870 186.780 ;
        RECT 247.150 186.610 247.320 186.780 ;
        RECT 247.600 186.610 247.770 186.780 ;
        RECT 248.050 186.610 248.220 186.780 ;
        RECT 248.500 186.610 248.670 186.780 ;
        RECT 249.350 186.610 249.520 186.780 ;
        RECT 249.800 186.610 249.970 186.780 ;
        RECT 250.250 186.610 250.420 186.780 ;
        RECT 250.700 186.610 250.870 186.780 ;
        RECT 251.150 186.610 251.320 186.780 ;
        RECT 251.600 186.610 251.770 186.780 ;
        RECT 252.050 186.610 252.220 186.780 ;
        RECT 252.500 186.610 252.670 186.780 ;
        RECT 252.950 186.610 253.120 186.780 ;
        RECT 253.400 186.610 253.570 186.780 ;
        RECT 253.850 186.610 254.020 186.780 ;
        RECT 254.300 186.610 254.470 186.780 ;
        RECT 254.750 186.610 254.920 186.780 ;
        RECT 255.200 186.610 255.370 186.780 ;
        RECT 256.050 186.610 256.220 186.780 ;
        RECT 256.500 186.610 256.670 186.780 ;
        RECT 256.950 186.610 257.120 186.780 ;
        RECT 257.400 186.610 257.570 186.780 ;
        RECT 257.850 186.610 258.020 186.780 ;
        RECT 258.300 186.610 258.470 186.780 ;
        RECT 258.750 186.610 258.920 186.780 ;
        RECT 259.200 186.610 259.370 186.780 ;
        RECT 259.650 186.610 259.820 186.780 ;
        RECT 260.100 186.610 260.270 186.780 ;
        RECT 260.550 186.610 260.720 186.780 ;
        RECT 261.000 186.610 261.170 186.780 ;
        RECT 261.450 186.610 261.620 186.780 ;
        RECT 261.900 186.610 262.070 186.780 ;
        RECT 66.385 180.625 66.555 180.795 ;
        RECT 95.930 179.615 97.900 182.305 ;
        RECT 209.970 185.810 210.140 185.980 ;
        RECT 210.420 185.810 210.590 185.980 ;
        RECT 210.870 185.810 211.040 185.980 ;
        RECT 211.320 185.810 211.490 185.980 ;
        RECT 211.770 185.810 211.940 185.980 ;
        RECT 212.220 185.810 212.390 185.980 ;
        RECT 212.670 185.810 212.840 185.980 ;
        RECT 213.120 185.810 213.290 185.980 ;
        RECT 213.570 185.810 213.740 185.980 ;
        RECT 214.020 185.810 214.190 185.980 ;
        RECT 214.470 185.810 214.640 185.980 ;
        RECT 216.670 185.810 216.840 185.980 ;
        RECT 217.120 185.810 217.290 185.980 ;
        RECT 217.570 185.810 217.740 185.980 ;
        RECT 218.020 185.810 218.190 185.980 ;
        RECT 218.470 185.810 218.640 185.980 ;
        RECT 218.920 185.810 219.090 185.980 ;
        RECT 219.370 185.810 219.540 185.980 ;
        RECT 219.820 185.810 219.990 185.980 ;
        RECT 220.270 185.810 220.440 185.980 ;
        RECT 220.720 185.810 220.890 185.980 ;
        RECT 221.170 185.810 221.340 185.980 ;
        RECT 223.370 185.810 223.540 185.980 ;
        RECT 223.820 185.810 223.990 185.980 ;
        RECT 224.270 185.810 224.440 185.980 ;
        RECT 224.720 185.810 224.890 185.980 ;
        RECT 225.170 185.810 225.340 185.980 ;
        RECT 225.620 185.810 225.790 185.980 ;
        RECT 226.070 185.810 226.240 185.980 ;
        RECT 226.520 185.810 226.690 185.980 ;
        RECT 226.970 185.810 227.140 185.980 ;
        RECT 227.420 185.810 227.590 185.980 ;
        RECT 227.870 185.810 228.040 185.980 ;
        RECT 230.070 185.810 230.240 185.980 ;
        RECT 230.520 185.810 230.690 185.980 ;
        RECT 230.970 185.810 231.140 185.980 ;
        RECT 231.420 185.810 231.590 185.980 ;
        RECT 231.870 185.810 232.040 185.980 ;
        RECT 232.320 185.810 232.490 185.980 ;
        RECT 232.770 185.810 232.940 185.980 ;
        RECT 233.220 185.810 233.390 185.980 ;
        RECT 233.670 185.810 233.840 185.980 ;
        RECT 234.120 185.810 234.290 185.980 ;
        RECT 234.570 185.810 234.740 185.980 ;
        RECT 236.770 185.810 236.940 185.980 ;
        RECT 237.220 185.810 237.390 185.980 ;
        RECT 237.670 185.810 237.840 185.980 ;
        RECT 238.120 185.810 238.290 185.980 ;
        RECT 238.570 185.810 238.740 185.980 ;
        RECT 239.020 185.810 239.190 185.980 ;
        RECT 239.470 185.810 239.640 185.980 ;
        RECT 239.920 185.810 240.090 185.980 ;
        RECT 240.370 185.810 240.540 185.980 ;
        RECT 240.820 185.810 240.990 185.980 ;
        RECT 241.270 185.810 241.440 185.980 ;
        RECT 243.470 185.810 243.640 185.980 ;
        RECT 243.920 185.810 244.090 185.980 ;
        RECT 244.370 185.810 244.540 185.980 ;
        RECT 244.820 185.810 244.990 185.980 ;
        RECT 245.270 185.810 245.440 185.980 ;
        RECT 245.720 185.810 245.890 185.980 ;
        RECT 246.170 185.810 246.340 185.980 ;
        RECT 246.620 185.810 246.790 185.980 ;
        RECT 247.070 185.810 247.240 185.980 ;
        RECT 247.520 185.810 247.690 185.980 ;
        RECT 247.970 185.810 248.140 185.980 ;
        RECT 250.170 185.810 250.340 185.980 ;
        RECT 250.620 185.810 250.790 185.980 ;
        RECT 251.070 185.810 251.240 185.980 ;
        RECT 251.520 185.810 251.690 185.980 ;
        RECT 251.970 185.810 252.140 185.980 ;
        RECT 252.420 185.810 252.590 185.980 ;
        RECT 252.870 185.810 253.040 185.980 ;
        RECT 253.320 185.810 253.490 185.980 ;
        RECT 253.770 185.810 253.940 185.980 ;
        RECT 254.220 185.810 254.390 185.980 ;
        RECT 254.670 185.810 254.840 185.980 ;
        RECT 256.870 185.810 257.040 185.980 ;
        RECT 257.320 185.810 257.490 185.980 ;
        RECT 257.770 185.810 257.940 185.980 ;
        RECT 258.220 185.810 258.390 185.980 ;
        RECT 258.670 185.810 258.840 185.980 ;
        RECT 259.120 185.810 259.290 185.980 ;
        RECT 259.570 185.810 259.740 185.980 ;
        RECT 260.020 185.810 260.190 185.980 ;
        RECT 260.470 185.810 260.640 185.980 ;
        RECT 260.920 185.810 261.090 185.980 ;
        RECT 261.370 185.810 261.540 185.980 ;
        RECT 60.875 178.875 61.045 179.045 ;
        RECT 61.875 178.875 62.045 179.045 ;
        RECT 62.875 178.875 63.045 179.045 ;
        RECT 63.875 178.875 64.045 179.045 ;
        RECT 64.875 178.875 65.045 179.045 ;
        RECT 65.875 178.875 66.045 179.045 ;
        RECT 69.305 178.875 69.475 179.045 ;
        RECT 70.305 178.875 70.475 179.045 ;
        RECT 71.305 178.875 71.475 179.045 ;
        RECT 72.305 178.875 72.475 179.045 ;
        RECT 73.305 178.875 73.475 179.045 ;
        RECT 74.305 178.875 74.475 179.045 ;
        RECT 75.305 178.875 75.475 179.045 ;
        RECT 76.305 178.875 76.475 179.045 ;
        RECT 77.305 178.875 77.475 179.045 ;
        RECT 78.305 178.875 78.475 179.045 ;
        RECT 79.305 178.875 79.475 179.045 ;
        RECT 83.025 178.875 83.195 179.045 ;
        RECT 84.025 178.875 84.195 179.045 ;
        RECT 85.025 178.875 85.195 179.045 ;
        RECT 86.025 178.875 86.195 179.045 ;
        RECT 87.025 178.875 87.195 179.045 ;
        RECT 88.025 178.875 88.195 179.045 ;
        RECT 89.025 178.875 89.195 179.045 ;
        RECT 90.025 178.875 90.195 179.045 ;
        RECT 91.025 178.875 91.195 179.045 ;
        RECT 92.025 178.875 92.195 179.045 ;
        RECT 93.025 178.875 93.195 179.045 ;
        RECT 96.755 178.875 96.925 179.045 ;
        RECT 97.755 178.875 97.925 179.045 ;
        RECT 98.755 178.875 98.925 179.045 ;
        RECT 99.755 178.875 99.925 179.045 ;
        RECT 100.755 178.875 100.925 179.045 ;
        RECT 101.755 178.875 101.925 179.045 ;
        RECT 102.755 178.875 102.925 179.045 ;
        RECT 103.755 178.875 103.925 179.045 ;
        RECT 104.755 178.875 104.925 179.045 ;
        RECT 105.755 178.875 105.925 179.045 ;
        RECT 106.755 178.875 106.925 179.045 ;
        RECT 107.755 178.875 107.925 179.045 ;
        RECT 108.755 178.875 108.925 179.045 ;
        RECT 109.755 178.875 109.925 179.045 ;
        RECT 113.405 178.875 113.575 179.045 ;
        RECT 114.405 178.875 114.575 179.045 ;
        RECT 115.405 178.875 115.575 179.045 ;
        RECT 116.405 178.875 116.575 179.045 ;
        RECT 117.405 178.875 117.575 179.045 ;
        RECT 118.405 178.875 118.575 179.045 ;
        RECT 119.405 178.875 119.575 179.045 ;
        RECT 120.405 178.875 120.575 179.045 ;
        RECT 121.405 178.875 121.575 179.045 ;
        RECT 122.405 178.875 122.575 179.045 ;
        RECT 123.405 178.875 123.575 179.045 ;
        RECT 128.005 178.875 128.175 179.045 ;
        RECT 130.005 178.875 130.175 179.045 ;
        RECT 132.005 178.875 132.175 179.045 ;
        RECT 134.005 178.875 134.175 179.045 ;
        RECT 136.005 178.875 136.175 179.045 ;
        RECT 138.005 178.875 138.175 179.045 ;
        RECT 140.005 178.875 140.175 179.045 ;
        RECT 142.005 178.875 142.175 179.045 ;
        RECT 144.005 178.875 144.175 179.045 ;
        RECT 146.005 178.875 146.175 179.045 ;
        RECT 150.555 178.875 150.725 179.045 ;
        RECT 152.555 178.875 152.725 179.045 ;
        RECT 154.555 178.875 154.725 179.045 ;
        RECT 156.555 178.875 156.725 179.045 ;
        RECT 158.555 178.875 158.725 179.045 ;
        RECT 160.555 178.875 160.725 179.045 ;
        RECT 162.555 178.875 162.725 179.045 ;
        RECT 164.555 178.875 164.725 179.045 ;
        RECT 166.555 178.875 166.725 179.045 ;
        RECT 168.555 178.875 168.725 179.045 ;
        RECT 170.555 178.875 170.725 179.045 ;
        RECT 172.555 178.875 172.725 179.045 ;
        RECT 174.555 178.875 174.725 179.045 ;
        RECT 176.555 178.875 176.725 179.045 ;
        RECT 178.555 178.875 178.725 179.045 ;
        RECT 180.555 178.875 180.725 179.045 ;
        RECT 182.555 178.875 182.725 179.045 ;
        RECT 184.555 178.875 184.725 179.045 ;
        RECT 188.275 178.875 188.445 179.045 ;
        RECT 190.275 178.875 190.445 179.045 ;
        RECT 192.275 178.875 192.445 179.045 ;
        RECT 194.275 178.875 194.445 179.045 ;
        RECT 196.275 178.875 196.445 179.045 ;
        RECT 198.275 178.875 198.445 179.045 ;
        RECT 200.275 178.875 200.445 179.045 ;
        RECT 209.835 178.875 210.005 179.045 ;
        RECT 210.835 178.875 211.005 179.045 ;
        RECT 211.835 178.875 212.005 179.045 ;
        RECT 212.835 178.875 213.005 179.045 ;
        RECT 213.835 178.875 214.005 179.045 ;
        RECT 214.835 178.875 215.005 179.045 ;
        RECT 215.835 178.875 216.005 179.045 ;
        RECT 216.835 178.875 217.005 179.045 ;
        RECT 217.835 178.875 218.005 179.045 ;
        RECT 218.835 178.875 219.005 179.045 ;
        RECT 219.835 178.875 220.005 179.045 ;
        RECT 220.835 178.875 221.005 179.045 ;
        RECT 221.835 178.875 222.005 179.045 ;
        RECT 222.835 178.875 223.005 179.045 ;
        RECT 223.835 178.875 224.005 179.045 ;
        RECT 224.835 178.875 225.005 179.045 ;
        RECT 225.835 178.875 226.005 179.045 ;
        RECT 226.835 178.875 227.005 179.045 ;
        RECT 227.835 178.875 228.005 179.045 ;
        RECT 228.835 178.875 229.005 179.045 ;
        RECT 229.835 178.875 230.005 179.045 ;
        RECT 230.835 178.875 231.005 179.045 ;
        RECT 231.835 178.875 232.005 179.045 ;
        RECT 232.835 178.875 233.005 179.045 ;
        RECT 233.835 178.875 234.005 179.045 ;
        RECT 234.835 178.875 235.005 179.045 ;
        RECT 235.835 178.875 236.005 179.045 ;
        RECT 236.835 178.875 237.005 179.045 ;
        RECT 237.835 178.875 238.005 179.045 ;
        RECT 238.835 178.875 239.005 179.045 ;
        RECT 239.835 178.875 240.005 179.045 ;
        RECT 240.835 178.875 241.005 179.045 ;
        RECT 241.835 178.875 242.005 179.045 ;
        RECT 242.835 178.875 243.005 179.045 ;
        RECT 243.835 178.875 244.005 179.045 ;
        RECT 244.835 178.875 245.005 179.045 ;
        RECT 245.835 178.875 246.005 179.045 ;
        RECT 246.835 178.875 247.005 179.045 ;
        RECT 247.835 178.875 248.005 179.045 ;
        RECT 248.835 178.875 249.005 179.045 ;
        RECT 249.835 178.875 250.005 179.045 ;
        RECT 250.835 178.875 251.005 179.045 ;
        RECT 251.835 178.875 252.005 179.045 ;
        RECT 252.835 178.875 253.005 179.045 ;
        RECT 253.835 178.875 254.005 179.045 ;
        RECT 254.835 178.875 255.005 179.045 ;
        RECT 255.835 178.875 256.005 179.045 ;
        RECT 256.835 178.875 257.005 179.045 ;
        RECT 257.835 178.875 258.005 179.045 ;
        RECT 258.835 178.875 259.005 179.045 ;
        RECT 259.835 178.875 260.005 179.045 ;
        RECT 260.835 178.875 261.005 179.045 ;
        RECT 261.835 178.875 262.005 179.045 ;
        RECT 209.150 167.810 209.320 167.980 ;
        RECT 209.600 167.810 209.770 167.980 ;
        RECT 210.050 167.810 210.220 167.980 ;
        RECT 210.500 167.810 210.670 167.980 ;
        RECT 210.950 167.810 211.120 167.980 ;
        RECT 211.400 167.810 211.570 167.980 ;
        RECT 211.850 167.810 212.020 167.980 ;
        RECT 212.300 167.810 212.470 167.980 ;
        RECT 212.750 167.810 212.920 167.980 ;
        RECT 213.200 167.810 213.370 167.980 ;
        RECT 213.650 167.810 213.820 167.980 ;
        RECT 214.100 167.810 214.270 167.980 ;
        RECT 214.550 167.810 214.720 167.980 ;
        RECT 215.000 167.810 215.170 167.980 ;
        RECT 215.850 167.810 216.020 167.980 ;
        RECT 216.300 167.810 216.470 167.980 ;
        RECT 216.750 167.810 216.920 167.980 ;
        RECT 217.200 167.810 217.370 167.980 ;
        RECT 217.650 167.810 217.820 167.980 ;
        RECT 218.100 167.810 218.270 167.980 ;
        RECT 218.550 167.810 218.720 167.980 ;
        RECT 219.000 167.810 219.170 167.980 ;
        RECT 219.450 167.810 219.620 167.980 ;
        RECT 219.900 167.810 220.070 167.980 ;
        RECT 220.350 167.810 220.520 167.980 ;
        RECT 220.800 167.810 220.970 167.980 ;
        RECT 221.250 167.810 221.420 167.980 ;
        RECT 221.700 167.810 221.870 167.980 ;
        RECT 222.550 167.810 222.720 167.980 ;
        RECT 223.000 167.810 223.170 167.980 ;
        RECT 223.450 167.810 223.620 167.980 ;
        RECT 223.900 167.810 224.070 167.980 ;
        RECT 224.350 167.810 224.520 167.980 ;
        RECT 224.800 167.810 224.970 167.980 ;
        RECT 225.250 167.810 225.420 167.980 ;
        RECT 225.700 167.810 225.870 167.980 ;
        RECT 226.150 167.810 226.320 167.980 ;
        RECT 226.600 167.810 226.770 167.980 ;
        RECT 227.050 167.810 227.220 167.980 ;
        RECT 227.500 167.810 227.670 167.980 ;
        RECT 227.950 167.810 228.120 167.980 ;
        RECT 228.400 167.810 228.570 167.980 ;
        RECT 229.250 167.810 229.420 167.980 ;
        RECT 229.700 167.810 229.870 167.980 ;
        RECT 230.150 167.810 230.320 167.980 ;
        RECT 230.600 167.810 230.770 167.980 ;
        RECT 231.050 167.810 231.220 167.980 ;
        RECT 231.500 167.810 231.670 167.980 ;
        RECT 231.950 167.810 232.120 167.980 ;
        RECT 232.400 167.810 232.570 167.980 ;
        RECT 232.850 167.810 233.020 167.980 ;
        RECT 233.300 167.810 233.470 167.980 ;
        RECT 233.750 167.810 233.920 167.980 ;
        RECT 234.200 167.810 234.370 167.980 ;
        RECT 234.650 167.810 234.820 167.980 ;
        RECT 235.100 167.810 235.270 167.980 ;
        RECT 235.950 167.810 236.120 167.980 ;
        RECT 236.400 167.810 236.570 167.980 ;
        RECT 236.850 167.810 237.020 167.980 ;
        RECT 237.300 167.810 237.470 167.980 ;
        RECT 237.750 167.810 237.920 167.980 ;
        RECT 238.200 167.810 238.370 167.980 ;
        RECT 238.650 167.810 238.820 167.980 ;
        RECT 239.100 167.810 239.270 167.980 ;
        RECT 239.550 167.810 239.720 167.980 ;
        RECT 240.000 167.810 240.170 167.980 ;
        RECT 240.450 167.810 240.620 167.980 ;
        RECT 240.900 167.810 241.070 167.980 ;
        RECT 241.350 167.810 241.520 167.980 ;
        RECT 241.800 167.810 241.970 167.980 ;
        RECT 242.650 167.810 242.820 167.980 ;
        RECT 243.100 167.810 243.270 167.980 ;
        RECT 243.550 167.810 243.720 167.980 ;
        RECT 244.000 167.810 244.170 167.980 ;
        RECT 244.450 167.810 244.620 167.980 ;
        RECT 244.900 167.810 245.070 167.980 ;
        RECT 245.350 167.810 245.520 167.980 ;
        RECT 245.800 167.810 245.970 167.980 ;
        RECT 246.250 167.810 246.420 167.980 ;
        RECT 246.700 167.810 246.870 167.980 ;
        RECT 247.150 167.810 247.320 167.980 ;
        RECT 247.600 167.810 247.770 167.980 ;
        RECT 248.050 167.810 248.220 167.980 ;
        RECT 248.500 167.810 248.670 167.980 ;
        RECT 249.350 167.810 249.520 167.980 ;
        RECT 249.800 167.810 249.970 167.980 ;
        RECT 250.250 167.810 250.420 167.980 ;
        RECT 250.700 167.810 250.870 167.980 ;
        RECT 251.150 167.810 251.320 167.980 ;
        RECT 251.600 167.810 251.770 167.980 ;
        RECT 252.050 167.810 252.220 167.980 ;
        RECT 252.500 167.810 252.670 167.980 ;
        RECT 252.950 167.810 253.120 167.980 ;
        RECT 253.400 167.810 253.570 167.980 ;
        RECT 253.850 167.810 254.020 167.980 ;
        RECT 254.300 167.810 254.470 167.980 ;
        RECT 254.750 167.810 254.920 167.980 ;
        RECT 255.200 167.810 255.370 167.980 ;
        RECT 256.050 167.810 256.220 167.980 ;
        RECT 256.500 167.810 256.670 167.980 ;
        RECT 256.950 167.810 257.120 167.980 ;
        RECT 257.400 167.810 257.570 167.980 ;
        RECT 257.850 167.810 258.020 167.980 ;
        RECT 258.300 167.810 258.470 167.980 ;
        RECT 258.750 167.810 258.920 167.980 ;
        RECT 259.200 167.810 259.370 167.980 ;
        RECT 259.650 167.810 259.820 167.980 ;
        RECT 260.100 167.810 260.270 167.980 ;
        RECT 260.550 167.810 260.720 167.980 ;
        RECT 261.000 167.810 261.170 167.980 ;
        RECT 261.450 167.810 261.620 167.980 ;
        RECT 261.900 167.810 262.070 167.980 ;
        RECT 110.140 160.815 112.110 163.505 ;
        RECT 209.970 167.010 210.140 167.180 ;
        RECT 210.420 167.010 210.590 167.180 ;
        RECT 210.870 167.010 211.040 167.180 ;
        RECT 211.320 167.010 211.490 167.180 ;
        RECT 211.770 167.010 211.940 167.180 ;
        RECT 212.220 167.010 212.390 167.180 ;
        RECT 212.670 167.010 212.840 167.180 ;
        RECT 213.120 167.010 213.290 167.180 ;
        RECT 213.570 167.010 213.740 167.180 ;
        RECT 214.020 167.010 214.190 167.180 ;
        RECT 214.470 167.010 214.640 167.180 ;
        RECT 216.670 167.010 216.840 167.180 ;
        RECT 217.120 167.010 217.290 167.180 ;
        RECT 217.570 167.010 217.740 167.180 ;
        RECT 218.020 167.010 218.190 167.180 ;
        RECT 218.470 167.010 218.640 167.180 ;
        RECT 218.920 167.010 219.090 167.180 ;
        RECT 219.370 167.010 219.540 167.180 ;
        RECT 219.820 167.010 219.990 167.180 ;
        RECT 220.270 167.010 220.440 167.180 ;
        RECT 220.720 167.010 220.890 167.180 ;
        RECT 221.170 167.010 221.340 167.180 ;
        RECT 223.370 167.010 223.540 167.180 ;
        RECT 223.820 167.010 223.990 167.180 ;
        RECT 224.270 167.010 224.440 167.180 ;
        RECT 224.720 167.010 224.890 167.180 ;
        RECT 225.170 167.010 225.340 167.180 ;
        RECT 225.620 167.010 225.790 167.180 ;
        RECT 226.070 167.010 226.240 167.180 ;
        RECT 226.520 167.010 226.690 167.180 ;
        RECT 226.970 167.010 227.140 167.180 ;
        RECT 227.420 167.010 227.590 167.180 ;
        RECT 227.870 167.010 228.040 167.180 ;
        RECT 230.070 167.010 230.240 167.180 ;
        RECT 230.520 167.010 230.690 167.180 ;
        RECT 230.970 167.010 231.140 167.180 ;
        RECT 231.420 167.010 231.590 167.180 ;
        RECT 231.870 167.010 232.040 167.180 ;
        RECT 232.320 167.010 232.490 167.180 ;
        RECT 232.770 167.010 232.940 167.180 ;
        RECT 233.220 167.010 233.390 167.180 ;
        RECT 233.670 167.010 233.840 167.180 ;
        RECT 234.120 167.010 234.290 167.180 ;
        RECT 234.570 167.010 234.740 167.180 ;
        RECT 236.770 167.010 236.940 167.180 ;
        RECT 237.220 167.010 237.390 167.180 ;
        RECT 237.670 167.010 237.840 167.180 ;
        RECT 238.120 167.010 238.290 167.180 ;
        RECT 238.570 167.010 238.740 167.180 ;
        RECT 239.020 167.010 239.190 167.180 ;
        RECT 239.470 167.010 239.640 167.180 ;
        RECT 239.920 167.010 240.090 167.180 ;
        RECT 240.370 167.010 240.540 167.180 ;
        RECT 240.820 167.010 240.990 167.180 ;
        RECT 241.270 167.010 241.440 167.180 ;
        RECT 243.470 167.010 243.640 167.180 ;
        RECT 243.920 167.010 244.090 167.180 ;
        RECT 244.370 167.010 244.540 167.180 ;
        RECT 244.820 167.010 244.990 167.180 ;
        RECT 245.270 167.010 245.440 167.180 ;
        RECT 245.720 167.010 245.890 167.180 ;
        RECT 246.170 167.010 246.340 167.180 ;
        RECT 246.620 167.010 246.790 167.180 ;
        RECT 247.070 167.010 247.240 167.180 ;
        RECT 247.520 167.010 247.690 167.180 ;
        RECT 247.970 167.010 248.140 167.180 ;
        RECT 250.170 167.010 250.340 167.180 ;
        RECT 250.620 167.010 250.790 167.180 ;
        RECT 251.070 167.010 251.240 167.180 ;
        RECT 251.520 167.010 251.690 167.180 ;
        RECT 251.970 167.010 252.140 167.180 ;
        RECT 252.420 167.010 252.590 167.180 ;
        RECT 252.870 167.010 253.040 167.180 ;
        RECT 253.320 167.010 253.490 167.180 ;
        RECT 253.770 167.010 253.940 167.180 ;
        RECT 254.220 167.010 254.390 167.180 ;
        RECT 254.670 167.010 254.840 167.180 ;
        RECT 256.870 167.010 257.040 167.180 ;
        RECT 257.320 167.010 257.490 167.180 ;
        RECT 257.770 167.010 257.940 167.180 ;
        RECT 258.220 167.010 258.390 167.180 ;
        RECT 258.670 167.010 258.840 167.180 ;
        RECT 259.120 167.010 259.290 167.180 ;
        RECT 259.570 167.010 259.740 167.180 ;
        RECT 260.020 167.010 260.190 167.180 ;
        RECT 260.470 167.010 260.640 167.180 ;
        RECT 260.920 167.010 261.090 167.180 ;
        RECT 261.370 167.010 261.540 167.180 ;
        RECT 97.235 160.075 97.405 160.245 ;
        RECT 98.235 160.075 98.405 160.245 ;
        RECT 99.235 160.075 99.405 160.245 ;
        RECT 100.235 160.075 100.405 160.245 ;
        RECT 101.235 160.075 101.405 160.245 ;
        RECT 102.235 160.075 102.405 160.245 ;
        RECT 103.235 160.075 103.405 160.245 ;
        RECT 104.235 160.075 104.405 160.245 ;
        RECT 105.235 160.075 105.405 160.245 ;
        RECT 106.235 160.075 106.405 160.245 ;
        RECT 107.235 160.075 107.405 160.245 ;
        RECT 110.965 160.075 111.135 160.245 ;
        RECT 111.965 160.075 112.135 160.245 ;
        RECT 112.965 160.075 113.135 160.245 ;
        RECT 113.965 160.075 114.135 160.245 ;
        RECT 114.965 160.075 115.135 160.245 ;
        RECT 115.965 160.075 116.135 160.245 ;
        RECT 116.965 160.075 117.135 160.245 ;
        RECT 117.965 160.075 118.135 160.245 ;
        RECT 118.965 160.075 119.135 160.245 ;
        RECT 119.965 160.075 120.135 160.245 ;
        RECT 120.965 160.075 121.135 160.245 ;
        RECT 121.965 160.075 122.135 160.245 ;
        RECT 122.965 160.075 123.135 160.245 ;
        RECT 123.965 160.075 124.135 160.245 ;
        RECT 131.935 160.075 132.105 160.245 ;
        RECT 133.935 160.075 134.105 160.245 ;
        RECT 135.935 160.075 136.105 160.245 ;
        RECT 137.935 160.075 138.105 160.245 ;
        RECT 139.935 160.075 140.105 160.245 ;
        RECT 141.935 160.075 142.105 160.245 ;
        RECT 143.935 160.075 144.105 160.245 ;
        RECT 145.935 160.075 146.105 160.245 ;
        RECT 147.935 160.075 148.105 160.245 ;
        RECT 149.935 160.075 150.105 160.245 ;
        RECT 151.935 160.075 152.105 160.245 ;
        RECT 153.935 160.075 154.105 160.245 ;
        RECT 155.935 160.075 156.105 160.245 ;
        RECT 157.935 160.075 158.105 160.245 ;
        RECT 159.935 160.075 160.105 160.245 ;
        RECT 161.935 160.075 162.105 160.245 ;
        RECT 163.935 160.075 164.105 160.245 ;
        RECT 165.935 160.075 166.105 160.245 ;
        RECT 169.175 160.075 169.345 160.245 ;
        RECT 171.175 160.075 171.345 160.245 ;
        RECT 173.175 160.075 173.345 160.245 ;
        RECT 175.175 160.075 175.345 160.245 ;
        RECT 177.175 160.075 177.345 160.245 ;
        RECT 179.175 160.075 179.345 160.245 ;
        RECT 181.175 160.075 181.345 160.245 ;
        RECT 183.175 160.075 183.345 160.245 ;
        RECT 185.175 160.075 185.345 160.245 ;
        RECT 187.175 160.075 187.345 160.245 ;
        RECT 189.175 160.075 189.345 160.245 ;
        RECT 191.175 160.075 191.345 160.245 ;
        RECT 193.175 160.075 193.345 160.245 ;
        RECT 195.175 160.075 195.345 160.245 ;
        RECT 197.175 160.075 197.345 160.245 ;
        RECT 199.175 160.075 199.345 160.245 ;
        RECT 201.175 160.075 201.345 160.245 ;
        RECT 203.175 160.075 203.345 160.245 ;
        RECT 209.835 160.075 210.005 160.245 ;
        RECT 210.835 160.075 211.005 160.245 ;
        RECT 211.835 160.075 212.005 160.245 ;
        RECT 212.835 160.075 213.005 160.245 ;
        RECT 213.835 160.075 214.005 160.245 ;
        RECT 214.835 160.075 215.005 160.245 ;
        RECT 215.835 160.075 216.005 160.245 ;
        RECT 216.835 160.075 217.005 160.245 ;
        RECT 217.835 160.075 218.005 160.245 ;
        RECT 218.835 160.075 219.005 160.245 ;
        RECT 219.835 160.075 220.005 160.245 ;
        RECT 220.835 160.075 221.005 160.245 ;
        RECT 221.835 160.075 222.005 160.245 ;
        RECT 222.835 160.075 223.005 160.245 ;
        RECT 223.835 160.075 224.005 160.245 ;
        RECT 224.835 160.075 225.005 160.245 ;
        RECT 225.835 160.075 226.005 160.245 ;
        RECT 226.835 160.075 227.005 160.245 ;
        RECT 227.835 160.075 228.005 160.245 ;
        RECT 228.835 160.075 229.005 160.245 ;
        RECT 229.835 160.075 230.005 160.245 ;
        RECT 230.835 160.075 231.005 160.245 ;
        RECT 231.835 160.075 232.005 160.245 ;
        RECT 232.835 160.075 233.005 160.245 ;
        RECT 233.835 160.075 234.005 160.245 ;
        RECT 234.835 160.075 235.005 160.245 ;
        RECT 235.835 160.075 236.005 160.245 ;
        RECT 236.835 160.075 237.005 160.245 ;
        RECT 237.835 160.075 238.005 160.245 ;
        RECT 238.835 160.075 239.005 160.245 ;
        RECT 239.835 160.075 240.005 160.245 ;
        RECT 240.835 160.075 241.005 160.245 ;
        RECT 241.835 160.075 242.005 160.245 ;
        RECT 242.835 160.075 243.005 160.245 ;
        RECT 243.835 160.075 244.005 160.245 ;
        RECT 244.835 160.075 245.005 160.245 ;
        RECT 245.835 160.075 246.005 160.245 ;
        RECT 246.835 160.075 247.005 160.245 ;
        RECT 247.835 160.075 248.005 160.245 ;
        RECT 248.835 160.075 249.005 160.245 ;
        RECT 249.835 160.075 250.005 160.245 ;
        RECT 250.835 160.075 251.005 160.245 ;
        RECT 251.835 160.075 252.005 160.245 ;
        RECT 252.835 160.075 253.005 160.245 ;
        RECT 253.835 160.075 254.005 160.245 ;
        RECT 254.835 160.075 255.005 160.245 ;
        RECT 255.835 160.075 256.005 160.245 ;
        RECT 256.835 160.075 257.005 160.245 ;
        RECT 257.835 160.075 258.005 160.245 ;
        RECT 258.835 160.075 259.005 160.245 ;
        RECT 259.835 160.075 260.005 160.245 ;
        RECT 260.835 160.075 261.005 160.245 ;
        RECT 261.835 160.075 262.005 160.245 ;
        RECT 209.150 149.010 209.320 149.180 ;
        RECT 209.600 149.010 209.770 149.180 ;
        RECT 210.050 149.010 210.220 149.180 ;
        RECT 210.500 149.010 210.670 149.180 ;
        RECT 210.950 149.010 211.120 149.180 ;
        RECT 211.400 149.010 211.570 149.180 ;
        RECT 211.850 149.010 212.020 149.180 ;
        RECT 212.300 149.010 212.470 149.180 ;
        RECT 212.750 149.010 212.920 149.180 ;
        RECT 213.200 149.010 213.370 149.180 ;
        RECT 213.650 149.010 213.820 149.180 ;
        RECT 214.100 149.010 214.270 149.180 ;
        RECT 214.550 149.010 214.720 149.180 ;
        RECT 215.000 149.010 215.170 149.180 ;
        RECT 215.850 149.010 216.020 149.180 ;
        RECT 216.300 149.010 216.470 149.180 ;
        RECT 216.750 149.010 216.920 149.180 ;
        RECT 217.200 149.010 217.370 149.180 ;
        RECT 217.650 149.010 217.820 149.180 ;
        RECT 218.100 149.010 218.270 149.180 ;
        RECT 218.550 149.010 218.720 149.180 ;
        RECT 219.000 149.010 219.170 149.180 ;
        RECT 219.450 149.010 219.620 149.180 ;
        RECT 219.900 149.010 220.070 149.180 ;
        RECT 220.350 149.010 220.520 149.180 ;
        RECT 220.800 149.010 220.970 149.180 ;
        RECT 221.250 149.010 221.420 149.180 ;
        RECT 221.700 149.010 221.870 149.180 ;
        RECT 222.550 149.010 222.720 149.180 ;
        RECT 223.000 149.010 223.170 149.180 ;
        RECT 223.450 149.010 223.620 149.180 ;
        RECT 223.900 149.010 224.070 149.180 ;
        RECT 224.350 149.010 224.520 149.180 ;
        RECT 224.800 149.010 224.970 149.180 ;
        RECT 225.250 149.010 225.420 149.180 ;
        RECT 225.700 149.010 225.870 149.180 ;
        RECT 226.150 149.010 226.320 149.180 ;
        RECT 226.600 149.010 226.770 149.180 ;
        RECT 227.050 149.010 227.220 149.180 ;
        RECT 227.500 149.010 227.670 149.180 ;
        RECT 227.950 149.010 228.120 149.180 ;
        RECT 228.400 149.010 228.570 149.180 ;
        RECT 229.250 149.010 229.420 149.180 ;
        RECT 229.700 149.010 229.870 149.180 ;
        RECT 230.150 149.010 230.320 149.180 ;
        RECT 230.600 149.010 230.770 149.180 ;
        RECT 231.050 149.010 231.220 149.180 ;
        RECT 231.500 149.010 231.670 149.180 ;
        RECT 231.950 149.010 232.120 149.180 ;
        RECT 232.400 149.010 232.570 149.180 ;
        RECT 232.850 149.010 233.020 149.180 ;
        RECT 233.300 149.010 233.470 149.180 ;
        RECT 233.750 149.010 233.920 149.180 ;
        RECT 234.200 149.010 234.370 149.180 ;
        RECT 234.650 149.010 234.820 149.180 ;
        RECT 235.100 149.010 235.270 149.180 ;
        RECT 235.950 149.010 236.120 149.180 ;
        RECT 236.400 149.010 236.570 149.180 ;
        RECT 236.850 149.010 237.020 149.180 ;
        RECT 237.300 149.010 237.470 149.180 ;
        RECT 237.750 149.010 237.920 149.180 ;
        RECT 238.200 149.010 238.370 149.180 ;
        RECT 238.650 149.010 238.820 149.180 ;
        RECT 239.100 149.010 239.270 149.180 ;
        RECT 239.550 149.010 239.720 149.180 ;
        RECT 240.000 149.010 240.170 149.180 ;
        RECT 240.450 149.010 240.620 149.180 ;
        RECT 240.900 149.010 241.070 149.180 ;
        RECT 241.350 149.010 241.520 149.180 ;
        RECT 241.800 149.010 241.970 149.180 ;
        RECT 242.650 149.010 242.820 149.180 ;
        RECT 243.100 149.010 243.270 149.180 ;
        RECT 243.550 149.010 243.720 149.180 ;
        RECT 244.000 149.010 244.170 149.180 ;
        RECT 244.450 149.010 244.620 149.180 ;
        RECT 244.900 149.010 245.070 149.180 ;
        RECT 245.350 149.010 245.520 149.180 ;
        RECT 245.800 149.010 245.970 149.180 ;
        RECT 246.250 149.010 246.420 149.180 ;
        RECT 246.700 149.010 246.870 149.180 ;
        RECT 247.150 149.010 247.320 149.180 ;
        RECT 247.600 149.010 247.770 149.180 ;
        RECT 248.050 149.010 248.220 149.180 ;
        RECT 248.500 149.010 248.670 149.180 ;
        RECT 249.350 149.010 249.520 149.180 ;
        RECT 249.800 149.010 249.970 149.180 ;
        RECT 250.250 149.010 250.420 149.180 ;
        RECT 250.700 149.010 250.870 149.180 ;
        RECT 251.150 149.010 251.320 149.180 ;
        RECT 251.600 149.010 251.770 149.180 ;
        RECT 252.050 149.010 252.220 149.180 ;
        RECT 252.500 149.010 252.670 149.180 ;
        RECT 252.950 149.010 253.120 149.180 ;
        RECT 253.400 149.010 253.570 149.180 ;
        RECT 253.850 149.010 254.020 149.180 ;
        RECT 254.300 149.010 254.470 149.180 ;
        RECT 254.750 149.010 254.920 149.180 ;
        RECT 255.200 149.010 255.370 149.180 ;
        RECT 256.050 149.010 256.220 149.180 ;
        RECT 256.500 149.010 256.670 149.180 ;
        RECT 256.950 149.010 257.120 149.180 ;
        RECT 257.400 149.010 257.570 149.180 ;
        RECT 257.850 149.010 258.020 149.180 ;
        RECT 258.300 149.010 258.470 149.180 ;
        RECT 258.750 149.010 258.920 149.180 ;
        RECT 259.200 149.010 259.370 149.180 ;
        RECT 259.650 149.010 259.820 149.180 ;
        RECT 260.100 149.010 260.270 149.180 ;
        RECT 260.550 149.010 260.720 149.180 ;
        RECT 261.000 149.010 261.170 149.180 ;
        RECT 261.450 149.010 261.620 149.180 ;
        RECT 261.900 149.010 262.070 149.180 ;
        RECT 209.970 148.210 210.140 148.380 ;
        RECT 210.420 148.210 210.590 148.380 ;
        RECT 210.870 148.210 211.040 148.380 ;
        RECT 211.320 148.210 211.490 148.380 ;
        RECT 211.770 148.210 211.940 148.380 ;
        RECT 212.220 148.210 212.390 148.380 ;
        RECT 212.670 148.210 212.840 148.380 ;
        RECT 213.120 148.210 213.290 148.380 ;
        RECT 213.570 148.210 213.740 148.380 ;
        RECT 214.020 148.210 214.190 148.380 ;
        RECT 214.470 148.210 214.640 148.380 ;
        RECT 216.670 148.210 216.840 148.380 ;
        RECT 217.120 148.210 217.290 148.380 ;
        RECT 217.570 148.210 217.740 148.380 ;
        RECT 218.020 148.210 218.190 148.380 ;
        RECT 218.470 148.210 218.640 148.380 ;
        RECT 218.920 148.210 219.090 148.380 ;
        RECT 219.370 148.210 219.540 148.380 ;
        RECT 219.820 148.210 219.990 148.380 ;
        RECT 220.270 148.210 220.440 148.380 ;
        RECT 220.720 148.210 220.890 148.380 ;
        RECT 221.170 148.210 221.340 148.380 ;
        RECT 223.370 148.210 223.540 148.380 ;
        RECT 223.820 148.210 223.990 148.380 ;
        RECT 224.270 148.210 224.440 148.380 ;
        RECT 224.720 148.210 224.890 148.380 ;
        RECT 225.170 148.210 225.340 148.380 ;
        RECT 225.620 148.210 225.790 148.380 ;
        RECT 226.070 148.210 226.240 148.380 ;
        RECT 226.520 148.210 226.690 148.380 ;
        RECT 226.970 148.210 227.140 148.380 ;
        RECT 227.420 148.210 227.590 148.380 ;
        RECT 227.870 148.210 228.040 148.380 ;
        RECT 230.070 148.210 230.240 148.380 ;
        RECT 230.520 148.210 230.690 148.380 ;
        RECT 230.970 148.210 231.140 148.380 ;
        RECT 231.420 148.210 231.590 148.380 ;
        RECT 231.870 148.210 232.040 148.380 ;
        RECT 232.320 148.210 232.490 148.380 ;
        RECT 232.770 148.210 232.940 148.380 ;
        RECT 233.220 148.210 233.390 148.380 ;
        RECT 233.670 148.210 233.840 148.380 ;
        RECT 234.120 148.210 234.290 148.380 ;
        RECT 234.570 148.210 234.740 148.380 ;
        RECT 236.770 148.210 236.940 148.380 ;
        RECT 237.220 148.210 237.390 148.380 ;
        RECT 237.670 148.210 237.840 148.380 ;
        RECT 238.120 148.210 238.290 148.380 ;
        RECT 238.570 148.210 238.740 148.380 ;
        RECT 239.020 148.210 239.190 148.380 ;
        RECT 239.470 148.210 239.640 148.380 ;
        RECT 239.920 148.210 240.090 148.380 ;
        RECT 240.370 148.210 240.540 148.380 ;
        RECT 240.820 148.210 240.990 148.380 ;
        RECT 241.270 148.210 241.440 148.380 ;
        RECT 243.470 148.210 243.640 148.380 ;
        RECT 243.920 148.210 244.090 148.380 ;
        RECT 244.370 148.210 244.540 148.380 ;
        RECT 244.820 148.210 244.990 148.380 ;
        RECT 245.270 148.210 245.440 148.380 ;
        RECT 245.720 148.210 245.890 148.380 ;
        RECT 246.170 148.210 246.340 148.380 ;
        RECT 246.620 148.210 246.790 148.380 ;
        RECT 247.070 148.210 247.240 148.380 ;
        RECT 247.520 148.210 247.690 148.380 ;
        RECT 247.970 148.210 248.140 148.380 ;
        RECT 250.170 148.210 250.340 148.380 ;
        RECT 250.620 148.210 250.790 148.380 ;
        RECT 251.070 148.210 251.240 148.380 ;
        RECT 251.520 148.210 251.690 148.380 ;
        RECT 251.970 148.210 252.140 148.380 ;
        RECT 252.420 148.210 252.590 148.380 ;
        RECT 252.870 148.210 253.040 148.380 ;
        RECT 253.320 148.210 253.490 148.380 ;
        RECT 253.770 148.210 253.940 148.380 ;
        RECT 254.220 148.210 254.390 148.380 ;
        RECT 254.670 148.210 254.840 148.380 ;
        RECT 256.870 148.210 257.040 148.380 ;
        RECT 257.320 148.210 257.490 148.380 ;
        RECT 257.770 148.210 257.940 148.380 ;
        RECT 258.220 148.210 258.390 148.380 ;
        RECT 258.670 148.210 258.840 148.380 ;
        RECT 259.120 148.210 259.290 148.380 ;
        RECT 259.570 148.210 259.740 148.380 ;
        RECT 260.020 148.210 260.190 148.380 ;
        RECT 260.470 148.210 260.640 148.380 ;
        RECT 260.920 148.210 261.090 148.380 ;
        RECT 261.370 148.210 261.540 148.380 ;
        RECT 83.515 141.275 83.685 141.445 ;
        RECT 84.515 141.275 84.685 141.445 ;
        RECT 85.515 141.275 85.685 141.445 ;
        RECT 86.515 141.275 86.685 141.445 ;
        RECT 87.515 141.275 87.685 141.445 ;
        RECT 88.515 141.275 88.685 141.445 ;
        RECT 89.515 141.275 89.685 141.445 ;
        RECT 90.515 141.275 90.685 141.445 ;
        RECT 91.515 141.275 91.685 141.445 ;
        RECT 92.515 141.275 92.685 141.445 ;
        RECT 93.515 141.275 93.685 141.445 ;
        RECT 97.235 141.275 97.405 141.445 ;
        RECT 98.235 141.275 98.405 141.445 ;
        RECT 99.235 141.275 99.405 141.445 ;
        RECT 100.235 141.275 100.405 141.445 ;
        RECT 101.235 141.275 101.405 141.445 ;
        RECT 102.235 141.275 102.405 141.445 ;
        RECT 103.235 141.275 103.405 141.445 ;
        RECT 104.235 141.275 104.405 141.445 ;
        RECT 105.235 141.275 105.405 141.445 ;
        RECT 106.235 141.275 106.405 141.445 ;
        RECT 107.235 141.275 107.405 141.445 ;
        RECT 110.955 141.275 111.125 141.445 ;
        RECT 111.955 141.275 112.125 141.445 ;
        RECT 112.955 141.275 113.125 141.445 ;
        RECT 113.955 141.275 114.125 141.445 ;
        RECT 114.955 141.275 115.125 141.445 ;
        RECT 115.955 141.275 116.125 141.445 ;
        RECT 116.955 141.275 117.125 141.445 ;
        RECT 117.955 141.275 118.125 141.445 ;
        RECT 118.955 141.275 119.125 141.445 ;
        RECT 119.955 141.275 120.125 141.445 ;
        RECT 120.955 141.275 121.125 141.445 ;
        RECT 136.925 141.275 137.095 141.445 ;
        RECT 137.925 141.275 138.095 141.445 ;
        RECT 138.925 141.275 139.095 141.445 ;
        RECT 139.925 141.275 140.095 141.445 ;
        RECT 140.925 141.275 141.095 141.445 ;
        RECT 141.925 141.275 142.095 141.445 ;
        RECT 142.925 141.275 143.095 141.445 ;
        RECT 143.925 141.275 144.095 141.445 ;
        RECT 144.925 141.275 145.095 141.445 ;
        RECT 145.925 141.275 146.095 141.445 ;
        RECT 146.925 141.275 147.095 141.445 ;
        RECT 150.555 141.275 150.725 141.445 ;
        RECT 152.555 141.275 152.725 141.445 ;
        RECT 154.555 141.275 154.725 141.445 ;
        RECT 156.555 141.275 156.725 141.445 ;
        RECT 158.555 141.275 158.725 141.445 ;
        RECT 160.555 141.275 160.725 141.445 ;
        RECT 162.555 141.275 162.725 141.445 ;
        RECT 164.555 141.275 164.725 141.445 ;
        RECT 166.555 141.275 166.725 141.445 ;
        RECT 168.555 141.275 168.725 141.445 ;
        RECT 170.555 141.275 170.725 141.445 ;
        RECT 172.555 141.275 172.725 141.445 ;
        RECT 174.555 141.275 174.725 141.445 ;
        RECT 176.555 141.275 176.725 141.445 ;
        RECT 178.555 141.275 178.725 141.445 ;
        RECT 180.555 141.275 180.725 141.445 ;
        RECT 182.555 141.275 182.725 141.445 ;
        RECT 184.555 141.275 184.725 141.445 ;
        RECT 188.275 141.275 188.445 141.445 ;
        RECT 190.275 141.275 190.445 141.445 ;
        RECT 192.275 141.275 192.445 141.445 ;
        RECT 194.275 141.275 194.445 141.445 ;
        RECT 196.275 141.275 196.445 141.445 ;
        RECT 198.275 141.275 198.445 141.445 ;
        RECT 200.275 141.275 200.445 141.445 ;
        RECT 209.835 141.275 210.005 141.445 ;
        RECT 210.835 141.275 211.005 141.445 ;
        RECT 211.835 141.275 212.005 141.445 ;
        RECT 212.835 141.275 213.005 141.445 ;
        RECT 213.835 141.275 214.005 141.445 ;
        RECT 214.835 141.275 215.005 141.445 ;
        RECT 215.835 141.275 216.005 141.445 ;
        RECT 216.835 141.275 217.005 141.445 ;
        RECT 217.835 141.275 218.005 141.445 ;
        RECT 218.835 141.275 219.005 141.445 ;
        RECT 219.835 141.275 220.005 141.445 ;
        RECT 220.835 141.275 221.005 141.445 ;
        RECT 221.835 141.275 222.005 141.445 ;
        RECT 222.835 141.275 223.005 141.445 ;
        RECT 223.835 141.275 224.005 141.445 ;
        RECT 224.835 141.275 225.005 141.445 ;
        RECT 225.835 141.275 226.005 141.445 ;
        RECT 226.835 141.275 227.005 141.445 ;
        RECT 227.835 141.275 228.005 141.445 ;
        RECT 228.835 141.275 229.005 141.445 ;
        RECT 229.835 141.275 230.005 141.445 ;
        RECT 230.835 141.275 231.005 141.445 ;
        RECT 231.835 141.275 232.005 141.445 ;
        RECT 232.835 141.275 233.005 141.445 ;
        RECT 233.835 141.275 234.005 141.445 ;
        RECT 234.835 141.275 235.005 141.445 ;
        RECT 235.835 141.275 236.005 141.445 ;
        RECT 236.835 141.275 237.005 141.445 ;
        RECT 237.835 141.275 238.005 141.445 ;
        RECT 238.835 141.275 239.005 141.445 ;
        RECT 239.835 141.275 240.005 141.445 ;
        RECT 240.835 141.275 241.005 141.445 ;
        RECT 241.835 141.275 242.005 141.445 ;
        RECT 242.835 141.275 243.005 141.445 ;
        RECT 243.835 141.275 244.005 141.445 ;
        RECT 244.835 141.275 245.005 141.445 ;
        RECT 245.835 141.275 246.005 141.445 ;
        RECT 246.835 141.275 247.005 141.445 ;
        RECT 247.835 141.275 248.005 141.445 ;
        RECT 248.835 141.275 249.005 141.445 ;
        RECT 249.835 141.275 250.005 141.445 ;
        RECT 250.835 141.275 251.005 141.445 ;
        RECT 251.835 141.275 252.005 141.445 ;
        RECT 252.835 141.275 253.005 141.445 ;
        RECT 253.835 141.275 254.005 141.445 ;
        RECT 254.835 141.275 255.005 141.445 ;
        RECT 255.835 141.275 256.005 141.445 ;
        RECT 256.835 141.275 257.005 141.445 ;
        RECT 257.835 141.275 258.005 141.445 ;
        RECT 258.835 141.275 259.005 141.445 ;
        RECT 259.835 141.275 260.005 141.445 ;
        RECT 260.835 141.275 261.005 141.445 ;
        RECT 261.835 141.275 262.005 141.445 ;
        RECT 129.440 129.275 129.610 129.445 ;
        RECT 129.440 128.915 129.610 129.085 ;
        RECT 129.440 128.555 129.610 128.725 ;
        RECT 129.440 128.195 129.610 128.365 ;
        RECT 129.440 127.835 129.610 128.005 ;
        RECT 129.440 127.475 129.610 127.645 ;
        RECT 129.440 127.115 129.610 127.285 ;
        RECT 129.440 126.755 129.610 126.925 ;
        RECT 129.440 126.395 129.610 126.565 ;
        RECT 129.440 126.035 129.610 126.205 ;
        RECT 129.440 125.675 129.610 125.845 ;
        RECT 134.020 129.275 134.190 129.445 ;
        RECT 134.020 128.915 134.190 129.085 ;
        RECT 134.020 128.555 134.190 128.725 ;
        RECT 134.020 128.195 134.190 128.365 ;
        RECT 134.020 127.835 134.190 128.005 ;
        RECT 134.020 127.475 134.190 127.645 ;
        RECT 134.020 127.115 134.190 127.285 ;
        RECT 134.020 126.755 134.190 126.925 ;
        RECT 134.020 126.395 134.190 126.565 ;
        RECT 134.020 126.035 134.190 126.205 ;
        RECT 134.020 125.675 134.190 125.845 ;
        RECT 138.600 129.275 138.770 129.445 ;
        RECT 138.600 128.915 138.770 129.085 ;
        RECT 138.600 128.555 138.770 128.725 ;
        RECT 138.600 128.195 138.770 128.365 ;
        RECT 138.600 127.835 138.770 128.005 ;
        RECT 138.600 127.475 138.770 127.645 ;
        RECT 138.600 127.115 138.770 127.285 ;
        RECT 138.600 126.755 138.770 126.925 ;
        RECT 138.600 126.395 138.770 126.565 ;
        RECT 138.600 126.035 138.770 126.205 ;
        RECT 138.600 125.675 138.770 125.845 ;
        RECT 143.180 129.275 143.350 129.445 ;
        RECT 143.180 128.915 143.350 129.085 ;
        RECT 143.180 128.555 143.350 128.725 ;
        RECT 143.180 128.195 143.350 128.365 ;
        RECT 143.180 127.835 143.350 128.005 ;
        RECT 143.180 127.475 143.350 127.645 ;
        RECT 143.180 127.115 143.350 127.285 ;
        RECT 143.180 126.755 143.350 126.925 ;
        RECT 143.180 126.395 143.350 126.565 ;
        RECT 143.180 126.035 143.350 126.205 ;
        RECT 143.180 125.675 143.350 125.845 ;
        RECT 147.760 129.275 147.930 129.445 ;
        RECT 147.760 128.915 147.930 129.085 ;
        RECT 147.760 128.555 147.930 128.725 ;
        RECT 147.760 128.195 147.930 128.365 ;
        RECT 147.760 127.835 147.930 128.005 ;
        RECT 147.760 127.475 147.930 127.645 ;
        RECT 147.760 127.115 147.930 127.285 ;
        RECT 147.760 126.755 147.930 126.925 ;
        RECT 147.760 126.395 147.930 126.565 ;
        RECT 147.760 126.035 147.930 126.205 ;
        RECT 147.760 125.675 147.930 125.845 ;
        RECT 112.915 122.475 113.085 122.645 ;
        RECT 113.915 122.475 114.085 122.645 ;
        RECT 114.915 122.475 115.085 122.645 ;
        RECT 115.915 122.475 116.085 122.645 ;
        RECT 116.915 122.475 117.085 122.645 ;
        RECT 117.915 122.475 118.085 122.645 ;
        RECT 118.915 122.475 119.085 122.645 ;
        RECT 119.915 122.475 120.085 122.645 ;
        RECT 120.915 122.475 121.085 122.645 ;
        RECT 121.915 122.475 122.085 122.645 ;
        RECT 122.915 122.475 123.085 122.645 ;
        RECT 128.005 122.475 128.175 122.645 ;
        RECT 130.005 122.475 130.175 122.645 ;
        RECT 132.005 122.475 132.175 122.645 ;
        RECT 134.005 122.475 134.175 122.645 ;
        RECT 136.005 122.475 136.175 122.645 ;
        RECT 138.005 122.475 138.175 122.645 ;
        RECT 140.005 122.475 140.175 122.645 ;
        RECT 142.005 122.475 142.175 122.645 ;
        RECT 144.005 122.475 144.175 122.645 ;
        RECT 146.005 122.475 146.175 122.645 ;
        RECT 150.555 122.475 150.725 122.645 ;
        RECT 152.555 122.475 152.725 122.645 ;
        RECT 154.555 122.475 154.725 122.645 ;
        RECT 156.555 122.475 156.725 122.645 ;
        RECT 158.555 122.475 158.725 122.645 ;
        RECT 160.555 122.475 160.725 122.645 ;
        RECT 162.555 122.475 162.725 122.645 ;
        RECT 164.555 122.475 164.725 122.645 ;
        RECT 166.555 122.475 166.725 122.645 ;
        RECT 168.555 122.475 168.725 122.645 ;
        RECT 170.555 122.475 170.725 122.645 ;
        RECT 172.555 122.475 172.725 122.645 ;
        RECT 174.555 122.475 174.725 122.645 ;
        RECT 176.555 122.475 176.725 122.645 ;
        RECT 178.555 122.475 178.725 122.645 ;
        RECT 180.555 122.475 180.725 122.645 ;
        RECT 182.555 122.475 182.725 122.645 ;
        RECT 184.555 122.475 184.725 122.645 ;
        RECT 187.885 122.475 188.055 122.645 ;
        RECT 188.885 122.475 189.055 122.645 ;
        RECT 189.885 122.475 190.055 122.645 ;
        RECT 190.885 122.475 191.055 122.645 ;
        RECT 191.885 122.475 192.055 122.645 ;
        RECT 192.885 122.475 193.055 122.645 ;
        RECT 193.885 122.475 194.055 122.645 ;
        RECT 194.885 122.475 195.055 122.645 ;
        RECT 195.885 122.475 196.055 122.645 ;
        RECT 196.885 122.475 197.055 122.645 ;
        RECT 197.885 122.475 198.055 122.645 ;
        RECT 201.605 122.475 201.775 122.645 ;
        RECT 202.605 122.475 202.775 122.645 ;
        RECT 203.605 122.475 203.775 122.645 ;
        RECT 204.605 122.475 204.775 122.645 ;
        RECT 205.605 122.475 205.775 122.645 ;
        RECT 206.605 122.475 206.775 122.645 ;
        RECT 207.605 122.475 207.775 122.645 ;
        RECT 208.605 122.475 208.775 122.645 ;
        RECT 209.605 122.475 209.775 122.645 ;
        RECT 210.605 122.475 210.775 122.645 ;
        RECT 211.605 122.475 211.775 122.645 ;
        RECT 215.325 122.475 215.495 122.645 ;
        RECT 216.325 122.475 216.495 122.645 ;
        RECT 217.325 122.475 217.495 122.645 ;
        RECT 218.325 122.475 218.495 122.645 ;
        RECT 219.325 122.475 219.495 122.645 ;
        RECT 220.325 122.475 220.495 122.645 ;
        RECT 221.325 122.475 221.495 122.645 ;
        RECT 222.325 122.475 222.495 122.645 ;
        RECT 223.325 122.475 223.495 122.645 ;
        RECT 224.325 122.475 224.495 122.645 ;
        RECT 225.325 122.475 225.495 122.645 ;
        RECT 229.045 122.475 229.215 122.645 ;
        RECT 230.045 122.475 230.215 122.645 ;
        RECT 231.045 122.475 231.215 122.645 ;
        RECT 232.045 122.475 232.215 122.645 ;
        RECT 233.045 122.475 233.215 122.645 ;
        RECT 234.045 122.475 234.215 122.645 ;
        RECT 235.045 122.475 235.215 122.645 ;
        RECT 236.045 122.475 236.215 122.645 ;
        RECT 237.045 122.475 237.215 122.645 ;
        RECT 238.045 122.475 238.215 122.645 ;
        RECT 239.045 122.475 239.215 122.645 ;
        RECT 242.765 122.475 242.935 122.645 ;
        RECT 243.765 122.475 243.935 122.645 ;
        RECT 244.765 122.475 244.935 122.645 ;
        RECT 245.765 122.475 245.935 122.645 ;
        RECT 246.765 122.475 246.935 122.645 ;
        RECT 247.765 122.475 247.935 122.645 ;
        RECT 248.765 122.475 248.935 122.645 ;
        RECT 249.765 122.475 249.935 122.645 ;
        RECT 250.765 122.475 250.935 122.645 ;
        RECT 251.765 122.475 251.935 122.645 ;
        RECT 252.765 122.475 252.935 122.645 ;
        RECT 120.265 103.675 120.435 103.845 ;
        RECT 121.265 103.675 121.435 103.845 ;
        RECT 122.265 103.675 122.435 103.845 ;
        RECT 123.265 103.675 123.435 103.845 ;
        RECT 124.265 103.675 124.435 103.845 ;
        RECT 125.265 103.675 125.435 103.845 ;
        RECT 126.265 103.675 126.435 103.845 ;
        RECT 127.265 103.675 127.435 103.845 ;
        RECT 128.265 103.675 128.435 103.845 ;
        RECT 129.265 103.675 129.435 103.845 ;
        RECT 130.265 103.675 130.435 103.845 ;
        RECT 136.925 103.675 137.095 103.845 ;
        RECT 137.925 103.675 138.095 103.845 ;
        RECT 138.925 103.675 139.095 103.845 ;
        RECT 139.925 103.675 140.095 103.845 ;
        RECT 140.925 103.675 141.095 103.845 ;
        RECT 141.925 103.675 142.095 103.845 ;
        RECT 142.925 103.675 143.095 103.845 ;
        RECT 143.925 103.675 144.095 103.845 ;
        RECT 144.925 103.675 145.095 103.845 ;
        RECT 145.925 103.675 146.095 103.845 ;
        RECT 146.925 103.675 147.095 103.845 ;
        RECT 150.645 103.675 150.815 103.845 ;
        RECT 151.645 103.675 151.815 103.845 ;
        RECT 152.645 103.675 152.815 103.845 ;
        RECT 153.645 103.675 153.815 103.845 ;
        RECT 154.645 103.675 154.815 103.845 ;
        RECT 155.645 103.675 155.815 103.845 ;
        RECT 156.645 103.675 156.815 103.845 ;
        RECT 157.645 103.675 157.815 103.845 ;
        RECT 158.645 103.675 158.815 103.845 ;
        RECT 159.645 103.675 159.815 103.845 ;
        RECT 160.645 103.675 160.815 103.845 ;
        RECT 166.815 103.675 166.985 103.845 ;
        RECT 167.815 103.675 167.985 103.845 ;
        RECT 168.815 103.675 168.985 103.845 ;
        RECT 169.815 103.675 169.985 103.845 ;
        RECT 170.815 103.675 170.985 103.845 ;
        RECT 171.815 103.675 171.985 103.845 ;
        RECT 172.815 103.675 172.985 103.845 ;
        RECT 173.815 103.675 173.985 103.845 ;
        RECT 174.815 103.675 174.985 103.845 ;
        RECT 175.815 103.675 175.985 103.845 ;
        RECT 176.815 103.675 176.985 103.845 ;
        RECT 187.885 103.675 188.055 103.845 ;
        RECT 188.885 103.675 189.055 103.845 ;
        RECT 189.885 103.675 190.055 103.845 ;
        RECT 190.885 103.675 191.055 103.845 ;
        RECT 191.885 103.675 192.055 103.845 ;
        RECT 192.885 103.675 193.055 103.845 ;
        RECT 193.885 103.675 194.055 103.845 ;
        RECT 194.885 103.675 195.055 103.845 ;
        RECT 195.885 103.675 196.055 103.845 ;
        RECT 196.885 103.675 197.055 103.845 ;
        RECT 197.885 103.675 198.055 103.845 ;
        RECT 201.605 103.675 201.775 103.845 ;
        RECT 202.605 103.675 202.775 103.845 ;
        RECT 203.605 103.675 203.775 103.845 ;
        RECT 204.605 103.675 204.775 103.845 ;
        RECT 205.605 103.675 205.775 103.845 ;
        RECT 206.605 103.675 206.775 103.845 ;
        RECT 207.605 103.675 207.775 103.845 ;
        RECT 208.605 103.675 208.775 103.845 ;
        RECT 209.605 103.675 209.775 103.845 ;
        RECT 210.605 103.675 210.775 103.845 ;
        RECT 211.605 103.675 211.775 103.845 ;
        RECT 242.765 103.675 242.935 103.845 ;
        RECT 243.765 103.675 243.935 103.845 ;
        RECT 244.765 103.675 244.935 103.845 ;
        RECT 245.765 103.675 245.935 103.845 ;
        RECT 246.765 103.675 246.935 103.845 ;
        RECT 247.765 103.675 247.935 103.845 ;
        RECT 248.765 103.675 248.935 103.845 ;
        RECT 249.765 103.675 249.935 103.845 ;
        RECT 250.765 103.675 250.935 103.845 ;
        RECT 251.765 103.675 251.935 103.845 ;
        RECT 252.765 103.675 252.935 103.845 ;
        RECT 125.065 84.875 125.235 85.045 ;
        RECT 127.065 84.875 127.235 85.045 ;
        RECT 129.065 84.875 129.235 85.045 ;
        RECT 131.065 84.875 131.235 85.045 ;
        RECT 133.065 84.875 133.235 85.045 ;
        RECT 135.065 84.875 135.235 85.045 ;
        RECT 137.065 84.875 137.235 85.045 ;
        RECT 139.065 84.875 139.235 85.045 ;
        RECT 141.065 84.875 141.235 85.045 ;
        RECT 143.065 84.875 143.235 85.045 ;
        RECT 145.065 84.875 145.235 85.045 ;
        RECT 147.065 84.875 147.235 85.045 ;
        RECT 149.065 84.875 149.235 85.045 ;
        RECT 151.065 84.875 151.235 85.045 ;
        RECT 153.065 84.875 153.235 85.045 ;
        RECT 155.065 84.875 155.235 85.045 ;
        RECT 157.065 84.875 157.235 85.045 ;
        RECT 159.065 84.875 159.235 85.045 ;
        RECT 161.065 84.875 161.235 85.045 ;
        RECT 163.065 84.875 163.235 85.045 ;
        RECT 165.065 84.875 165.235 85.045 ;
        RECT 167.065 84.875 167.235 85.045 ;
        RECT 169.065 84.875 169.235 85.045 ;
        RECT 171.065 84.875 171.235 85.045 ;
        RECT 173.065 84.875 173.235 85.045 ;
        RECT 175.065 84.875 175.235 85.045 ;
        RECT 177.065 84.875 177.235 85.045 ;
        RECT 179.065 84.875 179.235 85.045 ;
        RECT 181.065 84.875 181.235 85.045 ;
        RECT 183.065 84.875 183.235 85.045 ;
        RECT 185.065 84.875 185.235 85.045 ;
        RECT 187.065 84.875 187.235 85.045 ;
        RECT 189.065 84.875 189.235 85.045 ;
        RECT 191.065 84.875 191.235 85.045 ;
        RECT 193.065 84.875 193.235 85.045 ;
        RECT 195.065 84.875 195.235 85.045 ;
        RECT 197.065 84.875 197.235 85.045 ;
        RECT 199.065 84.875 199.235 85.045 ;
        RECT 201.065 84.875 201.235 85.045 ;
        RECT 203.065 84.875 203.235 85.045 ;
        RECT 205.065 84.875 205.235 85.045 ;
        RECT 207.065 84.875 207.235 85.045 ;
        RECT 209.065 84.875 209.235 85.045 ;
        RECT 211.065 84.875 211.235 85.045 ;
        RECT 213.065 84.875 213.235 85.045 ;
        RECT 215.065 84.875 215.235 85.045 ;
        RECT 217.065 84.875 217.235 85.045 ;
        RECT 219.065 84.875 219.235 85.045 ;
        RECT 221.065 84.875 221.235 85.045 ;
        RECT 223.065 84.875 223.235 85.045 ;
        RECT 225.065 84.875 225.235 85.045 ;
        RECT 227.065 84.875 227.235 85.045 ;
        RECT 229.065 84.875 229.235 85.045 ;
        RECT 231.065 84.875 231.235 85.045 ;
        RECT 233.065 84.875 233.235 85.045 ;
        RECT 235.065 84.875 235.235 85.045 ;
        RECT 237.065 84.875 237.235 85.045 ;
        RECT 239.065 84.875 239.235 85.045 ;
        RECT 241.065 84.875 241.235 85.045 ;
        RECT 243.065 84.875 243.235 85.045 ;
        RECT 245.065 84.875 245.235 85.045 ;
        RECT 247.065 84.875 247.235 85.045 ;
        RECT 249.065 84.875 249.235 85.045 ;
        RECT 251.065 84.875 251.235 85.045 ;
        RECT 253.065 84.875 253.235 85.045 ;
        RECT 255.065 84.875 255.235 85.045 ;
        RECT 257.065 84.875 257.235 85.045 ;
        RECT 259.065 84.875 259.235 85.045 ;
        RECT 261.065 84.875 261.235 85.045 ;
        RECT 220.225 66.075 220.395 66.245 ;
        RECT 221.225 66.075 221.395 66.245 ;
        RECT 222.225 66.075 222.395 66.245 ;
        RECT 223.225 66.075 223.395 66.245 ;
        RECT 224.225 66.075 224.395 66.245 ;
        RECT 225.225 66.075 225.395 66.245 ;
        RECT 226.225 66.075 226.395 66.245 ;
        RECT 227.225 66.075 227.395 66.245 ;
        RECT 228.225 66.075 228.395 66.245 ;
        RECT 229.225 66.075 229.395 66.245 ;
        RECT 230.225 66.075 230.395 66.245 ;
        RECT 233.945 66.075 234.115 66.245 ;
        RECT 234.945 66.075 235.115 66.245 ;
        RECT 235.945 66.075 236.115 66.245 ;
        RECT 236.945 66.075 237.115 66.245 ;
        RECT 237.945 66.075 238.115 66.245 ;
        RECT 238.945 66.075 239.115 66.245 ;
        RECT 239.945 66.075 240.115 66.245 ;
        RECT 240.945 66.075 241.115 66.245 ;
        RECT 241.945 66.075 242.115 66.245 ;
        RECT 242.945 66.075 243.115 66.245 ;
        RECT 243.945 66.075 244.115 66.245 ;
        RECT 247.665 66.075 247.835 66.245 ;
        RECT 248.665 66.075 248.835 66.245 ;
        RECT 249.665 66.075 249.835 66.245 ;
        RECT 250.665 66.075 250.835 66.245 ;
        RECT 251.665 66.075 251.835 66.245 ;
        RECT 252.665 66.075 252.835 66.245 ;
        RECT 253.665 66.075 253.835 66.245 ;
        RECT 254.665 66.075 254.835 66.245 ;
        RECT 255.665 66.075 255.835 66.245 ;
        RECT 256.665 66.075 256.835 66.245 ;
        RECT 257.665 66.075 257.835 66.245 ;
        RECT 219.735 47.275 219.905 47.445 ;
        RECT 220.735 47.275 220.905 47.445 ;
        RECT 221.735 47.275 221.905 47.445 ;
        RECT 222.735 47.275 222.905 47.445 ;
        RECT 223.735 47.275 223.905 47.445 ;
        RECT 224.735 47.275 224.905 47.445 ;
        RECT 225.735 47.275 225.905 47.445 ;
        RECT 226.735 47.275 226.905 47.445 ;
        RECT 227.735 47.275 227.905 47.445 ;
        RECT 228.735 47.275 228.905 47.445 ;
        RECT 229.735 47.275 229.905 47.445 ;
        RECT 233.455 47.275 233.625 47.445 ;
        RECT 234.455 47.275 234.625 47.445 ;
        RECT 235.455 47.275 235.625 47.445 ;
        RECT 236.455 47.275 236.625 47.445 ;
        RECT 237.455 47.275 237.625 47.445 ;
        RECT 238.455 47.275 238.625 47.445 ;
        RECT 239.455 47.275 239.625 47.445 ;
        RECT 240.455 47.275 240.625 47.445 ;
        RECT 241.455 47.275 241.625 47.445 ;
        RECT 242.455 47.275 242.625 47.445 ;
        RECT 243.455 47.275 243.625 47.445 ;
        RECT 247.175 47.275 247.345 47.445 ;
        RECT 248.175 47.275 248.345 47.445 ;
        RECT 249.175 47.275 249.345 47.445 ;
        RECT 250.175 47.275 250.345 47.445 ;
        RECT 251.175 47.275 251.345 47.445 ;
        RECT 252.175 47.275 252.345 47.445 ;
        RECT 253.175 47.275 253.345 47.445 ;
        RECT 254.175 47.275 254.345 47.445 ;
        RECT 255.175 47.275 255.345 47.445 ;
        RECT 256.175 47.275 256.345 47.445 ;
        RECT 257.175 47.275 257.345 47.445 ;
        RECT 236.555 29.215 238.525 31.905 ;
        RECT 223.655 28.475 223.825 28.645 ;
        RECT 224.655 28.475 224.825 28.645 ;
        RECT 225.655 28.475 225.825 28.645 ;
        RECT 226.655 28.475 226.825 28.645 ;
        RECT 227.655 28.475 227.825 28.645 ;
        RECT 228.655 28.475 228.825 28.645 ;
        RECT 229.655 28.475 229.825 28.645 ;
        RECT 230.655 28.475 230.825 28.645 ;
        RECT 231.655 28.475 231.825 28.645 ;
        RECT 232.655 28.475 232.825 28.645 ;
        RECT 233.655 28.475 233.825 28.645 ;
        RECT 237.375 28.475 237.545 28.645 ;
        RECT 238.375 28.475 238.545 28.645 ;
        RECT 239.375 28.475 239.545 28.645 ;
        RECT 240.375 28.475 240.545 28.645 ;
        RECT 241.375 28.475 241.545 28.645 ;
        RECT 242.375 28.475 242.545 28.645 ;
        RECT 243.375 28.475 243.545 28.645 ;
        RECT 244.375 28.475 244.545 28.645 ;
        RECT 245.375 28.475 245.545 28.645 ;
        RECT 246.375 28.475 246.545 28.645 ;
        RECT 247.375 28.475 247.545 28.645 ;
        RECT 251.095 28.475 251.265 28.645 ;
        RECT 252.095 28.475 252.265 28.645 ;
        RECT 253.095 28.475 253.265 28.645 ;
        RECT 254.095 28.475 254.265 28.645 ;
        RECT 255.095 28.475 255.265 28.645 ;
        RECT 256.095 28.475 256.265 28.645 ;
        RECT 257.095 28.475 257.265 28.645 ;
        RECT 258.095 28.475 258.265 28.645 ;
        RECT 259.095 28.475 259.265 28.645 ;
        RECT 260.095 28.475 260.265 28.645 ;
        RECT 261.095 28.475 261.265 28.645 ;
      LAYER met1 ;
        RECT 4.500 253.860 287.680 254.460 ;
        RECT 121.910 238.580 122.140 242.360 ;
        RECT 121.600 238.440 122.140 238.580 ;
        RECT 121.600 235.660 121.740 238.440 ;
        RECT 121.910 238.360 122.140 238.440 ;
        RECT 4.500 235.060 287.680 235.660 ;
        RECT 214.930 224.060 261.570 224.410 ;
        RECT 216.360 223.680 216.500 224.060 ;
        RECT 216.270 223.660 216.590 223.680 ;
        RECT 72.910 219.880 73.140 223.560 ;
        RECT 215.750 223.310 260.750 223.660 ;
        RECT 72.910 219.740 73.440 219.880 ;
        RECT 72.910 219.560 73.140 219.740 ;
        RECT 73.300 216.860 73.440 219.740 ;
        RECT 4.500 216.260 287.680 216.860 ;
        RECT 209.830 205.610 210.150 205.660 ;
        RECT 209.050 205.260 262.390 205.610 ;
        RECT 209.870 204.640 261.570 204.860 ;
        RECT 209.830 204.510 261.570 204.640 ;
        RECT 209.830 204.380 210.150 204.510 ;
        RECT 4.500 197.460 287.680 198.060 ;
        RECT 209.050 186.460 262.390 186.810 ;
        RECT 209.920 186.060 210.060 186.460 ;
        RECT 209.870 185.940 261.570 186.060 ;
        RECT 209.830 185.710 261.570 185.940 ;
        RECT 209.830 185.680 210.150 185.710 ;
        RECT 65.405 181.275 65.695 181.505 ;
        RECT 65.480 180.780 65.620 181.275 ;
        RECT 66.325 180.780 66.615 180.825 ;
        RECT 65.480 180.640 66.615 180.780 ;
        RECT 66.325 180.595 66.615 180.640 ;
        RECT 66.400 179.260 66.540 180.595 ;
        RECT 95.890 179.555 97.940 182.365 ;
        RECT 96.300 179.260 96.440 179.555 ;
        RECT 4.500 178.660 287.680 179.260 ;
        RECT 209.050 167.660 262.390 168.010 ;
        RECT 213.600 167.260 213.740 167.660 ;
        RECT 209.870 166.910 261.570 167.260 ;
        RECT 110.100 160.755 112.150 163.565 ;
        RECT 111.940 160.460 112.080 160.755 ;
        RECT 4.500 159.860 287.680 160.460 ;
        RECT 209.050 148.860 262.390 149.210 ;
        RECT 210.840 148.540 210.980 148.860 ;
        RECT 210.750 148.460 211.070 148.540 ;
        RECT 209.870 148.110 261.570 148.460 ;
        RECT 4.500 141.060 287.680 141.660 ;
        RECT 129.410 125.560 129.640 129.560 ;
        RECT 133.990 125.560 134.220 129.560 ;
        RECT 138.570 125.560 138.800 129.560 ;
        RECT 143.150 125.560 143.380 129.560 ;
        RECT 147.730 125.560 147.960 129.560 ;
        RECT 129.420 122.860 129.560 125.560 ;
        RECT 4.500 122.260 287.680 122.860 ;
        RECT 4.500 103.460 287.680 104.060 ;
        RECT 4.500 84.660 287.680 85.260 ;
        RECT 4.500 65.860 287.680 66.460 ;
        RECT 4.500 47.060 287.680 47.660 ;
        RECT 236.515 29.155 238.565 31.965 ;
        RECT 236.600 28.860 236.740 29.155 ;
        RECT 4.500 28.260 287.680 28.860 ;
      LAYER via ;
        RECT 4.610 253.870 12.550 254.450 ;
        RECT 279.630 253.870 287.570 254.450 ;
        RECT 4.610 235.070 12.550 235.650 ;
        RECT 88.420 235.320 88.680 235.580 ;
        RECT 279.630 235.070 287.570 235.650 ;
        RECT 216.300 223.420 216.560 223.680 ;
        RECT 4.610 216.270 12.550 216.850 ;
        RECT 41.500 216.280 41.760 216.540 ;
        RECT 216.300 216.280 216.560 216.540 ;
        RECT 279.630 216.270 287.570 216.850 ;
        RECT 209.860 205.400 210.120 205.660 ;
        RECT 209.860 204.380 210.120 204.640 ;
        RECT 4.610 197.470 12.550 198.050 ;
        RECT 77.380 197.580 77.640 197.840 ;
        RECT 209.860 197.580 210.120 197.840 ;
        RECT 279.630 197.470 287.570 198.050 ;
        RECT 209.860 185.680 210.120 185.940 ;
        RECT 4.610 178.670 12.550 179.250 ;
        RECT 209.860 178.880 210.120 179.140 ;
        RECT 279.630 178.670 287.570 179.250 ;
        RECT 209.400 167.660 209.660 167.920 ;
        RECT 4.610 159.870 12.550 160.450 ;
        RECT 279.630 159.870 287.570 160.450 ;
        RECT 210.780 148.280 211.040 148.540 ;
        RECT 4.610 141.070 12.550 141.650 ;
        RECT 210.780 141.140 211.040 141.400 ;
        RECT 279.630 141.070 287.570 141.650 ;
        RECT 4.610 122.270 12.550 122.850 ;
        RECT 279.630 122.270 287.570 122.850 ;
        RECT 4.610 103.470 12.550 104.050 ;
        RECT 279.630 103.470 287.570 104.050 ;
        RECT 4.610 84.670 12.550 85.250 ;
        RECT 279.630 84.670 287.570 85.250 ;
        RECT 4.610 65.870 12.550 66.450 ;
        RECT 279.630 65.870 287.570 66.450 ;
        RECT 4.610 47.070 12.550 47.650 ;
        RECT 279.630 47.070 287.570 47.650 ;
        RECT 4.610 28.270 12.550 28.850 ;
        RECT 279.630 28.270 287.570 28.850 ;
      LAYER met2 ;
        RECT 4.500 253.860 12.660 254.460 ;
        RECT 279.520 253.860 287.680 254.460 ;
        RECT 29.690 236.060 30.490 236.560 ;
        RECT 66.930 236.060 67.730 236.560 ;
        RECT 4.500 235.060 12.660 235.660 ;
        RECT 88.410 235.335 88.690 235.705 ;
        RECT 88.420 235.290 88.680 235.335 ;
        RECT 88.480 235.220 88.620 235.290 ;
        RECT 279.520 235.060 287.680 235.660 ;
        RECT 216.300 223.390 216.560 223.710 ;
        RECT 29.690 217.260 30.490 217.760 ;
        RECT 4.500 216.260 12.660 216.860 ;
        RECT 41.490 216.425 41.770 216.795 ;
        RECT 216.360 216.570 216.500 223.390 ;
        RECT 41.500 216.250 41.760 216.425 ;
        RECT 216.300 216.250 216.560 216.570 ;
        RECT 279.520 216.260 287.680 216.860 ;
        RECT 209.860 205.370 210.120 205.690 ;
        RECT 209.920 204.670 210.060 205.370 ;
        RECT 209.860 204.350 210.120 204.670 ;
        RECT 31.650 198.460 32.450 198.960 ;
        RECT 75.750 198.460 76.550 198.960 ;
        RECT 77.370 198.125 77.650 198.495 ;
        RECT 4.500 197.460 12.660 198.060 ;
        RECT 77.440 197.870 77.580 198.125 ;
        RECT 209.920 197.870 210.060 204.350 ;
        RECT 77.380 197.550 77.640 197.870 ;
        RECT 209.860 197.550 210.120 197.870 ;
        RECT 279.520 197.460 287.680 198.060 ;
        RECT 209.860 185.650 210.120 185.970 ;
        RECT 4.500 178.660 12.660 179.260 ;
        RECT 209.920 179.170 210.060 185.650 ;
        RECT 209.860 178.850 210.120 179.170 ;
        RECT 209.920 168.880 210.060 178.850 ;
        RECT 279.520 178.660 287.680 179.260 ;
        RECT 209.460 168.740 210.060 168.880 ;
        RECT 209.460 167.950 209.600 168.740 ;
        RECT 209.400 167.630 209.660 167.950 ;
        RECT 4.500 159.860 12.660 160.460 ;
        RECT 279.520 159.860 287.680 160.460 ;
        RECT 210.780 148.250 211.040 148.570 ;
        RECT 4.500 141.060 12.660 141.660 ;
        RECT 210.840 141.430 210.980 148.250 ;
        RECT 210.780 141.110 211.040 141.430 ;
        RECT 279.520 141.060 287.680 141.660 ;
        RECT 4.500 122.260 12.660 122.860 ;
        RECT 279.520 122.260 287.680 122.860 ;
        RECT 4.500 103.460 12.660 104.060 ;
        RECT 279.520 103.460 287.680 104.060 ;
        RECT 4.500 84.660 12.660 85.260 ;
        RECT 279.520 84.660 287.680 85.260 ;
        RECT 4.500 65.860 12.660 66.460 ;
        RECT 279.520 65.860 287.680 66.460 ;
        RECT 4.500 47.060 12.660 47.660 ;
        RECT 279.520 47.060 287.680 47.660 ;
        RECT 4.500 28.260 12.660 28.860 ;
        RECT 279.520 28.260 287.680 28.860 ;
      LAYER via2 ;
        RECT 4.640 254.020 4.920 254.300 ;
        RECT 5.040 254.020 5.320 254.300 ;
        RECT 5.440 254.020 5.720 254.300 ;
        RECT 5.840 254.020 6.120 254.300 ;
        RECT 6.240 254.020 6.520 254.300 ;
        RECT 6.640 254.020 6.920 254.300 ;
        RECT 7.040 254.020 7.320 254.300 ;
        RECT 7.440 254.020 7.720 254.300 ;
        RECT 7.840 254.020 8.120 254.300 ;
        RECT 8.240 254.020 8.520 254.300 ;
        RECT 8.640 254.020 8.920 254.300 ;
        RECT 9.040 254.020 9.320 254.300 ;
        RECT 9.440 254.020 9.720 254.300 ;
        RECT 9.840 254.020 10.120 254.300 ;
        RECT 10.240 254.020 10.520 254.300 ;
        RECT 10.640 254.020 10.920 254.300 ;
        RECT 11.040 254.020 11.320 254.300 ;
        RECT 11.440 254.020 11.720 254.300 ;
        RECT 11.840 254.020 12.120 254.300 ;
        RECT 12.240 254.020 12.520 254.300 ;
        RECT 279.660 254.020 279.940 254.300 ;
        RECT 280.060 254.020 280.340 254.300 ;
        RECT 280.460 254.020 280.740 254.300 ;
        RECT 280.860 254.020 281.140 254.300 ;
        RECT 281.260 254.020 281.540 254.300 ;
        RECT 281.660 254.020 281.940 254.300 ;
        RECT 282.060 254.020 282.340 254.300 ;
        RECT 282.460 254.020 282.740 254.300 ;
        RECT 282.860 254.020 283.140 254.300 ;
        RECT 283.260 254.020 283.540 254.300 ;
        RECT 283.660 254.020 283.940 254.300 ;
        RECT 284.060 254.020 284.340 254.300 ;
        RECT 284.460 254.020 284.740 254.300 ;
        RECT 284.860 254.020 285.140 254.300 ;
        RECT 285.260 254.020 285.540 254.300 ;
        RECT 285.660 254.020 285.940 254.300 ;
        RECT 286.060 254.020 286.340 254.300 ;
        RECT 286.460 254.020 286.740 254.300 ;
        RECT 286.860 254.020 287.140 254.300 ;
        RECT 287.260 254.020 287.540 254.300 ;
        RECT 29.950 236.170 30.230 236.450 ;
        RECT 67.190 236.170 67.470 236.450 ;
        RECT 4.640 235.220 4.920 235.500 ;
        RECT 5.040 235.220 5.320 235.500 ;
        RECT 5.440 235.220 5.720 235.500 ;
        RECT 5.840 235.220 6.120 235.500 ;
        RECT 6.240 235.220 6.520 235.500 ;
        RECT 6.640 235.220 6.920 235.500 ;
        RECT 7.040 235.220 7.320 235.500 ;
        RECT 7.440 235.220 7.720 235.500 ;
        RECT 7.840 235.220 8.120 235.500 ;
        RECT 8.240 235.220 8.520 235.500 ;
        RECT 8.640 235.220 8.920 235.500 ;
        RECT 9.040 235.220 9.320 235.500 ;
        RECT 9.440 235.220 9.720 235.500 ;
        RECT 9.840 235.220 10.120 235.500 ;
        RECT 10.240 235.220 10.520 235.500 ;
        RECT 10.640 235.220 10.920 235.500 ;
        RECT 11.040 235.220 11.320 235.500 ;
        RECT 11.440 235.220 11.720 235.500 ;
        RECT 11.840 235.220 12.120 235.500 ;
        RECT 12.240 235.220 12.520 235.500 ;
        RECT 88.410 235.380 88.690 235.660 ;
        RECT 279.660 235.220 279.940 235.500 ;
        RECT 280.060 235.220 280.340 235.500 ;
        RECT 280.460 235.220 280.740 235.500 ;
        RECT 280.860 235.220 281.140 235.500 ;
        RECT 281.260 235.220 281.540 235.500 ;
        RECT 281.660 235.220 281.940 235.500 ;
        RECT 282.060 235.220 282.340 235.500 ;
        RECT 282.460 235.220 282.740 235.500 ;
        RECT 282.860 235.220 283.140 235.500 ;
        RECT 283.260 235.220 283.540 235.500 ;
        RECT 283.660 235.220 283.940 235.500 ;
        RECT 284.060 235.220 284.340 235.500 ;
        RECT 284.460 235.220 284.740 235.500 ;
        RECT 284.860 235.220 285.140 235.500 ;
        RECT 285.260 235.220 285.540 235.500 ;
        RECT 285.660 235.220 285.940 235.500 ;
        RECT 286.060 235.220 286.340 235.500 ;
        RECT 286.460 235.220 286.740 235.500 ;
        RECT 286.860 235.220 287.140 235.500 ;
        RECT 287.260 235.220 287.540 235.500 ;
        RECT 29.950 217.370 30.230 217.650 ;
        RECT 4.640 216.420 4.920 216.700 ;
        RECT 5.040 216.420 5.320 216.700 ;
        RECT 5.440 216.420 5.720 216.700 ;
        RECT 5.840 216.420 6.120 216.700 ;
        RECT 6.240 216.420 6.520 216.700 ;
        RECT 6.640 216.420 6.920 216.700 ;
        RECT 7.040 216.420 7.320 216.700 ;
        RECT 7.440 216.420 7.720 216.700 ;
        RECT 7.840 216.420 8.120 216.700 ;
        RECT 8.240 216.420 8.520 216.700 ;
        RECT 8.640 216.420 8.920 216.700 ;
        RECT 9.040 216.420 9.320 216.700 ;
        RECT 9.440 216.420 9.720 216.700 ;
        RECT 9.840 216.420 10.120 216.700 ;
        RECT 10.240 216.420 10.520 216.700 ;
        RECT 10.640 216.420 10.920 216.700 ;
        RECT 11.040 216.420 11.320 216.700 ;
        RECT 11.440 216.420 11.720 216.700 ;
        RECT 11.840 216.420 12.120 216.700 ;
        RECT 12.240 216.420 12.520 216.700 ;
        RECT 41.490 216.470 41.770 216.750 ;
        RECT 279.660 216.420 279.940 216.700 ;
        RECT 280.060 216.420 280.340 216.700 ;
        RECT 280.460 216.420 280.740 216.700 ;
        RECT 280.860 216.420 281.140 216.700 ;
        RECT 281.260 216.420 281.540 216.700 ;
        RECT 281.660 216.420 281.940 216.700 ;
        RECT 282.060 216.420 282.340 216.700 ;
        RECT 282.460 216.420 282.740 216.700 ;
        RECT 282.860 216.420 283.140 216.700 ;
        RECT 283.260 216.420 283.540 216.700 ;
        RECT 283.660 216.420 283.940 216.700 ;
        RECT 284.060 216.420 284.340 216.700 ;
        RECT 284.460 216.420 284.740 216.700 ;
        RECT 284.860 216.420 285.140 216.700 ;
        RECT 285.260 216.420 285.540 216.700 ;
        RECT 285.660 216.420 285.940 216.700 ;
        RECT 286.060 216.420 286.340 216.700 ;
        RECT 286.460 216.420 286.740 216.700 ;
        RECT 286.860 216.420 287.140 216.700 ;
        RECT 287.260 216.420 287.540 216.700 ;
        RECT 31.910 198.570 32.190 198.850 ;
        RECT 76.010 198.570 76.290 198.850 ;
        RECT 77.370 198.170 77.650 198.450 ;
        RECT 4.640 197.620 4.920 197.900 ;
        RECT 5.040 197.620 5.320 197.900 ;
        RECT 5.440 197.620 5.720 197.900 ;
        RECT 5.840 197.620 6.120 197.900 ;
        RECT 6.240 197.620 6.520 197.900 ;
        RECT 6.640 197.620 6.920 197.900 ;
        RECT 7.040 197.620 7.320 197.900 ;
        RECT 7.440 197.620 7.720 197.900 ;
        RECT 7.840 197.620 8.120 197.900 ;
        RECT 8.240 197.620 8.520 197.900 ;
        RECT 8.640 197.620 8.920 197.900 ;
        RECT 9.040 197.620 9.320 197.900 ;
        RECT 9.440 197.620 9.720 197.900 ;
        RECT 9.840 197.620 10.120 197.900 ;
        RECT 10.240 197.620 10.520 197.900 ;
        RECT 10.640 197.620 10.920 197.900 ;
        RECT 11.040 197.620 11.320 197.900 ;
        RECT 11.440 197.620 11.720 197.900 ;
        RECT 11.840 197.620 12.120 197.900 ;
        RECT 12.240 197.620 12.520 197.900 ;
        RECT 279.660 197.620 279.940 197.900 ;
        RECT 280.060 197.620 280.340 197.900 ;
        RECT 280.460 197.620 280.740 197.900 ;
        RECT 280.860 197.620 281.140 197.900 ;
        RECT 281.260 197.620 281.540 197.900 ;
        RECT 281.660 197.620 281.940 197.900 ;
        RECT 282.060 197.620 282.340 197.900 ;
        RECT 282.460 197.620 282.740 197.900 ;
        RECT 282.860 197.620 283.140 197.900 ;
        RECT 283.260 197.620 283.540 197.900 ;
        RECT 283.660 197.620 283.940 197.900 ;
        RECT 284.060 197.620 284.340 197.900 ;
        RECT 284.460 197.620 284.740 197.900 ;
        RECT 284.860 197.620 285.140 197.900 ;
        RECT 285.260 197.620 285.540 197.900 ;
        RECT 285.660 197.620 285.940 197.900 ;
        RECT 286.060 197.620 286.340 197.900 ;
        RECT 286.460 197.620 286.740 197.900 ;
        RECT 286.860 197.620 287.140 197.900 ;
        RECT 287.260 197.620 287.540 197.900 ;
        RECT 4.640 178.820 4.920 179.100 ;
        RECT 5.040 178.820 5.320 179.100 ;
        RECT 5.440 178.820 5.720 179.100 ;
        RECT 5.840 178.820 6.120 179.100 ;
        RECT 6.240 178.820 6.520 179.100 ;
        RECT 6.640 178.820 6.920 179.100 ;
        RECT 7.040 178.820 7.320 179.100 ;
        RECT 7.440 178.820 7.720 179.100 ;
        RECT 7.840 178.820 8.120 179.100 ;
        RECT 8.240 178.820 8.520 179.100 ;
        RECT 8.640 178.820 8.920 179.100 ;
        RECT 9.040 178.820 9.320 179.100 ;
        RECT 9.440 178.820 9.720 179.100 ;
        RECT 9.840 178.820 10.120 179.100 ;
        RECT 10.240 178.820 10.520 179.100 ;
        RECT 10.640 178.820 10.920 179.100 ;
        RECT 11.040 178.820 11.320 179.100 ;
        RECT 11.440 178.820 11.720 179.100 ;
        RECT 11.840 178.820 12.120 179.100 ;
        RECT 12.240 178.820 12.520 179.100 ;
        RECT 279.660 178.820 279.940 179.100 ;
        RECT 280.060 178.820 280.340 179.100 ;
        RECT 280.460 178.820 280.740 179.100 ;
        RECT 280.860 178.820 281.140 179.100 ;
        RECT 281.260 178.820 281.540 179.100 ;
        RECT 281.660 178.820 281.940 179.100 ;
        RECT 282.060 178.820 282.340 179.100 ;
        RECT 282.460 178.820 282.740 179.100 ;
        RECT 282.860 178.820 283.140 179.100 ;
        RECT 283.260 178.820 283.540 179.100 ;
        RECT 283.660 178.820 283.940 179.100 ;
        RECT 284.060 178.820 284.340 179.100 ;
        RECT 284.460 178.820 284.740 179.100 ;
        RECT 284.860 178.820 285.140 179.100 ;
        RECT 285.260 178.820 285.540 179.100 ;
        RECT 285.660 178.820 285.940 179.100 ;
        RECT 286.060 178.820 286.340 179.100 ;
        RECT 286.460 178.820 286.740 179.100 ;
        RECT 286.860 178.820 287.140 179.100 ;
        RECT 287.260 178.820 287.540 179.100 ;
        RECT 4.640 160.020 4.920 160.300 ;
        RECT 5.040 160.020 5.320 160.300 ;
        RECT 5.440 160.020 5.720 160.300 ;
        RECT 5.840 160.020 6.120 160.300 ;
        RECT 6.240 160.020 6.520 160.300 ;
        RECT 6.640 160.020 6.920 160.300 ;
        RECT 7.040 160.020 7.320 160.300 ;
        RECT 7.440 160.020 7.720 160.300 ;
        RECT 7.840 160.020 8.120 160.300 ;
        RECT 8.240 160.020 8.520 160.300 ;
        RECT 8.640 160.020 8.920 160.300 ;
        RECT 9.040 160.020 9.320 160.300 ;
        RECT 9.440 160.020 9.720 160.300 ;
        RECT 9.840 160.020 10.120 160.300 ;
        RECT 10.240 160.020 10.520 160.300 ;
        RECT 10.640 160.020 10.920 160.300 ;
        RECT 11.040 160.020 11.320 160.300 ;
        RECT 11.440 160.020 11.720 160.300 ;
        RECT 11.840 160.020 12.120 160.300 ;
        RECT 12.240 160.020 12.520 160.300 ;
        RECT 279.660 160.020 279.940 160.300 ;
        RECT 280.060 160.020 280.340 160.300 ;
        RECT 280.460 160.020 280.740 160.300 ;
        RECT 280.860 160.020 281.140 160.300 ;
        RECT 281.260 160.020 281.540 160.300 ;
        RECT 281.660 160.020 281.940 160.300 ;
        RECT 282.060 160.020 282.340 160.300 ;
        RECT 282.460 160.020 282.740 160.300 ;
        RECT 282.860 160.020 283.140 160.300 ;
        RECT 283.260 160.020 283.540 160.300 ;
        RECT 283.660 160.020 283.940 160.300 ;
        RECT 284.060 160.020 284.340 160.300 ;
        RECT 284.460 160.020 284.740 160.300 ;
        RECT 284.860 160.020 285.140 160.300 ;
        RECT 285.260 160.020 285.540 160.300 ;
        RECT 285.660 160.020 285.940 160.300 ;
        RECT 286.060 160.020 286.340 160.300 ;
        RECT 286.460 160.020 286.740 160.300 ;
        RECT 286.860 160.020 287.140 160.300 ;
        RECT 287.260 160.020 287.540 160.300 ;
        RECT 4.640 141.220 4.920 141.500 ;
        RECT 5.040 141.220 5.320 141.500 ;
        RECT 5.440 141.220 5.720 141.500 ;
        RECT 5.840 141.220 6.120 141.500 ;
        RECT 6.240 141.220 6.520 141.500 ;
        RECT 6.640 141.220 6.920 141.500 ;
        RECT 7.040 141.220 7.320 141.500 ;
        RECT 7.440 141.220 7.720 141.500 ;
        RECT 7.840 141.220 8.120 141.500 ;
        RECT 8.240 141.220 8.520 141.500 ;
        RECT 8.640 141.220 8.920 141.500 ;
        RECT 9.040 141.220 9.320 141.500 ;
        RECT 9.440 141.220 9.720 141.500 ;
        RECT 9.840 141.220 10.120 141.500 ;
        RECT 10.240 141.220 10.520 141.500 ;
        RECT 10.640 141.220 10.920 141.500 ;
        RECT 11.040 141.220 11.320 141.500 ;
        RECT 11.440 141.220 11.720 141.500 ;
        RECT 11.840 141.220 12.120 141.500 ;
        RECT 12.240 141.220 12.520 141.500 ;
        RECT 279.660 141.220 279.940 141.500 ;
        RECT 280.060 141.220 280.340 141.500 ;
        RECT 280.460 141.220 280.740 141.500 ;
        RECT 280.860 141.220 281.140 141.500 ;
        RECT 281.260 141.220 281.540 141.500 ;
        RECT 281.660 141.220 281.940 141.500 ;
        RECT 282.060 141.220 282.340 141.500 ;
        RECT 282.460 141.220 282.740 141.500 ;
        RECT 282.860 141.220 283.140 141.500 ;
        RECT 283.260 141.220 283.540 141.500 ;
        RECT 283.660 141.220 283.940 141.500 ;
        RECT 284.060 141.220 284.340 141.500 ;
        RECT 284.460 141.220 284.740 141.500 ;
        RECT 284.860 141.220 285.140 141.500 ;
        RECT 285.260 141.220 285.540 141.500 ;
        RECT 285.660 141.220 285.940 141.500 ;
        RECT 286.060 141.220 286.340 141.500 ;
        RECT 286.460 141.220 286.740 141.500 ;
        RECT 286.860 141.220 287.140 141.500 ;
        RECT 287.260 141.220 287.540 141.500 ;
        RECT 4.640 122.420 4.920 122.700 ;
        RECT 5.040 122.420 5.320 122.700 ;
        RECT 5.440 122.420 5.720 122.700 ;
        RECT 5.840 122.420 6.120 122.700 ;
        RECT 6.240 122.420 6.520 122.700 ;
        RECT 6.640 122.420 6.920 122.700 ;
        RECT 7.040 122.420 7.320 122.700 ;
        RECT 7.440 122.420 7.720 122.700 ;
        RECT 7.840 122.420 8.120 122.700 ;
        RECT 8.240 122.420 8.520 122.700 ;
        RECT 8.640 122.420 8.920 122.700 ;
        RECT 9.040 122.420 9.320 122.700 ;
        RECT 9.440 122.420 9.720 122.700 ;
        RECT 9.840 122.420 10.120 122.700 ;
        RECT 10.240 122.420 10.520 122.700 ;
        RECT 10.640 122.420 10.920 122.700 ;
        RECT 11.040 122.420 11.320 122.700 ;
        RECT 11.440 122.420 11.720 122.700 ;
        RECT 11.840 122.420 12.120 122.700 ;
        RECT 12.240 122.420 12.520 122.700 ;
        RECT 279.660 122.420 279.940 122.700 ;
        RECT 280.060 122.420 280.340 122.700 ;
        RECT 280.460 122.420 280.740 122.700 ;
        RECT 280.860 122.420 281.140 122.700 ;
        RECT 281.260 122.420 281.540 122.700 ;
        RECT 281.660 122.420 281.940 122.700 ;
        RECT 282.060 122.420 282.340 122.700 ;
        RECT 282.460 122.420 282.740 122.700 ;
        RECT 282.860 122.420 283.140 122.700 ;
        RECT 283.260 122.420 283.540 122.700 ;
        RECT 283.660 122.420 283.940 122.700 ;
        RECT 284.060 122.420 284.340 122.700 ;
        RECT 284.460 122.420 284.740 122.700 ;
        RECT 284.860 122.420 285.140 122.700 ;
        RECT 285.260 122.420 285.540 122.700 ;
        RECT 285.660 122.420 285.940 122.700 ;
        RECT 286.060 122.420 286.340 122.700 ;
        RECT 286.460 122.420 286.740 122.700 ;
        RECT 286.860 122.420 287.140 122.700 ;
        RECT 287.260 122.420 287.540 122.700 ;
        RECT 4.640 103.620 4.920 103.900 ;
        RECT 5.040 103.620 5.320 103.900 ;
        RECT 5.440 103.620 5.720 103.900 ;
        RECT 5.840 103.620 6.120 103.900 ;
        RECT 6.240 103.620 6.520 103.900 ;
        RECT 6.640 103.620 6.920 103.900 ;
        RECT 7.040 103.620 7.320 103.900 ;
        RECT 7.440 103.620 7.720 103.900 ;
        RECT 7.840 103.620 8.120 103.900 ;
        RECT 8.240 103.620 8.520 103.900 ;
        RECT 8.640 103.620 8.920 103.900 ;
        RECT 9.040 103.620 9.320 103.900 ;
        RECT 9.440 103.620 9.720 103.900 ;
        RECT 9.840 103.620 10.120 103.900 ;
        RECT 10.240 103.620 10.520 103.900 ;
        RECT 10.640 103.620 10.920 103.900 ;
        RECT 11.040 103.620 11.320 103.900 ;
        RECT 11.440 103.620 11.720 103.900 ;
        RECT 11.840 103.620 12.120 103.900 ;
        RECT 12.240 103.620 12.520 103.900 ;
        RECT 279.660 103.620 279.940 103.900 ;
        RECT 280.060 103.620 280.340 103.900 ;
        RECT 280.460 103.620 280.740 103.900 ;
        RECT 280.860 103.620 281.140 103.900 ;
        RECT 281.260 103.620 281.540 103.900 ;
        RECT 281.660 103.620 281.940 103.900 ;
        RECT 282.060 103.620 282.340 103.900 ;
        RECT 282.460 103.620 282.740 103.900 ;
        RECT 282.860 103.620 283.140 103.900 ;
        RECT 283.260 103.620 283.540 103.900 ;
        RECT 283.660 103.620 283.940 103.900 ;
        RECT 284.060 103.620 284.340 103.900 ;
        RECT 284.460 103.620 284.740 103.900 ;
        RECT 284.860 103.620 285.140 103.900 ;
        RECT 285.260 103.620 285.540 103.900 ;
        RECT 285.660 103.620 285.940 103.900 ;
        RECT 286.060 103.620 286.340 103.900 ;
        RECT 286.460 103.620 286.740 103.900 ;
        RECT 286.860 103.620 287.140 103.900 ;
        RECT 287.260 103.620 287.540 103.900 ;
        RECT 4.640 84.820 4.920 85.100 ;
        RECT 5.040 84.820 5.320 85.100 ;
        RECT 5.440 84.820 5.720 85.100 ;
        RECT 5.840 84.820 6.120 85.100 ;
        RECT 6.240 84.820 6.520 85.100 ;
        RECT 6.640 84.820 6.920 85.100 ;
        RECT 7.040 84.820 7.320 85.100 ;
        RECT 7.440 84.820 7.720 85.100 ;
        RECT 7.840 84.820 8.120 85.100 ;
        RECT 8.240 84.820 8.520 85.100 ;
        RECT 8.640 84.820 8.920 85.100 ;
        RECT 9.040 84.820 9.320 85.100 ;
        RECT 9.440 84.820 9.720 85.100 ;
        RECT 9.840 84.820 10.120 85.100 ;
        RECT 10.240 84.820 10.520 85.100 ;
        RECT 10.640 84.820 10.920 85.100 ;
        RECT 11.040 84.820 11.320 85.100 ;
        RECT 11.440 84.820 11.720 85.100 ;
        RECT 11.840 84.820 12.120 85.100 ;
        RECT 12.240 84.820 12.520 85.100 ;
        RECT 279.660 84.820 279.940 85.100 ;
        RECT 280.060 84.820 280.340 85.100 ;
        RECT 280.460 84.820 280.740 85.100 ;
        RECT 280.860 84.820 281.140 85.100 ;
        RECT 281.260 84.820 281.540 85.100 ;
        RECT 281.660 84.820 281.940 85.100 ;
        RECT 282.060 84.820 282.340 85.100 ;
        RECT 282.460 84.820 282.740 85.100 ;
        RECT 282.860 84.820 283.140 85.100 ;
        RECT 283.260 84.820 283.540 85.100 ;
        RECT 283.660 84.820 283.940 85.100 ;
        RECT 284.060 84.820 284.340 85.100 ;
        RECT 284.460 84.820 284.740 85.100 ;
        RECT 284.860 84.820 285.140 85.100 ;
        RECT 285.260 84.820 285.540 85.100 ;
        RECT 285.660 84.820 285.940 85.100 ;
        RECT 286.060 84.820 286.340 85.100 ;
        RECT 286.460 84.820 286.740 85.100 ;
        RECT 286.860 84.820 287.140 85.100 ;
        RECT 287.260 84.820 287.540 85.100 ;
        RECT 4.640 66.020 4.920 66.300 ;
        RECT 5.040 66.020 5.320 66.300 ;
        RECT 5.440 66.020 5.720 66.300 ;
        RECT 5.840 66.020 6.120 66.300 ;
        RECT 6.240 66.020 6.520 66.300 ;
        RECT 6.640 66.020 6.920 66.300 ;
        RECT 7.040 66.020 7.320 66.300 ;
        RECT 7.440 66.020 7.720 66.300 ;
        RECT 7.840 66.020 8.120 66.300 ;
        RECT 8.240 66.020 8.520 66.300 ;
        RECT 8.640 66.020 8.920 66.300 ;
        RECT 9.040 66.020 9.320 66.300 ;
        RECT 9.440 66.020 9.720 66.300 ;
        RECT 9.840 66.020 10.120 66.300 ;
        RECT 10.240 66.020 10.520 66.300 ;
        RECT 10.640 66.020 10.920 66.300 ;
        RECT 11.040 66.020 11.320 66.300 ;
        RECT 11.440 66.020 11.720 66.300 ;
        RECT 11.840 66.020 12.120 66.300 ;
        RECT 12.240 66.020 12.520 66.300 ;
        RECT 279.660 66.020 279.940 66.300 ;
        RECT 280.060 66.020 280.340 66.300 ;
        RECT 280.460 66.020 280.740 66.300 ;
        RECT 280.860 66.020 281.140 66.300 ;
        RECT 281.260 66.020 281.540 66.300 ;
        RECT 281.660 66.020 281.940 66.300 ;
        RECT 282.060 66.020 282.340 66.300 ;
        RECT 282.460 66.020 282.740 66.300 ;
        RECT 282.860 66.020 283.140 66.300 ;
        RECT 283.260 66.020 283.540 66.300 ;
        RECT 283.660 66.020 283.940 66.300 ;
        RECT 284.060 66.020 284.340 66.300 ;
        RECT 284.460 66.020 284.740 66.300 ;
        RECT 284.860 66.020 285.140 66.300 ;
        RECT 285.260 66.020 285.540 66.300 ;
        RECT 285.660 66.020 285.940 66.300 ;
        RECT 286.060 66.020 286.340 66.300 ;
        RECT 286.460 66.020 286.740 66.300 ;
        RECT 286.860 66.020 287.140 66.300 ;
        RECT 287.260 66.020 287.540 66.300 ;
        RECT 4.640 47.220 4.920 47.500 ;
        RECT 5.040 47.220 5.320 47.500 ;
        RECT 5.440 47.220 5.720 47.500 ;
        RECT 5.840 47.220 6.120 47.500 ;
        RECT 6.240 47.220 6.520 47.500 ;
        RECT 6.640 47.220 6.920 47.500 ;
        RECT 7.040 47.220 7.320 47.500 ;
        RECT 7.440 47.220 7.720 47.500 ;
        RECT 7.840 47.220 8.120 47.500 ;
        RECT 8.240 47.220 8.520 47.500 ;
        RECT 8.640 47.220 8.920 47.500 ;
        RECT 9.040 47.220 9.320 47.500 ;
        RECT 9.440 47.220 9.720 47.500 ;
        RECT 9.840 47.220 10.120 47.500 ;
        RECT 10.240 47.220 10.520 47.500 ;
        RECT 10.640 47.220 10.920 47.500 ;
        RECT 11.040 47.220 11.320 47.500 ;
        RECT 11.440 47.220 11.720 47.500 ;
        RECT 11.840 47.220 12.120 47.500 ;
        RECT 12.240 47.220 12.520 47.500 ;
        RECT 279.660 47.220 279.940 47.500 ;
        RECT 280.060 47.220 280.340 47.500 ;
        RECT 280.460 47.220 280.740 47.500 ;
        RECT 280.860 47.220 281.140 47.500 ;
        RECT 281.260 47.220 281.540 47.500 ;
        RECT 281.660 47.220 281.940 47.500 ;
        RECT 282.060 47.220 282.340 47.500 ;
        RECT 282.460 47.220 282.740 47.500 ;
        RECT 282.860 47.220 283.140 47.500 ;
        RECT 283.260 47.220 283.540 47.500 ;
        RECT 283.660 47.220 283.940 47.500 ;
        RECT 284.060 47.220 284.340 47.500 ;
        RECT 284.460 47.220 284.740 47.500 ;
        RECT 284.860 47.220 285.140 47.500 ;
        RECT 285.260 47.220 285.540 47.500 ;
        RECT 285.660 47.220 285.940 47.500 ;
        RECT 286.060 47.220 286.340 47.500 ;
        RECT 286.460 47.220 286.740 47.500 ;
        RECT 286.860 47.220 287.140 47.500 ;
        RECT 287.260 47.220 287.540 47.500 ;
        RECT 4.640 28.420 4.920 28.700 ;
        RECT 5.040 28.420 5.320 28.700 ;
        RECT 5.440 28.420 5.720 28.700 ;
        RECT 5.840 28.420 6.120 28.700 ;
        RECT 6.240 28.420 6.520 28.700 ;
        RECT 6.640 28.420 6.920 28.700 ;
        RECT 7.040 28.420 7.320 28.700 ;
        RECT 7.440 28.420 7.720 28.700 ;
        RECT 7.840 28.420 8.120 28.700 ;
        RECT 8.240 28.420 8.520 28.700 ;
        RECT 8.640 28.420 8.920 28.700 ;
        RECT 9.040 28.420 9.320 28.700 ;
        RECT 9.440 28.420 9.720 28.700 ;
        RECT 9.840 28.420 10.120 28.700 ;
        RECT 10.240 28.420 10.520 28.700 ;
        RECT 10.640 28.420 10.920 28.700 ;
        RECT 11.040 28.420 11.320 28.700 ;
        RECT 11.440 28.420 11.720 28.700 ;
        RECT 11.840 28.420 12.120 28.700 ;
        RECT 12.240 28.420 12.520 28.700 ;
        RECT 279.660 28.420 279.940 28.700 ;
        RECT 280.060 28.420 280.340 28.700 ;
        RECT 280.460 28.420 280.740 28.700 ;
        RECT 280.860 28.420 281.140 28.700 ;
        RECT 281.260 28.420 281.540 28.700 ;
        RECT 281.660 28.420 281.940 28.700 ;
        RECT 282.060 28.420 282.340 28.700 ;
        RECT 282.460 28.420 282.740 28.700 ;
        RECT 282.860 28.420 283.140 28.700 ;
        RECT 283.260 28.420 283.540 28.700 ;
        RECT 283.660 28.420 283.940 28.700 ;
        RECT 284.060 28.420 284.340 28.700 ;
        RECT 284.460 28.420 284.740 28.700 ;
        RECT 284.860 28.420 285.140 28.700 ;
        RECT 285.260 28.420 285.540 28.700 ;
        RECT 285.660 28.420 285.940 28.700 ;
        RECT 286.060 28.420 286.340 28.700 ;
        RECT 286.460 28.420 286.740 28.700 ;
        RECT 286.860 28.420 287.140 28.700 ;
        RECT 287.260 28.420 287.540 28.700 ;
      LAYER met3 ;
        RECT 4.500 253.860 12.660 254.460 ;
        RECT 279.520 253.860 287.680 254.460 ;
        RECT 29.590 236.010 30.590 236.610 ;
        RECT 66.830 236.010 67.830 236.610 ;
        RECT 88.385 235.680 88.715 235.685 ;
        RECT 88.360 235.670 88.740 235.680 ;
        RECT 4.500 235.060 12.660 235.660 ;
        RECT 87.940 235.370 88.740 235.670 ;
        RECT 88.360 235.360 88.740 235.370 ;
        RECT 88.385 235.355 88.715 235.360 ;
        RECT 279.520 235.060 287.680 235.660 ;
        RECT 29.590 217.210 30.590 217.810 ;
        RECT 4.500 216.260 12.660 216.860 ;
        RECT 41.465 216.770 41.795 216.775 ;
        RECT 41.440 216.760 41.820 216.770 ;
        RECT 41.440 216.460 42.240 216.760 ;
        RECT 41.440 216.450 41.820 216.460 ;
        RECT 41.465 216.445 41.795 216.450 ;
        RECT 279.520 216.260 287.680 216.860 ;
        RECT 31.550 198.410 32.550 199.010 ;
        RECT 75.650 198.410 76.650 199.010 ;
        RECT 77.345 198.470 77.675 198.475 ;
        RECT 77.320 198.460 77.700 198.470 ;
        RECT 77.320 198.160 78.120 198.460 ;
        RECT 77.320 198.150 77.700 198.160 ;
        RECT 77.345 198.145 77.675 198.150 ;
        RECT 4.500 197.460 12.660 198.060 ;
        RECT 279.520 197.460 287.680 198.060 ;
        RECT 4.500 178.660 12.660 179.260 ;
        RECT 279.520 178.660 287.680 179.260 ;
        RECT 4.500 159.860 12.660 160.460 ;
        RECT 279.520 159.860 287.680 160.460 ;
        RECT 4.500 141.060 12.660 141.660 ;
        RECT 279.520 141.060 287.680 141.660 ;
        RECT 4.500 122.260 12.660 122.860 ;
        RECT 279.520 122.260 287.680 122.860 ;
        RECT 4.500 103.460 12.660 104.060 ;
        RECT 279.520 103.460 287.680 104.060 ;
        RECT 4.500 84.660 12.660 85.260 ;
        RECT 279.520 84.660 287.680 85.260 ;
        RECT 4.500 65.860 12.660 66.460 ;
        RECT 279.520 65.860 287.680 66.460 ;
        RECT 4.500 47.060 12.660 47.660 ;
        RECT 279.520 47.060 287.680 47.660 ;
        RECT 4.500 28.260 12.660 28.860 ;
        RECT 279.520 28.260 287.680 28.860 ;
      LAYER via3 ;
        RECT 4.620 254.000 4.940 254.320 ;
        RECT 5.020 254.000 5.340 254.320 ;
        RECT 5.420 254.000 5.740 254.320 ;
        RECT 5.820 254.000 6.140 254.320 ;
        RECT 6.220 254.000 6.540 254.320 ;
        RECT 6.620 254.000 6.940 254.320 ;
        RECT 7.020 254.000 7.340 254.320 ;
        RECT 7.420 254.000 7.740 254.320 ;
        RECT 7.820 254.000 8.140 254.320 ;
        RECT 8.220 254.000 8.540 254.320 ;
        RECT 8.620 254.000 8.940 254.320 ;
        RECT 9.020 254.000 9.340 254.320 ;
        RECT 9.420 254.000 9.740 254.320 ;
        RECT 9.820 254.000 10.140 254.320 ;
        RECT 10.220 254.000 10.540 254.320 ;
        RECT 10.620 254.000 10.940 254.320 ;
        RECT 11.020 254.000 11.340 254.320 ;
        RECT 11.420 254.000 11.740 254.320 ;
        RECT 11.820 254.000 12.140 254.320 ;
        RECT 12.220 254.000 12.540 254.320 ;
        RECT 279.640 254.000 279.960 254.320 ;
        RECT 280.040 254.000 280.360 254.320 ;
        RECT 280.440 254.000 280.760 254.320 ;
        RECT 280.840 254.000 281.160 254.320 ;
        RECT 281.240 254.000 281.560 254.320 ;
        RECT 281.640 254.000 281.960 254.320 ;
        RECT 282.040 254.000 282.360 254.320 ;
        RECT 282.440 254.000 282.760 254.320 ;
        RECT 282.840 254.000 283.160 254.320 ;
        RECT 283.240 254.000 283.560 254.320 ;
        RECT 283.640 254.000 283.960 254.320 ;
        RECT 284.040 254.000 284.360 254.320 ;
        RECT 284.440 254.000 284.760 254.320 ;
        RECT 284.840 254.000 285.160 254.320 ;
        RECT 285.240 254.000 285.560 254.320 ;
        RECT 285.640 254.000 285.960 254.320 ;
        RECT 286.040 254.000 286.360 254.320 ;
        RECT 286.440 254.000 286.760 254.320 ;
        RECT 286.840 254.000 287.160 254.320 ;
        RECT 287.240 254.000 287.560 254.320 ;
        RECT 29.730 236.150 30.050 236.470 ;
        RECT 30.130 236.150 30.450 236.470 ;
        RECT 66.970 236.150 67.290 236.470 ;
        RECT 67.370 236.150 67.690 236.470 ;
        RECT 4.620 235.200 4.940 235.520 ;
        RECT 5.020 235.200 5.340 235.520 ;
        RECT 5.420 235.200 5.740 235.520 ;
        RECT 5.820 235.200 6.140 235.520 ;
        RECT 6.220 235.200 6.540 235.520 ;
        RECT 6.620 235.200 6.940 235.520 ;
        RECT 7.020 235.200 7.340 235.520 ;
        RECT 7.420 235.200 7.740 235.520 ;
        RECT 7.820 235.200 8.140 235.520 ;
        RECT 8.220 235.200 8.540 235.520 ;
        RECT 8.620 235.200 8.940 235.520 ;
        RECT 9.020 235.200 9.340 235.520 ;
        RECT 9.420 235.200 9.740 235.520 ;
        RECT 9.820 235.200 10.140 235.520 ;
        RECT 10.220 235.200 10.540 235.520 ;
        RECT 10.620 235.200 10.940 235.520 ;
        RECT 11.020 235.200 11.340 235.520 ;
        RECT 11.420 235.200 11.740 235.520 ;
        RECT 11.820 235.200 12.140 235.520 ;
        RECT 12.220 235.200 12.540 235.520 ;
        RECT 88.390 235.360 88.710 235.680 ;
        RECT 279.640 235.200 279.960 235.520 ;
        RECT 280.040 235.200 280.360 235.520 ;
        RECT 280.440 235.200 280.760 235.520 ;
        RECT 280.840 235.200 281.160 235.520 ;
        RECT 281.240 235.200 281.560 235.520 ;
        RECT 281.640 235.200 281.960 235.520 ;
        RECT 282.040 235.200 282.360 235.520 ;
        RECT 282.440 235.200 282.760 235.520 ;
        RECT 282.840 235.200 283.160 235.520 ;
        RECT 283.240 235.200 283.560 235.520 ;
        RECT 283.640 235.200 283.960 235.520 ;
        RECT 284.040 235.200 284.360 235.520 ;
        RECT 284.440 235.200 284.760 235.520 ;
        RECT 284.840 235.200 285.160 235.520 ;
        RECT 285.240 235.200 285.560 235.520 ;
        RECT 285.640 235.200 285.960 235.520 ;
        RECT 286.040 235.200 286.360 235.520 ;
        RECT 286.440 235.200 286.760 235.520 ;
        RECT 286.840 235.200 287.160 235.520 ;
        RECT 287.240 235.200 287.560 235.520 ;
        RECT 29.730 217.350 30.050 217.670 ;
        RECT 30.130 217.350 30.450 217.670 ;
        RECT 4.620 216.400 4.940 216.720 ;
        RECT 5.020 216.400 5.340 216.720 ;
        RECT 5.420 216.400 5.740 216.720 ;
        RECT 5.820 216.400 6.140 216.720 ;
        RECT 6.220 216.400 6.540 216.720 ;
        RECT 6.620 216.400 6.940 216.720 ;
        RECT 7.020 216.400 7.340 216.720 ;
        RECT 7.420 216.400 7.740 216.720 ;
        RECT 7.820 216.400 8.140 216.720 ;
        RECT 8.220 216.400 8.540 216.720 ;
        RECT 8.620 216.400 8.940 216.720 ;
        RECT 9.020 216.400 9.340 216.720 ;
        RECT 9.420 216.400 9.740 216.720 ;
        RECT 9.820 216.400 10.140 216.720 ;
        RECT 10.220 216.400 10.540 216.720 ;
        RECT 10.620 216.400 10.940 216.720 ;
        RECT 11.020 216.400 11.340 216.720 ;
        RECT 11.420 216.400 11.740 216.720 ;
        RECT 11.820 216.400 12.140 216.720 ;
        RECT 12.220 216.400 12.540 216.720 ;
        RECT 41.470 216.450 41.790 216.770 ;
        RECT 279.640 216.400 279.960 216.720 ;
        RECT 280.040 216.400 280.360 216.720 ;
        RECT 280.440 216.400 280.760 216.720 ;
        RECT 280.840 216.400 281.160 216.720 ;
        RECT 281.240 216.400 281.560 216.720 ;
        RECT 281.640 216.400 281.960 216.720 ;
        RECT 282.040 216.400 282.360 216.720 ;
        RECT 282.440 216.400 282.760 216.720 ;
        RECT 282.840 216.400 283.160 216.720 ;
        RECT 283.240 216.400 283.560 216.720 ;
        RECT 283.640 216.400 283.960 216.720 ;
        RECT 284.040 216.400 284.360 216.720 ;
        RECT 284.440 216.400 284.760 216.720 ;
        RECT 284.840 216.400 285.160 216.720 ;
        RECT 285.240 216.400 285.560 216.720 ;
        RECT 285.640 216.400 285.960 216.720 ;
        RECT 286.040 216.400 286.360 216.720 ;
        RECT 286.440 216.400 286.760 216.720 ;
        RECT 286.840 216.400 287.160 216.720 ;
        RECT 287.240 216.400 287.560 216.720 ;
        RECT 31.690 198.550 32.010 198.870 ;
        RECT 32.090 198.550 32.410 198.870 ;
        RECT 75.790 198.550 76.110 198.870 ;
        RECT 76.190 198.550 76.510 198.870 ;
        RECT 77.350 198.150 77.670 198.470 ;
        RECT 4.620 197.600 4.940 197.920 ;
        RECT 5.020 197.600 5.340 197.920 ;
        RECT 5.420 197.600 5.740 197.920 ;
        RECT 5.820 197.600 6.140 197.920 ;
        RECT 6.220 197.600 6.540 197.920 ;
        RECT 6.620 197.600 6.940 197.920 ;
        RECT 7.020 197.600 7.340 197.920 ;
        RECT 7.420 197.600 7.740 197.920 ;
        RECT 7.820 197.600 8.140 197.920 ;
        RECT 8.220 197.600 8.540 197.920 ;
        RECT 8.620 197.600 8.940 197.920 ;
        RECT 9.020 197.600 9.340 197.920 ;
        RECT 9.420 197.600 9.740 197.920 ;
        RECT 9.820 197.600 10.140 197.920 ;
        RECT 10.220 197.600 10.540 197.920 ;
        RECT 10.620 197.600 10.940 197.920 ;
        RECT 11.020 197.600 11.340 197.920 ;
        RECT 11.420 197.600 11.740 197.920 ;
        RECT 11.820 197.600 12.140 197.920 ;
        RECT 12.220 197.600 12.540 197.920 ;
        RECT 279.640 197.600 279.960 197.920 ;
        RECT 280.040 197.600 280.360 197.920 ;
        RECT 280.440 197.600 280.760 197.920 ;
        RECT 280.840 197.600 281.160 197.920 ;
        RECT 281.240 197.600 281.560 197.920 ;
        RECT 281.640 197.600 281.960 197.920 ;
        RECT 282.040 197.600 282.360 197.920 ;
        RECT 282.440 197.600 282.760 197.920 ;
        RECT 282.840 197.600 283.160 197.920 ;
        RECT 283.240 197.600 283.560 197.920 ;
        RECT 283.640 197.600 283.960 197.920 ;
        RECT 284.040 197.600 284.360 197.920 ;
        RECT 284.440 197.600 284.760 197.920 ;
        RECT 284.840 197.600 285.160 197.920 ;
        RECT 285.240 197.600 285.560 197.920 ;
        RECT 285.640 197.600 285.960 197.920 ;
        RECT 286.040 197.600 286.360 197.920 ;
        RECT 286.440 197.600 286.760 197.920 ;
        RECT 286.840 197.600 287.160 197.920 ;
        RECT 287.240 197.600 287.560 197.920 ;
        RECT 4.620 178.800 4.940 179.120 ;
        RECT 5.020 178.800 5.340 179.120 ;
        RECT 5.420 178.800 5.740 179.120 ;
        RECT 5.820 178.800 6.140 179.120 ;
        RECT 6.220 178.800 6.540 179.120 ;
        RECT 6.620 178.800 6.940 179.120 ;
        RECT 7.020 178.800 7.340 179.120 ;
        RECT 7.420 178.800 7.740 179.120 ;
        RECT 7.820 178.800 8.140 179.120 ;
        RECT 8.220 178.800 8.540 179.120 ;
        RECT 8.620 178.800 8.940 179.120 ;
        RECT 9.020 178.800 9.340 179.120 ;
        RECT 9.420 178.800 9.740 179.120 ;
        RECT 9.820 178.800 10.140 179.120 ;
        RECT 10.220 178.800 10.540 179.120 ;
        RECT 10.620 178.800 10.940 179.120 ;
        RECT 11.020 178.800 11.340 179.120 ;
        RECT 11.420 178.800 11.740 179.120 ;
        RECT 11.820 178.800 12.140 179.120 ;
        RECT 12.220 178.800 12.540 179.120 ;
        RECT 279.640 178.800 279.960 179.120 ;
        RECT 280.040 178.800 280.360 179.120 ;
        RECT 280.440 178.800 280.760 179.120 ;
        RECT 280.840 178.800 281.160 179.120 ;
        RECT 281.240 178.800 281.560 179.120 ;
        RECT 281.640 178.800 281.960 179.120 ;
        RECT 282.040 178.800 282.360 179.120 ;
        RECT 282.440 178.800 282.760 179.120 ;
        RECT 282.840 178.800 283.160 179.120 ;
        RECT 283.240 178.800 283.560 179.120 ;
        RECT 283.640 178.800 283.960 179.120 ;
        RECT 284.040 178.800 284.360 179.120 ;
        RECT 284.440 178.800 284.760 179.120 ;
        RECT 284.840 178.800 285.160 179.120 ;
        RECT 285.240 178.800 285.560 179.120 ;
        RECT 285.640 178.800 285.960 179.120 ;
        RECT 286.040 178.800 286.360 179.120 ;
        RECT 286.440 178.800 286.760 179.120 ;
        RECT 286.840 178.800 287.160 179.120 ;
        RECT 287.240 178.800 287.560 179.120 ;
        RECT 4.620 160.000 4.940 160.320 ;
        RECT 5.020 160.000 5.340 160.320 ;
        RECT 5.420 160.000 5.740 160.320 ;
        RECT 5.820 160.000 6.140 160.320 ;
        RECT 6.220 160.000 6.540 160.320 ;
        RECT 6.620 160.000 6.940 160.320 ;
        RECT 7.020 160.000 7.340 160.320 ;
        RECT 7.420 160.000 7.740 160.320 ;
        RECT 7.820 160.000 8.140 160.320 ;
        RECT 8.220 160.000 8.540 160.320 ;
        RECT 8.620 160.000 8.940 160.320 ;
        RECT 9.020 160.000 9.340 160.320 ;
        RECT 9.420 160.000 9.740 160.320 ;
        RECT 9.820 160.000 10.140 160.320 ;
        RECT 10.220 160.000 10.540 160.320 ;
        RECT 10.620 160.000 10.940 160.320 ;
        RECT 11.020 160.000 11.340 160.320 ;
        RECT 11.420 160.000 11.740 160.320 ;
        RECT 11.820 160.000 12.140 160.320 ;
        RECT 12.220 160.000 12.540 160.320 ;
        RECT 279.640 160.000 279.960 160.320 ;
        RECT 280.040 160.000 280.360 160.320 ;
        RECT 280.440 160.000 280.760 160.320 ;
        RECT 280.840 160.000 281.160 160.320 ;
        RECT 281.240 160.000 281.560 160.320 ;
        RECT 281.640 160.000 281.960 160.320 ;
        RECT 282.040 160.000 282.360 160.320 ;
        RECT 282.440 160.000 282.760 160.320 ;
        RECT 282.840 160.000 283.160 160.320 ;
        RECT 283.240 160.000 283.560 160.320 ;
        RECT 283.640 160.000 283.960 160.320 ;
        RECT 284.040 160.000 284.360 160.320 ;
        RECT 284.440 160.000 284.760 160.320 ;
        RECT 284.840 160.000 285.160 160.320 ;
        RECT 285.240 160.000 285.560 160.320 ;
        RECT 285.640 160.000 285.960 160.320 ;
        RECT 286.040 160.000 286.360 160.320 ;
        RECT 286.440 160.000 286.760 160.320 ;
        RECT 286.840 160.000 287.160 160.320 ;
        RECT 287.240 160.000 287.560 160.320 ;
        RECT 4.620 141.200 4.940 141.520 ;
        RECT 5.020 141.200 5.340 141.520 ;
        RECT 5.420 141.200 5.740 141.520 ;
        RECT 5.820 141.200 6.140 141.520 ;
        RECT 6.220 141.200 6.540 141.520 ;
        RECT 6.620 141.200 6.940 141.520 ;
        RECT 7.020 141.200 7.340 141.520 ;
        RECT 7.420 141.200 7.740 141.520 ;
        RECT 7.820 141.200 8.140 141.520 ;
        RECT 8.220 141.200 8.540 141.520 ;
        RECT 8.620 141.200 8.940 141.520 ;
        RECT 9.020 141.200 9.340 141.520 ;
        RECT 9.420 141.200 9.740 141.520 ;
        RECT 9.820 141.200 10.140 141.520 ;
        RECT 10.220 141.200 10.540 141.520 ;
        RECT 10.620 141.200 10.940 141.520 ;
        RECT 11.020 141.200 11.340 141.520 ;
        RECT 11.420 141.200 11.740 141.520 ;
        RECT 11.820 141.200 12.140 141.520 ;
        RECT 12.220 141.200 12.540 141.520 ;
        RECT 279.640 141.200 279.960 141.520 ;
        RECT 280.040 141.200 280.360 141.520 ;
        RECT 280.440 141.200 280.760 141.520 ;
        RECT 280.840 141.200 281.160 141.520 ;
        RECT 281.240 141.200 281.560 141.520 ;
        RECT 281.640 141.200 281.960 141.520 ;
        RECT 282.040 141.200 282.360 141.520 ;
        RECT 282.440 141.200 282.760 141.520 ;
        RECT 282.840 141.200 283.160 141.520 ;
        RECT 283.240 141.200 283.560 141.520 ;
        RECT 283.640 141.200 283.960 141.520 ;
        RECT 284.040 141.200 284.360 141.520 ;
        RECT 284.440 141.200 284.760 141.520 ;
        RECT 284.840 141.200 285.160 141.520 ;
        RECT 285.240 141.200 285.560 141.520 ;
        RECT 285.640 141.200 285.960 141.520 ;
        RECT 286.040 141.200 286.360 141.520 ;
        RECT 286.440 141.200 286.760 141.520 ;
        RECT 286.840 141.200 287.160 141.520 ;
        RECT 287.240 141.200 287.560 141.520 ;
        RECT 4.620 122.400 4.940 122.720 ;
        RECT 5.020 122.400 5.340 122.720 ;
        RECT 5.420 122.400 5.740 122.720 ;
        RECT 5.820 122.400 6.140 122.720 ;
        RECT 6.220 122.400 6.540 122.720 ;
        RECT 6.620 122.400 6.940 122.720 ;
        RECT 7.020 122.400 7.340 122.720 ;
        RECT 7.420 122.400 7.740 122.720 ;
        RECT 7.820 122.400 8.140 122.720 ;
        RECT 8.220 122.400 8.540 122.720 ;
        RECT 8.620 122.400 8.940 122.720 ;
        RECT 9.020 122.400 9.340 122.720 ;
        RECT 9.420 122.400 9.740 122.720 ;
        RECT 9.820 122.400 10.140 122.720 ;
        RECT 10.220 122.400 10.540 122.720 ;
        RECT 10.620 122.400 10.940 122.720 ;
        RECT 11.020 122.400 11.340 122.720 ;
        RECT 11.420 122.400 11.740 122.720 ;
        RECT 11.820 122.400 12.140 122.720 ;
        RECT 12.220 122.400 12.540 122.720 ;
        RECT 279.640 122.400 279.960 122.720 ;
        RECT 280.040 122.400 280.360 122.720 ;
        RECT 280.440 122.400 280.760 122.720 ;
        RECT 280.840 122.400 281.160 122.720 ;
        RECT 281.240 122.400 281.560 122.720 ;
        RECT 281.640 122.400 281.960 122.720 ;
        RECT 282.040 122.400 282.360 122.720 ;
        RECT 282.440 122.400 282.760 122.720 ;
        RECT 282.840 122.400 283.160 122.720 ;
        RECT 283.240 122.400 283.560 122.720 ;
        RECT 283.640 122.400 283.960 122.720 ;
        RECT 284.040 122.400 284.360 122.720 ;
        RECT 284.440 122.400 284.760 122.720 ;
        RECT 284.840 122.400 285.160 122.720 ;
        RECT 285.240 122.400 285.560 122.720 ;
        RECT 285.640 122.400 285.960 122.720 ;
        RECT 286.040 122.400 286.360 122.720 ;
        RECT 286.440 122.400 286.760 122.720 ;
        RECT 286.840 122.400 287.160 122.720 ;
        RECT 287.240 122.400 287.560 122.720 ;
        RECT 4.620 103.600 4.940 103.920 ;
        RECT 5.020 103.600 5.340 103.920 ;
        RECT 5.420 103.600 5.740 103.920 ;
        RECT 5.820 103.600 6.140 103.920 ;
        RECT 6.220 103.600 6.540 103.920 ;
        RECT 6.620 103.600 6.940 103.920 ;
        RECT 7.020 103.600 7.340 103.920 ;
        RECT 7.420 103.600 7.740 103.920 ;
        RECT 7.820 103.600 8.140 103.920 ;
        RECT 8.220 103.600 8.540 103.920 ;
        RECT 8.620 103.600 8.940 103.920 ;
        RECT 9.020 103.600 9.340 103.920 ;
        RECT 9.420 103.600 9.740 103.920 ;
        RECT 9.820 103.600 10.140 103.920 ;
        RECT 10.220 103.600 10.540 103.920 ;
        RECT 10.620 103.600 10.940 103.920 ;
        RECT 11.020 103.600 11.340 103.920 ;
        RECT 11.420 103.600 11.740 103.920 ;
        RECT 11.820 103.600 12.140 103.920 ;
        RECT 12.220 103.600 12.540 103.920 ;
        RECT 279.640 103.600 279.960 103.920 ;
        RECT 280.040 103.600 280.360 103.920 ;
        RECT 280.440 103.600 280.760 103.920 ;
        RECT 280.840 103.600 281.160 103.920 ;
        RECT 281.240 103.600 281.560 103.920 ;
        RECT 281.640 103.600 281.960 103.920 ;
        RECT 282.040 103.600 282.360 103.920 ;
        RECT 282.440 103.600 282.760 103.920 ;
        RECT 282.840 103.600 283.160 103.920 ;
        RECT 283.240 103.600 283.560 103.920 ;
        RECT 283.640 103.600 283.960 103.920 ;
        RECT 284.040 103.600 284.360 103.920 ;
        RECT 284.440 103.600 284.760 103.920 ;
        RECT 284.840 103.600 285.160 103.920 ;
        RECT 285.240 103.600 285.560 103.920 ;
        RECT 285.640 103.600 285.960 103.920 ;
        RECT 286.040 103.600 286.360 103.920 ;
        RECT 286.440 103.600 286.760 103.920 ;
        RECT 286.840 103.600 287.160 103.920 ;
        RECT 287.240 103.600 287.560 103.920 ;
        RECT 4.620 84.800 4.940 85.120 ;
        RECT 5.020 84.800 5.340 85.120 ;
        RECT 5.420 84.800 5.740 85.120 ;
        RECT 5.820 84.800 6.140 85.120 ;
        RECT 6.220 84.800 6.540 85.120 ;
        RECT 6.620 84.800 6.940 85.120 ;
        RECT 7.020 84.800 7.340 85.120 ;
        RECT 7.420 84.800 7.740 85.120 ;
        RECT 7.820 84.800 8.140 85.120 ;
        RECT 8.220 84.800 8.540 85.120 ;
        RECT 8.620 84.800 8.940 85.120 ;
        RECT 9.020 84.800 9.340 85.120 ;
        RECT 9.420 84.800 9.740 85.120 ;
        RECT 9.820 84.800 10.140 85.120 ;
        RECT 10.220 84.800 10.540 85.120 ;
        RECT 10.620 84.800 10.940 85.120 ;
        RECT 11.020 84.800 11.340 85.120 ;
        RECT 11.420 84.800 11.740 85.120 ;
        RECT 11.820 84.800 12.140 85.120 ;
        RECT 12.220 84.800 12.540 85.120 ;
        RECT 279.640 84.800 279.960 85.120 ;
        RECT 280.040 84.800 280.360 85.120 ;
        RECT 280.440 84.800 280.760 85.120 ;
        RECT 280.840 84.800 281.160 85.120 ;
        RECT 281.240 84.800 281.560 85.120 ;
        RECT 281.640 84.800 281.960 85.120 ;
        RECT 282.040 84.800 282.360 85.120 ;
        RECT 282.440 84.800 282.760 85.120 ;
        RECT 282.840 84.800 283.160 85.120 ;
        RECT 283.240 84.800 283.560 85.120 ;
        RECT 283.640 84.800 283.960 85.120 ;
        RECT 284.040 84.800 284.360 85.120 ;
        RECT 284.440 84.800 284.760 85.120 ;
        RECT 284.840 84.800 285.160 85.120 ;
        RECT 285.240 84.800 285.560 85.120 ;
        RECT 285.640 84.800 285.960 85.120 ;
        RECT 286.040 84.800 286.360 85.120 ;
        RECT 286.440 84.800 286.760 85.120 ;
        RECT 286.840 84.800 287.160 85.120 ;
        RECT 287.240 84.800 287.560 85.120 ;
        RECT 4.620 66.000 4.940 66.320 ;
        RECT 5.020 66.000 5.340 66.320 ;
        RECT 5.420 66.000 5.740 66.320 ;
        RECT 5.820 66.000 6.140 66.320 ;
        RECT 6.220 66.000 6.540 66.320 ;
        RECT 6.620 66.000 6.940 66.320 ;
        RECT 7.020 66.000 7.340 66.320 ;
        RECT 7.420 66.000 7.740 66.320 ;
        RECT 7.820 66.000 8.140 66.320 ;
        RECT 8.220 66.000 8.540 66.320 ;
        RECT 8.620 66.000 8.940 66.320 ;
        RECT 9.020 66.000 9.340 66.320 ;
        RECT 9.420 66.000 9.740 66.320 ;
        RECT 9.820 66.000 10.140 66.320 ;
        RECT 10.220 66.000 10.540 66.320 ;
        RECT 10.620 66.000 10.940 66.320 ;
        RECT 11.020 66.000 11.340 66.320 ;
        RECT 11.420 66.000 11.740 66.320 ;
        RECT 11.820 66.000 12.140 66.320 ;
        RECT 12.220 66.000 12.540 66.320 ;
        RECT 279.640 66.000 279.960 66.320 ;
        RECT 280.040 66.000 280.360 66.320 ;
        RECT 280.440 66.000 280.760 66.320 ;
        RECT 280.840 66.000 281.160 66.320 ;
        RECT 281.240 66.000 281.560 66.320 ;
        RECT 281.640 66.000 281.960 66.320 ;
        RECT 282.040 66.000 282.360 66.320 ;
        RECT 282.440 66.000 282.760 66.320 ;
        RECT 282.840 66.000 283.160 66.320 ;
        RECT 283.240 66.000 283.560 66.320 ;
        RECT 283.640 66.000 283.960 66.320 ;
        RECT 284.040 66.000 284.360 66.320 ;
        RECT 284.440 66.000 284.760 66.320 ;
        RECT 284.840 66.000 285.160 66.320 ;
        RECT 285.240 66.000 285.560 66.320 ;
        RECT 285.640 66.000 285.960 66.320 ;
        RECT 286.040 66.000 286.360 66.320 ;
        RECT 286.440 66.000 286.760 66.320 ;
        RECT 286.840 66.000 287.160 66.320 ;
        RECT 287.240 66.000 287.560 66.320 ;
        RECT 4.620 47.200 4.940 47.520 ;
        RECT 5.020 47.200 5.340 47.520 ;
        RECT 5.420 47.200 5.740 47.520 ;
        RECT 5.820 47.200 6.140 47.520 ;
        RECT 6.220 47.200 6.540 47.520 ;
        RECT 6.620 47.200 6.940 47.520 ;
        RECT 7.020 47.200 7.340 47.520 ;
        RECT 7.420 47.200 7.740 47.520 ;
        RECT 7.820 47.200 8.140 47.520 ;
        RECT 8.220 47.200 8.540 47.520 ;
        RECT 8.620 47.200 8.940 47.520 ;
        RECT 9.020 47.200 9.340 47.520 ;
        RECT 9.420 47.200 9.740 47.520 ;
        RECT 9.820 47.200 10.140 47.520 ;
        RECT 10.220 47.200 10.540 47.520 ;
        RECT 10.620 47.200 10.940 47.520 ;
        RECT 11.020 47.200 11.340 47.520 ;
        RECT 11.420 47.200 11.740 47.520 ;
        RECT 11.820 47.200 12.140 47.520 ;
        RECT 12.220 47.200 12.540 47.520 ;
        RECT 279.640 47.200 279.960 47.520 ;
        RECT 280.040 47.200 280.360 47.520 ;
        RECT 280.440 47.200 280.760 47.520 ;
        RECT 280.840 47.200 281.160 47.520 ;
        RECT 281.240 47.200 281.560 47.520 ;
        RECT 281.640 47.200 281.960 47.520 ;
        RECT 282.040 47.200 282.360 47.520 ;
        RECT 282.440 47.200 282.760 47.520 ;
        RECT 282.840 47.200 283.160 47.520 ;
        RECT 283.240 47.200 283.560 47.520 ;
        RECT 283.640 47.200 283.960 47.520 ;
        RECT 284.040 47.200 284.360 47.520 ;
        RECT 284.440 47.200 284.760 47.520 ;
        RECT 284.840 47.200 285.160 47.520 ;
        RECT 285.240 47.200 285.560 47.520 ;
        RECT 285.640 47.200 285.960 47.520 ;
        RECT 286.040 47.200 286.360 47.520 ;
        RECT 286.440 47.200 286.760 47.520 ;
        RECT 286.840 47.200 287.160 47.520 ;
        RECT 287.240 47.200 287.560 47.520 ;
        RECT 4.620 28.400 4.940 28.720 ;
        RECT 5.020 28.400 5.340 28.720 ;
        RECT 5.420 28.400 5.740 28.720 ;
        RECT 5.820 28.400 6.140 28.720 ;
        RECT 6.220 28.400 6.540 28.720 ;
        RECT 6.620 28.400 6.940 28.720 ;
        RECT 7.020 28.400 7.340 28.720 ;
        RECT 7.420 28.400 7.740 28.720 ;
        RECT 7.820 28.400 8.140 28.720 ;
        RECT 8.220 28.400 8.540 28.720 ;
        RECT 8.620 28.400 8.940 28.720 ;
        RECT 9.020 28.400 9.340 28.720 ;
        RECT 9.420 28.400 9.740 28.720 ;
        RECT 9.820 28.400 10.140 28.720 ;
        RECT 10.220 28.400 10.540 28.720 ;
        RECT 10.620 28.400 10.940 28.720 ;
        RECT 11.020 28.400 11.340 28.720 ;
        RECT 11.420 28.400 11.740 28.720 ;
        RECT 11.820 28.400 12.140 28.720 ;
        RECT 12.220 28.400 12.540 28.720 ;
        RECT 279.640 28.400 279.960 28.720 ;
        RECT 280.040 28.400 280.360 28.720 ;
        RECT 280.440 28.400 280.760 28.720 ;
        RECT 280.840 28.400 281.160 28.720 ;
        RECT 281.240 28.400 281.560 28.720 ;
        RECT 281.640 28.400 281.960 28.720 ;
        RECT 282.040 28.400 282.360 28.720 ;
        RECT 282.440 28.400 282.760 28.720 ;
        RECT 282.840 28.400 283.160 28.720 ;
        RECT 283.240 28.400 283.560 28.720 ;
        RECT 283.640 28.400 283.960 28.720 ;
        RECT 284.040 28.400 284.360 28.720 ;
        RECT 284.440 28.400 284.760 28.720 ;
        RECT 284.840 28.400 285.160 28.720 ;
        RECT 285.240 28.400 285.560 28.720 ;
        RECT 285.640 28.400 285.960 28.720 ;
        RECT 286.040 28.400 286.360 28.720 ;
        RECT 286.440 28.400 286.760 28.720 ;
        RECT 286.840 28.400 287.160 28.720 ;
        RECT 287.240 28.400 287.560 28.720 ;
      LAYER met4 ;
        RECT 4.500 0.000 12.660 282.880 ;
        RECT 30.280 242.915 31.880 243.010 ;
        RECT 33.880 242.915 35.480 243.010 ;
        RECT 37.480 242.915 39.080 243.010 ;
        RECT 41.080 242.915 42.680 243.010 ;
        RECT 44.680 242.915 46.280 243.010 ;
        RECT 48.280 242.915 49.880 243.010 ;
        RECT 51.880 242.915 53.480 243.010 ;
        RECT 55.480 242.915 57.080 243.010 ;
        RECT 59.080 242.915 60.680 243.010 ;
        RECT 62.680 242.915 64.280 243.010 ;
        RECT 30.280 241.305 31.890 242.915 ;
        RECT 33.875 241.305 35.485 242.915 ;
        RECT 37.470 241.305 39.080 242.915 ;
        RECT 41.065 241.305 42.680 242.915 ;
        RECT 44.660 241.305 46.280 242.915 ;
        RECT 48.255 241.305 49.880 242.915 ;
        RECT 51.850 241.305 53.480 242.915 ;
        RECT 55.445 241.305 57.080 242.915 ;
        RECT 59.040 241.305 60.680 242.915 ;
        RECT 62.635 241.305 64.280 242.915 ;
        RECT 30.280 239.415 31.880 241.305 ;
        RECT 33.880 239.415 35.480 241.305 ;
        RECT 37.480 239.415 39.080 241.305 ;
        RECT 41.080 239.415 42.680 241.305 ;
        RECT 44.680 239.415 46.280 241.305 ;
        RECT 48.280 239.415 49.880 241.305 ;
        RECT 51.880 239.415 53.480 241.305 ;
        RECT 55.480 239.415 57.080 241.305 ;
        RECT 59.080 239.415 60.680 241.305 ;
        RECT 62.680 239.415 64.280 241.305 ;
        RECT 30.280 237.805 31.890 239.415 ;
        RECT 33.875 237.805 35.485 239.415 ;
        RECT 37.470 237.805 39.080 239.415 ;
        RECT 41.065 237.805 42.680 239.415 ;
        RECT 44.660 237.805 46.280 239.415 ;
        RECT 48.255 237.805 49.880 239.415 ;
        RECT 51.850 237.805 53.480 239.415 ;
        RECT 55.445 237.805 57.080 239.415 ;
        RECT 59.040 237.805 60.680 239.415 ;
        RECT 62.635 237.805 64.280 239.415 ;
        RECT 30.280 236.610 31.880 237.805 ;
        RECT 33.880 236.610 35.480 237.805 ;
        RECT 37.480 236.610 39.080 237.805 ;
        RECT 41.080 236.610 42.680 237.805 ;
        RECT 44.680 236.610 46.280 237.805 ;
        RECT 48.280 236.610 49.880 237.805 ;
        RECT 51.880 236.610 53.480 237.805 ;
        RECT 55.480 236.610 57.080 237.805 ;
        RECT 59.080 236.610 60.680 237.805 ;
        RECT 62.680 236.610 64.280 237.805 ;
        RECT 67.520 242.915 69.120 243.010 ;
        RECT 71.120 242.915 72.720 243.010 ;
        RECT 74.720 242.915 76.320 243.010 ;
        RECT 78.320 242.915 79.920 243.010 ;
        RECT 81.920 242.915 83.520 243.010 ;
        RECT 85.520 242.915 87.120 243.010 ;
        RECT 89.120 242.915 90.720 243.010 ;
        RECT 92.720 242.915 94.320 243.010 ;
        RECT 96.320 242.915 97.920 243.010 ;
        RECT 99.920 242.915 101.520 243.010 ;
        RECT 67.520 241.305 69.130 242.915 ;
        RECT 71.115 241.305 72.725 242.915 ;
        RECT 74.710 241.305 76.320 242.915 ;
        RECT 78.305 241.305 79.920 242.915 ;
        RECT 81.900 241.305 83.520 242.915 ;
        RECT 85.495 241.305 87.120 242.915 ;
        RECT 89.090 241.305 90.720 242.915 ;
        RECT 92.685 241.305 94.320 242.915 ;
        RECT 96.280 241.305 97.920 242.915 ;
        RECT 99.875 241.305 101.520 242.915 ;
        RECT 67.520 239.415 69.120 241.305 ;
        RECT 71.120 239.415 72.720 241.305 ;
        RECT 74.720 239.415 76.320 241.305 ;
        RECT 78.320 239.415 79.920 241.305 ;
        RECT 81.920 239.415 83.520 241.305 ;
        RECT 85.520 239.415 87.120 241.305 ;
        RECT 89.120 239.415 90.720 241.305 ;
        RECT 92.720 239.415 94.320 241.305 ;
        RECT 96.320 239.415 97.920 241.305 ;
        RECT 99.920 239.415 101.520 241.305 ;
        RECT 67.520 237.805 69.130 239.415 ;
        RECT 71.115 237.805 72.725 239.415 ;
        RECT 74.710 237.805 76.320 239.415 ;
        RECT 78.305 237.805 79.920 239.415 ;
        RECT 81.900 237.805 83.520 239.415 ;
        RECT 85.495 237.805 87.120 239.415 ;
        RECT 89.090 237.805 90.720 239.415 ;
        RECT 92.685 237.805 94.320 239.415 ;
        RECT 96.280 237.805 97.920 239.415 ;
        RECT 99.875 237.805 101.520 239.415 ;
        RECT 67.520 236.610 69.120 237.805 ;
        RECT 71.120 236.610 72.720 237.805 ;
        RECT 74.720 236.610 76.320 237.805 ;
        RECT 78.320 236.610 79.920 237.805 ;
        RECT 81.920 236.610 83.520 237.805 ;
        RECT 85.520 236.610 87.120 237.805 ;
        RECT 89.120 236.610 90.720 237.805 ;
        RECT 92.720 236.610 94.320 237.805 ;
        RECT 96.320 236.610 97.920 237.805 ;
        RECT 99.920 236.610 101.520 237.805 ;
        RECT 29.590 236.010 65.430 236.610 ;
        RECT 66.830 236.010 102.670 236.610 ;
        RECT 64.940 235.060 65.240 236.010 ;
        RECT 67.010 235.060 67.310 236.010 ;
        RECT 88.400 235.685 88.700 236.010 ;
        RECT 88.385 235.355 88.715 235.685 ;
        RECT 64.940 234.760 67.310 235.060 ;
        RECT 30.280 224.115 31.880 224.210 ;
        RECT 33.880 224.115 35.480 224.210 ;
        RECT 37.480 224.115 39.080 224.210 ;
        RECT 41.080 224.115 42.680 224.210 ;
        RECT 44.680 224.115 46.280 224.210 ;
        RECT 48.280 224.115 49.880 224.210 ;
        RECT 51.880 224.115 53.480 224.210 ;
        RECT 55.480 224.115 57.080 224.210 ;
        RECT 59.080 224.115 60.680 224.210 ;
        RECT 62.680 224.115 64.280 224.210 ;
        RECT 30.280 222.505 31.890 224.115 ;
        RECT 33.875 222.505 35.485 224.115 ;
        RECT 37.470 222.505 39.080 224.115 ;
        RECT 41.065 222.505 42.680 224.115 ;
        RECT 44.660 222.505 46.280 224.115 ;
        RECT 48.255 222.505 49.880 224.115 ;
        RECT 51.850 222.505 53.480 224.115 ;
        RECT 55.445 222.505 57.080 224.115 ;
        RECT 59.040 222.505 60.680 224.115 ;
        RECT 62.635 222.505 64.280 224.115 ;
        RECT 30.280 220.615 31.880 222.505 ;
        RECT 33.880 220.615 35.480 222.505 ;
        RECT 37.480 220.615 39.080 222.505 ;
        RECT 41.080 220.615 42.680 222.505 ;
        RECT 44.680 220.615 46.280 222.505 ;
        RECT 48.280 220.615 49.880 222.505 ;
        RECT 51.880 220.615 53.480 222.505 ;
        RECT 55.480 220.615 57.080 222.505 ;
        RECT 59.080 220.615 60.680 222.505 ;
        RECT 62.680 220.615 64.280 222.505 ;
        RECT 30.280 219.005 31.890 220.615 ;
        RECT 33.875 219.005 35.485 220.615 ;
        RECT 37.470 219.005 39.080 220.615 ;
        RECT 41.065 219.005 42.680 220.615 ;
        RECT 44.660 219.005 46.280 220.615 ;
        RECT 48.255 219.005 49.880 220.615 ;
        RECT 51.850 219.005 53.480 220.615 ;
        RECT 55.445 219.005 57.080 220.615 ;
        RECT 59.040 219.005 60.680 220.615 ;
        RECT 62.635 219.005 64.280 220.615 ;
        RECT 30.280 217.810 31.880 219.005 ;
        RECT 33.880 217.810 35.480 219.005 ;
        RECT 37.480 217.810 39.080 219.005 ;
        RECT 41.080 217.810 42.680 219.005 ;
        RECT 44.680 217.810 46.280 219.005 ;
        RECT 48.280 217.810 49.880 219.005 ;
        RECT 51.880 217.810 53.480 219.005 ;
        RECT 55.480 217.810 57.080 219.005 ;
        RECT 59.080 217.810 60.680 219.005 ;
        RECT 62.680 217.810 64.280 219.005 ;
        RECT 29.590 217.210 65.430 217.810 ;
        RECT 33.200 205.410 33.500 217.210 ;
        RECT 41.480 216.775 41.780 217.210 ;
        RECT 41.465 216.445 41.795 216.775 ;
        RECT 32.240 205.315 33.840 205.410 ;
        RECT 35.840 205.315 37.440 205.410 ;
        RECT 39.440 205.315 41.040 205.410 ;
        RECT 43.040 205.315 44.640 205.410 ;
        RECT 46.640 205.315 48.240 205.410 ;
        RECT 50.240 205.315 51.840 205.410 ;
        RECT 53.840 205.315 55.440 205.410 ;
        RECT 57.440 205.315 59.040 205.410 ;
        RECT 61.040 205.315 62.640 205.410 ;
        RECT 64.640 205.315 66.240 205.410 ;
        RECT 32.240 203.705 33.850 205.315 ;
        RECT 35.835 203.705 37.445 205.315 ;
        RECT 39.430 203.705 41.040 205.315 ;
        RECT 43.025 203.705 44.640 205.315 ;
        RECT 46.620 203.705 48.240 205.315 ;
        RECT 50.215 203.705 51.840 205.315 ;
        RECT 53.810 203.705 55.440 205.315 ;
        RECT 57.405 203.705 59.040 205.315 ;
        RECT 61.000 203.705 62.640 205.315 ;
        RECT 64.595 203.705 66.240 205.315 ;
        RECT 32.240 201.815 33.840 203.705 ;
        RECT 35.840 201.815 37.440 203.705 ;
        RECT 39.440 201.815 41.040 203.705 ;
        RECT 43.040 201.815 44.640 203.705 ;
        RECT 46.640 201.815 48.240 203.705 ;
        RECT 50.240 201.815 51.840 203.705 ;
        RECT 53.840 201.815 55.440 203.705 ;
        RECT 57.440 201.815 59.040 203.705 ;
        RECT 61.040 201.815 62.640 203.705 ;
        RECT 64.640 201.815 66.240 203.705 ;
        RECT 32.240 200.205 33.850 201.815 ;
        RECT 35.835 200.205 37.445 201.815 ;
        RECT 39.430 200.205 41.040 201.815 ;
        RECT 43.025 200.205 44.640 201.815 ;
        RECT 46.620 200.205 48.240 201.815 ;
        RECT 50.215 200.205 51.840 201.815 ;
        RECT 53.810 200.205 55.440 201.815 ;
        RECT 57.405 200.205 59.040 201.815 ;
        RECT 61.000 200.205 62.640 201.815 ;
        RECT 64.595 200.205 66.240 201.815 ;
        RECT 32.240 199.010 33.840 200.205 ;
        RECT 35.840 199.010 37.440 200.205 ;
        RECT 39.440 199.010 41.040 200.205 ;
        RECT 43.040 199.010 44.640 200.205 ;
        RECT 46.640 199.010 48.240 200.205 ;
        RECT 50.240 199.010 51.840 200.205 ;
        RECT 53.840 199.010 55.440 200.205 ;
        RECT 57.440 199.010 59.040 200.205 ;
        RECT 61.040 199.010 62.640 200.205 ;
        RECT 64.640 199.010 66.240 200.205 ;
        RECT 76.340 205.315 77.940 205.410 ;
        RECT 79.940 205.315 81.540 205.410 ;
        RECT 83.540 205.315 85.140 205.410 ;
        RECT 87.140 205.315 88.740 205.410 ;
        RECT 90.740 205.315 92.340 205.410 ;
        RECT 94.340 205.315 95.940 205.410 ;
        RECT 97.940 205.315 99.540 205.410 ;
        RECT 101.540 205.315 103.140 205.410 ;
        RECT 105.140 205.315 106.740 205.410 ;
        RECT 108.740 205.315 110.340 205.410 ;
        RECT 76.340 203.705 77.950 205.315 ;
        RECT 79.935 203.705 81.545 205.315 ;
        RECT 83.530 203.705 85.140 205.315 ;
        RECT 87.125 203.705 88.740 205.315 ;
        RECT 90.720 203.705 92.340 205.315 ;
        RECT 94.315 203.705 95.940 205.315 ;
        RECT 97.910 203.705 99.540 205.315 ;
        RECT 101.505 203.705 103.140 205.315 ;
        RECT 105.100 203.705 106.740 205.315 ;
        RECT 108.695 203.705 110.340 205.315 ;
        RECT 76.340 201.815 77.940 203.705 ;
        RECT 79.940 201.815 81.540 203.705 ;
        RECT 83.540 201.815 85.140 203.705 ;
        RECT 87.140 201.815 88.740 203.705 ;
        RECT 90.740 201.815 92.340 203.705 ;
        RECT 94.340 201.815 95.940 203.705 ;
        RECT 97.940 201.815 99.540 203.705 ;
        RECT 101.540 201.815 103.140 203.705 ;
        RECT 105.140 201.815 106.740 203.705 ;
        RECT 108.740 201.815 110.340 203.705 ;
        RECT 76.340 200.205 77.950 201.815 ;
        RECT 79.935 200.205 81.545 201.815 ;
        RECT 83.530 200.205 85.140 201.815 ;
        RECT 87.125 200.205 88.740 201.815 ;
        RECT 90.720 200.205 92.340 201.815 ;
        RECT 94.315 200.205 95.940 201.815 ;
        RECT 97.910 200.205 99.540 201.815 ;
        RECT 101.505 200.205 103.140 201.815 ;
        RECT 105.100 200.205 106.740 201.815 ;
        RECT 108.695 200.205 110.340 201.815 ;
        RECT 76.340 199.010 77.940 200.205 ;
        RECT 79.940 199.010 81.540 200.205 ;
        RECT 83.540 199.010 85.140 200.205 ;
        RECT 87.140 199.010 88.740 200.205 ;
        RECT 90.740 199.010 92.340 200.205 ;
        RECT 94.340 199.010 95.940 200.205 ;
        RECT 97.940 199.010 99.540 200.205 ;
        RECT 101.540 199.010 103.140 200.205 ;
        RECT 105.140 199.010 106.740 200.205 ;
        RECT 108.740 199.010 110.340 200.205 ;
        RECT 31.550 198.410 67.390 199.010 ;
        RECT 75.650 198.410 111.490 199.010 ;
        RECT 77.345 198.145 77.675 198.410 ;
        RECT 279.520 0.000 287.680 282.880 ;
      LAYER via4 ;
        RECT 4.790 270.770 12.370 278.350 ;
        RECT 279.810 270.770 287.390 278.350 ;
        RECT 4.790 4.370 12.370 11.950 ;
        RECT 279.810 4.370 287.390 11.950 ;
      LAYER met5 ;
        RECT 0.000 270.480 292.560 278.640 ;
        RECT 0.000 4.080 292.560 12.240 ;
    END
  END VSS
  PIN VDD
    ANTENNAGATEAREA 154.800003 ;
    ANTENNADIFFAREA 211.013992 ;
    PORT
      LAYER nwell ;
        RECT 123.660 243.895 262.190 245.060 ;
        RECT 123.660 236.830 262.195 243.895 ;
        RECT 124.145 236.825 262.195 236.830 ;
        RECT 74.660 225.095 213.190 226.260 ;
        RECT 74.660 218.030 213.195 225.095 ;
        RECT 75.145 218.025 213.195 218.030 ;
        RECT 112.880 206.295 141.490 207.460 ;
        RECT 146.200 206.295 174.810 207.460 ;
        RECT 112.880 199.230 141.495 206.295 ;
        RECT 146.200 199.230 174.815 206.295 ;
        RECT 113.365 199.225 141.495 199.230 ;
        RECT 146.685 199.225 174.815 199.230 ;
        RECT 186.870 187.495 201.740 188.660 ;
        RECT 186.870 180.430 201.745 187.495 ;
        RECT 187.355 180.425 201.745 180.430 ;
        RECT 186.870 149.895 201.740 151.060 ;
        RECT 186.870 142.830 201.745 149.895 ;
        RECT 187.355 142.825 201.745 142.830 ;
        RECT 123.660 93.495 262.190 94.660 ;
        RECT 123.660 86.430 262.195 93.495 ;
        RECT 124.145 86.425 262.195 86.430 ;
      LAYER li1 ;
        RECT 29.590 244.610 65.430 244.910 ;
        RECT 66.830 244.610 102.670 244.910 ;
        RECT 104.160 244.610 116.360 244.910 ;
        RECT 119.100 244.610 122.170 244.910 ;
        RECT 123.660 244.610 262.190 244.910 ;
        RECT 123.800 243.560 124.100 244.610 ;
        RECT 129.040 244.210 129.840 244.610 ;
        RECT 135.540 244.210 136.340 244.610 ;
        RECT 142.040 244.210 142.840 244.610 ;
        RECT 148.540 244.210 149.340 244.610 ;
        RECT 155.040 244.210 155.840 244.610 ;
        RECT 161.540 244.210 162.340 244.610 ;
        RECT 168.040 244.210 168.840 244.610 ;
        RECT 174.540 244.210 175.340 244.610 ;
        RECT 181.040 244.210 181.840 244.610 ;
        RECT 187.540 244.210 188.340 244.610 ;
        RECT 194.040 244.210 194.840 244.610 ;
        RECT 200.540 244.210 201.340 244.610 ;
        RECT 207.040 244.210 207.840 244.610 ;
        RECT 213.540 244.210 214.340 244.610 ;
        RECT 220.040 244.210 220.840 244.610 ;
        RECT 226.540 244.210 227.340 244.610 ;
        RECT 233.040 244.210 233.840 244.610 ;
        RECT 239.540 244.210 240.340 244.610 ;
        RECT 246.040 244.210 246.840 244.610 ;
        RECT 252.540 244.210 253.340 244.610 ;
        RECT 124.450 243.810 262.190 244.010 ;
        RECT 126.675 237.115 126.845 243.810 ;
        RECT 131.255 237.115 131.425 243.810 ;
        RECT 135.835 237.115 136.005 243.810 ;
        RECT 140.415 237.115 140.585 243.810 ;
        RECT 144.995 237.115 145.165 243.810 ;
        RECT 149.575 237.115 149.745 243.810 ;
        RECT 154.155 237.115 154.325 243.810 ;
        RECT 158.735 237.115 158.905 243.810 ;
        RECT 163.315 237.115 163.485 243.810 ;
        RECT 167.895 237.115 168.065 243.810 ;
        RECT 172.475 237.115 172.645 243.810 ;
        RECT 177.055 237.115 177.225 243.810 ;
        RECT 181.635 237.115 181.805 243.810 ;
        RECT 186.215 237.115 186.385 243.810 ;
        RECT 190.795 237.115 190.965 243.810 ;
        RECT 195.375 237.115 195.545 243.810 ;
        RECT 199.955 237.115 200.125 243.810 ;
        RECT 204.535 237.115 204.705 243.810 ;
        RECT 209.115 237.115 209.285 243.810 ;
        RECT 213.695 237.115 213.865 243.810 ;
        RECT 218.275 237.115 218.445 243.810 ;
        RECT 222.855 237.115 223.025 243.810 ;
        RECT 227.435 237.115 227.605 243.810 ;
        RECT 232.015 237.115 232.185 243.810 ;
        RECT 236.595 237.115 236.765 243.810 ;
        RECT 241.175 237.115 241.345 243.810 ;
        RECT 245.755 237.115 245.925 243.810 ;
        RECT 250.335 237.115 250.505 243.810 ;
        RECT 254.915 237.115 255.085 243.810 ;
        RECT 259.495 237.115 259.665 243.810 ;
        RECT 29.590 225.810 65.430 226.110 ;
        RECT 70.100 225.810 73.170 226.110 ;
        RECT 74.660 225.810 213.190 226.110 ;
        RECT 214.800 225.810 261.700 226.110 ;
        RECT 74.800 224.760 75.100 225.810 ;
        RECT 80.040 225.410 80.840 225.810 ;
        RECT 86.540 225.410 87.340 225.810 ;
        RECT 93.040 225.410 93.840 225.810 ;
        RECT 99.540 225.410 100.340 225.810 ;
        RECT 106.040 225.410 106.840 225.810 ;
        RECT 112.540 225.410 113.340 225.810 ;
        RECT 119.040 225.410 119.840 225.810 ;
        RECT 125.540 225.410 126.340 225.810 ;
        RECT 132.040 225.410 132.840 225.810 ;
        RECT 138.540 225.410 139.340 225.810 ;
        RECT 145.040 225.410 145.840 225.810 ;
        RECT 151.540 225.410 152.340 225.810 ;
        RECT 158.040 225.410 158.840 225.810 ;
        RECT 164.540 225.410 165.340 225.810 ;
        RECT 171.040 225.410 171.840 225.810 ;
        RECT 177.540 225.410 178.340 225.810 ;
        RECT 184.040 225.410 184.840 225.810 ;
        RECT 190.540 225.410 191.340 225.810 ;
        RECT 197.040 225.410 197.840 225.810 ;
        RECT 203.540 225.410 204.340 225.810 ;
        RECT 75.450 225.010 213.190 225.210 ;
        RECT 77.675 218.315 77.845 225.010 ;
        RECT 82.255 218.315 82.425 225.010 ;
        RECT 86.835 218.315 87.005 225.010 ;
        RECT 91.415 218.315 91.585 225.010 ;
        RECT 95.995 218.315 96.165 225.010 ;
        RECT 100.575 218.315 100.745 225.010 ;
        RECT 105.155 218.315 105.325 225.010 ;
        RECT 109.735 218.315 109.905 225.010 ;
        RECT 114.315 218.315 114.485 225.010 ;
        RECT 118.895 218.315 119.065 225.010 ;
        RECT 123.475 218.315 123.645 225.010 ;
        RECT 128.055 218.315 128.225 225.010 ;
        RECT 132.635 218.315 132.805 225.010 ;
        RECT 137.215 218.315 137.385 225.010 ;
        RECT 141.795 218.315 141.965 225.010 ;
        RECT 146.375 218.315 146.545 225.010 ;
        RECT 150.955 218.315 151.125 225.010 ;
        RECT 155.535 218.315 155.705 225.010 ;
        RECT 160.115 218.315 160.285 225.010 ;
        RECT 164.695 218.315 164.865 225.010 ;
        RECT 169.275 218.315 169.445 225.010 ;
        RECT 173.855 218.315 174.025 225.010 ;
        RECT 178.435 218.315 178.605 225.010 ;
        RECT 183.015 218.315 183.185 225.010 ;
        RECT 187.595 218.315 187.765 225.010 ;
        RECT 192.175 218.315 192.345 225.010 ;
        RECT 196.755 218.315 196.925 225.010 ;
        RECT 201.335 218.315 201.505 225.010 ;
        RECT 205.915 218.315 206.085 225.010 ;
        RECT 210.495 218.315 210.665 225.010 ;
        RECT 31.550 207.010 67.390 207.310 ;
        RECT 75.650 207.010 111.490 207.310 ;
        RECT 112.880 207.010 141.490 207.310 ;
        RECT 146.200 207.010 174.810 207.310 ;
        RECT 185.890 207.010 207.280 207.310 ;
        RECT 208.920 207.010 262.520 207.310 ;
        RECT 113.020 205.960 113.320 207.010 ;
        RECT 118.260 206.610 119.060 207.010 ;
        RECT 124.760 206.610 125.560 207.010 ;
        RECT 131.260 206.610 132.060 207.010 ;
        RECT 113.670 206.210 141.490 206.410 ;
        RECT 115.895 199.515 116.065 206.210 ;
        RECT 120.475 199.515 120.645 206.210 ;
        RECT 124.345 206.125 124.515 206.210 ;
        RECT 125.055 199.515 125.225 206.210 ;
        RECT 129.635 199.515 129.805 206.210 ;
        RECT 134.215 199.515 134.385 206.210 ;
        RECT 138.795 199.515 138.965 206.210 ;
        RECT 146.340 205.960 146.640 207.010 ;
        RECT 151.580 206.610 152.380 207.010 ;
        RECT 158.080 206.610 158.880 207.010 ;
        RECT 164.580 206.610 165.380 207.010 ;
        RECT 146.990 206.210 174.810 206.410 ;
        RECT 149.215 199.515 149.385 206.210 ;
        RECT 153.795 199.515 153.965 206.210 ;
        RECT 158.375 199.515 158.545 206.210 ;
        RECT 162.955 199.515 163.125 206.210 ;
        RECT 167.535 199.515 167.705 206.210 ;
        RECT 172.115 199.515 172.285 206.210 ;
        RECT 113.370 198.475 141.490 198.580 ;
        RECT 113.370 198.305 141.535 198.475 ;
        RECT 113.370 198.280 141.490 198.305 ;
        RECT 59.960 188.210 66.660 188.510 ;
        RECT 68.390 188.210 80.590 188.510 ;
        RECT 82.110 188.210 94.310 188.510 ;
        RECT 95.840 188.210 110.900 188.510 ;
        RECT 112.490 188.210 124.690 188.510 ;
        RECT 126.600 188.210 147.990 188.510 ;
        RECT 149.640 188.210 185.480 188.510 ;
        RECT 186.870 188.210 201.740 188.510 ;
        RECT 208.920 188.210 262.520 188.510 ;
        RECT 187.010 187.160 187.310 188.210 ;
        RECT 192.250 187.810 193.050 188.210 ;
        RECT 187.660 187.410 201.740 187.610 ;
        RECT 189.885 180.715 190.055 187.410 ;
        RECT 194.465 180.715 194.635 187.410 ;
        RECT 199.045 180.715 199.215 187.410 ;
        RECT 96.320 169.410 108.520 169.710 ;
        RECT 110.050 169.410 125.110 169.710 ;
        RECT 131.020 169.410 166.860 169.710 ;
        RECT 168.260 169.410 204.100 169.710 ;
        RECT 208.920 169.410 262.520 169.710 ;
        RECT 82.600 150.610 94.800 150.910 ;
        RECT 96.320 150.610 108.520 150.910 ;
        RECT 110.040 150.610 122.240 150.910 ;
        RECT 136.010 150.610 148.210 150.910 ;
        RECT 149.640 150.610 185.480 150.910 ;
        RECT 186.870 150.610 201.740 150.910 ;
        RECT 208.920 150.610 262.520 150.910 ;
        RECT 187.010 149.560 187.310 150.610 ;
        RECT 192.250 150.210 193.050 150.610 ;
        RECT 187.660 149.995 201.740 150.010 ;
        RECT 187.660 149.825 201.795 149.995 ;
        RECT 187.660 149.810 201.740 149.825 ;
        RECT 189.885 143.115 190.055 149.810 ;
        RECT 194.465 143.115 194.635 149.810 ;
        RECT 199.045 143.115 199.215 149.810 ;
        RECT 112.000 131.810 124.200 132.110 ;
        RECT 126.600 131.810 147.990 132.110 ;
        RECT 149.640 131.810 185.480 132.110 ;
        RECT 186.970 131.810 199.170 132.110 ;
        RECT 200.690 131.810 212.890 132.110 ;
        RECT 214.410 131.810 226.610 132.110 ;
        RECT 228.130 131.810 240.330 132.110 ;
        RECT 241.850 131.810 254.050 132.110 ;
        RECT 119.350 113.010 131.550 113.310 ;
        RECT 136.010 113.010 148.210 113.310 ;
        RECT 149.730 113.010 161.930 113.310 ;
        RECT 165.900 113.010 178.100 113.310 ;
        RECT 186.970 113.010 199.170 113.310 ;
        RECT 200.690 113.010 212.890 113.310 ;
        RECT 241.850 113.010 254.050 113.310 ;
        RECT 123.660 94.210 262.190 94.510 ;
        RECT 123.800 93.160 124.100 94.210 ;
        RECT 129.040 93.810 129.840 94.210 ;
        RECT 135.540 93.810 136.340 94.210 ;
        RECT 142.040 93.810 142.840 94.210 ;
        RECT 148.540 93.810 149.340 94.210 ;
        RECT 155.040 93.810 155.840 94.210 ;
        RECT 161.540 93.810 162.340 94.210 ;
        RECT 168.040 93.810 168.840 94.210 ;
        RECT 174.540 93.810 175.340 94.210 ;
        RECT 181.040 93.810 181.840 94.210 ;
        RECT 187.540 93.810 188.340 94.210 ;
        RECT 194.040 93.810 194.840 94.210 ;
        RECT 200.540 93.810 201.340 94.210 ;
        RECT 207.040 93.810 207.840 94.210 ;
        RECT 213.540 93.810 214.340 94.210 ;
        RECT 220.040 93.810 220.840 94.210 ;
        RECT 226.540 93.810 227.340 94.210 ;
        RECT 233.040 93.810 233.840 94.210 ;
        RECT 239.540 93.810 240.340 94.210 ;
        RECT 246.040 93.810 246.840 94.210 ;
        RECT 252.540 93.810 253.340 94.210 ;
        RECT 124.450 93.410 262.190 93.610 ;
        RECT 126.675 86.715 126.845 93.410 ;
        RECT 131.255 86.715 131.425 93.410 ;
        RECT 135.835 86.715 136.005 93.410 ;
        RECT 140.415 86.715 140.585 93.410 ;
        RECT 144.995 86.715 145.165 93.410 ;
        RECT 149.575 86.715 149.745 93.410 ;
        RECT 154.155 86.715 154.325 93.410 ;
        RECT 158.735 86.715 158.905 93.410 ;
        RECT 163.315 86.715 163.485 93.410 ;
        RECT 167.895 86.715 168.065 93.410 ;
        RECT 172.475 86.715 172.645 93.410 ;
        RECT 177.055 86.715 177.225 93.410 ;
        RECT 181.635 86.715 181.805 93.410 ;
        RECT 186.215 86.715 186.385 93.410 ;
        RECT 190.795 86.715 190.965 93.410 ;
        RECT 195.375 86.715 195.545 93.410 ;
        RECT 199.955 86.715 200.125 93.410 ;
        RECT 204.535 86.715 204.705 93.410 ;
        RECT 209.115 86.715 209.285 93.410 ;
        RECT 213.695 86.715 213.865 93.410 ;
        RECT 218.275 86.715 218.445 93.410 ;
        RECT 222.855 86.715 223.025 93.410 ;
        RECT 227.435 86.715 227.605 93.410 ;
        RECT 232.015 86.715 232.185 93.410 ;
        RECT 236.595 86.715 236.765 93.410 ;
        RECT 241.175 86.715 241.345 93.410 ;
        RECT 245.755 86.715 245.925 93.410 ;
        RECT 250.335 86.715 250.505 93.410 ;
        RECT 254.915 86.715 255.085 93.410 ;
        RECT 259.495 86.715 259.665 93.410 ;
        RECT 219.310 75.410 231.510 75.710 ;
        RECT 233.030 75.410 245.230 75.710 ;
        RECT 246.750 75.410 258.950 75.710 ;
        RECT 218.820 56.610 231.020 56.910 ;
        RECT 232.540 56.610 244.740 56.910 ;
        RECT 246.260 56.610 258.460 56.910 ;
        RECT 222.740 37.810 234.940 38.110 ;
        RECT 236.460 37.810 248.660 38.110 ;
        RECT 250.180 37.810 262.380 38.110 ;
      LAYER mcon ;
        RECT 30.505 244.675 30.675 244.845 ;
        RECT 32.505 244.675 32.675 244.845 ;
        RECT 34.505 244.675 34.675 244.845 ;
        RECT 36.505 244.675 36.675 244.845 ;
        RECT 38.505 244.675 38.675 244.845 ;
        RECT 40.505 244.675 40.675 244.845 ;
        RECT 42.505 244.675 42.675 244.845 ;
        RECT 44.505 244.675 44.675 244.845 ;
        RECT 46.505 244.675 46.675 244.845 ;
        RECT 48.505 244.675 48.675 244.845 ;
        RECT 50.505 244.675 50.675 244.845 ;
        RECT 52.505 244.675 52.675 244.845 ;
        RECT 54.505 244.675 54.675 244.845 ;
        RECT 56.505 244.675 56.675 244.845 ;
        RECT 58.505 244.675 58.675 244.845 ;
        RECT 60.505 244.675 60.675 244.845 ;
        RECT 62.505 244.675 62.675 244.845 ;
        RECT 64.505 244.675 64.675 244.845 ;
        RECT 67.745 244.675 67.915 244.845 ;
        RECT 69.745 244.675 69.915 244.845 ;
        RECT 71.745 244.675 71.915 244.845 ;
        RECT 73.745 244.675 73.915 244.845 ;
        RECT 75.745 244.675 75.915 244.845 ;
        RECT 77.745 244.675 77.915 244.845 ;
        RECT 79.745 244.675 79.915 244.845 ;
        RECT 81.745 244.675 81.915 244.845 ;
        RECT 83.745 244.675 83.915 244.845 ;
        RECT 85.745 244.675 85.915 244.845 ;
        RECT 87.745 244.675 87.915 244.845 ;
        RECT 89.745 244.675 89.915 244.845 ;
        RECT 91.745 244.675 91.915 244.845 ;
        RECT 93.745 244.675 93.915 244.845 ;
        RECT 95.745 244.675 95.915 244.845 ;
        RECT 97.745 244.675 97.915 244.845 ;
        RECT 99.745 244.675 99.915 244.845 ;
        RECT 101.745 244.675 101.915 244.845 ;
        RECT 105.075 244.675 105.245 244.845 ;
        RECT 106.075 244.675 106.245 244.845 ;
        RECT 107.075 244.675 107.245 244.845 ;
        RECT 108.075 244.675 108.245 244.845 ;
        RECT 109.075 244.675 109.245 244.845 ;
        RECT 110.075 244.675 110.245 244.845 ;
        RECT 111.075 244.675 111.245 244.845 ;
        RECT 112.075 244.675 112.245 244.845 ;
        RECT 113.075 244.675 113.245 244.845 ;
        RECT 114.075 244.675 114.245 244.845 ;
        RECT 115.075 244.675 115.245 244.845 ;
        RECT 120.505 244.675 120.675 244.845 ;
        RECT 125.065 244.675 125.235 244.845 ;
        RECT 127.065 244.675 127.235 244.845 ;
        RECT 129.065 244.675 129.235 244.845 ;
        RECT 131.065 244.675 131.235 244.845 ;
        RECT 133.065 244.675 133.235 244.845 ;
        RECT 135.065 244.675 135.235 244.845 ;
        RECT 137.065 244.675 137.235 244.845 ;
        RECT 139.065 244.675 139.235 244.845 ;
        RECT 141.065 244.675 141.235 244.845 ;
        RECT 143.065 244.675 143.235 244.845 ;
        RECT 145.065 244.675 145.235 244.845 ;
        RECT 147.065 244.675 147.235 244.845 ;
        RECT 149.065 244.675 149.235 244.845 ;
        RECT 151.065 244.675 151.235 244.845 ;
        RECT 153.065 244.675 153.235 244.845 ;
        RECT 155.065 244.675 155.235 244.845 ;
        RECT 157.065 244.675 157.235 244.845 ;
        RECT 159.065 244.675 159.235 244.845 ;
        RECT 161.065 244.675 161.235 244.845 ;
        RECT 163.065 244.675 163.235 244.845 ;
        RECT 165.065 244.675 165.235 244.845 ;
        RECT 167.065 244.675 167.235 244.845 ;
        RECT 169.065 244.675 169.235 244.845 ;
        RECT 171.065 244.675 171.235 244.845 ;
        RECT 173.065 244.675 173.235 244.845 ;
        RECT 175.065 244.675 175.235 244.845 ;
        RECT 177.065 244.675 177.235 244.845 ;
        RECT 179.065 244.675 179.235 244.845 ;
        RECT 181.065 244.675 181.235 244.845 ;
        RECT 183.065 244.675 183.235 244.845 ;
        RECT 185.065 244.675 185.235 244.845 ;
        RECT 187.065 244.675 187.235 244.845 ;
        RECT 189.065 244.675 189.235 244.845 ;
        RECT 191.065 244.675 191.235 244.845 ;
        RECT 193.065 244.675 193.235 244.845 ;
        RECT 195.065 244.675 195.235 244.845 ;
        RECT 197.065 244.675 197.235 244.845 ;
        RECT 199.065 244.675 199.235 244.845 ;
        RECT 201.065 244.675 201.235 244.845 ;
        RECT 203.065 244.675 203.235 244.845 ;
        RECT 205.065 244.675 205.235 244.845 ;
        RECT 207.065 244.675 207.235 244.845 ;
        RECT 209.065 244.675 209.235 244.845 ;
        RECT 211.065 244.675 211.235 244.845 ;
        RECT 213.065 244.675 213.235 244.845 ;
        RECT 215.065 244.675 215.235 244.845 ;
        RECT 217.065 244.675 217.235 244.845 ;
        RECT 219.065 244.675 219.235 244.845 ;
        RECT 221.065 244.675 221.235 244.845 ;
        RECT 223.065 244.675 223.235 244.845 ;
        RECT 225.065 244.675 225.235 244.845 ;
        RECT 227.065 244.675 227.235 244.845 ;
        RECT 229.065 244.675 229.235 244.845 ;
        RECT 231.065 244.675 231.235 244.845 ;
        RECT 233.065 244.675 233.235 244.845 ;
        RECT 235.065 244.675 235.235 244.845 ;
        RECT 237.065 244.675 237.235 244.845 ;
        RECT 239.065 244.675 239.235 244.845 ;
        RECT 241.065 244.675 241.235 244.845 ;
        RECT 243.065 244.675 243.235 244.845 ;
        RECT 245.065 244.675 245.235 244.845 ;
        RECT 247.065 244.675 247.235 244.845 ;
        RECT 249.065 244.675 249.235 244.845 ;
        RECT 251.065 244.675 251.235 244.845 ;
        RECT 253.065 244.675 253.235 244.845 ;
        RECT 255.065 244.675 255.235 244.845 ;
        RECT 257.065 244.675 257.235 244.845 ;
        RECT 259.065 244.675 259.235 244.845 ;
        RECT 261.065 244.675 261.235 244.845 ;
        RECT 126.675 243.335 126.845 243.505 ;
        RECT 126.675 242.975 126.845 243.145 ;
        RECT 126.675 242.615 126.845 242.785 ;
        RECT 126.675 242.255 126.845 242.425 ;
        RECT 126.675 241.895 126.845 242.065 ;
        RECT 126.675 241.535 126.845 241.705 ;
        RECT 126.675 241.175 126.845 241.345 ;
        RECT 126.675 240.815 126.845 240.985 ;
        RECT 126.675 240.455 126.845 240.625 ;
        RECT 126.675 240.095 126.845 240.265 ;
        RECT 126.675 239.735 126.845 239.905 ;
        RECT 126.675 239.375 126.845 239.545 ;
        RECT 126.675 239.015 126.845 239.185 ;
        RECT 126.675 238.655 126.845 238.825 ;
        RECT 126.675 238.295 126.845 238.465 ;
        RECT 126.675 237.935 126.845 238.105 ;
        RECT 126.675 237.575 126.845 237.745 ;
        RECT 126.675 237.215 126.845 237.385 ;
        RECT 131.255 243.335 131.425 243.505 ;
        RECT 131.255 242.975 131.425 243.145 ;
        RECT 131.255 242.615 131.425 242.785 ;
        RECT 131.255 242.255 131.425 242.425 ;
        RECT 131.255 241.895 131.425 242.065 ;
        RECT 131.255 241.535 131.425 241.705 ;
        RECT 131.255 241.175 131.425 241.345 ;
        RECT 131.255 240.815 131.425 240.985 ;
        RECT 131.255 240.455 131.425 240.625 ;
        RECT 131.255 240.095 131.425 240.265 ;
        RECT 131.255 239.735 131.425 239.905 ;
        RECT 131.255 239.375 131.425 239.545 ;
        RECT 131.255 239.015 131.425 239.185 ;
        RECT 131.255 238.655 131.425 238.825 ;
        RECT 131.255 238.295 131.425 238.465 ;
        RECT 131.255 237.935 131.425 238.105 ;
        RECT 131.255 237.575 131.425 237.745 ;
        RECT 131.255 237.215 131.425 237.385 ;
        RECT 135.835 243.335 136.005 243.505 ;
        RECT 135.835 242.975 136.005 243.145 ;
        RECT 135.835 242.615 136.005 242.785 ;
        RECT 135.835 242.255 136.005 242.425 ;
        RECT 135.835 241.895 136.005 242.065 ;
        RECT 135.835 241.535 136.005 241.705 ;
        RECT 135.835 241.175 136.005 241.345 ;
        RECT 135.835 240.815 136.005 240.985 ;
        RECT 135.835 240.455 136.005 240.625 ;
        RECT 135.835 240.095 136.005 240.265 ;
        RECT 135.835 239.735 136.005 239.905 ;
        RECT 135.835 239.375 136.005 239.545 ;
        RECT 135.835 239.015 136.005 239.185 ;
        RECT 135.835 238.655 136.005 238.825 ;
        RECT 135.835 238.295 136.005 238.465 ;
        RECT 135.835 237.935 136.005 238.105 ;
        RECT 135.835 237.575 136.005 237.745 ;
        RECT 135.835 237.215 136.005 237.385 ;
        RECT 140.415 243.335 140.585 243.505 ;
        RECT 140.415 242.975 140.585 243.145 ;
        RECT 140.415 242.615 140.585 242.785 ;
        RECT 140.415 242.255 140.585 242.425 ;
        RECT 140.415 241.895 140.585 242.065 ;
        RECT 140.415 241.535 140.585 241.705 ;
        RECT 140.415 241.175 140.585 241.345 ;
        RECT 140.415 240.815 140.585 240.985 ;
        RECT 140.415 240.455 140.585 240.625 ;
        RECT 140.415 240.095 140.585 240.265 ;
        RECT 140.415 239.735 140.585 239.905 ;
        RECT 140.415 239.375 140.585 239.545 ;
        RECT 140.415 239.015 140.585 239.185 ;
        RECT 140.415 238.655 140.585 238.825 ;
        RECT 140.415 238.295 140.585 238.465 ;
        RECT 140.415 237.935 140.585 238.105 ;
        RECT 140.415 237.575 140.585 237.745 ;
        RECT 140.415 237.215 140.585 237.385 ;
        RECT 144.995 243.335 145.165 243.505 ;
        RECT 144.995 242.975 145.165 243.145 ;
        RECT 144.995 242.615 145.165 242.785 ;
        RECT 144.995 242.255 145.165 242.425 ;
        RECT 144.995 241.895 145.165 242.065 ;
        RECT 144.995 241.535 145.165 241.705 ;
        RECT 144.995 241.175 145.165 241.345 ;
        RECT 144.995 240.815 145.165 240.985 ;
        RECT 144.995 240.455 145.165 240.625 ;
        RECT 144.995 240.095 145.165 240.265 ;
        RECT 144.995 239.735 145.165 239.905 ;
        RECT 144.995 239.375 145.165 239.545 ;
        RECT 144.995 239.015 145.165 239.185 ;
        RECT 144.995 238.655 145.165 238.825 ;
        RECT 144.995 238.295 145.165 238.465 ;
        RECT 144.995 237.935 145.165 238.105 ;
        RECT 144.995 237.575 145.165 237.745 ;
        RECT 144.995 237.215 145.165 237.385 ;
        RECT 149.575 243.335 149.745 243.505 ;
        RECT 149.575 242.975 149.745 243.145 ;
        RECT 149.575 242.615 149.745 242.785 ;
        RECT 149.575 242.255 149.745 242.425 ;
        RECT 149.575 241.895 149.745 242.065 ;
        RECT 149.575 241.535 149.745 241.705 ;
        RECT 149.575 241.175 149.745 241.345 ;
        RECT 149.575 240.815 149.745 240.985 ;
        RECT 149.575 240.455 149.745 240.625 ;
        RECT 149.575 240.095 149.745 240.265 ;
        RECT 149.575 239.735 149.745 239.905 ;
        RECT 149.575 239.375 149.745 239.545 ;
        RECT 149.575 239.015 149.745 239.185 ;
        RECT 149.575 238.655 149.745 238.825 ;
        RECT 149.575 238.295 149.745 238.465 ;
        RECT 149.575 237.935 149.745 238.105 ;
        RECT 149.575 237.575 149.745 237.745 ;
        RECT 149.575 237.215 149.745 237.385 ;
        RECT 154.155 243.335 154.325 243.505 ;
        RECT 154.155 242.975 154.325 243.145 ;
        RECT 154.155 242.615 154.325 242.785 ;
        RECT 154.155 242.255 154.325 242.425 ;
        RECT 154.155 241.895 154.325 242.065 ;
        RECT 154.155 241.535 154.325 241.705 ;
        RECT 154.155 241.175 154.325 241.345 ;
        RECT 154.155 240.815 154.325 240.985 ;
        RECT 154.155 240.455 154.325 240.625 ;
        RECT 154.155 240.095 154.325 240.265 ;
        RECT 154.155 239.735 154.325 239.905 ;
        RECT 154.155 239.375 154.325 239.545 ;
        RECT 154.155 239.015 154.325 239.185 ;
        RECT 154.155 238.655 154.325 238.825 ;
        RECT 154.155 238.295 154.325 238.465 ;
        RECT 154.155 237.935 154.325 238.105 ;
        RECT 154.155 237.575 154.325 237.745 ;
        RECT 154.155 237.215 154.325 237.385 ;
        RECT 158.735 243.335 158.905 243.505 ;
        RECT 158.735 242.975 158.905 243.145 ;
        RECT 158.735 242.615 158.905 242.785 ;
        RECT 158.735 242.255 158.905 242.425 ;
        RECT 158.735 241.895 158.905 242.065 ;
        RECT 158.735 241.535 158.905 241.705 ;
        RECT 158.735 241.175 158.905 241.345 ;
        RECT 158.735 240.815 158.905 240.985 ;
        RECT 158.735 240.455 158.905 240.625 ;
        RECT 158.735 240.095 158.905 240.265 ;
        RECT 158.735 239.735 158.905 239.905 ;
        RECT 158.735 239.375 158.905 239.545 ;
        RECT 158.735 239.015 158.905 239.185 ;
        RECT 158.735 238.655 158.905 238.825 ;
        RECT 158.735 238.295 158.905 238.465 ;
        RECT 158.735 237.935 158.905 238.105 ;
        RECT 158.735 237.575 158.905 237.745 ;
        RECT 158.735 237.215 158.905 237.385 ;
        RECT 163.315 243.335 163.485 243.505 ;
        RECT 163.315 242.975 163.485 243.145 ;
        RECT 163.315 242.615 163.485 242.785 ;
        RECT 163.315 242.255 163.485 242.425 ;
        RECT 163.315 241.895 163.485 242.065 ;
        RECT 163.315 241.535 163.485 241.705 ;
        RECT 163.315 241.175 163.485 241.345 ;
        RECT 163.315 240.815 163.485 240.985 ;
        RECT 163.315 240.455 163.485 240.625 ;
        RECT 163.315 240.095 163.485 240.265 ;
        RECT 163.315 239.735 163.485 239.905 ;
        RECT 163.315 239.375 163.485 239.545 ;
        RECT 163.315 239.015 163.485 239.185 ;
        RECT 163.315 238.655 163.485 238.825 ;
        RECT 163.315 238.295 163.485 238.465 ;
        RECT 163.315 237.935 163.485 238.105 ;
        RECT 163.315 237.575 163.485 237.745 ;
        RECT 163.315 237.215 163.485 237.385 ;
        RECT 167.895 243.335 168.065 243.505 ;
        RECT 167.895 242.975 168.065 243.145 ;
        RECT 167.895 242.615 168.065 242.785 ;
        RECT 167.895 242.255 168.065 242.425 ;
        RECT 167.895 241.895 168.065 242.065 ;
        RECT 167.895 241.535 168.065 241.705 ;
        RECT 167.895 241.175 168.065 241.345 ;
        RECT 167.895 240.815 168.065 240.985 ;
        RECT 167.895 240.455 168.065 240.625 ;
        RECT 167.895 240.095 168.065 240.265 ;
        RECT 167.895 239.735 168.065 239.905 ;
        RECT 167.895 239.375 168.065 239.545 ;
        RECT 167.895 239.015 168.065 239.185 ;
        RECT 167.895 238.655 168.065 238.825 ;
        RECT 167.895 238.295 168.065 238.465 ;
        RECT 167.895 237.935 168.065 238.105 ;
        RECT 167.895 237.575 168.065 237.745 ;
        RECT 167.895 237.215 168.065 237.385 ;
        RECT 172.475 243.335 172.645 243.505 ;
        RECT 172.475 242.975 172.645 243.145 ;
        RECT 172.475 242.615 172.645 242.785 ;
        RECT 172.475 242.255 172.645 242.425 ;
        RECT 172.475 241.895 172.645 242.065 ;
        RECT 172.475 241.535 172.645 241.705 ;
        RECT 172.475 241.175 172.645 241.345 ;
        RECT 172.475 240.815 172.645 240.985 ;
        RECT 172.475 240.455 172.645 240.625 ;
        RECT 172.475 240.095 172.645 240.265 ;
        RECT 172.475 239.735 172.645 239.905 ;
        RECT 172.475 239.375 172.645 239.545 ;
        RECT 172.475 239.015 172.645 239.185 ;
        RECT 172.475 238.655 172.645 238.825 ;
        RECT 172.475 238.295 172.645 238.465 ;
        RECT 172.475 237.935 172.645 238.105 ;
        RECT 172.475 237.575 172.645 237.745 ;
        RECT 172.475 237.215 172.645 237.385 ;
        RECT 177.055 243.335 177.225 243.505 ;
        RECT 177.055 242.975 177.225 243.145 ;
        RECT 177.055 242.615 177.225 242.785 ;
        RECT 177.055 242.255 177.225 242.425 ;
        RECT 177.055 241.895 177.225 242.065 ;
        RECT 177.055 241.535 177.225 241.705 ;
        RECT 177.055 241.175 177.225 241.345 ;
        RECT 177.055 240.815 177.225 240.985 ;
        RECT 177.055 240.455 177.225 240.625 ;
        RECT 177.055 240.095 177.225 240.265 ;
        RECT 177.055 239.735 177.225 239.905 ;
        RECT 177.055 239.375 177.225 239.545 ;
        RECT 177.055 239.015 177.225 239.185 ;
        RECT 177.055 238.655 177.225 238.825 ;
        RECT 177.055 238.295 177.225 238.465 ;
        RECT 177.055 237.935 177.225 238.105 ;
        RECT 177.055 237.575 177.225 237.745 ;
        RECT 177.055 237.215 177.225 237.385 ;
        RECT 181.635 243.335 181.805 243.505 ;
        RECT 181.635 242.975 181.805 243.145 ;
        RECT 181.635 242.615 181.805 242.785 ;
        RECT 181.635 242.255 181.805 242.425 ;
        RECT 181.635 241.895 181.805 242.065 ;
        RECT 181.635 241.535 181.805 241.705 ;
        RECT 181.635 241.175 181.805 241.345 ;
        RECT 181.635 240.815 181.805 240.985 ;
        RECT 181.635 240.455 181.805 240.625 ;
        RECT 181.635 240.095 181.805 240.265 ;
        RECT 181.635 239.735 181.805 239.905 ;
        RECT 181.635 239.375 181.805 239.545 ;
        RECT 181.635 239.015 181.805 239.185 ;
        RECT 181.635 238.655 181.805 238.825 ;
        RECT 181.635 238.295 181.805 238.465 ;
        RECT 181.635 237.935 181.805 238.105 ;
        RECT 181.635 237.575 181.805 237.745 ;
        RECT 181.635 237.215 181.805 237.385 ;
        RECT 186.215 243.335 186.385 243.505 ;
        RECT 186.215 242.975 186.385 243.145 ;
        RECT 186.215 242.615 186.385 242.785 ;
        RECT 186.215 242.255 186.385 242.425 ;
        RECT 186.215 241.895 186.385 242.065 ;
        RECT 186.215 241.535 186.385 241.705 ;
        RECT 186.215 241.175 186.385 241.345 ;
        RECT 186.215 240.815 186.385 240.985 ;
        RECT 186.215 240.455 186.385 240.625 ;
        RECT 186.215 240.095 186.385 240.265 ;
        RECT 186.215 239.735 186.385 239.905 ;
        RECT 186.215 239.375 186.385 239.545 ;
        RECT 186.215 239.015 186.385 239.185 ;
        RECT 186.215 238.655 186.385 238.825 ;
        RECT 186.215 238.295 186.385 238.465 ;
        RECT 186.215 237.935 186.385 238.105 ;
        RECT 186.215 237.575 186.385 237.745 ;
        RECT 186.215 237.215 186.385 237.385 ;
        RECT 190.795 243.335 190.965 243.505 ;
        RECT 190.795 242.975 190.965 243.145 ;
        RECT 190.795 242.615 190.965 242.785 ;
        RECT 190.795 242.255 190.965 242.425 ;
        RECT 190.795 241.895 190.965 242.065 ;
        RECT 190.795 241.535 190.965 241.705 ;
        RECT 190.795 241.175 190.965 241.345 ;
        RECT 190.795 240.815 190.965 240.985 ;
        RECT 190.795 240.455 190.965 240.625 ;
        RECT 190.795 240.095 190.965 240.265 ;
        RECT 190.795 239.735 190.965 239.905 ;
        RECT 190.795 239.375 190.965 239.545 ;
        RECT 190.795 239.015 190.965 239.185 ;
        RECT 190.795 238.655 190.965 238.825 ;
        RECT 190.795 238.295 190.965 238.465 ;
        RECT 190.795 237.935 190.965 238.105 ;
        RECT 190.795 237.575 190.965 237.745 ;
        RECT 190.795 237.215 190.965 237.385 ;
        RECT 195.375 243.335 195.545 243.505 ;
        RECT 195.375 242.975 195.545 243.145 ;
        RECT 195.375 242.615 195.545 242.785 ;
        RECT 195.375 242.255 195.545 242.425 ;
        RECT 195.375 241.895 195.545 242.065 ;
        RECT 195.375 241.535 195.545 241.705 ;
        RECT 195.375 241.175 195.545 241.345 ;
        RECT 195.375 240.815 195.545 240.985 ;
        RECT 195.375 240.455 195.545 240.625 ;
        RECT 195.375 240.095 195.545 240.265 ;
        RECT 195.375 239.735 195.545 239.905 ;
        RECT 195.375 239.375 195.545 239.545 ;
        RECT 195.375 239.015 195.545 239.185 ;
        RECT 195.375 238.655 195.545 238.825 ;
        RECT 195.375 238.295 195.545 238.465 ;
        RECT 195.375 237.935 195.545 238.105 ;
        RECT 195.375 237.575 195.545 237.745 ;
        RECT 195.375 237.215 195.545 237.385 ;
        RECT 199.955 243.335 200.125 243.505 ;
        RECT 199.955 242.975 200.125 243.145 ;
        RECT 199.955 242.615 200.125 242.785 ;
        RECT 199.955 242.255 200.125 242.425 ;
        RECT 199.955 241.895 200.125 242.065 ;
        RECT 199.955 241.535 200.125 241.705 ;
        RECT 199.955 241.175 200.125 241.345 ;
        RECT 199.955 240.815 200.125 240.985 ;
        RECT 199.955 240.455 200.125 240.625 ;
        RECT 199.955 240.095 200.125 240.265 ;
        RECT 199.955 239.735 200.125 239.905 ;
        RECT 199.955 239.375 200.125 239.545 ;
        RECT 199.955 239.015 200.125 239.185 ;
        RECT 199.955 238.655 200.125 238.825 ;
        RECT 199.955 238.295 200.125 238.465 ;
        RECT 199.955 237.935 200.125 238.105 ;
        RECT 199.955 237.575 200.125 237.745 ;
        RECT 199.955 237.215 200.125 237.385 ;
        RECT 204.535 243.335 204.705 243.505 ;
        RECT 204.535 242.975 204.705 243.145 ;
        RECT 204.535 242.615 204.705 242.785 ;
        RECT 204.535 242.255 204.705 242.425 ;
        RECT 204.535 241.895 204.705 242.065 ;
        RECT 204.535 241.535 204.705 241.705 ;
        RECT 204.535 241.175 204.705 241.345 ;
        RECT 204.535 240.815 204.705 240.985 ;
        RECT 204.535 240.455 204.705 240.625 ;
        RECT 204.535 240.095 204.705 240.265 ;
        RECT 204.535 239.735 204.705 239.905 ;
        RECT 204.535 239.375 204.705 239.545 ;
        RECT 204.535 239.015 204.705 239.185 ;
        RECT 204.535 238.655 204.705 238.825 ;
        RECT 204.535 238.295 204.705 238.465 ;
        RECT 204.535 237.935 204.705 238.105 ;
        RECT 204.535 237.575 204.705 237.745 ;
        RECT 204.535 237.215 204.705 237.385 ;
        RECT 209.115 243.335 209.285 243.505 ;
        RECT 209.115 242.975 209.285 243.145 ;
        RECT 209.115 242.615 209.285 242.785 ;
        RECT 209.115 242.255 209.285 242.425 ;
        RECT 209.115 241.895 209.285 242.065 ;
        RECT 209.115 241.535 209.285 241.705 ;
        RECT 209.115 241.175 209.285 241.345 ;
        RECT 209.115 240.815 209.285 240.985 ;
        RECT 209.115 240.455 209.285 240.625 ;
        RECT 209.115 240.095 209.285 240.265 ;
        RECT 209.115 239.735 209.285 239.905 ;
        RECT 209.115 239.375 209.285 239.545 ;
        RECT 209.115 239.015 209.285 239.185 ;
        RECT 209.115 238.655 209.285 238.825 ;
        RECT 209.115 238.295 209.285 238.465 ;
        RECT 209.115 237.935 209.285 238.105 ;
        RECT 209.115 237.575 209.285 237.745 ;
        RECT 209.115 237.215 209.285 237.385 ;
        RECT 213.695 243.335 213.865 243.505 ;
        RECT 213.695 242.975 213.865 243.145 ;
        RECT 213.695 242.615 213.865 242.785 ;
        RECT 213.695 242.255 213.865 242.425 ;
        RECT 213.695 241.895 213.865 242.065 ;
        RECT 213.695 241.535 213.865 241.705 ;
        RECT 213.695 241.175 213.865 241.345 ;
        RECT 213.695 240.815 213.865 240.985 ;
        RECT 213.695 240.455 213.865 240.625 ;
        RECT 213.695 240.095 213.865 240.265 ;
        RECT 213.695 239.735 213.865 239.905 ;
        RECT 213.695 239.375 213.865 239.545 ;
        RECT 213.695 239.015 213.865 239.185 ;
        RECT 213.695 238.655 213.865 238.825 ;
        RECT 213.695 238.295 213.865 238.465 ;
        RECT 213.695 237.935 213.865 238.105 ;
        RECT 213.695 237.575 213.865 237.745 ;
        RECT 213.695 237.215 213.865 237.385 ;
        RECT 218.275 243.335 218.445 243.505 ;
        RECT 218.275 242.975 218.445 243.145 ;
        RECT 218.275 242.615 218.445 242.785 ;
        RECT 218.275 242.255 218.445 242.425 ;
        RECT 218.275 241.895 218.445 242.065 ;
        RECT 218.275 241.535 218.445 241.705 ;
        RECT 218.275 241.175 218.445 241.345 ;
        RECT 218.275 240.815 218.445 240.985 ;
        RECT 218.275 240.455 218.445 240.625 ;
        RECT 218.275 240.095 218.445 240.265 ;
        RECT 218.275 239.735 218.445 239.905 ;
        RECT 218.275 239.375 218.445 239.545 ;
        RECT 218.275 239.015 218.445 239.185 ;
        RECT 218.275 238.655 218.445 238.825 ;
        RECT 218.275 238.295 218.445 238.465 ;
        RECT 218.275 237.935 218.445 238.105 ;
        RECT 218.275 237.575 218.445 237.745 ;
        RECT 218.275 237.215 218.445 237.385 ;
        RECT 222.855 243.335 223.025 243.505 ;
        RECT 222.855 242.975 223.025 243.145 ;
        RECT 222.855 242.615 223.025 242.785 ;
        RECT 222.855 242.255 223.025 242.425 ;
        RECT 222.855 241.895 223.025 242.065 ;
        RECT 222.855 241.535 223.025 241.705 ;
        RECT 222.855 241.175 223.025 241.345 ;
        RECT 222.855 240.815 223.025 240.985 ;
        RECT 222.855 240.455 223.025 240.625 ;
        RECT 222.855 240.095 223.025 240.265 ;
        RECT 222.855 239.735 223.025 239.905 ;
        RECT 222.855 239.375 223.025 239.545 ;
        RECT 222.855 239.015 223.025 239.185 ;
        RECT 222.855 238.655 223.025 238.825 ;
        RECT 222.855 238.295 223.025 238.465 ;
        RECT 222.855 237.935 223.025 238.105 ;
        RECT 222.855 237.575 223.025 237.745 ;
        RECT 222.855 237.215 223.025 237.385 ;
        RECT 227.435 243.335 227.605 243.505 ;
        RECT 227.435 242.975 227.605 243.145 ;
        RECT 227.435 242.615 227.605 242.785 ;
        RECT 227.435 242.255 227.605 242.425 ;
        RECT 227.435 241.895 227.605 242.065 ;
        RECT 227.435 241.535 227.605 241.705 ;
        RECT 227.435 241.175 227.605 241.345 ;
        RECT 227.435 240.815 227.605 240.985 ;
        RECT 227.435 240.455 227.605 240.625 ;
        RECT 227.435 240.095 227.605 240.265 ;
        RECT 227.435 239.735 227.605 239.905 ;
        RECT 227.435 239.375 227.605 239.545 ;
        RECT 227.435 239.015 227.605 239.185 ;
        RECT 227.435 238.655 227.605 238.825 ;
        RECT 227.435 238.295 227.605 238.465 ;
        RECT 227.435 237.935 227.605 238.105 ;
        RECT 227.435 237.575 227.605 237.745 ;
        RECT 227.435 237.215 227.605 237.385 ;
        RECT 232.015 243.335 232.185 243.505 ;
        RECT 232.015 242.975 232.185 243.145 ;
        RECT 232.015 242.615 232.185 242.785 ;
        RECT 232.015 242.255 232.185 242.425 ;
        RECT 232.015 241.895 232.185 242.065 ;
        RECT 232.015 241.535 232.185 241.705 ;
        RECT 232.015 241.175 232.185 241.345 ;
        RECT 232.015 240.815 232.185 240.985 ;
        RECT 232.015 240.455 232.185 240.625 ;
        RECT 232.015 240.095 232.185 240.265 ;
        RECT 232.015 239.735 232.185 239.905 ;
        RECT 232.015 239.375 232.185 239.545 ;
        RECT 232.015 239.015 232.185 239.185 ;
        RECT 232.015 238.655 232.185 238.825 ;
        RECT 232.015 238.295 232.185 238.465 ;
        RECT 232.015 237.935 232.185 238.105 ;
        RECT 232.015 237.575 232.185 237.745 ;
        RECT 232.015 237.215 232.185 237.385 ;
        RECT 236.595 243.335 236.765 243.505 ;
        RECT 236.595 242.975 236.765 243.145 ;
        RECT 236.595 242.615 236.765 242.785 ;
        RECT 236.595 242.255 236.765 242.425 ;
        RECT 236.595 241.895 236.765 242.065 ;
        RECT 236.595 241.535 236.765 241.705 ;
        RECT 236.595 241.175 236.765 241.345 ;
        RECT 236.595 240.815 236.765 240.985 ;
        RECT 236.595 240.455 236.765 240.625 ;
        RECT 236.595 240.095 236.765 240.265 ;
        RECT 236.595 239.735 236.765 239.905 ;
        RECT 236.595 239.375 236.765 239.545 ;
        RECT 236.595 239.015 236.765 239.185 ;
        RECT 236.595 238.655 236.765 238.825 ;
        RECT 236.595 238.295 236.765 238.465 ;
        RECT 236.595 237.935 236.765 238.105 ;
        RECT 236.595 237.575 236.765 237.745 ;
        RECT 236.595 237.215 236.765 237.385 ;
        RECT 241.175 243.335 241.345 243.505 ;
        RECT 241.175 242.975 241.345 243.145 ;
        RECT 241.175 242.615 241.345 242.785 ;
        RECT 241.175 242.255 241.345 242.425 ;
        RECT 241.175 241.895 241.345 242.065 ;
        RECT 241.175 241.535 241.345 241.705 ;
        RECT 241.175 241.175 241.345 241.345 ;
        RECT 241.175 240.815 241.345 240.985 ;
        RECT 241.175 240.455 241.345 240.625 ;
        RECT 241.175 240.095 241.345 240.265 ;
        RECT 241.175 239.735 241.345 239.905 ;
        RECT 241.175 239.375 241.345 239.545 ;
        RECT 241.175 239.015 241.345 239.185 ;
        RECT 241.175 238.655 241.345 238.825 ;
        RECT 241.175 238.295 241.345 238.465 ;
        RECT 241.175 237.935 241.345 238.105 ;
        RECT 241.175 237.575 241.345 237.745 ;
        RECT 241.175 237.215 241.345 237.385 ;
        RECT 245.755 243.335 245.925 243.505 ;
        RECT 245.755 242.975 245.925 243.145 ;
        RECT 245.755 242.615 245.925 242.785 ;
        RECT 245.755 242.255 245.925 242.425 ;
        RECT 245.755 241.895 245.925 242.065 ;
        RECT 245.755 241.535 245.925 241.705 ;
        RECT 245.755 241.175 245.925 241.345 ;
        RECT 245.755 240.815 245.925 240.985 ;
        RECT 245.755 240.455 245.925 240.625 ;
        RECT 245.755 240.095 245.925 240.265 ;
        RECT 245.755 239.735 245.925 239.905 ;
        RECT 245.755 239.375 245.925 239.545 ;
        RECT 245.755 239.015 245.925 239.185 ;
        RECT 245.755 238.655 245.925 238.825 ;
        RECT 245.755 238.295 245.925 238.465 ;
        RECT 245.755 237.935 245.925 238.105 ;
        RECT 245.755 237.575 245.925 237.745 ;
        RECT 245.755 237.215 245.925 237.385 ;
        RECT 250.335 243.335 250.505 243.505 ;
        RECT 250.335 242.975 250.505 243.145 ;
        RECT 250.335 242.615 250.505 242.785 ;
        RECT 250.335 242.255 250.505 242.425 ;
        RECT 250.335 241.895 250.505 242.065 ;
        RECT 250.335 241.535 250.505 241.705 ;
        RECT 250.335 241.175 250.505 241.345 ;
        RECT 250.335 240.815 250.505 240.985 ;
        RECT 250.335 240.455 250.505 240.625 ;
        RECT 250.335 240.095 250.505 240.265 ;
        RECT 250.335 239.735 250.505 239.905 ;
        RECT 250.335 239.375 250.505 239.545 ;
        RECT 250.335 239.015 250.505 239.185 ;
        RECT 250.335 238.655 250.505 238.825 ;
        RECT 250.335 238.295 250.505 238.465 ;
        RECT 250.335 237.935 250.505 238.105 ;
        RECT 250.335 237.575 250.505 237.745 ;
        RECT 250.335 237.215 250.505 237.385 ;
        RECT 254.915 243.335 255.085 243.505 ;
        RECT 254.915 242.975 255.085 243.145 ;
        RECT 254.915 242.615 255.085 242.785 ;
        RECT 254.915 242.255 255.085 242.425 ;
        RECT 254.915 241.895 255.085 242.065 ;
        RECT 254.915 241.535 255.085 241.705 ;
        RECT 254.915 241.175 255.085 241.345 ;
        RECT 254.915 240.815 255.085 240.985 ;
        RECT 254.915 240.455 255.085 240.625 ;
        RECT 254.915 240.095 255.085 240.265 ;
        RECT 254.915 239.735 255.085 239.905 ;
        RECT 254.915 239.375 255.085 239.545 ;
        RECT 254.915 239.015 255.085 239.185 ;
        RECT 254.915 238.655 255.085 238.825 ;
        RECT 254.915 238.295 255.085 238.465 ;
        RECT 254.915 237.935 255.085 238.105 ;
        RECT 254.915 237.575 255.085 237.745 ;
        RECT 254.915 237.215 255.085 237.385 ;
        RECT 259.495 243.335 259.665 243.505 ;
        RECT 259.495 242.975 259.665 243.145 ;
        RECT 259.495 242.615 259.665 242.785 ;
        RECT 259.495 242.255 259.665 242.425 ;
        RECT 259.495 241.895 259.665 242.065 ;
        RECT 259.495 241.535 259.665 241.705 ;
        RECT 259.495 241.175 259.665 241.345 ;
        RECT 259.495 240.815 259.665 240.985 ;
        RECT 259.495 240.455 259.665 240.625 ;
        RECT 259.495 240.095 259.665 240.265 ;
        RECT 259.495 239.735 259.665 239.905 ;
        RECT 259.495 239.375 259.665 239.545 ;
        RECT 259.495 239.015 259.665 239.185 ;
        RECT 259.495 238.655 259.665 238.825 ;
        RECT 259.495 238.295 259.665 238.465 ;
        RECT 259.495 237.935 259.665 238.105 ;
        RECT 259.495 237.575 259.665 237.745 ;
        RECT 259.495 237.215 259.665 237.385 ;
        RECT 30.505 225.875 30.675 226.045 ;
        RECT 32.505 225.875 32.675 226.045 ;
        RECT 34.505 225.875 34.675 226.045 ;
        RECT 36.505 225.875 36.675 226.045 ;
        RECT 38.505 225.875 38.675 226.045 ;
        RECT 40.505 225.875 40.675 226.045 ;
        RECT 42.505 225.875 42.675 226.045 ;
        RECT 44.505 225.875 44.675 226.045 ;
        RECT 46.505 225.875 46.675 226.045 ;
        RECT 48.505 225.875 48.675 226.045 ;
        RECT 50.505 225.875 50.675 226.045 ;
        RECT 52.505 225.875 52.675 226.045 ;
        RECT 54.505 225.875 54.675 226.045 ;
        RECT 56.505 225.875 56.675 226.045 ;
        RECT 58.505 225.875 58.675 226.045 ;
        RECT 60.505 225.875 60.675 226.045 ;
        RECT 62.505 225.875 62.675 226.045 ;
        RECT 64.505 225.875 64.675 226.045 ;
        RECT 71.505 225.875 71.675 226.045 ;
        RECT 76.065 225.875 76.235 226.045 ;
        RECT 78.065 225.875 78.235 226.045 ;
        RECT 80.065 225.875 80.235 226.045 ;
        RECT 82.065 225.875 82.235 226.045 ;
        RECT 84.065 225.875 84.235 226.045 ;
        RECT 86.065 225.875 86.235 226.045 ;
        RECT 88.065 225.875 88.235 226.045 ;
        RECT 90.065 225.875 90.235 226.045 ;
        RECT 92.065 225.875 92.235 226.045 ;
        RECT 94.065 225.875 94.235 226.045 ;
        RECT 96.065 225.875 96.235 226.045 ;
        RECT 98.065 225.875 98.235 226.045 ;
        RECT 100.065 225.875 100.235 226.045 ;
        RECT 102.065 225.875 102.235 226.045 ;
        RECT 104.065 225.875 104.235 226.045 ;
        RECT 106.065 225.875 106.235 226.045 ;
        RECT 108.065 225.875 108.235 226.045 ;
        RECT 110.065 225.875 110.235 226.045 ;
        RECT 112.065 225.875 112.235 226.045 ;
        RECT 114.065 225.875 114.235 226.045 ;
        RECT 116.065 225.875 116.235 226.045 ;
        RECT 118.065 225.875 118.235 226.045 ;
        RECT 120.065 225.875 120.235 226.045 ;
        RECT 122.065 225.875 122.235 226.045 ;
        RECT 124.065 225.875 124.235 226.045 ;
        RECT 126.065 225.875 126.235 226.045 ;
        RECT 128.065 225.875 128.235 226.045 ;
        RECT 130.065 225.875 130.235 226.045 ;
        RECT 132.065 225.875 132.235 226.045 ;
        RECT 134.065 225.875 134.235 226.045 ;
        RECT 136.065 225.875 136.235 226.045 ;
        RECT 138.065 225.875 138.235 226.045 ;
        RECT 140.065 225.875 140.235 226.045 ;
        RECT 142.065 225.875 142.235 226.045 ;
        RECT 144.065 225.875 144.235 226.045 ;
        RECT 146.065 225.875 146.235 226.045 ;
        RECT 148.065 225.875 148.235 226.045 ;
        RECT 150.065 225.875 150.235 226.045 ;
        RECT 152.065 225.875 152.235 226.045 ;
        RECT 154.065 225.875 154.235 226.045 ;
        RECT 156.065 225.875 156.235 226.045 ;
        RECT 158.065 225.875 158.235 226.045 ;
        RECT 160.065 225.875 160.235 226.045 ;
        RECT 162.065 225.875 162.235 226.045 ;
        RECT 164.065 225.875 164.235 226.045 ;
        RECT 166.065 225.875 166.235 226.045 ;
        RECT 168.065 225.875 168.235 226.045 ;
        RECT 170.065 225.875 170.235 226.045 ;
        RECT 172.065 225.875 172.235 226.045 ;
        RECT 174.065 225.875 174.235 226.045 ;
        RECT 176.065 225.875 176.235 226.045 ;
        RECT 178.065 225.875 178.235 226.045 ;
        RECT 180.065 225.875 180.235 226.045 ;
        RECT 182.065 225.875 182.235 226.045 ;
        RECT 184.065 225.875 184.235 226.045 ;
        RECT 186.065 225.875 186.235 226.045 ;
        RECT 188.065 225.875 188.235 226.045 ;
        RECT 190.065 225.875 190.235 226.045 ;
        RECT 192.065 225.875 192.235 226.045 ;
        RECT 194.065 225.875 194.235 226.045 ;
        RECT 196.065 225.875 196.235 226.045 ;
        RECT 198.065 225.875 198.235 226.045 ;
        RECT 200.065 225.875 200.235 226.045 ;
        RECT 202.065 225.875 202.235 226.045 ;
        RECT 204.065 225.875 204.235 226.045 ;
        RECT 206.065 225.875 206.235 226.045 ;
        RECT 208.065 225.875 208.235 226.045 ;
        RECT 210.065 225.875 210.235 226.045 ;
        RECT 212.065 225.875 212.235 226.045 ;
        RECT 215.715 225.875 215.885 226.045 ;
        RECT 216.715 225.875 216.885 226.045 ;
        RECT 217.715 225.875 217.885 226.045 ;
        RECT 218.715 225.875 218.885 226.045 ;
        RECT 219.715 225.875 219.885 226.045 ;
        RECT 220.715 225.875 220.885 226.045 ;
        RECT 221.715 225.875 221.885 226.045 ;
        RECT 222.715 225.875 222.885 226.045 ;
        RECT 223.715 225.875 223.885 226.045 ;
        RECT 224.715 225.875 224.885 226.045 ;
        RECT 225.715 225.875 225.885 226.045 ;
        RECT 226.715 225.875 226.885 226.045 ;
        RECT 227.715 225.875 227.885 226.045 ;
        RECT 228.715 225.875 228.885 226.045 ;
        RECT 229.715 225.875 229.885 226.045 ;
        RECT 230.715 225.875 230.885 226.045 ;
        RECT 231.715 225.875 231.885 226.045 ;
        RECT 232.715 225.875 232.885 226.045 ;
        RECT 233.715 225.875 233.885 226.045 ;
        RECT 234.715 225.875 234.885 226.045 ;
        RECT 235.715 225.875 235.885 226.045 ;
        RECT 236.715 225.875 236.885 226.045 ;
        RECT 237.715 225.875 237.885 226.045 ;
        RECT 238.715 225.875 238.885 226.045 ;
        RECT 239.715 225.875 239.885 226.045 ;
        RECT 240.715 225.875 240.885 226.045 ;
        RECT 241.715 225.875 241.885 226.045 ;
        RECT 242.715 225.875 242.885 226.045 ;
        RECT 243.715 225.875 243.885 226.045 ;
        RECT 244.715 225.875 244.885 226.045 ;
        RECT 245.715 225.875 245.885 226.045 ;
        RECT 246.715 225.875 246.885 226.045 ;
        RECT 247.715 225.875 247.885 226.045 ;
        RECT 248.715 225.875 248.885 226.045 ;
        RECT 249.715 225.875 249.885 226.045 ;
        RECT 250.715 225.875 250.885 226.045 ;
        RECT 251.715 225.875 251.885 226.045 ;
        RECT 252.715 225.875 252.885 226.045 ;
        RECT 253.715 225.875 253.885 226.045 ;
        RECT 254.715 225.875 254.885 226.045 ;
        RECT 255.715 225.875 255.885 226.045 ;
        RECT 256.715 225.875 256.885 226.045 ;
        RECT 257.715 225.875 257.885 226.045 ;
        RECT 258.715 225.875 258.885 226.045 ;
        RECT 259.715 225.875 259.885 226.045 ;
        RECT 260.715 225.875 260.885 226.045 ;
        RECT 77.675 224.535 77.845 224.705 ;
        RECT 77.675 224.175 77.845 224.345 ;
        RECT 77.675 223.815 77.845 223.985 ;
        RECT 77.675 223.455 77.845 223.625 ;
        RECT 77.675 223.095 77.845 223.265 ;
        RECT 77.675 222.735 77.845 222.905 ;
        RECT 77.675 222.375 77.845 222.545 ;
        RECT 77.675 222.015 77.845 222.185 ;
        RECT 77.675 221.655 77.845 221.825 ;
        RECT 77.675 221.295 77.845 221.465 ;
        RECT 77.675 220.935 77.845 221.105 ;
        RECT 77.675 220.575 77.845 220.745 ;
        RECT 77.675 220.215 77.845 220.385 ;
        RECT 77.675 219.855 77.845 220.025 ;
        RECT 77.675 219.495 77.845 219.665 ;
        RECT 77.675 219.135 77.845 219.305 ;
        RECT 77.675 218.775 77.845 218.945 ;
        RECT 77.675 218.415 77.845 218.585 ;
        RECT 82.255 224.535 82.425 224.705 ;
        RECT 82.255 224.175 82.425 224.345 ;
        RECT 82.255 223.815 82.425 223.985 ;
        RECT 82.255 223.455 82.425 223.625 ;
        RECT 82.255 223.095 82.425 223.265 ;
        RECT 82.255 222.735 82.425 222.905 ;
        RECT 82.255 222.375 82.425 222.545 ;
        RECT 82.255 222.015 82.425 222.185 ;
        RECT 82.255 221.655 82.425 221.825 ;
        RECT 82.255 221.295 82.425 221.465 ;
        RECT 82.255 220.935 82.425 221.105 ;
        RECT 82.255 220.575 82.425 220.745 ;
        RECT 82.255 220.215 82.425 220.385 ;
        RECT 82.255 219.855 82.425 220.025 ;
        RECT 82.255 219.495 82.425 219.665 ;
        RECT 82.255 219.135 82.425 219.305 ;
        RECT 82.255 218.775 82.425 218.945 ;
        RECT 82.255 218.415 82.425 218.585 ;
        RECT 86.835 224.535 87.005 224.705 ;
        RECT 86.835 224.175 87.005 224.345 ;
        RECT 86.835 223.815 87.005 223.985 ;
        RECT 86.835 223.455 87.005 223.625 ;
        RECT 86.835 223.095 87.005 223.265 ;
        RECT 86.835 222.735 87.005 222.905 ;
        RECT 86.835 222.375 87.005 222.545 ;
        RECT 86.835 222.015 87.005 222.185 ;
        RECT 86.835 221.655 87.005 221.825 ;
        RECT 86.835 221.295 87.005 221.465 ;
        RECT 86.835 220.935 87.005 221.105 ;
        RECT 86.835 220.575 87.005 220.745 ;
        RECT 86.835 220.215 87.005 220.385 ;
        RECT 86.835 219.855 87.005 220.025 ;
        RECT 86.835 219.495 87.005 219.665 ;
        RECT 86.835 219.135 87.005 219.305 ;
        RECT 86.835 218.775 87.005 218.945 ;
        RECT 86.835 218.415 87.005 218.585 ;
        RECT 91.415 224.535 91.585 224.705 ;
        RECT 91.415 224.175 91.585 224.345 ;
        RECT 91.415 223.815 91.585 223.985 ;
        RECT 91.415 223.455 91.585 223.625 ;
        RECT 91.415 223.095 91.585 223.265 ;
        RECT 91.415 222.735 91.585 222.905 ;
        RECT 91.415 222.375 91.585 222.545 ;
        RECT 91.415 222.015 91.585 222.185 ;
        RECT 91.415 221.655 91.585 221.825 ;
        RECT 91.415 221.295 91.585 221.465 ;
        RECT 91.415 220.935 91.585 221.105 ;
        RECT 91.415 220.575 91.585 220.745 ;
        RECT 91.415 220.215 91.585 220.385 ;
        RECT 91.415 219.855 91.585 220.025 ;
        RECT 91.415 219.495 91.585 219.665 ;
        RECT 91.415 219.135 91.585 219.305 ;
        RECT 91.415 218.775 91.585 218.945 ;
        RECT 91.415 218.415 91.585 218.585 ;
        RECT 95.995 224.535 96.165 224.705 ;
        RECT 95.995 224.175 96.165 224.345 ;
        RECT 95.995 223.815 96.165 223.985 ;
        RECT 95.995 223.455 96.165 223.625 ;
        RECT 95.995 223.095 96.165 223.265 ;
        RECT 95.995 222.735 96.165 222.905 ;
        RECT 95.995 222.375 96.165 222.545 ;
        RECT 95.995 222.015 96.165 222.185 ;
        RECT 95.995 221.655 96.165 221.825 ;
        RECT 95.995 221.295 96.165 221.465 ;
        RECT 95.995 220.935 96.165 221.105 ;
        RECT 95.995 220.575 96.165 220.745 ;
        RECT 95.995 220.215 96.165 220.385 ;
        RECT 95.995 219.855 96.165 220.025 ;
        RECT 95.995 219.495 96.165 219.665 ;
        RECT 95.995 219.135 96.165 219.305 ;
        RECT 95.995 218.775 96.165 218.945 ;
        RECT 95.995 218.415 96.165 218.585 ;
        RECT 100.575 224.535 100.745 224.705 ;
        RECT 100.575 224.175 100.745 224.345 ;
        RECT 100.575 223.815 100.745 223.985 ;
        RECT 100.575 223.455 100.745 223.625 ;
        RECT 100.575 223.095 100.745 223.265 ;
        RECT 100.575 222.735 100.745 222.905 ;
        RECT 100.575 222.375 100.745 222.545 ;
        RECT 100.575 222.015 100.745 222.185 ;
        RECT 100.575 221.655 100.745 221.825 ;
        RECT 100.575 221.295 100.745 221.465 ;
        RECT 100.575 220.935 100.745 221.105 ;
        RECT 100.575 220.575 100.745 220.745 ;
        RECT 100.575 220.215 100.745 220.385 ;
        RECT 100.575 219.855 100.745 220.025 ;
        RECT 100.575 219.495 100.745 219.665 ;
        RECT 100.575 219.135 100.745 219.305 ;
        RECT 100.575 218.775 100.745 218.945 ;
        RECT 100.575 218.415 100.745 218.585 ;
        RECT 105.155 224.535 105.325 224.705 ;
        RECT 105.155 224.175 105.325 224.345 ;
        RECT 105.155 223.815 105.325 223.985 ;
        RECT 105.155 223.455 105.325 223.625 ;
        RECT 105.155 223.095 105.325 223.265 ;
        RECT 105.155 222.735 105.325 222.905 ;
        RECT 105.155 222.375 105.325 222.545 ;
        RECT 105.155 222.015 105.325 222.185 ;
        RECT 105.155 221.655 105.325 221.825 ;
        RECT 105.155 221.295 105.325 221.465 ;
        RECT 105.155 220.935 105.325 221.105 ;
        RECT 105.155 220.575 105.325 220.745 ;
        RECT 105.155 220.215 105.325 220.385 ;
        RECT 105.155 219.855 105.325 220.025 ;
        RECT 105.155 219.495 105.325 219.665 ;
        RECT 105.155 219.135 105.325 219.305 ;
        RECT 105.155 218.775 105.325 218.945 ;
        RECT 105.155 218.415 105.325 218.585 ;
        RECT 109.735 224.535 109.905 224.705 ;
        RECT 109.735 224.175 109.905 224.345 ;
        RECT 109.735 223.815 109.905 223.985 ;
        RECT 109.735 223.455 109.905 223.625 ;
        RECT 109.735 223.095 109.905 223.265 ;
        RECT 109.735 222.735 109.905 222.905 ;
        RECT 109.735 222.375 109.905 222.545 ;
        RECT 109.735 222.015 109.905 222.185 ;
        RECT 109.735 221.655 109.905 221.825 ;
        RECT 109.735 221.295 109.905 221.465 ;
        RECT 109.735 220.935 109.905 221.105 ;
        RECT 109.735 220.575 109.905 220.745 ;
        RECT 109.735 220.215 109.905 220.385 ;
        RECT 109.735 219.855 109.905 220.025 ;
        RECT 109.735 219.495 109.905 219.665 ;
        RECT 109.735 219.135 109.905 219.305 ;
        RECT 109.735 218.775 109.905 218.945 ;
        RECT 109.735 218.415 109.905 218.585 ;
        RECT 114.315 224.535 114.485 224.705 ;
        RECT 114.315 224.175 114.485 224.345 ;
        RECT 114.315 223.815 114.485 223.985 ;
        RECT 114.315 223.455 114.485 223.625 ;
        RECT 114.315 223.095 114.485 223.265 ;
        RECT 114.315 222.735 114.485 222.905 ;
        RECT 114.315 222.375 114.485 222.545 ;
        RECT 114.315 222.015 114.485 222.185 ;
        RECT 114.315 221.655 114.485 221.825 ;
        RECT 114.315 221.295 114.485 221.465 ;
        RECT 114.315 220.935 114.485 221.105 ;
        RECT 114.315 220.575 114.485 220.745 ;
        RECT 114.315 220.215 114.485 220.385 ;
        RECT 114.315 219.855 114.485 220.025 ;
        RECT 114.315 219.495 114.485 219.665 ;
        RECT 114.315 219.135 114.485 219.305 ;
        RECT 114.315 218.775 114.485 218.945 ;
        RECT 114.315 218.415 114.485 218.585 ;
        RECT 118.895 224.535 119.065 224.705 ;
        RECT 118.895 224.175 119.065 224.345 ;
        RECT 118.895 223.815 119.065 223.985 ;
        RECT 118.895 223.455 119.065 223.625 ;
        RECT 118.895 223.095 119.065 223.265 ;
        RECT 118.895 222.735 119.065 222.905 ;
        RECT 118.895 222.375 119.065 222.545 ;
        RECT 118.895 222.015 119.065 222.185 ;
        RECT 118.895 221.655 119.065 221.825 ;
        RECT 118.895 221.295 119.065 221.465 ;
        RECT 118.895 220.935 119.065 221.105 ;
        RECT 118.895 220.575 119.065 220.745 ;
        RECT 118.895 220.215 119.065 220.385 ;
        RECT 118.895 219.855 119.065 220.025 ;
        RECT 118.895 219.495 119.065 219.665 ;
        RECT 118.895 219.135 119.065 219.305 ;
        RECT 118.895 218.775 119.065 218.945 ;
        RECT 118.895 218.415 119.065 218.585 ;
        RECT 123.475 224.535 123.645 224.705 ;
        RECT 123.475 224.175 123.645 224.345 ;
        RECT 123.475 223.815 123.645 223.985 ;
        RECT 123.475 223.455 123.645 223.625 ;
        RECT 123.475 223.095 123.645 223.265 ;
        RECT 123.475 222.735 123.645 222.905 ;
        RECT 123.475 222.375 123.645 222.545 ;
        RECT 123.475 222.015 123.645 222.185 ;
        RECT 123.475 221.655 123.645 221.825 ;
        RECT 123.475 221.295 123.645 221.465 ;
        RECT 123.475 220.935 123.645 221.105 ;
        RECT 123.475 220.575 123.645 220.745 ;
        RECT 123.475 220.215 123.645 220.385 ;
        RECT 123.475 219.855 123.645 220.025 ;
        RECT 123.475 219.495 123.645 219.665 ;
        RECT 123.475 219.135 123.645 219.305 ;
        RECT 123.475 218.775 123.645 218.945 ;
        RECT 123.475 218.415 123.645 218.585 ;
        RECT 128.055 224.535 128.225 224.705 ;
        RECT 128.055 224.175 128.225 224.345 ;
        RECT 128.055 223.815 128.225 223.985 ;
        RECT 128.055 223.455 128.225 223.625 ;
        RECT 128.055 223.095 128.225 223.265 ;
        RECT 128.055 222.735 128.225 222.905 ;
        RECT 128.055 222.375 128.225 222.545 ;
        RECT 128.055 222.015 128.225 222.185 ;
        RECT 128.055 221.655 128.225 221.825 ;
        RECT 128.055 221.295 128.225 221.465 ;
        RECT 128.055 220.935 128.225 221.105 ;
        RECT 128.055 220.575 128.225 220.745 ;
        RECT 128.055 220.215 128.225 220.385 ;
        RECT 128.055 219.855 128.225 220.025 ;
        RECT 128.055 219.495 128.225 219.665 ;
        RECT 128.055 219.135 128.225 219.305 ;
        RECT 128.055 218.775 128.225 218.945 ;
        RECT 128.055 218.415 128.225 218.585 ;
        RECT 132.635 224.535 132.805 224.705 ;
        RECT 132.635 224.175 132.805 224.345 ;
        RECT 132.635 223.815 132.805 223.985 ;
        RECT 132.635 223.455 132.805 223.625 ;
        RECT 132.635 223.095 132.805 223.265 ;
        RECT 132.635 222.735 132.805 222.905 ;
        RECT 132.635 222.375 132.805 222.545 ;
        RECT 132.635 222.015 132.805 222.185 ;
        RECT 132.635 221.655 132.805 221.825 ;
        RECT 132.635 221.295 132.805 221.465 ;
        RECT 132.635 220.935 132.805 221.105 ;
        RECT 132.635 220.575 132.805 220.745 ;
        RECT 132.635 220.215 132.805 220.385 ;
        RECT 132.635 219.855 132.805 220.025 ;
        RECT 132.635 219.495 132.805 219.665 ;
        RECT 132.635 219.135 132.805 219.305 ;
        RECT 132.635 218.775 132.805 218.945 ;
        RECT 132.635 218.415 132.805 218.585 ;
        RECT 137.215 224.535 137.385 224.705 ;
        RECT 137.215 224.175 137.385 224.345 ;
        RECT 137.215 223.815 137.385 223.985 ;
        RECT 137.215 223.455 137.385 223.625 ;
        RECT 137.215 223.095 137.385 223.265 ;
        RECT 137.215 222.735 137.385 222.905 ;
        RECT 137.215 222.375 137.385 222.545 ;
        RECT 137.215 222.015 137.385 222.185 ;
        RECT 137.215 221.655 137.385 221.825 ;
        RECT 137.215 221.295 137.385 221.465 ;
        RECT 137.215 220.935 137.385 221.105 ;
        RECT 137.215 220.575 137.385 220.745 ;
        RECT 137.215 220.215 137.385 220.385 ;
        RECT 137.215 219.855 137.385 220.025 ;
        RECT 137.215 219.495 137.385 219.665 ;
        RECT 137.215 219.135 137.385 219.305 ;
        RECT 137.215 218.775 137.385 218.945 ;
        RECT 137.215 218.415 137.385 218.585 ;
        RECT 141.795 224.535 141.965 224.705 ;
        RECT 141.795 224.175 141.965 224.345 ;
        RECT 141.795 223.815 141.965 223.985 ;
        RECT 141.795 223.455 141.965 223.625 ;
        RECT 141.795 223.095 141.965 223.265 ;
        RECT 141.795 222.735 141.965 222.905 ;
        RECT 141.795 222.375 141.965 222.545 ;
        RECT 141.795 222.015 141.965 222.185 ;
        RECT 141.795 221.655 141.965 221.825 ;
        RECT 141.795 221.295 141.965 221.465 ;
        RECT 141.795 220.935 141.965 221.105 ;
        RECT 141.795 220.575 141.965 220.745 ;
        RECT 141.795 220.215 141.965 220.385 ;
        RECT 141.795 219.855 141.965 220.025 ;
        RECT 141.795 219.495 141.965 219.665 ;
        RECT 141.795 219.135 141.965 219.305 ;
        RECT 141.795 218.775 141.965 218.945 ;
        RECT 141.795 218.415 141.965 218.585 ;
        RECT 146.375 224.535 146.545 224.705 ;
        RECT 146.375 224.175 146.545 224.345 ;
        RECT 146.375 223.815 146.545 223.985 ;
        RECT 146.375 223.455 146.545 223.625 ;
        RECT 146.375 223.095 146.545 223.265 ;
        RECT 146.375 222.735 146.545 222.905 ;
        RECT 146.375 222.375 146.545 222.545 ;
        RECT 146.375 222.015 146.545 222.185 ;
        RECT 146.375 221.655 146.545 221.825 ;
        RECT 146.375 221.295 146.545 221.465 ;
        RECT 146.375 220.935 146.545 221.105 ;
        RECT 146.375 220.575 146.545 220.745 ;
        RECT 146.375 220.215 146.545 220.385 ;
        RECT 146.375 219.855 146.545 220.025 ;
        RECT 146.375 219.495 146.545 219.665 ;
        RECT 146.375 219.135 146.545 219.305 ;
        RECT 146.375 218.775 146.545 218.945 ;
        RECT 146.375 218.415 146.545 218.585 ;
        RECT 150.955 224.535 151.125 224.705 ;
        RECT 150.955 224.175 151.125 224.345 ;
        RECT 150.955 223.815 151.125 223.985 ;
        RECT 150.955 223.455 151.125 223.625 ;
        RECT 150.955 223.095 151.125 223.265 ;
        RECT 150.955 222.735 151.125 222.905 ;
        RECT 150.955 222.375 151.125 222.545 ;
        RECT 150.955 222.015 151.125 222.185 ;
        RECT 150.955 221.655 151.125 221.825 ;
        RECT 150.955 221.295 151.125 221.465 ;
        RECT 150.955 220.935 151.125 221.105 ;
        RECT 150.955 220.575 151.125 220.745 ;
        RECT 150.955 220.215 151.125 220.385 ;
        RECT 150.955 219.855 151.125 220.025 ;
        RECT 150.955 219.495 151.125 219.665 ;
        RECT 150.955 219.135 151.125 219.305 ;
        RECT 150.955 218.775 151.125 218.945 ;
        RECT 150.955 218.415 151.125 218.585 ;
        RECT 155.535 224.535 155.705 224.705 ;
        RECT 155.535 224.175 155.705 224.345 ;
        RECT 155.535 223.815 155.705 223.985 ;
        RECT 155.535 223.455 155.705 223.625 ;
        RECT 155.535 223.095 155.705 223.265 ;
        RECT 155.535 222.735 155.705 222.905 ;
        RECT 155.535 222.375 155.705 222.545 ;
        RECT 155.535 222.015 155.705 222.185 ;
        RECT 155.535 221.655 155.705 221.825 ;
        RECT 155.535 221.295 155.705 221.465 ;
        RECT 155.535 220.935 155.705 221.105 ;
        RECT 155.535 220.575 155.705 220.745 ;
        RECT 155.535 220.215 155.705 220.385 ;
        RECT 155.535 219.855 155.705 220.025 ;
        RECT 155.535 219.495 155.705 219.665 ;
        RECT 155.535 219.135 155.705 219.305 ;
        RECT 155.535 218.775 155.705 218.945 ;
        RECT 155.535 218.415 155.705 218.585 ;
        RECT 160.115 224.535 160.285 224.705 ;
        RECT 160.115 224.175 160.285 224.345 ;
        RECT 160.115 223.815 160.285 223.985 ;
        RECT 160.115 223.455 160.285 223.625 ;
        RECT 160.115 223.095 160.285 223.265 ;
        RECT 160.115 222.735 160.285 222.905 ;
        RECT 160.115 222.375 160.285 222.545 ;
        RECT 160.115 222.015 160.285 222.185 ;
        RECT 160.115 221.655 160.285 221.825 ;
        RECT 160.115 221.295 160.285 221.465 ;
        RECT 160.115 220.935 160.285 221.105 ;
        RECT 160.115 220.575 160.285 220.745 ;
        RECT 160.115 220.215 160.285 220.385 ;
        RECT 160.115 219.855 160.285 220.025 ;
        RECT 160.115 219.495 160.285 219.665 ;
        RECT 160.115 219.135 160.285 219.305 ;
        RECT 160.115 218.775 160.285 218.945 ;
        RECT 160.115 218.415 160.285 218.585 ;
        RECT 164.695 224.535 164.865 224.705 ;
        RECT 164.695 224.175 164.865 224.345 ;
        RECT 164.695 223.815 164.865 223.985 ;
        RECT 164.695 223.455 164.865 223.625 ;
        RECT 164.695 223.095 164.865 223.265 ;
        RECT 164.695 222.735 164.865 222.905 ;
        RECT 164.695 222.375 164.865 222.545 ;
        RECT 164.695 222.015 164.865 222.185 ;
        RECT 164.695 221.655 164.865 221.825 ;
        RECT 164.695 221.295 164.865 221.465 ;
        RECT 164.695 220.935 164.865 221.105 ;
        RECT 164.695 220.575 164.865 220.745 ;
        RECT 164.695 220.215 164.865 220.385 ;
        RECT 164.695 219.855 164.865 220.025 ;
        RECT 164.695 219.495 164.865 219.665 ;
        RECT 164.695 219.135 164.865 219.305 ;
        RECT 164.695 218.775 164.865 218.945 ;
        RECT 164.695 218.415 164.865 218.585 ;
        RECT 169.275 224.535 169.445 224.705 ;
        RECT 169.275 224.175 169.445 224.345 ;
        RECT 169.275 223.815 169.445 223.985 ;
        RECT 169.275 223.455 169.445 223.625 ;
        RECT 169.275 223.095 169.445 223.265 ;
        RECT 169.275 222.735 169.445 222.905 ;
        RECT 169.275 222.375 169.445 222.545 ;
        RECT 169.275 222.015 169.445 222.185 ;
        RECT 169.275 221.655 169.445 221.825 ;
        RECT 169.275 221.295 169.445 221.465 ;
        RECT 169.275 220.935 169.445 221.105 ;
        RECT 169.275 220.575 169.445 220.745 ;
        RECT 169.275 220.215 169.445 220.385 ;
        RECT 169.275 219.855 169.445 220.025 ;
        RECT 169.275 219.495 169.445 219.665 ;
        RECT 169.275 219.135 169.445 219.305 ;
        RECT 169.275 218.775 169.445 218.945 ;
        RECT 169.275 218.415 169.445 218.585 ;
        RECT 173.855 224.535 174.025 224.705 ;
        RECT 173.855 224.175 174.025 224.345 ;
        RECT 173.855 223.815 174.025 223.985 ;
        RECT 173.855 223.455 174.025 223.625 ;
        RECT 173.855 223.095 174.025 223.265 ;
        RECT 173.855 222.735 174.025 222.905 ;
        RECT 173.855 222.375 174.025 222.545 ;
        RECT 173.855 222.015 174.025 222.185 ;
        RECT 173.855 221.655 174.025 221.825 ;
        RECT 173.855 221.295 174.025 221.465 ;
        RECT 173.855 220.935 174.025 221.105 ;
        RECT 173.855 220.575 174.025 220.745 ;
        RECT 173.855 220.215 174.025 220.385 ;
        RECT 173.855 219.855 174.025 220.025 ;
        RECT 173.855 219.495 174.025 219.665 ;
        RECT 173.855 219.135 174.025 219.305 ;
        RECT 173.855 218.775 174.025 218.945 ;
        RECT 173.855 218.415 174.025 218.585 ;
        RECT 178.435 224.535 178.605 224.705 ;
        RECT 178.435 224.175 178.605 224.345 ;
        RECT 178.435 223.815 178.605 223.985 ;
        RECT 178.435 223.455 178.605 223.625 ;
        RECT 178.435 223.095 178.605 223.265 ;
        RECT 178.435 222.735 178.605 222.905 ;
        RECT 178.435 222.375 178.605 222.545 ;
        RECT 178.435 222.015 178.605 222.185 ;
        RECT 178.435 221.655 178.605 221.825 ;
        RECT 178.435 221.295 178.605 221.465 ;
        RECT 178.435 220.935 178.605 221.105 ;
        RECT 178.435 220.575 178.605 220.745 ;
        RECT 178.435 220.215 178.605 220.385 ;
        RECT 178.435 219.855 178.605 220.025 ;
        RECT 178.435 219.495 178.605 219.665 ;
        RECT 178.435 219.135 178.605 219.305 ;
        RECT 178.435 218.775 178.605 218.945 ;
        RECT 178.435 218.415 178.605 218.585 ;
        RECT 183.015 224.535 183.185 224.705 ;
        RECT 183.015 224.175 183.185 224.345 ;
        RECT 183.015 223.815 183.185 223.985 ;
        RECT 183.015 223.455 183.185 223.625 ;
        RECT 183.015 223.095 183.185 223.265 ;
        RECT 183.015 222.735 183.185 222.905 ;
        RECT 183.015 222.375 183.185 222.545 ;
        RECT 183.015 222.015 183.185 222.185 ;
        RECT 183.015 221.655 183.185 221.825 ;
        RECT 183.015 221.295 183.185 221.465 ;
        RECT 183.015 220.935 183.185 221.105 ;
        RECT 183.015 220.575 183.185 220.745 ;
        RECT 183.015 220.215 183.185 220.385 ;
        RECT 183.015 219.855 183.185 220.025 ;
        RECT 183.015 219.495 183.185 219.665 ;
        RECT 183.015 219.135 183.185 219.305 ;
        RECT 183.015 218.775 183.185 218.945 ;
        RECT 183.015 218.415 183.185 218.585 ;
        RECT 187.595 224.535 187.765 224.705 ;
        RECT 187.595 224.175 187.765 224.345 ;
        RECT 187.595 223.815 187.765 223.985 ;
        RECT 187.595 223.455 187.765 223.625 ;
        RECT 187.595 223.095 187.765 223.265 ;
        RECT 187.595 222.735 187.765 222.905 ;
        RECT 187.595 222.375 187.765 222.545 ;
        RECT 187.595 222.015 187.765 222.185 ;
        RECT 187.595 221.655 187.765 221.825 ;
        RECT 187.595 221.295 187.765 221.465 ;
        RECT 187.595 220.935 187.765 221.105 ;
        RECT 187.595 220.575 187.765 220.745 ;
        RECT 187.595 220.215 187.765 220.385 ;
        RECT 187.595 219.855 187.765 220.025 ;
        RECT 187.595 219.495 187.765 219.665 ;
        RECT 187.595 219.135 187.765 219.305 ;
        RECT 187.595 218.775 187.765 218.945 ;
        RECT 187.595 218.415 187.765 218.585 ;
        RECT 192.175 224.535 192.345 224.705 ;
        RECT 192.175 224.175 192.345 224.345 ;
        RECT 192.175 223.815 192.345 223.985 ;
        RECT 192.175 223.455 192.345 223.625 ;
        RECT 192.175 223.095 192.345 223.265 ;
        RECT 192.175 222.735 192.345 222.905 ;
        RECT 192.175 222.375 192.345 222.545 ;
        RECT 192.175 222.015 192.345 222.185 ;
        RECT 192.175 221.655 192.345 221.825 ;
        RECT 192.175 221.295 192.345 221.465 ;
        RECT 192.175 220.935 192.345 221.105 ;
        RECT 192.175 220.575 192.345 220.745 ;
        RECT 192.175 220.215 192.345 220.385 ;
        RECT 192.175 219.855 192.345 220.025 ;
        RECT 192.175 219.495 192.345 219.665 ;
        RECT 192.175 219.135 192.345 219.305 ;
        RECT 192.175 218.775 192.345 218.945 ;
        RECT 192.175 218.415 192.345 218.585 ;
        RECT 196.755 224.535 196.925 224.705 ;
        RECT 196.755 224.175 196.925 224.345 ;
        RECT 196.755 223.815 196.925 223.985 ;
        RECT 196.755 223.455 196.925 223.625 ;
        RECT 196.755 223.095 196.925 223.265 ;
        RECT 196.755 222.735 196.925 222.905 ;
        RECT 196.755 222.375 196.925 222.545 ;
        RECT 196.755 222.015 196.925 222.185 ;
        RECT 196.755 221.655 196.925 221.825 ;
        RECT 196.755 221.295 196.925 221.465 ;
        RECT 196.755 220.935 196.925 221.105 ;
        RECT 196.755 220.575 196.925 220.745 ;
        RECT 196.755 220.215 196.925 220.385 ;
        RECT 196.755 219.855 196.925 220.025 ;
        RECT 196.755 219.495 196.925 219.665 ;
        RECT 196.755 219.135 196.925 219.305 ;
        RECT 196.755 218.775 196.925 218.945 ;
        RECT 196.755 218.415 196.925 218.585 ;
        RECT 201.335 224.535 201.505 224.705 ;
        RECT 201.335 224.175 201.505 224.345 ;
        RECT 201.335 223.815 201.505 223.985 ;
        RECT 201.335 223.455 201.505 223.625 ;
        RECT 201.335 223.095 201.505 223.265 ;
        RECT 201.335 222.735 201.505 222.905 ;
        RECT 201.335 222.375 201.505 222.545 ;
        RECT 201.335 222.015 201.505 222.185 ;
        RECT 201.335 221.655 201.505 221.825 ;
        RECT 201.335 221.295 201.505 221.465 ;
        RECT 201.335 220.935 201.505 221.105 ;
        RECT 201.335 220.575 201.505 220.745 ;
        RECT 201.335 220.215 201.505 220.385 ;
        RECT 201.335 219.855 201.505 220.025 ;
        RECT 201.335 219.495 201.505 219.665 ;
        RECT 201.335 219.135 201.505 219.305 ;
        RECT 201.335 218.775 201.505 218.945 ;
        RECT 201.335 218.415 201.505 218.585 ;
        RECT 205.915 224.535 206.085 224.705 ;
        RECT 205.915 224.175 206.085 224.345 ;
        RECT 205.915 223.815 206.085 223.985 ;
        RECT 205.915 223.455 206.085 223.625 ;
        RECT 205.915 223.095 206.085 223.265 ;
        RECT 205.915 222.735 206.085 222.905 ;
        RECT 205.915 222.375 206.085 222.545 ;
        RECT 205.915 222.015 206.085 222.185 ;
        RECT 205.915 221.655 206.085 221.825 ;
        RECT 205.915 221.295 206.085 221.465 ;
        RECT 205.915 220.935 206.085 221.105 ;
        RECT 205.915 220.575 206.085 220.745 ;
        RECT 205.915 220.215 206.085 220.385 ;
        RECT 205.915 219.855 206.085 220.025 ;
        RECT 205.915 219.495 206.085 219.665 ;
        RECT 205.915 219.135 206.085 219.305 ;
        RECT 205.915 218.775 206.085 218.945 ;
        RECT 205.915 218.415 206.085 218.585 ;
        RECT 210.495 224.535 210.665 224.705 ;
        RECT 210.495 224.175 210.665 224.345 ;
        RECT 210.495 223.815 210.665 223.985 ;
        RECT 210.495 223.455 210.665 223.625 ;
        RECT 210.495 223.095 210.665 223.265 ;
        RECT 210.495 222.735 210.665 222.905 ;
        RECT 210.495 222.375 210.665 222.545 ;
        RECT 210.495 222.015 210.665 222.185 ;
        RECT 210.495 221.655 210.665 221.825 ;
        RECT 210.495 221.295 210.665 221.465 ;
        RECT 210.495 220.935 210.665 221.105 ;
        RECT 210.495 220.575 210.665 220.745 ;
        RECT 210.495 220.215 210.665 220.385 ;
        RECT 210.495 219.855 210.665 220.025 ;
        RECT 210.495 219.495 210.665 219.665 ;
        RECT 210.495 219.135 210.665 219.305 ;
        RECT 210.495 218.775 210.665 218.945 ;
        RECT 210.495 218.415 210.665 218.585 ;
        RECT 32.465 207.075 32.635 207.245 ;
        RECT 34.465 207.075 34.635 207.245 ;
        RECT 36.465 207.075 36.635 207.245 ;
        RECT 38.465 207.075 38.635 207.245 ;
        RECT 40.465 207.075 40.635 207.245 ;
        RECT 42.465 207.075 42.635 207.245 ;
        RECT 44.465 207.075 44.635 207.245 ;
        RECT 46.465 207.075 46.635 207.245 ;
        RECT 48.465 207.075 48.635 207.245 ;
        RECT 50.465 207.075 50.635 207.245 ;
        RECT 52.465 207.075 52.635 207.245 ;
        RECT 54.465 207.075 54.635 207.245 ;
        RECT 56.465 207.075 56.635 207.245 ;
        RECT 58.465 207.075 58.635 207.245 ;
        RECT 60.465 207.075 60.635 207.245 ;
        RECT 62.465 207.075 62.635 207.245 ;
        RECT 64.465 207.075 64.635 207.245 ;
        RECT 66.465 207.075 66.635 207.245 ;
        RECT 76.565 207.075 76.735 207.245 ;
        RECT 78.565 207.075 78.735 207.245 ;
        RECT 80.565 207.075 80.735 207.245 ;
        RECT 82.565 207.075 82.735 207.245 ;
        RECT 84.565 207.075 84.735 207.245 ;
        RECT 86.565 207.075 86.735 207.245 ;
        RECT 88.565 207.075 88.735 207.245 ;
        RECT 90.565 207.075 90.735 207.245 ;
        RECT 92.565 207.075 92.735 207.245 ;
        RECT 94.565 207.075 94.735 207.245 ;
        RECT 96.565 207.075 96.735 207.245 ;
        RECT 98.565 207.075 98.735 207.245 ;
        RECT 100.565 207.075 100.735 207.245 ;
        RECT 102.565 207.075 102.735 207.245 ;
        RECT 104.565 207.075 104.735 207.245 ;
        RECT 106.565 207.075 106.735 207.245 ;
        RECT 108.565 207.075 108.735 207.245 ;
        RECT 110.565 207.075 110.735 207.245 ;
        RECT 114.285 207.075 114.455 207.245 ;
        RECT 116.285 207.075 116.455 207.245 ;
        RECT 118.285 207.075 118.455 207.245 ;
        RECT 120.285 207.075 120.455 207.245 ;
        RECT 122.285 207.075 122.455 207.245 ;
        RECT 124.285 207.075 124.455 207.245 ;
        RECT 126.285 207.075 126.455 207.245 ;
        RECT 128.285 207.075 128.455 207.245 ;
        RECT 130.285 207.075 130.455 207.245 ;
        RECT 132.285 207.075 132.455 207.245 ;
        RECT 134.285 207.075 134.455 207.245 ;
        RECT 136.285 207.075 136.455 207.245 ;
        RECT 138.285 207.075 138.455 207.245 ;
        RECT 140.285 207.075 140.455 207.245 ;
        RECT 147.605 207.075 147.775 207.245 ;
        RECT 149.605 207.075 149.775 207.245 ;
        RECT 151.605 207.075 151.775 207.245 ;
        RECT 153.605 207.075 153.775 207.245 ;
        RECT 155.605 207.075 155.775 207.245 ;
        RECT 157.605 207.075 157.775 207.245 ;
        RECT 159.605 207.075 159.775 207.245 ;
        RECT 161.605 207.075 161.775 207.245 ;
        RECT 163.605 207.075 163.775 207.245 ;
        RECT 165.605 207.075 165.775 207.245 ;
        RECT 167.605 207.075 167.775 207.245 ;
        RECT 169.605 207.075 169.775 207.245 ;
        RECT 171.605 207.075 171.775 207.245 ;
        RECT 173.605 207.075 173.775 207.245 ;
        RECT 187.295 207.075 187.465 207.245 ;
        RECT 189.295 207.075 189.465 207.245 ;
        RECT 191.295 207.075 191.465 207.245 ;
        RECT 193.295 207.075 193.465 207.245 ;
        RECT 195.295 207.075 195.465 207.245 ;
        RECT 197.295 207.075 197.465 207.245 ;
        RECT 199.295 207.075 199.465 207.245 ;
        RECT 201.295 207.075 201.465 207.245 ;
        RECT 203.295 207.075 203.465 207.245 ;
        RECT 205.295 207.075 205.465 207.245 ;
        RECT 209.835 207.075 210.005 207.245 ;
        RECT 210.835 207.075 211.005 207.245 ;
        RECT 211.835 207.075 212.005 207.245 ;
        RECT 212.835 207.075 213.005 207.245 ;
        RECT 213.835 207.075 214.005 207.245 ;
        RECT 214.835 207.075 215.005 207.245 ;
        RECT 215.835 207.075 216.005 207.245 ;
        RECT 216.835 207.075 217.005 207.245 ;
        RECT 217.835 207.075 218.005 207.245 ;
        RECT 218.835 207.075 219.005 207.245 ;
        RECT 219.835 207.075 220.005 207.245 ;
        RECT 220.835 207.075 221.005 207.245 ;
        RECT 221.835 207.075 222.005 207.245 ;
        RECT 222.835 207.075 223.005 207.245 ;
        RECT 223.835 207.075 224.005 207.245 ;
        RECT 224.835 207.075 225.005 207.245 ;
        RECT 225.835 207.075 226.005 207.245 ;
        RECT 226.835 207.075 227.005 207.245 ;
        RECT 227.835 207.075 228.005 207.245 ;
        RECT 228.835 207.075 229.005 207.245 ;
        RECT 229.835 207.075 230.005 207.245 ;
        RECT 230.835 207.075 231.005 207.245 ;
        RECT 231.835 207.075 232.005 207.245 ;
        RECT 232.835 207.075 233.005 207.245 ;
        RECT 233.835 207.075 234.005 207.245 ;
        RECT 234.835 207.075 235.005 207.245 ;
        RECT 235.835 207.075 236.005 207.245 ;
        RECT 236.835 207.075 237.005 207.245 ;
        RECT 237.835 207.075 238.005 207.245 ;
        RECT 238.835 207.075 239.005 207.245 ;
        RECT 239.835 207.075 240.005 207.245 ;
        RECT 240.835 207.075 241.005 207.245 ;
        RECT 241.835 207.075 242.005 207.245 ;
        RECT 242.835 207.075 243.005 207.245 ;
        RECT 243.835 207.075 244.005 207.245 ;
        RECT 244.835 207.075 245.005 207.245 ;
        RECT 245.835 207.075 246.005 207.245 ;
        RECT 246.835 207.075 247.005 207.245 ;
        RECT 247.835 207.075 248.005 207.245 ;
        RECT 248.835 207.075 249.005 207.245 ;
        RECT 249.835 207.075 250.005 207.245 ;
        RECT 250.835 207.075 251.005 207.245 ;
        RECT 251.835 207.075 252.005 207.245 ;
        RECT 252.835 207.075 253.005 207.245 ;
        RECT 253.835 207.075 254.005 207.245 ;
        RECT 254.835 207.075 255.005 207.245 ;
        RECT 255.835 207.075 256.005 207.245 ;
        RECT 256.835 207.075 257.005 207.245 ;
        RECT 257.835 207.075 258.005 207.245 ;
        RECT 258.835 207.075 259.005 207.245 ;
        RECT 259.835 207.075 260.005 207.245 ;
        RECT 260.835 207.075 261.005 207.245 ;
        RECT 261.835 207.075 262.005 207.245 ;
        RECT 115.895 205.735 116.065 205.905 ;
        RECT 115.895 205.375 116.065 205.545 ;
        RECT 115.895 205.015 116.065 205.185 ;
        RECT 115.895 204.655 116.065 204.825 ;
        RECT 115.895 204.295 116.065 204.465 ;
        RECT 115.895 203.935 116.065 204.105 ;
        RECT 115.895 203.575 116.065 203.745 ;
        RECT 115.895 203.215 116.065 203.385 ;
        RECT 115.895 202.855 116.065 203.025 ;
        RECT 115.895 202.495 116.065 202.665 ;
        RECT 115.895 202.135 116.065 202.305 ;
        RECT 115.895 201.775 116.065 201.945 ;
        RECT 115.895 201.415 116.065 201.585 ;
        RECT 115.895 201.055 116.065 201.225 ;
        RECT 115.895 200.695 116.065 200.865 ;
        RECT 115.895 200.335 116.065 200.505 ;
        RECT 115.895 199.975 116.065 200.145 ;
        RECT 115.895 199.615 116.065 199.785 ;
        RECT 120.475 205.735 120.645 205.905 ;
        RECT 120.475 205.375 120.645 205.545 ;
        RECT 120.475 205.015 120.645 205.185 ;
        RECT 120.475 204.655 120.645 204.825 ;
        RECT 120.475 204.295 120.645 204.465 ;
        RECT 120.475 203.935 120.645 204.105 ;
        RECT 120.475 203.575 120.645 203.745 ;
        RECT 120.475 203.215 120.645 203.385 ;
        RECT 120.475 202.855 120.645 203.025 ;
        RECT 120.475 202.495 120.645 202.665 ;
        RECT 120.475 202.135 120.645 202.305 ;
        RECT 120.475 201.775 120.645 201.945 ;
        RECT 120.475 201.415 120.645 201.585 ;
        RECT 120.475 201.055 120.645 201.225 ;
        RECT 120.475 200.695 120.645 200.865 ;
        RECT 120.475 200.335 120.645 200.505 ;
        RECT 120.475 199.975 120.645 200.145 ;
        RECT 120.475 199.615 120.645 199.785 ;
        RECT 125.055 205.735 125.225 205.905 ;
        RECT 125.055 205.375 125.225 205.545 ;
        RECT 125.055 205.015 125.225 205.185 ;
        RECT 125.055 204.655 125.225 204.825 ;
        RECT 125.055 204.295 125.225 204.465 ;
        RECT 125.055 203.935 125.225 204.105 ;
        RECT 125.055 203.575 125.225 203.745 ;
        RECT 125.055 203.215 125.225 203.385 ;
        RECT 125.055 202.855 125.225 203.025 ;
        RECT 125.055 202.495 125.225 202.665 ;
        RECT 125.055 202.135 125.225 202.305 ;
        RECT 125.055 201.775 125.225 201.945 ;
        RECT 125.055 201.415 125.225 201.585 ;
        RECT 125.055 201.055 125.225 201.225 ;
        RECT 125.055 200.695 125.225 200.865 ;
        RECT 125.055 200.335 125.225 200.505 ;
        RECT 125.055 199.975 125.225 200.145 ;
        RECT 125.055 199.615 125.225 199.785 ;
        RECT 129.635 205.735 129.805 205.905 ;
        RECT 129.635 205.375 129.805 205.545 ;
        RECT 129.635 205.015 129.805 205.185 ;
        RECT 129.635 204.655 129.805 204.825 ;
        RECT 129.635 204.295 129.805 204.465 ;
        RECT 129.635 203.935 129.805 204.105 ;
        RECT 129.635 203.575 129.805 203.745 ;
        RECT 129.635 203.215 129.805 203.385 ;
        RECT 129.635 202.855 129.805 203.025 ;
        RECT 129.635 202.495 129.805 202.665 ;
        RECT 129.635 202.135 129.805 202.305 ;
        RECT 129.635 201.775 129.805 201.945 ;
        RECT 129.635 201.415 129.805 201.585 ;
        RECT 129.635 201.055 129.805 201.225 ;
        RECT 129.635 200.695 129.805 200.865 ;
        RECT 129.635 200.335 129.805 200.505 ;
        RECT 129.635 199.975 129.805 200.145 ;
        RECT 129.635 199.615 129.805 199.785 ;
        RECT 134.215 205.735 134.385 205.905 ;
        RECT 134.215 205.375 134.385 205.545 ;
        RECT 134.215 205.015 134.385 205.185 ;
        RECT 134.215 204.655 134.385 204.825 ;
        RECT 134.215 204.295 134.385 204.465 ;
        RECT 134.215 203.935 134.385 204.105 ;
        RECT 134.215 203.575 134.385 203.745 ;
        RECT 134.215 203.215 134.385 203.385 ;
        RECT 134.215 202.855 134.385 203.025 ;
        RECT 134.215 202.495 134.385 202.665 ;
        RECT 134.215 202.135 134.385 202.305 ;
        RECT 134.215 201.775 134.385 201.945 ;
        RECT 134.215 201.415 134.385 201.585 ;
        RECT 134.215 201.055 134.385 201.225 ;
        RECT 134.215 200.695 134.385 200.865 ;
        RECT 134.215 200.335 134.385 200.505 ;
        RECT 134.215 199.975 134.385 200.145 ;
        RECT 134.215 199.615 134.385 199.785 ;
        RECT 138.795 205.735 138.965 205.905 ;
        RECT 138.795 205.375 138.965 205.545 ;
        RECT 138.795 205.015 138.965 205.185 ;
        RECT 138.795 204.655 138.965 204.825 ;
        RECT 138.795 204.295 138.965 204.465 ;
        RECT 138.795 203.935 138.965 204.105 ;
        RECT 138.795 203.575 138.965 203.745 ;
        RECT 138.795 203.215 138.965 203.385 ;
        RECT 138.795 202.855 138.965 203.025 ;
        RECT 138.795 202.495 138.965 202.665 ;
        RECT 138.795 202.135 138.965 202.305 ;
        RECT 138.795 201.775 138.965 201.945 ;
        RECT 138.795 201.415 138.965 201.585 ;
        RECT 138.795 201.055 138.965 201.225 ;
        RECT 138.795 200.695 138.965 200.865 ;
        RECT 138.795 200.335 138.965 200.505 ;
        RECT 138.795 199.975 138.965 200.145 ;
        RECT 138.795 199.615 138.965 199.785 ;
        RECT 149.215 205.735 149.385 205.905 ;
        RECT 149.215 205.375 149.385 205.545 ;
        RECT 149.215 205.015 149.385 205.185 ;
        RECT 149.215 204.655 149.385 204.825 ;
        RECT 149.215 204.295 149.385 204.465 ;
        RECT 149.215 203.935 149.385 204.105 ;
        RECT 149.215 203.575 149.385 203.745 ;
        RECT 149.215 203.215 149.385 203.385 ;
        RECT 149.215 202.855 149.385 203.025 ;
        RECT 149.215 202.495 149.385 202.665 ;
        RECT 149.215 202.135 149.385 202.305 ;
        RECT 149.215 201.775 149.385 201.945 ;
        RECT 149.215 201.415 149.385 201.585 ;
        RECT 149.215 201.055 149.385 201.225 ;
        RECT 149.215 200.695 149.385 200.865 ;
        RECT 149.215 200.335 149.385 200.505 ;
        RECT 149.215 199.975 149.385 200.145 ;
        RECT 149.215 199.615 149.385 199.785 ;
        RECT 153.795 205.735 153.965 205.905 ;
        RECT 153.795 205.375 153.965 205.545 ;
        RECT 153.795 205.015 153.965 205.185 ;
        RECT 153.795 204.655 153.965 204.825 ;
        RECT 153.795 204.295 153.965 204.465 ;
        RECT 153.795 203.935 153.965 204.105 ;
        RECT 153.795 203.575 153.965 203.745 ;
        RECT 153.795 203.215 153.965 203.385 ;
        RECT 153.795 202.855 153.965 203.025 ;
        RECT 153.795 202.495 153.965 202.665 ;
        RECT 153.795 202.135 153.965 202.305 ;
        RECT 153.795 201.775 153.965 201.945 ;
        RECT 153.795 201.415 153.965 201.585 ;
        RECT 153.795 201.055 153.965 201.225 ;
        RECT 153.795 200.695 153.965 200.865 ;
        RECT 153.795 200.335 153.965 200.505 ;
        RECT 153.795 199.975 153.965 200.145 ;
        RECT 153.795 199.615 153.965 199.785 ;
        RECT 158.375 205.735 158.545 205.905 ;
        RECT 158.375 205.375 158.545 205.545 ;
        RECT 158.375 205.015 158.545 205.185 ;
        RECT 158.375 204.655 158.545 204.825 ;
        RECT 158.375 204.295 158.545 204.465 ;
        RECT 158.375 203.935 158.545 204.105 ;
        RECT 158.375 203.575 158.545 203.745 ;
        RECT 158.375 203.215 158.545 203.385 ;
        RECT 158.375 202.855 158.545 203.025 ;
        RECT 158.375 202.495 158.545 202.665 ;
        RECT 158.375 202.135 158.545 202.305 ;
        RECT 158.375 201.775 158.545 201.945 ;
        RECT 158.375 201.415 158.545 201.585 ;
        RECT 158.375 201.055 158.545 201.225 ;
        RECT 158.375 200.695 158.545 200.865 ;
        RECT 158.375 200.335 158.545 200.505 ;
        RECT 158.375 199.975 158.545 200.145 ;
        RECT 158.375 199.615 158.545 199.785 ;
        RECT 162.955 205.735 163.125 205.905 ;
        RECT 162.955 205.375 163.125 205.545 ;
        RECT 162.955 205.015 163.125 205.185 ;
        RECT 162.955 204.655 163.125 204.825 ;
        RECT 162.955 204.295 163.125 204.465 ;
        RECT 162.955 203.935 163.125 204.105 ;
        RECT 162.955 203.575 163.125 203.745 ;
        RECT 162.955 203.215 163.125 203.385 ;
        RECT 162.955 202.855 163.125 203.025 ;
        RECT 162.955 202.495 163.125 202.665 ;
        RECT 162.955 202.135 163.125 202.305 ;
        RECT 162.955 201.775 163.125 201.945 ;
        RECT 162.955 201.415 163.125 201.585 ;
        RECT 162.955 201.055 163.125 201.225 ;
        RECT 162.955 200.695 163.125 200.865 ;
        RECT 162.955 200.335 163.125 200.505 ;
        RECT 162.955 199.975 163.125 200.145 ;
        RECT 162.955 199.615 163.125 199.785 ;
        RECT 167.535 205.735 167.705 205.905 ;
        RECT 167.535 205.375 167.705 205.545 ;
        RECT 167.535 205.015 167.705 205.185 ;
        RECT 167.535 204.655 167.705 204.825 ;
        RECT 167.535 204.295 167.705 204.465 ;
        RECT 167.535 203.935 167.705 204.105 ;
        RECT 167.535 203.575 167.705 203.745 ;
        RECT 167.535 203.215 167.705 203.385 ;
        RECT 167.535 202.855 167.705 203.025 ;
        RECT 167.535 202.495 167.705 202.665 ;
        RECT 167.535 202.135 167.705 202.305 ;
        RECT 167.535 201.775 167.705 201.945 ;
        RECT 167.535 201.415 167.705 201.585 ;
        RECT 167.535 201.055 167.705 201.225 ;
        RECT 167.535 200.695 167.705 200.865 ;
        RECT 167.535 200.335 167.705 200.505 ;
        RECT 167.535 199.975 167.705 200.145 ;
        RECT 167.535 199.615 167.705 199.785 ;
        RECT 172.115 205.735 172.285 205.905 ;
        RECT 172.115 205.375 172.285 205.545 ;
        RECT 172.115 205.015 172.285 205.185 ;
        RECT 172.115 204.655 172.285 204.825 ;
        RECT 172.115 204.295 172.285 204.465 ;
        RECT 172.115 203.935 172.285 204.105 ;
        RECT 172.115 203.575 172.285 203.745 ;
        RECT 172.115 203.215 172.285 203.385 ;
        RECT 172.115 202.855 172.285 203.025 ;
        RECT 172.115 202.495 172.285 202.665 ;
        RECT 172.115 202.135 172.285 202.305 ;
        RECT 172.115 201.775 172.285 201.945 ;
        RECT 172.115 201.415 172.285 201.585 ;
        RECT 172.115 201.055 172.285 201.225 ;
        RECT 172.115 200.695 172.285 200.865 ;
        RECT 172.115 200.335 172.285 200.505 ;
        RECT 172.115 199.975 172.285 200.145 ;
        RECT 172.115 199.615 172.285 199.785 ;
        RECT 141.365 198.305 141.535 198.475 ;
        RECT 60.875 188.275 61.045 188.445 ;
        RECT 61.875 188.275 62.045 188.445 ;
        RECT 62.875 188.275 63.045 188.445 ;
        RECT 63.875 188.275 64.045 188.445 ;
        RECT 64.875 188.275 65.045 188.445 ;
        RECT 65.875 188.275 66.045 188.445 ;
        RECT 69.305 188.275 69.475 188.445 ;
        RECT 70.305 188.275 70.475 188.445 ;
        RECT 71.305 188.275 71.475 188.445 ;
        RECT 72.305 188.275 72.475 188.445 ;
        RECT 73.305 188.275 73.475 188.445 ;
        RECT 74.305 188.275 74.475 188.445 ;
        RECT 75.305 188.275 75.475 188.445 ;
        RECT 76.305 188.275 76.475 188.445 ;
        RECT 77.305 188.275 77.475 188.445 ;
        RECT 78.305 188.275 78.475 188.445 ;
        RECT 79.305 188.275 79.475 188.445 ;
        RECT 83.025 188.275 83.195 188.445 ;
        RECT 84.025 188.275 84.195 188.445 ;
        RECT 85.025 188.275 85.195 188.445 ;
        RECT 86.025 188.275 86.195 188.445 ;
        RECT 87.025 188.275 87.195 188.445 ;
        RECT 88.025 188.275 88.195 188.445 ;
        RECT 89.025 188.275 89.195 188.445 ;
        RECT 90.025 188.275 90.195 188.445 ;
        RECT 91.025 188.275 91.195 188.445 ;
        RECT 92.025 188.275 92.195 188.445 ;
        RECT 93.025 188.275 93.195 188.445 ;
        RECT 96.755 188.275 96.925 188.445 ;
        RECT 97.755 188.275 97.925 188.445 ;
        RECT 98.755 188.275 98.925 188.445 ;
        RECT 99.755 188.275 99.925 188.445 ;
        RECT 100.755 188.275 100.925 188.445 ;
        RECT 101.755 188.275 101.925 188.445 ;
        RECT 102.755 188.275 102.925 188.445 ;
        RECT 103.755 188.275 103.925 188.445 ;
        RECT 104.755 188.275 104.925 188.445 ;
        RECT 105.755 188.275 105.925 188.445 ;
        RECT 106.755 188.275 106.925 188.445 ;
        RECT 107.755 188.275 107.925 188.445 ;
        RECT 108.755 188.275 108.925 188.445 ;
        RECT 109.755 188.275 109.925 188.445 ;
        RECT 113.405 188.275 113.575 188.445 ;
        RECT 114.405 188.275 114.575 188.445 ;
        RECT 115.405 188.275 115.575 188.445 ;
        RECT 116.405 188.275 116.575 188.445 ;
        RECT 117.405 188.275 117.575 188.445 ;
        RECT 118.405 188.275 118.575 188.445 ;
        RECT 119.405 188.275 119.575 188.445 ;
        RECT 120.405 188.275 120.575 188.445 ;
        RECT 121.405 188.275 121.575 188.445 ;
        RECT 122.405 188.275 122.575 188.445 ;
        RECT 123.405 188.275 123.575 188.445 ;
        RECT 128.005 188.275 128.175 188.445 ;
        RECT 130.005 188.275 130.175 188.445 ;
        RECT 132.005 188.275 132.175 188.445 ;
        RECT 134.005 188.275 134.175 188.445 ;
        RECT 136.005 188.275 136.175 188.445 ;
        RECT 138.005 188.275 138.175 188.445 ;
        RECT 140.005 188.275 140.175 188.445 ;
        RECT 142.005 188.275 142.175 188.445 ;
        RECT 144.005 188.275 144.175 188.445 ;
        RECT 146.005 188.275 146.175 188.445 ;
        RECT 150.555 188.275 150.725 188.445 ;
        RECT 152.555 188.275 152.725 188.445 ;
        RECT 154.555 188.275 154.725 188.445 ;
        RECT 156.555 188.275 156.725 188.445 ;
        RECT 158.555 188.275 158.725 188.445 ;
        RECT 160.555 188.275 160.725 188.445 ;
        RECT 162.555 188.275 162.725 188.445 ;
        RECT 164.555 188.275 164.725 188.445 ;
        RECT 166.555 188.275 166.725 188.445 ;
        RECT 168.555 188.275 168.725 188.445 ;
        RECT 170.555 188.275 170.725 188.445 ;
        RECT 172.555 188.275 172.725 188.445 ;
        RECT 174.555 188.275 174.725 188.445 ;
        RECT 176.555 188.275 176.725 188.445 ;
        RECT 178.555 188.275 178.725 188.445 ;
        RECT 180.555 188.275 180.725 188.445 ;
        RECT 182.555 188.275 182.725 188.445 ;
        RECT 184.555 188.275 184.725 188.445 ;
        RECT 188.275 188.275 188.445 188.445 ;
        RECT 190.275 188.275 190.445 188.445 ;
        RECT 192.275 188.275 192.445 188.445 ;
        RECT 194.275 188.275 194.445 188.445 ;
        RECT 196.275 188.275 196.445 188.445 ;
        RECT 198.275 188.275 198.445 188.445 ;
        RECT 200.275 188.275 200.445 188.445 ;
        RECT 209.835 188.275 210.005 188.445 ;
        RECT 210.835 188.275 211.005 188.445 ;
        RECT 211.835 188.275 212.005 188.445 ;
        RECT 212.835 188.275 213.005 188.445 ;
        RECT 213.835 188.275 214.005 188.445 ;
        RECT 214.835 188.275 215.005 188.445 ;
        RECT 215.835 188.275 216.005 188.445 ;
        RECT 216.835 188.275 217.005 188.445 ;
        RECT 217.835 188.275 218.005 188.445 ;
        RECT 218.835 188.275 219.005 188.445 ;
        RECT 219.835 188.275 220.005 188.445 ;
        RECT 220.835 188.275 221.005 188.445 ;
        RECT 221.835 188.275 222.005 188.445 ;
        RECT 222.835 188.275 223.005 188.445 ;
        RECT 223.835 188.275 224.005 188.445 ;
        RECT 224.835 188.275 225.005 188.445 ;
        RECT 225.835 188.275 226.005 188.445 ;
        RECT 226.835 188.275 227.005 188.445 ;
        RECT 227.835 188.275 228.005 188.445 ;
        RECT 228.835 188.275 229.005 188.445 ;
        RECT 229.835 188.275 230.005 188.445 ;
        RECT 230.835 188.275 231.005 188.445 ;
        RECT 231.835 188.275 232.005 188.445 ;
        RECT 232.835 188.275 233.005 188.445 ;
        RECT 233.835 188.275 234.005 188.445 ;
        RECT 234.835 188.275 235.005 188.445 ;
        RECT 235.835 188.275 236.005 188.445 ;
        RECT 236.835 188.275 237.005 188.445 ;
        RECT 237.835 188.275 238.005 188.445 ;
        RECT 238.835 188.275 239.005 188.445 ;
        RECT 239.835 188.275 240.005 188.445 ;
        RECT 240.835 188.275 241.005 188.445 ;
        RECT 241.835 188.275 242.005 188.445 ;
        RECT 242.835 188.275 243.005 188.445 ;
        RECT 243.835 188.275 244.005 188.445 ;
        RECT 244.835 188.275 245.005 188.445 ;
        RECT 245.835 188.275 246.005 188.445 ;
        RECT 246.835 188.275 247.005 188.445 ;
        RECT 247.835 188.275 248.005 188.445 ;
        RECT 248.835 188.275 249.005 188.445 ;
        RECT 249.835 188.275 250.005 188.445 ;
        RECT 250.835 188.275 251.005 188.445 ;
        RECT 251.835 188.275 252.005 188.445 ;
        RECT 252.835 188.275 253.005 188.445 ;
        RECT 253.835 188.275 254.005 188.445 ;
        RECT 254.835 188.275 255.005 188.445 ;
        RECT 255.835 188.275 256.005 188.445 ;
        RECT 256.835 188.275 257.005 188.445 ;
        RECT 257.835 188.275 258.005 188.445 ;
        RECT 258.835 188.275 259.005 188.445 ;
        RECT 259.835 188.275 260.005 188.445 ;
        RECT 260.835 188.275 261.005 188.445 ;
        RECT 261.835 188.275 262.005 188.445 ;
        RECT 187.825 187.425 187.995 187.595 ;
        RECT 189.885 186.935 190.055 187.105 ;
        RECT 189.885 186.575 190.055 186.745 ;
        RECT 189.885 186.215 190.055 186.385 ;
        RECT 189.885 185.855 190.055 186.025 ;
        RECT 189.885 185.495 190.055 185.665 ;
        RECT 189.885 185.135 190.055 185.305 ;
        RECT 189.885 184.775 190.055 184.945 ;
        RECT 189.885 184.415 190.055 184.585 ;
        RECT 189.885 184.055 190.055 184.225 ;
        RECT 189.885 183.695 190.055 183.865 ;
        RECT 189.885 183.335 190.055 183.505 ;
        RECT 189.885 182.975 190.055 183.145 ;
        RECT 189.885 182.615 190.055 182.785 ;
        RECT 189.885 182.255 190.055 182.425 ;
        RECT 189.885 181.895 190.055 182.065 ;
        RECT 189.885 181.535 190.055 181.705 ;
        RECT 189.885 181.175 190.055 181.345 ;
        RECT 189.885 180.815 190.055 180.985 ;
        RECT 194.465 186.935 194.635 187.105 ;
        RECT 194.465 186.575 194.635 186.745 ;
        RECT 194.465 186.215 194.635 186.385 ;
        RECT 194.465 185.855 194.635 186.025 ;
        RECT 194.465 185.495 194.635 185.665 ;
        RECT 194.465 185.135 194.635 185.305 ;
        RECT 194.465 184.775 194.635 184.945 ;
        RECT 194.465 184.415 194.635 184.585 ;
        RECT 194.465 184.055 194.635 184.225 ;
        RECT 194.465 183.695 194.635 183.865 ;
        RECT 194.465 183.335 194.635 183.505 ;
        RECT 194.465 182.975 194.635 183.145 ;
        RECT 194.465 182.615 194.635 182.785 ;
        RECT 194.465 182.255 194.635 182.425 ;
        RECT 194.465 181.895 194.635 182.065 ;
        RECT 194.465 181.535 194.635 181.705 ;
        RECT 194.465 181.175 194.635 181.345 ;
        RECT 194.465 180.815 194.635 180.985 ;
        RECT 199.045 186.935 199.215 187.105 ;
        RECT 199.045 186.575 199.215 186.745 ;
        RECT 199.045 186.215 199.215 186.385 ;
        RECT 199.045 185.855 199.215 186.025 ;
        RECT 199.045 185.495 199.215 185.665 ;
        RECT 199.045 185.135 199.215 185.305 ;
        RECT 199.045 184.775 199.215 184.945 ;
        RECT 199.045 184.415 199.215 184.585 ;
        RECT 199.045 184.055 199.215 184.225 ;
        RECT 199.045 183.695 199.215 183.865 ;
        RECT 199.045 183.335 199.215 183.505 ;
        RECT 199.045 182.975 199.215 183.145 ;
        RECT 199.045 182.615 199.215 182.785 ;
        RECT 199.045 182.255 199.215 182.425 ;
        RECT 199.045 181.895 199.215 182.065 ;
        RECT 199.045 181.535 199.215 181.705 ;
        RECT 199.045 181.175 199.215 181.345 ;
        RECT 199.045 180.815 199.215 180.985 ;
        RECT 97.235 169.475 97.405 169.645 ;
        RECT 98.235 169.475 98.405 169.645 ;
        RECT 99.235 169.475 99.405 169.645 ;
        RECT 100.235 169.475 100.405 169.645 ;
        RECT 101.235 169.475 101.405 169.645 ;
        RECT 102.235 169.475 102.405 169.645 ;
        RECT 103.235 169.475 103.405 169.645 ;
        RECT 104.235 169.475 104.405 169.645 ;
        RECT 105.235 169.475 105.405 169.645 ;
        RECT 106.235 169.475 106.405 169.645 ;
        RECT 107.235 169.475 107.405 169.645 ;
        RECT 110.965 169.475 111.135 169.645 ;
        RECT 111.965 169.475 112.135 169.645 ;
        RECT 112.965 169.475 113.135 169.645 ;
        RECT 113.965 169.475 114.135 169.645 ;
        RECT 114.965 169.475 115.135 169.645 ;
        RECT 115.965 169.475 116.135 169.645 ;
        RECT 116.965 169.475 117.135 169.645 ;
        RECT 117.965 169.475 118.135 169.645 ;
        RECT 118.965 169.475 119.135 169.645 ;
        RECT 119.965 169.475 120.135 169.645 ;
        RECT 120.965 169.475 121.135 169.645 ;
        RECT 121.965 169.475 122.135 169.645 ;
        RECT 122.965 169.475 123.135 169.645 ;
        RECT 123.965 169.475 124.135 169.645 ;
        RECT 131.935 169.475 132.105 169.645 ;
        RECT 133.935 169.475 134.105 169.645 ;
        RECT 135.935 169.475 136.105 169.645 ;
        RECT 137.935 169.475 138.105 169.645 ;
        RECT 139.935 169.475 140.105 169.645 ;
        RECT 141.935 169.475 142.105 169.645 ;
        RECT 143.935 169.475 144.105 169.645 ;
        RECT 145.935 169.475 146.105 169.645 ;
        RECT 147.935 169.475 148.105 169.645 ;
        RECT 149.935 169.475 150.105 169.645 ;
        RECT 151.935 169.475 152.105 169.645 ;
        RECT 153.935 169.475 154.105 169.645 ;
        RECT 155.935 169.475 156.105 169.645 ;
        RECT 157.935 169.475 158.105 169.645 ;
        RECT 159.935 169.475 160.105 169.645 ;
        RECT 161.935 169.475 162.105 169.645 ;
        RECT 163.935 169.475 164.105 169.645 ;
        RECT 165.935 169.475 166.105 169.645 ;
        RECT 169.175 169.475 169.345 169.645 ;
        RECT 171.175 169.475 171.345 169.645 ;
        RECT 173.175 169.475 173.345 169.645 ;
        RECT 175.175 169.475 175.345 169.645 ;
        RECT 177.175 169.475 177.345 169.645 ;
        RECT 179.175 169.475 179.345 169.645 ;
        RECT 181.175 169.475 181.345 169.645 ;
        RECT 183.175 169.475 183.345 169.645 ;
        RECT 185.175 169.475 185.345 169.645 ;
        RECT 187.175 169.475 187.345 169.645 ;
        RECT 189.175 169.475 189.345 169.645 ;
        RECT 191.175 169.475 191.345 169.645 ;
        RECT 193.175 169.475 193.345 169.645 ;
        RECT 195.175 169.475 195.345 169.645 ;
        RECT 197.175 169.475 197.345 169.645 ;
        RECT 199.175 169.475 199.345 169.645 ;
        RECT 201.175 169.475 201.345 169.645 ;
        RECT 203.175 169.475 203.345 169.645 ;
        RECT 209.835 169.475 210.005 169.645 ;
        RECT 210.835 169.475 211.005 169.645 ;
        RECT 211.835 169.475 212.005 169.645 ;
        RECT 212.835 169.475 213.005 169.645 ;
        RECT 213.835 169.475 214.005 169.645 ;
        RECT 214.835 169.475 215.005 169.645 ;
        RECT 215.835 169.475 216.005 169.645 ;
        RECT 216.835 169.475 217.005 169.645 ;
        RECT 217.835 169.475 218.005 169.645 ;
        RECT 218.835 169.475 219.005 169.645 ;
        RECT 219.835 169.475 220.005 169.645 ;
        RECT 220.835 169.475 221.005 169.645 ;
        RECT 221.835 169.475 222.005 169.645 ;
        RECT 222.835 169.475 223.005 169.645 ;
        RECT 223.835 169.475 224.005 169.645 ;
        RECT 224.835 169.475 225.005 169.645 ;
        RECT 225.835 169.475 226.005 169.645 ;
        RECT 226.835 169.475 227.005 169.645 ;
        RECT 227.835 169.475 228.005 169.645 ;
        RECT 228.835 169.475 229.005 169.645 ;
        RECT 229.835 169.475 230.005 169.645 ;
        RECT 230.835 169.475 231.005 169.645 ;
        RECT 231.835 169.475 232.005 169.645 ;
        RECT 232.835 169.475 233.005 169.645 ;
        RECT 233.835 169.475 234.005 169.645 ;
        RECT 234.835 169.475 235.005 169.645 ;
        RECT 235.835 169.475 236.005 169.645 ;
        RECT 236.835 169.475 237.005 169.645 ;
        RECT 237.835 169.475 238.005 169.645 ;
        RECT 238.835 169.475 239.005 169.645 ;
        RECT 239.835 169.475 240.005 169.645 ;
        RECT 240.835 169.475 241.005 169.645 ;
        RECT 241.835 169.475 242.005 169.645 ;
        RECT 242.835 169.475 243.005 169.645 ;
        RECT 243.835 169.475 244.005 169.645 ;
        RECT 244.835 169.475 245.005 169.645 ;
        RECT 245.835 169.475 246.005 169.645 ;
        RECT 246.835 169.475 247.005 169.645 ;
        RECT 247.835 169.475 248.005 169.645 ;
        RECT 248.835 169.475 249.005 169.645 ;
        RECT 249.835 169.475 250.005 169.645 ;
        RECT 250.835 169.475 251.005 169.645 ;
        RECT 251.835 169.475 252.005 169.645 ;
        RECT 252.835 169.475 253.005 169.645 ;
        RECT 253.835 169.475 254.005 169.645 ;
        RECT 254.835 169.475 255.005 169.645 ;
        RECT 255.835 169.475 256.005 169.645 ;
        RECT 256.835 169.475 257.005 169.645 ;
        RECT 257.835 169.475 258.005 169.645 ;
        RECT 258.835 169.475 259.005 169.645 ;
        RECT 259.835 169.475 260.005 169.645 ;
        RECT 260.835 169.475 261.005 169.645 ;
        RECT 261.835 169.475 262.005 169.645 ;
        RECT 83.515 150.675 83.685 150.845 ;
        RECT 84.515 150.675 84.685 150.845 ;
        RECT 85.515 150.675 85.685 150.845 ;
        RECT 86.515 150.675 86.685 150.845 ;
        RECT 87.515 150.675 87.685 150.845 ;
        RECT 88.515 150.675 88.685 150.845 ;
        RECT 89.515 150.675 89.685 150.845 ;
        RECT 90.515 150.675 90.685 150.845 ;
        RECT 91.515 150.675 91.685 150.845 ;
        RECT 92.515 150.675 92.685 150.845 ;
        RECT 93.515 150.675 93.685 150.845 ;
        RECT 97.235 150.675 97.405 150.845 ;
        RECT 98.235 150.675 98.405 150.845 ;
        RECT 99.235 150.675 99.405 150.845 ;
        RECT 100.235 150.675 100.405 150.845 ;
        RECT 101.235 150.675 101.405 150.845 ;
        RECT 102.235 150.675 102.405 150.845 ;
        RECT 103.235 150.675 103.405 150.845 ;
        RECT 104.235 150.675 104.405 150.845 ;
        RECT 105.235 150.675 105.405 150.845 ;
        RECT 106.235 150.675 106.405 150.845 ;
        RECT 107.235 150.675 107.405 150.845 ;
        RECT 110.955 150.675 111.125 150.845 ;
        RECT 111.955 150.675 112.125 150.845 ;
        RECT 112.955 150.675 113.125 150.845 ;
        RECT 113.955 150.675 114.125 150.845 ;
        RECT 114.955 150.675 115.125 150.845 ;
        RECT 115.955 150.675 116.125 150.845 ;
        RECT 116.955 150.675 117.125 150.845 ;
        RECT 117.955 150.675 118.125 150.845 ;
        RECT 118.955 150.675 119.125 150.845 ;
        RECT 119.955 150.675 120.125 150.845 ;
        RECT 120.955 150.675 121.125 150.845 ;
        RECT 136.925 150.675 137.095 150.845 ;
        RECT 137.925 150.675 138.095 150.845 ;
        RECT 138.925 150.675 139.095 150.845 ;
        RECT 139.925 150.675 140.095 150.845 ;
        RECT 140.925 150.675 141.095 150.845 ;
        RECT 141.925 150.675 142.095 150.845 ;
        RECT 142.925 150.675 143.095 150.845 ;
        RECT 143.925 150.675 144.095 150.845 ;
        RECT 144.925 150.675 145.095 150.845 ;
        RECT 145.925 150.675 146.095 150.845 ;
        RECT 146.925 150.675 147.095 150.845 ;
        RECT 150.555 150.675 150.725 150.845 ;
        RECT 152.555 150.675 152.725 150.845 ;
        RECT 154.555 150.675 154.725 150.845 ;
        RECT 156.555 150.675 156.725 150.845 ;
        RECT 158.555 150.675 158.725 150.845 ;
        RECT 160.555 150.675 160.725 150.845 ;
        RECT 162.555 150.675 162.725 150.845 ;
        RECT 164.555 150.675 164.725 150.845 ;
        RECT 166.555 150.675 166.725 150.845 ;
        RECT 168.555 150.675 168.725 150.845 ;
        RECT 170.555 150.675 170.725 150.845 ;
        RECT 172.555 150.675 172.725 150.845 ;
        RECT 174.555 150.675 174.725 150.845 ;
        RECT 176.555 150.675 176.725 150.845 ;
        RECT 178.555 150.675 178.725 150.845 ;
        RECT 180.555 150.675 180.725 150.845 ;
        RECT 182.555 150.675 182.725 150.845 ;
        RECT 184.555 150.675 184.725 150.845 ;
        RECT 188.275 150.675 188.445 150.845 ;
        RECT 190.275 150.675 190.445 150.845 ;
        RECT 192.275 150.675 192.445 150.845 ;
        RECT 194.275 150.675 194.445 150.845 ;
        RECT 196.275 150.675 196.445 150.845 ;
        RECT 198.275 150.675 198.445 150.845 ;
        RECT 200.275 150.675 200.445 150.845 ;
        RECT 209.835 150.675 210.005 150.845 ;
        RECT 210.835 150.675 211.005 150.845 ;
        RECT 211.835 150.675 212.005 150.845 ;
        RECT 212.835 150.675 213.005 150.845 ;
        RECT 213.835 150.675 214.005 150.845 ;
        RECT 214.835 150.675 215.005 150.845 ;
        RECT 215.835 150.675 216.005 150.845 ;
        RECT 216.835 150.675 217.005 150.845 ;
        RECT 217.835 150.675 218.005 150.845 ;
        RECT 218.835 150.675 219.005 150.845 ;
        RECT 219.835 150.675 220.005 150.845 ;
        RECT 220.835 150.675 221.005 150.845 ;
        RECT 221.835 150.675 222.005 150.845 ;
        RECT 222.835 150.675 223.005 150.845 ;
        RECT 223.835 150.675 224.005 150.845 ;
        RECT 224.835 150.675 225.005 150.845 ;
        RECT 225.835 150.675 226.005 150.845 ;
        RECT 226.835 150.675 227.005 150.845 ;
        RECT 227.835 150.675 228.005 150.845 ;
        RECT 228.835 150.675 229.005 150.845 ;
        RECT 229.835 150.675 230.005 150.845 ;
        RECT 230.835 150.675 231.005 150.845 ;
        RECT 231.835 150.675 232.005 150.845 ;
        RECT 232.835 150.675 233.005 150.845 ;
        RECT 233.835 150.675 234.005 150.845 ;
        RECT 234.835 150.675 235.005 150.845 ;
        RECT 235.835 150.675 236.005 150.845 ;
        RECT 236.835 150.675 237.005 150.845 ;
        RECT 237.835 150.675 238.005 150.845 ;
        RECT 238.835 150.675 239.005 150.845 ;
        RECT 239.835 150.675 240.005 150.845 ;
        RECT 240.835 150.675 241.005 150.845 ;
        RECT 241.835 150.675 242.005 150.845 ;
        RECT 242.835 150.675 243.005 150.845 ;
        RECT 243.835 150.675 244.005 150.845 ;
        RECT 244.835 150.675 245.005 150.845 ;
        RECT 245.835 150.675 246.005 150.845 ;
        RECT 246.835 150.675 247.005 150.845 ;
        RECT 247.835 150.675 248.005 150.845 ;
        RECT 248.835 150.675 249.005 150.845 ;
        RECT 249.835 150.675 250.005 150.845 ;
        RECT 250.835 150.675 251.005 150.845 ;
        RECT 251.835 150.675 252.005 150.845 ;
        RECT 252.835 150.675 253.005 150.845 ;
        RECT 253.835 150.675 254.005 150.845 ;
        RECT 254.835 150.675 255.005 150.845 ;
        RECT 255.835 150.675 256.005 150.845 ;
        RECT 256.835 150.675 257.005 150.845 ;
        RECT 257.835 150.675 258.005 150.845 ;
        RECT 258.835 150.675 259.005 150.845 ;
        RECT 259.835 150.675 260.005 150.845 ;
        RECT 260.835 150.675 261.005 150.845 ;
        RECT 261.835 150.675 262.005 150.845 ;
        RECT 201.625 149.825 201.795 149.995 ;
        RECT 189.885 149.335 190.055 149.505 ;
        RECT 189.885 148.975 190.055 149.145 ;
        RECT 189.885 148.615 190.055 148.785 ;
        RECT 189.885 148.255 190.055 148.425 ;
        RECT 189.885 147.895 190.055 148.065 ;
        RECT 189.885 147.535 190.055 147.705 ;
        RECT 189.885 147.175 190.055 147.345 ;
        RECT 189.885 146.815 190.055 146.985 ;
        RECT 189.885 146.455 190.055 146.625 ;
        RECT 189.885 146.095 190.055 146.265 ;
        RECT 189.885 145.735 190.055 145.905 ;
        RECT 189.885 145.375 190.055 145.545 ;
        RECT 189.885 145.015 190.055 145.185 ;
        RECT 189.885 144.655 190.055 144.825 ;
        RECT 189.885 144.295 190.055 144.465 ;
        RECT 189.885 143.935 190.055 144.105 ;
        RECT 189.885 143.575 190.055 143.745 ;
        RECT 189.885 143.215 190.055 143.385 ;
        RECT 194.465 149.335 194.635 149.505 ;
        RECT 194.465 148.975 194.635 149.145 ;
        RECT 194.465 148.615 194.635 148.785 ;
        RECT 194.465 148.255 194.635 148.425 ;
        RECT 194.465 147.895 194.635 148.065 ;
        RECT 194.465 147.535 194.635 147.705 ;
        RECT 194.465 147.175 194.635 147.345 ;
        RECT 194.465 146.815 194.635 146.985 ;
        RECT 194.465 146.455 194.635 146.625 ;
        RECT 194.465 146.095 194.635 146.265 ;
        RECT 194.465 145.735 194.635 145.905 ;
        RECT 194.465 145.375 194.635 145.545 ;
        RECT 194.465 145.015 194.635 145.185 ;
        RECT 194.465 144.655 194.635 144.825 ;
        RECT 194.465 144.295 194.635 144.465 ;
        RECT 194.465 143.935 194.635 144.105 ;
        RECT 194.465 143.575 194.635 143.745 ;
        RECT 194.465 143.215 194.635 143.385 ;
        RECT 199.045 149.335 199.215 149.505 ;
        RECT 199.045 148.975 199.215 149.145 ;
        RECT 199.045 148.615 199.215 148.785 ;
        RECT 199.045 148.255 199.215 148.425 ;
        RECT 199.045 147.895 199.215 148.065 ;
        RECT 199.045 147.535 199.215 147.705 ;
        RECT 199.045 147.175 199.215 147.345 ;
        RECT 199.045 146.815 199.215 146.985 ;
        RECT 199.045 146.455 199.215 146.625 ;
        RECT 199.045 146.095 199.215 146.265 ;
        RECT 199.045 145.735 199.215 145.905 ;
        RECT 199.045 145.375 199.215 145.545 ;
        RECT 199.045 145.015 199.215 145.185 ;
        RECT 199.045 144.655 199.215 144.825 ;
        RECT 199.045 144.295 199.215 144.465 ;
        RECT 199.045 143.935 199.215 144.105 ;
        RECT 199.045 143.575 199.215 143.745 ;
        RECT 199.045 143.215 199.215 143.385 ;
        RECT 112.915 131.875 113.085 132.045 ;
        RECT 113.915 131.875 114.085 132.045 ;
        RECT 114.915 131.875 115.085 132.045 ;
        RECT 115.915 131.875 116.085 132.045 ;
        RECT 116.915 131.875 117.085 132.045 ;
        RECT 117.915 131.875 118.085 132.045 ;
        RECT 118.915 131.875 119.085 132.045 ;
        RECT 119.915 131.875 120.085 132.045 ;
        RECT 120.915 131.875 121.085 132.045 ;
        RECT 121.915 131.875 122.085 132.045 ;
        RECT 122.915 131.875 123.085 132.045 ;
        RECT 128.005 131.875 128.175 132.045 ;
        RECT 130.005 131.875 130.175 132.045 ;
        RECT 132.005 131.875 132.175 132.045 ;
        RECT 134.005 131.875 134.175 132.045 ;
        RECT 136.005 131.875 136.175 132.045 ;
        RECT 138.005 131.875 138.175 132.045 ;
        RECT 140.005 131.875 140.175 132.045 ;
        RECT 142.005 131.875 142.175 132.045 ;
        RECT 144.005 131.875 144.175 132.045 ;
        RECT 146.005 131.875 146.175 132.045 ;
        RECT 150.555 131.875 150.725 132.045 ;
        RECT 152.555 131.875 152.725 132.045 ;
        RECT 154.555 131.875 154.725 132.045 ;
        RECT 156.555 131.875 156.725 132.045 ;
        RECT 158.555 131.875 158.725 132.045 ;
        RECT 160.555 131.875 160.725 132.045 ;
        RECT 162.555 131.875 162.725 132.045 ;
        RECT 164.555 131.875 164.725 132.045 ;
        RECT 166.555 131.875 166.725 132.045 ;
        RECT 168.555 131.875 168.725 132.045 ;
        RECT 170.555 131.875 170.725 132.045 ;
        RECT 172.555 131.875 172.725 132.045 ;
        RECT 174.555 131.875 174.725 132.045 ;
        RECT 176.555 131.875 176.725 132.045 ;
        RECT 178.555 131.875 178.725 132.045 ;
        RECT 180.555 131.875 180.725 132.045 ;
        RECT 182.555 131.875 182.725 132.045 ;
        RECT 184.555 131.875 184.725 132.045 ;
        RECT 187.885 131.875 188.055 132.045 ;
        RECT 188.885 131.875 189.055 132.045 ;
        RECT 189.885 131.875 190.055 132.045 ;
        RECT 190.885 131.875 191.055 132.045 ;
        RECT 191.885 131.875 192.055 132.045 ;
        RECT 192.885 131.875 193.055 132.045 ;
        RECT 193.885 131.875 194.055 132.045 ;
        RECT 194.885 131.875 195.055 132.045 ;
        RECT 195.885 131.875 196.055 132.045 ;
        RECT 196.885 131.875 197.055 132.045 ;
        RECT 197.885 131.875 198.055 132.045 ;
        RECT 201.605 131.875 201.775 132.045 ;
        RECT 202.605 131.875 202.775 132.045 ;
        RECT 203.605 131.875 203.775 132.045 ;
        RECT 204.605 131.875 204.775 132.045 ;
        RECT 205.605 131.875 205.775 132.045 ;
        RECT 206.605 131.875 206.775 132.045 ;
        RECT 207.605 131.875 207.775 132.045 ;
        RECT 208.605 131.875 208.775 132.045 ;
        RECT 209.605 131.875 209.775 132.045 ;
        RECT 210.605 131.875 210.775 132.045 ;
        RECT 211.605 131.875 211.775 132.045 ;
        RECT 215.325 131.875 215.495 132.045 ;
        RECT 216.325 131.875 216.495 132.045 ;
        RECT 217.325 131.875 217.495 132.045 ;
        RECT 218.325 131.875 218.495 132.045 ;
        RECT 219.325 131.875 219.495 132.045 ;
        RECT 220.325 131.875 220.495 132.045 ;
        RECT 221.325 131.875 221.495 132.045 ;
        RECT 222.325 131.875 222.495 132.045 ;
        RECT 223.325 131.875 223.495 132.045 ;
        RECT 224.325 131.875 224.495 132.045 ;
        RECT 225.325 131.875 225.495 132.045 ;
        RECT 229.045 131.875 229.215 132.045 ;
        RECT 230.045 131.875 230.215 132.045 ;
        RECT 231.045 131.875 231.215 132.045 ;
        RECT 232.045 131.875 232.215 132.045 ;
        RECT 233.045 131.875 233.215 132.045 ;
        RECT 234.045 131.875 234.215 132.045 ;
        RECT 235.045 131.875 235.215 132.045 ;
        RECT 236.045 131.875 236.215 132.045 ;
        RECT 237.045 131.875 237.215 132.045 ;
        RECT 238.045 131.875 238.215 132.045 ;
        RECT 239.045 131.875 239.215 132.045 ;
        RECT 242.765 131.875 242.935 132.045 ;
        RECT 243.765 131.875 243.935 132.045 ;
        RECT 244.765 131.875 244.935 132.045 ;
        RECT 245.765 131.875 245.935 132.045 ;
        RECT 246.765 131.875 246.935 132.045 ;
        RECT 247.765 131.875 247.935 132.045 ;
        RECT 248.765 131.875 248.935 132.045 ;
        RECT 249.765 131.875 249.935 132.045 ;
        RECT 250.765 131.875 250.935 132.045 ;
        RECT 251.765 131.875 251.935 132.045 ;
        RECT 252.765 131.875 252.935 132.045 ;
        RECT 120.265 113.075 120.435 113.245 ;
        RECT 121.265 113.075 121.435 113.245 ;
        RECT 122.265 113.075 122.435 113.245 ;
        RECT 123.265 113.075 123.435 113.245 ;
        RECT 124.265 113.075 124.435 113.245 ;
        RECT 125.265 113.075 125.435 113.245 ;
        RECT 126.265 113.075 126.435 113.245 ;
        RECT 127.265 113.075 127.435 113.245 ;
        RECT 128.265 113.075 128.435 113.245 ;
        RECT 129.265 113.075 129.435 113.245 ;
        RECT 130.265 113.075 130.435 113.245 ;
        RECT 136.925 113.075 137.095 113.245 ;
        RECT 137.925 113.075 138.095 113.245 ;
        RECT 138.925 113.075 139.095 113.245 ;
        RECT 139.925 113.075 140.095 113.245 ;
        RECT 140.925 113.075 141.095 113.245 ;
        RECT 141.925 113.075 142.095 113.245 ;
        RECT 142.925 113.075 143.095 113.245 ;
        RECT 143.925 113.075 144.095 113.245 ;
        RECT 144.925 113.075 145.095 113.245 ;
        RECT 145.925 113.075 146.095 113.245 ;
        RECT 146.925 113.075 147.095 113.245 ;
        RECT 150.645 113.075 150.815 113.245 ;
        RECT 151.645 113.075 151.815 113.245 ;
        RECT 152.645 113.075 152.815 113.245 ;
        RECT 153.645 113.075 153.815 113.245 ;
        RECT 154.645 113.075 154.815 113.245 ;
        RECT 155.645 113.075 155.815 113.245 ;
        RECT 156.645 113.075 156.815 113.245 ;
        RECT 157.645 113.075 157.815 113.245 ;
        RECT 158.645 113.075 158.815 113.245 ;
        RECT 159.645 113.075 159.815 113.245 ;
        RECT 160.645 113.075 160.815 113.245 ;
        RECT 166.815 113.075 166.985 113.245 ;
        RECT 167.815 113.075 167.985 113.245 ;
        RECT 168.815 113.075 168.985 113.245 ;
        RECT 169.815 113.075 169.985 113.245 ;
        RECT 170.815 113.075 170.985 113.245 ;
        RECT 171.815 113.075 171.985 113.245 ;
        RECT 172.815 113.075 172.985 113.245 ;
        RECT 173.815 113.075 173.985 113.245 ;
        RECT 174.815 113.075 174.985 113.245 ;
        RECT 175.815 113.075 175.985 113.245 ;
        RECT 176.815 113.075 176.985 113.245 ;
        RECT 187.885 113.075 188.055 113.245 ;
        RECT 188.885 113.075 189.055 113.245 ;
        RECT 189.885 113.075 190.055 113.245 ;
        RECT 190.885 113.075 191.055 113.245 ;
        RECT 191.885 113.075 192.055 113.245 ;
        RECT 192.885 113.075 193.055 113.245 ;
        RECT 193.885 113.075 194.055 113.245 ;
        RECT 194.885 113.075 195.055 113.245 ;
        RECT 195.885 113.075 196.055 113.245 ;
        RECT 196.885 113.075 197.055 113.245 ;
        RECT 197.885 113.075 198.055 113.245 ;
        RECT 201.605 113.075 201.775 113.245 ;
        RECT 202.605 113.075 202.775 113.245 ;
        RECT 203.605 113.075 203.775 113.245 ;
        RECT 204.605 113.075 204.775 113.245 ;
        RECT 205.605 113.075 205.775 113.245 ;
        RECT 206.605 113.075 206.775 113.245 ;
        RECT 207.605 113.075 207.775 113.245 ;
        RECT 208.605 113.075 208.775 113.245 ;
        RECT 209.605 113.075 209.775 113.245 ;
        RECT 210.605 113.075 210.775 113.245 ;
        RECT 211.605 113.075 211.775 113.245 ;
        RECT 242.765 113.075 242.935 113.245 ;
        RECT 243.765 113.075 243.935 113.245 ;
        RECT 244.765 113.075 244.935 113.245 ;
        RECT 245.765 113.075 245.935 113.245 ;
        RECT 246.765 113.075 246.935 113.245 ;
        RECT 247.765 113.075 247.935 113.245 ;
        RECT 248.765 113.075 248.935 113.245 ;
        RECT 249.765 113.075 249.935 113.245 ;
        RECT 250.765 113.075 250.935 113.245 ;
        RECT 251.765 113.075 251.935 113.245 ;
        RECT 252.765 113.075 252.935 113.245 ;
        RECT 125.065 94.275 125.235 94.445 ;
        RECT 127.065 94.275 127.235 94.445 ;
        RECT 129.065 94.275 129.235 94.445 ;
        RECT 131.065 94.275 131.235 94.445 ;
        RECT 133.065 94.275 133.235 94.445 ;
        RECT 135.065 94.275 135.235 94.445 ;
        RECT 137.065 94.275 137.235 94.445 ;
        RECT 139.065 94.275 139.235 94.445 ;
        RECT 141.065 94.275 141.235 94.445 ;
        RECT 143.065 94.275 143.235 94.445 ;
        RECT 145.065 94.275 145.235 94.445 ;
        RECT 147.065 94.275 147.235 94.445 ;
        RECT 149.065 94.275 149.235 94.445 ;
        RECT 151.065 94.275 151.235 94.445 ;
        RECT 153.065 94.275 153.235 94.445 ;
        RECT 155.065 94.275 155.235 94.445 ;
        RECT 157.065 94.275 157.235 94.445 ;
        RECT 159.065 94.275 159.235 94.445 ;
        RECT 161.065 94.275 161.235 94.445 ;
        RECT 163.065 94.275 163.235 94.445 ;
        RECT 165.065 94.275 165.235 94.445 ;
        RECT 167.065 94.275 167.235 94.445 ;
        RECT 169.065 94.275 169.235 94.445 ;
        RECT 171.065 94.275 171.235 94.445 ;
        RECT 173.065 94.275 173.235 94.445 ;
        RECT 175.065 94.275 175.235 94.445 ;
        RECT 177.065 94.275 177.235 94.445 ;
        RECT 179.065 94.275 179.235 94.445 ;
        RECT 181.065 94.275 181.235 94.445 ;
        RECT 183.065 94.275 183.235 94.445 ;
        RECT 185.065 94.275 185.235 94.445 ;
        RECT 187.065 94.275 187.235 94.445 ;
        RECT 189.065 94.275 189.235 94.445 ;
        RECT 191.065 94.275 191.235 94.445 ;
        RECT 193.065 94.275 193.235 94.445 ;
        RECT 195.065 94.275 195.235 94.445 ;
        RECT 197.065 94.275 197.235 94.445 ;
        RECT 199.065 94.275 199.235 94.445 ;
        RECT 201.065 94.275 201.235 94.445 ;
        RECT 203.065 94.275 203.235 94.445 ;
        RECT 205.065 94.275 205.235 94.445 ;
        RECT 207.065 94.275 207.235 94.445 ;
        RECT 209.065 94.275 209.235 94.445 ;
        RECT 211.065 94.275 211.235 94.445 ;
        RECT 213.065 94.275 213.235 94.445 ;
        RECT 215.065 94.275 215.235 94.445 ;
        RECT 217.065 94.275 217.235 94.445 ;
        RECT 219.065 94.275 219.235 94.445 ;
        RECT 221.065 94.275 221.235 94.445 ;
        RECT 223.065 94.275 223.235 94.445 ;
        RECT 225.065 94.275 225.235 94.445 ;
        RECT 227.065 94.275 227.235 94.445 ;
        RECT 229.065 94.275 229.235 94.445 ;
        RECT 231.065 94.275 231.235 94.445 ;
        RECT 233.065 94.275 233.235 94.445 ;
        RECT 235.065 94.275 235.235 94.445 ;
        RECT 237.065 94.275 237.235 94.445 ;
        RECT 239.065 94.275 239.235 94.445 ;
        RECT 241.065 94.275 241.235 94.445 ;
        RECT 243.065 94.275 243.235 94.445 ;
        RECT 245.065 94.275 245.235 94.445 ;
        RECT 247.065 94.275 247.235 94.445 ;
        RECT 249.065 94.275 249.235 94.445 ;
        RECT 251.065 94.275 251.235 94.445 ;
        RECT 253.065 94.275 253.235 94.445 ;
        RECT 255.065 94.275 255.235 94.445 ;
        RECT 257.065 94.275 257.235 94.445 ;
        RECT 259.065 94.275 259.235 94.445 ;
        RECT 261.065 94.275 261.235 94.445 ;
        RECT 126.675 92.935 126.845 93.105 ;
        RECT 126.675 92.575 126.845 92.745 ;
        RECT 126.675 92.215 126.845 92.385 ;
        RECT 126.675 91.855 126.845 92.025 ;
        RECT 126.675 91.495 126.845 91.665 ;
        RECT 126.675 91.135 126.845 91.305 ;
        RECT 126.675 90.775 126.845 90.945 ;
        RECT 126.675 90.415 126.845 90.585 ;
        RECT 126.675 90.055 126.845 90.225 ;
        RECT 126.675 89.695 126.845 89.865 ;
        RECT 126.675 89.335 126.845 89.505 ;
        RECT 126.675 88.975 126.845 89.145 ;
        RECT 126.675 88.615 126.845 88.785 ;
        RECT 126.675 88.255 126.845 88.425 ;
        RECT 126.675 87.895 126.845 88.065 ;
        RECT 126.675 87.535 126.845 87.705 ;
        RECT 126.675 87.175 126.845 87.345 ;
        RECT 126.675 86.815 126.845 86.985 ;
        RECT 131.255 92.935 131.425 93.105 ;
        RECT 131.255 92.575 131.425 92.745 ;
        RECT 131.255 92.215 131.425 92.385 ;
        RECT 131.255 91.855 131.425 92.025 ;
        RECT 131.255 91.495 131.425 91.665 ;
        RECT 131.255 91.135 131.425 91.305 ;
        RECT 131.255 90.775 131.425 90.945 ;
        RECT 131.255 90.415 131.425 90.585 ;
        RECT 131.255 90.055 131.425 90.225 ;
        RECT 131.255 89.695 131.425 89.865 ;
        RECT 131.255 89.335 131.425 89.505 ;
        RECT 131.255 88.975 131.425 89.145 ;
        RECT 131.255 88.615 131.425 88.785 ;
        RECT 131.255 88.255 131.425 88.425 ;
        RECT 131.255 87.895 131.425 88.065 ;
        RECT 131.255 87.535 131.425 87.705 ;
        RECT 131.255 87.175 131.425 87.345 ;
        RECT 131.255 86.815 131.425 86.985 ;
        RECT 135.835 92.935 136.005 93.105 ;
        RECT 135.835 92.575 136.005 92.745 ;
        RECT 135.835 92.215 136.005 92.385 ;
        RECT 135.835 91.855 136.005 92.025 ;
        RECT 135.835 91.495 136.005 91.665 ;
        RECT 135.835 91.135 136.005 91.305 ;
        RECT 135.835 90.775 136.005 90.945 ;
        RECT 135.835 90.415 136.005 90.585 ;
        RECT 135.835 90.055 136.005 90.225 ;
        RECT 135.835 89.695 136.005 89.865 ;
        RECT 135.835 89.335 136.005 89.505 ;
        RECT 135.835 88.975 136.005 89.145 ;
        RECT 135.835 88.615 136.005 88.785 ;
        RECT 135.835 88.255 136.005 88.425 ;
        RECT 135.835 87.895 136.005 88.065 ;
        RECT 135.835 87.535 136.005 87.705 ;
        RECT 135.835 87.175 136.005 87.345 ;
        RECT 135.835 86.815 136.005 86.985 ;
        RECT 140.415 92.935 140.585 93.105 ;
        RECT 140.415 92.575 140.585 92.745 ;
        RECT 140.415 92.215 140.585 92.385 ;
        RECT 140.415 91.855 140.585 92.025 ;
        RECT 140.415 91.495 140.585 91.665 ;
        RECT 140.415 91.135 140.585 91.305 ;
        RECT 140.415 90.775 140.585 90.945 ;
        RECT 140.415 90.415 140.585 90.585 ;
        RECT 140.415 90.055 140.585 90.225 ;
        RECT 140.415 89.695 140.585 89.865 ;
        RECT 140.415 89.335 140.585 89.505 ;
        RECT 140.415 88.975 140.585 89.145 ;
        RECT 140.415 88.615 140.585 88.785 ;
        RECT 140.415 88.255 140.585 88.425 ;
        RECT 140.415 87.895 140.585 88.065 ;
        RECT 140.415 87.535 140.585 87.705 ;
        RECT 140.415 87.175 140.585 87.345 ;
        RECT 140.415 86.815 140.585 86.985 ;
        RECT 144.995 92.935 145.165 93.105 ;
        RECT 144.995 92.575 145.165 92.745 ;
        RECT 144.995 92.215 145.165 92.385 ;
        RECT 144.995 91.855 145.165 92.025 ;
        RECT 144.995 91.495 145.165 91.665 ;
        RECT 144.995 91.135 145.165 91.305 ;
        RECT 144.995 90.775 145.165 90.945 ;
        RECT 144.995 90.415 145.165 90.585 ;
        RECT 144.995 90.055 145.165 90.225 ;
        RECT 144.995 89.695 145.165 89.865 ;
        RECT 144.995 89.335 145.165 89.505 ;
        RECT 144.995 88.975 145.165 89.145 ;
        RECT 144.995 88.615 145.165 88.785 ;
        RECT 144.995 88.255 145.165 88.425 ;
        RECT 144.995 87.895 145.165 88.065 ;
        RECT 144.995 87.535 145.165 87.705 ;
        RECT 144.995 87.175 145.165 87.345 ;
        RECT 144.995 86.815 145.165 86.985 ;
        RECT 149.575 92.935 149.745 93.105 ;
        RECT 149.575 92.575 149.745 92.745 ;
        RECT 149.575 92.215 149.745 92.385 ;
        RECT 149.575 91.855 149.745 92.025 ;
        RECT 149.575 91.495 149.745 91.665 ;
        RECT 149.575 91.135 149.745 91.305 ;
        RECT 149.575 90.775 149.745 90.945 ;
        RECT 149.575 90.415 149.745 90.585 ;
        RECT 149.575 90.055 149.745 90.225 ;
        RECT 149.575 89.695 149.745 89.865 ;
        RECT 149.575 89.335 149.745 89.505 ;
        RECT 149.575 88.975 149.745 89.145 ;
        RECT 149.575 88.615 149.745 88.785 ;
        RECT 149.575 88.255 149.745 88.425 ;
        RECT 149.575 87.895 149.745 88.065 ;
        RECT 149.575 87.535 149.745 87.705 ;
        RECT 149.575 87.175 149.745 87.345 ;
        RECT 149.575 86.815 149.745 86.985 ;
        RECT 154.155 92.935 154.325 93.105 ;
        RECT 154.155 92.575 154.325 92.745 ;
        RECT 154.155 92.215 154.325 92.385 ;
        RECT 154.155 91.855 154.325 92.025 ;
        RECT 154.155 91.495 154.325 91.665 ;
        RECT 154.155 91.135 154.325 91.305 ;
        RECT 154.155 90.775 154.325 90.945 ;
        RECT 154.155 90.415 154.325 90.585 ;
        RECT 154.155 90.055 154.325 90.225 ;
        RECT 154.155 89.695 154.325 89.865 ;
        RECT 154.155 89.335 154.325 89.505 ;
        RECT 154.155 88.975 154.325 89.145 ;
        RECT 154.155 88.615 154.325 88.785 ;
        RECT 154.155 88.255 154.325 88.425 ;
        RECT 154.155 87.895 154.325 88.065 ;
        RECT 154.155 87.535 154.325 87.705 ;
        RECT 154.155 87.175 154.325 87.345 ;
        RECT 154.155 86.815 154.325 86.985 ;
        RECT 158.735 92.935 158.905 93.105 ;
        RECT 158.735 92.575 158.905 92.745 ;
        RECT 158.735 92.215 158.905 92.385 ;
        RECT 158.735 91.855 158.905 92.025 ;
        RECT 158.735 91.495 158.905 91.665 ;
        RECT 158.735 91.135 158.905 91.305 ;
        RECT 158.735 90.775 158.905 90.945 ;
        RECT 158.735 90.415 158.905 90.585 ;
        RECT 158.735 90.055 158.905 90.225 ;
        RECT 158.735 89.695 158.905 89.865 ;
        RECT 158.735 89.335 158.905 89.505 ;
        RECT 158.735 88.975 158.905 89.145 ;
        RECT 158.735 88.615 158.905 88.785 ;
        RECT 158.735 88.255 158.905 88.425 ;
        RECT 158.735 87.895 158.905 88.065 ;
        RECT 158.735 87.535 158.905 87.705 ;
        RECT 158.735 87.175 158.905 87.345 ;
        RECT 158.735 86.815 158.905 86.985 ;
        RECT 163.315 92.935 163.485 93.105 ;
        RECT 163.315 92.575 163.485 92.745 ;
        RECT 163.315 92.215 163.485 92.385 ;
        RECT 163.315 91.855 163.485 92.025 ;
        RECT 163.315 91.495 163.485 91.665 ;
        RECT 163.315 91.135 163.485 91.305 ;
        RECT 163.315 90.775 163.485 90.945 ;
        RECT 163.315 90.415 163.485 90.585 ;
        RECT 163.315 90.055 163.485 90.225 ;
        RECT 163.315 89.695 163.485 89.865 ;
        RECT 163.315 89.335 163.485 89.505 ;
        RECT 163.315 88.975 163.485 89.145 ;
        RECT 163.315 88.615 163.485 88.785 ;
        RECT 163.315 88.255 163.485 88.425 ;
        RECT 163.315 87.895 163.485 88.065 ;
        RECT 163.315 87.535 163.485 87.705 ;
        RECT 163.315 87.175 163.485 87.345 ;
        RECT 163.315 86.815 163.485 86.985 ;
        RECT 167.895 92.935 168.065 93.105 ;
        RECT 167.895 92.575 168.065 92.745 ;
        RECT 167.895 92.215 168.065 92.385 ;
        RECT 167.895 91.855 168.065 92.025 ;
        RECT 167.895 91.495 168.065 91.665 ;
        RECT 167.895 91.135 168.065 91.305 ;
        RECT 167.895 90.775 168.065 90.945 ;
        RECT 167.895 90.415 168.065 90.585 ;
        RECT 167.895 90.055 168.065 90.225 ;
        RECT 167.895 89.695 168.065 89.865 ;
        RECT 167.895 89.335 168.065 89.505 ;
        RECT 167.895 88.975 168.065 89.145 ;
        RECT 167.895 88.615 168.065 88.785 ;
        RECT 167.895 88.255 168.065 88.425 ;
        RECT 167.895 87.895 168.065 88.065 ;
        RECT 167.895 87.535 168.065 87.705 ;
        RECT 167.895 87.175 168.065 87.345 ;
        RECT 167.895 86.815 168.065 86.985 ;
        RECT 172.475 92.935 172.645 93.105 ;
        RECT 172.475 92.575 172.645 92.745 ;
        RECT 172.475 92.215 172.645 92.385 ;
        RECT 172.475 91.855 172.645 92.025 ;
        RECT 172.475 91.495 172.645 91.665 ;
        RECT 172.475 91.135 172.645 91.305 ;
        RECT 172.475 90.775 172.645 90.945 ;
        RECT 172.475 90.415 172.645 90.585 ;
        RECT 172.475 90.055 172.645 90.225 ;
        RECT 172.475 89.695 172.645 89.865 ;
        RECT 172.475 89.335 172.645 89.505 ;
        RECT 172.475 88.975 172.645 89.145 ;
        RECT 172.475 88.615 172.645 88.785 ;
        RECT 172.475 88.255 172.645 88.425 ;
        RECT 172.475 87.895 172.645 88.065 ;
        RECT 172.475 87.535 172.645 87.705 ;
        RECT 172.475 87.175 172.645 87.345 ;
        RECT 172.475 86.815 172.645 86.985 ;
        RECT 177.055 92.935 177.225 93.105 ;
        RECT 177.055 92.575 177.225 92.745 ;
        RECT 177.055 92.215 177.225 92.385 ;
        RECT 177.055 91.855 177.225 92.025 ;
        RECT 177.055 91.495 177.225 91.665 ;
        RECT 177.055 91.135 177.225 91.305 ;
        RECT 177.055 90.775 177.225 90.945 ;
        RECT 177.055 90.415 177.225 90.585 ;
        RECT 177.055 90.055 177.225 90.225 ;
        RECT 177.055 89.695 177.225 89.865 ;
        RECT 177.055 89.335 177.225 89.505 ;
        RECT 177.055 88.975 177.225 89.145 ;
        RECT 177.055 88.615 177.225 88.785 ;
        RECT 177.055 88.255 177.225 88.425 ;
        RECT 177.055 87.895 177.225 88.065 ;
        RECT 177.055 87.535 177.225 87.705 ;
        RECT 177.055 87.175 177.225 87.345 ;
        RECT 177.055 86.815 177.225 86.985 ;
        RECT 181.635 92.935 181.805 93.105 ;
        RECT 181.635 92.575 181.805 92.745 ;
        RECT 181.635 92.215 181.805 92.385 ;
        RECT 181.635 91.855 181.805 92.025 ;
        RECT 181.635 91.495 181.805 91.665 ;
        RECT 181.635 91.135 181.805 91.305 ;
        RECT 181.635 90.775 181.805 90.945 ;
        RECT 181.635 90.415 181.805 90.585 ;
        RECT 181.635 90.055 181.805 90.225 ;
        RECT 181.635 89.695 181.805 89.865 ;
        RECT 181.635 89.335 181.805 89.505 ;
        RECT 181.635 88.975 181.805 89.145 ;
        RECT 181.635 88.615 181.805 88.785 ;
        RECT 181.635 88.255 181.805 88.425 ;
        RECT 181.635 87.895 181.805 88.065 ;
        RECT 181.635 87.535 181.805 87.705 ;
        RECT 181.635 87.175 181.805 87.345 ;
        RECT 181.635 86.815 181.805 86.985 ;
        RECT 186.215 92.935 186.385 93.105 ;
        RECT 186.215 92.575 186.385 92.745 ;
        RECT 186.215 92.215 186.385 92.385 ;
        RECT 186.215 91.855 186.385 92.025 ;
        RECT 186.215 91.495 186.385 91.665 ;
        RECT 186.215 91.135 186.385 91.305 ;
        RECT 186.215 90.775 186.385 90.945 ;
        RECT 186.215 90.415 186.385 90.585 ;
        RECT 186.215 90.055 186.385 90.225 ;
        RECT 186.215 89.695 186.385 89.865 ;
        RECT 186.215 89.335 186.385 89.505 ;
        RECT 186.215 88.975 186.385 89.145 ;
        RECT 186.215 88.615 186.385 88.785 ;
        RECT 186.215 88.255 186.385 88.425 ;
        RECT 186.215 87.895 186.385 88.065 ;
        RECT 186.215 87.535 186.385 87.705 ;
        RECT 186.215 87.175 186.385 87.345 ;
        RECT 186.215 86.815 186.385 86.985 ;
        RECT 190.795 92.935 190.965 93.105 ;
        RECT 190.795 92.575 190.965 92.745 ;
        RECT 190.795 92.215 190.965 92.385 ;
        RECT 190.795 91.855 190.965 92.025 ;
        RECT 190.795 91.495 190.965 91.665 ;
        RECT 190.795 91.135 190.965 91.305 ;
        RECT 190.795 90.775 190.965 90.945 ;
        RECT 190.795 90.415 190.965 90.585 ;
        RECT 190.795 90.055 190.965 90.225 ;
        RECT 190.795 89.695 190.965 89.865 ;
        RECT 190.795 89.335 190.965 89.505 ;
        RECT 190.795 88.975 190.965 89.145 ;
        RECT 190.795 88.615 190.965 88.785 ;
        RECT 190.795 88.255 190.965 88.425 ;
        RECT 190.795 87.895 190.965 88.065 ;
        RECT 190.795 87.535 190.965 87.705 ;
        RECT 190.795 87.175 190.965 87.345 ;
        RECT 190.795 86.815 190.965 86.985 ;
        RECT 195.375 92.935 195.545 93.105 ;
        RECT 195.375 92.575 195.545 92.745 ;
        RECT 195.375 92.215 195.545 92.385 ;
        RECT 195.375 91.855 195.545 92.025 ;
        RECT 195.375 91.495 195.545 91.665 ;
        RECT 195.375 91.135 195.545 91.305 ;
        RECT 195.375 90.775 195.545 90.945 ;
        RECT 195.375 90.415 195.545 90.585 ;
        RECT 195.375 90.055 195.545 90.225 ;
        RECT 195.375 89.695 195.545 89.865 ;
        RECT 195.375 89.335 195.545 89.505 ;
        RECT 195.375 88.975 195.545 89.145 ;
        RECT 195.375 88.615 195.545 88.785 ;
        RECT 195.375 88.255 195.545 88.425 ;
        RECT 195.375 87.895 195.545 88.065 ;
        RECT 195.375 87.535 195.545 87.705 ;
        RECT 195.375 87.175 195.545 87.345 ;
        RECT 195.375 86.815 195.545 86.985 ;
        RECT 199.955 92.935 200.125 93.105 ;
        RECT 199.955 92.575 200.125 92.745 ;
        RECT 199.955 92.215 200.125 92.385 ;
        RECT 199.955 91.855 200.125 92.025 ;
        RECT 199.955 91.495 200.125 91.665 ;
        RECT 199.955 91.135 200.125 91.305 ;
        RECT 199.955 90.775 200.125 90.945 ;
        RECT 199.955 90.415 200.125 90.585 ;
        RECT 199.955 90.055 200.125 90.225 ;
        RECT 199.955 89.695 200.125 89.865 ;
        RECT 199.955 89.335 200.125 89.505 ;
        RECT 199.955 88.975 200.125 89.145 ;
        RECT 199.955 88.615 200.125 88.785 ;
        RECT 199.955 88.255 200.125 88.425 ;
        RECT 199.955 87.895 200.125 88.065 ;
        RECT 199.955 87.535 200.125 87.705 ;
        RECT 199.955 87.175 200.125 87.345 ;
        RECT 199.955 86.815 200.125 86.985 ;
        RECT 204.535 92.935 204.705 93.105 ;
        RECT 204.535 92.575 204.705 92.745 ;
        RECT 204.535 92.215 204.705 92.385 ;
        RECT 204.535 91.855 204.705 92.025 ;
        RECT 204.535 91.495 204.705 91.665 ;
        RECT 204.535 91.135 204.705 91.305 ;
        RECT 204.535 90.775 204.705 90.945 ;
        RECT 204.535 90.415 204.705 90.585 ;
        RECT 204.535 90.055 204.705 90.225 ;
        RECT 204.535 89.695 204.705 89.865 ;
        RECT 204.535 89.335 204.705 89.505 ;
        RECT 204.535 88.975 204.705 89.145 ;
        RECT 204.535 88.615 204.705 88.785 ;
        RECT 204.535 88.255 204.705 88.425 ;
        RECT 204.535 87.895 204.705 88.065 ;
        RECT 204.535 87.535 204.705 87.705 ;
        RECT 204.535 87.175 204.705 87.345 ;
        RECT 204.535 86.815 204.705 86.985 ;
        RECT 209.115 92.935 209.285 93.105 ;
        RECT 209.115 92.575 209.285 92.745 ;
        RECT 209.115 92.215 209.285 92.385 ;
        RECT 209.115 91.855 209.285 92.025 ;
        RECT 209.115 91.495 209.285 91.665 ;
        RECT 209.115 91.135 209.285 91.305 ;
        RECT 209.115 90.775 209.285 90.945 ;
        RECT 209.115 90.415 209.285 90.585 ;
        RECT 209.115 90.055 209.285 90.225 ;
        RECT 209.115 89.695 209.285 89.865 ;
        RECT 209.115 89.335 209.285 89.505 ;
        RECT 209.115 88.975 209.285 89.145 ;
        RECT 209.115 88.615 209.285 88.785 ;
        RECT 209.115 88.255 209.285 88.425 ;
        RECT 209.115 87.895 209.285 88.065 ;
        RECT 209.115 87.535 209.285 87.705 ;
        RECT 209.115 87.175 209.285 87.345 ;
        RECT 209.115 86.815 209.285 86.985 ;
        RECT 213.695 92.935 213.865 93.105 ;
        RECT 213.695 92.575 213.865 92.745 ;
        RECT 213.695 92.215 213.865 92.385 ;
        RECT 213.695 91.855 213.865 92.025 ;
        RECT 213.695 91.495 213.865 91.665 ;
        RECT 213.695 91.135 213.865 91.305 ;
        RECT 213.695 90.775 213.865 90.945 ;
        RECT 213.695 90.415 213.865 90.585 ;
        RECT 213.695 90.055 213.865 90.225 ;
        RECT 213.695 89.695 213.865 89.865 ;
        RECT 213.695 89.335 213.865 89.505 ;
        RECT 213.695 88.975 213.865 89.145 ;
        RECT 213.695 88.615 213.865 88.785 ;
        RECT 213.695 88.255 213.865 88.425 ;
        RECT 213.695 87.895 213.865 88.065 ;
        RECT 213.695 87.535 213.865 87.705 ;
        RECT 213.695 87.175 213.865 87.345 ;
        RECT 213.695 86.815 213.865 86.985 ;
        RECT 218.275 92.935 218.445 93.105 ;
        RECT 218.275 92.575 218.445 92.745 ;
        RECT 218.275 92.215 218.445 92.385 ;
        RECT 218.275 91.855 218.445 92.025 ;
        RECT 218.275 91.495 218.445 91.665 ;
        RECT 218.275 91.135 218.445 91.305 ;
        RECT 218.275 90.775 218.445 90.945 ;
        RECT 218.275 90.415 218.445 90.585 ;
        RECT 218.275 90.055 218.445 90.225 ;
        RECT 218.275 89.695 218.445 89.865 ;
        RECT 218.275 89.335 218.445 89.505 ;
        RECT 218.275 88.975 218.445 89.145 ;
        RECT 218.275 88.615 218.445 88.785 ;
        RECT 218.275 88.255 218.445 88.425 ;
        RECT 218.275 87.895 218.445 88.065 ;
        RECT 218.275 87.535 218.445 87.705 ;
        RECT 218.275 87.175 218.445 87.345 ;
        RECT 218.275 86.815 218.445 86.985 ;
        RECT 222.855 92.935 223.025 93.105 ;
        RECT 222.855 92.575 223.025 92.745 ;
        RECT 222.855 92.215 223.025 92.385 ;
        RECT 222.855 91.855 223.025 92.025 ;
        RECT 222.855 91.495 223.025 91.665 ;
        RECT 222.855 91.135 223.025 91.305 ;
        RECT 222.855 90.775 223.025 90.945 ;
        RECT 222.855 90.415 223.025 90.585 ;
        RECT 222.855 90.055 223.025 90.225 ;
        RECT 222.855 89.695 223.025 89.865 ;
        RECT 222.855 89.335 223.025 89.505 ;
        RECT 222.855 88.975 223.025 89.145 ;
        RECT 222.855 88.615 223.025 88.785 ;
        RECT 222.855 88.255 223.025 88.425 ;
        RECT 222.855 87.895 223.025 88.065 ;
        RECT 222.855 87.535 223.025 87.705 ;
        RECT 222.855 87.175 223.025 87.345 ;
        RECT 222.855 86.815 223.025 86.985 ;
        RECT 227.435 92.935 227.605 93.105 ;
        RECT 227.435 92.575 227.605 92.745 ;
        RECT 227.435 92.215 227.605 92.385 ;
        RECT 227.435 91.855 227.605 92.025 ;
        RECT 227.435 91.495 227.605 91.665 ;
        RECT 227.435 91.135 227.605 91.305 ;
        RECT 227.435 90.775 227.605 90.945 ;
        RECT 227.435 90.415 227.605 90.585 ;
        RECT 227.435 90.055 227.605 90.225 ;
        RECT 227.435 89.695 227.605 89.865 ;
        RECT 227.435 89.335 227.605 89.505 ;
        RECT 227.435 88.975 227.605 89.145 ;
        RECT 227.435 88.615 227.605 88.785 ;
        RECT 227.435 88.255 227.605 88.425 ;
        RECT 227.435 87.895 227.605 88.065 ;
        RECT 227.435 87.535 227.605 87.705 ;
        RECT 227.435 87.175 227.605 87.345 ;
        RECT 227.435 86.815 227.605 86.985 ;
        RECT 232.015 92.935 232.185 93.105 ;
        RECT 232.015 92.575 232.185 92.745 ;
        RECT 232.015 92.215 232.185 92.385 ;
        RECT 232.015 91.855 232.185 92.025 ;
        RECT 232.015 91.495 232.185 91.665 ;
        RECT 232.015 91.135 232.185 91.305 ;
        RECT 232.015 90.775 232.185 90.945 ;
        RECT 232.015 90.415 232.185 90.585 ;
        RECT 232.015 90.055 232.185 90.225 ;
        RECT 232.015 89.695 232.185 89.865 ;
        RECT 232.015 89.335 232.185 89.505 ;
        RECT 232.015 88.975 232.185 89.145 ;
        RECT 232.015 88.615 232.185 88.785 ;
        RECT 232.015 88.255 232.185 88.425 ;
        RECT 232.015 87.895 232.185 88.065 ;
        RECT 232.015 87.535 232.185 87.705 ;
        RECT 232.015 87.175 232.185 87.345 ;
        RECT 232.015 86.815 232.185 86.985 ;
        RECT 236.595 92.935 236.765 93.105 ;
        RECT 236.595 92.575 236.765 92.745 ;
        RECT 236.595 92.215 236.765 92.385 ;
        RECT 236.595 91.855 236.765 92.025 ;
        RECT 236.595 91.495 236.765 91.665 ;
        RECT 236.595 91.135 236.765 91.305 ;
        RECT 236.595 90.775 236.765 90.945 ;
        RECT 236.595 90.415 236.765 90.585 ;
        RECT 236.595 90.055 236.765 90.225 ;
        RECT 236.595 89.695 236.765 89.865 ;
        RECT 236.595 89.335 236.765 89.505 ;
        RECT 236.595 88.975 236.765 89.145 ;
        RECT 236.595 88.615 236.765 88.785 ;
        RECT 236.595 88.255 236.765 88.425 ;
        RECT 236.595 87.895 236.765 88.065 ;
        RECT 236.595 87.535 236.765 87.705 ;
        RECT 236.595 87.175 236.765 87.345 ;
        RECT 236.595 86.815 236.765 86.985 ;
        RECT 241.175 92.935 241.345 93.105 ;
        RECT 241.175 92.575 241.345 92.745 ;
        RECT 241.175 92.215 241.345 92.385 ;
        RECT 241.175 91.855 241.345 92.025 ;
        RECT 241.175 91.495 241.345 91.665 ;
        RECT 241.175 91.135 241.345 91.305 ;
        RECT 241.175 90.775 241.345 90.945 ;
        RECT 241.175 90.415 241.345 90.585 ;
        RECT 241.175 90.055 241.345 90.225 ;
        RECT 241.175 89.695 241.345 89.865 ;
        RECT 241.175 89.335 241.345 89.505 ;
        RECT 241.175 88.975 241.345 89.145 ;
        RECT 241.175 88.615 241.345 88.785 ;
        RECT 241.175 88.255 241.345 88.425 ;
        RECT 241.175 87.895 241.345 88.065 ;
        RECT 241.175 87.535 241.345 87.705 ;
        RECT 241.175 87.175 241.345 87.345 ;
        RECT 241.175 86.815 241.345 86.985 ;
        RECT 245.755 92.935 245.925 93.105 ;
        RECT 245.755 92.575 245.925 92.745 ;
        RECT 245.755 92.215 245.925 92.385 ;
        RECT 245.755 91.855 245.925 92.025 ;
        RECT 245.755 91.495 245.925 91.665 ;
        RECT 245.755 91.135 245.925 91.305 ;
        RECT 245.755 90.775 245.925 90.945 ;
        RECT 245.755 90.415 245.925 90.585 ;
        RECT 245.755 90.055 245.925 90.225 ;
        RECT 245.755 89.695 245.925 89.865 ;
        RECT 245.755 89.335 245.925 89.505 ;
        RECT 245.755 88.975 245.925 89.145 ;
        RECT 245.755 88.615 245.925 88.785 ;
        RECT 245.755 88.255 245.925 88.425 ;
        RECT 245.755 87.895 245.925 88.065 ;
        RECT 245.755 87.535 245.925 87.705 ;
        RECT 245.755 87.175 245.925 87.345 ;
        RECT 245.755 86.815 245.925 86.985 ;
        RECT 250.335 92.935 250.505 93.105 ;
        RECT 250.335 92.575 250.505 92.745 ;
        RECT 250.335 92.215 250.505 92.385 ;
        RECT 250.335 91.855 250.505 92.025 ;
        RECT 250.335 91.495 250.505 91.665 ;
        RECT 250.335 91.135 250.505 91.305 ;
        RECT 250.335 90.775 250.505 90.945 ;
        RECT 250.335 90.415 250.505 90.585 ;
        RECT 250.335 90.055 250.505 90.225 ;
        RECT 250.335 89.695 250.505 89.865 ;
        RECT 250.335 89.335 250.505 89.505 ;
        RECT 250.335 88.975 250.505 89.145 ;
        RECT 250.335 88.615 250.505 88.785 ;
        RECT 250.335 88.255 250.505 88.425 ;
        RECT 250.335 87.895 250.505 88.065 ;
        RECT 250.335 87.535 250.505 87.705 ;
        RECT 250.335 87.175 250.505 87.345 ;
        RECT 250.335 86.815 250.505 86.985 ;
        RECT 254.915 92.935 255.085 93.105 ;
        RECT 254.915 92.575 255.085 92.745 ;
        RECT 254.915 92.215 255.085 92.385 ;
        RECT 254.915 91.855 255.085 92.025 ;
        RECT 254.915 91.495 255.085 91.665 ;
        RECT 254.915 91.135 255.085 91.305 ;
        RECT 254.915 90.775 255.085 90.945 ;
        RECT 254.915 90.415 255.085 90.585 ;
        RECT 254.915 90.055 255.085 90.225 ;
        RECT 254.915 89.695 255.085 89.865 ;
        RECT 254.915 89.335 255.085 89.505 ;
        RECT 254.915 88.975 255.085 89.145 ;
        RECT 254.915 88.615 255.085 88.785 ;
        RECT 254.915 88.255 255.085 88.425 ;
        RECT 254.915 87.895 255.085 88.065 ;
        RECT 254.915 87.535 255.085 87.705 ;
        RECT 254.915 87.175 255.085 87.345 ;
        RECT 254.915 86.815 255.085 86.985 ;
        RECT 259.495 92.935 259.665 93.105 ;
        RECT 259.495 92.575 259.665 92.745 ;
        RECT 259.495 92.215 259.665 92.385 ;
        RECT 259.495 91.855 259.665 92.025 ;
        RECT 259.495 91.495 259.665 91.665 ;
        RECT 259.495 91.135 259.665 91.305 ;
        RECT 259.495 90.775 259.665 90.945 ;
        RECT 259.495 90.415 259.665 90.585 ;
        RECT 259.495 90.055 259.665 90.225 ;
        RECT 259.495 89.695 259.665 89.865 ;
        RECT 259.495 89.335 259.665 89.505 ;
        RECT 259.495 88.975 259.665 89.145 ;
        RECT 259.495 88.615 259.665 88.785 ;
        RECT 259.495 88.255 259.665 88.425 ;
        RECT 259.495 87.895 259.665 88.065 ;
        RECT 259.495 87.535 259.665 87.705 ;
        RECT 259.495 87.175 259.665 87.345 ;
        RECT 259.495 86.815 259.665 86.985 ;
        RECT 220.225 75.475 220.395 75.645 ;
        RECT 221.225 75.475 221.395 75.645 ;
        RECT 222.225 75.475 222.395 75.645 ;
        RECT 223.225 75.475 223.395 75.645 ;
        RECT 224.225 75.475 224.395 75.645 ;
        RECT 225.225 75.475 225.395 75.645 ;
        RECT 226.225 75.475 226.395 75.645 ;
        RECT 227.225 75.475 227.395 75.645 ;
        RECT 228.225 75.475 228.395 75.645 ;
        RECT 229.225 75.475 229.395 75.645 ;
        RECT 230.225 75.475 230.395 75.645 ;
        RECT 233.945 75.475 234.115 75.645 ;
        RECT 234.945 75.475 235.115 75.645 ;
        RECT 235.945 75.475 236.115 75.645 ;
        RECT 236.945 75.475 237.115 75.645 ;
        RECT 237.945 75.475 238.115 75.645 ;
        RECT 238.945 75.475 239.115 75.645 ;
        RECT 239.945 75.475 240.115 75.645 ;
        RECT 240.945 75.475 241.115 75.645 ;
        RECT 241.945 75.475 242.115 75.645 ;
        RECT 242.945 75.475 243.115 75.645 ;
        RECT 243.945 75.475 244.115 75.645 ;
        RECT 247.665 75.475 247.835 75.645 ;
        RECT 248.665 75.475 248.835 75.645 ;
        RECT 249.665 75.475 249.835 75.645 ;
        RECT 250.665 75.475 250.835 75.645 ;
        RECT 251.665 75.475 251.835 75.645 ;
        RECT 252.665 75.475 252.835 75.645 ;
        RECT 253.665 75.475 253.835 75.645 ;
        RECT 254.665 75.475 254.835 75.645 ;
        RECT 255.665 75.475 255.835 75.645 ;
        RECT 256.665 75.475 256.835 75.645 ;
        RECT 257.665 75.475 257.835 75.645 ;
        RECT 219.735 56.675 219.905 56.845 ;
        RECT 220.735 56.675 220.905 56.845 ;
        RECT 221.735 56.675 221.905 56.845 ;
        RECT 222.735 56.675 222.905 56.845 ;
        RECT 223.735 56.675 223.905 56.845 ;
        RECT 224.735 56.675 224.905 56.845 ;
        RECT 225.735 56.675 225.905 56.845 ;
        RECT 226.735 56.675 226.905 56.845 ;
        RECT 227.735 56.675 227.905 56.845 ;
        RECT 228.735 56.675 228.905 56.845 ;
        RECT 229.735 56.675 229.905 56.845 ;
        RECT 233.455 56.675 233.625 56.845 ;
        RECT 234.455 56.675 234.625 56.845 ;
        RECT 235.455 56.675 235.625 56.845 ;
        RECT 236.455 56.675 236.625 56.845 ;
        RECT 237.455 56.675 237.625 56.845 ;
        RECT 238.455 56.675 238.625 56.845 ;
        RECT 239.455 56.675 239.625 56.845 ;
        RECT 240.455 56.675 240.625 56.845 ;
        RECT 241.455 56.675 241.625 56.845 ;
        RECT 242.455 56.675 242.625 56.845 ;
        RECT 243.455 56.675 243.625 56.845 ;
        RECT 247.175 56.675 247.345 56.845 ;
        RECT 248.175 56.675 248.345 56.845 ;
        RECT 249.175 56.675 249.345 56.845 ;
        RECT 250.175 56.675 250.345 56.845 ;
        RECT 251.175 56.675 251.345 56.845 ;
        RECT 252.175 56.675 252.345 56.845 ;
        RECT 253.175 56.675 253.345 56.845 ;
        RECT 254.175 56.675 254.345 56.845 ;
        RECT 255.175 56.675 255.345 56.845 ;
        RECT 256.175 56.675 256.345 56.845 ;
        RECT 257.175 56.675 257.345 56.845 ;
        RECT 223.655 37.875 223.825 38.045 ;
        RECT 224.655 37.875 224.825 38.045 ;
        RECT 225.655 37.875 225.825 38.045 ;
        RECT 226.655 37.875 226.825 38.045 ;
        RECT 227.655 37.875 227.825 38.045 ;
        RECT 228.655 37.875 228.825 38.045 ;
        RECT 229.655 37.875 229.825 38.045 ;
        RECT 230.655 37.875 230.825 38.045 ;
        RECT 231.655 37.875 231.825 38.045 ;
        RECT 232.655 37.875 232.825 38.045 ;
        RECT 233.655 37.875 233.825 38.045 ;
        RECT 237.375 37.875 237.545 38.045 ;
        RECT 238.375 37.875 238.545 38.045 ;
        RECT 239.375 37.875 239.545 38.045 ;
        RECT 240.375 37.875 240.545 38.045 ;
        RECT 241.375 37.875 241.545 38.045 ;
        RECT 242.375 37.875 242.545 38.045 ;
        RECT 243.375 37.875 243.545 38.045 ;
        RECT 244.375 37.875 244.545 38.045 ;
        RECT 245.375 37.875 245.545 38.045 ;
        RECT 246.375 37.875 246.545 38.045 ;
        RECT 247.375 37.875 247.545 38.045 ;
        RECT 251.095 37.875 251.265 38.045 ;
        RECT 252.095 37.875 252.265 38.045 ;
        RECT 253.095 37.875 253.265 38.045 ;
        RECT 254.095 37.875 254.265 38.045 ;
        RECT 255.095 37.875 255.265 38.045 ;
        RECT 256.095 37.875 256.265 38.045 ;
        RECT 257.095 37.875 257.265 38.045 ;
        RECT 258.095 37.875 258.265 38.045 ;
        RECT 259.095 37.875 259.265 38.045 ;
        RECT 260.095 37.875 260.265 38.045 ;
        RECT 261.095 37.875 261.265 38.045 ;
      LAYER met1 ;
        RECT 16.740 244.460 275.440 245.060 ;
        RECT 126.660 243.585 126.800 244.460 ;
        RECT 126.645 237.135 126.875 243.585 ;
        RECT 131.225 237.135 131.455 243.585 ;
        RECT 135.805 237.135 136.035 243.585 ;
        RECT 140.385 237.135 140.615 243.585 ;
        RECT 144.965 237.135 145.195 243.585 ;
        RECT 149.545 237.135 149.775 243.585 ;
        RECT 154.125 237.135 154.355 243.585 ;
        RECT 158.705 237.135 158.935 243.585 ;
        RECT 163.285 237.135 163.515 243.585 ;
        RECT 167.865 237.135 168.095 243.585 ;
        RECT 172.445 237.135 172.675 243.585 ;
        RECT 177.025 237.135 177.255 243.585 ;
        RECT 181.605 237.135 181.835 243.585 ;
        RECT 186.185 237.135 186.415 243.585 ;
        RECT 190.765 237.135 190.995 243.585 ;
        RECT 195.345 237.135 195.575 243.585 ;
        RECT 199.925 237.135 200.155 243.585 ;
        RECT 204.505 237.135 204.735 243.585 ;
        RECT 209.085 237.135 209.315 243.585 ;
        RECT 213.665 237.135 213.895 243.585 ;
        RECT 218.245 237.135 218.475 243.585 ;
        RECT 222.825 237.135 223.055 243.585 ;
        RECT 227.405 237.135 227.635 243.585 ;
        RECT 231.985 237.135 232.215 243.585 ;
        RECT 236.565 237.135 236.795 243.585 ;
        RECT 241.145 237.135 241.375 243.585 ;
        RECT 245.725 237.135 245.955 243.585 ;
        RECT 250.305 237.135 250.535 243.585 ;
        RECT 254.885 237.135 255.115 243.585 ;
        RECT 259.465 237.135 259.695 243.585 ;
        RECT 16.740 225.660 275.440 226.260 ;
        RECT 128.040 224.785 128.180 225.660 ;
        RECT 77.645 218.335 77.875 224.785 ;
        RECT 82.225 218.335 82.455 224.785 ;
        RECT 86.805 218.335 87.035 224.785 ;
        RECT 91.385 218.335 91.615 224.785 ;
        RECT 95.965 218.335 96.195 224.785 ;
        RECT 100.545 218.335 100.775 224.785 ;
        RECT 105.125 218.335 105.355 224.785 ;
        RECT 109.705 218.335 109.935 224.785 ;
        RECT 114.285 218.335 114.515 224.785 ;
        RECT 118.865 218.335 119.095 224.785 ;
        RECT 123.445 218.335 123.675 224.785 ;
        RECT 128.025 218.335 128.255 224.785 ;
        RECT 132.605 218.335 132.835 224.785 ;
        RECT 137.185 218.335 137.415 224.785 ;
        RECT 141.765 218.335 141.995 224.785 ;
        RECT 146.345 218.335 146.575 224.785 ;
        RECT 150.925 218.335 151.155 224.785 ;
        RECT 155.505 218.335 155.735 224.785 ;
        RECT 160.085 218.335 160.315 224.785 ;
        RECT 164.665 218.335 164.895 224.785 ;
        RECT 169.245 218.335 169.475 224.785 ;
        RECT 173.825 218.335 174.055 224.785 ;
        RECT 178.405 218.335 178.635 224.785 ;
        RECT 182.985 218.335 183.215 224.785 ;
        RECT 187.565 218.335 187.795 224.785 ;
        RECT 192.145 218.335 192.375 224.785 ;
        RECT 196.725 218.335 196.955 224.785 ;
        RECT 201.305 218.335 201.535 224.785 ;
        RECT 205.885 218.335 206.115 224.785 ;
        RECT 210.465 218.335 210.695 224.785 ;
        RECT 16.740 206.860 275.440 207.460 ;
        RECT 124.360 206.325 124.500 206.860 ;
        RECT 124.285 206.095 124.575 206.325 ;
        RECT 163.000 205.985 163.140 206.860 ;
        RECT 115.865 199.535 116.095 205.985 ;
        RECT 120.445 199.535 120.675 205.985 ;
        RECT 125.025 199.535 125.255 205.985 ;
        RECT 129.605 199.535 129.835 205.985 ;
        RECT 134.185 199.535 134.415 205.985 ;
        RECT 138.765 199.535 138.995 205.985 ;
        RECT 149.185 199.820 149.415 205.985 ;
        RECT 147.360 199.680 149.415 199.820 ;
        RECT 147.360 198.800 147.500 199.680 ;
        RECT 149.185 199.535 149.415 199.680 ;
        RECT 153.765 199.535 153.995 205.985 ;
        RECT 158.345 199.535 158.575 205.985 ;
        RECT 162.925 199.535 163.155 205.985 ;
        RECT 167.505 199.535 167.735 205.985 ;
        RECT 172.085 199.535 172.315 205.985 ;
        RECT 141.380 198.660 147.500 198.800 ;
        RECT 141.380 198.505 141.520 198.660 ;
        RECT 141.305 198.275 141.595 198.505 ;
        RECT 16.740 188.060 275.440 188.660 ;
        RECT 187.840 187.625 187.980 188.060 ;
        RECT 187.765 187.395 188.055 187.625 ;
        RECT 189.855 180.735 190.085 187.185 ;
        RECT 194.435 180.735 194.665 187.185 ;
        RECT 199.015 180.735 199.245 187.185 ;
        RECT 16.740 169.260 275.440 169.860 ;
        RECT 16.740 150.460 275.440 151.060 ;
        RECT 201.640 150.025 201.780 150.460 ;
        RECT 201.565 149.795 201.855 150.025 ;
        RECT 189.855 143.135 190.085 149.585 ;
        RECT 194.435 143.135 194.665 149.585 ;
        RECT 199.015 143.135 199.245 149.585 ;
        RECT 16.740 131.660 275.440 132.260 ;
        RECT 16.740 112.860 275.440 113.460 ;
        RECT 16.740 94.060 275.440 94.660 ;
        RECT 126.660 93.185 126.800 94.060 ;
        RECT 126.645 86.735 126.875 93.185 ;
        RECT 131.225 86.735 131.455 93.185 ;
        RECT 135.805 86.735 136.035 93.185 ;
        RECT 140.385 86.735 140.615 93.185 ;
        RECT 144.965 86.735 145.195 93.185 ;
        RECT 149.545 86.735 149.775 93.185 ;
        RECT 154.125 86.735 154.355 93.185 ;
        RECT 158.705 86.735 158.935 93.185 ;
        RECT 163.285 86.735 163.515 93.185 ;
        RECT 167.865 86.735 168.095 93.185 ;
        RECT 172.445 86.735 172.675 93.185 ;
        RECT 177.025 86.735 177.255 93.185 ;
        RECT 181.605 86.735 181.835 93.185 ;
        RECT 186.185 86.735 186.415 93.185 ;
        RECT 190.765 86.735 190.995 93.185 ;
        RECT 195.345 86.735 195.575 93.185 ;
        RECT 199.925 86.735 200.155 93.185 ;
        RECT 204.505 86.735 204.735 93.185 ;
        RECT 209.085 86.735 209.315 93.185 ;
        RECT 213.665 86.735 213.895 93.185 ;
        RECT 218.245 86.735 218.475 93.185 ;
        RECT 222.825 86.735 223.055 93.185 ;
        RECT 227.405 86.735 227.635 93.185 ;
        RECT 231.985 86.735 232.215 93.185 ;
        RECT 236.565 86.735 236.795 93.185 ;
        RECT 241.145 86.735 241.375 93.185 ;
        RECT 245.725 86.735 245.955 93.185 ;
        RECT 250.305 86.735 250.535 93.185 ;
        RECT 254.885 86.735 255.115 93.185 ;
        RECT 259.465 86.735 259.695 93.185 ;
        RECT 16.740 75.260 275.440 75.860 ;
        RECT 16.740 56.460 275.440 57.060 ;
        RECT 16.740 37.660 275.440 38.260 ;
      LAYER via ;
        RECT 16.850 244.470 24.790 245.050 ;
        RECT 267.390 244.470 275.330 245.050 ;
        RECT 16.850 225.670 24.790 226.250 ;
        RECT 267.390 225.670 275.330 226.250 ;
        RECT 16.850 206.870 24.790 207.450 ;
        RECT 267.390 206.870 275.330 207.450 ;
        RECT 16.850 188.070 24.790 188.650 ;
        RECT 167.080 188.060 167.340 188.320 ;
        RECT 267.390 188.070 275.330 188.650 ;
        RECT 16.850 169.270 24.790 169.850 ;
        RECT 167.080 169.360 167.340 169.620 ;
        RECT 267.390 169.270 275.330 169.850 ;
        RECT 16.850 150.470 24.790 151.050 ;
        RECT 167.080 150.660 167.340 150.920 ;
        RECT 267.390 150.470 275.330 151.050 ;
        RECT 16.850 131.670 24.790 132.250 ;
        RECT 167.080 131.960 167.340 132.220 ;
        RECT 267.390 131.670 275.330 132.250 ;
        RECT 16.850 112.870 24.790 113.450 ;
        RECT 267.390 112.870 275.330 113.450 ;
        RECT 16.850 94.070 24.790 94.650 ;
        RECT 267.390 94.070 275.330 94.650 ;
        RECT 16.850 75.270 24.790 75.850 ;
        RECT 267.390 75.270 275.330 75.850 ;
        RECT 16.850 56.470 24.790 57.050 ;
        RECT 267.390 56.470 275.330 57.050 ;
        RECT 16.850 37.670 24.790 38.250 ;
        RECT 267.390 37.670 275.330 38.250 ;
      LAYER met2 ;
        RECT 16.740 244.460 24.900 245.060 ;
        RECT 267.280 244.460 275.440 245.060 ;
        RECT 16.740 225.660 24.900 226.260 ;
        RECT 267.280 225.660 275.440 226.260 ;
        RECT 16.740 206.860 24.900 207.460 ;
        RECT 267.280 206.860 275.440 207.460 ;
        RECT 16.740 188.060 24.900 188.660 ;
        RECT 167.080 188.125 167.340 188.350 ;
        RECT 167.070 187.755 167.350 188.125 ;
        RECT 267.280 188.060 275.440 188.660 ;
        RECT 149.630 186.810 150.630 187.210 ;
        RECT 16.740 169.260 24.900 169.860 ;
        RECT 167.070 168.845 167.350 169.650 ;
        RECT 267.280 169.260 275.440 169.860 ;
        RECT 131.010 168.010 132.010 168.410 ;
        RECT 168.250 168.010 169.250 168.410 ;
        RECT 16.740 150.460 24.900 151.060 ;
        RECT 167.080 150.915 167.340 150.950 ;
        RECT 167.070 150.545 167.350 150.915 ;
        RECT 167.140 150.465 167.280 150.545 ;
        RECT 267.280 150.460 275.440 151.060 ;
        RECT 149.630 149.210 150.630 149.610 ;
        RECT 16.740 131.660 24.900 132.260 ;
        RECT 167.080 132.005 167.340 132.250 ;
        RECT 167.070 131.635 167.350 132.005 ;
        RECT 267.280 131.660 275.440 132.260 ;
        RECT 149.630 130.410 150.630 130.810 ;
        RECT 16.740 112.860 24.900 113.460 ;
        RECT 267.280 112.860 275.440 113.460 ;
        RECT 16.740 94.060 24.900 94.660 ;
        RECT 267.280 94.060 275.440 94.660 ;
        RECT 16.740 75.260 24.900 75.860 ;
        RECT 267.280 75.260 275.440 75.860 ;
        RECT 16.740 56.460 24.900 57.060 ;
        RECT 267.280 56.460 275.440 57.060 ;
        RECT 16.740 37.660 24.900 38.260 ;
        RECT 267.280 37.660 275.440 38.260 ;
      LAYER via2 ;
        RECT 16.880 244.620 17.160 244.900 ;
        RECT 17.280 244.620 17.560 244.900 ;
        RECT 17.680 244.620 17.960 244.900 ;
        RECT 18.080 244.620 18.360 244.900 ;
        RECT 18.480 244.620 18.760 244.900 ;
        RECT 18.880 244.620 19.160 244.900 ;
        RECT 19.280 244.620 19.560 244.900 ;
        RECT 19.680 244.620 19.960 244.900 ;
        RECT 20.080 244.620 20.360 244.900 ;
        RECT 20.480 244.620 20.760 244.900 ;
        RECT 20.880 244.620 21.160 244.900 ;
        RECT 21.280 244.620 21.560 244.900 ;
        RECT 21.680 244.620 21.960 244.900 ;
        RECT 22.080 244.620 22.360 244.900 ;
        RECT 22.480 244.620 22.760 244.900 ;
        RECT 22.880 244.620 23.160 244.900 ;
        RECT 23.280 244.620 23.560 244.900 ;
        RECT 23.680 244.620 23.960 244.900 ;
        RECT 24.080 244.620 24.360 244.900 ;
        RECT 24.480 244.620 24.760 244.900 ;
        RECT 267.420 244.620 267.700 244.900 ;
        RECT 267.820 244.620 268.100 244.900 ;
        RECT 268.220 244.620 268.500 244.900 ;
        RECT 268.620 244.620 268.900 244.900 ;
        RECT 269.020 244.620 269.300 244.900 ;
        RECT 269.420 244.620 269.700 244.900 ;
        RECT 269.820 244.620 270.100 244.900 ;
        RECT 270.220 244.620 270.500 244.900 ;
        RECT 270.620 244.620 270.900 244.900 ;
        RECT 271.020 244.620 271.300 244.900 ;
        RECT 271.420 244.620 271.700 244.900 ;
        RECT 271.820 244.620 272.100 244.900 ;
        RECT 272.220 244.620 272.500 244.900 ;
        RECT 272.620 244.620 272.900 244.900 ;
        RECT 273.020 244.620 273.300 244.900 ;
        RECT 273.420 244.620 273.700 244.900 ;
        RECT 273.820 244.620 274.100 244.900 ;
        RECT 274.220 244.620 274.500 244.900 ;
        RECT 274.620 244.620 274.900 244.900 ;
        RECT 275.020 244.620 275.300 244.900 ;
        RECT 16.880 225.820 17.160 226.100 ;
        RECT 17.280 225.820 17.560 226.100 ;
        RECT 17.680 225.820 17.960 226.100 ;
        RECT 18.080 225.820 18.360 226.100 ;
        RECT 18.480 225.820 18.760 226.100 ;
        RECT 18.880 225.820 19.160 226.100 ;
        RECT 19.280 225.820 19.560 226.100 ;
        RECT 19.680 225.820 19.960 226.100 ;
        RECT 20.080 225.820 20.360 226.100 ;
        RECT 20.480 225.820 20.760 226.100 ;
        RECT 20.880 225.820 21.160 226.100 ;
        RECT 21.280 225.820 21.560 226.100 ;
        RECT 21.680 225.820 21.960 226.100 ;
        RECT 22.080 225.820 22.360 226.100 ;
        RECT 22.480 225.820 22.760 226.100 ;
        RECT 22.880 225.820 23.160 226.100 ;
        RECT 23.280 225.820 23.560 226.100 ;
        RECT 23.680 225.820 23.960 226.100 ;
        RECT 24.080 225.820 24.360 226.100 ;
        RECT 24.480 225.820 24.760 226.100 ;
        RECT 267.420 225.820 267.700 226.100 ;
        RECT 267.820 225.820 268.100 226.100 ;
        RECT 268.220 225.820 268.500 226.100 ;
        RECT 268.620 225.820 268.900 226.100 ;
        RECT 269.020 225.820 269.300 226.100 ;
        RECT 269.420 225.820 269.700 226.100 ;
        RECT 269.820 225.820 270.100 226.100 ;
        RECT 270.220 225.820 270.500 226.100 ;
        RECT 270.620 225.820 270.900 226.100 ;
        RECT 271.020 225.820 271.300 226.100 ;
        RECT 271.420 225.820 271.700 226.100 ;
        RECT 271.820 225.820 272.100 226.100 ;
        RECT 272.220 225.820 272.500 226.100 ;
        RECT 272.620 225.820 272.900 226.100 ;
        RECT 273.020 225.820 273.300 226.100 ;
        RECT 273.420 225.820 273.700 226.100 ;
        RECT 273.820 225.820 274.100 226.100 ;
        RECT 274.220 225.820 274.500 226.100 ;
        RECT 274.620 225.820 274.900 226.100 ;
        RECT 275.020 225.820 275.300 226.100 ;
        RECT 16.880 207.020 17.160 207.300 ;
        RECT 17.280 207.020 17.560 207.300 ;
        RECT 17.680 207.020 17.960 207.300 ;
        RECT 18.080 207.020 18.360 207.300 ;
        RECT 18.480 207.020 18.760 207.300 ;
        RECT 18.880 207.020 19.160 207.300 ;
        RECT 19.280 207.020 19.560 207.300 ;
        RECT 19.680 207.020 19.960 207.300 ;
        RECT 20.080 207.020 20.360 207.300 ;
        RECT 20.480 207.020 20.760 207.300 ;
        RECT 20.880 207.020 21.160 207.300 ;
        RECT 21.280 207.020 21.560 207.300 ;
        RECT 21.680 207.020 21.960 207.300 ;
        RECT 22.080 207.020 22.360 207.300 ;
        RECT 22.480 207.020 22.760 207.300 ;
        RECT 22.880 207.020 23.160 207.300 ;
        RECT 23.280 207.020 23.560 207.300 ;
        RECT 23.680 207.020 23.960 207.300 ;
        RECT 24.080 207.020 24.360 207.300 ;
        RECT 24.480 207.020 24.760 207.300 ;
        RECT 267.420 207.020 267.700 207.300 ;
        RECT 267.820 207.020 268.100 207.300 ;
        RECT 268.220 207.020 268.500 207.300 ;
        RECT 268.620 207.020 268.900 207.300 ;
        RECT 269.020 207.020 269.300 207.300 ;
        RECT 269.420 207.020 269.700 207.300 ;
        RECT 269.820 207.020 270.100 207.300 ;
        RECT 270.220 207.020 270.500 207.300 ;
        RECT 270.620 207.020 270.900 207.300 ;
        RECT 271.020 207.020 271.300 207.300 ;
        RECT 271.420 207.020 271.700 207.300 ;
        RECT 271.820 207.020 272.100 207.300 ;
        RECT 272.220 207.020 272.500 207.300 ;
        RECT 272.620 207.020 272.900 207.300 ;
        RECT 273.020 207.020 273.300 207.300 ;
        RECT 273.420 207.020 273.700 207.300 ;
        RECT 273.820 207.020 274.100 207.300 ;
        RECT 274.220 207.020 274.500 207.300 ;
        RECT 274.620 207.020 274.900 207.300 ;
        RECT 275.020 207.020 275.300 207.300 ;
        RECT 16.880 188.220 17.160 188.500 ;
        RECT 17.280 188.220 17.560 188.500 ;
        RECT 17.680 188.220 17.960 188.500 ;
        RECT 18.080 188.220 18.360 188.500 ;
        RECT 18.480 188.220 18.760 188.500 ;
        RECT 18.880 188.220 19.160 188.500 ;
        RECT 19.280 188.220 19.560 188.500 ;
        RECT 19.680 188.220 19.960 188.500 ;
        RECT 20.080 188.220 20.360 188.500 ;
        RECT 20.480 188.220 20.760 188.500 ;
        RECT 20.880 188.220 21.160 188.500 ;
        RECT 21.280 188.220 21.560 188.500 ;
        RECT 21.680 188.220 21.960 188.500 ;
        RECT 22.080 188.220 22.360 188.500 ;
        RECT 22.480 188.220 22.760 188.500 ;
        RECT 22.880 188.220 23.160 188.500 ;
        RECT 23.280 188.220 23.560 188.500 ;
        RECT 23.680 188.220 23.960 188.500 ;
        RECT 24.080 188.220 24.360 188.500 ;
        RECT 24.480 188.220 24.760 188.500 ;
        RECT 267.420 188.220 267.700 188.500 ;
        RECT 267.820 188.220 268.100 188.500 ;
        RECT 268.220 188.220 268.500 188.500 ;
        RECT 268.620 188.220 268.900 188.500 ;
        RECT 269.020 188.220 269.300 188.500 ;
        RECT 269.420 188.220 269.700 188.500 ;
        RECT 269.820 188.220 270.100 188.500 ;
        RECT 270.220 188.220 270.500 188.500 ;
        RECT 270.620 188.220 270.900 188.500 ;
        RECT 271.020 188.220 271.300 188.500 ;
        RECT 271.420 188.220 271.700 188.500 ;
        RECT 271.820 188.220 272.100 188.500 ;
        RECT 272.220 188.220 272.500 188.500 ;
        RECT 272.620 188.220 272.900 188.500 ;
        RECT 273.020 188.220 273.300 188.500 ;
        RECT 273.420 188.220 273.700 188.500 ;
        RECT 273.820 188.220 274.100 188.500 ;
        RECT 274.220 188.220 274.500 188.500 ;
        RECT 274.620 188.220 274.900 188.500 ;
        RECT 275.020 188.220 275.300 188.500 ;
        RECT 167.070 187.800 167.350 188.080 ;
        RECT 149.790 186.870 150.070 187.150 ;
        RECT 150.190 186.870 150.470 187.150 ;
        RECT 16.880 169.420 17.160 169.700 ;
        RECT 17.280 169.420 17.560 169.700 ;
        RECT 17.680 169.420 17.960 169.700 ;
        RECT 18.080 169.420 18.360 169.700 ;
        RECT 18.480 169.420 18.760 169.700 ;
        RECT 18.880 169.420 19.160 169.700 ;
        RECT 19.280 169.420 19.560 169.700 ;
        RECT 19.680 169.420 19.960 169.700 ;
        RECT 20.080 169.420 20.360 169.700 ;
        RECT 20.480 169.420 20.760 169.700 ;
        RECT 20.880 169.420 21.160 169.700 ;
        RECT 21.280 169.420 21.560 169.700 ;
        RECT 21.680 169.420 21.960 169.700 ;
        RECT 22.080 169.420 22.360 169.700 ;
        RECT 22.480 169.420 22.760 169.700 ;
        RECT 22.880 169.420 23.160 169.700 ;
        RECT 23.280 169.420 23.560 169.700 ;
        RECT 23.680 169.420 23.960 169.700 ;
        RECT 24.080 169.420 24.360 169.700 ;
        RECT 24.480 169.420 24.760 169.700 ;
        RECT 267.420 169.420 267.700 169.700 ;
        RECT 267.820 169.420 268.100 169.700 ;
        RECT 268.220 169.420 268.500 169.700 ;
        RECT 268.620 169.420 268.900 169.700 ;
        RECT 269.020 169.420 269.300 169.700 ;
        RECT 269.420 169.420 269.700 169.700 ;
        RECT 269.820 169.420 270.100 169.700 ;
        RECT 270.220 169.420 270.500 169.700 ;
        RECT 270.620 169.420 270.900 169.700 ;
        RECT 271.020 169.420 271.300 169.700 ;
        RECT 271.420 169.420 271.700 169.700 ;
        RECT 271.820 169.420 272.100 169.700 ;
        RECT 272.220 169.420 272.500 169.700 ;
        RECT 272.620 169.420 272.900 169.700 ;
        RECT 273.020 169.420 273.300 169.700 ;
        RECT 273.420 169.420 273.700 169.700 ;
        RECT 273.820 169.420 274.100 169.700 ;
        RECT 274.220 169.420 274.500 169.700 ;
        RECT 274.620 169.420 274.900 169.700 ;
        RECT 275.020 169.420 275.300 169.700 ;
        RECT 167.070 168.890 167.350 169.170 ;
        RECT 131.170 168.070 131.450 168.350 ;
        RECT 131.570 168.070 131.850 168.350 ;
        RECT 168.410 168.070 168.690 168.350 ;
        RECT 168.810 168.070 169.090 168.350 ;
        RECT 16.880 150.620 17.160 150.900 ;
        RECT 17.280 150.620 17.560 150.900 ;
        RECT 17.680 150.620 17.960 150.900 ;
        RECT 18.080 150.620 18.360 150.900 ;
        RECT 18.480 150.620 18.760 150.900 ;
        RECT 18.880 150.620 19.160 150.900 ;
        RECT 19.280 150.620 19.560 150.900 ;
        RECT 19.680 150.620 19.960 150.900 ;
        RECT 20.080 150.620 20.360 150.900 ;
        RECT 20.480 150.620 20.760 150.900 ;
        RECT 20.880 150.620 21.160 150.900 ;
        RECT 21.280 150.620 21.560 150.900 ;
        RECT 21.680 150.620 21.960 150.900 ;
        RECT 22.080 150.620 22.360 150.900 ;
        RECT 22.480 150.620 22.760 150.900 ;
        RECT 22.880 150.620 23.160 150.900 ;
        RECT 23.280 150.620 23.560 150.900 ;
        RECT 23.680 150.620 23.960 150.900 ;
        RECT 24.080 150.620 24.360 150.900 ;
        RECT 24.480 150.620 24.760 150.900 ;
        RECT 167.070 150.590 167.350 150.870 ;
        RECT 267.420 150.620 267.700 150.900 ;
        RECT 267.820 150.620 268.100 150.900 ;
        RECT 268.220 150.620 268.500 150.900 ;
        RECT 268.620 150.620 268.900 150.900 ;
        RECT 269.020 150.620 269.300 150.900 ;
        RECT 269.420 150.620 269.700 150.900 ;
        RECT 269.820 150.620 270.100 150.900 ;
        RECT 270.220 150.620 270.500 150.900 ;
        RECT 270.620 150.620 270.900 150.900 ;
        RECT 271.020 150.620 271.300 150.900 ;
        RECT 271.420 150.620 271.700 150.900 ;
        RECT 271.820 150.620 272.100 150.900 ;
        RECT 272.220 150.620 272.500 150.900 ;
        RECT 272.620 150.620 272.900 150.900 ;
        RECT 273.020 150.620 273.300 150.900 ;
        RECT 273.420 150.620 273.700 150.900 ;
        RECT 273.820 150.620 274.100 150.900 ;
        RECT 274.220 150.620 274.500 150.900 ;
        RECT 274.620 150.620 274.900 150.900 ;
        RECT 275.020 150.620 275.300 150.900 ;
        RECT 149.790 149.270 150.070 149.550 ;
        RECT 150.190 149.270 150.470 149.550 ;
        RECT 16.880 131.820 17.160 132.100 ;
        RECT 17.280 131.820 17.560 132.100 ;
        RECT 17.680 131.820 17.960 132.100 ;
        RECT 18.080 131.820 18.360 132.100 ;
        RECT 18.480 131.820 18.760 132.100 ;
        RECT 18.880 131.820 19.160 132.100 ;
        RECT 19.280 131.820 19.560 132.100 ;
        RECT 19.680 131.820 19.960 132.100 ;
        RECT 20.080 131.820 20.360 132.100 ;
        RECT 20.480 131.820 20.760 132.100 ;
        RECT 20.880 131.820 21.160 132.100 ;
        RECT 21.280 131.820 21.560 132.100 ;
        RECT 21.680 131.820 21.960 132.100 ;
        RECT 22.080 131.820 22.360 132.100 ;
        RECT 22.480 131.820 22.760 132.100 ;
        RECT 22.880 131.820 23.160 132.100 ;
        RECT 23.280 131.820 23.560 132.100 ;
        RECT 23.680 131.820 23.960 132.100 ;
        RECT 24.080 131.820 24.360 132.100 ;
        RECT 24.480 131.820 24.760 132.100 ;
        RECT 167.070 131.680 167.350 131.960 ;
        RECT 267.420 131.820 267.700 132.100 ;
        RECT 267.820 131.820 268.100 132.100 ;
        RECT 268.220 131.820 268.500 132.100 ;
        RECT 268.620 131.820 268.900 132.100 ;
        RECT 269.020 131.820 269.300 132.100 ;
        RECT 269.420 131.820 269.700 132.100 ;
        RECT 269.820 131.820 270.100 132.100 ;
        RECT 270.220 131.820 270.500 132.100 ;
        RECT 270.620 131.820 270.900 132.100 ;
        RECT 271.020 131.820 271.300 132.100 ;
        RECT 271.420 131.820 271.700 132.100 ;
        RECT 271.820 131.820 272.100 132.100 ;
        RECT 272.220 131.820 272.500 132.100 ;
        RECT 272.620 131.820 272.900 132.100 ;
        RECT 273.020 131.820 273.300 132.100 ;
        RECT 273.420 131.820 273.700 132.100 ;
        RECT 273.820 131.820 274.100 132.100 ;
        RECT 274.220 131.820 274.500 132.100 ;
        RECT 274.620 131.820 274.900 132.100 ;
        RECT 275.020 131.820 275.300 132.100 ;
        RECT 149.790 130.470 150.070 130.750 ;
        RECT 150.190 130.470 150.470 130.750 ;
        RECT 16.880 113.020 17.160 113.300 ;
        RECT 17.280 113.020 17.560 113.300 ;
        RECT 17.680 113.020 17.960 113.300 ;
        RECT 18.080 113.020 18.360 113.300 ;
        RECT 18.480 113.020 18.760 113.300 ;
        RECT 18.880 113.020 19.160 113.300 ;
        RECT 19.280 113.020 19.560 113.300 ;
        RECT 19.680 113.020 19.960 113.300 ;
        RECT 20.080 113.020 20.360 113.300 ;
        RECT 20.480 113.020 20.760 113.300 ;
        RECT 20.880 113.020 21.160 113.300 ;
        RECT 21.280 113.020 21.560 113.300 ;
        RECT 21.680 113.020 21.960 113.300 ;
        RECT 22.080 113.020 22.360 113.300 ;
        RECT 22.480 113.020 22.760 113.300 ;
        RECT 22.880 113.020 23.160 113.300 ;
        RECT 23.280 113.020 23.560 113.300 ;
        RECT 23.680 113.020 23.960 113.300 ;
        RECT 24.080 113.020 24.360 113.300 ;
        RECT 24.480 113.020 24.760 113.300 ;
        RECT 267.420 113.020 267.700 113.300 ;
        RECT 267.820 113.020 268.100 113.300 ;
        RECT 268.220 113.020 268.500 113.300 ;
        RECT 268.620 113.020 268.900 113.300 ;
        RECT 269.020 113.020 269.300 113.300 ;
        RECT 269.420 113.020 269.700 113.300 ;
        RECT 269.820 113.020 270.100 113.300 ;
        RECT 270.220 113.020 270.500 113.300 ;
        RECT 270.620 113.020 270.900 113.300 ;
        RECT 271.020 113.020 271.300 113.300 ;
        RECT 271.420 113.020 271.700 113.300 ;
        RECT 271.820 113.020 272.100 113.300 ;
        RECT 272.220 113.020 272.500 113.300 ;
        RECT 272.620 113.020 272.900 113.300 ;
        RECT 273.020 113.020 273.300 113.300 ;
        RECT 273.420 113.020 273.700 113.300 ;
        RECT 273.820 113.020 274.100 113.300 ;
        RECT 274.220 113.020 274.500 113.300 ;
        RECT 274.620 113.020 274.900 113.300 ;
        RECT 275.020 113.020 275.300 113.300 ;
        RECT 16.880 94.220 17.160 94.500 ;
        RECT 17.280 94.220 17.560 94.500 ;
        RECT 17.680 94.220 17.960 94.500 ;
        RECT 18.080 94.220 18.360 94.500 ;
        RECT 18.480 94.220 18.760 94.500 ;
        RECT 18.880 94.220 19.160 94.500 ;
        RECT 19.280 94.220 19.560 94.500 ;
        RECT 19.680 94.220 19.960 94.500 ;
        RECT 20.080 94.220 20.360 94.500 ;
        RECT 20.480 94.220 20.760 94.500 ;
        RECT 20.880 94.220 21.160 94.500 ;
        RECT 21.280 94.220 21.560 94.500 ;
        RECT 21.680 94.220 21.960 94.500 ;
        RECT 22.080 94.220 22.360 94.500 ;
        RECT 22.480 94.220 22.760 94.500 ;
        RECT 22.880 94.220 23.160 94.500 ;
        RECT 23.280 94.220 23.560 94.500 ;
        RECT 23.680 94.220 23.960 94.500 ;
        RECT 24.080 94.220 24.360 94.500 ;
        RECT 24.480 94.220 24.760 94.500 ;
        RECT 267.420 94.220 267.700 94.500 ;
        RECT 267.820 94.220 268.100 94.500 ;
        RECT 268.220 94.220 268.500 94.500 ;
        RECT 268.620 94.220 268.900 94.500 ;
        RECT 269.020 94.220 269.300 94.500 ;
        RECT 269.420 94.220 269.700 94.500 ;
        RECT 269.820 94.220 270.100 94.500 ;
        RECT 270.220 94.220 270.500 94.500 ;
        RECT 270.620 94.220 270.900 94.500 ;
        RECT 271.020 94.220 271.300 94.500 ;
        RECT 271.420 94.220 271.700 94.500 ;
        RECT 271.820 94.220 272.100 94.500 ;
        RECT 272.220 94.220 272.500 94.500 ;
        RECT 272.620 94.220 272.900 94.500 ;
        RECT 273.020 94.220 273.300 94.500 ;
        RECT 273.420 94.220 273.700 94.500 ;
        RECT 273.820 94.220 274.100 94.500 ;
        RECT 274.220 94.220 274.500 94.500 ;
        RECT 274.620 94.220 274.900 94.500 ;
        RECT 275.020 94.220 275.300 94.500 ;
        RECT 16.880 75.420 17.160 75.700 ;
        RECT 17.280 75.420 17.560 75.700 ;
        RECT 17.680 75.420 17.960 75.700 ;
        RECT 18.080 75.420 18.360 75.700 ;
        RECT 18.480 75.420 18.760 75.700 ;
        RECT 18.880 75.420 19.160 75.700 ;
        RECT 19.280 75.420 19.560 75.700 ;
        RECT 19.680 75.420 19.960 75.700 ;
        RECT 20.080 75.420 20.360 75.700 ;
        RECT 20.480 75.420 20.760 75.700 ;
        RECT 20.880 75.420 21.160 75.700 ;
        RECT 21.280 75.420 21.560 75.700 ;
        RECT 21.680 75.420 21.960 75.700 ;
        RECT 22.080 75.420 22.360 75.700 ;
        RECT 22.480 75.420 22.760 75.700 ;
        RECT 22.880 75.420 23.160 75.700 ;
        RECT 23.280 75.420 23.560 75.700 ;
        RECT 23.680 75.420 23.960 75.700 ;
        RECT 24.080 75.420 24.360 75.700 ;
        RECT 24.480 75.420 24.760 75.700 ;
        RECT 267.420 75.420 267.700 75.700 ;
        RECT 267.820 75.420 268.100 75.700 ;
        RECT 268.220 75.420 268.500 75.700 ;
        RECT 268.620 75.420 268.900 75.700 ;
        RECT 269.020 75.420 269.300 75.700 ;
        RECT 269.420 75.420 269.700 75.700 ;
        RECT 269.820 75.420 270.100 75.700 ;
        RECT 270.220 75.420 270.500 75.700 ;
        RECT 270.620 75.420 270.900 75.700 ;
        RECT 271.020 75.420 271.300 75.700 ;
        RECT 271.420 75.420 271.700 75.700 ;
        RECT 271.820 75.420 272.100 75.700 ;
        RECT 272.220 75.420 272.500 75.700 ;
        RECT 272.620 75.420 272.900 75.700 ;
        RECT 273.020 75.420 273.300 75.700 ;
        RECT 273.420 75.420 273.700 75.700 ;
        RECT 273.820 75.420 274.100 75.700 ;
        RECT 274.220 75.420 274.500 75.700 ;
        RECT 274.620 75.420 274.900 75.700 ;
        RECT 275.020 75.420 275.300 75.700 ;
        RECT 16.880 56.620 17.160 56.900 ;
        RECT 17.280 56.620 17.560 56.900 ;
        RECT 17.680 56.620 17.960 56.900 ;
        RECT 18.080 56.620 18.360 56.900 ;
        RECT 18.480 56.620 18.760 56.900 ;
        RECT 18.880 56.620 19.160 56.900 ;
        RECT 19.280 56.620 19.560 56.900 ;
        RECT 19.680 56.620 19.960 56.900 ;
        RECT 20.080 56.620 20.360 56.900 ;
        RECT 20.480 56.620 20.760 56.900 ;
        RECT 20.880 56.620 21.160 56.900 ;
        RECT 21.280 56.620 21.560 56.900 ;
        RECT 21.680 56.620 21.960 56.900 ;
        RECT 22.080 56.620 22.360 56.900 ;
        RECT 22.480 56.620 22.760 56.900 ;
        RECT 22.880 56.620 23.160 56.900 ;
        RECT 23.280 56.620 23.560 56.900 ;
        RECT 23.680 56.620 23.960 56.900 ;
        RECT 24.080 56.620 24.360 56.900 ;
        RECT 24.480 56.620 24.760 56.900 ;
        RECT 267.420 56.620 267.700 56.900 ;
        RECT 267.820 56.620 268.100 56.900 ;
        RECT 268.220 56.620 268.500 56.900 ;
        RECT 268.620 56.620 268.900 56.900 ;
        RECT 269.020 56.620 269.300 56.900 ;
        RECT 269.420 56.620 269.700 56.900 ;
        RECT 269.820 56.620 270.100 56.900 ;
        RECT 270.220 56.620 270.500 56.900 ;
        RECT 270.620 56.620 270.900 56.900 ;
        RECT 271.020 56.620 271.300 56.900 ;
        RECT 271.420 56.620 271.700 56.900 ;
        RECT 271.820 56.620 272.100 56.900 ;
        RECT 272.220 56.620 272.500 56.900 ;
        RECT 272.620 56.620 272.900 56.900 ;
        RECT 273.020 56.620 273.300 56.900 ;
        RECT 273.420 56.620 273.700 56.900 ;
        RECT 273.820 56.620 274.100 56.900 ;
        RECT 274.220 56.620 274.500 56.900 ;
        RECT 274.620 56.620 274.900 56.900 ;
        RECT 275.020 56.620 275.300 56.900 ;
        RECT 16.880 37.820 17.160 38.100 ;
        RECT 17.280 37.820 17.560 38.100 ;
        RECT 17.680 37.820 17.960 38.100 ;
        RECT 18.080 37.820 18.360 38.100 ;
        RECT 18.480 37.820 18.760 38.100 ;
        RECT 18.880 37.820 19.160 38.100 ;
        RECT 19.280 37.820 19.560 38.100 ;
        RECT 19.680 37.820 19.960 38.100 ;
        RECT 20.080 37.820 20.360 38.100 ;
        RECT 20.480 37.820 20.760 38.100 ;
        RECT 20.880 37.820 21.160 38.100 ;
        RECT 21.280 37.820 21.560 38.100 ;
        RECT 21.680 37.820 21.960 38.100 ;
        RECT 22.080 37.820 22.360 38.100 ;
        RECT 22.480 37.820 22.760 38.100 ;
        RECT 22.880 37.820 23.160 38.100 ;
        RECT 23.280 37.820 23.560 38.100 ;
        RECT 23.680 37.820 23.960 38.100 ;
        RECT 24.080 37.820 24.360 38.100 ;
        RECT 24.480 37.820 24.760 38.100 ;
        RECT 267.420 37.820 267.700 38.100 ;
        RECT 267.820 37.820 268.100 38.100 ;
        RECT 268.220 37.820 268.500 38.100 ;
        RECT 268.620 37.820 268.900 38.100 ;
        RECT 269.020 37.820 269.300 38.100 ;
        RECT 269.420 37.820 269.700 38.100 ;
        RECT 269.820 37.820 270.100 38.100 ;
        RECT 270.220 37.820 270.500 38.100 ;
        RECT 270.620 37.820 270.900 38.100 ;
        RECT 271.020 37.820 271.300 38.100 ;
        RECT 271.420 37.820 271.700 38.100 ;
        RECT 271.820 37.820 272.100 38.100 ;
        RECT 272.220 37.820 272.500 38.100 ;
        RECT 272.620 37.820 272.900 38.100 ;
        RECT 273.020 37.820 273.300 38.100 ;
        RECT 273.420 37.820 273.700 38.100 ;
        RECT 273.820 37.820 274.100 38.100 ;
        RECT 274.220 37.820 274.500 38.100 ;
        RECT 274.620 37.820 274.900 38.100 ;
        RECT 275.020 37.820 275.300 38.100 ;
      LAYER met3 ;
        RECT 16.740 244.460 24.900 245.060 ;
        RECT 267.280 244.460 275.440 245.060 ;
        RECT 16.740 225.660 24.900 226.260 ;
        RECT 267.280 225.660 275.440 226.260 ;
        RECT 16.740 206.860 24.900 207.460 ;
        RECT 267.280 206.860 275.440 207.460 ;
        RECT 16.740 188.060 24.900 188.660 ;
        RECT 167.045 188.100 167.375 188.105 ;
        RECT 167.020 188.090 167.400 188.100 ;
        RECT 166.600 187.790 167.400 188.090 ;
        RECT 267.280 188.060 275.440 188.660 ;
        RECT 167.020 187.780 167.400 187.790 ;
        RECT 167.045 187.775 167.375 187.780 ;
        RECT 149.630 180.710 185.490 187.210 ;
        RECT 16.740 169.260 24.900 169.860 ;
        RECT 267.280 169.260 275.440 169.860 ;
        RECT 166.330 169.180 166.710 169.190 ;
        RECT 167.045 169.180 167.375 169.195 ;
        RECT 170.470 169.180 170.850 169.190 ;
        RECT 166.330 168.880 170.850 169.180 ;
        RECT 166.330 168.870 166.710 168.880 ;
        RECT 167.045 168.865 167.375 168.880 ;
        RECT 170.470 168.870 170.850 168.880 ;
        RECT 131.010 161.910 166.870 168.410 ;
        RECT 168.250 161.910 204.110 168.410 ;
        RECT 16.740 150.460 24.900 151.060 ;
        RECT 167.045 150.890 167.375 150.895 ;
        RECT 167.020 150.880 167.400 150.890 ;
        RECT 166.600 150.580 167.400 150.880 ;
        RECT 167.020 150.570 167.400 150.580 ;
        RECT 167.045 150.565 167.375 150.570 ;
        RECT 267.280 150.460 275.440 151.060 ;
        RECT 149.630 143.110 185.490 149.610 ;
        RECT 16.740 131.660 24.900 132.260 ;
        RECT 167.045 131.980 167.375 131.985 ;
        RECT 167.020 131.970 167.400 131.980 ;
        RECT 166.600 131.670 167.400 131.970 ;
        RECT 167.020 131.660 167.400 131.670 ;
        RECT 267.280 131.660 275.440 132.260 ;
        RECT 167.045 131.655 167.375 131.660 ;
        RECT 149.630 124.310 185.490 130.810 ;
        RECT 16.740 112.860 24.900 113.460 ;
        RECT 267.280 112.860 275.440 113.460 ;
        RECT 16.740 94.060 24.900 94.660 ;
        RECT 267.280 94.060 275.440 94.660 ;
        RECT 16.740 75.260 24.900 75.860 ;
        RECT 267.280 75.260 275.440 75.860 ;
        RECT 16.740 56.460 24.900 57.060 ;
        RECT 267.280 56.460 275.440 57.060 ;
        RECT 16.740 37.660 24.900 38.260 ;
        RECT 267.280 37.660 275.440 38.260 ;
      LAYER via3 ;
        RECT 16.860 244.600 17.180 244.920 ;
        RECT 17.260 244.600 17.580 244.920 ;
        RECT 17.660 244.600 17.980 244.920 ;
        RECT 18.060 244.600 18.380 244.920 ;
        RECT 18.460 244.600 18.780 244.920 ;
        RECT 18.860 244.600 19.180 244.920 ;
        RECT 19.260 244.600 19.580 244.920 ;
        RECT 19.660 244.600 19.980 244.920 ;
        RECT 20.060 244.600 20.380 244.920 ;
        RECT 20.460 244.600 20.780 244.920 ;
        RECT 20.860 244.600 21.180 244.920 ;
        RECT 21.260 244.600 21.580 244.920 ;
        RECT 21.660 244.600 21.980 244.920 ;
        RECT 22.060 244.600 22.380 244.920 ;
        RECT 22.460 244.600 22.780 244.920 ;
        RECT 22.860 244.600 23.180 244.920 ;
        RECT 23.260 244.600 23.580 244.920 ;
        RECT 23.660 244.600 23.980 244.920 ;
        RECT 24.060 244.600 24.380 244.920 ;
        RECT 24.460 244.600 24.780 244.920 ;
        RECT 267.400 244.600 267.720 244.920 ;
        RECT 267.800 244.600 268.120 244.920 ;
        RECT 268.200 244.600 268.520 244.920 ;
        RECT 268.600 244.600 268.920 244.920 ;
        RECT 269.000 244.600 269.320 244.920 ;
        RECT 269.400 244.600 269.720 244.920 ;
        RECT 269.800 244.600 270.120 244.920 ;
        RECT 270.200 244.600 270.520 244.920 ;
        RECT 270.600 244.600 270.920 244.920 ;
        RECT 271.000 244.600 271.320 244.920 ;
        RECT 271.400 244.600 271.720 244.920 ;
        RECT 271.800 244.600 272.120 244.920 ;
        RECT 272.200 244.600 272.520 244.920 ;
        RECT 272.600 244.600 272.920 244.920 ;
        RECT 273.000 244.600 273.320 244.920 ;
        RECT 273.400 244.600 273.720 244.920 ;
        RECT 273.800 244.600 274.120 244.920 ;
        RECT 274.200 244.600 274.520 244.920 ;
        RECT 274.600 244.600 274.920 244.920 ;
        RECT 275.000 244.600 275.320 244.920 ;
        RECT 16.860 225.800 17.180 226.120 ;
        RECT 17.260 225.800 17.580 226.120 ;
        RECT 17.660 225.800 17.980 226.120 ;
        RECT 18.060 225.800 18.380 226.120 ;
        RECT 18.460 225.800 18.780 226.120 ;
        RECT 18.860 225.800 19.180 226.120 ;
        RECT 19.260 225.800 19.580 226.120 ;
        RECT 19.660 225.800 19.980 226.120 ;
        RECT 20.060 225.800 20.380 226.120 ;
        RECT 20.460 225.800 20.780 226.120 ;
        RECT 20.860 225.800 21.180 226.120 ;
        RECT 21.260 225.800 21.580 226.120 ;
        RECT 21.660 225.800 21.980 226.120 ;
        RECT 22.060 225.800 22.380 226.120 ;
        RECT 22.460 225.800 22.780 226.120 ;
        RECT 22.860 225.800 23.180 226.120 ;
        RECT 23.260 225.800 23.580 226.120 ;
        RECT 23.660 225.800 23.980 226.120 ;
        RECT 24.060 225.800 24.380 226.120 ;
        RECT 24.460 225.800 24.780 226.120 ;
        RECT 267.400 225.800 267.720 226.120 ;
        RECT 267.800 225.800 268.120 226.120 ;
        RECT 268.200 225.800 268.520 226.120 ;
        RECT 268.600 225.800 268.920 226.120 ;
        RECT 269.000 225.800 269.320 226.120 ;
        RECT 269.400 225.800 269.720 226.120 ;
        RECT 269.800 225.800 270.120 226.120 ;
        RECT 270.200 225.800 270.520 226.120 ;
        RECT 270.600 225.800 270.920 226.120 ;
        RECT 271.000 225.800 271.320 226.120 ;
        RECT 271.400 225.800 271.720 226.120 ;
        RECT 271.800 225.800 272.120 226.120 ;
        RECT 272.200 225.800 272.520 226.120 ;
        RECT 272.600 225.800 272.920 226.120 ;
        RECT 273.000 225.800 273.320 226.120 ;
        RECT 273.400 225.800 273.720 226.120 ;
        RECT 273.800 225.800 274.120 226.120 ;
        RECT 274.200 225.800 274.520 226.120 ;
        RECT 274.600 225.800 274.920 226.120 ;
        RECT 275.000 225.800 275.320 226.120 ;
        RECT 16.860 207.000 17.180 207.320 ;
        RECT 17.260 207.000 17.580 207.320 ;
        RECT 17.660 207.000 17.980 207.320 ;
        RECT 18.060 207.000 18.380 207.320 ;
        RECT 18.460 207.000 18.780 207.320 ;
        RECT 18.860 207.000 19.180 207.320 ;
        RECT 19.260 207.000 19.580 207.320 ;
        RECT 19.660 207.000 19.980 207.320 ;
        RECT 20.060 207.000 20.380 207.320 ;
        RECT 20.460 207.000 20.780 207.320 ;
        RECT 20.860 207.000 21.180 207.320 ;
        RECT 21.260 207.000 21.580 207.320 ;
        RECT 21.660 207.000 21.980 207.320 ;
        RECT 22.060 207.000 22.380 207.320 ;
        RECT 22.460 207.000 22.780 207.320 ;
        RECT 22.860 207.000 23.180 207.320 ;
        RECT 23.260 207.000 23.580 207.320 ;
        RECT 23.660 207.000 23.980 207.320 ;
        RECT 24.060 207.000 24.380 207.320 ;
        RECT 24.460 207.000 24.780 207.320 ;
        RECT 267.400 207.000 267.720 207.320 ;
        RECT 267.800 207.000 268.120 207.320 ;
        RECT 268.200 207.000 268.520 207.320 ;
        RECT 268.600 207.000 268.920 207.320 ;
        RECT 269.000 207.000 269.320 207.320 ;
        RECT 269.400 207.000 269.720 207.320 ;
        RECT 269.800 207.000 270.120 207.320 ;
        RECT 270.200 207.000 270.520 207.320 ;
        RECT 270.600 207.000 270.920 207.320 ;
        RECT 271.000 207.000 271.320 207.320 ;
        RECT 271.400 207.000 271.720 207.320 ;
        RECT 271.800 207.000 272.120 207.320 ;
        RECT 272.200 207.000 272.520 207.320 ;
        RECT 272.600 207.000 272.920 207.320 ;
        RECT 273.000 207.000 273.320 207.320 ;
        RECT 273.400 207.000 273.720 207.320 ;
        RECT 273.800 207.000 274.120 207.320 ;
        RECT 274.200 207.000 274.520 207.320 ;
        RECT 274.600 207.000 274.920 207.320 ;
        RECT 275.000 207.000 275.320 207.320 ;
        RECT 16.860 188.200 17.180 188.520 ;
        RECT 17.260 188.200 17.580 188.520 ;
        RECT 17.660 188.200 17.980 188.520 ;
        RECT 18.060 188.200 18.380 188.520 ;
        RECT 18.460 188.200 18.780 188.520 ;
        RECT 18.860 188.200 19.180 188.520 ;
        RECT 19.260 188.200 19.580 188.520 ;
        RECT 19.660 188.200 19.980 188.520 ;
        RECT 20.060 188.200 20.380 188.520 ;
        RECT 20.460 188.200 20.780 188.520 ;
        RECT 20.860 188.200 21.180 188.520 ;
        RECT 21.260 188.200 21.580 188.520 ;
        RECT 21.660 188.200 21.980 188.520 ;
        RECT 22.060 188.200 22.380 188.520 ;
        RECT 22.460 188.200 22.780 188.520 ;
        RECT 22.860 188.200 23.180 188.520 ;
        RECT 23.260 188.200 23.580 188.520 ;
        RECT 23.660 188.200 23.980 188.520 ;
        RECT 24.060 188.200 24.380 188.520 ;
        RECT 24.460 188.200 24.780 188.520 ;
        RECT 267.400 188.200 267.720 188.520 ;
        RECT 267.800 188.200 268.120 188.520 ;
        RECT 268.200 188.200 268.520 188.520 ;
        RECT 268.600 188.200 268.920 188.520 ;
        RECT 269.000 188.200 269.320 188.520 ;
        RECT 269.400 188.200 269.720 188.520 ;
        RECT 269.800 188.200 270.120 188.520 ;
        RECT 270.200 188.200 270.520 188.520 ;
        RECT 270.600 188.200 270.920 188.520 ;
        RECT 271.000 188.200 271.320 188.520 ;
        RECT 271.400 188.200 271.720 188.520 ;
        RECT 271.800 188.200 272.120 188.520 ;
        RECT 272.200 188.200 272.520 188.520 ;
        RECT 272.600 188.200 272.920 188.520 ;
        RECT 273.000 188.200 273.320 188.520 ;
        RECT 273.400 188.200 273.720 188.520 ;
        RECT 273.800 188.200 274.120 188.520 ;
        RECT 274.200 188.200 274.520 188.520 ;
        RECT 274.600 188.200 274.920 188.520 ;
        RECT 275.000 188.200 275.320 188.520 ;
        RECT 167.050 187.780 167.370 188.100 ;
        RECT 152.710 186.750 153.030 187.070 ;
        RECT 156.305 186.750 156.625 187.070 ;
        RECT 159.900 186.750 160.220 187.070 ;
        RECT 163.495 186.750 163.815 187.070 ;
        RECT 167.090 186.750 167.410 187.070 ;
        RECT 170.685 186.750 171.005 187.070 ;
        RECT 174.280 186.750 174.600 187.070 ;
        RECT 177.875 186.750 178.195 187.070 ;
        RECT 181.470 186.750 181.790 187.070 ;
        RECT 185.065 186.750 185.385 187.070 ;
        RECT 152.710 186.350 153.030 186.670 ;
        RECT 156.305 186.350 156.625 186.670 ;
        RECT 159.900 186.350 160.220 186.670 ;
        RECT 163.495 186.350 163.815 186.670 ;
        RECT 167.090 186.350 167.410 186.670 ;
        RECT 170.685 186.350 171.005 186.670 ;
        RECT 174.280 186.350 174.600 186.670 ;
        RECT 177.875 186.350 178.195 186.670 ;
        RECT 181.470 186.350 181.790 186.670 ;
        RECT 185.065 186.350 185.385 186.670 ;
        RECT 152.710 185.950 153.030 186.270 ;
        RECT 156.305 185.950 156.625 186.270 ;
        RECT 159.900 185.950 160.220 186.270 ;
        RECT 163.495 185.950 163.815 186.270 ;
        RECT 167.090 185.950 167.410 186.270 ;
        RECT 170.685 185.950 171.005 186.270 ;
        RECT 174.280 185.950 174.600 186.270 ;
        RECT 177.875 185.950 178.195 186.270 ;
        RECT 181.470 185.950 181.790 186.270 ;
        RECT 185.065 185.950 185.385 186.270 ;
        RECT 152.710 185.550 153.030 185.870 ;
        RECT 156.305 185.550 156.625 185.870 ;
        RECT 159.900 185.550 160.220 185.870 ;
        RECT 163.495 185.550 163.815 185.870 ;
        RECT 167.090 185.550 167.410 185.870 ;
        RECT 170.685 185.550 171.005 185.870 ;
        RECT 174.280 185.550 174.600 185.870 ;
        RECT 177.875 185.550 178.195 185.870 ;
        RECT 181.470 185.550 181.790 185.870 ;
        RECT 185.065 185.550 185.385 185.870 ;
        RECT 152.710 185.150 153.030 185.470 ;
        RECT 156.305 185.150 156.625 185.470 ;
        RECT 159.900 185.150 160.220 185.470 ;
        RECT 163.495 185.150 163.815 185.470 ;
        RECT 167.090 185.150 167.410 185.470 ;
        RECT 170.685 185.150 171.005 185.470 ;
        RECT 174.280 185.150 174.600 185.470 ;
        RECT 177.875 185.150 178.195 185.470 ;
        RECT 181.470 185.150 181.790 185.470 ;
        RECT 185.065 185.150 185.385 185.470 ;
        RECT 152.710 184.750 153.030 185.070 ;
        RECT 156.305 184.750 156.625 185.070 ;
        RECT 159.900 184.750 160.220 185.070 ;
        RECT 163.495 184.750 163.815 185.070 ;
        RECT 167.090 184.750 167.410 185.070 ;
        RECT 170.685 184.750 171.005 185.070 ;
        RECT 174.280 184.750 174.600 185.070 ;
        RECT 177.875 184.750 178.195 185.070 ;
        RECT 181.470 184.750 181.790 185.070 ;
        RECT 185.065 184.750 185.385 185.070 ;
        RECT 152.710 184.350 153.030 184.670 ;
        RECT 156.305 184.350 156.625 184.670 ;
        RECT 159.900 184.350 160.220 184.670 ;
        RECT 163.495 184.350 163.815 184.670 ;
        RECT 167.090 184.350 167.410 184.670 ;
        RECT 170.685 184.350 171.005 184.670 ;
        RECT 174.280 184.350 174.600 184.670 ;
        RECT 177.875 184.350 178.195 184.670 ;
        RECT 181.470 184.350 181.790 184.670 ;
        RECT 185.065 184.350 185.385 184.670 ;
        RECT 152.710 183.250 153.030 183.570 ;
        RECT 156.305 183.250 156.625 183.570 ;
        RECT 159.900 183.250 160.220 183.570 ;
        RECT 163.495 183.250 163.815 183.570 ;
        RECT 167.090 183.250 167.410 183.570 ;
        RECT 170.685 183.250 171.005 183.570 ;
        RECT 174.280 183.250 174.600 183.570 ;
        RECT 177.875 183.250 178.195 183.570 ;
        RECT 181.470 183.250 181.790 183.570 ;
        RECT 185.065 183.250 185.385 183.570 ;
        RECT 152.710 182.850 153.030 183.170 ;
        RECT 156.305 182.850 156.625 183.170 ;
        RECT 159.900 182.850 160.220 183.170 ;
        RECT 163.495 182.850 163.815 183.170 ;
        RECT 167.090 182.850 167.410 183.170 ;
        RECT 170.685 182.850 171.005 183.170 ;
        RECT 174.280 182.850 174.600 183.170 ;
        RECT 177.875 182.850 178.195 183.170 ;
        RECT 181.470 182.850 181.790 183.170 ;
        RECT 185.065 182.850 185.385 183.170 ;
        RECT 152.710 182.450 153.030 182.770 ;
        RECT 156.305 182.450 156.625 182.770 ;
        RECT 159.900 182.450 160.220 182.770 ;
        RECT 163.495 182.450 163.815 182.770 ;
        RECT 167.090 182.450 167.410 182.770 ;
        RECT 170.685 182.450 171.005 182.770 ;
        RECT 174.280 182.450 174.600 182.770 ;
        RECT 177.875 182.450 178.195 182.770 ;
        RECT 181.470 182.450 181.790 182.770 ;
        RECT 185.065 182.450 185.385 182.770 ;
        RECT 152.710 182.050 153.030 182.370 ;
        RECT 156.305 182.050 156.625 182.370 ;
        RECT 159.900 182.050 160.220 182.370 ;
        RECT 163.495 182.050 163.815 182.370 ;
        RECT 167.090 182.050 167.410 182.370 ;
        RECT 170.685 182.050 171.005 182.370 ;
        RECT 174.280 182.050 174.600 182.370 ;
        RECT 177.875 182.050 178.195 182.370 ;
        RECT 181.470 182.050 181.790 182.370 ;
        RECT 185.065 182.050 185.385 182.370 ;
        RECT 152.710 181.650 153.030 181.970 ;
        RECT 156.305 181.650 156.625 181.970 ;
        RECT 159.900 181.650 160.220 181.970 ;
        RECT 163.495 181.650 163.815 181.970 ;
        RECT 167.090 181.650 167.410 181.970 ;
        RECT 170.685 181.650 171.005 181.970 ;
        RECT 174.280 181.650 174.600 181.970 ;
        RECT 177.875 181.650 178.195 181.970 ;
        RECT 181.470 181.650 181.790 181.970 ;
        RECT 185.065 181.650 185.385 181.970 ;
        RECT 152.710 181.250 153.030 181.570 ;
        RECT 156.305 181.250 156.625 181.570 ;
        RECT 159.900 181.250 160.220 181.570 ;
        RECT 163.495 181.250 163.815 181.570 ;
        RECT 167.090 181.250 167.410 181.570 ;
        RECT 170.685 181.250 171.005 181.570 ;
        RECT 174.280 181.250 174.600 181.570 ;
        RECT 177.875 181.250 178.195 181.570 ;
        RECT 181.470 181.250 181.790 181.570 ;
        RECT 185.065 181.250 185.385 181.570 ;
        RECT 152.710 180.850 153.030 181.170 ;
        RECT 156.305 180.850 156.625 181.170 ;
        RECT 159.900 180.850 160.220 181.170 ;
        RECT 163.495 180.850 163.815 181.170 ;
        RECT 167.090 180.850 167.410 181.170 ;
        RECT 170.685 180.850 171.005 181.170 ;
        RECT 174.280 180.850 174.600 181.170 ;
        RECT 177.875 180.850 178.195 181.170 ;
        RECT 181.470 180.850 181.790 181.170 ;
        RECT 185.065 180.850 185.385 181.170 ;
        RECT 16.860 169.400 17.180 169.720 ;
        RECT 17.260 169.400 17.580 169.720 ;
        RECT 17.660 169.400 17.980 169.720 ;
        RECT 18.060 169.400 18.380 169.720 ;
        RECT 18.460 169.400 18.780 169.720 ;
        RECT 18.860 169.400 19.180 169.720 ;
        RECT 19.260 169.400 19.580 169.720 ;
        RECT 19.660 169.400 19.980 169.720 ;
        RECT 20.060 169.400 20.380 169.720 ;
        RECT 20.460 169.400 20.780 169.720 ;
        RECT 20.860 169.400 21.180 169.720 ;
        RECT 21.260 169.400 21.580 169.720 ;
        RECT 21.660 169.400 21.980 169.720 ;
        RECT 22.060 169.400 22.380 169.720 ;
        RECT 22.460 169.400 22.780 169.720 ;
        RECT 22.860 169.400 23.180 169.720 ;
        RECT 23.260 169.400 23.580 169.720 ;
        RECT 23.660 169.400 23.980 169.720 ;
        RECT 24.060 169.400 24.380 169.720 ;
        RECT 24.460 169.400 24.780 169.720 ;
        RECT 267.400 169.400 267.720 169.720 ;
        RECT 267.800 169.400 268.120 169.720 ;
        RECT 268.200 169.400 268.520 169.720 ;
        RECT 268.600 169.400 268.920 169.720 ;
        RECT 269.000 169.400 269.320 169.720 ;
        RECT 269.400 169.400 269.720 169.720 ;
        RECT 269.800 169.400 270.120 169.720 ;
        RECT 270.200 169.400 270.520 169.720 ;
        RECT 270.600 169.400 270.920 169.720 ;
        RECT 271.000 169.400 271.320 169.720 ;
        RECT 271.400 169.400 271.720 169.720 ;
        RECT 271.800 169.400 272.120 169.720 ;
        RECT 272.200 169.400 272.520 169.720 ;
        RECT 272.600 169.400 272.920 169.720 ;
        RECT 273.000 169.400 273.320 169.720 ;
        RECT 273.400 169.400 273.720 169.720 ;
        RECT 273.800 169.400 274.120 169.720 ;
        RECT 274.200 169.400 274.520 169.720 ;
        RECT 274.600 169.400 274.920 169.720 ;
        RECT 275.000 169.400 275.320 169.720 ;
        RECT 166.360 168.870 166.680 169.190 ;
        RECT 170.500 168.870 170.820 169.190 ;
        RECT 134.090 167.950 134.410 168.270 ;
        RECT 137.685 167.950 138.005 168.270 ;
        RECT 141.280 167.950 141.600 168.270 ;
        RECT 144.875 167.950 145.195 168.270 ;
        RECT 148.470 167.950 148.790 168.270 ;
        RECT 152.065 167.950 152.385 168.270 ;
        RECT 155.660 167.950 155.980 168.270 ;
        RECT 159.255 167.950 159.575 168.270 ;
        RECT 162.850 167.950 163.170 168.270 ;
        RECT 166.445 167.950 166.765 168.270 ;
        RECT 134.090 167.550 134.410 167.870 ;
        RECT 137.685 167.550 138.005 167.870 ;
        RECT 141.280 167.550 141.600 167.870 ;
        RECT 144.875 167.550 145.195 167.870 ;
        RECT 148.470 167.550 148.790 167.870 ;
        RECT 152.065 167.550 152.385 167.870 ;
        RECT 155.660 167.550 155.980 167.870 ;
        RECT 159.255 167.550 159.575 167.870 ;
        RECT 162.850 167.550 163.170 167.870 ;
        RECT 166.445 167.550 166.765 167.870 ;
        RECT 134.090 167.150 134.410 167.470 ;
        RECT 137.685 167.150 138.005 167.470 ;
        RECT 141.280 167.150 141.600 167.470 ;
        RECT 144.875 167.150 145.195 167.470 ;
        RECT 148.470 167.150 148.790 167.470 ;
        RECT 152.065 167.150 152.385 167.470 ;
        RECT 155.660 167.150 155.980 167.470 ;
        RECT 159.255 167.150 159.575 167.470 ;
        RECT 162.850 167.150 163.170 167.470 ;
        RECT 166.445 167.150 166.765 167.470 ;
        RECT 134.090 166.750 134.410 167.070 ;
        RECT 137.685 166.750 138.005 167.070 ;
        RECT 141.280 166.750 141.600 167.070 ;
        RECT 144.875 166.750 145.195 167.070 ;
        RECT 148.470 166.750 148.790 167.070 ;
        RECT 152.065 166.750 152.385 167.070 ;
        RECT 155.660 166.750 155.980 167.070 ;
        RECT 159.255 166.750 159.575 167.070 ;
        RECT 162.850 166.750 163.170 167.070 ;
        RECT 166.445 166.750 166.765 167.070 ;
        RECT 134.090 166.350 134.410 166.670 ;
        RECT 137.685 166.350 138.005 166.670 ;
        RECT 141.280 166.350 141.600 166.670 ;
        RECT 144.875 166.350 145.195 166.670 ;
        RECT 148.470 166.350 148.790 166.670 ;
        RECT 152.065 166.350 152.385 166.670 ;
        RECT 155.660 166.350 155.980 166.670 ;
        RECT 159.255 166.350 159.575 166.670 ;
        RECT 162.850 166.350 163.170 166.670 ;
        RECT 166.445 166.350 166.765 166.670 ;
        RECT 134.090 165.950 134.410 166.270 ;
        RECT 137.685 165.950 138.005 166.270 ;
        RECT 141.280 165.950 141.600 166.270 ;
        RECT 144.875 165.950 145.195 166.270 ;
        RECT 148.470 165.950 148.790 166.270 ;
        RECT 152.065 165.950 152.385 166.270 ;
        RECT 155.660 165.950 155.980 166.270 ;
        RECT 159.255 165.950 159.575 166.270 ;
        RECT 162.850 165.950 163.170 166.270 ;
        RECT 166.445 165.950 166.765 166.270 ;
        RECT 134.090 165.550 134.410 165.870 ;
        RECT 137.685 165.550 138.005 165.870 ;
        RECT 141.280 165.550 141.600 165.870 ;
        RECT 144.875 165.550 145.195 165.870 ;
        RECT 148.470 165.550 148.790 165.870 ;
        RECT 152.065 165.550 152.385 165.870 ;
        RECT 155.660 165.550 155.980 165.870 ;
        RECT 159.255 165.550 159.575 165.870 ;
        RECT 162.850 165.550 163.170 165.870 ;
        RECT 166.445 165.550 166.765 165.870 ;
        RECT 134.090 164.450 134.410 164.770 ;
        RECT 137.685 164.450 138.005 164.770 ;
        RECT 141.280 164.450 141.600 164.770 ;
        RECT 144.875 164.450 145.195 164.770 ;
        RECT 148.470 164.450 148.790 164.770 ;
        RECT 152.065 164.450 152.385 164.770 ;
        RECT 155.660 164.450 155.980 164.770 ;
        RECT 159.255 164.450 159.575 164.770 ;
        RECT 162.850 164.450 163.170 164.770 ;
        RECT 166.445 164.450 166.765 164.770 ;
        RECT 134.090 164.050 134.410 164.370 ;
        RECT 137.685 164.050 138.005 164.370 ;
        RECT 141.280 164.050 141.600 164.370 ;
        RECT 144.875 164.050 145.195 164.370 ;
        RECT 148.470 164.050 148.790 164.370 ;
        RECT 152.065 164.050 152.385 164.370 ;
        RECT 155.660 164.050 155.980 164.370 ;
        RECT 159.255 164.050 159.575 164.370 ;
        RECT 162.850 164.050 163.170 164.370 ;
        RECT 166.445 164.050 166.765 164.370 ;
        RECT 134.090 163.650 134.410 163.970 ;
        RECT 137.685 163.650 138.005 163.970 ;
        RECT 141.280 163.650 141.600 163.970 ;
        RECT 144.875 163.650 145.195 163.970 ;
        RECT 148.470 163.650 148.790 163.970 ;
        RECT 152.065 163.650 152.385 163.970 ;
        RECT 155.660 163.650 155.980 163.970 ;
        RECT 159.255 163.650 159.575 163.970 ;
        RECT 162.850 163.650 163.170 163.970 ;
        RECT 166.445 163.650 166.765 163.970 ;
        RECT 134.090 163.250 134.410 163.570 ;
        RECT 137.685 163.250 138.005 163.570 ;
        RECT 141.280 163.250 141.600 163.570 ;
        RECT 144.875 163.250 145.195 163.570 ;
        RECT 148.470 163.250 148.790 163.570 ;
        RECT 152.065 163.250 152.385 163.570 ;
        RECT 155.660 163.250 155.980 163.570 ;
        RECT 159.255 163.250 159.575 163.570 ;
        RECT 162.850 163.250 163.170 163.570 ;
        RECT 166.445 163.250 166.765 163.570 ;
        RECT 134.090 162.850 134.410 163.170 ;
        RECT 137.685 162.850 138.005 163.170 ;
        RECT 141.280 162.850 141.600 163.170 ;
        RECT 144.875 162.850 145.195 163.170 ;
        RECT 148.470 162.850 148.790 163.170 ;
        RECT 152.065 162.850 152.385 163.170 ;
        RECT 155.660 162.850 155.980 163.170 ;
        RECT 159.255 162.850 159.575 163.170 ;
        RECT 162.850 162.850 163.170 163.170 ;
        RECT 166.445 162.850 166.765 163.170 ;
        RECT 134.090 162.450 134.410 162.770 ;
        RECT 137.685 162.450 138.005 162.770 ;
        RECT 141.280 162.450 141.600 162.770 ;
        RECT 144.875 162.450 145.195 162.770 ;
        RECT 148.470 162.450 148.790 162.770 ;
        RECT 152.065 162.450 152.385 162.770 ;
        RECT 155.660 162.450 155.980 162.770 ;
        RECT 159.255 162.450 159.575 162.770 ;
        RECT 162.850 162.450 163.170 162.770 ;
        RECT 166.445 162.450 166.765 162.770 ;
        RECT 134.090 162.050 134.410 162.370 ;
        RECT 137.685 162.050 138.005 162.370 ;
        RECT 141.280 162.050 141.600 162.370 ;
        RECT 144.875 162.050 145.195 162.370 ;
        RECT 148.470 162.050 148.790 162.370 ;
        RECT 152.065 162.050 152.385 162.370 ;
        RECT 155.660 162.050 155.980 162.370 ;
        RECT 159.255 162.050 159.575 162.370 ;
        RECT 162.850 162.050 163.170 162.370 ;
        RECT 166.445 162.050 166.765 162.370 ;
        RECT 171.330 167.950 171.650 168.270 ;
        RECT 174.925 167.950 175.245 168.270 ;
        RECT 178.520 167.950 178.840 168.270 ;
        RECT 182.115 167.950 182.435 168.270 ;
        RECT 185.710 167.950 186.030 168.270 ;
        RECT 189.305 167.950 189.625 168.270 ;
        RECT 192.900 167.950 193.220 168.270 ;
        RECT 196.495 167.950 196.815 168.270 ;
        RECT 200.090 167.950 200.410 168.270 ;
        RECT 203.685 167.950 204.005 168.270 ;
        RECT 171.330 167.550 171.650 167.870 ;
        RECT 174.925 167.550 175.245 167.870 ;
        RECT 178.520 167.550 178.840 167.870 ;
        RECT 182.115 167.550 182.435 167.870 ;
        RECT 185.710 167.550 186.030 167.870 ;
        RECT 189.305 167.550 189.625 167.870 ;
        RECT 192.900 167.550 193.220 167.870 ;
        RECT 196.495 167.550 196.815 167.870 ;
        RECT 200.090 167.550 200.410 167.870 ;
        RECT 203.685 167.550 204.005 167.870 ;
        RECT 171.330 167.150 171.650 167.470 ;
        RECT 174.925 167.150 175.245 167.470 ;
        RECT 178.520 167.150 178.840 167.470 ;
        RECT 182.115 167.150 182.435 167.470 ;
        RECT 185.710 167.150 186.030 167.470 ;
        RECT 189.305 167.150 189.625 167.470 ;
        RECT 192.900 167.150 193.220 167.470 ;
        RECT 196.495 167.150 196.815 167.470 ;
        RECT 200.090 167.150 200.410 167.470 ;
        RECT 203.685 167.150 204.005 167.470 ;
        RECT 171.330 166.750 171.650 167.070 ;
        RECT 174.925 166.750 175.245 167.070 ;
        RECT 178.520 166.750 178.840 167.070 ;
        RECT 182.115 166.750 182.435 167.070 ;
        RECT 185.710 166.750 186.030 167.070 ;
        RECT 189.305 166.750 189.625 167.070 ;
        RECT 192.900 166.750 193.220 167.070 ;
        RECT 196.495 166.750 196.815 167.070 ;
        RECT 200.090 166.750 200.410 167.070 ;
        RECT 203.685 166.750 204.005 167.070 ;
        RECT 171.330 166.350 171.650 166.670 ;
        RECT 174.925 166.350 175.245 166.670 ;
        RECT 178.520 166.350 178.840 166.670 ;
        RECT 182.115 166.350 182.435 166.670 ;
        RECT 185.710 166.350 186.030 166.670 ;
        RECT 189.305 166.350 189.625 166.670 ;
        RECT 192.900 166.350 193.220 166.670 ;
        RECT 196.495 166.350 196.815 166.670 ;
        RECT 200.090 166.350 200.410 166.670 ;
        RECT 203.685 166.350 204.005 166.670 ;
        RECT 171.330 165.950 171.650 166.270 ;
        RECT 174.925 165.950 175.245 166.270 ;
        RECT 178.520 165.950 178.840 166.270 ;
        RECT 182.115 165.950 182.435 166.270 ;
        RECT 185.710 165.950 186.030 166.270 ;
        RECT 189.305 165.950 189.625 166.270 ;
        RECT 192.900 165.950 193.220 166.270 ;
        RECT 196.495 165.950 196.815 166.270 ;
        RECT 200.090 165.950 200.410 166.270 ;
        RECT 203.685 165.950 204.005 166.270 ;
        RECT 171.330 165.550 171.650 165.870 ;
        RECT 174.925 165.550 175.245 165.870 ;
        RECT 178.520 165.550 178.840 165.870 ;
        RECT 182.115 165.550 182.435 165.870 ;
        RECT 185.710 165.550 186.030 165.870 ;
        RECT 189.305 165.550 189.625 165.870 ;
        RECT 192.900 165.550 193.220 165.870 ;
        RECT 196.495 165.550 196.815 165.870 ;
        RECT 200.090 165.550 200.410 165.870 ;
        RECT 203.685 165.550 204.005 165.870 ;
        RECT 171.330 164.450 171.650 164.770 ;
        RECT 174.925 164.450 175.245 164.770 ;
        RECT 178.520 164.450 178.840 164.770 ;
        RECT 182.115 164.450 182.435 164.770 ;
        RECT 185.710 164.450 186.030 164.770 ;
        RECT 189.305 164.450 189.625 164.770 ;
        RECT 192.900 164.450 193.220 164.770 ;
        RECT 196.495 164.450 196.815 164.770 ;
        RECT 200.090 164.450 200.410 164.770 ;
        RECT 203.685 164.450 204.005 164.770 ;
        RECT 171.330 164.050 171.650 164.370 ;
        RECT 174.925 164.050 175.245 164.370 ;
        RECT 178.520 164.050 178.840 164.370 ;
        RECT 182.115 164.050 182.435 164.370 ;
        RECT 185.710 164.050 186.030 164.370 ;
        RECT 189.305 164.050 189.625 164.370 ;
        RECT 192.900 164.050 193.220 164.370 ;
        RECT 196.495 164.050 196.815 164.370 ;
        RECT 200.090 164.050 200.410 164.370 ;
        RECT 203.685 164.050 204.005 164.370 ;
        RECT 171.330 163.650 171.650 163.970 ;
        RECT 174.925 163.650 175.245 163.970 ;
        RECT 178.520 163.650 178.840 163.970 ;
        RECT 182.115 163.650 182.435 163.970 ;
        RECT 185.710 163.650 186.030 163.970 ;
        RECT 189.305 163.650 189.625 163.970 ;
        RECT 192.900 163.650 193.220 163.970 ;
        RECT 196.495 163.650 196.815 163.970 ;
        RECT 200.090 163.650 200.410 163.970 ;
        RECT 203.685 163.650 204.005 163.970 ;
        RECT 171.330 163.250 171.650 163.570 ;
        RECT 174.925 163.250 175.245 163.570 ;
        RECT 178.520 163.250 178.840 163.570 ;
        RECT 182.115 163.250 182.435 163.570 ;
        RECT 185.710 163.250 186.030 163.570 ;
        RECT 189.305 163.250 189.625 163.570 ;
        RECT 192.900 163.250 193.220 163.570 ;
        RECT 196.495 163.250 196.815 163.570 ;
        RECT 200.090 163.250 200.410 163.570 ;
        RECT 203.685 163.250 204.005 163.570 ;
        RECT 171.330 162.850 171.650 163.170 ;
        RECT 174.925 162.850 175.245 163.170 ;
        RECT 178.520 162.850 178.840 163.170 ;
        RECT 182.115 162.850 182.435 163.170 ;
        RECT 185.710 162.850 186.030 163.170 ;
        RECT 189.305 162.850 189.625 163.170 ;
        RECT 192.900 162.850 193.220 163.170 ;
        RECT 196.495 162.850 196.815 163.170 ;
        RECT 200.090 162.850 200.410 163.170 ;
        RECT 203.685 162.850 204.005 163.170 ;
        RECT 171.330 162.450 171.650 162.770 ;
        RECT 174.925 162.450 175.245 162.770 ;
        RECT 178.520 162.450 178.840 162.770 ;
        RECT 182.115 162.450 182.435 162.770 ;
        RECT 185.710 162.450 186.030 162.770 ;
        RECT 189.305 162.450 189.625 162.770 ;
        RECT 192.900 162.450 193.220 162.770 ;
        RECT 196.495 162.450 196.815 162.770 ;
        RECT 200.090 162.450 200.410 162.770 ;
        RECT 203.685 162.450 204.005 162.770 ;
        RECT 171.330 162.050 171.650 162.370 ;
        RECT 174.925 162.050 175.245 162.370 ;
        RECT 178.520 162.050 178.840 162.370 ;
        RECT 182.115 162.050 182.435 162.370 ;
        RECT 185.710 162.050 186.030 162.370 ;
        RECT 189.305 162.050 189.625 162.370 ;
        RECT 192.900 162.050 193.220 162.370 ;
        RECT 196.495 162.050 196.815 162.370 ;
        RECT 200.090 162.050 200.410 162.370 ;
        RECT 203.685 162.050 204.005 162.370 ;
        RECT 16.860 150.600 17.180 150.920 ;
        RECT 17.260 150.600 17.580 150.920 ;
        RECT 17.660 150.600 17.980 150.920 ;
        RECT 18.060 150.600 18.380 150.920 ;
        RECT 18.460 150.600 18.780 150.920 ;
        RECT 18.860 150.600 19.180 150.920 ;
        RECT 19.260 150.600 19.580 150.920 ;
        RECT 19.660 150.600 19.980 150.920 ;
        RECT 20.060 150.600 20.380 150.920 ;
        RECT 20.460 150.600 20.780 150.920 ;
        RECT 20.860 150.600 21.180 150.920 ;
        RECT 21.260 150.600 21.580 150.920 ;
        RECT 21.660 150.600 21.980 150.920 ;
        RECT 22.060 150.600 22.380 150.920 ;
        RECT 22.460 150.600 22.780 150.920 ;
        RECT 22.860 150.600 23.180 150.920 ;
        RECT 23.260 150.600 23.580 150.920 ;
        RECT 23.660 150.600 23.980 150.920 ;
        RECT 24.060 150.600 24.380 150.920 ;
        RECT 24.460 150.600 24.780 150.920 ;
        RECT 167.050 150.570 167.370 150.890 ;
        RECT 267.400 150.600 267.720 150.920 ;
        RECT 267.800 150.600 268.120 150.920 ;
        RECT 268.200 150.600 268.520 150.920 ;
        RECT 268.600 150.600 268.920 150.920 ;
        RECT 269.000 150.600 269.320 150.920 ;
        RECT 269.400 150.600 269.720 150.920 ;
        RECT 269.800 150.600 270.120 150.920 ;
        RECT 270.200 150.600 270.520 150.920 ;
        RECT 270.600 150.600 270.920 150.920 ;
        RECT 271.000 150.600 271.320 150.920 ;
        RECT 271.400 150.600 271.720 150.920 ;
        RECT 271.800 150.600 272.120 150.920 ;
        RECT 272.200 150.600 272.520 150.920 ;
        RECT 272.600 150.600 272.920 150.920 ;
        RECT 273.000 150.600 273.320 150.920 ;
        RECT 273.400 150.600 273.720 150.920 ;
        RECT 273.800 150.600 274.120 150.920 ;
        RECT 274.200 150.600 274.520 150.920 ;
        RECT 274.600 150.600 274.920 150.920 ;
        RECT 275.000 150.600 275.320 150.920 ;
        RECT 152.710 149.150 153.030 149.470 ;
        RECT 156.305 149.150 156.625 149.470 ;
        RECT 159.900 149.150 160.220 149.470 ;
        RECT 163.495 149.150 163.815 149.470 ;
        RECT 167.090 149.150 167.410 149.470 ;
        RECT 170.685 149.150 171.005 149.470 ;
        RECT 174.280 149.150 174.600 149.470 ;
        RECT 177.875 149.150 178.195 149.470 ;
        RECT 181.470 149.150 181.790 149.470 ;
        RECT 185.065 149.150 185.385 149.470 ;
        RECT 152.710 148.750 153.030 149.070 ;
        RECT 156.305 148.750 156.625 149.070 ;
        RECT 159.900 148.750 160.220 149.070 ;
        RECT 163.495 148.750 163.815 149.070 ;
        RECT 167.090 148.750 167.410 149.070 ;
        RECT 170.685 148.750 171.005 149.070 ;
        RECT 174.280 148.750 174.600 149.070 ;
        RECT 177.875 148.750 178.195 149.070 ;
        RECT 181.470 148.750 181.790 149.070 ;
        RECT 185.065 148.750 185.385 149.070 ;
        RECT 152.710 148.350 153.030 148.670 ;
        RECT 156.305 148.350 156.625 148.670 ;
        RECT 159.900 148.350 160.220 148.670 ;
        RECT 163.495 148.350 163.815 148.670 ;
        RECT 167.090 148.350 167.410 148.670 ;
        RECT 170.685 148.350 171.005 148.670 ;
        RECT 174.280 148.350 174.600 148.670 ;
        RECT 177.875 148.350 178.195 148.670 ;
        RECT 181.470 148.350 181.790 148.670 ;
        RECT 185.065 148.350 185.385 148.670 ;
        RECT 152.710 147.950 153.030 148.270 ;
        RECT 156.305 147.950 156.625 148.270 ;
        RECT 159.900 147.950 160.220 148.270 ;
        RECT 163.495 147.950 163.815 148.270 ;
        RECT 167.090 147.950 167.410 148.270 ;
        RECT 170.685 147.950 171.005 148.270 ;
        RECT 174.280 147.950 174.600 148.270 ;
        RECT 177.875 147.950 178.195 148.270 ;
        RECT 181.470 147.950 181.790 148.270 ;
        RECT 185.065 147.950 185.385 148.270 ;
        RECT 152.710 147.550 153.030 147.870 ;
        RECT 156.305 147.550 156.625 147.870 ;
        RECT 159.900 147.550 160.220 147.870 ;
        RECT 163.495 147.550 163.815 147.870 ;
        RECT 167.090 147.550 167.410 147.870 ;
        RECT 170.685 147.550 171.005 147.870 ;
        RECT 174.280 147.550 174.600 147.870 ;
        RECT 177.875 147.550 178.195 147.870 ;
        RECT 181.470 147.550 181.790 147.870 ;
        RECT 185.065 147.550 185.385 147.870 ;
        RECT 152.710 147.150 153.030 147.470 ;
        RECT 156.305 147.150 156.625 147.470 ;
        RECT 159.900 147.150 160.220 147.470 ;
        RECT 163.495 147.150 163.815 147.470 ;
        RECT 167.090 147.150 167.410 147.470 ;
        RECT 170.685 147.150 171.005 147.470 ;
        RECT 174.280 147.150 174.600 147.470 ;
        RECT 177.875 147.150 178.195 147.470 ;
        RECT 181.470 147.150 181.790 147.470 ;
        RECT 185.065 147.150 185.385 147.470 ;
        RECT 152.710 146.750 153.030 147.070 ;
        RECT 156.305 146.750 156.625 147.070 ;
        RECT 159.900 146.750 160.220 147.070 ;
        RECT 163.495 146.750 163.815 147.070 ;
        RECT 167.090 146.750 167.410 147.070 ;
        RECT 170.685 146.750 171.005 147.070 ;
        RECT 174.280 146.750 174.600 147.070 ;
        RECT 177.875 146.750 178.195 147.070 ;
        RECT 181.470 146.750 181.790 147.070 ;
        RECT 185.065 146.750 185.385 147.070 ;
        RECT 152.710 145.650 153.030 145.970 ;
        RECT 156.305 145.650 156.625 145.970 ;
        RECT 159.900 145.650 160.220 145.970 ;
        RECT 163.495 145.650 163.815 145.970 ;
        RECT 167.090 145.650 167.410 145.970 ;
        RECT 170.685 145.650 171.005 145.970 ;
        RECT 174.280 145.650 174.600 145.970 ;
        RECT 177.875 145.650 178.195 145.970 ;
        RECT 181.470 145.650 181.790 145.970 ;
        RECT 185.065 145.650 185.385 145.970 ;
        RECT 152.710 145.250 153.030 145.570 ;
        RECT 156.305 145.250 156.625 145.570 ;
        RECT 159.900 145.250 160.220 145.570 ;
        RECT 163.495 145.250 163.815 145.570 ;
        RECT 167.090 145.250 167.410 145.570 ;
        RECT 170.685 145.250 171.005 145.570 ;
        RECT 174.280 145.250 174.600 145.570 ;
        RECT 177.875 145.250 178.195 145.570 ;
        RECT 181.470 145.250 181.790 145.570 ;
        RECT 185.065 145.250 185.385 145.570 ;
        RECT 152.710 144.850 153.030 145.170 ;
        RECT 156.305 144.850 156.625 145.170 ;
        RECT 159.900 144.850 160.220 145.170 ;
        RECT 163.495 144.850 163.815 145.170 ;
        RECT 167.090 144.850 167.410 145.170 ;
        RECT 170.685 144.850 171.005 145.170 ;
        RECT 174.280 144.850 174.600 145.170 ;
        RECT 177.875 144.850 178.195 145.170 ;
        RECT 181.470 144.850 181.790 145.170 ;
        RECT 185.065 144.850 185.385 145.170 ;
        RECT 152.710 144.450 153.030 144.770 ;
        RECT 156.305 144.450 156.625 144.770 ;
        RECT 159.900 144.450 160.220 144.770 ;
        RECT 163.495 144.450 163.815 144.770 ;
        RECT 167.090 144.450 167.410 144.770 ;
        RECT 170.685 144.450 171.005 144.770 ;
        RECT 174.280 144.450 174.600 144.770 ;
        RECT 177.875 144.450 178.195 144.770 ;
        RECT 181.470 144.450 181.790 144.770 ;
        RECT 185.065 144.450 185.385 144.770 ;
        RECT 152.710 144.050 153.030 144.370 ;
        RECT 156.305 144.050 156.625 144.370 ;
        RECT 159.900 144.050 160.220 144.370 ;
        RECT 163.495 144.050 163.815 144.370 ;
        RECT 167.090 144.050 167.410 144.370 ;
        RECT 170.685 144.050 171.005 144.370 ;
        RECT 174.280 144.050 174.600 144.370 ;
        RECT 177.875 144.050 178.195 144.370 ;
        RECT 181.470 144.050 181.790 144.370 ;
        RECT 185.065 144.050 185.385 144.370 ;
        RECT 152.710 143.650 153.030 143.970 ;
        RECT 156.305 143.650 156.625 143.970 ;
        RECT 159.900 143.650 160.220 143.970 ;
        RECT 163.495 143.650 163.815 143.970 ;
        RECT 167.090 143.650 167.410 143.970 ;
        RECT 170.685 143.650 171.005 143.970 ;
        RECT 174.280 143.650 174.600 143.970 ;
        RECT 177.875 143.650 178.195 143.970 ;
        RECT 181.470 143.650 181.790 143.970 ;
        RECT 185.065 143.650 185.385 143.970 ;
        RECT 152.710 143.250 153.030 143.570 ;
        RECT 156.305 143.250 156.625 143.570 ;
        RECT 159.900 143.250 160.220 143.570 ;
        RECT 163.495 143.250 163.815 143.570 ;
        RECT 167.090 143.250 167.410 143.570 ;
        RECT 170.685 143.250 171.005 143.570 ;
        RECT 174.280 143.250 174.600 143.570 ;
        RECT 177.875 143.250 178.195 143.570 ;
        RECT 181.470 143.250 181.790 143.570 ;
        RECT 185.065 143.250 185.385 143.570 ;
        RECT 16.860 131.800 17.180 132.120 ;
        RECT 17.260 131.800 17.580 132.120 ;
        RECT 17.660 131.800 17.980 132.120 ;
        RECT 18.060 131.800 18.380 132.120 ;
        RECT 18.460 131.800 18.780 132.120 ;
        RECT 18.860 131.800 19.180 132.120 ;
        RECT 19.260 131.800 19.580 132.120 ;
        RECT 19.660 131.800 19.980 132.120 ;
        RECT 20.060 131.800 20.380 132.120 ;
        RECT 20.460 131.800 20.780 132.120 ;
        RECT 20.860 131.800 21.180 132.120 ;
        RECT 21.260 131.800 21.580 132.120 ;
        RECT 21.660 131.800 21.980 132.120 ;
        RECT 22.060 131.800 22.380 132.120 ;
        RECT 22.460 131.800 22.780 132.120 ;
        RECT 22.860 131.800 23.180 132.120 ;
        RECT 23.260 131.800 23.580 132.120 ;
        RECT 23.660 131.800 23.980 132.120 ;
        RECT 24.060 131.800 24.380 132.120 ;
        RECT 24.460 131.800 24.780 132.120 ;
        RECT 167.050 131.660 167.370 131.980 ;
        RECT 267.400 131.800 267.720 132.120 ;
        RECT 267.800 131.800 268.120 132.120 ;
        RECT 268.200 131.800 268.520 132.120 ;
        RECT 268.600 131.800 268.920 132.120 ;
        RECT 269.000 131.800 269.320 132.120 ;
        RECT 269.400 131.800 269.720 132.120 ;
        RECT 269.800 131.800 270.120 132.120 ;
        RECT 270.200 131.800 270.520 132.120 ;
        RECT 270.600 131.800 270.920 132.120 ;
        RECT 271.000 131.800 271.320 132.120 ;
        RECT 271.400 131.800 271.720 132.120 ;
        RECT 271.800 131.800 272.120 132.120 ;
        RECT 272.200 131.800 272.520 132.120 ;
        RECT 272.600 131.800 272.920 132.120 ;
        RECT 273.000 131.800 273.320 132.120 ;
        RECT 273.400 131.800 273.720 132.120 ;
        RECT 273.800 131.800 274.120 132.120 ;
        RECT 274.200 131.800 274.520 132.120 ;
        RECT 274.600 131.800 274.920 132.120 ;
        RECT 275.000 131.800 275.320 132.120 ;
        RECT 152.710 130.350 153.030 130.670 ;
        RECT 156.305 130.350 156.625 130.670 ;
        RECT 159.900 130.350 160.220 130.670 ;
        RECT 163.495 130.350 163.815 130.670 ;
        RECT 167.090 130.350 167.410 130.670 ;
        RECT 170.685 130.350 171.005 130.670 ;
        RECT 174.280 130.350 174.600 130.670 ;
        RECT 177.875 130.350 178.195 130.670 ;
        RECT 181.470 130.350 181.790 130.670 ;
        RECT 185.065 130.350 185.385 130.670 ;
        RECT 152.710 129.950 153.030 130.270 ;
        RECT 156.305 129.950 156.625 130.270 ;
        RECT 159.900 129.950 160.220 130.270 ;
        RECT 163.495 129.950 163.815 130.270 ;
        RECT 167.090 129.950 167.410 130.270 ;
        RECT 170.685 129.950 171.005 130.270 ;
        RECT 174.280 129.950 174.600 130.270 ;
        RECT 177.875 129.950 178.195 130.270 ;
        RECT 181.470 129.950 181.790 130.270 ;
        RECT 185.065 129.950 185.385 130.270 ;
        RECT 152.710 129.550 153.030 129.870 ;
        RECT 156.305 129.550 156.625 129.870 ;
        RECT 159.900 129.550 160.220 129.870 ;
        RECT 163.495 129.550 163.815 129.870 ;
        RECT 167.090 129.550 167.410 129.870 ;
        RECT 170.685 129.550 171.005 129.870 ;
        RECT 174.280 129.550 174.600 129.870 ;
        RECT 177.875 129.550 178.195 129.870 ;
        RECT 181.470 129.550 181.790 129.870 ;
        RECT 185.065 129.550 185.385 129.870 ;
        RECT 152.710 129.150 153.030 129.470 ;
        RECT 156.305 129.150 156.625 129.470 ;
        RECT 159.900 129.150 160.220 129.470 ;
        RECT 163.495 129.150 163.815 129.470 ;
        RECT 167.090 129.150 167.410 129.470 ;
        RECT 170.685 129.150 171.005 129.470 ;
        RECT 174.280 129.150 174.600 129.470 ;
        RECT 177.875 129.150 178.195 129.470 ;
        RECT 181.470 129.150 181.790 129.470 ;
        RECT 185.065 129.150 185.385 129.470 ;
        RECT 152.710 128.750 153.030 129.070 ;
        RECT 156.305 128.750 156.625 129.070 ;
        RECT 159.900 128.750 160.220 129.070 ;
        RECT 163.495 128.750 163.815 129.070 ;
        RECT 167.090 128.750 167.410 129.070 ;
        RECT 170.685 128.750 171.005 129.070 ;
        RECT 174.280 128.750 174.600 129.070 ;
        RECT 177.875 128.750 178.195 129.070 ;
        RECT 181.470 128.750 181.790 129.070 ;
        RECT 185.065 128.750 185.385 129.070 ;
        RECT 152.710 128.350 153.030 128.670 ;
        RECT 156.305 128.350 156.625 128.670 ;
        RECT 159.900 128.350 160.220 128.670 ;
        RECT 163.495 128.350 163.815 128.670 ;
        RECT 167.090 128.350 167.410 128.670 ;
        RECT 170.685 128.350 171.005 128.670 ;
        RECT 174.280 128.350 174.600 128.670 ;
        RECT 177.875 128.350 178.195 128.670 ;
        RECT 181.470 128.350 181.790 128.670 ;
        RECT 185.065 128.350 185.385 128.670 ;
        RECT 152.710 127.950 153.030 128.270 ;
        RECT 156.305 127.950 156.625 128.270 ;
        RECT 159.900 127.950 160.220 128.270 ;
        RECT 163.495 127.950 163.815 128.270 ;
        RECT 167.090 127.950 167.410 128.270 ;
        RECT 170.685 127.950 171.005 128.270 ;
        RECT 174.280 127.950 174.600 128.270 ;
        RECT 177.875 127.950 178.195 128.270 ;
        RECT 181.470 127.950 181.790 128.270 ;
        RECT 185.065 127.950 185.385 128.270 ;
        RECT 152.710 126.850 153.030 127.170 ;
        RECT 156.305 126.850 156.625 127.170 ;
        RECT 159.900 126.850 160.220 127.170 ;
        RECT 163.495 126.850 163.815 127.170 ;
        RECT 167.090 126.850 167.410 127.170 ;
        RECT 170.685 126.850 171.005 127.170 ;
        RECT 174.280 126.850 174.600 127.170 ;
        RECT 177.875 126.850 178.195 127.170 ;
        RECT 181.470 126.850 181.790 127.170 ;
        RECT 185.065 126.850 185.385 127.170 ;
        RECT 152.710 126.450 153.030 126.770 ;
        RECT 156.305 126.450 156.625 126.770 ;
        RECT 159.900 126.450 160.220 126.770 ;
        RECT 163.495 126.450 163.815 126.770 ;
        RECT 167.090 126.450 167.410 126.770 ;
        RECT 170.685 126.450 171.005 126.770 ;
        RECT 174.280 126.450 174.600 126.770 ;
        RECT 177.875 126.450 178.195 126.770 ;
        RECT 181.470 126.450 181.790 126.770 ;
        RECT 185.065 126.450 185.385 126.770 ;
        RECT 152.710 126.050 153.030 126.370 ;
        RECT 156.305 126.050 156.625 126.370 ;
        RECT 159.900 126.050 160.220 126.370 ;
        RECT 163.495 126.050 163.815 126.370 ;
        RECT 167.090 126.050 167.410 126.370 ;
        RECT 170.685 126.050 171.005 126.370 ;
        RECT 174.280 126.050 174.600 126.370 ;
        RECT 177.875 126.050 178.195 126.370 ;
        RECT 181.470 126.050 181.790 126.370 ;
        RECT 185.065 126.050 185.385 126.370 ;
        RECT 152.710 125.650 153.030 125.970 ;
        RECT 156.305 125.650 156.625 125.970 ;
        RECT 159.900 125.650 160.220 125.970 ;
        RECT 163.495 125.650 163.815 125.970 ;
        RECT 167.090 125.650 167.410 125.970 ;
        RECT 170.685 125.650 171.005 125.970 ;
        RECT 174.280 125.650 174.600 125.970 ;
        RECT 177.875 125.650 178.195 125.970 ;
        RECT 181.470 125.650 181.790 125.970 ;
        RECT 185.065 125.650 185.385 125.970 ;
        RECT 152.710 125.250 153.030 125.570 ;
        RECT 156.305 125.250 156.625 125.570 ;
        RECT 159.900 125.250 160.220 125.570 ;
        RECT 163.495 125.250 163.815 125.570 ;
        RECT 167.090 125.250 167.410 125.570 ;
        RECT 170.685 125.250 171.005 125.570 ;
        RECT 174.280 125.250 174.600 125.570 ;
        RECT 177.875 125.250 178.195 125.570 ;
        RECT 181.470 125.250 181.790 125.570 ;
        RECT 185.065 125.250 185.385 125.570 ;
        RECT 152.710 124.850 153.030 125.170 ;
        RECT 156.305 124.850 156.625 125.170 ;
        RECT 159.900 124.850 160.220 125.170 ;
        RECT 163.495 124.850 163.815 125.170 ;
        RECT 167.090 124.850 167.410 125.170 ;
        RECT 170.685 124.850 171.005 125.170 ;
        RECT 174.280 124.850 174.600 125.170 ;
        RECT 177.875 124.850 178.195 125.170 ;
        RECT 181.470 124.850 181.790 125.170 ;
        RECT 185.065 124.850 185.385 125.170 ;
        RECT 152.710 124.450 153.030 124.770 ;
        RECT 156.305 124.450 156.625 124.770 ;
        RECT 159.900 124.450 160.220 124.770 ;
        RECT 163.495 124.450 163.815 124.770 ;
        RECT 167.090 124.450 167.410 124.770 ;
        RECT 170.685 124.450 171.005 124.770 ;
        RECT 174.280 124.450 174.600 124.770 ;
        RECT 177.875 124.450 178.195 124.770 ;
        RECT 181.470 124.450 181.790 124.770 ;
        RECT 185.065 124.450 185.385 124.770 ;
        RECT 16.860 113.000 17.180 113.320 ;
        RECT 17.260 113.000 17.580 113.320 ;
        RECT 17.660 113.000 17.980 113.320 ;
        RECT 18.060 113.000 18.380 113.320 ;
        RECT 18.460 113.000 18.780 113.320 ;
        RECT 18.860 113.000 19.180 113.320 ;
        RECT 19.260 113.000 19.580 113.320 ;
        RECT 19.660 113.000 19.980 113.320 ;
        RECT 20.060 113.000 20.380 113.320 ;
        RECT 20.460 113.000 20.780 113.320 ;
        RECT 20.860 113.000 21.180 113.320 ;
        RECT 21.260 113.000 21.580 113.320 ;
        RECT 21.660 113.000 21.980 113.320 ;
        RECT 22.060 113.000 22.380 113.320 ;
        RECT 22.460 113.000 22.780 113.320 ;
        RECT 22.860 113.000 23.180 113.320 ;
        RECT 23.260 113.000 23.580 113.320 ;
        RECT 23.660 113.000 23.980 113.320 ;
        RECT 24.060 113.000 24.380 113.320 ;
        RECT 24.460 113.000 24.780 113.320 ;
        RECT 267.400 113.000 267.720 113.320 ;
        RECT 267.800 113.000 268.120 113.320 ;
        RECT 268.200 113.000 268.520 113.320 ;
        RECT 268.600 113.000 268.920 113.320 ;
        RECT 269.000 113.000 269.320 113.320 ;
        RECT 269.400 113.000 269.720 113.320 ;
        RECT 269.800 113.000 270.120 113.320 ;
        RECT 270.200 113.000 270.520 113.320 ;
        RECT 270.600 113.000 270.920 113.320 ;
        RECT 271.000 113.000 271.320 113.320 ;
        RECT 271.400 113.000 271.720 113.320 ;
        RECT 271.800 113.000 272.120 113.320 ;
        RECT 272.200 113.000 272.520 113.320 ;
        RECT 272.600 113.000 272.920 113.320 ;
        RECT 273.000 113.000 273.320 113.320 ;
        RECT 273.400 113.000 273.720 113.320 ;
        RECT 273.800 113.000 274.120 113.320 ;
        RECT 274.200 113.000 274.520 113.320 ;
        RECT 274.600 113.000 274.920 113.320 ;
        RECT 275.000 113.000 275.320 113.320 ;
        RECT 16.860 94.200 17.180 94.520 ;
        RECT 17.260 94.200 17.580 94.520 ;
        RECT 17.660 94.200 17.980 94.520 ;
        RECT 18.060 94.200 18.380 94.520 ;
        RECT 18.460 94.200 18.780 94.520 ;
        RECT 18.860 94.200 19.180 94.520 ;
        RECT 19.260 94.200 19.580 94.520 ;
        RECT 19.660 94.200 19.980 94.520 ;
        RECT 20.060 94.200 20.380 94.520 ;
        RECT 20.460 94.200 20.780 94.520 ;
        RECT 20.860 94.200 21.180 94.520 ;
        RECT 21.260 94.200 21.580 94.520 ;
        RECT 21.660 94.200 21.980 94.520 ;
        RECT 22.060 94.200 22.380 94.520 ;
        RECT 22.460 94.200 22.780 94.520 ;
        RECT 22.860 94.200 23.180 94.520 ;
        RECT 23.260 94.200 23.580 94.520 ;
        RECT 23.660 94.200 23.980 94.520 ;
        RECT 24.060 94.200 24.380 94.520 ;
        RECT 24.460 94.200 24.780 94.520 ;
        RECT 267.400 94.200 267.720 94.520 ;
        RECT 267.800 94.200 268.120 94.520 ;
        RECT 268.200 94.200 268.520 94.520 ;
        RECT 268.600 94.200 268.920 94.520 ;
        RECT 269.000 94.200 269.320 94.520 ;
        RECT 269.400 94.200 269.720 94.520 ;
        RECT 269.800 94.200 270.120 94.520 ;
        RECT 270.200 94.200 270.520 94.520 ;
        RECT 270.600 94.200 270.920 94.520 ;
        RECT 271.000 94.200 271.320 94.520 ;
        RECT 271.400 94.200 271.720 94.520 ;
        RECT 271.800 94.200 272.120 94.520 ;
        RECT 272.200 94.200 272.520 94.520 ;
        RECT 272.600 94.200 272.920 94.520 ;
        RECT 273.000 94.200 273.320 94.520 ;
        RECT 273.400 94.200 273.720 94.520 ;
        RECT 273.800 94.200 274.120 94.520 ;
        RECT 274.200 94.200 274.520 94.520 ;
        RECT 274.600 94.200 274.920 94.520 ;
        RECT 275.000 94.200 275.320 94.520 ;
        RECT 16.860 75.400 17.180 75.720 ;
        RECT 17.260 75.400 17.580 75.720 ;
        RECT 17.660 75.400 17.980 75.720 ;
        RECT 18.060 75.400 18.380 75.720 ;
        RECT 18.460 75.400 18.780 75.720 ;
        RECT 18.860 75.400 19.180 75.720 ;
        RECT 19.260 75.400 19.580 75.720 ;
        RECT 19.660 75.400 19.980 75.720 ;
        RECT 20.060 75.400 20.380 75.720 ;
        RECT 20.460 75.400 20.780 75.720 ;
        RECT 20.860 75.400 21.180 75.720 ;
        RECT 21.260 75.400 21.580 75.720 ;
        RECT 21.660 75.400 21.980 75.720 ;
        RECT 22.060 75.400 22.380 75.720 ;
        RECT 22.460 75.400 22.780 75.720 ;
        RECT 22.860 75.400 23.180 75.720 ;
        RECT 23.260 75.400 23.580 75.720 ;
        RECT 23.660 75.400 23.980 75.720 ;
        RECT 24.060 75.400 24.380 75.720 ;
        RECT 24.460 75.400 24.780 75.720 ;
        RECT 267.400 75.400 267.720 75.720 ;
        RECT 267.800 75.400 268.120 75.720 ;
        RECT 268.200 75.400 268.520 75.720 ;
        RECT 268.600 75.400 268.920 75.720 ;
        RECT 269.000 75.400 269.320 75.720 ;
        RECT 269.400 75.400 269.720 75.720 ;
        RECT 269.800 75.400 270.120 75.720 ;
        RECT 270.200 75.400 270.520 75.720 ;
        RECT 270.600 75.400 270.920 75.720 ;
        RECT 271.000 75.400 271.320 75.720 ;
        RECT 271.400 75.400 271.720 75.720 ;
        RECT 271.800 75.400 272.120 75.720 ;
        RECT 272.200 75.400 272.520 75.720 ;
        RECT 272.600 75.400 272.920 75.720 ;
        RECT 273.000 75.400 273.320 75.720 ;
        RECT 273.400 75.400 273.720 75.720 ;
        RECT 273.800 75.400 274.120 75.720 ;
        RECT 274.200 75.400 274.520 75.720 ;
        RECT 274.600 75.400 274.920 75.720 ;
        RECT 275.000 75.400 275.320 75.720 ;
        RECT 16.860 56.600 17.180 56.920 ;
        RECT 17.260 56.600 17.580 56.920 ;
        RECT 17.660 56.600 17.980 56.920 ;
        RECT 18.060 56.600 18.380 56.920 ;
        RECT 18.460 56.600 18.780 56.920 ;
        RECT 18.860 56.600 19.180 56.920 ;
        RECT 19.260 56.600 19.580 56.920 ;
        RECT 19.660 56.600 19.980 56.920 ;
        RECT 20.060 56.600 20.380 56.920 ;
        RECT 20.460 56.600 20.780 56.920 ;
        RECT 20.860 56.600 21.180 56.920 ;
        RECT 21.260 56.600 21.580 56.920 ;
        RECT 21.660 56.600 21.980 56.920 ;
        RECT 22.060 56.600 22.380 56.920 ;
        RECT 22.460 56.600 22.780 56.920 ;
        RECT 22.860 56.600 23.180 56.920 ;
        RECT 23.260 56.600 23.580 56.920 ;
        RECT 23.660 56.600 23.980 56.920 ;
        RECT 24.060 56.600 24.380 56.920 ;
        RECT 24.460 56.600 24.780 56.920 ;
        RECT 267.400 56.600 267.720 56.920 ;
        RECT 267.800 56.600 268.120 56.920 ;
        RECT 268.200 56.600 268.520 56.920 ;
        RECT 268.600 56.600 268.920 56.920 ;
        RECT 269.000 56.600 269.320 56.920 ;
        RECT 269.400 56.600 269.720 56.920 ;
        RECT 269.800 56.600 270.120 56.920 ;
        RECT 270.200 56.600 270.520 56.920 ;
        RECT 270.600 56.600 270.920 56.920 ;
        RECT 271.000 56.600 271.320 56.920 ;
        RECT 271.400 56.600 271.720 56.920 ;
        RECT 271.800 56.600 272.120 56.920 ;
        RECT 272.200 56.600 272.520 56.920 ;
        RECT 272.600 56.600 272.920 56.920 ;
        RECT 273.000 56.600 273.320 56.920 ;
        RECT 273.400 56.600 273.720 56.920 ;
        RECT 273.800 56.600 274.120 56.920 ;
        RECT 274.200 56.600 274.520 56.920 ;
        RECT 274.600 56.600 274.920 56.920 ;
        RECT 275.000 56.600 275.320 56.920 ;
        RECT 16.860 37.800 17.180 38.120 ;
        RECT 17.260 37.800 17.580 38.120 ;
        RECT 17.660 37.800 17.980 38.120 ;
        RECT 18.060 37.800 18.380 38.120 ;
        RECT 18.460 37.800 18.780 38.120 ;
        RECT 18.860 37.800 19.180 38.120 ;
        RECT 19.260 37.800 19.580 38.120 ;
        RECT 19.660 37.800 19.980 38.120 ;
        RECT 20.060 37.800 20.380 38.120 ;
        RECT 20.460 37.800 20.780 38.120 ;
        RECT 20.860 37.800 21.180 38.120 ;
        RECT 21.260 37.800 21.580 38.120 ;
        RECT 21.660 37.800 21.980 38.120 ;
        RECT 22.060 37.800 22.380 38.120 ;
        RECT 22.460 37.800 22.780 38.120 ;
        RECT 22.860 37.800 23.180 38.120 ;
        RECT 23.260 37.800 23.580 38.120 ;
        RECT 23.660 37.800 23.980 38.120 ;
        RECT 24.060 37.800 24.380 38.120 ;
        RECT 24.460 37.800 24.780 38.120 ;
        RECT 267.400 37.800 267.720 38.120 ;
        RECT 267.800 37.800 268.120 38.120 ;
        RECT 268.200 37.800 268.520 38.120 ;
        RECT 268.600 37.800 268.920 38.120 ;
        RECT 269.000 37.800 269.320 38.120 ;
        RECT 269.400 37.800 269.720 38.120 ;
        RECT 269.800 37.800 270.120 38.120 ;
        RECT 270.200 37.800 270.520 38.120 ;
        RECT 270.600 37.800 270.920 38.120 ;
        RECT 271.000 37.800 271.320 38.120 ;
        RECT 271.400 37.800 271.720 38.120 ;
        RECT 271.800 37.800 272.120 38.120 ;
        RECT 272.200 37.800 272.520 38.120 ;
        RECT 272.600 37.800 272.920 38.120 ;
        RECT 273.000 37.800 273.320 38.120 ;
        RECT 273.400 37.800 273.720 38.120 ;
        RECT 273.800 37.800 274.120 38.120 ;
        RECT 274.200 37.800 274.520 38.120 ;
        RECT 274.600 37.800 274.920 38.120 ;
        RECT 275.000 37.800 275.320 38.120 ;
      LAYER met4 ;
        RECT 16.740 0.000 24.900 282.880 ;
        RECT 167.045 187.775 167.375 188.105 ;
        RECT 167.060 187.150 167.360 187.775 ;
        RECT 152.630 184.270 153.110 187.150 ;
        RECT 156.225 184.270 156.705 187.150 ;
        RECT 159.820 184.270 160.300 187.150 ;
        RECT 163.415 184.270 163.895 187.150 ;
        RECT 167.010 184.270 167.490 187.150 ;
        RECT 170.605 184.270 171.085 187.150 ;
        RECT 174.200 184.270 174.680 187.150 ;
        RECT 177.795 184.270 178.275 187.150 ;
        RECT 181.390 184.270 181.870 187.150 ;
        RECT 184.985 184.270 185.465 187.150 ;
        RECT 152.630 180.770 153.110 183.650 ;
        RECT 156.225 180.770 156.705 183.650 ;
        RECT 159.820 180.770 160.300 183.650 ;
        RECT 163.415 180.770 163.895 183.650 ;
        RECT 167.010 180.770 167.490 183.650 ;
        RECT 170.605 180.770 171.085 183.650 ;
        RECT 174.200 180.770 174.680 183.650 ;
        RECT 177.795 180.770 178.275 183.650 ;
        RECT 181.390 180.770 181.870 183.650 ;
        RECT 184.985 180.770 185.465 183.650 ;
        RECT 166.355 168.865 166.685 169.195 ;
        RECT 170.495 169.180 170.825 169.195 ;
        RECT 170.495 168.880 171.670 169.180 ;
        RECT 170.495 168.865 170.825 168.880 ;
        RECT 166.370 168.350 166.670 168.865 ;
        RECT 171.370 168.350 171.670 168.880 ;
        RECT 134.010 165.470 134.490 168.350 ;
        RECT 137.605 165.470 138.085 168.350 ;
        RECT 141.200 165.470 141.680 168.350 ;
        RECT 144.795 165.470 145.275 168.350 ;
        RECT 148.390 165.470 148.870 168.350 ;
        RECT 151.985 165.470 152.465 168.350 ;
        RECT 155.580 165.470 156.060 168.350 ;
        RECT 159.175 165.470 159.655 168.350 ;
        RECT 162.770 165.470 163.250 168.350 ;
        RECT 166.365 165.470 166.845 168.350 ;
        RECT 171.250 165.470 171.730 168.350 ;
        RECT 174.845 165.470 175.325 168.350 ;
        RECT 178.440 165.470 178.920 168.350 ;
        RECT 182.035 165.470 182.515 168.350 ;
        RECT 185.630 165.470 186.110 168.350 ;
        RECT 189.225 165.470 189.705 168.350 ;
        RECT 192.820 165.470 193.300 168.350 ;
        RECT 196.415 165.470 196.895 168.350 ;
        RECT 200.010 165.470 200.490 168.350 ;
        RECT 203.605 165.470 204.085 168.350 ;
        RECT 134.010 161.970 134.490 164.850 ;
        RECT 137.605 161.970 138.085 164.850 ;
        RECT 141.200 161.970 141.680 164.850 ;
        RECT 144.795 161.970 145.275 164.850 ;
        RECT 148.390 161.970 148.870 164.850 ;
        RECT 151.985 161.970 152.465 164.850 ;
        RECT 155.580 161.970 156.060 164.850 ;
        RECT 159.175 161.970 159.655 164.850 ;
        RECT 162.770 161.970 163.250 164.850 ;
        RECT 166.365 161.970 166.845 164.850 ;
        RECT 171.250 161.970 171.730 164.850 ;
        RECT 174.845 161.970 175.325 164.850 ;
        RECT 178.440 161.970 178.920 164.850 ;
        RECT 182.035 161.970 182.515 164.850 ;
        RECT 185.630 161.970 186.110 164.850 ;
        RECT 189.225 161.970 189.705 164.850 ;
        RECT 192.820 161.970 193.300 164.850 ;
        RECT 196.415 161.970 196.895 164.850 ;
        RECT 200.010 161.970 200.490 164.850 ;
        RECT 203.605 161.970 204.085 164.850 ;
        RECT 167.045 150.565 167.375 150.895 ;
        RECT 167.060 149.550 167.360 150.565 ;
        RECT 152.630 146.670 153.110 149.550 ;
        RECT 156.225 146.670 156.705 149.550 ;
        RECT 159.820 146.670 160.300 149.550 ;
        RECT 163.415 146.670 163.895 149.550 ;
        RECT 167.010 146.670 167.490 149.550 ;
        RECT 170.605 146.670 171.085 149.550 ;
        RECT 174.200 146.670 174.680 149.550 ;
        RECT 177.795 146.670 178.275 149.550 ;
        RECT 181.390 146.670 181.870 149.550 ;
        RECT 184.985 146.670 185.465 149.550 ;
        RECT 152.630 143.170 153.110 146.050 ;
        RECT 156.225 143.170 156.705 146.050 ;
        RECT 159.820 143.170 160.300 146.050 ;
        RECT 163.415 143.170 163.895 146.050 ;
        RECT 167.010 143.170 167.490 146.050 ;
        RECT 170.605 143.170 171.085 146.050 ;
        RECT 174.200 143.170 174.680 146.050 ;
        RECT 177.795 143.170 178.275 146.050 ;
        RECT 181.390 143.170 181.870 146.050 ;
        RECT 184.985 143.170 185.465 146.050 ;
        RECT 167.045 131.655 167.375 131.985 ;
        RECT 167.060 130.750 167.360 131.655 ;
        RECT 152.630 127.870 153.110 130.750 ;
        RECT 156.225 127.870 156.705 130.750 ;
        RECT 159.820 127.870 160.300 130.750 ;
        RECT 163.415 127.870 163.895 130.750 ;
        RECT 167.010 127.870 167.490 130.750 ;
        RECT 170.605 127.870 171.085 130.750 ;
        RECT 174.200 127.870 174.680 130.750 ;
        RECT 177.795 127.870 178.275 130.750 ;
        RECT 181.390 127.870 181.870 130.750 ;
        RECT 184.985 127.870 185.465 130.750 ;
        RECT 152.630 124.370 153.110 127.250 ;
        RECT 156.225 124.370 156.705 127.250 ;
        RECT 159.820 124.370 160.300 127.250 ;
        RECT 163.415 124.370 163.895 127.250 ;
        RECT 167.010 124.370 167.490 127.250 ;
        RECT 170.605 124.370 171.085 127.250 ;
        RECT 174.200 124.370 174.680 127.250 ;
        RECT 177.795 124.370 178.275 127.250 ;
        RECT 181.390 124.370 181.870 127.250 ;
        RECT 184.985 124.370 185.465 127.250 ;
        RECT 267.280 0.000 275.440 282.880 ;
      LAYER via4 ;
        RECT 17.030 258.530 24.610 266.110 ;
        RECT 267.570 258.530 275.150 266.110 ;
        RECT 17.030 16.610 24.610 24.190 ;
        RECT 267.570 16.610 275.150 24.190 ;
      LAYER met5 ;
        RECT 0.000 258.240 292.560 266.400 ;
        RECT 0.000 16.320 292.560 24.480 ;
    END
  END VDD
  OBS
      LAYER pwell ;
        RECT 119.460 238.230 122.300 242.490 ;
        RECT 70.460 219.430 73.300 223.690 ;
        RECT 186.250 200.630 207.410 204.890 ;
        RECT 126.960 181.830 148.120 186.090 ;
        RECT 126.960 125.430 148.120 129.690 ;
      LAYER li1 ;
        RECT 104.160 240.735 106.320 243.585 ;
        RECT 104.160 235.935 106.320 238.785 ;
        RECT 114.200 235.935 116.360 243.585 ;
        RECT 119.650 238.630 119.820 242.380 ;
        RECT 119.645 238.340 119.820 238.630 ;
        RECT 119.645 237.510 119.815 238.340 ;
        RECT 119.590 237.210 122.170 237.510 ;
        RECT 119.990 236.080 122.170 236.380 ;
        RECT 147.345 236.180 147.515 236.215 ;
        RECT 120.205 236.045 120.375 236.080 ;
        RECT 124.150 235.880 262.190 236.180 ;
        RECT 70.650 219.830 70.820 223.580 ;
        RECT 70.645 219.540 70.820 219.830 ;
        RECT 70.645 218.710 70.815 219.540 ;
        RECT 216.415 219.525 219.885 222.995 ;
        RECT 223.115 219.525 226.585 222.995 ;
        RECT 229.815 219.525 233.285 222.995 ;
        RECT 236.515 219.525 239.985 222.995 ;
        RECT 243.215 219.525 246.685 222.995 ;
        RECT 249.915 219.525 253.385 222.995 ;
        RECT 256.615 219.525 260.085 222.995 ;
        RECT 70.590 218.410 73.170 218.710 ;
        RECT 71.905 218.365 72.075 218.410 ;
        RECT 70.990 217.280 73.170 217.580 ;
        RECT 75.150 217.080 213.190 217.380 ;
        RECT 186.380 206.210 207.280 206.510 ;
        RECT 146.925 199.110 147.095 206.005 ;
        RECT 151.505 199.110 151.675 206.005 ;
        RECT 156.085 199.110 156.255 206.005 ;
        RECT 160.665 199.110 160.835 206.005 ;
        RECT 165.245 199.110 165.415 206.005 ;
        RECT 169.825 199.110 169.995 206.005 ;
        RECT 174.405 199.110 174.575 206.005 ;
        RECT 188.725 204.780 188.895 206.210 ;
        RECT 193.305 204.780 193.475 206.210 ;
        RECT 197.885 204.780 198.055 206.210 ;
        RECT 202.465 204.780 202.635 206.210 ;
        RECT 207.045 204.780 207.215 206.210 ;
        RECT 186.440 201.030 186.610 204.780 ;
        RECT 188.725 204.690 188.900 204.780 ;
        RECT 186.435 200.740 186.610 201.030 ;
        RECT 188.730 200.740 188.900 204.690 ;
        RECT 191.020 201.030 191.190 204.780 ;
        RECT 193.305 204.690 193.480 204.780 ;
        RECT 191.015 200.740 191.190 201.030 ;
        RECT 193.310 200.740 193.480 204.690 ;
        RECT 195.600 201.030 195.770 204.780 ;
        RECT 197.885 204.690 198.060 204.780 ;
        RECT 195.595 200.740 195.770 201.030 ;
        RECT 197.890 200.740 198.060 204.690 ;
        RECT 200.180 201.030 200.350 204.780 ;
        RECT 202.465 204.690 202.640 204.780 ;
        RECT 200.175 200.740 200.350 201.030 ;
        RECT 202.470 200.740 202.640 204.690 ;
        RECT 204.760 201.030 204.930 204.780 ;
        RECT 207.045 204.690 207.220 204.780 ;
        RECT 204.755 200.740 204.930 201.030 ;
        RECT 207.050 200.740 207.220 204.690 ;
        RECT 186.435 200.410 186.605 200.740 ;
        RECT 191.015 200.410 191.185 200.740 ;
        RECT 195.595 200.410 195.765 200.740 ;
        RECT 200.175 200.410 200.345 200.740 ;
        RECT 204.755 200.410 204.925 200.740 ;
        RECT 210.535 200.725 214.005 204.195 ;
        RECT 217.235 200.725 220.705 204.195 ;
        RECT 223.935 200.725 227.405 204.195 ;
        RECT 230.635 200.725 234.105 204.195 ;
        RECT 237.335 200.725 240.805 204.195 ;
        RECT 244.035 200.725 247.505 204.195 ;
        RECT 250.735 200.725 254.205 204.195 ;
        RECT 257.435 200.725 260.905 204.195 ;
        RECT 186.380 200.110 207.280 200.410 ;
        RECT 146.690 198.810 174.810 199.110 ;
        RECT 146.690 198.280 174.810 198.580 ;
        RECT 127.090 187.410 147.990 187.710 ;
        RECT 68.390 184.335 70.550 187.185 ;
        RECT 68.390 179.535 70.550 182.385 ;
        RECT 78.430 179.535 80.590 187.185 ;
        RECT 82.110 184.335 84.270 187.185 ;
        RECT 82.110 179.535 84.270 182.385 ;
        RECT 92.150 179.535 94.310 187.185 ;
        RECT 95.835 184.335 97.995 187.185 ;
        RECT 108.745 179.535 110.905 187.185 ;
        RECT 112.490 184.335 114.650 187.185 ;
        RECT 112.490 179.535 114.650 182.385 ;
        RECT 122.530 179.535 124.690 187.185 ;
        RECT 129.435 185.980 129.605 187.410 ;
        RECT 134.015 185.980 134.185 187.410 ;
        RECT 138.595 185.980 138.765 187.410 ;
        RECT 143.175 185.980 143.345 187.410 ;
        RECT 147.755 185.980 147.925 187.410 ;
        RECT 127.150 182.230 127.320 185.980 ;
        RECT 129.435 185.890 129.610 185.980 ;
        RECT 127.145 181.940 127.320 182.230 ;
        RECT 129.440 181.940 129.610 185.890 ;
        RECT 131.730 182.230 131.900 185.980 ;
        RECT 134.015 185.890 134.190 185.980 ;
        RECT 131.725 181.940 131.900 182.230 ;
        RECT 134.020 181.940 134.190 185.890 ;
        RECT 136.310 182.230 136.480 185.980 ;
        RECT 138.595 185.890 138.770 185.980 ;
        RECT 136.305 181.940 136.480 182.230 ;
        RECT 138.600 181.940 138.770 185.890 ;
        RECT 140.890 182.230 141.060 185.980 ;
        RECT 143.175 185.890 143.350 185.980 ;
        RECT 140.885 181.940 141.060 182.230 ;
        RECT 143.180 181.940 143.350 185.890 ;
        RECT 145.470 182.230 145.640 185.980 ;
        RECT 147.755 185.890 147.930 185.980 ;
        RECT 145.465 181.940 145.640 182.230 ;
        RECT 147.760 181.940 147.930 185.890 ;
        RECT 127.145 181.610 127.315 181.940 ;
        RECT 131.725 181.610 131.895 181.940 ;
        RECT 136.305 181.610 136.475 181.940 ;
        RECT 140.885 181.610 141.055 181.940 ;
        RECT 145.465 181.610 145.635 181.940 ;
        RECT 127.090 181.310 147.990 181.610 ;
        RECT 187.595 180.310 187.765 187.205 ;
        RECT 192.175 180.310 192.345 187.205 ;
        RECT 196.755 180.310 196.925 187.205 ;
        RECT 201.335 180.310 201.505 187.205 ;
        RECT 210.535 181.925 214.005 185.395 ;
        RECT 217.235 181.925 220.705 185.395 ;
        RECT 223.935 181.925 227.405 185.395 ;
        RECT 230.635 181.925 234.105 185.395 ;
        RECT 237.335 181.925 240.805 185.395 ;
        RECT 244.035 181.925 247.505 185.395 ;
        RECT 250.735 181.925 254.205 185.395 ;
        RECT 257.435 181.925 260.905 185.395 ;
        RECT 187.360 180.010 201.740 180.310 ;
        RECT 187.360 179.480 201.740 179.780 ;
        RECT 96.320 165.535 98.480 168.385 ;
        RECT 96.320 160.735 98.480 163.585 ;
        RECT 106.360 160.735 108.520 168.385 ;
        RECT 110.045 165.535 112.205 168.385 ;
        RECT 122.955 160.735 125.115 168.385 ;
        RECT 210.535 163.125 214.005 166.595 ;
        RECT 217.235 163.125 220.705 166.595 ;
        RECT 223.935 163.125 227.405 166.595 ;
        RECT 230.635 163.125 234.105 166.595 ;
        RECT 237.335 163.125 240.805 166.595 ;
        RECT 244.035 163.125 247.505 166.595 ;
        RECT 250.735 163.125 254.205 166.595 ;
        RECT 257.435 163.125 260.905 166.595 ;
        RECT 82.600 146.735 84.760 149.585 ;
        RECT 82.600 141.935 84.760 144.785 ;
        RECT 92.640 141.935 94.800 149.585 ;
        RECT 96.320 146.735 98.480 149.585 ;
        RECT 96.320 141.935 98.480 144.785 ;
        RECT 106.360 141.935 108.520 149.585 ;
        RECT 110.040 141.935 112.200 144.785 ;
        RECT 120.080 141.935 122.240 149.585 ;
        RECT 136.010 146.735 138.170 149.585 ;
        RECT 136.010 141.935 138.170 144.785 ;
        RECT 146.050 141.935 148.210 149.585 ;
        RECT 187.595 142.710 187.765 149.605 ;
        RECT 192.175 142.710 192.345 149.605 ;
        RECT 192.885 142.710 193.055 142.715 ;
        RECT 196.755 142.710 196.925 149.605 ;
        RECT 201.335 142.710 201.505 149.605 ;
        RECT 210.535 144.325 214.005 147.795 ;
        RECT 217.235 144.325 220.705 147.795 ;
        RECT 223.935 144.325 227.405 147.795 ;
        RECT 230.635 144.325 234.105 147.795 ;
        RECT 237.335 144.325 240.805 147.795 ;
        RECT 244.035 144.325 247.505 147.795 ;
        RECT 250.735 144.325 254.205 147.795 ;
        RECT 257.435 144.325 260.905 147.795 ;
        RECT 187.360 142.410 201.740 142.710 ;
        RECT 187.360 141.880 201.740 142.180 ;
        RECT 192.885 141.865 193.055 141.880 ;
        RECT 112.000 127.935 114.160 130.785 ;
        RECT 112.000 123.135 114.160 125.985 ;
        RECT 122.040 123.135 124.200 130.785 ;
        RECT 127.150 125.830 127.320 129.580 ;
        RECT 131.730 125.830 131.900 129.580 ;
        RECT 136.310 125.830 136.480 129.580 ;
        RECT 140.890 125.830 141.060 129.580 ;
        RECT 145.470 125.830 145.640 129.580 ;
        RECT 186.970 127.935 189.130 130.785 ;
        RECT 127.145 125.540 127.320 125.830 ;
        RECT 131.725 125.540 131.900 125.830 ;
        RECT 136.305 125.540 136.480 125.830 ;
        RECT 140.885 125.540 141.060 125.830 ;
        RECT 145.465 125.540 145.640 125.830 ;
        RECT 127.145 125.210 127.315 125.540 ;
        RECT 131.725 125.210 131.895 125.540 ;
        RECT 136.305 125.210 136.475 125.540 ;
        RECT 140.885 125.210 141.055 125.540 ;
        RECT 145.465 125.210 145.635 125.540 ;
        RECT 127.090 124.910 147.990 125.210 ;
        RECT 186.970 123.135 189.130 125.985 ;
        RECT 197.010 123.135 199.170 130.785 ;
        RECT 200.690 127.935 202.850 130.785 ;
        RECT 200.690 123.135 202.850 125.985 ;
        RECT 210.730 123.135 212.890 130.785 ;
        RECT 214.410 127.935 216.570 130.785 ;
        RECT 214.410 123.135 216.570 125.985 ;
        RECT 224.450 123.135 226.610 130.785 ;
        RECT 228.130 127.935 230.290 130.785 ;
        RECT 238.170 123.135 240.330 130.785 ;
        RECT 241.850 127.935 244.010 130.785 ;
        RECT 241.850 123.135 244.010 125.985 ;
        RECT 251.890 123.135 254.050 130.785 ;
        RECT 119.350 109.135 121.510 111.985 ;
        RECT 119.350 104.335 121.510 107.185 ;
        RECT 129.390 104.335 131.550 111.985 ;
        RECT 136.010 109.135 138.170 111.985 ;
        RECT 136.010 104.335 138.170 107.185 ;
        RECT 146.050 104.335 148.210 111.985 ;
        RECT 149.730 109.135 151.890 111.985 ;
        RECT 149.730 104.335 151.890 107.185 ;
        RECT 159.770 104.335 161.930 111.985 ;
        RECT 165.900 109.135 168.060 111.985 ;
        RECT 165.900 104.335 168.060 107.185 ;
        RECT 175.940 104.335 178.100 111.985 ;
        RECT 186.970 109.135 189.130 111.985 ;
        RECT 186.970 104.335 189.130 107.185 ;
        RECT 197.010 104.335 199.170 111.985 ;
        RECT 200.690 109.135 202.850 111.985 ;
        RECT 200.690 104.335 202.850 107.185 ;
        RECT 210.730 104.335 212.890 111.985 ;
        RECT 241.850 104.335 244.010 107.185 ;
        RECT 251.890 104.335 254.050 111.985 ;
        RECT 124.150 85.480 262.190 85.780 ;
        RECT 219.310 71.535 221.470 74.385 ;
        RECT 219.310 66.735 221.470 69.585 ;
        RECT 229.350 66.735 231.510 74.385 ;
        RECT 233.030 71.535 235.190 74.385 ;
        RECT 233.030 66.735 235.190 69.585 ;
        RECT 243.070 66.735 245.230 74.385 ;
        RECT 246.750 71.535 248.910 74.385 ;
        RECT 246.750 66.735 248.910 69.585 ;
        RECT 256.790 66.735 258.950 74.385 ;
        RECT 218.820 47.935 220.980 50.785 ;
        RECT 228.860 47.935 231.020 55.585 ;
        RECT 232.540 52.735 234.700 55.585 ;
        RECT 232.540 47.935 234.700 50.785 ;
        RECT 242.580 47.935 244.740 55.585 ;
        RECT 246.260 52.735 248.420 55.585 ;
        RECT 246.260 47.935 248.420 50.785 ;
        RECT 256.300 47.935 258.460 55.585 ;
        RECT 222.740 33.935 224.900 36.785 ;
        RECT 222.740 29.135 224.900 31.985 ;
        RECT 232.780 29.135 234.940 36.785 ;
        RECT 236.460 33.935 238.620 36.785 ;
        RECT 246.500 29.135 248.660 36.785 ;
        RECT 250.180 33.935 252.340 36.785 ;
        RECT 250.180 29.135 252.340 31.985 ;
        RECT 260.220 29.135 262.380 36.785 ;
      LAYER mcon ;
        RECT 104.255 240.815 106.225 243.505 ;
        RECT 114.290 240.815 116.260 243.505 ;
        RECT 104.255 236.015 106.225 238.705 ;
        RECT 114.290 236.015 116.260 238.705 ;
        RECT 119.650 242.075 119.820 242.245 ;
        RECT 119.650 241.715 119.820 241.885 ;
        RECT 119.650 241.355 119.820 241.525 ;
        RECT 119.650 240.995 119.820 241.165 ;
        RECT 119.650 240.635 119.820 240.805 ;
        RECT 119.650 240.275 119.820 240.445 ;
        RECT 119.650 239.915 119.820 240.085 ;
        RECT 119.650 239.555 119.820 239.725 ;
        RECT 119.650 239.195 119.820 239.365 ;
        RECT 119.650 238.835 119.820 239.005 ;
        RECT 119.650 238.475 119.820 238.645 ;
        RECT 147.345 236.045 147.515 236.215 ;
        RECT 70.650 223.275 70.820 223.445 ;
        RECT 70.650 222.915 70.820 223.085 ;
        RECT 70.650 222.555 70.820 222.725 ;
        RECT 70.650 222.195 70.820 222.365 ;
        RECT 70.650 221.835 70.820 222.005 ;
        RECT 70.650 221.475 70.820 221.645 ;
        RECT 70.650 221.115 70.820 221.285 ;
        RECT 70.650 220.755 70.820 220.925 ;
        RECT 70.650 220.395 70.820 220.565 ;
        RECT 70.650 220.035 70.820 220.205 ;
        RECT 70.650 219.675 70.820 219.845 ;
        RECT 216.780 222.390 216.950 222.560 ;
        RECT 217.280 222.390 217.450 222.560 ;
        RECT 217.780 222.390 217.950 222.560 ;
        RECT 218.280 222.390 218.450 222.560 ;
        RECT 218.780 222.390 218.950 222.560 ;
        RECT 219.280 222.390 219.450 222.560 ;
        RECT 216.780 221.890 216.950 222.060 ;
        RECT 217.280 221.890 217.450 222.060 ;
        RECT 217.780 221.890 217.950 222.060 ;
        RECT 218.280 221.890 218.450 222.060 ;
        RECT 218.780 221.890 218.950 222.060 ;
        RECT 219.280 221.890 219.450 222.060 ;
        RECT 216.780 221.390 216.950 221.560 ;
        RECT 217.280 221.390 217.450 221.560 ;
        RECT 217.780 221.390 217.950 221.560 ;
        RECT 218.280 221.390 218.450 221.560 ;
        RECT 218.780 221.390 218.950 221.560 ;
        RECT 219.280 221.390 219.450 221.560 ;
        RECT 216.780 220.890 216.950 221.060 ;
        RECT 217.280 220.890 217.450 221.060 ;
        RECT 217.780 220.890 217.950 221.060 ;
        RECT 218.280 220.890 218.450 221.060 ;
        RECT 218.780 220.890 218.950 221.060 ;
        RECT 219.280 220.890 219.450 221.060 ;
        RECT 216.780 220.390 216.950 220.560 ;
        RECT 217.280 220.390 217.450 220.560 ;
        RECT 217.780 220.390 217.950 220.560 ;
        RECT 218.280 220.390 218.450 220.560 ;
        RECT 218.780 220.390 218.950 220.560 ;
        RECT 219.280 220.390 219.450 220.560 ;
        RECT 216.780 219.890 216.950 220.060 ;
        RECT 217.280 219.890 217.450 220.060 ;
        RECT 217.780 219.890 217.950 220.060 ;
        RECT 218.280 219.890 218.450 220.060 ;
        RECT 218.780 219.890 218.950 220.060 ;
        RECT 219.280 219.890 219.450 220.060 ;
        RECT 223.480 222.390 223.650 222.560 ;
        RECT 223.980 222.390 224.150 222.560 ;
        RECT 224.480 222.390 224.650 222.560 ;
        RECT 224.980 222.390 225.150 222.560 ;
        RECT 225.480 222.390 225.650 222.560 ;
        RECT 225.980 222.390 226.150 222.560 ;
        RECT 223.480 221.890 223.650 222.060 ;
        RECT 223.980 221.890 224.150 222.060 ;
        RECT 224.480 221.890 224.650 222.060 ;
        RECT 224.980 221.890 225.150 222.060 ;
        RECT 225.480 221.890 225.650 222.060 ;
        RECT 225.980 221.890 226.150 222.060 ;
        RECT 223.480 221.390 223.650 221.560 ;
        RECT 223.980 221.390 224.150 221.560 ;
        RECT 224.480 221.390 224.650 221.560 ;
        RECT 224.980 221.390 225.150 221.560 ;
        RECT 225.480 221.390 225.650 221.560 ;
        RECT 225.980 221.390 226.150 221.560 ;
        RECT 223.480 220.890 223.650 221.060 ;
        RECT 223.980 220.890 224.150 221.060 ;
        RECT 224.480 220.890 224.650 221.060 ;
        RECT 224.980 220.890 225.150 221.060 ;
        RECT 225.480 220.890 225.650 221.060 ;
        RECT 225.980 220.890 226.150 221.060 ;
        RECT 223.480 220.390 223.650 220.560 ;
        RECT 223.980 220.390 224.150 220.560 ;
        RECT 224.480 220.390 224.650 220.560 ;
        RECT 224.980 220.390 225.150 220.560 ;
        RECT 225.480 220.390 225.650 220.560 ;
        RECT 225.980 220.390 226.150 220.560 ;
        RECT 223.480 219.890 223.650 220.060 ;
        RECT 223.980 219.890 224.150 220.060 ;
        RECT 224.480 219.890 224.650 220.060 ;
        RECT 224.980 219.890 225.150 220.060 ;
        RECT 225.480 219.890 225.650 220.060 ;
        RECT 225.980 219.890 226.150 220.060 ;
        RECT 230.180 222.390 230.350 222.560 ;
        RECT 230.680 222.390 230.850 222.560 ;
        RECT 231.180 222.390 231.350 222.560 ;
        RECT 231.680 222.390 231.850 222.560 ;
        RECT 232.180 222.390 232.350 222.560 ;
        RECT 232.680 222.390 232.850 222.560 ;
        RECT 230.180 221.890 230.350 222.060 ;
        RECT 230.680 221.890 230.850 222.060 ;
        RECT 231.180 221.890 231.350 222.060 ;
        RECT 231.680 221.890 231.850 222.060 ;
        RECT 232.180 221.890 232.350 222.060 ;
        RECT 232.680 221.890 232.850 222.060 ;
        RECT 230.180 221.390 230.350 221.560 ;
        RECT 230.680 221.390 230.850 221.560 ;
        RECT 231.180 221.390 231.350 221.560 ;
        RECT 231.680 221.390 231.850 221.560 ;
        RECT 232.180 221.390 232.350 221.560 ;
        RECT 232.680 221.390 232.850 221.560 ;
        RECT 230.180 220.890 230.350 221.060 ;
        RECT 230.680 220.890 230.850 221.060 ;
        RECT 231.180 220.890 231.350 221.060 ;
        RECT 231.680 220.890 231.850 221.060 ;
        RECT 232.180 220.890 232.350 221.060 ;
        RECT 232.680 220.890 232.850 221.060 ;
        RECT 230.180 220.390 230.350 220.560 ;
        RECT 230.680 220.390 230.850 220.560 ;
        RECT 231.180 220.390 231.350 220.560 ;
        RECT 231.680 220.390 231.850 220.560 ;
        RECT 232.180 220.390 232.350 220.560 ;
        RECT 232.680 220.390 232.850 220.560 ;
        RECT 230.180 219.890 230.350 220.060 ;
        RECT 230.680 219.890 230.850 220.060 ;
        RECT 231.180 219.890 231.350 220.060 ;
        RECT 231.680 219.890 231.850 220.060 ;
        RECT 232.180 219.890 232.350 220.060 ;
        RECT 232.680 219.890 232.850 220.060 ;
        RECT 236.880 222.390 237.050 222.560 ;
        RECT 237.380 222.390 237.550 222.560 ;
        RECT 237.880 222.390 238.050 222.560 ;
        RECT 238.380 222.390 238.550 222.560 ;
        RECT 238.880 222.390 239.050 222.560 ;
        RECT 239.380 222.390 239.550 222.560 ;
        RECT 236.880 221.890 237.050 222.060 ;
        RECT 237.380 221.890 237.550 222.060 ;
        RECT 237.880 221.890 238.050 222.060 ;
        RECT 238.380 221.890 238.550 222.060 ;
        RECT 238.880 221.890 239.050 222.060 ;
        RECT 239.380 221.890 239.550 222.060 ;
        RECT 236.880 221.390 237.050 221.560 ;
        RECT 237.380 221.390 237.550 221.560 ;
        RECT 237.880 221.390 238.050 221.560 ;
        RECT 238.380 221.390 238.550 221.560 ;
        RECT 238.880 221.390 239.050 221.560 ;
        RECT 239.380 221.390 239.550 221.560 ;
        RECT 236.880 220.890 237.050 221.060 ;
        RECT 237.380 220.890 237.550 221.060 ;
        RECT 237.880 220.890 238.050 221.060 ;
        RECT 238.380 220.890 238.550 221.060 ;
        RECT 238.880 220.890 239.050 221.060 ;
        RECT 239.380 220.890 239.550 221.060 ;
        RECT 236.880 220.390 237.050 220.560 ;
        RECT 237.380 220.390 237.550 220.560 ;
        RECT 237.880 220.390 238.050 220.560 ;
        RECT 238.380 220.390 238.550 220.560 ;
        RECT 238.880 220.390 239.050 220.560 ;
        RECT 239.380 220.390 239.550 220.560 ;
        RECT 236.880 219.890 237.050 220.060 ;
        RECT 237.380 219.890 237.550 220.060 ;
        RECT 237.880 219.890 238.050 220.060 ;
        RECT 238.380 219.890 238.550 220.060 ;
        RECT 238.880 219.890 239.050 220.060 ;
        RECT 239.380 219.890 239.550 220.060 ;
        RECT 243.580 222.390 243.750 222.560 ;
        RECT 244.080 222.390 244.250 222.560 ;
        RECT 244.580 222.390 244.750 222.560 ;
        RECT 245.080 222.390 245.250 222.560 ;
        RECT 245.580 222.390 245.750 222.560 ;
        RECT 246.080 222.390 246.250 222.560 ;
        RECT 243.580 221.890 243.750 222.060 ;
        RECT 244.080 221.890 244.250 222.060 ;
        RECT 244.580 221.890 244.750 222.060 ;
        RECT 245.080 221.890 245.250 222.060 ;
        RECT 245.580 221.890 245.750 222.060 ;
        RECT 246.080 221.890 246.250 222.060 ;
        RECT 243.580 221.390 243.750 221.560 ;
        RECT 244.080 221.390 244.250 221.560 ;
        RECT 244.580 221.390 244.750 221.560 ;
        RECT 245.080 221.390 245.250 221.560 ;
        RECT 245.580 221.390 245.750 221.560 ;
        RECT 246.080 221.390 246.250 221.560 ;
        RECT 243.580 220.890 243.750 221.060 ;
        RECT 244.080 220.890 244.250 221.060 ;
        RECT 244.580 220.890 244.750 221.060 ;
        RECT 245.080 220.890 245.250 221.060 ;
        RECT 245.580 220.890 245.750 221.060 ;
        RECT 246.080 220.890 246.250 221.060 ;
        RECT 243.580 220.390 243.750 220.560 ;
        RECT 244.080 220.390 244.250 220.560 ;
        RECT 244.580 220.390 244.750 220.560 ;
        RECT 245.080 220.390 245.250 220.560 ;
        RECT 245.580 220.390 245.750 220.560 ;
        RECT 246.080 220.390 246.250 220.560 ;
        RECT 243.580 219.890 243.750 220.060 ;
        RECT 244.080 219.890 244.250 220.060 ;
        RECT 244.580 219.890 244.750 220.060 ;
        RECT 245.080 219.890 245.250 220.060 ;
        RECT 245.580 219.890 245.750 220.060 ;
        RECT 246.080 219.890 246.250 220.060 ;
        RECT 250.280 222.390 250.450 222.560 ;
        RECT 250.780 222.390 250.950 222.560 ;
        RECT 251.280 222.390 251.450 222.560 ;
        RECT 251.780 222.390 251.950 222.560 ;
        RECT 252.280 222.390 252.450 222.560 ;
        RECT 252.780 222.390 252.950 222.560 ;
        RECT 250.280 221.890 250.450 222.060 ;
        RECT 250.780 221.890 250.950 222.060 ;
        RECT 251.280 221.890 251.450 222.060 ;
        RECT 251.780 221.890 251.950 222.060 ;
        RECT 252.280 221.890 252.450 222.060 ;
        RECT 252.780 221.890 252.950 222.060 ;
        RECT 250.280 221.390 250.450 221.560 ;
        RECT 250.780 221.390 250.950 221.560 ;
        RECT 251.280 221.390 251.450 221.560 ;
        RECT 251.780 221.390 251.950 221.560 ;
        RECT 252.280 221.390 252.450 221.560 ;
        RECT 252.780 221.390 252.950 221.560 ;
        RECT 250.280 220.890 250.450 221.060 ;
        RECT 250.780 220.890 250.950 221.060 ;
        RECT 251.280 220.890 251.450 221.060 ;
        RECT 251.780 220.890 251.950 221.060 ;
        RECT 252.280 220.890 252.450 221.060 ;
        RECT 252.780 220.890 252.950 221.060 ;
        RECT 250.280 220.390 250.450 220.560 ;
        RECT 250.780 220.390 250.950 220.560 ;
        RECT 251.280 220.390 251.450 220.560 ;
        RECT 251.780 220.390 251.950 220.560 ;
        RECT 252.280 220.390 252.450 220.560 ;
        RECT 252.780 220.390 252.950 220.560 ;
        RECT 250.280 219.890 250.450 220.060 ;
        RECT 250.780 219.890 250.950 220.060 ;
        RECT 251.280 219.890 251.450 220.060 ;
        RECT 251.780 219.890 251.950 220.060 ;
        RECT 252.280 219.890 252.450 220.060 ;
        RECT 252.780 219.890 252.950 220.060 ;
        RECT 256.980 222.390 257.150 222.560 ;
        RECT 257.480 222.390 257.650 222.560 ;
        RECT 257.980 222.390 258.150 222.560 ;
        RECT 258.480 222.390 258.650 222.560 ;
        RECT 258.980 222.390 259.150 222.560 ;
        RECT 259.480 222.390 259.650 222.560 ;
        RECT 256.980 221.890 257.150 222.060 ;
        RECT 257.480 221.890 257.650 222.060 ;
        RECT 257.980 221.890 258.150 222.060 ;
        RECT 258.480 221.890 258.650 222.060 ;
        RECT 258.980 221.890 259.150 222.060 ;
        RECT 259.480 221.890 259.650 222.060 ;
        RECT 256.980 221.390 257.150 221.560 ;
        RECT 257.480 221.390 257.650 221.560 ;
        RECT 257.980 221.390 258.150 221.560 ;
        RECT 258.480 221.390 258.650 221.560 ;
        RECT 258.980 221.390 259.150 221.560 ;
        RECT 259.480 221.390 259.650 221.560 ;
        RECT 256.980 220.890 257.150 221.060 ;
        RECT 257.480 220.890 257.650 221.060 ;
        RECT 257.980 220.890 258.150 221.060 ;
        RECT 258.480 220.890 258.650 221.060 ;
        RECT 258.980 220.890 259.150 221.060 ;
        RECT 259.480 220.890 259.650 221.060 ;
        RECT 256.980 220.390 257.150 220.560 ;
        RECT 257.480 220.390 257.650 220.560 ;
        RECT 257.980 220.390 258.150 220.560 ;
        RECT 258.480 220.390 258.650 220.560 ;
        RECT 258.980 220.390 259.150 220.560 ;
        RECT 259.480 220.390 259.650 220.560 ;
        RECT 256.980 219.890 257.150 220.060 ;
        RECT 257.480 219.890 257.650 220.060 ;
        RECT 257.980 219.890 258.150 220.060 ;
        RECT 258.480 219.890 258.650 220.060 ;
        RECT 258.980 219.890 259.150 220.060 ;
        RECT 259.480 219.890 259.650 220.060 ;
        RECT 72.825 217.345 72.995 217.515 ;
        RECT 147.345 217.175 147.515 217.345 ;
        RECT 146.925 205.735 147.095 205.905 ;
        RECT 146.925 205.375 147.095 205.545 ;
        RECT 146.925 205.015 147.095 205.185 ;
        RECT 146.925 204.655 147.095 204.825 ;
        RECT 146.925 204.295 147.095 204.465 ;
        RECT 146.925 203.935 147.095 204.105 ;
        RECT 146.925 203.575 147.095 203.745 ;
        RECT 146.925 203.215 147.095 203.385 ;
        RECT 146.925 202.855 147.095 203.025 ;
        RECT 146.925 202.495 147.095 202.665 ;
        RECT 146.925 202.135 147.095 202.305 ;
        RECT 146.925 201.775 147.095 201.945 ;
        RECT 146.925 201.415 147.095 201.585 ;
        RECT 146.925 201.055 147.095 201.225 ;
        RECT 146.925 200.695 147.095 200.865 ;
        RECT 146.925 200.335 147.095 200.505 ;
        RECT 146.925 199.975 147.095 200.145 ;
        RECT 146.925 199.615 147.095 199.785 ;
        RECT 151.505 205.735 151.675 205.905 ;
        RECT 151.505 205.375 151.675 205.545 ;
        RECT 151.505 205.015 151.675 205.185 ;
        RECT 151.505 204.655 151.675 204.825 ;
        RECT 151.505 204.295 151.675 204.465 ;
        RECT 151.505 203.935 151.675 204.105 ;
        RECT 151.505 203.575 151.675 203.745 ;
        RECT 151.505 203.215 151.675 203.385 ;
        RECT 151.505 202.855 151.675 203.025 ;
        RECT 151.505 202.495 151.675 202.665 ;
        RECT 151.505 202.135 151.675 202.305 ;
        RECT 151.505 201.775 151.675 201.945 ;
        RECT 151.505 201.415 151.675 201.585 ;
        RECT 151.505 201.055 151.675 201.225 ;
        RECT 151.505 200.695 151.675 200.865 ;
        RECT 151.505 200.335 151.675 200.505 ;
        RECT 151.505 199.975 151.675 200.145 ;
        RECT 151.505 199.615 151.675 199.785 ;
        RECT 156.085 205.735 156.255 205.905 ;
        RECT 156.085 205.375 156.255 205.545 ;
        RECT 156.085 205.015 156.255 205.185 ;
        RECT 156.085 204.655 156.255 204.825 ;
        RECT 156.085 204.295 156.255 204.465 ;
        RECT 156.085 203.935 156.255 204.105 ;
        RECT 156.085 203.575 156.255 203.745 ;
        RECT 156.085 203.215 156.255 203.385 ;
        RECT 156.085 202.855 156.255 203.025 ;
        RECT 156.085 202.495 156.255 202.665 ;
        RECT 156.085 202.135 156.255 202.305 ;
        RECT 156.085 201.775 156.255 201.945 ;
        RECT 156.085 201.415 156.255 201.585 ;
        RECT 156.085 201.055 156.255 201.225 ;
        RECT 156.085 200.695 156.255 200.865 ;
        RECT 156.085 200.335 156.255 200.505 ;
        RECT 156.085 199.975 156.255 200.145 ;
        RECT 156.085 199.615 156.255 199.785 ;
        RECT 160.665 205.735 160.835 205.905 ;
        RECT 160.665 205.375 160.835 205.545 ;
        RECT 160.665 205.015 160.835 205.185 ;
        RECT 160.665 204.655 160.835 204.825 ;
        RECT 160.665 204.295 160.835 204.465 ;
        RECT 160.665 203.935 160.835 204.105 ;
        RECT 160.665 203.575 160.835 203.745 ;
        RECT 160.665 203.215 160.835 203.385 ;
        RECT 160.665 202.855 160.835 203.025 ;
        RECT 160.665 202.495 160.835 202.665 ;
        RECT 160.665 202.135 160.835 202.305 ;
        RECT 160.665 201.775 160.835 201.945 ;
        RECT 160.665 201.415 160.835 201.585 ;
        RECT 160.665 201.055 160.835 201.225 ;
        RECT 160.665 200.695 160.835 200.865 ;
        RECT 160.665 200.335 160.835 200.505 ;
        RECT 160.665 199.975 160.835 200.145 ;
        RECT 160.665 199.615 160.835 199.785 ;
        RECT 165.245 205.735 165.415 205.905 ;
        RECT 165.245 205.375 165.415 205.545 ;
        RECT 165.245 205.015 165.415 205.185 ;
        RECT 165.245 204.655 165.415 204.825 ;
        RECT 165.245 204.295 165.415 204.465 ;
        RECT 165.245 203.935 165.415 204.105 ;
        RECT 165.245 203.575 165.415 203.745 ;
        RECT 165.245 203.215 165.415 203.385 ;
        RECT 165.245 202.855 165.415 203.025 ;
        RECT 165.245 202.495 165.415 202.665 ;
        RECT 165.245 202.135 165.415 202.305 ;
        RECT 165.245 201.775 165.415 201.945 ;
        RECT 165.245 201.415 165.415 201.585 ;
        RECT 165.245 201.055 165.415 201.225 ;
        RECT 165.245 200.695 165.415 200.865 ;
        RECT 165.245 200.335 165.415 200.505 ;
        RECT 165.245 199.975 165.415 200.145 ;
        RECT 165.245 199.615 165.415 199.785 ;
        RECT 169.825 205.735 169.995 205.905 ;
        RECT 169.825 205.375 169.995 205.545 ;
        RECT 169.825 205.015 169.995 205.185 ;
        RECT 169.825 204.655 169.995 204.825 ;
        RECT 169.825 204.295 169.995 204.465 ;
        RECT 169.825 203.935 169.995 204.105 ;
        RECT 169.825 203.575 169.995 203.745 ;
        RECT 169.825 203.215 169.995 203.385 ;
        RECT 169.825 202.855 169.995 203.025 ;
        RECT 169.825 202.495 169.995 202.665 ;
        RECT 169.825 202.135 169.995 202.305 ;
        RECT 169.825 201.775 169.995 201.945 ;
        RECT 169.825 201.415 169.995 201.585 ;
        RECT 169.825 201.055 169.995 201.225 ;
        RECT 169.825 200.695 169.995 200.865 ;
        RECT 169.825 200.335 169.995 200.505 ;
        RECT 169.825 199.975 169.995 200.145 ;
        RECT 169.825 199.615 169.995 199.785 ;
        RECT 174.405 205.735 174.575 205.905 ;
        RECT 174.405 205.375 174.575 205.545 ;
        RECT 174.405 205.015 174.575 205.185 ;
        RECT 174.405 204.655 174.575 204.825 ;
        RECT 174.405 204.295 174.575 204.465 ;
        RECT 174.405 203.935 174.575 204.105 ;
        RECT 174.405 203.575 174.575 203.745 ;
        RECT 174.405 203.215 174.575 203.385 ;
        RECT 174.405 202.855 174.575 203.025 ;
        RECT 174.405 202.495 174.575 202.665 ;
        RECT 174.405 202.135 174.575 202.305 ;
        RECT 174.405 201.775 174.575 201.945 ;
        RECT 174.405 201.415 174.575 201.585 ;
        RECT 174.405 201.055 174.575 201.225 ;
        RECT 186.440 204.475 186.610 204.645 ;
        RECT 186.440 204.115 186.610 204.285 ;
        RECT 186.440 203.755 186.610 203.925 ;
        RECT 186.440 203.395 186.610 203.565 ;
        RECT 186.440 203.035 186.610 203.205 ;
        RECT 186.440 202.675 186.610 202.845 ;
        RECT 186.440 202.315 186.610 202.485 ;
        RECT 186.440 201.955 186.610 202.125 ;
        RECT 186.440 201.595 186.610 201.765 ;
        RECT 186.440 201.235 186.610 201.405 ;
        RECT 174.405 200.695 174.575 200.865 ;
        RECT 174.405 200.335 174.575 200.505 ;
        RECT 186.440 200.875 186.610 201.045 ;
        RECT 188.730 204.475 188.900 204.645 ;
        RECT 188.730 204.115 188.900 204.285 ;
        RECT 188.730 203.755 188.900 203.925 ;
        RECT 188.730 203.395 188.900 203.565 ;
        RECT 188.730 203.035 188.900 203.205 ;
        RECT 188.730 202.675 188.900 202.845 ;
        RECT 188.730 202.315 188.900 202.485 ;
        RECT 188.730 201.955 188.900 202.125 ;
        RECT 188.730 201.595 188.900 201.765 ;
        RECT 188.730 201.235 188.900 201.405 ;
        RECT 188.730 200.875 188.900 201.045 ;
        RECT 191.020 204.475 191.190 204.645 ;
        RECT 191.020 204.115 191.190 204.285 ;
        RECT 191.020 203.755 191.190 203.925 ;
        RECT 191.020 203.395 191.190 203.565 ;
        RECT 191.020 203.035 191.190 203.205 ;
        RECT 191.020 202.675 191.190 202.845 ;
        RECT 191.020 202.315 191.190 202.485 ;
        RECT 191.020 201.955 191.190 202.125 ;
        RECT 191.020 201.595 191.190 201.765 ;
        RECT 191.020 201.235 191.190 201.405 ;
        RECT 191.020 200.875 191.190 201.045 ;
        RECT 193.310 204.475 193.480 204.645 ;
        RECT 193.310 204.115 193.480 204.285 ;
        RECT 193.310 203.755 193.480 203.925 ;
        RECT 193.310 203.395 193.480 203.565 ;
        RECT 193.310 203.035 193.480 203.205 ;
        RECT 193.310 202.675 193.480 202.845 ;
        RECT 193.310 202.315 193.480 202.485 ;
        RECT 193.310 201.955 193.480 202.125 ;
        RECT 193.310 201.595 193.480 201.765 ;
        RECT 193.310 201.235 193.480 201.405 ;
        RECT 193.310 200.875 193.480 201.045 ;
        RECT 195.600 204.475 195.770 204.645 ;
        RECT 195.600 204.115 195.770 204.285 ;
        RECT 195.600 203.755 195.770 203.925 ;
        RECT 195.600 203.395 195.770 203.565 ;
        RECT 195.600 203.035 195.770 203.205 ;
        RECT 195.600 202.675 195.770 202.845 ;
        RECT 195.600 202.315 195.770 202.485 ;
        RECT 195.600 201.955 195.770 202.125 ;
        RECT 195.600 201.595 195.770 201.765 ;
        RECT 195.600 201.235 195.770 201.405 ;
        RECT 195.600 200.875 195.770 201.045 ;
        RECT 197.890 204.475 198.060 204.645 ;
        RECT 197.890 204.115 198.060 204.285 ;
        RECT 197.890 203.755 198.060 203.925 ;
        RECT 197.890 203.395 198.060 203.565 ;
        RECT 197.890 203.035 198.060 203.205 ;
        RECT 197.890 202.675 198.060 202.845 ;
        RECT 197.890 202.315 198.060 202.485 ;
        RECT 197.890 201.955 198.060 202.125 ;
        RECT 197.890 201.595 198.060 201.765 ;
        RECT 197.890 201.235 198.060 201.405 ;
        RECT 197.890 200.875 198.060 201.045 ;
        RECT 200.180 204.475 200.350 204.645 ;
        RECT 200.180 204.115 200.350 204.285 ;
        RECT 200.180 203.755 200.350 203.925 ;
        RECT 200.180 203.395 200.350 203.565 ;
        RECT 200.180 203.035 200.350 203.205 ;
        RECT 200.180 202.675 200.350 202.845 ;
        RECT 200.180 202.315 200.350 202.485 ;
        RECT 200.180 201.955 200.350 202.125 ;
        RECT 200.180 201.595 200.350 201.765 ;
        RECT 200.180 201.235 200.350 201.405 ;
        RECT 200.180 200.875 200.350 201.045 ;
        RECT 202.470 204.475 202.640 204.645 ;
        RECT 202.470 204.115 202.640 204.285 ;
        RECT 202.470 203.755 202.640 203.925 ;
        RECT 202.470 203.395 202.640 203.565 ;
        RECT 202.470 203.035 202.640 203.205 ;
        RECT 202.470 202.675 202.640 202.845 ;
        RECT 202.470 202.315 202.640 202.485 ;
        RECT 202.470 201.955 202.640 202.125 ;
        RECT 202.470 201.595 202.640 201.765 ;
        RECT 202.470 201.235 202.640 201.405 ;
        RECT 202.470 200.875 202.640 201.045 ;
        RECT 204.760 204.475 204.930 204.645 ;
        RECT 204.760 204.115 204.930 204.285 ;
        RECT 204.760 203.755 204.930 203.925 ;
        RECT 204.760 203.395 204.930 203.565 ;
        RECT 204.760 203.035 204.930 203.205 ;
        RECT 204.760 202.675 204.930 202.845 ;
        RECT 204.760 202.315 204.930 202.485 ;
        RECT 204.760 201.955 204.930 202.125 ;
        RECT 204.760 201.595 204.930 201.765 ;
        RECT 204.760 201.235 204.930 201.405 ;
        RECT 204.760 200.875 204.930 201.045 ;
        RECT 207.050 204.475 207.220 204.645 ;
        RECT 207.050 204.115 207.220 204.285 ;
        RECT 207.050 203.755 207.220 203.925 ;
        RECT 207.050 203.395 207.220 203.565 ;
        RECT 207.050 203.035 207.220 203.205 ;
        RECT 207.050 202.675 207.220 202.845 ;
        RECT 207.050 202.315 207.220 202.485 ;
        RECT 207.050 201.955 207.220 202.125 ;
        RECT 207.050 201.595 207.220 201.765 ;
        RECT 207.050 201.235 207.220 201.405 ;
        RECT 207.050 200.875 207.220 201.045 ;
        RECT 210.900 203.590 211.070 203.760 ;
        RECT 211.400 203.590 211.570 203.760 ;
        RECT 211.900 203.590 212.070 203.760 ;
        RECT 212.400 203.590 212.570 203.760 ;
        RECT 212.900 203.590 213.070 203.760 ;
        RECT 213.400 203.590 213.570 203.760 ;
        RECT 210.900 203.090 211.070 203.260 ;
        RECT 211.400 203.090 211.570 203.260 ;
        RECT 211.900 203.090 212.070 203.260 ;
        RECT 212.400 203.090 212.570 203.260 ;
        RECT 212.900 203.090 213.070 203.260 ;
        RECT 213.400 203.090 213.570 203.260 ;
        RECT 210.900 202.590 211.070 202.760 ;
        RECT 211.400 202.590 211.570 202.760 ;
        RECT 211.900 202.590 212.070 202.760 ;
        RECT 212.400 202.590 212.570 202.760 ;
        RECT 212.900 202.590 213.070 202.760 ;
        RECT 213.400 202.590 213.570 202.760 ;
        RECT 210.900 202.090 211.070 202.260 ;
        RECT 211.400 202.090 211.570 202.260 ;
        RECT 211.900 202.090 212.070 202.260 ;
        RECT 212.400 202.090 212.570 202.260 ;
        RECT 212.900 202.090 213.070 202.260 ;
        RECT 213.400 202.090 213.570 202.260 ;
        RECT 210.900 201.590 211.070 201.760 ;
        RECT 211.400 201.590 211.570 201.760 ;
        RECT 211.900 201.590 212.070 201.760 ;
        RECT 212.400 201.590 212.570 201.760 ;
        RECT 212.900 201.590 213.070 201.760 ;
        RECT 213.400 201.590 213.570 201.760 ;
        RECT 210.900 201.090 211.070 201.260 ;
        RECT 211.400 201.090 211.570 201.260 ;
        RECT 211.900 201.090 212.070 201.260 ;
        RECT 212.400 201.090 212.570 201.260 ;
        RECT 212.900 201.090 213.070 201.260 ;
        RECT 213.400 201.090 213.570 201.260 ;
        RECT 217.600 203.590 217.770 203.760 ;
        RECT 218.100 203.590 218.270 203.760 ;
        RECT 218.600 203.590 218.770 203.760 ;
        RECT 219.100 203.590 219.270 203.760 ;
        RECT 219.600 203.590 219.770 203.760 ;
        RECT 220.100 203.590 220.270 203.760 ;
        RECT 217.600 203.090 217.770 203.260 ;
        RECT 218.100 203.090 218.270 203.260 ;
        RECT 218.600 203.090 218.770 203.260 ;
        RECT 219.100 203.090 219.270 203.260 ;
        RECT 219.600 203.090 219.770 203.260 ;
        RECT 220.100 203.090 220.270 203.260 ;
        RECT 217.600 202.590 217.770 202.760 ;
        RECT 218.100 202.590 218.270 202.760 ;
        RECT 218.600 202.590 218.770 202.760 ;
        RECT 219.100 202.590 219.270 202.760 ;
        RECT 219.600 202.590 219.770 202.760 ;
        RECT 220.100 202.590 220.270 202.760 ;
        RECT 217.600 202.090 217.770 202.260 ;
        RECT 218.100 202.090 218.270 202.260 ;
        RECT 218.600 202.090 218.770 202.260 ;
        RECT 219.100 202.090 219.270 202.260 ;
        RECT 219.600 202.090 219.770 202.260 ;
        RECT 220.100 202.090 220.270 202.260 ;
        RECT 217.600 201.590 217.770 201.760 ;
        RECT 218.100 201.590 218.270 201.760 ;
        RECT 218.600 201.590 218.770 201.760 ;
        RECT 219.100 201.590 219.270 201.760 ;
        RECT 219.600 201.590 219.770 201.760 ;
        RECT 220.100 201.590 220.270 201.760 ;
        RECT 217.600 201.090 217.770 201.260 ;
        RECT 218.100 201.090 218.270 201.260 ;
        RECT 218.600 201.090 218.770 201.260 ;
        RECT 219.100 201.090 219.270 201.260 ;
        RECT 219.600 201.090 219.770 201.260 ;
        RECT 220.100 201.090 220.270 201.260 ;
        RECT 224.300 203.590 224.470 203.760 ;
        RECT 224.800 203.590 224.970 203.760 ;
        RECT 225.300 203.590 225.470 203.760 ;
        RECT 225.800 203.590 225.970 203.760 ;
        RECT 226.300 203.590 226.470 203.760 ;
        RECT 226.800 203.590 226.970 203.760 ;
        RECT 224.300 203.090 224.470 203.260 ;
        RECT 224.800 203.090 224.970 203.260 ;
        RECT 225.300 203.090 225.470 203.260 ;
        RECT 225.800 203.090 225.970 203.260 ;
        RECT 226.300 203.090 226.470 203.260 ;
        RECT 226.800 203.090 226.970 203.260 ;
        RECT 224.300 202.590 224.470 202.760 ;
        RECT 224.800 202.590 224.970 202.760 ;
        RECT 225.300 202.590 225.470 202.760 ;
        RECT 225.800 202.590 225.970 202.760 ;
        RECT 226.300 202.590 226.470 202.760 ;
        RECT 226.800 202.590 226.970 202.760 ;
        RECT 224.300 202.090 224.470 202.260 ;
        RECT 224.800 202.090 224.970 202.260 ;
        RECT 225.300 202.090 225.470 202.260 ;
        RECT 225.800 202.090 225.970 202.260 ;
        RECT 226.300 202.090 226.470 202.260 ;
        RECT 226.800 202.090 226.970 202.260 ;
        RECT 224.300 201.590 224.470 201.760 ;
        RECT 224.800 201.590 224.970 201.760 ;
        RECT 225.300 201.590 225.470 201.760 ;
        RECT 225.800 201.590 225.970 201.760 ;
        RECT 226.300 201.590 226.470 201.760 ;
        RECT 226.800 201.590 226.970 201.760 ;
        RECT 224.300 201.090 224.470 201.260 ;
        RECT 224.800 201.090 224.970 201.260 ;
        RECT 225.300 201.090 225.470 201.260 ;
        RECT 225.800 201.090 225.970 201.260 ;
        RECT 226.300 201.090 226.470 201.260 ;
        RECT 226.800 201.090 226.970 201.260 ;
        RECT 231.000 203.590 231.170 203.760 ;
        RECT 231.500 203.590 231.670 203.760 ;
        RECT 232.000 203.590 232.170 203.760 ;
        RECT 232.500 203.590 232.670 203.760 ;
        RECT 233.000 203.590 233.170 203.760 ;
        RECT 233.500 203.590 233.670 203.760 ;
        RECT 231.000 203.090 231.170 203.260 ;
        RECT 231.500 203.090 231.670 203.260 ;
        RECT 232.000 203.090 232.170 203.260 ;
        RECT 232.500 203.090 232.670 203.260 ;
        RECT 233.000 203.090 233.170 203.260 ;
        RECT 233.500 203.090 233.670 203.260 ;
        RECT 231.000 202.590 231.170 202.760 ;
        RECT 231.500 202.590 231.670 202.760 ;
        RECT 232.000 202.590 232.170 202.760 ;
        RECT 232.500 202.590 232.670 202.760 ;
        RECT 233.000 202.590 233.170 202.760 ;
        RECT 233.500 202.590 233.670 202.760 ;
        RECT 231.000 202.090 231.170 202.260 ;
        RECT 231.500 202.090 231.670 202.260 ;
        RECT 232.000 202.090 232.170 202.260 ;
        RECT 232.500 202.090 232.670 202.260 ;
        RECT 233.000 202.090 233.170 202.260 ;
        RECT 233.500 202.090 233.670 202.260 ;
        RECT 231.000 201.590 231.170 201.760 ;
        RECT 231.500 201.590 231.670 201.760 ;
        RECT 232.000 201.590 232.170 201.760 ;
        RECT 232.500 201.590 232.670 201.760 ;
        RECT 233.000 201.590 233.170 201.760 ;
        RECT 233.500 201.590 233.670 201.760 ;
        RECT 231.000 201.090 231.170 201.260 ;
        RECT 231.500 201.090 231.670 201.260 ;
        RECT 232.000 201.090 232.170 201.260 ;
        RECT 232.500 201.090 232.670 201.260 ;
        RECT 233.000 201.090 233.170 201.260 ;
        RECT 233.500 201.090 233.670 201.260 ;
        RECT 237.700 203.590 237.870 203.760 ;
        RECT 238.200 203.590 238.370 203.760 ;
        RECT 238.700 203.590 238.870 203.760 ;
        RECT 239.200 203.590 239.370 203.760 ;
        RECT 239.700 203.590 239.870 203.760 ;
        RECT 240.200 203.590 240.370 203.760 ;
        RECT 237.700 203.090 237.870 203.260 ;
        RECT 238.200 203.090 238.370 203.260 ;
        RECT 238.700 203.090 238.870 203.260 ;
        RECT 239.200 203.090 239.370 203.260 ;
        RECT 239.700 203.090 239.870 203.260 ;
        RECT 240.200 203.090 240.370 203.260 ;
        RECT 237.700 202.590 237.870 202.760 ;
        RECT 238.200 202.590 238.370 202.760 ;
        RECT 238.700 202.590 238.870 202.760 ;
        RECT 239.200 202.590 239.370 202.760 ;
        RECT 239.700 202.590 239.870 202.760 ;
        RECT 240.200 202.590 240.370 202.760 ;
        RECT 237.700 202.090 237.870 202.260 ;
        RECT 238.200 202.090 238.370 202.260 ;
        RECT 238.700 202.090 238.870 202.260 ;
        RECT 239.200 202.090 239.370 202.260 ;
        RECT 239.700 202.090 239.870 202.260 ;
        RECT 240.200 202.090 240.370 202.260 ;
        RECT 237.700 201.590 237.870 201.760 ;
        RECT 238.200 201.590 238.370 201.760 ;
        RECT 238.700 201.590 238.870 201.760 ;
        RECT 239.200 201.590 239.370 201.760 ;
        RECT 239.700 201.590 239.870 201.760 ;
        RECT 240.200 201.590 240.370 201.760 ;
        RECT 237.700 201.090 237.870 201.260 ;
        RECT 238.200 201.090 238.370 201.260 ;
        RECT 238.700 201.090 238.870 201.260 ;
        RECT 239.200 201.090 239.370 201.260 ;
        RECT 239.700 201.090 239.870 201.260 ;
        RECT 240.200 201.090 240.370 201.260 ;
        RECT 244.400 203.590 244.570 203.760 ;
        RECT 244.900 203.590 245.070 203.760 ;
        RECT 245.400 203.590 245.570 203.760 ;
        RECT 245.900 203.590 246.070 203.760 ;
        RECT 246.400 203.590 246.570 203.760 ;
        RECT 246.900 203.590 247.070 203.760 ;
        RECT 244.400 203.090 244.570 203.260 ;
        RECT 244.900 203.090 245.070 203.260 ;
        RECT 245.400 203.090 245.570 203.260 ;
        RECT 245.900 203.090 246.070 203.260 ;
        RECT 246.400 203.090 246.570 203.260 ;
        RECT 246.900 203.090 247.070 203.260 ;
        RECT 244.400 202.590 244.570 202.760 ;
        RECT 244.900 202.590 245.070 202.760 ;
        RECT 245.400 202.590 245.570 202.760 ;
        RECT 245.900 202.590 246.070 202.760 ;
        RECT 246.400 202.590 246.570 202.760 ;
        RECT 246.900 202.590 247.070 202.760 ;
        RECT 244.400 202.090 244.570 202.260 ;
        RECT 244.900 202.090 245.070 202.260 ;
        RECT 245.400 202.090 245.570 202.260 ;
        RECT 245.900 202.090 246.070 202.260 ;
        RECT 246.400 202.090 246.570 202.260 ;
        RECT 246.900 202.090 247.070 202.260 ;
        RECT 244.400 201.590 244.570 201.760 ;
        RECT 244.900 201.590 245.070 201.760 ;
        RECT 245.400 201.590 245.570 201.760 ;
        RECT 245.900 201.590 246.070 201.760 ;
        RECT 246.400 201.590 246.570 201.760 ;
        RECT 246.900 201.590 247.070 201.760 ;
        RECT 244.400 201.090 244.570 201.260 ;
        RECT 244.900 201.090 245.070 201.260 ;
        RECT 245.400 201.090 245.570 201.260 ;
        RECT 245.900 201.090 246.070 201.260 ;
        RECT 246.400 201.090 246.570 201.260 ;
        RECT 246.900 201.090 247.070 201.260 ;
        RECT 251.100 203.590 251.270 203.760 ;
        RECT 251.600 203.590 251.770 203.760 ;
        RECT 252.100 203.590 252.270 203.760 ;
        RECT 252.600 203.590 252.770 203.760 ;
        RECT 253.100 203.590 253.270 203.760 ;
        RECT 253.600 203.590 253.770 203.760 ;
        RECT 251.100 203.090 251.270 203.260 ;
        RECT 251.600 203.090 251.770 203.260 ;
        RECT 252.100 203.090 252.270 203.260 ;
        RECT 252.600 203.090 252.770 203.260 ;
        RECT 253.100 203.090 253.270 203.260 ;
        RECT 253.600 203.090 253.770 203.260 ;
        RECT 251.100 202.590 251.270 202.760 ;
        RECT 251.600 202.590 251.770 202.760 ;
        RECT 252.100 202.590 252.270 202.760 ;
        RECT 252.600 202.590 252.770 202.760 ;
        RECT 253.100 202.590 253.270 202.760 ;
        RECT 253.600 202.590 253.770 202.760 ;
        RECT 251.100 202.090 251.270 202.260 ;
        RECT 251.600 202.090 251.770 202.260 ;
        RECT 252.100 202.090 252.270 202.260 ;
        RECT 252.600 202.090 252.770 202.260 ;
        RECT 253.100 202.090 253.270 202.260 ;
        RECT 253.600 202.090 253.770 202.260 ;
        RECT 251.100 201.590 251.270 201.760 ;
        RECT 251.600 201.590 251.770 201.760 ;
        RECT 252.100 201.590 252.270 201.760 ;
        RECT 252.600 201.590 252.770 201.760 ;
        RECT 253.100 201.590 253.270 201.760 ;
        RECT 253.600 201.590 253.770 201.760 ;
        RECT 251.100 201.090 251.270 201.260 ;
        RECT 251.600 201.090 251.770 201.260 ;
        RECT 252.100 201.090 252.270 201.260 ;
        RECT 252.600 201.090 252.770 201.260 ;
        RECT 253.100 201.090 253.270 201.260 ;
        RECT 253.600 201.090 253.770 201.260 ;
        RECT 257.800 203.590 257.970 203.760 ;
        RECT 258.300 203.590 258.470 203.760 ;
        RECT 258.800 203.590 258.970 203.760 ;
        RECT 259.300 203.590 259.470 203.760 ;
        RECT 259.800 203.590 259.970 203.760 ;
        RECT 260.300 203.590 260.470 203.760 ;
        RECT 257.800 203.090 257.970 203.260 ;
        RECT 258.300 203.090 258.470 203.260 ;
        RECT 258.800 203.090 258.970 203.260 ;
        RECT 259.300 203.090 259.470 203.260 ;
        RECT 259.800 203.090 259.970 203.260 ;
        RECT 260.300 203.090 260.470 203.260 ;
        RECT 257.800 202.590 257.970 202.760 ;
        RECT 258.300 202.590 258.470 202.760 ;
        RECT 258.800 202.590 258.970 202.760 ;
        RECT 259.300 202.590 259.470 202.760 ;
        RECT 259.800 202.590 259.970 202.760 ;
        RECT 260.300 202.590 260.470 202.760 ;
        RECT 257.800 202.090 257.970 202.260 ;
        RECT 258.300 202.090 258.470 202.260 ;
        RECT 258.800 202.090 258.970 202.260 ;
        RECT 259.300 202.090 259.470 202.260 ;
        RECT 259.800 202.090 259.970 202.260 ;
        RECT 260.300 202.090 260.470 202.260 ;
        RECT 257.800 201.590 257.970 201.760 ;
        RECT 258.300 201.590 258.470 201.760 ;
        RECT 258.800 201.590 258.970 201.760 ;
        RECT 259.300 201.590 259.470 201.760 ;
        RECT 259.800 201.590 259.970 201.760 ;
        RECT 260.300 201.590 260.470 201.760 ;
        RECT 257.800 201.090 257.970 201.260 ;
        RECT 258.300 201.090 258.470 201.260 ;
        RECT 258.800 201.090 258.970 201.260 ;
        RECT 259.300 201.090 259.470 201.260 ;
        RECT 259.800 201.090 259.970 201.260 ;
        RECT 260.300 201.090 260.470 201.260 ;
        RECT 174.405 199.975 174.575 200.145 ;
        RECT 174.405 199.615 174.575 199.785 ;
        RECT 147.345 198.305 147.515 198.475 ;
        RECT 68.485 184.415 70.455 187.105 ;
        RECT 78.520 184.415 80.490 187.105 ;
        RECT 68.485 179.615 70.455 182.305 ;
        RECT 82.205 184.415 84.175 187.105 ;
        RECT 92.240 184.415 94.210 187.105 ;
        RECT 78.520 179.615 80.490 182.305 ;
        RECT 82.205 179.615 84.175 182.305 ;
        RECT 95.930 184.415 97.900 187.105 ;
        RECT 108.835 184.415 110.805 187.105 ;
        RECT 92.240 179.615 94.210 182.305 ;
        RECT 112.585 184.415 114.555 187.105 ;
        RECT 122.620 184.415 124.590 187.105 ;
        RECT 187.595 186.935 187.765 187.105 ;
        RECT 187.595 186.575 187.765 186.745 ;
        RECT 187.595 186.215 187.765 186.385 ;
        RECT 108.835 179.615 110.805 182.305 ;
        RECT 112.585 179.615 114.555 182.305 ;
        RECT 122.620 179.615 124.590 182.305 ;
        RECT 127.150 185.675 127.320 185.845 ;
        RECT 127.150 185.315 127.320 185.485 ;
        RECT 127.150 184.955 127.320 185.125 ;
        RECT 127.150 184.595 127.320 184.765 ;
        RECT 127.150 184.235 127.320 184.405 ;
        RECT 127.150 183.875 127.320 184.045 ;
        RECT 127.150 183.515 127.320 183.685 ;
        RECT 127.150 183.155 127.320 183.325 ;
        RECT 127.150 182.795 127.320 182.965 ;
        RECT 127.150 182.435 127.320 182.605 ;
        RECT 127.150 182.075 127.320 182.245 ;
        RECT 129.440 185.675 129.610 185.845 ;
        RECT 129.440 185.315 129.610 185.485 ;
        RECT 129.440 184.955 129.610 185.125 ;
        RECT 129.440 184.595 129.610 184.765 ;
        RECT 129.440 184.235 129.610 184.405 ;
        RECT 129.440 183.875 129.610 184.045 ;
        RECT 129.440 183.515 129.610 183.685 ;
        RECT 129.440 183.155 129.610 183.325 ;
        RECT 129.440 182.795 129.610 182.965 ;
        RECT 129.440 182.435 129.610 182.605 ;
        RECT 129.440 182.075 129.610 182.245 ;
        RECT 131.730 185.675 131.900 185.845 ;
        RECT 131.730 185.315 131.900 185.485 ;
        RECT 131.730 184.955 131.900 185.125 ;
        RECT 131.730 184.595 131.900 184.765 ;
        RECT 131.730 184.235 131.900 184.405 ;
        RECT 131.730 183.875 131.900 184.045 ;
        RECT 131.730 183.515 131.900 183.685 ;
        RECT 131.730 183.155 131.900 183.325 ;
        RECT 131.730 182.795 131.900 182.965 ;
        RECT 131.730 182.435 131.900 182.605 ;
        RECT 131.730 182.075 131.900 182.245 ;
        RECT 134.020 185.675 134.190 185.845 ;
        RECT 134.020 185.315 134.190 185.485 ;
        RECT 134.020 184.955 134.190 185.125 ;
        RECT 134.020 184.595 134.190 184.765 ;
        RECT 134.020 184.235 134.190 184.405 ;
        RECT 134.020 183.875 134.190 184.045 ;
        RECT 134.020 183.515 134.190 183.685 ;
        RECT 134.020 183.155 134.190 183.325 ;
        RECT 134.020 182.795 134.190 182.965 ;
        RECT 134.020 182.435 134.190 182.605 ;
        RECT 134.020 182.075 134.190 182.245 ;
        RECT 136.310 185.675 136.480 185.845 ;
        RECT 136.310 185.315 136.480 185.485 ;
        RECT 136.310 184.955 136.480 185.125 ;
        RECT 136.310 184.595 136.480 184.765 ;
        RECT 136.310 184.235 136.480 184.405 ;
        RECT 136.310 183.875 136.480 184.045 ;
        RECT 136.310 183.515 136.480 183.685 ;
        RECT 136.310 183.155 136.480 183.325 ;
        RECT 136.310 182.795 136.480 182.965 ;
        RECT 136.310 182.435 136.480 182.605 ;
        RECT 136.310 182.075 136.480 182.245 ;
        RECT 138.600 185.675 138.770 185.845 ;
        RECT 138.600 185.315 138.770 185.485 ;
        RECT 138.600 184.955 138.770 185.125 ;
        RECT 138.600 184.595 138.770 184.765 ;
        RECT 138.600 184.235 138.770 184.405 ;
        RECT 138.600 183.875 138.770 184.045 ;
        RECT 138.600 183.515 138.770 183.685 ;
        RECT 138.600 183.155 138.770 183.325 ;
        RECT 138.600 182.795 138.770 182.965 ;
        RECT 138.600 182.435 138.770 182.605 ;
        RECT 138.600 182.075 138.770 182.245 ;
        RECT 140.890 185.675 141.060 185.845 ;
        RECT 140.890 185.315 141.060 185.485 ;
        RECT 140.890 184.955 141.060 185.125 ;
        RECT 140.890 184.595 141.060 184.765 ;
        RECT 140.890 184.235 141.060 184.405 ;
        RECT 140.890 183.875 141.060 184.045 ;
        RECT 140.890 183.515 141.060 183.685 ;
        RECT 140.890 183.155 141.060 183.325 ;
        RECT 140.890 182.795 141.060 182.965 ;
        RECT 140.890 182.435 141.060 182.605 ;
        RECT 140.890 182.075 141.060 182.245 ;
        RECT 143.180 185.675 143.350 185.845 ;
        RECT 143.180 185.315 143.350 185.485 ;
        RECT 143.180 184.955 143.350 185.125 ;
        RECT 143.180 184.595 143.350 184.765 ;
        RECT 143.180 184.235 143.350 184.405 ;
        RECT 143.180 183.875 143.350 184.045 ;
        RECT 143.180 183.515 143.350 183.685 ;
        RECT 143.180 183.155 143.350 183.325 ;
        RECT 143.180 182.795 143.350 182.965 ;
        RECT 143.180 182.435 143.350 182.605 ;
        RECT 143.180 182.075 143.350 182.245 ;
        RECT 145.470 185.675 145.640 185.845 ;
        RECT 145.470 185.315 145.640 185.485 ;
        RECT 145.470 184.955 145.640 185.125 ;
        RECT 145.470 184.595 145.640 184.765 ;
        RECT 145.470 184.235 145.640 184.405 ;
        RECT 145.470 183.875 145.640 184.045 ;
        RECT 145.470 183.515 145.640 183.685 ;
        RECT 145.470 183.155 145.640 183.325 ;
        RECT 145.470 182.795 145.640 182.965 ;
        RECT 145.470 182.435 145.640 182.605 ;
        RECT 145.470 182.075 145.640 182.245 ;
        RECT 147.760 185.675 147.930 185.845 ;
        RECT 147.760 185.315 147.930 185.485 ;
        RECT 147.760 184.955 147.930 185.125 ;
        RECT 147.760 184.595 147.930 184.765 ;
        RECT 147.760 184.235 147.930 184.405 ;
        RECT 147.760 183.875 147.930 184.045 ;
        RECT 147.760 183.515 147.930 183.685 ;
        RECT 147.760 183.155 147.930 183.325 ;
        RECT 147.760 182.795 147.930 182.965 ;
        RECT 147.760 182.435 147.930 182.605 ;
        RECT 147.760 182.075 147.930 182.245 ;
        RECT 187.595 185.855 187.765 186.025 ;
        RECT 187.595 185.495 187.765 185.665 ;
        RECT 187.595 185.135 187.765 185.305 ;
        RECT 187.595 184.775 187.765 184.945 ;
        RECT 187.595 184.415 187.765 184.585 ;
        RECT 187.595 184.055 187.765 184.225 ;
        RECT 187.595 183.695 187.765 183.865 ;
        RECT 187.595 183.335 187.765 183.505 ;
        RECT 187.595 182.975 187.765 183.145 ;
        RECT 187.595 182.615 187.765 182.785 ;
        RECT 187.595 182.255 187.765 182.425 ;
        RECT 187.595 181.895 187.765 182.065 ;
        RECT 187.595 181.535 187.765 181.705 ;
        RECT 187.595 181.175 187.765 181.345 ;
        RECT 187.595 180.815 187.765 180.985 ;
        RECT 192.175 186.935 192.345 187.105 ;
        RECT 192.175 186.575 192.345 186.745 ;
        RECT 192.175 186.215 192.345 186.385 ;
        RECT 192.175 185.855 192.345 186.025 ;
        RECT 192.175 185.495 192.345 185.665 ;
        RECT 192.175 185.135 192.345 185.305 ;
        RECT 192.175 184.775 192.345 184.945 ;
        RECT 192.175 184.415 192.345 184.585 ;
        RECT 192.175 184.055 192.345 184.225 ;
        RECT 192.175 183.695 192.345 183.865 ;
        RECT 192.175 183.335 192.345 183.505 ;
        RECT 192.175 182.975 192.345 183.145 ;
        RECT 192.175 182.615 192.345 182.785 ;
        RECT 192.175 182.255 192.345 182.425 ;
        RECT 192.175 181.895 192.345 182.065 ;
        RECT 192.175 181.535 192.345 181.705 ;
        RECT 192.175 181.175 192.345 181.345 ;
        RECT 192.175 180.815 192.345 180.985 ;
        RECT 196.755 186.935 196.925 187.105 ;
        RECT 196.755 186.575 196.925 186.745 ;
        RECT 196.755 186.215 196.925 186.385 ;
        RECT 196.755 185.855 196.925 186.025 ;
        RECT 196.755 185.495 196.925 185.665 ;
        RECT 196.755 185.135 196.925 185.305 ;
        RECT 196.755 184.775 196.925 184.945 ;
        RECT 196.755 184.415 196.925 184.585 ;
        RECT 196.755 184.055 196.925 184.225 ;
        RECT 196.755 183.695 196.925 183.865 ;
        RECT 196.755 183.335 196.925 183.505 ;
        RECT 196.755 182.975 196.925 183.145 ;
        RECT 196.755 182.615 196.925 182.785 ;
        RECT 196.755 182.255 196.925 182.425 ;
        RECT 196.755 181.895 196.925 182.065 ;
        RECT 196.755 181.535 196.925 181.705 ;
        RECT 196.755 181.175 196.925 181.345 ;
        RECT 196.755 180.815 196.925 180.985 ;
        RECT 201.335 186.935 201.505 187.105 ;
        RECT 201.335 186.575 201.505 186.745 ;
        RECT 201.335 186.215 201.505 186.385 ;
        RECT 201.335 185.855 201.505 186.025 ;
        RECT 201.335 185.495 201.505 185.665 ;
        RECT 201.335 185.135 201.505 185.305 ;
        RECT 201.335 184.775 201.505 184.945 ;
        RECT 201.335 184.415 201.505 184.585 ;
        RECT 201.335 184.055 201.505 184.225 ;
        RECT 201.335 183.695 201.505 183.865 ;
        RECT 201.335 183.335 201.505 183.505 ;
        RECT 201.335 182.975 201.505 183.145 ;
        RECT 201.335 182.615 201.505 182.785 ;
        RECT 201.335 182.255 201.505 182.425 ;
        RECT 201.335 181.895 201.505 182.065 ;
        RECT 210.900 184.790 211.070 184.960 ;
        RECT 211.400 184.790 211.570 184.960 ;
        RECT 211.900 184.790 212.070 184.960 ;
        RECT 212.400 184.790 212.570 184.960 ;
        RECT 212.900 184.790 213.070 184.960 ;
        RECT 213.400 184.790 213.570 184.960 ;
        RECT 210.900 184.290 211.070 184.460 ;
        RECT 211.400 184.290 211.570 184.460 ;
        RECT 211.900 184.290 212.070 184.460 ;
        RECT 212.400 184.290 212.570 184.460 ;
        RECT 212.900 184.290 213.070 184.460 ;
        RECT 213.400 184.290 213.570 184.460 ;
        RECT 210.900 183.790 211.070 183.960 ;
        RECT 211.400 183.790 211.570 183.960 ;
        RECT 211.900 183.790 212.070 183.960 ;
        RECT 212.400 183.790 212.570 183.960 ;
        RECT 212.900 183.790 213.070 183.960 ;
        RECT 213.400 183.790 213.570 183.960 ;
        RECT 210.900 183.290 211.070 183.460 ;
        RECT 211.400 183.290 211.570 183.460 ;
        RECT 211.900 183.290 212.070 183.460 ;
        RECT 212.400 183.290 212.570 183.460 ;
        RECT 212.900 183.290 213.070 183.460 ;
        RECT 213.400 183.290 213.570 183.460 ;
        RECT 210.900 182.790 211.070 182.960 ;
        RECT 211.400 182.790 211.570 182.960 ;
        RECT 211.900 182.790 212.070 182.960 ;
        RECT 212.400 182.790 212.570 182.960 ;
        RECT 212.900 182.790 213.070 182.960 ;
        RECT 213.400 182.790 213.570 182.960 ;
        RECT 210.900 182.290 211.070 182.460 ;
        RECT 211.400 182.290 211.570 182.460 ;
        RECT 211.900 182.290 212.070 182.460 ;
        RECT 212.400 182.290 212.570 182.460 ;
        RECT 212.900 182.290 213.070 182.460 ;
        RECT 213.400 182.290 213.570 182.460 ;
        RECT 217.600 184.790 217.770 184.960 ;
        RECT 218.100 184.790 218.270 184.960 ;
        RECT 218.600 184.790 218.770 184.960 ;
        RECT 219.100 184.790 219.270 184.960 ;
        RECT 219.600 184.790 219.770 184.960 ;
        RECT 220.100 184.790 220.270 184.960 ;
        RECT 217.600 184.290 217.770 184.460 ;
        RECT 218.100 184.290 218.270 184.460 ;
        RECT 218.600 184.290 218.770 184.460 ;
        RECT 219.100 184.290 219.270 184.460 ;
        RECT 219.600 184.290 219.770 184.460 ;
        RECT 220.100 184.290 220.270 184.460 ;
        RECT 217.600 183.790 217.770 183.960 ;
        RECT 218.100 183.790 218.270 183.960 ;
        RECT 218.600 183.790 218.770 183.960 ;
        RECT 219.100 183.790 219.270 183.960 ;
        RECT 219.600 183.790 219.770 183.960 ;
        RECT 220.100 183.790 220.270 183.960 ;
        RECT 217.600 183.290 217.770 183.460 ;
        RECT 218.100 183.290 218.270 183.460 ;
        RECT 218.600 183.290 218.770 183.460 ;
        RECT 219.100 183.290 219.270 183.460 ;
        RECT 219.600 183.290 219.770 183.460 ;
        RECT 220.100 183.290 220.270 183.460 ;
        RECT 217.600 182.790 217.770 182.960 ;
        RECT 218.100 182.790 218.270 182.960 ;
        RECT 218.600 182.790 218.770 182.960 ;
        RECT 219.100 182.790 219.270 182.960 ;
        RECT 219.600 182.790 219.770 182.960 ;
        RECT 220.100 182.790 220.270 182.960 ;
        RECT 217.600 182.290 217.770 182.460 ;
        RECT 218.100 182.290 218.270 182.460 ;
        RECT 218.600 182.290 218.770 182.460 ;
        RECT 219.100 182.290 219.270 182.460 ;
        RECT 219.600 182.290 219.770 182.460 ;
        RECT 220.100 182.290 220.270 182.460 ;
        RECT 224.300 184.790 224.470 184.960 ;
        RECT 224.800 184.790 224.970 184.960 ;
        RECT 225.300 184.790 225.470 184.960 ;
        RECT 225.800 184.790 225.970 184.960 ;
        RECT 226.300 184.790 226.470 184.960 ;
        RECT 226.800 184.790 226.970 184.960 ;
        RECT 224.300 184.290 224.470 184.460 ;
        RECT 224.800 184.290 224.970 184.460 ;
        RECT 225.300 184.290 225.470 184.460 ;
        RECT 225.800 184.290 225.970 184.460 ;
        RECT 226.300 184.290 226.470 184.460 ;
        RECT 226.800 184.290 226.970 184.460 ;
        RECT 224.300 183.790 224.470 183.960 ;
        RECT 224.800 183.790 224.970 183.960 ;
        RECT 225.300 183.790 225.470 183.960 ;
        RECT 225.800 183.790 225.970 183.960 ;
        RECT 226.300 183.790 226.470 183.960 ;
        RECT 226.800 183.790 226.970 183.960 ;
        RECT 224.300 183.290 224.470 183.460 ;
        RECT 224.800 183.290 224.970 183.460 ;
        RECT 225.300 183.290 225.470 183.460 ;
        RECT 225.800 183.290 225.970 183.460 ;
        RECT 226.300 183.290 226.470 183.460 ;
        RECT 226.800 183.290 226.970 183.460 ;
        RECT 224.300 182.790 224.470 182.960 ;
        RECT 224.800 182.790 224.970 182.960 ;
        RECT 225.300 182.790 225.470 182.960 ;
        RECT 225.800 182.790 225.970 182.960 ;
        RECT 226.300 182.790 226.470 182.960 ;
        RECT 226.800 182.790 226.970 182.960 ;
        RECT 224.300 182.290 224.470 182.460 ;
        RECT 224.800 182.290 224.970 182.460 ;
        RECT 225.300 182.290 225.470 182.460 ;
        RECT 225.800 182.290 225.970 182.460 ;
        RECT 226.300 182.290 226.470 182.460 ;
        RECT 226.800 182.290 226.970 182.460 ;
        RECT 231.000 184.790 231.170 184.960 ;
        RECT 231.500 184.790 231.670 184.960 ;
        RECT 232.000 184.790 232.170 184.960 ;
        RECT 232.500 184.790 232.670 184.960 ;
        RECT 233.000 184.790 233.170 184.960 ;
        RECT 233.500 184.790 233.670 184.960 ;
        RECT 231.000 184.290 231.170 184.460 ;
        RECT 231.500 184.290 231.670 184.460 ;
        RECT 232.000 184.290 232.170 184.460 ;
        RECT 232.500 184.290 232.670 184.460 ;
        RECT 233.000 184.290 233.170 184.460 ;
        RECT 233.500 184.290 233.670 184.460 ;
        RECT 231.000 183.790 231.170 183.960 ;
        RECT 231.500 183.790 231.670 183.960 ;
        RECT 232.000 183.790 232.170 183.960 ;
        RECT 232.500 183.790 232.670 183.960 ;
        RECT 233.000 183.790 233.170 183.960 ;
        RECT 233.500 183.790 233.670 183.960 ;
        RECT 231.000 183.290 231.170 183.460 ;
        RECT 231.500 183.290 231.670 183.460 ;
        RECT 232.000 183.290 232.170 183.460 ;
        RECT 232.500 183.290 232.670 183.460 ;
        RECT 233.000 183.290 233.170 183.460 ;
        RECT 233.500 183.290 233.670 183.460 ;
        RECT 231.000 182.790 231.170 182.960 ;
        RECT 231.500 182.790 231.670 182.960 ;
        RECT 232.000 182.790 232.170 182.960 ;
        RECT 232.500 182.790 232.670 182.960 ;
        RECT 233.000 182.790 233.170 182.960 ;
        RECT 233.500 182.790 233.670 182.960 ;
        RECT 231.000 182.290 231.170 182.460 ;
        RECT 231.500 182.290 231.670 182.460 ;
        RECT 232.000 182.290 232.170 182.460 ;
        RECT 232.500 182.290 232.670 182.460 ;
        RECT 233.000 182.290 233.170 182.460 ;
        RECT 233.500 182.290 233.670 182.460 ;
        RECT 237.700 184.790 237.870 184.960 ;
        RECT 238.200 184.790 238.370 184.960 ;
        RECT 238.700 184.790 238.870 184.960 ;
        RECT 239.200 184.790 239.370 184.960 ;
        RECT 239.700 184.790 239.870 184.960 ;
        RECT 240.200 184.790 240.370 184.960 ;
        RECT 237.700 184.290 237.870 184.460 ;
        RECT 238.200 184.290 238.370 184.460 ;
        RECT 238.700 184.290 238.870 184.460 ;
        RECT 239.200 184.290 239.370 184.460 ;
        RECT 239.700 184.290 239.870 184.460 ;
        RECT 240.200 184.290 240.370 184.460 ;
        RECT 237.700 183.790 237.870 183.960 ;
        RECT 238.200 183.790 238.370 183.960 ;
        RECT 238.700 183.790 238.870 183.960 ;
        RECT 239.200 183.790 239.370 183.960 ;
        RECT 239.700 183.790 239.870 183.960 ;
        RECT 240.200 183.790 240.370 183.960 ;
        RECT 237.700 183.290 237.870 183.460 ;
        RECT 238.200 183.290 238.370 183.460 ;
        RECT 238.700 183.290 238.870 183.460 ;
        RECT 239.200 183.290 239.370 183.460 ;
        RECT 239.700 183.290 239.870 183.460 ;
        RECT 240.200 183.290 240.370 183.460 ;
        RECT 237.700 182.790 237.870 182.960 ;
        RECT 238.200 182.790 238.370 182.960 ;
        RECT 238.700 182.790 238.870 182.960 ;
        RECT 239.200 182.790 239.370 182.960 ;
        RECT 239.700 182.790 239.870 182.960 ;
        RECT 240.200 182.790 240.370 182.960 ;
        RECT 237.700 182.290 237.870 182.460 ;
        RECT 238.200 182.290 238.370 182.460 ;
        RECT 238.700 182.290 238.870 182.460 ;
        RECT 239.200 182.290 239.370 182.460 ;
        RECT 239.700 182.290 239.870 182.460 ;
        RECT 240.200 182.290 240.370 182.460 ;
        RECT 244.400 184.790 244.570 184.960 ;
        RECT 244.900 184.790 245.070 184.960 ;
        RECT 245.400 184.790 245.570 184.960 ;
        RECT 245.900 184.790 246.070 184.960 ;
        RECT 246.400 184.790 246.570 184.960 ;
        RECT 246.900 184.790 247.070 184.960 ;
        RECT 244.400 184.290 244.570 184.460 ;
        RECT 244.900 184.290 245.070 184.460 ;
        RECT 245.400 184.290 245.570 184.460 ;
        RECT 245.900 184.290 246.070 184.460 ;
        RECT 246.400 184.290 246.570 184.460 ;
        RECT 246.900 184.290 247.070 184.460 ;
        RECT 244.400 183.790 244.570 183.960 ;
        RECT 244.900 183.790 245.070 183.960 ;
        RECT 245.400 183.790 245.570 183.960 ;
        RECT 245.900 183.790 246.070 183.960 ;
        RECT 246.400 183.790 246.570 183.960 ;
        RECT 246.900 183.790 247.070 183.960 ;
        RECT 244.400 183.290 244.570 183.460 ;
        RECT 244.900 183.290 245.070 183.460 ;
        RECT 245.400 183.290 245.570 183.460 ;
        RECT 245.900 183.290 246.070 183.460 ;
        RECT 246.400 183.290 246.570 183.460 ;
        RECT 246.900 183.290 247.070 183.460 ;
        RECT 244.400 182.790 244.570 182.960 ;
        RECT 244.900 182.790 245.070 182.960 ;
        RECT 245.400 182.790 245.570 182.960 ;
        RECT 245.900 182.790 246.070 182.960 ;
        RECT 246.400 182.790 246.570 182.960 ;
        RECT 246.900 182.790 247.070 182.960 ;
        RECT 244.400 182.290 244.570 182.460 ;
        RECT 244.900 182.290 245.070 182.460 ;
        RECT 245.400 182.290 245.570 182.460 ;
        RECT 245.900 182.290 246.070 182.460 ;
        RECT 246.400 182.290 246.570 182.460 ;
        RECT 246.900 182.290 247.070 182.460 ;
        RECT 251.100 184.790 251.270 184.960 ;
        RECT 251.600 184.790 251.770 184.960 ;
        RECT 252.100 184.790 252.270 184.960 ;
        RECT 252.600 184.790 252.770 184.960 ;
        RECT 253.100 184.790 253.270 184.960 ;
        RECT 253.600 184.790 253.770 184.960 ;
        RECT 251.100 184.290 251.270 184.460 ;
        RECT 251.600 184.290 251.770 184.460 ;
        RECT 252.100 184.290 252.270 184.460 ;
        RECT 252.600 184.290 252.770 184.460 ;
        RECT 253.100 184.290 253.270 184.460 ;
        RECT 253.600 184.290 253.770 184.460 ;
        RECT 251.100 183.790 251.270 183.960 ;
        RECT 251.600 183.790 251.770 183.960 ;
        RECT 252.100 183.790 252.270 183.960 ;
        RECT 252.600 183.790 252.770 183.960 ;
        RECT 253.100 183.790 253.270 183.960 ;
        RECT 253.600 183.790 253.770 183.960 ;
        RECT 251.100 183.290 251.270 183.460 ;
        RECT 251.600 183.290 251.770 183.460 ;
        RECT 252.100 183.290 252.270 183.460 ;
        RECT 252.600 183.290 252.770 183.460 ;
        RECT 253.100 183.290 253.270 183.460 ;
        RECT 253.600 183.290 253.770 183.460 ;
        RECT 251.100 182.790 251.270 182.960 ;
        RECT 251.600 182.790 251.770 182.960 ;
        RECT 252.100 182.790 252.270 182.960 ;
        RECT 252.600 182.790 252.770 182.960 ;
        RECT 253.100 182.790 253.270 182.960 ;
        RECT 253.600 182.790 253.770 182.960 ;
        RECT 251.100 182.290 251.270 182.460 ;
        RECT 251.600 182.290 251.770 182.460 ;
        RECT 252.100 182.290 252.270 182.460 ;
        RECT 252.600 182.290 252.770 182.460 ;
        RECT 253.100 182.290 253.270 182.460 ;
        RECT 253.600 182.290 253.770 182.460 ;
        RECT 257.800 184.790 257.970 184.960 ;
        RECT 258.300 184.790 258.470 184.960 ;
        RECT 258.800 184.790 258.970 184.960 ;
        RECT 259.300 184.790 259.470 184.960 ;
        RECT 259.800 184.790 259.970 184.960 ;
        RECT 260.300 184.790 260.470 184.960 ;
        RECT 257.800 184.290 257.970 184.460 ;
        RECT 258.300 184.290 258.470 184.460 ;
        RECT 258.800 184.290 258.970 184.460 ;
        RECT 259.300 184.290 259.470 184.460 ;
        RECT 259.800 184.290 259.970 184.460 ;
        RECT 260.300 184.290 260.470 184.460 ;
        RECT 257.800 183.790 257.970 183.960 ;
        RECT 258.300 183.790 258.470 183.960 ;
        RECT 258.800 183.790 258.970 183.960 ;
        RECT 259.300 183.790 259.470 183.960 ;
        RECT 259.800 183.790 259.970 183.960 ;
        RECT 260.300 183.790 260.470 183.960 ;
        RECT 257.800 183.290 257.970 183.460 ;
        RECT 258.300 183.290 258.470 183.460 ;
        RECT 258.800 183.290 258.970 183.460 ;
        RECT 259.300 183.290 259.470 183.460 ;
        RECT 259.800 183.290 259.970 183.460 ;
        RECT 260.300 183.290 260.470 183.460 ;
        RECT 257.800 182.790 257.970 182.960 ;
        RECT 258.300 182.790 258.470 182.960 ;
        RECT 258.800 182.790 258.970 182.960 ;
        RECT 259.300 182.790 259.470 182.960 ;
        RECT 259.800 182.790 259.970 182.960 ;
        RECT 260.300 182.790 260.470 182.960 ;
        RECT 257.800 182.290 257.970 182.460 ;
        RECT 258.300 182.290 258.470 182.460 ;
        RECT 258.800 182.290 258.970 182.460 ;
        RECT 259.300 182.290 259.470 182.460 ;
        RECT 259.800 182.290 259.970 182.460 ;
        RECT 260.300 182.290 260.470 182.460 ;
        RECT 201.335 181.535 201.505 181.705 ;
        RECT 201.335 181.175 201.505 181.345 ;
        RECT 201.335 180.815 201.505 180.985 ;
        RECT 187.825 180.115 187.995 180.285 ;
        RECT 192.885 179.605 193.055 179.775 ;
        RECT 96.415 165.615 98.385 168.305 ;
        RECT 106.450 165.615 108.420 168.305 ;
        RECT 96.415 160.815 98.385 163.505 ;
        RECT 110.140 165.615 112.110 168.305 ;
        RECT 123.045 165.615 125.015 168.305 ;
        RECT 106.450 160.815 108.420 163.505 ;
        RECT 123.045 160.815 125.015 163.505 ;
        RECT 210.900 165.990 211.070 166.160 ;
        RECT 211.400 165.990 211.570 166.160 ;
        RECT 211.900 165.990 212.070 166.160 ;
        RECT 212.400 165.990 212.570 166.160 ;
        RECT 212.900 165.990 213.070 166.160 ;
        RECT 213.400 165.990 213.570 166.160 ;
        RECT 210.900 165.490 211.070 165.660 ;
        RECT 211.400 165.490 211.570 165.660 ;
        RECT 211.900 165.490 212.070 165.660 ;
        RECT 212.400 165.490 212.570 165.660 ;
        RECT 212.900 165.490 213.070 165.660 ;
        RECT 213.400 165.490 213.570 165.660 ;
        RECT 210.900 164.990 211.070 165.160 ;
        RECT 211.400 164.990 211.570 165.160 ;
        RECT 211.900 164.990 212.070 165.160 ;
        RECT 212.400 164.990 212.570 165.160 ;
        RECT 212.900 164.990 213.070 165.160 ;
        RECT 213.400 164.990 213.570 165.160 ;
        RECT 210.900 164.490 211.070 164.660 ;
        RECT 211.400 164.490 211.570 164.660 ;
        RECT 211.900 164.490 212.070 164.660 ;
        RECT 212.400 164.490 212.570 164.660 ;
        RECT 212.900 164.490 213.070 164.660 ;
        RECT 213.400 164.490 213.570 164.660 ;
        RECT 210.900 163.990 211.070 164.160 ;
        RECT 211.400 163.990 211.570 164.160 ;
        RECT 211.900 163.990 212.070 164.160 ;
        RECT 212.400 163.990 212.570 164.160 ;
        RECT 212.900 163.990 213.070 164.160 ;
        RECT 213.400 163.990 213.570 164.160 ;
        RECT 210.900 163.490 211.070 163.660 ;
        RECT 211.400 163.490 211.570 163.660 ;
        RECT 211.900 163.490 212.070 163.660 ;
        RECT 212.400 163.490 212.570 163.660 ;
        RECT 212.900 163.490 213.070 163.660 ;
        RECT 213.400 163.490 213.570 163.660 ;
        RECT 217.600 165.990 217.770 166.160 ;
        RECT 218.100 165.990 218.270 166.160 ;
        RECT 218.600 165.990 218.770 166.160 ;
        RECT 219.100 165.990 219.270 166.160 ;
        RECT 219.600 165.990 219.770 166.160 ;
        RECT 220.100 165.990 220.270 166.160 ;
        RECT 217.600 165.490 217.770 165.660 ;
        RECT 218.100 165.490 218.270 165.660 ;
        RECT 218.600 165.490 218.770 165.660 ;
        RECT 219.100 165.490 219.270 165.660 ;
        RECT 219.600 165.490 219.770 165.660 ;
        RECT 220.100 165.490 220.270 165.660 ;
        RECT 217.600 164.990 217.770 165.160 ;
        RECT 218.100 164.990 218.270 165.160 ;
        RECT 218.600 164.990 218.770 165.160 ;
        RECT 219.100 164.990 219.270 165.160 ;
        RECT 219.600 164.990 219.770 165.160 ;
        RECT 220.100 164.990 220.270 165.160 ;
        RECT 217.600 164.490 217.770 164.660 ;
        RECT 218.100 164.490 218.270 164.660 ;
        RECT 218.600 164.490 218.770 164.660 ;
        RECT 219.100 164.490 219.270 164.660 ;
        RECT 219.600 164.490 219.770 164.660 ;
        RECT 220.100 164.490 220.270 164.660 ;
        RECT 217.600 163.990 217.770 164.160 ;
        RECT 218.100 163.990 218.270 164.160 ;
        RECT 218.600 163.990 218.770 164.160 ;
        RECT 219.100 163.990 219.270 164.160 ;
        RECT 219.600 163.990 219.770 164.160 ;
        RECT 220.100 163.990 220.270 164.160 ;
        RECT 217.600 163.490 217.770 163.660 ;
        RECT 218.100 163.490 218.270 163.660 ;
        RECT 218.600 163.490 218.770 163.660 ;
        RECT 219.100 163.490 219.270 163.660 ;
        RECT 219.600 163.490 219.770 163.660 ;
        RECT 220.100 163.490 220.270 163.660 ;
        RECT 224.300 165.990 224.470 166.160 ;
        RECT 224.800 165.990 224.970 166.160 ;
        RECT 225.300 165.990 225.470 166.160 ;
        RECT 225.800 165.990 225.970 166.160 ;
        RECT 226.300 165.990 226.470 166.160 ;
        RECT 226.800 165.990 226.970 166.160 ;
        RECT 224.300 165.490 224.470 165.660 ;
        RECT 224.800 165.490 224.970 165.660 ;
        RECT 225.300 165.490 225.470 165.660 ;
        RECT 225.800 165.490 225.970 165.660 ;
        RECT 226.300 165.490 226.470 165.660 ;
        RECT 226.800 165.490 226.970 165.660 ;
        RECT 224.300 164.990 224.470 165.160 ;
        RECT 224.800 164.990 224.970 165.160 ;
        RECT 225.300 164.990 225.470 165.160 ;
        RECT 225.800 164.990 225.970 165.160 ;
        RECT 226.300 164.990 226.470 165.160 ;
        RECT 226.800 164.990 226.970 165.160 ;
        RECT 224.300 164.490 224.470 164.660 ;
        RECT 224.800 164.490 224.970 164.660 ;
        RECT 225.300 164.490 225.470 164.660 ;
        RECT 225.800 164.490 225.970 164.660 ;
        RECT 226.300 164.490 226.470 164.660 ;
        RECT 226.800 164.490 226.970 164.660 ;
        RECT 224.300 163.990 224.470 164.160 ;
        RECT 224.800 163.990 224.970 164.160 ;
        RECT 225.300 163.990 225.470 164.160 ;
        RECT 225.800 163.990 225.970 164.160 ;
        RECT 226.300 163.990 226.470 164.160 ;
        RECT 226.800 163.990 226.970 164.160 ;
        RECT 224.300 163.490 224.470 163.660 ;
        RECT 224.800 163.490 224.970 163.660 ;
        RECT 225.300 163.490 225.470 163.660 ;
        RECT 225.800 163.490 225.970 163.660 ;
        RECT 226.300 163.490 226.470 163.660 ;
        RECT 226.800 163.490 226.970 163.660 ;
        RECT 231.000 165.990 231.170 166.160 ;
        RECT 231.500 165.990 231.670 166.160 ;
        RECT 232.000 165.990 232.170 166.160 ;
        RECT 232.500 165.990 232.670 166.160 ;
        RECT 233.000 165.990 233.170 166.160 ;
        RECT 233.500 165.990 233.670 166.160 ;
        RECT 231.000 165.490 231.170 165.660 ;
        RECT 231.500 165.490 231.670 165.660 ;
        RECT 232.000 165.490 232.170 165.660 ;
        RECT 232.500 165.490 232.670 165.660 ;
        RECT 233.000 165.490 233.170 165.660 ;
        RECT 233.500 165.490 233.670 165.660 ;
        RECT 231.000 164.990 231.170 165.160 ;
        RECT 231.500 164.990 231.670 165.160 ;
        RECT 232.000 164.990 232.170 165.160 ;
        RECT 232.500 164.990 232.670 165.160 ;
        RECT 233.000 164.990 233.170 165.160 ;
        RECT 233.500 164.990 233.670 165.160 ;
        RECT 231.000 164.490 231.170 164.660 ;
        RECT 231.500 164.490 231.670 164.660 ;
        RECT 232.000 164.490 232.170 164.660 ;
        RECT 232.500 164.490 232.670 164.660 ;
        RECT 233.000 164.490 233.170 164.660 ;
        RECT 233.500 164.490 233.670 164.660 ;
        RECT 231.000 163.990 231.170 164.160 ;
        RECT 231.500 163.990 231.670 164.160 ;
        RECT 232.000 163.990 232.170 164.160 ;
        RECT 232.500 163.990 232.670 164.160 ;
        RECT 233.000 163.990 233.170 164.160 ;
        RECT 233.500 163.990 233.670 164.160 ;
        RECT 231.000 163.490 231.170 163.660 ;
        RECT 231.500 163.490 231.670 163.660 ;
        RECT 232.000 163.490 232.170 163.660 ;
        RECT 232.500 163.490 232.670 163.660 ;
        RECT 233.000 163.490 233.170 163.660 ;
        RECT 233.500 163.490 233.670 163.660 ;
        RECT 237.700 165.990 237.870 166.160 ;
        RECT 238.200 165.990 238.370 166.160 ;
        RECT 238.700 165.990 238.870 166.160 ;
        RECT 239.200 165.990 239.370 166.160 ;
        RECT 239.700 165.990 239.870 166.160 ;
        RECT 240.200 165.990 240.370 166.160 ;
        RECT 237.700 165.490 237.870 165.660 ;
        RECT 238.200 165.490 238.370 165.660 ;
        RECT 238.700 165.490 238.870 165.660 ;
        RECT 239.200 165.490 239.370 165.660 ;
        RECT 239.700 165.490 239.870 165.660 ;
        RECT 240.200 165.490 240.370 165.660 ;
        RECT 237.700 164.990 237.870 165.160 ;
        RECT 238.200 164.990 238.370 165.160 ;
        RECT 238.700 164.990 238.870 165.160 ;
        RECT 239.200 164.990 239.370 165.160 ;
        RECT 239.700 164.990 239.870 165.160 ;
        RECT 240.200 164.990 240.370 165.160 ;
        RECT 237.700 164.490 237.870 164.660 ;
        RECT 238.200 164.490 238.370 164.660 ;
        RECT 238.700 164.490 238.870 164.660 ;
        RECT 239.200 164.490 239.370 164.660 ;
        RECT 239.700 164.490 239.870 164.660 ;
        RECT 240.200 164.490 240.370 164.660 ;
        RECT 237.700 163.990 237.870 164.160 ;
        RECT 238.200 163.990 238.370 164.160 ;
        RECT 238.700 163.990 238.870 164.160 ;
        RECT 239.200 163.990 239.370 164.160 ;
        RECT 239.700 163.990 239.870 164.160 ;
        RECT 240.200 163.990 240.370 164.160 ;
        RECT 237.700 163.490 237.870 163.660 ;
        RECT 238.200 163.490 238.370 163.660 ;
        RECT 238.700 163.490 238.870 163.660 ;
        RECT 239.200 163.490 239.370 163.660 ;
        RECT 239.700 163.490 239.870 163.660 ;
        RECT 240.200 163.490 240.370 163.660 ;
        RECT 244.400 165.990 244.570 166.160 ;
        RECT 244.900 165.990 245.070 166.160 ;
        RECT 245.400 165.990 245.570 166.160 ;
        RECT 245.900 165.990 246.070 166.160 ;
        RECT 246.400 165.990 246.570 166.160 ;
        RECT 246.900 165.990 247.070 166.160 ;
        RECT 244.400 165.490 244.570 165.660 ;
        RECT 244.900 165.490 245.070 165.660 ;
        RECT 245.400 165.490 245.570 165.660 ;
        RECT 245.900 165.490 246.070 165.660 ;
        RECT 246.400 165.490 246.570 165.660 ;
        RECT 246.900 165.490 247.070 165.660 ;
        RECT 244.400 164.990 244.570 165.160 ;
        RECT 244.900 164.990 245.070 165.160 ;
        RECT 245.400 164.990 245.570 165.160 ;
        RECT 245.900 164.990 246.070 165.160 ;
        RECT 246.400 164.990 246.570 165.160 ;
        RECT 246.900 164.990 247.070 165.160 ;
        RECT 244.400 164.490 244.570 164.660 ;
        RECT 244.900 164.490 245.070 164.660 ;
        RECT 245.400 164.490 245.570 164.660 ;
        RECT 245.900 164.490 246.070 164.660 ;
        RECT 246.400 164.490 246.570 164.660 ;
        RECT 246.900 164.490 247.070 164.660 ;
        RECT 244.400 163.990 244.570 164.160 ;
        RECT 244.900 163.990 245.070 164.160 ;
        RECT 245.400 163.990 245.570 164.160 ;
        RECT 245.900 163.990 246.070 164.160 ;
        RECT 246.400 163.990 246.570 164.160 ;
        RECT 246.900 163.990 247.070 164.160 ;
        RECT 244.400 163.490 244.570 163.660 ;
        RECT 244.900 163.490 245.070 163.660 ;
        RECT 245.400 163.490 245.570 163.660 ;
        RECT 245.900 163.490 246.070 163.660 ;
        RECT 246.400 163.490 246.570 163.660 ;
        RECT 246.900 163.490 247.070 163.660 ;
        RECT 251.100 165.990 251.270 166.160 ;
        RECT 251.600 165.990 251.770 166.160 ;
        RECT 252.100 165.990 252.270 166.160 ;
        RECT 252.600 165.990 252.770 166.160 ;
        RECT 253.100 165.990 253.270 166.160 ;
        RECT 253.600 165.990 253.770 166.160 ;
        RECT 251.100 165.490 251.270 165.660 ;
        RECT 251.600 165.490 251.770 165.660 ;
        RECT 252.100 165.490 252.270 165.660 ;
        RECT 252.600 165.490 252.770 165.660 ;
        RECT 253.100 165.490 253.270 165.660 ;
        RECT 253.600 165.490 253.770 165.660 ;
        RECT 251.100 164.990 251.270 165.160 ;
        RECT 251.600 164.990 251.770 165.160 ;
        RECT 252.100 164.990 252.270 165.160 ;
        RECT 252.600 164.990 252.770 165.160 ;
        RECT 253.100 164.990 253.270 165.160 ;
        RECT 253.600 164.990 253.770 165.160 ;
        RECT 251.100 164.490 251.270 164.660 ;
        RECT 251.600 164.490 251.770 164.660 ;
        RECT 252.100 164.490 252.270 164.660 ;
        RECT 252.600 164.490 252.770 164.660 ;
        RECT 253.100 164.490 253.270 164.660 ;
        RECT 253.600 164.490 253.770 164.660 ;
        RECT 251.100 163.990 251.270 164.160 ;
        RECT 251.600 163.990 251.770 164.160 ;
        RECT 252.100 163.990 252.270 164.160 ;
        RECT 252.600 163.990 252.770 164.160 ;
        RECT 253.100 163.990 253.270 164.160 ;
        RECT 253.600 163.990 253.770 164.160 ;
        RECT 251.100 163.490 251.270 163.660 ;
        RECT 251.600 163.490 251.770 163.660 ;
        RECT 252.100 163.490 252.270 163.660 ;
        RECT 252.600 163.490 252.770 163.660 ;
        RECT 253.100 163.490 253.270 163.660 ;
        RECT 253.600 163.490 253.770 163.660 ;
        RECT 257.800 165.990 257.970 166.160 ;
        RECT 258.300 165.990 258.470 166.160 ;
        RECT 258.800 165.990 258.970 166.160 ;
        RECT 259.300 165.990 259.470 166.160 ;
        RECT 259.800 165.990 259.970 166.160 ;
        RECT 260.300 165.990 260.470 166.160 ;
        RECT 257.800 165.490 257.970 165.660 ;
        RECT 258.300 165.490 258.470 165.660 ;
        RECT 258.800 165.490 258.970 165.660 ;
        RECT 259.300 165.490 259.470 165.660 ;
        RECT 259.800 165.490 259.970 165.660 ;
        RECT 260.300 165.490 260.470 165.660 ;
        RECT 257.800 164.990 257.970 165.160 ;
        RECT 258.300 164.990 258.470 165.160 ;
        RECT 258.800 164.990 258.970 165.160 ;
        RECT 259.300 164.990 259.470 165.160 ;
        RECT 259.800 164.990 259.970 165.160 ;
        RECT 260.300 164.990 260.470 165.160 ;
        RECT 257.800 164.490 257.970 164.660 ;
        RECT 258.300 164.490 258.470 164.660 ;
        RECT 258.800 164.490 258.970 164.660 ;
        RECT 259.300 164.490 259.470 164.660 ;
        RECT 259.800 164.490 259.970 164.660 ;
        RECT 260.300 164.490 260.470 164.660 ;
        RECT 257.800 163.990 257.970 164.160 ;
        RECT 258.300 163.990 258.470 164.160 ;
        RECT 258.800 163.990 258.970 164.160 ;
        RECT 259.300 163.990 259.470 164.160 ;
        RECT 259.800 163.990 259.970 164.160 ;
        RECT 260.300 163.990 260.470 164.160 ;
        RECT 257.800 163.490 257.970 163.660 ;
        RECT 258.300 163.490 258.470 163.660 ;
        RECT 258.800 163.490 258.970 163.660 ;
        RECT 259.300 163.490 259.470 163.660 ;
        RECT 259.800 163.490 259.970 163.660 ;
        RECT 260.300 163.490 260.470 163.660 ;
        RECT 82.695 146.815 84.665 149.505 ;
        RECT 92.730 146.815 94.700 149.505 ;
        RECT 82.695 142.015 84.665 144.705 ;
        RECT 96.415 146.815 98.385 149.505 ;
        RECT 106.450 146.815 108.420 149.505 ;
        RECT 92.730 142.015 94.700 144.705 ;
        RECT 96.415 142.015 98.385 144.705 ;
        RECT 120.170 146.815 122.140 149.505 ;
        RECT 106.450 142.015 108.420 144.705 ;
        RECT 110.135 142.015 112.105 144.705 ;
        RECT 136.105 146.815 138.075 149.505 ;
        RECT 146.140 146.815 148.110 149.505 ;
        RECT 120.170 142.015 122.140 144.705 ;
        RECT 136.105 142.015 138.075 144.705 ;
        RECT 146.140 142.015 148.110 144.705 ;
        RECT 187.595 149.335 187.765 149.505 ;
        RECT 187.595 148.975 187.765 149.145 ;
        RECT 187.595 148.615 187.765 148.785 ;
        RECT 187.595 148.255 187.765 148.425 ;
        RECT 187.595 147.895 187.765 148.065 ;
        RECT 187.595 147.535 187.765 147.705 ;
        RECT 187.595 147.175 187.765 147.345 ;
        RECT 187.595 146.815 187.765 146.985 ;
        RECT 187.595 146.455 187.765 146.625 ;
        RECT 187.595 146.095 187.765 146.265 ;
        RECT 187.595 145.735 187.765 145.905 ;
        RECT 187.595 145.375 187.765 145.545 ;
        RECT 187.595 145.015 187.765 145.185 ;
        RECT 187.595 144.655 187.765 144.825 ;
        RECT 187.595 144.295 187.765 144.465 ;
        RECT 187.595 143.935 187.765 144.105 ;
        RECT 187.595 143.575 187.765 143.745 ;
        RECT 187.595 143.215 187.765 143.385 ;
        RECT 192.175 149.335 192.345 149.505 ;
        RECT 192.175 148.975 192.345 149.145 ;
        RECT 192.175 148.615 192.345 148.785 ;
        RECT 192.175 148.255 192.345 148.425 ;
        RECT 192.175 147.895 192.345 148.065 ;
        RECT 192.175 147.535 192.345 147.705 ;
        RECT 192.175 147.175 192.345 147.345 ;
        RECT 192.175 146.815 192.345 146.985 ;
        RECT 192.175 146.455 192.345 146.625 ;
        RECT 192.175 146.095 192.345 146.265 ;
        RECT 192.175 145.735 192.345 145.905 ;
        RECT 192.175 145.375 192.345 145.545 ;
        RECT 192.175 145.015 192.345 145.185 ;
        RECT 192.175 144.655 192.345 144.825 ;
        RECT 192.175 144.295 192.345 144.465 ;
        RECT 192.175 143.935 192.345 144.105 ;
        RECT 192.175 143.575 192.345 143.745 ;
        RECT 192.175 143.215 192.345 143.385 ;
        RECT 196.755 149.335 196.925 149.505 ;
        RECT 196.755 148.975 196.925 149.145 ;
        RECT 196.755 148.615 196.925 148.785 ;
        RECT 196.755 148.255 196.925 148.425 ;
        RECT 196.755 147.895 196.925 148.065 ;
        RECT 196.755 147.535 196.925 147.705 ;
        RECT 196.755 147.175 196.925 147.345 ;
        RECT 196.755 146.815 196.925 146.985 ;
        RECT 196.755 146.455 196.925 146.625 ;
        RECT 196.755 146.095 196.925 146.265 ;
        RECT 196.755 145.735 196.925 145.905 ;
        RECT 196.755 145.375 196.925 145.545 ;
        RECT 196.755 145.015 196.925 145.185 ;
        RECT 196.755 144.655 196.925 144.825 ;
        RECT 196.755 144.295 196.925 144.465 ;
        RECT 196.755 143.935 196.925 144.105 ;
        RECT 196.755 143.575 196.925 143.745 ;
        RECT 196.755 143.215 196.925 143.385 ;
        RECT 192.885 142.545 193.055 142.715 ;
        RECT 201.335 149.335 201.505 149.505 ;
        RECT 201.335 148.975 201.505 149.145 ;
        RECT 201.335 148.615 201.505 148.785 ;
        RECT 201.335 148.255 201.505 148.425 ;
        RECT 201.335 147.895 201.505 148.065 ;
        RECT 201.335 147.535 201.505 147.705 ;
        RECT 201.335 147.175 201.505 147.345 ;
        RECT 201.335 146.815 201.505 146.985 ;
        RECT 201.335 146.455 201.505 146.625 ;
        RECT 201.335 146.095 201.505 146.265 ;
        RECT 201.335 145.735 201.505 145.905 ;
        RECT 201.335 145.375 201.505 145.545 ;
        RECT 201.335 145.015 201.505 145.185 ;
        RECT 201.335 144.655 201.505 144.825 ;
        RECT 201.335 144.295 201.505 144.465 ;
        RECT 210.900 147.190 211.070 147.360 ;
        RECT 211.400 147.190 211.570 147.360 ;
        RECT 211.900 147.190 212.070 147.360 ;
        RECT 212.400 147.190 212.570 147.360 ;
        RECT 212.900 147.190 213.070 147.360 ;
        RECT 213.400 147.190 213.570 147.360 ;
        RECT 210.900 146.690 211.070 146.860 ;
        RECT 211.400 146.690 211.570 146.860 ;
        RECT 211.900 146.690 212.070 146.860 ;
        RECT 212.400 146.690 212.570 146.860 ;
        RECT 212.900 146.690 213.070 146.860 ;
        RECT 213.400 146.690 213.570 146.860 ;
        RECT 210.900 146.190 211.070 146.360 ;
        RECT 211.400 146.190 211.570 146.360 ;
        RECT 211.900 146.190 212.070 146.360 ;
        RECT 212.400 146.190 212.570 146.360 ;
        RECT 212.900 146.190 213.070 146.360 ;
        RECT 213.400 146.190 213.570 146.360 ;
        RECT 210.900 145.690 211.070 145.860 ;
        RECT 211.400 145.690 211.570 145.860 ;
        RECT 211.900 145.690 212.070 145.860 ;
        RECT 212.400 145.690 212.570 145.860 ;
        RECT 212.900 145.690 213.070 145.860 ;
        RECT 213.400 145.690 213.570 145.860 ;
        RECT 210.900 145.190 211.070 145.360 ;
        RECT 211.400 145.190 211.570 145.360 ;
        RECT 211.900 145.190 212.070 145.360 ;
        RECT 212.400 145.190 212.570 145.360 ;
        RECT 212.900 145.190 213.070 145.360 ;
        RECT 213.400 145.190 213.570 145.360 ;
        RECT 210.900 144.690 211.070 144.860 ;
        RECT 211.400 144.690 211.570 144.860 ;
        RECT 211.900 144.690 212.070 144.860 ;
        RECT 212.400 144.690 212.570 144.860 ;
        RECT 212.900 144.690 213.070 144.860 ;
        RECT 213.400 144.690 213.570 144.860 ;
        RECT 217.600 147.190 217.770 147.360 ;
        RECT 218.100 147.190 218.270 147.360 ;
        RECT 218.600 147.190 218.770 147.360 ;
        RECT 219.100 147.190 219.270 147.360 ;
        RECT 219.600 147.190 219.770 147.360 ;
        RECT 220.100 147.190 220.270 147.360 ;
        RECT 217.600 146.690 217.770 146.860 ;
        RECT 218.100 146.690 218.270 146.860 ;
        RECT 218.600 146.690 218.770 146.860 ;
        RECT 219.100 146.690 219.270 146.860 ;
        RECT 219.600 146.690 219.770 146.860 ;
        RECT 220.100 146.690 220.270 146.860 ;
        RECT 217.600 146.190 217.770 146.360 ;
        RECT 218.100 146.190 218.270 146.360 ;
        RECT 218.600 146.190 218.770 146.360 ;
        RECT 219.100 146.190 219.270 146.360 ;
        RECT 219.600 146.190 219.770 146.360 ;
        RECT 220.100 146.190 220.270 146.360 ;
        RECT 217.600 145.690 217.770 145.860 ;
        RECT 218.100 145.690 218.270 145.860 ;
        RECT 218.600 145.690 218.770 145.860 ;
        RECT 219.100 145.690 219.270 145.860 ;
        RECT 219.600 145.690 219.770 145.860 ;
        RECT 220.100 145.690 220.270 145.860 ;
        RECT 217.600 145.190 217.770 145.360 ;
        RECT 218.100 145.190 218.270 145.360 ;
        RECT 218.600 145.190 218.770 145.360 ;
        RECT 219.100 145.190 219.270 145.360 ;
        RECT 219.600 145.190 219.770 145.360 ;
        RECT 220.100 145.190 220.270 145.360 ;
        RECT 217.600 144.690 217.770 144.860 ;
        RECT 218.100 144.690 218.270 144.860 ;
        RECT 218.600 144.690 218.770 144.860 ;
        RECT 219.100 144.690 219.270 144.860 ;
        RECT 219.600 144.690 219.770 144.860 ;
        RECT 220.100 144.690 220.270 144.860 ;
        RECT 224.300 147.190 224.470 147.360 ;
        RECT 224.800 147.190 224.970 147.360 ;
        RECT 225.300 147.190 225.470 147.360 ;
        RECT 225.800 147.190 225.970 147.360 ;
        RECT 226.300 147.190 226.470 147.360 ;
        RECT 226.800 147.190 226.970 147.360 ;
        RECT 224.300 146.690 224.470 146.860 ;
        RECT 224.800 146.690 224.970 146.860 ;
        RECT 225.300 146.690 225.470 146.860 ;
        RECT 225.800 146.690 225.970 146.860 ;
        RECT 226.300 146.690 226.470 146.860 ;
        RECT 226.800 146.690 226.970 146.860 ;
        RECT 224.300 146.190 224.470 146.360 ;
        RECT 224.800 146.190 224.970 146.360 ;
        RECT 225.300 146.190 225.470 146.360 ;
        RECT 225.800 146.190 225.970 146.360 ;
        RECT 226.300 146.190 226.470 146.360 ;
        RECT 226.800 146.190 226.970 146.360 ;
        RECT 224.300 145.690 224.470 145.860 ;
        RECT 224.800 145.690 224.970 145.860 ;
        RECT 225.300 145.690 225.470 145.860 ;
        RECT 225.800 145.690 225.970 145.860 ;
        RECT 226.300 145.690 226.470 145.860 ;
        RECT 226.800 145.690 226.970 145.860 ;
        RECT 224.300 145.190 224.470 145.360 ;
        RECT 224.800 145.190 224.970 145.360 ;
        RECT 225.300 145.190 225.470 145.360 ;
        RECT 225.800 145.190 225.970 145.360 ;
        RECT 226.300 145.190 226.470 145.360 ;
        RECT 226.800 145.190 226.970 145.360 ;
        RECT 224.300 144.690 224.470 144.860 ;
        RECT 224.800 144.690 224.970 144.860 ;
        RECT 225.300 144.690 225.470 144.860 ;
        RECT 225.800 144.690 225.970 144.860 ;
        RECT 226.300 144.690 226.470 144.860 ;
        RECT 226.800 144.690 226.970 144.860 ;
        RECT 231.000 147.190 231.170 147.360 ;
        RECT 231.500 147.190 231.670 147.360 ;
        RECT 232.000 147.190 232.170 147.360 ;
        RECT 232.500 147.190 232.670 147.360 ;
        RECT 233.000 147.190 233.170 147.360 ;
        RECT 233.500 147.190 233.670 147.360 ;
        RECT 231.000 146.690 231.170 146.860 ;
        RECT 231.500 146.690 231.670 146.860 ;
        RECT 232.000 146.690 232.170 146.860 ;
        RECT 232.500 146.690 232.670 146.860 ;
        RECT 233.000 146.690 233.170 146.860 ;
        RECT 233.500 146.690 233.670 146.860 ;
        RECT 231.000 146.190 231.170 146.360 ;
        RECT 231.500 146.190 231.670 146.360 ;
        RECT 232.000 146.190 232.170 146.360 ;
        RECT 232.500 146.190 232.670 146.360 ;
        RECT 233.000 146.190 233.170 146.360 ;
        RECT 233.500 146.190 233.670 146.360 ;
        RECT 231.000 145.690 231.170 145.860 ;
        RECT 231.500 145.690 231.670 145.860 ;
        RECT 232.000 145.690 232.170 145.860 ;
        RECT 232.500 145.690 232.670 145.860 ;
        RECT 233.000 145.690 233.170 145.860 ;
        RECT 233.500 145.690 233.670 145.860 ;
        RECT 231.000 145.190 231.170 145.360 ;
        RECT 231.500 145.190 231.670 145.360 ;
        RECT 232.000 145.190 232.170 145.360 ;
        RECT 232.500 145.190 232.670 145.360 ;
        RECT 233.000 145.190 233.170 145.360 ;
        RECT 233.500 145.190 233.670 145.360 ;
        RECT 231.000 144.690 231.170 144.860 ;
        RECT 231.500 144.690 231.670 144.860 ;
        RECT 232.000 144.690 232.170 144.860 ;
        RECT 232.500 144.690 232.670 144.860 ;
        RECT 233.000 144.690 233.170 144.860 ;
        RECT 233.500 144.690 233.670 144.860 ;
        RECT 237.700 147.190 237.870 147.360 ;
        RECT 238.200 147.190 238.370 147.360 ;
        RECT 238.700 147.190 238.870 147.360 ;
        RECT 239.200 147.190 239.370 147.360 ;
        RECT 239.700 147.190 239.870 147.360 ;
        RECT 240.200 147.190 240.370 147.360 ;
        RECT 237.700 146.690 237.870 146.860 ;
        RECT 238.200 146.690 238.370 146.860 ;
        RECT 238.700 146.690 238.870 146.860 ;
        RECT 239.200 146.690 239.370 146.860 ;
        RECT 239.700 146.690 239.870 146.860 ;
        RECT 240.200 146.690 240.370 146.860 ;
        RECT 237.700 146.190 237.870 146.360 ;
        RECT 238.200 146.190 238.370 146.360 ;
        RECT 238.700 146.190 238.870 146.360 ;
        RECT 239.200 146.190 239.370 146.360 ;
        RECT 239.700 146.190 239.870 146.360 ;
        RECT 240.200 146.190 240.370 146.360 ;
        RECT 237.700 145.690 237.870 145.860 ;
        RECT 238.200 145.690 238.370 145.860 ;
        RECT 238.700 145.690 238.870 145.860 ;
        RECT 239.200 145.690 239.370 145.860 ;
        RECT 239.700 145.690 239.870 145.860 ;
        RECT 240.200 145.690 240.370 145.860 ;
        RECT 237.700 145.190 237.870 145.360 ;
        RECT 238.200 145.190 238.370 145.360 ;
        RECT 238.700 145.190 238.870 145.360 ;
        RECT 239.200 145.190 239.370 145.360 ;
        RECT 239.700 145.190 239.870 145.360 ;
        RECT 240.200 145.190 240.370 145.360 ;
        RECT 237.700 144.690 237.870 144.860 ;
        RECT 238.200 144.690 238.370 144.860 ;
        RECT 238.700 144.690 238.870 144.860 ;
        RECT 239.200 144.690 239.370 144.860 ;
        RECT 239.700 144.690 239.870 144.860 ;
        RECT 240.200 144.690 240.370 144.860 ;
        RECT 244.400 147.190 244.570 147.360 ;
        RECT 244.900 147.190 245.070 147.360 ;
        RECT 245.400 147.190 245.570 147.360 ;
        RECT 245.900 147.190 246.070 147.360 ;
        RECT 246.400 147.190 246.570 147.360 ;
        RECT 246.900 147.190 247.070 147.360 ;
        RECT 244.400 146.690 244.570 146.860 ;
        RECT 244.900 146.690 245.070 146.860 ;
        RECT 245.400 146.690 245.570 146.860 ;
        RECT 245.900 146.690 246.070 146.860 ;
        RECT 246.400 146.690 246.570 146.860 ;
        RECT 246.900 146.690 247.070 146.860 ;
        RECT 244.400 146.190 244.570 146.360 ;
        RECT 244.900 146.190 245.070 146.360 ;
        RECT 245.400 146.190 245.570 146.360 ;
        RECT 245.900 146.190 246.070 146.360 ;
        RECT 246.400 146.190 246.570 146.360 ;
        RECT 246.900 146.190 247.070 146.360 ;
        RECT 244.400 145.690 244.570 145.860 ;
        RECT 244.900 145.690 245.070 145.860 ;
        RECT 245.400 145.690 245.570 145.860 ;
        RECT 245.900 145.690 246.070 145.860 ;
        RECT 246.400 145.690 246.570 145.860 ;
        RECT 246.900 145.690 247.070 145.860 ;
        RECT 244.400 145.190 244.570 145.360 ;
        RECT 244.900 145.190 245.070 145.360 ;
        RECT 245.400 145.190 245.570 145.360 ;
        RECT 245.900 145.190 246.070 145.360 ;
        RECT 246.400 145.190 246.570 145.360 ;
        RECT 246.900 145.190 247.070 145.360 ;
        RECT 244.400 144.690 244.570 144.860 ;
        RECT 244.900 144.690 245.070 144.860 ;
        RECT 245.400 144.690 245.570 144.860 ;
        RECT 245.900 144.690 246.070 144.860 ;
        RECT 246.400 144.690 246.570 144.860 ;
        RECT 246.900 144.690 247.070 144.860 ;
        RECT 251.100 147.190 251.270 147.360 ;
        RECT 251.600 147.190 251.770 147.360 ;
        RECT 252.100 147.190 252.270 147.360 ;
        RECT 252.600 147.190 252.770 147.360 ;
        RECT 253.100 147.190 253.270 147.360 ;
        RECT 253.600 147.190 253.770 147.360 ;
        RECT 251.100 146.690 251.270 146.860 ;
        RECT 251.600 146.690 251.770 146.860 ;
        RECT 252.100 146.690 252.270 146.860 ;
        RECT 252.600 146.690 252.770 146.860 ;
        RECT 253.100 146.690 253.270 146.860 ;
        RECT 253.600 146.690 253.770 146.860 ;
        RECT 251.100 146.190 251.270 146.360 ;
        RECT 251.600 146.190 251.770 146.360 ;
        RECT 252.100 146.190 252.270 146.360 ;
        RECT 252.600 146.190 252.770 146.360 ;
        RECT 253.100 146.190 253.270 146.360 ;
        RECT 253.600 146.190 253.770 146.360 ;
        RECT 251.100 145.690 251.270 145.860 ;
        RECT 251.600 145.690 251.770 145.860 ;
        RECT 252.100 145.690 252.270 145.860 ;
        RECT 252.600 145.690 252.770 145.860 ;
        RECT 253.100 145.690 253.270 145.860 ;
        RECT 253.600 145.690 253.770 145.860 ;
        RECT 251.100 145.190 251.270 145.360 ;
        RECT 251.600 145.190 251.770 145.360 ;
        RECT 252.100 145.190 252.270 145.360 ;
        RECT 252.600 145.190 252.770 145.360 ;
        RECT 253.100 145.190 253.270 145.360 ;
        RECT 253.600 145.190 253.770 145.360 ;
        RECT 251.100 144.690 251.270 144.860 ;
        RECT 251.600 144.690 251.770 144.860 ;
        RECT 252.100 144.690 252.270 144.860 ;
        RECT 252.600 144.690 252.770 144.860 ;
        RECT 253.100 144.690 253.270 144.860 ;
        RECT 253.600 144.690 253.770 144.860 ;
        RECT 257.800 147.190 257.970 147.360 ;
        RECT 258.300 147.190 258.470 147.360 ;
        RECT 258.800 147.190 258.970 147.360 ;
        RECT 259.300 147.190 259.470 147.360 ;
        RECT 259.800 147.190 259.970 147.360 ;
        RECT 260.300 147.190 260.470 147.360 ;
        RECT 257.800 146.690 257.970 146.860 ;
        RECT 258.300 146.690 258.470 146.860 ;
        RECT 258.800 146.690 258.970 146.860 ;
        RECT 259.300 146.690 259.470 146.860 ;
        RECT 259.800 146.690 259.970 146.860 ;
        RECT 260.300 146.690 260.470 146.860 ;
        RECT 257.800 146.190 257.970 146.360 ;
        RECT 258.300 146.190 258.470 146.360 ;
        RECT 258.800 146.190 258.970 146.360 ;
        RECT 259.300 146.190 259.470 146.360 ;
        RECT 259.800 146.190 259.970 146.360 ;
        RECT 260.300 146.190 260.470 146.360 ;
        RECT 257.800 145.690 257.970 145.860 ;
        RECT 258.300 145.690 258.470 145.860 ;
        RECT 258.800 145.690 258.970 145.860 ;
        RECT 259.300 145.690 259.470 145.860 ;
        RECT 259.800 145.690 259.970 145.860 ;
        RECT 260.300 145.690 260.470 145.860 ;
        RECT 257.800 145.190 257.970 145.360 ;
        RECT 258.300 145.190 258.470 145.360 ;
        RECT 258.800 145.190 258.970 145.360 ;
        RECT 259.300 145.190 259.470 145.360 ;
        RECT 259.800 145.190 259.970 145.360 ;
        RECT 260.300 145.190 260.470 145.360 ;
        RECT 257.800 144.690 257.970 144.860 ;
        RECT 258.300 144.690 258.470 144.860 ;
        RECT 258.800 144.690 258.970 144.860 ;
        RECT 259.300 144.690 259.470 144.860 ;
        RECT 259.800 144.690 259.970 144.860 ;
        RECT 260.300 144.690 260.470 144.860 ;
        RECT 201.335 143.935 201.505 144.105 ;
        RECT 201.335 143.575 201.505 143.745 ;
        RECT 201.335 143.215 201.505 143.385 ;
        RECT 112.095 128.015 114.065 130.705 ;
        RECT 122.130 128.015 124.100 130.705 ;
        RECT 112.095 123.215 114.065 125.905 ;
        RECT 122.130 123.215 124.100 125.905 ;
        RECT 127.150 129.275 127.320 129.445 ;
        RECT 127.150 128.915 127.320 129.085 ;
        RECT 127.150 128.555 127.320 128.725 ;
        RECT 127.150 128.195 127.320 128.365 ;
        RECT 127.150 127.835 127.320 128.005 ;
        RECT 127.150 127.475 127.320 127.645 ;
        RECT 127.150 127.115 127.320 127.285 ;
        RECT 127.150 126.755 127.320 126.925 ;
        RECT 127.150 126.395 127.320 126.565 ;
        RECT 127.150 126.035 127.320 126.205 ;
        RECT 127.150 125.675 127.320 125.845 ;
        RECT 131.730 129.275 131.900 129.445 ;
        RECT 131.730 128.915 131.900 129.085 ;
        RECT 131.730 128.555 131.900 128.725 ;
        RECT 131.730 128.195 131.900 128.365 ;
        RECT 131.730 127.835 131.900 128.005 ;
        RECT 131.730 127.475 131.900 127.645 ;
        RECT 131.730 127.115 131.900 127.285 ;
        RECT 131.730 126.755 131.900 126.925 ;
        RECT 131.730 126.395 131.900 126.565 ;
        RECT 131.730 126.035 131.900 126.205 ;
        RECT 131.730 125.675 131.900 125.845 ;
        RECT 136.310 129.275 136.480 129.445 ;
        RECT 136.310 128.915 136.480 129.085 ;
        RECT 136.310 128.555 136.480 128.725 ;
        RECT 136.310 128.195 136.480 128.365 ;
        RECT 136.310 127.835 136.480 128.005 ;
        RECT 136.310 127.475 136.480 127.645 ;
        RECT 136.310 127.115 136.480 127.285 ;
        RECT 136.310 126.755 136.480 126.925 ;
        RECT 136.310 126.395 136.480 126.565 ;
        RECT 136.310 126.035 136.480 126.205 ;
        RECT 136.310 125.675 136.480 125.845 ;
        RECT 140.890 129.275 141.060 129.445 ;
        RECT 140.890 128.915 141.060 129.085 ;
        RECT 140.890 128.555 141.060 128.725 ;
        RECT 140.890 128.195 141.060 128.365 ;
        RECT 140.890 127.835 141.060 128.005 ;
        RECT 140.890 127.475 141.060 127.645 ;
        RECT 140.890 127.115 141.060 127.285 ;
        RECT 140.890 126.755 141.060 126.925 ;
        RECT 140.890 126.395 141.060 126.565 ;
        RECT 140.890 126.035 141.060 126.205 ;
        RECT 140.890 125.675 141.060 125.845 ;
        RECT 145.470 129.275 145.640 129.445 ;
        RECT 145.470 128.915 145.640 129.085 ;
        RECT 145.470 128.555 145.640 128.725 ;
        RECT 145.470 128.195 145.640 128.365 ;
        RECT 145.470 127.835 145.640 128.005 ;
        RECT 187.065 128.015 189.035 130.705 ;
        RECT 197.100 128.015 199.070 130.705 ;
        RECT 145.470 127.475 145.640 127.645 ;
        RECT 145.470 127.115 145.640 127.285 ;
        RECT 145.470 126.755 145.640 126.925 ;
        RECT 145.470 126.395 145.640 126.565 ;
        RECT 145.470 126.035 145.640 126.205 ;
        RECT 145.470 125.675 145.640 125.845 ;
        RECT 187.065 123.215 189.035 125.905 ;
        RECT 200.785 128.015 202.755 130.705 ;
        RECT 210.820 128.015 212.790 130.705 ;
        RECT 197.100 123.215 199.070 125.905 ;
        RECT 200.785 123.215 202.755 125.905 ;
        RECT 214.505 128.015 216.475 130.705 ;
        RECT 224.540 128.015 226.510 130.705 ;
        RECT 210.820 123.215 212.790 125.905 ;
        RECT 214.505 123.215 216.475 125.905 ;
        RECT 228.225 128.015 230.195 130.705 ;
        RECT 238.260 128.015 240.230 130.705 ;
        RECT 224.540 123.215 226.510 125.905 ;
        RECT 241.945 128.015 243.915 130.705 ;
        RECT 251.980 128.015 253.950 130.705 ;
        RECT 238.260 123.215 240.230 125.905 ;
        RECT 241.945 123.215 243.915 125.905 ;
        RECT 251.980 123.215 253.950 125.905 ;
        RECT 119.445 109.215 121.415 111.905 ;
        RECT 129.480 109.215 131.450 111.905 ;
        RECT 119.445 104.415 121.415 107.105 ;
        RECT 136.105 109.215 138.075 111.905 ;
        RECT 146.140 109.215 148.110 111.905 ;
        RECT 129.480 104.415 131.450 107.105 ;
        RECT 136.105 104.415 138.075 107.105 ;
        RECT 149.825 109.215 151.795 111.905 ;
        RECT 159.860 109.215 161.830 111.905 ;
        RECT 146.140 104.415 148.110 107.105 ;
        RECT 149.825 104.415 151.795 107.105 ;
        RECT 165.995 109.215 167.965 111.905 ;
        RECT 176.030 109.215 178.000 111.905 ;
        RECT 159.860 104.415 161.830 107.105 ;
        RECT 165.995 104.415 167.965 107.105 ;
        RECT 187.065 109.215 189.035 111.905 ;
        RECT 197.100 109.215 199.070 111.905 ;
        RECT 176.030 104.415 178.000 107.105 ;
        RECT 187.065 104.415 189.035 107.105 ;
        RECT 200.785 109.215 202.755 111.905 ;
        RECT 210.820 109.215 212.790 111.905 ;
        RECT 197.100 104.415 199.070 107.105 ;
        RECT 200.785 104.415 202.755 107.105 ;
        RECT 251.980 109.215 253.950 111.905 ;
        RECT 210.820 104.415 212.790 107.105 ;
        RECT 241.945 104.415 243.915 107.105 ;
        RECT 251.980 104.415 253.950 107.105 ;
        RECT 127.105 85.595 127.275 85.765 ;
        RECT 219.405 71.615 221.375 74.305 ;
        RECT 229.440 71.615 231.410 74.305 ;
        RECT 219.405 66.815 221.375 69.505 ;
        RECT 233.125 71.615 235.095 74.305 ;
        RECT 243.160 71.615 245.130 74.305 ;
        RECT 229.440 66.815 231.410 69.505 ;
        RECT 233.125 66.815 235.095 69.505 ;
        RECT 246.845 71.615 248.815 74.305 ;
        RECT 256.880 71.615 258.850 74.305 ;
        RECT 243.160 66.815 245.130 69.505 ;
        RECT 246.845 66.815 248.815 69.505 ;
        RECT 256.880 66.815 258.850 69.505 ;
        RECT 228.950 52.815 230.920 55.505 ;
        RECT 218.915 48.015 220.885 50.705 ;
        RECT 232.635 52.815 234.605 55.505 ;
        RECT 242.670 52.815 244.640 55.505 ;
        RECT 228.950 48.015 230.920 50.705 ;
        RECT 232.635 48.015 234.605 50.705 ;
        RECT 246.355 52.815 248.325 55.505 ;
        RECT 256.390 52.815 258.360 55.505 ;
        RECT 242.670 48.015 244.640 50.705 ;
        RECT 246.355 48.015 248.325 50.705 ;
        RECT 256.390 48.015 258.360 50.705 ;
        RECT 222.835 34.015 224.805 36.705 ;
        RECT 232.870 34.015 234.840 36.705 ;
        RECT 222.835 29.215 224.805 31.905 ;
        RECT 236.555 34.015 238.525 36.705 ;
        RECT 246.590 34.015 248.560 36.705 ;
        RECT 232.870 29.215 234.840 31.905 ;
        RECT 250.275 34.015 252.245 36.705 ;
        RECT 260.310 34.015 262.280 36.705 ;
        RECT 246.590 29.215 248.560 31.905 ;
        RECT 250.275 29.215 252.245 31.905 ;
        RECT 260.310 29.215 262.280 31.905 ;
      LAYER met1 ;
        RECT 104.215 240.755 106.265 243.565 ;
        RECT 114.255 240.755 116.305 243.565 ;
        RECT 105.040 240.340 105.180 240.755 ;
        RECT 104.950 240.080 105.270 240.340 ;
        RECT 97.130 236.540 97.450 236.600 ;
        RECT 104.215 236.540 106.265 238.765 ;
        RECT 97.130 236.400 106.265 236.540 ;
        RECT 97.130 236.340 97.450 236.400 ;
        RECT 104.215 235.955 106.265 236.400 ;
        RECT 114.200 235.935 116.360 240.755 ;
        RECT 119.620 238.580 119.850 242.360 ;
        RECT 119.620 238.440 120.360 238.580 ;
        RECT 119.620 238.360 119.850 238.440 ;
        RECT 118.750 236.200 119.070 236.260 ;
        RECT 120.220 236.245 120.360 238.440 ;
        RECT 120.145 236.200 120.435 236.245 ;
        RECT 147.270 236.200 147.590 236.260 ;
        RECT 118.750 236.060 120.435 236.200 ;
        RECT 146.995 236.060 147.590 236.200 ;
        RECT 118.750 236.000 119.070 236.060 ;
        RECT 120.145 236.015 120.435 236.060 ;
        RECT 147.270 236.000 147.590 236.060 ;
        RECT 70.620 219.560 70.850 223.560 ;
        RECT 216.620 219.730 259.880 222.790 ;
        RECT 220.500 219.260 220.640 219.730 ;
        RECT 220.410 219.000 220.730 219.260 ;
        RECT 71.830 218.520 72.150 218.580 ;
        RECT 71.555 218.380 72.150 218.520 ;
        RECT 71.830 218.320 72.150 218.380 ;
        RECT 72.750 217.500 73.070 217.560 ;
        RECT 72.475 217.360 73.070 217.500 ;
        RECT 72.750 217.300 73.070 217.360 ;
        RECT 147.270 217.330 147.590 217.390 ;
        RECT 146.995 217.190 147.590 217.330 ;
        RECT 147.270 217.130 147.590 217.190 ;
        RECT 141.750 199.820 142.070 199.880 ;
        RECT 146.895 199.820 147.125 205.985 ;
        RECT 141.750 199.680 147.125 199.820 ;
        RECT 141.750 199.620 142.070 199.680 ;
        RECT 146.895 199.535 147.125 199.680 ;
        RECT 151.475 199.535 151.705 205.985 ;
        RECT 156.055 199.535 156.285 205.985 ;
        RECT 160.635 199.535 160.865 205.985 ;
        RECT 165.215 199.535 165.445 205.985 ;
        RECT 169.795 199.535 170.025 205.985 ;
        RECT 174.375 199.535 174.605 205.985 ;
        RECT 186.410 200.760 186.640 204.760 ;
        RECT 188.700 200.760 188.930 204.760 ;
        RECT 190.990 201.180 191.220 204.760 ;
        RECT 192.810 201.180 193.130 201.240 ;
        RECT 190.990 201.040 193.130 201.180 ;
        RECT 190.990 200.760 191.220 201.040 ;
        RECT 192.810 200.980 193.130 201.040 ;
        RECT 193.280 200.760 193.510 204.760 ;
        RECT 195.570 200.760 195.800 204.760 ;
        RECT 197.860 200.760 198.090 204.760 ;
        RECT 200.150 200.760 200.380 204.760 ;
        RECT 202.440 200.760 202.670 204.760 ;
        RECT 204.730 200.760 204.960 204.760 ;
        RECT 207.020 200.760 207.250 204.760 ;
        RECT 210.740 200.930 260.700 203.990 ;
        RECT 179.010 200.500 179.330 200.560 ;
        RECT 188.760 200.500 188.900 200.760 ;
        RECT 179.010 200.360 188.900 200.500 ;
        RECT 179.010 200.300 179.330 200.360 ;
        RECT 118.750 199.140 119.070 199.200 ;
        RECT 118.750 199.000 139.680 199.140 ;
        RECT 118.750 198.940 119.070 199.000 ;
        RECT 139.540 198.800 139.680 199.000 ;
        RECT 140.830 198.800 141.150 198.860 ;
        RECT 139.540 198.660 141.150 198.800 ;
        RECT 140.830 198.600 141.150 198.660 ;
        RECT 147.270 198.460 147.590 198.520 ;
        RECT 146.995 198.320 147.590 198.460 ;
        RECT 147.270 198.260 147.590 198.320 ;
        RECT 71.830 190.440 72.150 190.700 ;
        RECT 71.920 190.300 72.060 190.440 ;
        RECT 128.870 190.300 129.190 190.360 ;
        RECT 71.920 190.160 129.190 190.300 ;
        RECT 128.870 190.100 129.190 190.160 ;
        RECT 172.110 189.960 172.430 190.020 ;
        RECT 179.010 189.960 179.330 190.020 ;
        RECT 172.110 189.820 179.330 189.960 ;
        RECT 172.110 189.760 172.430 189.820 ;
        RECT 179.010 189.760 179.330 189.820 ;
        RECT 111.390 187.580 111.710 187.640 ;
        RECT 108.260 187.440 111.710 187.580 ;
        RECT 68.445 184.520 70.495 187.165 ;
        RECT 77.810 184.520 78.130 184.580 ;
        RECT 68.445 184.380 78.130 184.520 ;
        RECT 68.445 184.355 70.495 184.380 ;
        RECT 77.810 184.320 78.130 184.380 ;
        RECT 78.485 184.355 80.535 187.165 ;
        RECT 82.165 184.355 84.215 187.165 ;
        RECT 92.205 184.355 94.255 187.165 ;
        RECT 95.890 186.900 97.940 187.165 ;
        RECT 108.260 186.900 108.400 187.440 ;
        RECT 111.390 187.380 111.710 187.440 ;
        RECT 95.890 186.760 108.400 186.900 ;
        RECT 95.890 184.355 97.940 186.760 ;
        RECT 108.800 184.355 110.850 187.165 ;
        RECT 111.850 184.520 112.170 184.580 ;
        RECT 112.545 184.520 114.595 187.165 ;
        RECT 111.850 184.380 114.595 184.520 ;
        RECT 68.445 179.555 70.495 182.365 ;
        RECT 78.430 179.535 80.590 184.355 ;
        RECT 82.870 184.320 83.190 184.355 ;
        RECT 81.030 182.140 81.350 182.200 ;
        RECT 82.165 182.140 84.215 182.365 ;
        RECT 81.030 182.000 84.215 182.140 ;
        RECT 81.030 181.940 81.350 182.000 ;
        RECT 82.165 179.555 84.215 182.000 ;
        RECT 92.150 179.535 94.310 184.355 ;
        RECT 108.745 179.535 110.905 184.355 ;
        RECT 111.850 184.320 112.170 184.380 ;
        RECT 112.545 184.355 114.595 184.380 ;
        RECT 122.585 184.355 124.635 187.165 ;
        RECT 111.390 182.140 111.710 182.200 ;
        RECT 112.545 182.140 114.595 182.365 ;
        RECT 111.390 182.000 114.595 182.140 ;
        RECT 111.390 181.940 111.710 182.000 ;
        RECT 112.545 179.555 114.595 182.000 ;
        RECT 122.530 179.535 124.690 184.355 ;
        RECT 127.120 181.960 127.350 185.960 ;
        RECT 128.870 185.880 129.190 185.940 ;
        RECT 129.410 185.880 129.640 185.960 ;
        RECT 128.870 185.740 129.640 185.880 ;
        RECT 128.870 185.680 129.190 185.740 ;
        RECT 129.410 181.960 129.640 185.740 ;
        RECT 131.700 181.960 131.930 185.960 ;
        RECT 133.990 181.960 134.220 185.960 ;
        RECT 136.280 181.960 136.510 185.960 ;
        RECT 138.570 181.960 138.800 185.960 ;
        RECT 140.860 181.960 141.090 185.960 ;
        RECT 143.150 181.960 143.380 185.960 ;
        RECT 145.440 184.860 145.670 185.960 ;
        RECT 147.730 185.880 147.960 185.960 ;
        RECT 172.110 185.880 172.430 185.940 ;
        RECT 147.730 185.740 172.430 185.880 ;
        RECT 147.270 184.860 147.590 184.920 ;
        RECT 145.440 184.720 147.590 184.860 ;
        RECT 145.440 181.960 145.670 184.720 ;
        RECT 147.270 184.660 147.590 184.720 ;
        RECT 147.730 181.960 147.960 185.740 ;
        RECT 172.110 185.680 172.430 185.740 ;
        RECT 187.565 180.735 187.795 187.185 ;
        RECT 192.145 180.735 192.375 187.185 ;
        RECT 196.725 180.735 196.955 187.185 ;
        RECT 201.305 180.735 201.535 187.185 ;
        RECT 210.740 182.130 260.700 185.190 ;
        RECT 187.765 180.160 188.055 180.315 ;
        RECT 187.750 179.900 188.070 180.160 ;
        RECT 192.810 179.760 193.130 179.820 ;
        RECT 192.535 179.620 193.130 179.760 ;
        RECT 192.810 179.560 193.130 179.620 ;
        RECT 96.375 165.555 98.425 168.365 ;
        RECT 106.415 165.555 108.465 168.365 ;
        RECT 110.100 165.820 112.150 168.365 ;
        RECT 122.430 165.820 122.750 165.880 ;
        RECT 110.100 165.680 122.750 165.820 ;
        RECT 110.100 165.555 112.150 165.680 ;
        RECT 122.430 165.620 122.750 165.680 ;
        RECT 123.010 165.555 125.060 168.365 ;
        RECT 82.870 163.440 83.190 163.500 ;
        RECT 96.375 163.440 98.425 163.565 ;
        RECT 82.870 163.300 98.425 163.440 ;
        RECT 82.870 163.240 83.190 163.300 ;
        RECT 96.375 160.755 98.425 163.300 ;
        RECT 106.360 160.735 108.520 165.555 ;
        RECT 122.955 160.735 125.115 165.555 ;
        RECT 210.740 163.330 260.700 166.390 ;
        RECT 211.210 163.240 211.530 163.330 ;
        RECT 104.490 150.180 104.810 150.240 ;
        RECT 111.850 150.180 112.170 150.240 ;
        RECT 104.490 150.040 112.170 150.180 ;
        RECT 104.490 149.980 104.810 150.040 ;
        RECT 111.850 149.980 112.170 150.040 ;
        RECT 82.655 146.755 84.705 149.565 ;
        RECT 92.695 146.755 94.745 149.565 ;
        RECT 95.290 147.120 95.610 147.180 ;
        RECT 96.375 147.120 98.425 149.565 ;
        RECT 95.290 146.980 98.425 147.120 ;
        RECT 95.290 146.920 95.610 146.980 ;
        RECT 96.375 146.755 98.425 146.980 ;
        RECT 106.415 146.755 108.465 149.565 ;
        RECT 120.135 146.755 122.185 149.565 ;
        RECT 136.065 146.755 138.115 149.565 ;
        RECT 146.105 146.755 148.155 149.565 ;
        RECT 82.655 144.740 84.705 144.765 ;
        RECT 92.070 144.740 92.390 144.800 ;
        RECT 82.655 144.600 92.390 144.740 ;
        RECT 82.655 141.955 84.705 144.600 ;
        RECT 92.070 144.540 92.390 144.600 ;
        RECT 92.640 141.935 94.800 146.755 ;
        RECT 96.375 144.740 98.425 144.765 ;
        RECT 104.490 144.740 104.810 144.800 ;
        RECT 96.375 144.600 104.810 144.740 ;
        RECT 96.375 141.955 98.425 144.600 ;
        RECT 104.490 144.540 104.810 144.600 ;
        RECT 106.360 141.935 108.520 146.755 ;
        RECT 108.660 144.740 108.920 144.830 ;
        RECT 110.095 144.740 112.145 144.765 ;
        RECT 108.660 144.600 112.145 144.740 ;
        RECT 108.660 144.510 108.920 144.600 ;
        RECT 110.095 141.955 112.145 144.600 ;
        RECT 120.080 141.935 122.240 146.755 ;
        RECT 122.430 144.740 122.750 144.800 ;
        RECT 136.065 144.740 138.115 144.765 ;
        RECT 122.430 144.600 138.115 144.740 ;
        RECT 122.430 144.540 122.750 144.600 ;
        RECT 136.065 141.955 138.115 144.600 ;
        RECT 146.050 141.935 148.210 146.755 ;
        RECT 187.565 143.135 187.795 149.585 ;
        RECT 192.145 143.135 192.375 149.585 ;
        RECT 196.725 143.135 196.955 149.585 ;
        RECT 201.305 143.135 201.535 149.585 ;
        RECT 210.740 144.530 260.700 147.590 ;
        RECT 192.825 142.515 193.115 142.745 ;
        RECT 192.900 142.080 193.040 142.515 ;
        RECT 192.810 142.020 193.130 142.080 ;
        RECT 192.535 141.880 193.130 142.020 ;
        RECT 192.810 141.820 193.130 141.880 ;
        RECT 199.710 131.140 200.030 131.200 ;
        RECT 188.760 131.000 200.030 131.140 ;
        RECT 188.760 130.765 188.900 131.000 ;
        RECT 199.710 130.940 200.030 131.000 ;
        RECT 207.160 131.000 228.460 131.140 ;
        RECT 207.160 130.860 207.300 131.000 ;
        RECT 69.530 129.440 69.850 129.500 ;
        RECT 112.055 129.440 114.105 130.765 ;
        RECT 69.530 129.300 114.105 129.440 ;
        RECT 69.530 129.240 69.850 129.300 ;
        RECT 112.055 127.955 114.105 129.300 ;
        RECT 122.095 127.955 124.145 130.765 ;
        RECT 112.055 123.320 114.105 125.965 ;
        RECT 114.610 123.320 114.930 123.380 ;
        RECT 112.055 123.180 114.930 123.320 ;
        RECT 112.055 123.155 114.105 123.180 ;
        RECT 114.610 123.120 114.930 123.180 ;
        RECT 122.040 123.135 124.200 127.955 ;
        RECT 127.120 125.760 127.350 129.560 ;
        RECT 127.030 125.500 127.350 125.760 ;
        RECT 131.700 125.560 131.930 129.560 ;
        RECT 136.280 125.560 136.510 129.560 ;
        RECT 140.860 125.560 141.090 129.560 ;
        RECT 145.440 128.760 145.670 129.560 ;
        RECT 147.270 128.760 147.590 128.820 ;
        RECT 145.440 128.620 147.590 128.760 ;
        RECT 145.440 125.560 145.670 128.620 ;
        RECT 147.270 128.560 147.590 128.620 ;
        RECT 187.025 127.955 189.075 130.765 ;
        RECT 197.065 127.955 199.115 130.765 ;
        RECT 200.745 128.140 202.795 130.765 ;
        RECT 207.070 130.600 207.390 130.860 ;
        RECT 228.320 130.765 228.460 131.000 ;
        RECT 200.630 127.955 202.795 128.140 ;
        RECT 210.785 127.955 212.835 130.765 ;
        RECT 213.510 128.420 213.830 128.480 ;
        RECT 214.465 128.420 216.515 130.765 ;
        RECT 213.510 128.280 216.515 128.420 ;
        RECT 213.510 128.220 213.830 128.280 ;
        RECT 214.465 127.955 216.515 128.280 ;
        RECT 224.505 127.955 226.555 130.765 ;
        RECT 228.185 127.955 230.235 130.765 ;
        RECT 238.225 127.955 240.275 130.765 ;
        RECT 241.905 127.955 243.955 130.765 ;
        RECT 251.945 127.955 253.995 130.765 ;
        RECT 187.025 123.380 189.075 125.965 ;
        RECT 186.830 123.155 189.075 123.380 ;
        RECT 186.830 123.120 187.150 123.155 ;
        RECT 197.010 123.135 199.170 127.955 ;
        RECT 200.630 127.880 200.950 127.955 ;
        RECT 199.710 125.700 200.030 125.760 ;
        RECT 200.745 125.700 202.795 125.965 ;
        RECT 199.710 125.560 202.795 125.700 ;
        RECT 199.710 125.500 200.030 125.560 ;
        RECT 200.745 123.155 202.795 125.560 ;
        RECT 210.730 123.135 212.890 127.955 ;
        RECT 214.465 123.380 216.515 125.965 ;
        RECT 214.430 123.155 216.515 123.380 ;
        RECT 214.430 123.120 214.750 123.155 ;
        RECT 224.450 123.135 226.610 127.955 ;
        RECT 238.170 123.135 240.330 127.955 ;
        RECT 242.950 127.880 243.270 127.955 ;
        RECT 241.905 123.155 243.955 125.965 ;
        RECT 251.890 123.135 254.050 127.955 ;
        RECT 191.430 120.940 191.750 121.000 ;
        RECT 214.430 120.940 214.750 121.000 ;
        RECT 191.430 120.800 214.750 120.940 ;
        RECT 191.430 120.740 191.750 120.800 ;
        RECT 214.430 120.740 214.750 120.800 ;
        RECT 154.630 117.200 154.950 117.260 ;
        RECT 186.830 117.200 187.150 117.260 ;
        RECT 154.630 117.060 187.150 117.200 ;
        RECT 154.630 117.000 154.950 117.060 ;
        RECT 186.830 117.000 187.150 117.060 ;
        RECT 174.870 112.440 175.190 112.500 ;
        RECT 200.630 112.440 200.950 112.500 ;
        RECT 213.510 112.440 213.830 112.500 ;
        RECT 174.870 112.300 200.950 112.440 ;
        RECT 174.870 112.240 175.190 112.300 ;
        RECT 200.630 112.240 200.950 112.300 ;
        RECT 202.560 112.300 213.830 112.440 ;
        RECT 202.560 111.965 202.700 112.300 ;
        RECT 213.510 112.240 213.830 112.300 ;
        RECT 114.610 111.760 114.930 111.820 ;
        RECT 119.405 111.760 121.455 111.965 ;
        RECT 114.610 111.620 121.455 111.760 ;
        RECT 114.610 111.560 114.930 111.620 ;
        RECT 119.405 109.155 121.455 111.620 ;
        RECT 129.445 109.155 131.495 111.965 ;
        RECT 136.065 109.380 138.115 111.965 ;
        RECT 145.430 109.380 145.750 109.440 ;
        RECT 136.065 109.240 145.750 109.380 ;
        RECT 136.065 109.155 138.115 109.240 ;
        RECT 145.430 109.180 145.750 109.240 ;
        RECT 146.105 109.155 148.155 111.965 ;
        RECT 149.785 111.760 151.835 111.965 ;
        RECT 154.630 111.760 154.950 111.820 ;
        RECT 149.785 111.620 154.950 111.760 ;
        RECT 149.785 109.155 151.835 111.620 ;
        RECT 154.630 111.560 154.950 111.620 ;
        RECT 159.825 109.155 161.875 111.965 ;
        RECT 165.955 109.380 168.005 111.965 ;
        RECT 175.330 109.380 175.650 109.440 ;
        RECT 165.955 109.240 175.650 109.380 ;
        RECT 165.955 109.155 168.005 109.240 ;
        RECT 175.330 109.180 175.650 109.240 ;
        RECT 175.995 109.155 178.045 111.965 ;
        RECT 187.025 111.760 189.075 111.965 ;
        RECT 191.430 111.760 191.750 111.820 ;
        RECT 187.025 111.620 191.750 111.760 ;
        RECT 187.025 109.155 189.075 111.620 ;
        RECT 191.430 111.560 191.750 111.620 ;
        RECT 197.065 109.155 199.115 111.965 ;
        RECT 200.745 109.155 202.795 111.965 ;
        RECT 210.785 109.155 212.835 111.965 ;
        RECT 251.945 109.155 253.995 111.965 ;
        RECT 83.330 107.000 83.650 107.060 ;
        RECT 119.405 107.000 121.455 107.165 ;
        RECT 83.330 106.860 121.455 107.000 ;
        RECT 83.330 106.800 83.650 106.860 ;
        RECT 119.405 104.355 121.455 106.860 ;
        RECT 129.390 104.335 131.550 109.155 ;
        RECT 136.065 104.355 138.115 107.165 ;
        RECT 146.050 104.335 148.210 109.155 ;
        RECT 148.650 107.000 148.970 107.060 ;
        RECT 149.785 107.000 151.835 107.165 ;
        RECT 148.650 106.860 151.835 107.000 ;
        RECT 148.650 106.800 148.970 106.860 ;
        RECT 149.785 104.355 151.835 106.860 ;
        RECT 159.770 104.335 161.930 109.155 ;
        RECT 165.955 107.000 168.005 107.165 ;
        RECT 174.870 107.000 175.190 107.060 ;
        RECT 165.955 106.860 175.190 107.000 ;
        RECT 165.955 104.355 168.005 106.860 ;
        RECT 174.870 106.800 175.190 106.860 ;
        RECT 175.940 104.335 178.100 109.155 ;
        RECT 178.550 107.000 178.870 107.060 ;
        RECT 187.025 107.000 189.075 107.165 ;
        RECT 178.550 106.860 189.075 107.000 ;
        RECT 178.550 106.800 178.870 106.860 ;
        RECT 187.025 104.355 189.075 106.860 ;
        RECT 197.010 104.335 199.170 109.155 ;
        RECT 200.745 107.000 202.795 107.165 ;
        RECT 207.070 107.000 207.390 107.060 ;
        RECT 200.745 106.860 207.390 107.000 ;
        RECT 200.745 104.355 202.795 106.860 ;
        RECT 207.070 106.800 207.390 106.860 ;
        RECT 210.730 104.335 212.890 109.155 ;
        RECT 241.905 104.355 243.955 107.165 ;
        RECT 251.890 104.335 254.050 109.155 ;
        RECT 127.030 85.720 127.350 85.980 ;
        RECT 127.045 85.565 127.335 85.720 ;
        RECT 245.250 75.040 245.570 75.100 ;
        RECT 220.960 74.900 245.570 75.040 ;
        RECT 220.960 74.365 221.100 74.900 ;
        RECT 245.250 74.840 245.570 74.900 ;
        RECT 221.880 74.560 245.480 74.700 ;
        RECT 221.880 74.420 222.020 74.560 ;
        RECT 219.365 71.555 221.415 74.365 ;
        RECT 221.790 74.160 222.110 74.420 ;
        RECT 229.405 71.555 231.455 74.365 ;
        RECT 233.085 71.555 235.135 74.365 ;
        RECT 243.125 71.555 245.175 74.365 ;
        RECT 245.340 74.360 245.480 74.560 ;
        RECT 246.805 74.360 248.855 74.365 ;
        RECT 245.340 74.220 248.855 74.360 ;
        RECT 246.805 71.555 248.855 74.220 ;
        RECT 256.845 71.555 258.895 74.365 ;
        RECT 219.365 69.320 221.415 69.565 ;
        RECT 219.365 69.060 221.650 69.320 ;
        RECT 219.365 66.755 221.415 69.060 ;
        RECT 229.350 66.735 231.510 71.555 ;
        RECT 233.290 71.440 233.610 71.555 ;
        RECT 233.085 66.755 235.135 69.565 ;
        RECT 234.670 66.680 234.990 66.755 ;
        RECT 243.070 66.735 245.230 71.555 ;
        RECT 246.805 66.755 248.855 69.565 ;
        RECT 247.550 66.680 247.870 66.755 ;
        RECT 256.790 66.735 258.950 71.555 ;
        RECT 223.630 56.000 223.950 56.060 ;
        RECT 234.670 56.000 234.990 56.060 ;
        RECT 223.630 55.860 231.680 56.000 ;
        RECT 223.630 55.800 223.950 55.860 ;
        RECT 228.915 52.755 230.965 55.565 ;
        RECT 231.540 55.320 231.680 55.860 ;
        RECT 234.670 55.860 245.020 56.000 ;
        RECT 234.670 55.800 234.990 55.860 ;
        RECT 232.595 55.320 234.645 55.565 ;
        RECT 231.540 55.180 234.645 55.320 ;
        RECT 232.595 52.755 234.645 55.180 ;
        RECT 242.635 52.755 244.685 55.565 ;
        RECT 244.880 55.320 245.020 55.860 ;
        RECT 246.315 55.320 248.365 55.565 ;
        RECT 244.880 55.180 248.365 55.320 ;
        RECT 246.315 52.755 248.365 55.180 ;
        RECT 256.355 52.755 258.405 55.565 ;
        RECT 218.875 48.180 220.925 50.765 ;
        RECT 228.230 48.180 228.550 48.240 ;
        RECT 218.875 48.040 228.550 48.180 ;
        RECT 218.875 47.955 220.925 48.040 ;
        RECT 228.230 47.980 228.550 48.040 ;
        RECT 228.860 47.935 231.020 52.755 ;
        RECT 232.595 47.955 234.645 50.765 ;
        RECT 242.580 47.935 244.740 52.755 ;
        RECT 245.250 50.560 245.570 50.620 ;
        RECT 246.315 50.560 248.365 50.765 ;
        RECT 245.250 50.420 248.365 50.560 ;
        RECT 245.250 50.360 245.570 50.420 ;
        RECT 246.315 47.955 248.365 50.420 ;
        RECT 256.300 47.935 258.460 52.755 ;
        RECT 228.230 46.820 228.550 46.880 ;
        RECT 249.390 46.820 249.710 46.880 ;
        RECT 228.230 46.680 249.710 46.820 ;
        RECT 228.230 46.620 228.550 46.680 ;
        RECT 249.390 46.620 249.710 46.680 ;
        RECT 248.930 37.300 249.250 37.360 ;
        RECT 232.460 37.160 249.250 37.300 ;
        RECT 222.795 36.620 224.845 36.765 ;
        RECT 232.460 36.620 232.600 37.160 ;
        RECT 248.930 37.100 249.250 37.160 ;
        RECT 222.795 36.480 232.600 36.620 ;
        RECT 222.795 33.955 224.845 36.480 ;
        RECT 232.835 33.955 234.885 36.765 ;
        RECT 236.515 36.620 238.565 36.765 ;
        RECT 245.710 36.620 246.030 36.680 ;
        RECT 236.515 36.480 246.030 36.620 ;
        RECT 236.515 33.955 238.565 36.480 ;
        RECT 245.710 36.420 246.030 36.480 ;
        RECT 246.555 33.955 248.605 36.765 ;
        RECT 249.390 36.620 249.710 36.680 ;
        RECT 250.235 36.620 252.285 36.765 ;
        RECT 249.390 36.480 252.285 36.620 ;
        RECT 249.390 36.420 249.710 36.480 ;
        RECT 250.235 33.955 252.285 36.480 ;
        RECT 260.275 33.955 262.325 36.765 ;
        RECT 222.795 29.155 224.845 31.965 ;
        RECT 232.780 29.135 234.940 33.955 ;
        RECT 246.500 29.135 248.660 33.955 ;
        RECT 248.930 31.860 249.250 31.920 ;
        RECT 250.235 31.860 252.285 31.965 ;
        RECT 248.930 31.720 252.285 31.860 ;
        RECT 248.930 31.660 249.250 31.720 ;
        RECT 250.235 29.155 252.285 31.720 ;
        RECT 260.220 29.135 262.380 33.955 ;
      LAYER via ;
        RECT 104.980 240.080 105.240 240.340 ;
        RECT 97.160 236.340 97.420 236.600 ;
        RECT 118.780 236.000 119.040 236.260 ;
        RECT 147.300 236.000 147.560 236.260 ;
        RECT 220.440 219.000 220.700 219.260 ;
        RECT 71.860 218.320 72.120 218.580 ;
        RECT 72.780 217.300 73.040 217.560 ;
        RECT 147.300 217.130 147.560 217.390 ;
        RECT 141.780 199.620 142.040 199.880 ;
        RECT 192.840 200.980 193.100 201.240 ;
        RECT 220.440 203.700 220.700 203.960 ;
        RECT 210.780 200.980 211.040 201.240 ;
        RECT 179.040 200.300 179.300 200.560 ;
        RECT 118.780 198.940 119.040 199.200 ;
        RECT 140.860 198.600 141.120 198.860 ;
        RECT 147.300 198.260 147.560 198.520 ;
        RECT 71.860 190.440 72.120 190.700 ;
        RECT 128.900 190.100 129.160 190.360 ;
        RECT 172.140 189.760 172.400 190.020 ;
        RECT 179.040 189.760 179.300 190.020 ;
        RECT 77.840 184.320 78.100 184.580 ;
        RECT 69.560 179.560 69.820 179.820 ;
        RECT 82.900 184.320 83.160 184.580 ;
        RECT 111.420 187.380 111.680 187.640 ;
        RECT 81.060 181.940 81.320 182.200 ;
        RECT 111.880 184.320 112.140 184.580 ;
        RECT 111.420 181.940 111.680 182.200 ;
        RECT 128.900 185.680 129.160 185.940 ;
        RECT 147.300 184.660 147.560 184.920 ;
        RECT 172.140 185.680 172.400 185.940 ;
        RECT 210.780 182.280 211.040 182.540 ;
        RECT 187.780 179.900 188.040 180.160 ;
        RECT 192.840 179.560 193.100 179.820 ;
        RECT 97.160 168.000 97.420 168.260 ;
        RECT 122.460 165.620 122.720 165.880 ;
        RECT 210.780 165.960 211.040 166.220 ;
        RECT 82.900 163.240 83.160 163.500 ;
        RECT 211.240 163.240 211.500 163.500 ;
        RECT 104.520 149.980 104.780 150.240 ;
        RECT 111.880 149.980 112.140 150.240 ;
        RECT 83.360 146.920 83.620 147.180 ;
        RECT 95.320 146.920 95.580 147.180 ;
        RECT 137.180 146.920 137.440 147.180 ;
        RECT 92.100 144.540 92.360 144.800 ;
        RECT 104.520 144.540 104.780 144.800 ;
        RECT 108.660 144.540 108.920 144.800 ;
        RECT 122.460 144.540 122.720 144.800 ;
        RECT 211.240 147.260 211.500 147.520 ;
        RECT 242.060 144.540 242.320 144.800 ;
        RECT 192.840 141.820 193.100 142.080 ;
        RECT 199.740 130.940 200.000 131.200 ;
        RECT 69.560 129.240 69.820 129.500 ;
        RECT 114.640 123.120 114.900 123.380 ;
        RECT 127.060 125.500 127.320 125.760 ;
        RECT 147.300 128.560 147.560 128.820 ;
        RECT 207.100 130.600 207.360 130.860 ;
        RECT 186.860 123.120 187.120 123.380 ;
        RECT 200.660 127.880 200.920 128.140 ;
        RECT 213.540 128.220 213.800 128.480 ;
        RECT 199.740 125.500 200.000 125.760 ;
        RECT 214.460 123.120 214.720 123.380 ;
        RECT 242.980 127.880 243.240 128.140 ;
        RECT 242.060 125.500 242.320 125.760 ;
        RECT 191.460 120.740 191.720 121.000 ;
        RECT 214.460 120.740 214.720 121.000 ;
        RECT 154.660 117.000 154.920 117.260 ;
        RECT 186.860 117.000 187.120 117.260 ;
        RECT 174.900 112.240 175.160 112.500 ;
        RECT 200.660 112.240 200.920 112.500 ;
        RECT 213.540 112.240 213.800 112.500 ;
        RECT 114.640 111.560 114.900 111.820 ;
        RECT 145.460 109.180 145.720 109.440 ;
        RECT 154.660 111.560 154.920 111.820 ;
        RECT 175.360 109.180 175.620 109.440 ;
        RECT 191.460 111.560 191.720 111.820 ;
        RECT 83.360 106.800 83.620 107.060 ;
        RECT 137.180 106.800 137.440 107.060 ;
        RECT 148.680 106.800 148.940 107.060 ;
        RECT 174.900 106.800 175.160 107.060 ;
        RECT 178.580 106.800 178.840 107.060 ;
        RECT 207.100 106.800 207.360 107.060 ;
        RECT 242.980 106.800 243.240 107.060 ;
        RECT 127.060 85.720 127.320 85.980 ;
        RECT 245.280 74.840 245.540 75.100 ;
        RECT 221.820 74.160 222.080 74.420 ;
        RECT 221.360 69.060 221.620 69.320 ;
        RECT 233.320 71.440 233.580 71.700 ;
        RECT 234.700 66.680 234.960 66.940 ;
        RECT 247.580 66.680 247.840 66.940 ;
        RECT 223.660 55.800 223.920 56.060 ;
        RECT 234.700 55.800 234.960 56.060 ;
        RECT 228.260 47.980 228.520 48.240 ;
        RECT 233.320 50.360 233.580 50.620 ;
        RECT 245.280 50.360 245.540 50.620 ;
        RECT 228.260 46.620 228.520 46.880 ;
        RECT 249.420 46.620 249.680 46.880 ;
        RECT 248.960 37.100 249.220 37.360 ;
        RECT 245.740 36.420 246.000 36.680 ;
        RECT 249.420 36.420 249.680 36.680 ;
        RECT 223.660 31.660 223.920 31.920 ;
        RECT 248.960 31.660 249.220 31.920 ;
      LAYER met2 ;
        RECT 104.980 240.050 105.240 240.370 ;
        RECT 97.160 236.310 97.420 236.630 ;
        RECT 71.860 218.290 72.120 218.610 ;
        RECT 71.920 190.730 72.060 218.290 ;
        RECT 72.780 217.405 73.040 217.590 ;
        RECT 72.770 217.035 73.050 217.405 ;
        RECT 71.860 190.410 72.120 190.730 ;
        RECT 77.840 184.520 78.100 184.610 ;
        RECT 77.840 184.380 81.260 184.520 ;
        RECT 77.840 184.290 78.100 184.380 ;
        RECT 81.120 182.230 81.260 184.380 ;
        RECT 82.900 184.290 83.160 184.610 ;
        RECT 81.060 181.910 81.320 182.230 ;
        RECT 69.560 179.530 69.820 179.850 ;
        RECT 69.620 129.530 69.760 179.530 ;
        RECT 82.960 163.530 83.100 184.290 ;
        RECT 97.220 168.290 97.360 236.310 ;
        RECT 97.160 167.970 97.420 168.290 ;
        RECT 82.900 163.210 83.160 163.530 ;
        RECT 104.520 149.950 104.780 150.270 ;
        RECT 83.360 146.890 83.620 147.210 ;
        RECT 95.320 147.120 95.580 147.210 ;
        RECT 92.160 146.980 95.580 147.120 ;
        RECT 69.560 129.210 69.820 129.530 ;
        RECT 83.420 107.090 83.560 146.890 ;
        RECT 92.160 144.830 92.300 146.980 ;
        RECT 95.320 146.890 95.580 146.980 ;
        RECT 104.580 144.830 104.720 149.950 ;
        RECT 105.040 145.760 105.180 240.050 ;
        RECT 118.780 235.970 119.040 236.290 ;
        RECT 147.300 235.970 147.560 236.290 ;
        RECT 118.840 217.405 118.980 235.970 ;
        RECT 147.360 217.420 147.500 235.970 ;
        RECT 220.440 218.970 220.700 219.290 ;
        RECT 118.770 217.035 119.050 217.405 ;
        RECT 147.300 217.100 147.560 217.420 ;
        RECT 118.840 199.230 118.980 217.035 ;
        RECT 141.780 199.590 142.040 199.910 ;
        RECT 118.780 198.910 119.040 199.230 ;
        RECT 140.860 198.800 141.120 198.890 ;
        RECT 141.840 198.800 141.980 199.590 ;
        RECT 140.860 198.660 141.980 198.800 ;
        RECT 140.860 198.570 141.120 198.660 ;
        RECT 147.360 198.550 147.500 217.100 ;
        RECT 220.500 203.990 220.640 218.970 ;
        RECT 220.440 203.670 220.700 203.990 ;
        RECT 192.840 200.950 193.100 201.270 ;
        RECT 210.780 200.950 211.040 201.270 ;
        RECT 179.040 200.270 179.300 200.590 ;
        RECT 147.300 198.230 147.560 198.550 ;
        RECT 128.900 190.070 129.160 190.390 ;
        RECT 111.420 187.350 111.680 187.670 ;
        RECT 111.480 182.230 111.620 187.350 ;
        RECT 128.960 185.970 129.100 190.070 ;
        RECT 128.900 185.650 129.160 185.970 ;
        RECT 147.360 185.075 147.500 198.230 ;
        RECT 179.100 190.050 179.240 200.270 ;
        RECT 172.140 189.730 172.400 190.050 ;
        RECT 179.040 189.730 179.300 190.050 ;
        RECT 172.200 185.970 172.340 189.730 ;
        RECT 172.140 185.650 172.400 185.970 ;
        RECT 147.290 184.705 147.570 185.075 ;
        RECT 147.300 184.630 147.560 184.705 ;
        RECT 111.880 184.290 112.140 184.610 ;
        RECT 147.360 184.590 147.500 184.630 ;
        RECT 111.420 181.910 111.680 182.230 ;
        RECT 111.940 150.270 112.080 184.290 ;
        RECT 149.740 179.660 150.540 180.160 ;
        RECT 187.770 179.825 188.050 180.195 ;
        RECT 192.900 179.850 193.040 200.950 ;
        RECT 210.840 182.570 210.980 200.950 ;
        RECT 210.780 182.250 211.040 182.570 ;
        RECT 187.840 179.710 187.980 179.825 ;
        RECT 192.840 179.530 193.100 179.850 ;
        RECT 122.460 165.590 122.720 165.910 ;
        RECT 111.880 149.950 112.140 150.270 ;
        RECT 105.040 145.620 108.860 145.760 ;
        RECT 108.720 144.830 108.860 145.620 ;
        RECT 122.520 144.830 122.660 165.590 ;
        RECT 131.120 160.860 131.920 161.360 ;
        RECT 168.360 160.860 169.160 161.360 ;
        RECT 137.180 146.890 137.440 147.210 ;
        RECT 92.100 144.510 92.360 144.830 ;
        RECT 104.520 144.510 104.780 144.830 ;
        RECT 108.660 144.510 108.920 144.830 ;
        RECT 122.460 144.510 122.720 144.830 ;
        RECT 127.060 125.470 127.320 125.790 ;
        RECT 114.640 123.090 114.900 123.410 ;
        RECT 114.700 111.850 114.840 123.090 ;
        RECT 114.640 111.530 114.900 111.850 ;
        RECT 83.360 106.770 83.620 107.090 ;
        RECT 127.120 86.010 127.260 125.470 ;
        RECT 137.240 107.090 137.380 146.890 ;
        RECT 149.740 142.060 150.540 142.560 ;
        RECT 192.900 142.110 193.040 179.530 ;
        RECT 210.840 166.250 210.980 182.250 ;
        RECT 210.780 165.930 211.040 166.250 ;
        RECT 211.240 163.210 211.500 163.530 ;
        RECT 211.300 147.550 211.440 163.210 ;
        RECT 211.240 147.230 211.500 147.550 ;
        RECT 242.060 144.510 242.320 144.830 ;
        RECT 192.840 141.790 193.100 142.110 ;
        RECT 199.740 130.910 200.000 131.230 ;
        RECT 147.290 128.585 147.570 128.955 ;
        RECT 147.300 128.530 147.560 128.585 ;
        RECT 147.360 128.470 147.500 128.530 ;
        RECT 199.800 125.790 199.940 130.910 ;
        RECT 207.100 130.570 207.360 130.890 ;
        RECT 200.660 127.850 200.920 128.170 ;
        RECT 199.740 125.470 200.000 125.790 ;
        RECT 149.740 123.260 150.540 123.760 ;
        RECT 186.860 123.090 187.120 123.410 ;
        RECT 186.920 117.290 187.060 123.090 ;
        RECT 191.460 120.710 191.720 121.030 ;
        RECT 154.660 116.970 154.920 117.290 ;
        RECT 186.860 116.970 187.120 117.290 ;
        RECT 154.720 111.850 154.860 116.970 ;
        RECT 174.900 112.210 175.160 112.530 ;
        RECT 154.660 111.530 154.920 111.850 ;
        RECT 145.460 109.150 145.720 109.470 ;
        RECT 137.180 106.770 137.440 107.090 ;
        RECT 145.520 107.000 145.660 109.150 ;
        RECT 174.960 107.090 175.100 112.210 ;
        RECT 191.520 111.850 191.660 120.710 ;
        RECT 200.720 112.530 200.860 127.850 ;
        RECT 200.660 112.210 200.920 112.530 ;
        RECT 191.460 111.530 191.720 111.850 ;
        RECT 175.360 109.150 175.620 109.470 ;
        RECT 148.680 107.000 148.940 107.090 ;
        RECT 145.520 106.860 148.940 107.000 ;
        RECT 148.680 106.770 148.940 106.860 ;
        RECT 174.900 106.770 175.160 107.090 ;
        RECT 175.420 107.000 175.560 109.150 ;
        RECT 207.160 107.090 207.300 130.570 ;
        RECT 213.540 128.190 213.800 128.510 ;
        RECT 213.600 112.530 213.740 128.190 ;
        RECT 242.120 125.790 242.260 144.510 ;
        RECT 242.980 127.850 243.240 128.170 ;
        RECT 242.060 125.470 242.320 125.790 ;
        RECT 214.460 123.090 214.720 123.410 ;
        RECT 214.520 121.030 214.660 123.090 ;
        RECT 214.460 120.710 214.720 121.030 ;
        RECT 213.540 112.210 213.800 112.530 ;
        RECT 243.040 107.090 243.180 127.850 ;
        RECT 178.580 107.000 178.840 107.090 ;
        RECT 175.420 106.860 178.840 107.000 ;
        RECT 178.580 106.770 178.840 106.860 ;
        RECT 207.100 106.770 207.360 107.090 ;
        RECT 242.980 106.770 243.240 107.090 ;
        RECT 127.060 85.690 127.320 86.010 ;
        RECT 245.280 74.810 245.540 75.130 ;
        RECT 221.820 74.360 222.080 74.450 ;
        RECT 221.420 74.220 222.080 74.360 ;
        RECT 221.420 69.350 221.560 74.220 ;
        RECT 221.820 74.130 222.080 74.220 ;
        RECT 233.320 71.410 233.580 71.730 ;
        RECT 221.360 69.030 221.620 69.350 ;
        RECT 223.660 55.770 223.920 56.090 ;
        RECT 223.720 31.950 223.860 55.770 ;
        RECT 233.380 50.650 233.520 71.410 ;
        RECT 234.700 66.650 234.960 66.970 ;
        RECT 234.760 56.090 234.900 66.650 ;
        RECT 234.700 55.770 234.960 56.090 ;
        RECT 245.340 50.650 245.480 74.810 ;
        RECT 247.580 66.650 247.840 66.970 ;
        RECT 233.320 50.330 233.580 50.650 ;
        RECT 245.280 50.330 245.540 50.650 ;
        RECT 228.260 47.950 228.520 48.270 ;
        RECT 228.320 46.910 228.460 47.950 ;
        RECT 228.260 46.590 228.520 46.910 ;
        RECT 247.640 37.640 247.780 66.650 ;
        RECT 249.420 46.590 249.680 46.910 ;
        RECT 245.800 37.500 247.780 37.640 ;
        RECT 245.800 36.710 245.940 37.500 ;
        RECT 248.960 37.070 249.220 37.390 ;
        RECT 245.740 36.390 246.000 36.710 ;
        RECT 249.020 31.950 249.160 37.070 ;
        RECT 249.480 36.710 249.620 46.590 ;
        RECT 249.420 36.390 249.680 36.710 ;
        RECT 223.660 31.630 223.920 31.950 ;
        RECT 248.960 31.630 249.220 31.950 ;
      LAYER via2 ;
        RECT 72.770 217.080 73.050 217.360 ;
        RECT 118.770 217.080 119.050 217.360 ;
        RECT 147.290 184.750 147.570 185.030 ;
        RECT 150.000 179.770 150.280 180.050 ;
        RECT 187.770 179.870 188.050 180.150 ;
        RECT 131.380 160.970 131.660 161.250 ;
        RECT 168.620 160.970 168.900 161.250 ;
        RECT 150.000 142.170 150.280 142.450 ;
        RECT 147.290 128.630 147.570 128.910 ;
        RECT 150.000 123.370 150.280 123.650 ;
      LAYER met3 ;
        RECT 72.745 217.370 73.075 217.385 ;
        RECT 118.745 217.370 119.075 217.385 ;
        RECT 72.745 217.070 119.075 217.370 ;
        RECT 72.745 217.055 73.075 217.070 ;
        RECT 118.745 217.055 119.075 217.070 ;
        RECT 147.265 185.040 147.595 185.055 ;
        RECT 148.390 185.040 148.770 185.050 ;
        RECT 147.265 184.740 148.770 185.040 ;
        RECT 147.265 184.725 147.595 184.740 ;
        RECT 148.390 184.730 148.770 184.740 ;
        RECT 149.640 179.610 150.640 180.210 ;
        RECT 187.745 180.170 188.075 180.175 ;
        RECT 187.720 180.160 188.100 180.170 ;
        RECT 187.300 179.860 188.100 180.160 ;
        RECT 187.720 179.850 188.100 179.860 ;
        RECT 187.745 179.845 188.075 179.850 ;
        RECT 131.020 160.810 132.020 161.410 ;
        RECT 168.260 160.810 169.260 161.410 ;
        RECT 149.640 142.010 150.640 142.610 ;
        RECT 147.265 128.920 147.595 128.935 ;
        RECT 148.390 128.920 148.770 128.930 ;
        RECT 147.265 128.620 148.770 128.920 ;
        RECT 147.265 128.605 147.595 128.620 ;
        RECT 148.390 128.610 148.770 128.620 ;
        RECT 149.640 123.210 150.640 123.810 ;
      LAYER via3 ;
        RECT 148.420 184.730 148.740 185.050 ;
        RECT 149.780 179.750 150.100 180.070 ;
        RECT 150.180 179.750 150.500 180.070 ;
        RECT 187.750 179.850 188.070 180.170 ;
        RECT 131.160 160.950 131.480 161.270 ;
        RECT 131.560 160.950 131.880 161.270 ;
        RECT 168.400 160.950 168.720 161.270 ;
        RECT 168.800 160.950 169.120 161.270 ;
        RECT 149.780 142.150 150.100 142.470 ;
        RECT 150.180 142.150 150.500 142.470 ;
        RECT 148.420 128.610 148.740 128.930 ;
        RECT 149.780 123.350 150.100 123.670 ;
        RECT 150.180 123.350 150.500 123.670 ;
      LAYER met4 ;
        RECT 150.330 186.515 151.930 186.610 ;
        RECT 153.930 186.515 155.530 186.610 ;
        RECT 157.530 186.515 159.130 186.610 ;
        RECT 161.130 186.515 162.730 186.610 ;
        RECT 164.730 186.515 166.330 186.610 ;
        RECT 168.330 186.515 169.930 186.610 ;
        RECT 171.930 186.515 173.530 186.610 ;
        RECT 175.530 186.515 177.130 186.610 ;
        RECT 179.130 186.515 180.730 186.610 ;
        RECT 182.730 186.515 184.330 186.610 ;
        RECT 148.415 185.040 148.745 185.055 ;
        RECT 150.330 185.040 151.940 186.515 ;
        RECT 148.415 184.905 151.940 185.040 ;
        RECT 153.925 184.905 155.535 186.515 ;
        RECT 157.520 184.905 159.130 186.515 ;
        RECT 161.115 184.905 162.730 186.515 ;
        RECT 164.710 184.905 166.330 186.515 ;
        RECT 168.305 184.905 169.930 186.515 ;
        RECT 171.900 184.905 173.530 186.515 ;
        RECT 175.495 184.905 177.130 186.515 ;
        RECT 179.090 184.905 180.730 186.515 ;
        RECT 182.685 184.905 184.330 186.515 ;
        RECT 148.415 184.740 151.930 184.905 ;
        RECT 148.415 184.725 148.745 184.740 ;
        RECT 150.330 183.015 151.930 184.740 ;
        RECT 153.930 183.015 155.530 184.905 ;
        RECT 157.530 183.015 159.130 184.905 ;
        RECT 161.130 183.015 162.730 184.905 ;
        RECT 164.730 183.015 166.330 184.905 ;
        RECT 168.330 183.015 169.930 184.905 ;
        RECT 171.930 183.015 173.530 184.905 ;
        RECT 175.530 183.015 177.130 184.905 ;
        RECT 179.130 183.015 180.730 184.905 ;
        RECT 182.730 183.015 184.330 184.905 ;
        RECT 150.330 181.405 151.940 183.015 ;
        RECT 153.925 181.405 155.535 183.015 ;
        RECT 157.520 181.405 159.130 183.015 ;
        RECT 161.115 181.405 162.730 183.015 ;
        RECT 164.710 181.405 166.330 183.015 ;
        RECT 168.305 181.405 169.930 183.015 ;
        RECT 171.900 181.405 173.530 183.015 ;
        RECT 175.495 181.405 177.130 183.015 ;
        RECT 179.090 181.405 180.730 183.015 ;
        RECT 182.685 181.405 184.330 183.015 ;
        RECT 150.330 180.210 151.930 181.405 ;
        RECT 153.930 180.210 155.530 181.405 ;
        RECT 157.530 180.210 159.130 181.405 ;
        RECT 161.130 180.210 162.730 181.405 ;
        RECT 164.730 180.210 166.330 181.405 ;
        RECT 168.330 180.210 169.930 181.405 ;
        RECT 171.930 180.210 173.530 181.405 ;
        RECT 175.530 180.210 177.130 181.405 ;
        RECT 179.130 180.210 180.730 181.405 ;
        RECT 182.730 180.210 184.330 181.405 ;
        RECT 149.640 179.610 185.480 180.210 ;
        RECT 187.745 179.845 188.075 180.175 ;
        RECT 164.990 167.810 165.290 179.610 ;
        RECT 187.760 167.810 188.060 179.845 ;
        RECT 131.710 167.715 133.310 167.810 ;
        RECT 135.310 167.715 136.910 167.810 ;
        RECT 138.910 167.715 140.510 167.810 ;
        RECT 142.510 167.715 144.110 167.810 ;
        RECT 146.110 167.715 147.710 167.810 ;
        RECT 149.710 167.715 151.310 167.810 ;
        RECT 153.310 167.715 154.910 167.810 ;
        RECT 156.910 167.715 158.510 167.810 ;
        RECT 160.510 167.715 162.110 167.810 ;
        RECT 164.110 167.715 165.710 167.810 ;
        RECT 131.710 166.105 133.320 167.715 ;
        RECT 135.305 166.105 136.915 167.715 ;
        RECT 138.900 166.105 140.510 167.715 ;
        RECT 142.495 166.105 144.110 167.715 ;
        RECT 146.090 166.105 147.710 167.715 ;
        RECT 149.685 166.105 151.310 167.715 ;
        RECT 153.280 166.105 154.910 167.715 ;
        RECT 156.875 166.105 158.510 167.715 ;
        RECT 160.470 166.105 162.110 167.715 ;
        RECT 164.065 166.105 165.710 167.715 ;
        RECT 131.710 164.215 133.310 166.105 ;
        RECT 135.310 164.215 136.910 166.105 ;
        RECT 138.910 164.215 140.510 166.105 ;
        RECT 142.510 164.215 144.110 166.105 ;
        RECT 146.110 164.215 147.710 166.105 ;
        RECT 149.710 164.215 151.310 166.105 ;
        RECT 153.310 164.215 154.910 166.105 ;
        RECT 156.910 164.215 158.510 166.105 ;
        RECT 160.510 164.215 162.110 166.105 ;
        RECT 164.110 164.215 165.710 166.105 ;
        RECT 131.710 162.605 133.320 164.215 ;
        RECT 135.305 162.605 136.915 164.215 ;
        RECT 138.900 162.605 140.510 164.215 ;
        RECT 142.495 162.605 144.110 164.215 ;
        RECT 146.090 162.605 147.710 164.215 ;
        RECT 149.685 162.605 151.310 164.215 ;
        RECT 153.280 162.605 154.910 164.215 ;
        RECT 156.875 162.605 158.510 164.215 ;
        RECT 160.470 162.605 162.110 164.215 ;
        RECT 164.065 162.605 165.710 164.215 ;
        RECT 131.710 161.410 133.310 162.605 ;
        RECT 135.310 161.410 136.910 162.605 ;
        RECT 138.910 161.410 140.510 162.605 ;
        RECT 142.510 161.410 144.110 162.605 ;
        RECT 146.110 161.410 147.710 162.605 ;
        RECT 149.710 161.410 151.310 162.605 ;
        RECT 153.310 161.410 154.910 162.605 ;
        RECT 156.910 161.410 158.510 162.605 ;
        RECT 160.510 161.410 162.110 162.605 ;
        RECT 164.110 161.410 165.710 162.605 ;
        RECT 168.950 167.715 170.550 167.810 ;
        RECT 172.550 167.715 174.150 167.810 ;
        RECT 176.150 167.715 177.750 167.810 ;
        RECT 179.750 167.715 181.350 167.810 ;
        RECT 183.350 167.715 184.950 167.810 ;
        RECT 186.950 167.715 188.550 167.810 ;
        RECT 190.550 167.715 192.150 167.810 ;
        RECT 194.150 167.715 195.750 167.810 ;
        RECT 197.750 167.715 199.350 167.810 ;
        RECT 201.350 167.715 202.950 167.810 ;
        RECT 168.950 166.105 170.560 167.715 ;
        RECT 172.545 166.105 174.155 167.715 ;
        RECT 176.140 166.105 177.750 167.715 ;
        RECT 179.735 166.105 181.350 167.715 ;
        RECT 183.330 166.105 184.950 167.715 ;
        RECT 186.925 166.105 188.550 167.715 ;
        RECT 190.520 166.105 192.150 167.715 ;
        RECT 194.115 166.105 195.750 167.715 ;
        RECT 197.710 166.105 199.350 167.715 ;
        RECT 201.305 166.105 202.950 167.715 ;
        RECT 168.950 164.215 170.550 166.105 ;
        RECT 172.550 164.215 174.150 166.105 ;
        RECT 176.150 164.215 177.750 166.105 ;
        RECT 179.750 164.215 181.350 166.105 ;
        RECT 183.350 164.215 184.950 166.105 ;
        RECT 186.950 164.215 188.550 166.105 ;
        RECT 190.550 164.215 192.150 166.105 ;
        RECT 194.150 164.215 195.750 166.105 ;
        RECT 197.750 164.215 199.350 166.105 ;
        RECT 201.350 164.215 202.950 166.105 ;
        RECT 168.950 162.605 170.560 164.215 ;
        RECT 172.545 162.605 174.155 164.215 ;
        RECT 176.140 162.605 177.750 164.215 ;
        RECT 179.735 162.605 181.350 164.215 ;
        RECT 183.330 162.605 184.950 164.215 ;
        RECT 186.925 162.605 188.550 164.215 ;
        RECT 190.520 162.605 192.150 164.215 ;
        RECT 194.115 162.605 195.750 164.215 ;
        RECT 197.710 162.605 199.350 164.215 ;
        RECT 201.305 162.605 202.950 164.215 ;
        RECT 168.950 161.410 170.550 162.605 ;
        RECT 172.550 161.410 174.150 162.605 ;
        RECT 176.150 161.410 177.750 162.605 ;
        RECT 179.750 161.410 181.350 162.605 ;
        RECT 183.350 161.410 184.950 162.605 ;
        RECT 186.950 161.410 188.550 162.605 ;
        RECT 190.550 161.410 192.150 162.605 ;
        RECT 194.150 161.410 195.750 162.605 ;
        RECT 197.750 161.410 199.350 162.605 ;
        RECT 201.350 161.410 202.950 162.605 ;
        RECT 131.020 161.250 166.860 161.410 ;
        RECT 168.260 161.250 204.100 161.410 ;
        RECT 131.020 160.950 204.100 161.250 ;
        RECT 131.020 160.810 166.860 160.950 ;
        RECT 168.260 160.810 204.100 160.950 ;
        RECT 169.130 149.010 169.430 160.810 ;
        RECT 150.330 148.915 151.930 149.010 ;
        RECT 153.930 148.915 155.530 149.010 ;
        RECT 157.530 148.915 159.130 149.010 ;
        RECT 161.130 148.915 162.730 149.010 ;
        RECT 164.730 148.915 166.330 149.010 ;
        RECT 168.330 148.915 169.930 149.010 ;
        RECT 171.930 148.915 173.530 149.010 ;
        RECT 175.530 148.915 177.130 149.010 ;
        RECT 179.130 148.915 180.730 149.010 ;
        RECT 182.730 148.915 184.330 149.010 ;
        RECT 150.330 147.305 151.940 148.915 ;
        RECT 153.925 147.305 155.535 148.915 ;
        RECT 157.520 147.305 159.130 148.915 ;
        RECT 161.115 147.305 162.730 148.915 ;
        RECT 164.710 147.305 166.330 148.915 ;
        RECT 168.305 147.305 169.930 148.915 ;
        RECT 171.900 147.305 173.530 148.915 ;
        RECT 175.495 147.305 177.130 148.915 ;
        RECT 179.090 147.305 180.730 148.915 ;
        RECT 182.685 147.305 184.330 148.915 ;
        RECT 150.330 145.415 151.930 147.305 ;
        RECT 153.930 145.415 155.530 147.305 ;
        RECT 157.530 145.415 159.130 147.305 ;
        RECT 161.130 145.415 162.730 147.305 ;
        RECT 164.730 145.415 166.330 147.305 ;
        RECT 168.330 145.415 169.930 147.305 ;
        RECT 171.930 145.415 173.530 147.305 ;
        RECT 175.530 145.415 177.130 147.305 ;
        RECT 179.130 145.415 180.730 147.305 ;
        RECT 182.730 145.415 184.330 147.305 ;
        RECT 150.330 143.805 151.940 145.415 ;
        RECT 153.925 143.805 155.535 145.415 ;
        RECT 157.520 143.805 159.130 145.415 ;
        RECT 161.115 143.805 162.730 145.415 ;
        RECT 164.710 143.805 166.330 145.415 ;
        RECT 168.305 143.805 169.930 145.415 ;
        RECT 171.900 143.805 173.530 145.415 ;
        RECT 175.495 143.805 177.130 145.415 ;
        RECT 179.090 143.805 180.730 145.415 ;
        RECT 182.685 143.805 184.330 145.415 ;
        RECT 150.330 142.610 151.930 143.805 ;
        RECT 153.930 142.610 155.530 143.805 ;
        RECT 157.530 142.610 159.130 143.805 ;
        RECT 161.130 142.610 162.730 143.805 ;
        RECT 164.730 142.610 166.330 143.805 ;
        RECT 168.330 142.610 169.930 143.805 ;
        RECT 171.930 142.610 173.530 143.805 ;
        RECT 175.530 142.610 177.130 143.805 ;
        RECT 179.130 142.610 180.730 143.805 ;
        RECT 182.730 142.610 184.330 143.805 ;
        RECT 149.640 142.010 185.480 142.610 ;
        RECT 158.090 130.210 158.390 142.010 ;
        RECT 150.330 130.115 151.930 130.210 ;
        RECT 153.930 130.115 155.530 130.210 ;
        RECT 157.530 130.115 159.130 130.210 ;
        RECT 161.130 130.115 162.730 130.210 ;
        RECT 164.730 130.115 166.330 130.210 ;
        RECT 168.330 130.115 169.930 130.210 ;
        RECT 171.930 130.115 173.530 130.210 ;
        RECT 175.530 130.115 177.130 130.210 ;
        RECT 179.130 130.115 180.730 130.210 ;
        RECT 182.730 130.115 184.330 130.210 ;
        RECT 148.415 128.920 148.745 128.935 ;
        RECT 150.330 128.920 151.940 130.115 ;
        RECT 148.415 128.620 151.940 128.920 ;
        RECT 148.415 128.605 148.745 128.620 ;
        RECT 150.330 128.505 151.940 128.620 ;
        RECT 153.925 128.505 155.535 130.115 ;
        RECT 157.520 128.505 159.130 130.115 ;
        RECT 161.115 128.505 162.730 130.115 ;
        RECT 164.710 128.505 166.330 130.115 ;
        RECT 168.305 128.505 169.930 130.115 ;
        RECT 171.900 128.505 173.530 130.115 ;
        RECT 175.495 128.505 177.130 130.115 ;
        RECT 179.090 128.505 180.730 130.115 ;
        RECT 182.685 128.505 184.330 130.115 ;
        RECT 150.330 126.615 151.930 128.505 ;
        RECT 153.930 126.615 155.530 128.505 ;
        RECT 157.530 126.615 159.130 128.505 ;
        RECT 161.130 126.615 162.730 128.505 ;
        RECT 164.730 126.615 166.330 128.505 ;
        RECT 168.330 126.615 169.930 128.505 ;
        RECT 171.930 126.615 173.530 128.505 ;
        RECT 175.530 126.615 177.130 128.505 ;
        RECT 179.130 126.615 180.730 128.505 ;
        RECT 182.730 126.615 184.330 128.505 ;
        RECT 150.330 125.005 151.940 126.615 ;
        RECT 153.925 125.005 155.535 126.615 ;
        RECT 157.520 125.005 159.130 126.615 ;
        RECT 161.115 125.005 162.730 126.615 ;
        RECT 164.710 125.005 166.330 126.615 ;
        RECT 168.305 125.005 169.930 126.615 ;
        RECT 171.900 125.005 173.530 126.615 ;
        RECT 175.495 125.005 177.130 126.615 ;
        RECT 179.090 125.005 180.730 126.615 ;
        RECT 182.685 125.005 184.330 126.615 ;
        RECT 150.330 123.810 151.930 125.005 ;
        RECT 153.930 123.810 155.530 125.005 ;
        RECT 157.530 123.810 159.130 125.005 ;
        RECT 161.130 123.810 162.730 125.005 ;
        RECT 164.730 123.810 166.330 125.005 ;
        RECT 168.330 123.810 169.930 125.005 ;
        RECT 171.930 123.810 173.530 125.005 ;
        RECT 175.530 123.810 177.130 125.005 ;
        RECT 179.130 123.810 180.730 125.005 ;
        RECT 182.730 123.810 184.330 125.005 ;
        RECT 149.640 123.210 185.480 123.810 ;
  END
END bgr_0
END LIBRARY

