* NGSPICE file created from sky130_asc_pfet_01v8_lvt_6.ext - technology: sky130A

.subckt sky130_asc_pfet_01v8_lvt_6 GATE SOURCE DRAIN VPWR VGND
X0 DRAIN GATE SOURCE w_130_1000# sky130_fd_pr__pfet_01v8_lvt ad=7.482e+12p pd=5.392e+07u as=5.6115e+12p ps=4.044e+07u w=6.45e+06u l=2e+06u
X1 SOURCE GATE DRAIN w_130_1000# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=6.45e+06u l=2e+06u
X2 SOURCE GATE DRAIN w_130_1000# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=6.45e+06u l=2e+06u
X3 DRAIN GATE SOURCE w_130_1000# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=6.45e+06u l=2e+06u
X4 SOURCE GATE DRAIN w_130_1000# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=6.45e+06u l=2e+06u
X5 DRAIN GATE SOURCE w_130_1000# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=6.45e+06u l=2e+06u
.ends

