magic
tech sky130A
magscale 1 2
timestamp 1652753014
<< pwell >>
rect 90 30 704 1426
<< nmoslvt >>
rect 246 600 646 1400
<< ndiff >>
rect 188 1388 246 1400
rect 188 612 200 1388
rect 234 612 246 1388
rect 188 600 246 612
rect 646 1388 704 1400
rect 646 612 658 1388
rect 692 612 704 1388
rect 646 600 704 612
<< ndiffc >>
rect 200 612 234 1388
rect 658 612 692 1388
<< psubdiff >>
rect 128 160 168 200
rect 128 80 168 120
<< psubdiffcont >>
rect 128 120 168 160
<< poly >>
rect 246 1400 646 1426
rect 246 574 646 600
rect 394 224 514 574
rect 268 204 704 224
rect 268 144 358 204
rect 418 144 704 204
rect 268 124 704 144
<< polycont >>
rect 358 144 418 204
<< locali >>
rect 90 1850 358 1910
rect 418 1850 704 1910
rect 188 1690 704 1750
rect 657 1404 691 1690
rect 200 1388 234 1404
rect 199 612 200 654
rect 657 1388 692 1404
rect 657 1386 658 1388
rect 199 596 234 612
rect 658 596 692 612
rect 199 430 233 596
rect 188 370 704 430
rect 118 160 178 240
rect 118 120 128 160
rect 168 120 178 160
rect 268 144 358 204
rect 418 144 704 204
rect 118 30 178 120
rect 90 -30 358 30
rect 418 -30 704 30
<< viali >>
rect 358 1850 418 1910
rect 200 612 234 1388
rect 658 612 692 1388
rect 358 -30 418 30
<< metal1 >>
rect 90 1910 704 1940
rect 90 1850 358 1910
rect 418 1850 704 1910
rect 90 1820 704 1850
rect 194 1388 240 1400
rect 194 612 200 1388
rect 234 612 240 1388
rect 194 600 240 612
rect 652 1388 698 1400
rect 652 612 658 1388
rect 692 612 698 1388
rect 652 600 698 612
rect 90 30 704 60
rect 90 -30 358 30
rect 418 -30 704 30
rect 90 -60 704 -30
<< labels >>
flabel metal1 188 1850 248 1910 1 FreeSans 800 0 0 0 VPWR
port 4 n power bidirectional
flabel metal1 188 -30 248 30 1 FreeSans 800 0 0 0 VGND
port 5 n ground bidirectional
flabel locali 644 1690 704 1750 1 FreeSans 800 0 0 0 SOURCE
port 2 n default bidirectional
flabel locali 644 370 704 430 1 FreeSans 800 0 0 0 DRAIN
port 3 n default bidirectional
flabel locali 644 144 704 204 1 FreeSans 800 0 0 0 GATE
port 1 n default bidirectional
<< properties >>
string FIXED_BBOX 0 0 794 1880
string LEFclass CORE
string LEFsite unitasc
<< end >>
