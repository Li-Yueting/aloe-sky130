* NGSPICE file created from bgr_top.ext - technology: sky130A

.subckt sky130_asc_res_xhigh_po_2p85_1 Rin Rout VPWR VGND a_2148_115#
X0 Rin a_2148_115# VGND sky130_fd_pr__res_xhigh_po w=2.85e+06u l=7.88e+06u
X1 Rout a_2148_115# VGND sky130_fd_pr__res_xhigh_po w=2.85e+06u l=7.88e+06u
C0 VPWR Rin 0.17fF
C1 a_2148_115# VPWR 0.17fF
C2 Rout Rin 0.12fF
C3 VPWR VGND 2.31fF
C4 Rout VGND 1.26fF
C5 Rin VGND 0.78fF
C6 a_2148_115# VGND 2.70fF
.ends

.subckt sky130_asc_pfet_01v8_lvt_60 GATE SOURCE DRAIN VGND VPWR VSUBS
X0 DRAIN GATE SOURCE VPWR sky130_fd_pr__pfet_01v8_lvt ad=5.79855e+13p pd=4.1788e+08u as=5.6115e+13p ps=4.044e+08u w=6.45e+06u l=2e+06u
X1 SOURCE GATE DRAIN VPWR sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=6.45e+06u l=2e+06u
X2 DRAIN GATE SOURCE VPWR sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=6.45e+06u l=2e+06u
X3 SOURCE GATE DRAIN VPWR sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=6.45e+06u l=2e+06u
X4 DRAIN GATE SOURCE VPWR sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=6.45e+06u l=2e+06u
X5 DRAIN GATE SOURCE VPWR sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=6.45e+06u l=2e+06u
X6 DRAIN GATE SOURCE VPWR sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=6.45e+06u l=2e+06u
X7 DRAIN GATE SOURCE VPWR sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=6.45e+06u l=2e+06u
X8 DRAIN GATE SOURCE VPWR sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=6.45e+06u l=2e+06u
X9 SOURCE GATE DRAIN VPWR sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=6.45e+06u l=2e+06u
X10 DRAIN GATE SOURCE VPWR sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=6.45e+06u l=2e+06u
X11 SOURCE GATE DRAIN VPWR sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=6.45e+06u l=2e+06u
X12 SOURCE GATE DRAIN VPWR sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=6.45e+06u l=2e+06u
X13 DRAIN GATE SOURCE VPWR sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=6.45e+06u l=2e+06u
X14 DRAIN GATE SOURCE VPWR sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=6.45e+06u l=2e+06u
X15 SOURCE GATE DRAIN VPWR sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=6.45e+06u l=2e+06u
X16 SOURCE GATE DRAIN VPWR sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=6.45e+06u l=2e+06u
X17 DRAIN GATE SOURCE VPWR sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=6.45e+06u l=2e+06u
X18 SOURCE GATE DRAIN VPWR sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=6.45e+06u l=2e+06u
X19 DRAIN GATE SOURCE VPWR sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=6.45e+06u l=2e+06u
X20 SOURCE GATE DRAIN VPWR sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=6.45e+06u l=2e+06u
X21 DRAIN GATE SOURCE VPWR sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=6.45e+06u l=2e+06u
X22 SOURCE GATE DRAIN VPWR sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=6.45e+06u l=2e+06u
X23 DRAIN GATE SOURCE VPWR sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=6.45e+06u l=2e+06u
X24 SOURCE GATE DRAIN VPWR sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=6.45e+06u l=2e+06u
X25 DRAIN GATE SOURCE VPWR sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=6.45e+06u l=2e+06u
X26 SOURCE GATE DRAIN VPWR sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=6.45e+06u l=2e+06u
X27 SOURCE GATE DRAIN VPWR sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=6.45e+06u l=2e+06u
X28 DRAIN GATE SOURCE VPWR sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=6.45e+06u l=2e+06u
X29 SOURCE GATE DRAIN VPWR sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=6.45e+06u l=2e+06u
X30 DRAIN GATE SOURCE VPWR sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=6.45e+06u l=2e+06u
X31 SOURCE GATE DRAIN VPWR sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=6.45e+06u l=2e+06u
X32 DRAIN GATE SOURCE VPWR sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=6.45e+06u l=2e+06u
X33 SOURCE GATE DRAIN VPWR sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=6.45e+06u l=2e+06u
X34 DRAIN GATE SOURCE VPWR sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=6.45e+06u l=2e+06u
X35 SOURCE GATE DRAIN VPWR sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=6.45e+06u l=2e+06u
X36 DRAIN GATE SOURCE VPWR sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=6.45e+06u l=2e+06u
X37 SOURCE GATE DRAIN VPWR sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=6.45e+06u l=2e+06u
X38 DRAIN GATE SOURCE VPWR sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=6.45e+06u l=2e+06u
X39 SOURCE GATE DRAIN VPWR sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=6.45e+06u l=2e+06u
X40 SOURCE GATE DRAIN VPWR sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=6.45e+06u l=2e+06u
X41 DRAIN GATE SOURCE VPWR sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=6.45e+06u l=2e+06u
X42 DRAIN GATE SOURCE VPWR sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=6.45e+06u l=2e+06u
X43 DRAIN GATE SOURCE VPWR sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=6.45e+06u l=2e+06u
X44 SOURCE GATE DRAIN VPWR sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=6.45e+06u l=2e+06u
X45 SOURCE GATE DRAIN VPWR sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=6.45e+06u l=2e+06u
X46 DRAIN GATE SOURCE VPWR sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=6.45e+06u l=2e+06u
X47 SOURCE GATE DRAIN VPWR sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=6.45e+06u l=2e+06u
X48 SOURCE GATE DRAIN VPWR sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=6.45e+06u l=2e+06u
X49 SOURCE GATE DRAIN VPWR sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=6.45e+06u l=2e+06u
X50 DRAIN GATE SOURCE VPWR sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=6.45e+06u l=2e+06u
X51 SOURCE GATE DRAIN VPWR sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=6.45e+06u l=2e+06u
X52 SOURCE GATE DRAIN VPWR sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=6.45e+06u l=2e+06u
X53 SOURCE GATE DRAIN VPWR sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=6.45e+06u l=2e+06u
X54 DRAIN GATE SOURCE VPWR sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=6.45e+06u l=2e+06u
X55 SOURCE GATE DRAIN VPWR sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=6.45e+06u l=2e+06u
X56 DRAIN GATE SOURCE VPWR sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=6.45e+06u l=2e+06u
X57 DRAIN GATE SOURCE VPWR sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=6.45e+06u l=2e+06u
X58 SOURCE GATE DRAIN VPWR sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=6.45e+06u l=2e+06u
X59 DRAIN GATE SOURCE VPWR sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=6.45e+06u l=2e+06u
C0 SOURCE VGND 0.32fF
C1 DRAIN VGND 5.28fF
C2 VPWR GATE 27.32fF
C3 SOURCE DRAIN 1.25fF
C4 GATE VGND 12.31fF
C5 VPWR SOURCE 22.83fF
C6 VPWR DRAIN 1.83fF
C7 SOURCE GATE 0.18fF
C8 GATE DRAIN 25.46fF
C9 VGND VSUBS 25.41fF
C10 SOURCE VSUBS 0.00fF
C11 DRAIN VSUBS 9.62fF
C12 GATE VSUBS 30.27fF
C13 VPWR VSUBS 142.65fF
.ends

.subckt sky130_asc_pnp_05v5_W3p40L3p40_7 Emitter Base Collector VPWR VGND
X0 Collector Base Emitter sky130_fd_pr__pnp_05v5_W3p40L3p40
X1 Collector Base Emitter sky130_fd_pr__pnp_05v5_W3p40L3p40
X2 Collector Base Emitter sky130_fd_pr__pnp_05v5_W3p40L3p40
X3 Collector Base Emitter sky130_fd_pr__pnp_05v5_W3p40L3p40
X4 Collector Base Emitter sky130_fd_pr__pnp_05v5_W3p40L3p40
X5 Collector Base Emitter sky130_fd_pr__pnp_05v5_W3p40L3p40
X6 Collector Base Emitter sky130_fd_pr__pnp_05v5_W3p40L3p40
C0 Base Emitter 18.67fF
C1 VGND Collector 9.81fF
C2 VPWR Collector 11.49fF
C3 Emitter Collector 9.06fF
C4 Base Collector 28.86fF
.ends

.subckt sky130_asc_res_xhigh_po_2p85_2 Rin Rout VPWR a_2723_115# VGND
X0 Rout a_2723_115# VGND sky130_fd_pr__res_xhigh_po w=2.85e+06u l=1.075e+07u
X1 Rin a_2723_115# VGND sky130_fd_pr__res_xhigh_po w=2.85e+06u l=1.075e+07u
C0 Rin Rout 0.12fF
C1 Rin VPWR 0.17fF
C2 a_2723_115# VPWR 0.17fF
C3 VPWR VGND 2.83fF
C4 Rout VGND 1.26fF
C5 Rin VGND 0.78fF
C6 a_2723_115# VGND 2.70fF
.ends

.subckt sky130_asc_pfet_01v8_lvt_12 GATE SOURCE DRAIN VGND VPWR VSUBS
X0 SOURCE GATE DRAIN VPWR sky130_fd_pr__pfet_01v8_lvt ad=1.1223e+13p pd=8.088e+07u as=1.30935e+13p ps=9.436e+07u w=6.45e+06u l=2e+06u
X1 DRAIN GATE SOURCE VPWR sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=6.45e+06u l=2e+06u
X2 DRAIN GATE SOURCE VPWR sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=6.45e+06u l=2e+06u
X3 SOURCE GATE DRAIN VPWR sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=6.45e+06u l=2e+06u
X4 SOURCE GATE DRAIN VPWR sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=6.45e+06u l=2e+06u
X5 DRAIN GATE SOURCE VPWR sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=6.45e+06u l=2e+06u
X6 SOURCE GATE DRAIN VPWR sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=6.45e+06u l=2e+06u
X7 DRAIN GATE SOURCE VPWR sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=6.45e+06u l=2e+06u
X8 DRAIN GATE SOURCE VPWR sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=6.45e+06u l=2e+06u
X9 SOURCE GATE DRAIN VPWR sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=6.45e+06u l=2e+06u
X10 SOURCE GATE DRAIN VPWR sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=6.45e+06u l=2e+06u
X11 DRAIN GATE SOURCE VPWR sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=6.45e+06u l=2e+06u
C0 GATE VGND 2.51fF
C1 SOURCE DRAIN 0.26fF
C2 VPWR GATE 5.46fF
C3 SOURCE VGND 0.06fF
C4 DRAIN VGND 1.08fF
C5 SOURCE VPWR 4.54fF
C6 SOURCE GATE 0.04fF
C7 VPWR DRAIN 0.42fF
C8 DRAIN GATE 5.17fF
C9 VGND VSUBS 5.31fF
C10 SOURCE VSUBS 0.00fF
C11 DRAIN VSUBS 1.99fF
C12 GATE VSUBS 6.20fF
C13 VPWR VSUBS 29.52fF
.ends

.subckt sky130_asc_nfet_01v8_lvt_9 GATE SOURCE DRAIN VPWR VGND
X0 SOURCE GATE DRAIN VGND sky130_fd_pr__nfet_01v8_lvt ad=4.35e+12p pd=3.29e+07u as=4.35e+12p ps=3.29e+07u w=3e+06u l=2e+06u
X1 SOURCE GATE DRAIN VGND sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=2e+06u
X2 DRAIN GATE SOURCE VGND sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=2e+06u
X3 SOURCE GATE DRAIN VGND sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=2e+06u
X4 SOURCE GATE DRAIN VGND sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=2e+06u
X5 DRAIN GATE SOURCE VGND sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=2e+06u
X6 DRAIN GATE SOURCE VGND sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=2e+06u
X7 SOURCE GATE DRAIN VGND sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=2e+06u
X8 DRAIN GATE SOURCE VGND sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=2e+06u
C0 VPWR SOURCE 1.38fF
C1 DRAIN SOURCE 0.04fF
C2 DRAIN GATE 2.90fF
C3 GATE SOURCE 0.01fF
C4 VPWR VGND 3.99fF
C5 SOURCE VGND 2.86fF
C6 DRAIN VGND 2.50fF
C7 GATE VGND 10.91fF
.ends

.subckt sky130_asc_pfet_01v8_lvt_6 GATE SOURCE DRAIN VGND VPWR VSUBS
X0 SOURCE GATE DRAIN VPWR sky130_fd_pr__pfet_01v8_lvt ad=5.6115e+12p pd=4.044e+07u as=7.482e+12p ps=5.392e+07u w=6.45e+06u l=2e+06u
X1 SOURCE GATE DRAIN VPWR sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=6.45e+06u l=2e+06u
X2 DRAIN GATE SOURCE VPWR sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=6.45e+06u l=2e+06u
X3 DRAIN GATE SOURCE VPWR sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=6.45e+06u l=2e+06u
X4 SOURCE GATE DRAIN VPWR sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=6.45e+06u l=2e+06u
X5 DRAIN GATE SOURCE VPWR sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=6.45e+06u l=2e+06u
C0 GATE SOURCE 0.02fF
C1 VPWR GATE 2.73fF
C2 SOURCE VGND 0.03fF
C3 DRAIN GATE 2.63fF
C4 DRAIN VGND 0.56fF
C5 VPWR SOURCE 2.27fF
C6 DRAIN SOURCE 0.14fF
C7 GATE VGND 1.28fF
C8 VPWR DRAIN 0.24fF
C9 VGND VSUBS 2.79fF
C10 SOURCE VSUBS 0.00fF
C11 DRAIN VSUBS 1.04fF
C12 GATE VSUBS 3.19fF
C13 VPWR VSUBS 15.38fF
.ends

.subckt sky130_asc_pnp_05v5_W3p40L3p40_1 Emitter Base Collector VPWR VGND
X0 Collector Base Emitter sky130_fd_pr__pnp_05v5_W3p40L3p40
C0 Base Emitter 1.55fF
C1 VGND Collector 1.50fF
C2 VPWR Collector 1.46fF
C3 Emitter Collector 0.40fF
C4 Base Collector 3.33fF
.ends

.subckt sky130_asc_cap_mim_m3_1 Cin Cout VPWR VGND VSUBS
X0 Cout Cin sky130_fd_pr__cap_mim_m3_1 l=2e+06u w=2e+06u
X1 Cout Cin sky130_fd_pr__cap_mim_m3_1 l=2e+06u w=2e+06u
X2 Cout Cin sky130_fd_pr__cap_mim_m3_1 l=2e+06u w=2e+06u
X3 Cout Cin sky130_fd_pr__cap_mim_m3_1 l=2e+06u w=2e+06u
X4 Cout Cin sky130_fd_pr__cap_mim_m3_1 l=2e+06u w=2e+06u
X5 Cout Cin sky130_fd_pr__cap_mim_m3_1 l=2e+06u w=2e+06u
X6 Cout Cin sky130_fd_pr__cap_mim_m3_1 l=2e+06u w=2e+06u
X7 Cout Cin sky130_fd_pr__cap_mim_m3_1 l=2e+06u w=2e+06u
X8 Cout Cin sky130_fd_pr__cap_mim_m3_1 l=2e+06u w=2e+06u
X9 Cout Cin sky130_fd_pr__cap_mim_m3_1 l=2e+06u w=2e+06u
X10 Cout Cin sky130_fd_pr__cap_mim_m3_1 l=2e+06u w=2e+06u
X11 Cout Cin sky130_fd_pr__cap_mim_m3_1 l=2e+06u w=2e+06u
X12 Cout Cin sky130_fd_pr__cap_mim_m3_1 l=2e+06u w=2e+06u
X13 Cout Cin sky130_fd_pr__cap_mim_m3_1 l=2e+06u w=2e+06u
X14 Cout Cin sky130_fd_pr__cap_mim_m3_1 l=2e+06u w=2e+06u
X15 Cout Cin sky130_fd_pr__cap_mim_m3_1 l=2e+06u w=2e+06u
X16 Cout Cin sky130_fd_pr__cap_mim_m3_1 l=2e+06u w=2e+06u
X17 Cout Cin sky130_fd_pr__cap_mim_m3_1 l=2e+06u w=2e+06u
X18 Cout Cin sky130_fd_pr__cap_mim_m3_1 l=2e+06u w=2e+06u
X19 Cout Cin sky130_fd_pr__cap_mim_m3_1 l=2e+06u w=2e+06u
C0 Cout Cin 28.31fF
C1 Cout VSUBS 2.81fF
C2 Cin VSUBS 6.38fF
C3 VGND VSUBS 6.63fF
C4 VPWR VSUBS 6.63fF
.ends

.subckt sky130_asc_pnp_05v5_W3p40L3p40_8 Emitter Base Collector VPWR VGND
X0 Collector Base Emitter sky130_fd_pr__pnp_05v5_W3p40L3p40
X1 Collector Base Emitter sky130_fd_pr__pnp_05v5_W3p40L3p40
X2 Collector Base Emitter sky130_fd_pr__pnp_05v5_W3p40L3p40
X3 Collector Base Emitter sky130_fd_pr__pnp_05v5_W3p40L3p40
X4 Collector Base Emitter sky130_fd_pr__pnp_05v5_W3p40L3p40
X5 Collector Base Emitter sky130_fd_pr__pnp_05v5_W3p40L3p40
X6 Collector Base Emitter sky130_fd_pr__pnp_05v5_W3p40L3p40
X7 Collector Base Emitter sky130_fd_pr__pnp_05v5_W3p40L3p40
C0 Base Emitter 21.50fF
C1 VGND Collector 11.20fF
C2 VPWR Collector 13.12fF
C3 Emitter Collector 10.49fF
C4 Base Collector 33.06fF
.ends

.subckt sky130_asc_nfet_01v8_lvt_1 GATE SOURCE DRAIN VPWR VGND
X0 SOURCE GATE DRAIN VGND sky130_fd_pr__nfet_01v8_lvt ad=1.16e+12p pd=8.58e+06u as=1.16e+12p ps=8.58e+06u w=4e+06u l=2e+06u
C0 VPWR SOURCE 0.17fF
C1 GATE DRAIN 0.18fF
C2 GATE SOURCE 0.00fF
C3 DRAIN SOURCE 0.01fF
C4 VPWR VGND 0.64fF
C5 SOURCE VGND 0.40fF
C6 DRAIN VGND 0.34fF
C7 GATE VGND 1.34fF
.ends

.subckt bgr_top porst va vb vbg VSS VDD
Xsky130_asc_res_xhigh_po_2p85_1_7 sky130_asc_res_xhigh_po_2p85_1_7/Rin sky130_asc_res_xhigh_po_2p85_1_6/Rin
+ VDD VSS sky130_asc_res_xhigh_po_2p85_1_7/a_2148_115# sky130_asc_res_xhigh_po_2p85_1
Xsky130_asc_res_xhigh_po_2p85_1_8 vbg sky130_asc_res_xhigh_po_2p85_1_7/Rin VDD VSS
+ sky130_asc_res_xhigh_po_2p85_1_8/a_2148_115# sky130_asc_res_xhigh_po_2p85_1
Xsky130_asc_res_xhigh_po_2p85_1_9 sky130_asc_res_xhigh_po_2p85_1_9/Rin sky130_asc_res_xhigh_po_2p85_2_0/Rin
+ VDD VSS sky130_asc_res_xhigh_po_2p85_1_9/a_2148_115# sky130_asc_res_xhigh_po_2p85_1
Xsky130_asc_pfet_01v8_lvt_60_0 sky130_asc_cap_mim_m3_1_4/Cout VDD vbg VSS VDD VSS
+ sky130_asc_pfet_01v8_lvt_60
Xsky130_asc_pfet_01v8_lvt_60_1 sky130_asc_cap_mim_m3_1_4/Cout VDD vb VSS VDD VSS sky130_asc_pfet_01v8_lvt_60
Xsky130_asc_pfet_01v8_lvt_60_2 sky130_asc_cap_mim_m3_1_4/Cout VDD va VSS VDD VSS sky130_asc_pfet_01v8_lvt_60
Xsky130_asc_res_xhigh_po_2p85_1_30 va sky130_asc_res_xhigh_po_2p85_1_29/Rin VDD VSS
+ sky130_asc_res_xhigh_po_2p85_1_30/a_2148_115# sky130_asc_res_xhigh_po_2p85_1
Xsky130_asc_res_xhigh_po_2p85_1_20 vb sky130_asc_res_xhigh_po_2p85_1_19/Rin VDD VSS
+ sky130_asc_res_xhigh_po_2p85_1_20/a_2148_115# sky130_asc_res_xhigh_po_2p85_1
Xsky130_asc_pnp_05v5_W3p40L3p40_7_0 sky130_asc_res_xhigh_po_2p85_1_19/Rout VSS VSS
+ VDD VSS sky130_asc_pnp_05v5_W3p40L3p40_7
Xsky130_asc_res_xhigh_po_2p85_1_10 sky130_asc_res_xhigh_po_2p85_1_10/Rin sky130_asc_res_xhigh_po_2p85_1_9/Rin
+ VDD VSS sky130_asc_res_xhigh_po_2p85_1_10/a_2148_115# sky130_asc_res_xhigh_po_2p85_1
Xsky130_asc_res_xhigh_po_2p85_1_21 sky130_asc_res_xhigh_po_2p85_1_21/Rin sky130_asc_res_xhigh_po_2p85_2_1/Rin
+ VDD VSS sky130_asc_res_xhigh_po_2p85_1_21/a_2148_115# sky130_asc_res_xhigh_po_2p85_1
Xsky130_asc_res_xhigh_po_2p85_2_0 sky130_asc_res_xhigh_po_2p85_2_0/Rin VSS VDD sky130_asc_res_xhigh_po_2p85_2_0/a_2723_115#
+ VSS sky130_asc_res_xhigh_po_2p85_2
Xsky130_asc_res_xhigh_po_2p85_1_11 sky130_asc_res_xhigh_po_2p85_1_11/Rin sky130_asc_res_xhigh_po_2p85_1_10/Rin
+ VDD VSS sky130_asc_res_xhigh_po_2p85_1_11/a_2148_115# sky130_asc_res_xhigh_po_2p85_1
Xsky130_asc_res_xhigh_po_2p85_1_22 sky130_asc_res_xhigh_po_2p85_1_22/Rin sky130_asc_res_xhigh_po_2p85_1_21/Rin
+ VDD VSS sky130_asc_res_xhigh_po_2p85_1_22/a_2148_115# sky130_asc_res_xhigh_po_2p85_1
Xsky130_asc_res_xhigh_po_2p85_2_1 sky130_asc_res_xhigh_po_2p85_2_1/Rin VSS VDD sky130_asc_res_xhigh_po_2p85_2_1/a_2723_115#
+ VSS sky130_asc_res_xhigh_po_2p85_2
Xsky130_asc_res_xhigh_po_2p85_1_12 sky130_asc_res_xhigh_po_2p85_1_12/Rin sky130_asc_res_xhigh_po_2p85_1_11/Rin
+ VDD VSS sky130_asc_res_xhigh_po_2p85_1_12/a_2148_115# sky130_asc_res_xhigh_po_2p85_1
Xsky130_asc_res_xhigh_po_2p85_1_23 sky130_asc_res_xhigh_po_2p85_1_23/Rin sky130_asc_res_xhigh_po_2p85_1_22/Rin
+ VDD VSS sky130_asc_res_xhigh_po_2p85_1_23/a_2148_115# sky130_asc_res_xhigh_po_2p85_1
Xsky130_asc_res_xhigh_po_2p85_1_13 sky130_asc_res_xhigh_po_2p85_1_13/Rin sky130_asc_res_xhigh_po_2p85_1_12/Rin
+ VDD VSS sky130_asc_res_xhigh_po_2p85_1_13/a_2148_115# sky130_asc_res_xhigh_po_2p85_1
Xsky130_asc_res_xhigh_po_2p85_1_24 sky130_asc_res_xhigh_po_2p85_1_24/Rin sky130_asc_res_xhigh_po_2p85_1_23/Rin
+ VDD VSS sky130_asc_res_xhigh_po_2p85_1_24/a_2148_115# sky130_asc_res_xhigh_po_2p85_1
Xsky130_asc_pfet_01v8_lvt_12_0 VDD VDD va VSS VDD VSS sky130_asc_pfet_01v8_lvt_12
Xsky130_asc_res_xhigh_po_2p85_1_14 sky130_asc_res_xhigh_po_2p85_1_14/Rin sky130_asc_res_xhigh_po_2p85_1_13/Rin
+ VDD VSS sky130_asc_res_xhigh_po_2p85_1_14/a_2148_115# sky130_asc_res_xhigh_po_2p85_1
Xsky130_asc_res_xhigh_po_2p85_1_25 sky130_asc_res_xhigh_po_2p85_1_25/Rin sky130_asc_res_xhigh_po_2p85_1_24/Rin
+ VDD VSS sky130_asc_res_xhigh_po_2p85_1_25/a_2148_115# sky130_asc_res_xhigh_po_2p85_1
Xsky130_asc_pfet_01v8_lvt_12_1 sky130_asc_cap_mim_m3_1_4/Cout VDD sky130_asc_nfet_01v8_lvt_1_1/GATE
+ VSS VDD VSS sky130_asc_pfet_01v8_lvt_12
Xsky130_asc_res_xhigh_po_2p85_1_15 sky130_asc_res_xhigh_po_2p85_1_15/Rin sky130_asc_res_xhigh_po_2p85_1_14/Rin
+ VDD VSS sky130_asc_res_xhigh_po_2p85_1_15/a_2148_115# sky130_asc_res_xhigh_po_2p85_1
Xsky130_asc_res_xhigh_po_2p85_1_26 sky130_asc_res_xhigh_po_2p85_1_26/Rin sky130_asc_res_xhigh_po_2p85_1_25/Rin
+ VDD VSS sky130_asc_res_xhigh_po_2p85_1_26/a_2148_115# sky130_asc_res_xhigh_po_2p85_1
Xsky130_asc_res_xhigh_po_2p85_1_16 sky130_asc_res_xhigh_po_2p85_1_18/Rin sky130_asc_res_xhigh_po_2p85_1_15/Rin
+ VDD VSS sky130_asc_res_xhigh_po_2p85_1_16/a_2148_115# sky130_asc_res_xhigh_po_2p85_1
Xsky130_asc_res_xhigh_po_2p85_1_27 sky130_asc_res_xhigh_po_2p85_1_27/Rin sky130_asc_res_xhigh_po_2p85_1_26/Rin
+ VDD VSS sky130_asc_res_xhigh_po_2p85_1_27/a_2148_115# sky130_asc_res_xhigh_po_2p85_1
Xsky130_asc_res_xhigh_po_2p85_1_17 sky130_asc_res_xhigh_po_2p85_1_17/Rin vb VDD VSS
+ sky130_asc_res_xhigh_po_2p85_1_17/a_2148_115# sky130_asc_res_xhigh_po_2p85_1
Xsky130_asc_res_xhigh_po_2p85_1_28 sky130_asc_res_xhigh_po_2p85_1_28/Rin sky130_asc_res_xhigh_po_2p85_1_27/Rin
+ VDD VSS sky130_asc_res_xhigh_po_2p85_1_28/a_2148_115# sky130_asc_res_xhigh_po_2p85_1
Xsky130_asc_nfet_01v8_lvt_9_0 porst VSS sky130_asc_cap_mim_m3_1_4/Cout VDD VSS sky130_asc_nfet_01v8_lvt_9
Xsky130_asc_res_xhigh_po_2p85_1_18 sky130_asc_res_xhigh_po_2p85_1_18/Rin sky130_asc_res_xhigh_po_2p85_1_17/Rin
+ VDD VSS sky130_asc_res_xhigh_po_2p85_1_18/a_2148_115# sky130_asc_res_xhigh_po_2p85_1
Xsky130_asc_res_xhigh_po_2p85_1_29 sky130_asc_res_xhigh_po_2p85_1_29/Rin sky130_asc_res_xhigh_po_2p85_1_28/Rin
+ VDD VSS sky130_asc_res_xhigh_po_2p85_1_29/a_2148_115# sky130_asc_res_xhigh_po_2p85_1
Xsky130_asc_pfet_01v8_lvt_6_0 sky130_asc_pfet_01v8_lvt_6_1/GATE VDD sky130_asc_cap_mim_m3_1_4/Cout
+ VSS VDD VSS sky130_asc_pfet_01v8_lvt_6
Xsky130_asc_nfet_01v8_lvt_9_1 va sky130_asc_nfet_01v8_lvt_1_1/DRAIN sky130_asc_cap_mim_m3_1_4/Cout
+ VDD VSS sky130_asc_nfet_01v8_lvt_9
Xsky130_asc_res_xhigh_po_2p85_1_19 sky130_asc_res_xhigh_po_2p85_1_19/Rin sky130_asc_res_xhigh_po_2p85_1_19/Rout
+ VDD VSS sky130_asc_res_xhigh_po_2p85_1_19/a_2148_115# sky130_asc_res_xhigh_po_2p85_1
Xsky130_asc_pfet_01v8_lvt_6_1 sky130_asc_pfet_01v8_lvt_6_1/GATE VDD sky130_asc_pfet_01v8_lvt_6_1/GATE
+ VSS VDD VSS sky130_asc_pfet_01v8_lvt_6
Xsky130_asc_pnp_05v5_W3p40L3p40_1_0 va VSS VSS VDD VSS sky130_asc_pnp_05v5_W3p40L3p40_1
Xsky130_asc_nfet_01v8_lvt_9_2 vb sky130_asc_nfet_01v8_lvt_1_1/DRAIN sky130_asc_pfet_01v8_lvt_6_1/GATE
+ VDD VSS sky130_asc_nfet_01v8_lvt_9
Xsky130_asc_cap_mim_m3_1_0 VDD sky130_asc_cap_mim_m3_1_4/Cout VDD VSS VSS sky130_asc_cap_mim_m3_1
Xsky130_asc_cap_mim_m3_1_1 VDD sky130_asc_cap_mim_m3_1_4/Cout VDD VSS VSS sky130_asc_cap_mim_m3_1
Xsky130_asc_pnp_05v5_W3p40L3p40_8_0 sky130_asc_res_xhigh_po_2p85_1_19/Rout VSS VSS
+ VDD VSS sky130_asc_pnp_05v5_W3p40L3p40_8
Xsky130_asc_cap_mim_m3_1_2 VDD sky130_asc_cap_mim_m3_1_4/Cout VDD VSS VSS sky130_asc_cap_mim_m3_1
Xsky130_asc_pnp_05v5_W3p40L3p40_8_1 sky130_asc_res_xhigh_po_2p85_1_19/Rout VSS VSS
+ VDD VSS sky130_asc_pnp_05v5_W3p40L3p40_8
Xsky130_asc_cap_mim_m3_1_3 VDD sky130_asc_cap_mim_m3_1_4/Cout VDD VSS VSS sky130_asc_cap_mim_m3_1
Xsky130_asc_pnp_05v5_W3p40L3p40_8_2 sky130_asc_res_xhigh_po_2p85_1_19/Rout VSS VSS
+ VDD VSS sky130_asc_pnp_05v5_W3p40L3p40_8
Xsky130_asc_cap_mim_m3_1_4 VDD sky130_asc_cap_mim_m3_1_4/Cout VDD VSS VSS sky130_asc_cap_mim_m3_1
Xsky130_asc_pnp_05v5_W3p40L3p40_8_3 sky130_asc_res_xhigh_po_2p85_1_19/Rout VSS VSS
+ VDD VSS sky130_asc_pnp_05v5_W3p40L3p40_8
Xsky130_asc_cap_mim_m3_1_5 va VSS VDD VSS VSS sky130_asc_cap_mim_m3_1
Xsky130_asc_res_xhigh_po_2p85_1_0 sky130_asc_res_xhigh_po_2p85_1_0/Rin VSS VDD VSS
+ sky130_asc_res_xhigh_po_2p85_1_0/a_2148_115# sky130_asc_res_xhigh_po_2p85_1
Xsky130_asc_cap_mim_m3_1_6 va VSS VDD VSS VSS sky130_asc_cap_mim_m3_1
Xsky130_asc_nfet_01v8_lvt_1_0 sky130_asc_nfet_01v8_lvt_1_1/GATE VSS sky130_asc_nfet_01v8_lvt_1_1/GATE
+ VDD VSS sky130_asc_nfet_01v8_lvt_1
Xsky130_asc_res_xhigh_po_2p85_1_1 sky130_asc_res_xhigh_po_2p85_1_1/Rin sky130_asc_res_xhigh_po_2p85_1_0/Rin
+ VDD VSS sky130_asc_res_xhigh_po_2p85_1_1/a_2148_115# sky130_asc_res_xhigh_po_2p85_1
Xsky130_asc_cap_mim_m3_1_7 va VSS VDD VSS VSS sky130_asc_cap_mim_m3_1
Xsky130_asc_nfet_01v8_lvt_1_1 sky130_asc_nfet_01v8_lvt_1_1/GATE VSS sky130_asc_nfet_01v8_lvt_1_1/DRAIN
+ VDD VSS sky130_asc_nfet_01v8_lvt_1
Xsky130_asc_res_xhigh_po_2p85_1_2 sky130_asc_res_xhigh_po_2p85_1_2/Rin sky130_asc_res_xhigh_po_2p85_1_1/Rin
+ VDD VSS sky130_asc_res_xhigh_po_2p85_1_2/a_2148_115# sky130_asc_res_xhigh_po_2p85_1
Xsky130_asc_cap_mim_m3_1_8 va VSS VDD VSS VSS sky130_asc_cap_mim_m3_1
Xsky130_asc_res_xhigh_po_2p85_1_3 sky130_asc_res_xhigh_po_2p85_1_3/Rin sky130_asc_res_xhigh_po_2p85_1_2/Rin
+ VDD VSS sky130_asc_res_xhigh_po_2p85_1_3/a_2148_115# sky130_asc_res_xhigh_po_2p85_1
Xsky130_asc_cap_mim_m3_1_9 va VSS VDD VSS VSS sky130_asc_cap_mim_m3_1
Xsky130_asc_res_xhigh_po_2p85_1_4 sky130_asc_res_xhigh_po_2p85_1_4/Rin sky130_asc_res_xhigh_po_2p85_1_3/Rin
+ VDD VSS sky130_asc_res_xhigh_po_2p85_1_4/a_2148_115# sky130_asc_res_xhigh_po_2p85_1
Xsky130_asc_res_xhigh_po_2p85_1_5 sky130_asc_res_xhigh_po_2p85_1_5/Rin sky130_asc_res_xhigh_po_2p85_1_4/Rin
+ VDD VSS sky130_asc_res_xhigh_po_2p85_1_5/a_2148_115# sky130_asc_res_xhigh_po_2p85_1
Xsky130_asc_res_xhigh_po_2p85_1_6 sky130_asc_res_xhigh_po_2p85_1_6/Rin sky130_asc_res_xhigh_po_2p85_1_5/Rin
+ VDD VSS sky130_asc_res_xhigh_po_2p85_1_6/a_2148_115# sky130_asc_res_xhigh_po_2p85_1
C0 sky130_asc_res_xhigh_po_2p85_1_10/Rin sky130_asc_res_xhigh_po_2p85_1_9/a_2148_115# 0.20fF
C1 sky130_asc_res_xhigh_po_2p85_2_0/Rin sky130_asc_res_xhigh_po_2p85_1_17/Rin 0.03fF
C2 VSS sky130_asc_res_xhigh_po_2p85_2_0/a_2723_115# 0.00fF
C3 sky130_asc_res_xhigh_po_2p85_2_0/Rin sky130_asc_cap_mim_m3_1_4/Cout 0.34fF
C4 sky130_asc_res_xhigh_po_2p85_2_0/Rin vb 0.07fF
C5 sky130_asc_res_xhigh_po_2p85_2_1/Rin sky130_asc_nfet_01v8_lvt_1_1/DRAIN 0.05fF
C6 VDD sky130_asc_res_xhigh_po_2p85_1_15/Rin 0.32fF
C7 sky130_asc_res_xhigh_po_2p85_1_0/Rin sky130_asc_res_xhigh_po_2p85_1_6/Rin 1.60fF
C8 sky130_asc_res_xhigh_po_2p85_1_9/Rin sky130_asc_res_xhigh_po_2p85_1_19/Rout 0.03fF
C9 VDD sky130_asc_res_xhigh_po_2p85_1_21/Rin 0.35fF
C10 sky130_asc_nfet_01v8_lvt_1_1/GATE sky130_asc_res_xhigh_po_2p85_1_22/Rin 0.47fF
C11 vbg sky130_asc_res_xhigh_po_2p85_1_3/Rin 0.03fF
C12 VDD vbg 0.42fF
C13 sky130_asc_res_xhigh_po_2p85_1_4/a_2148_115# sky130_asc_res_xhigh_po_2p85_1_5/Rin 0.62fF
C14 sky130_asc_res_xhigh_po_2p85_2_1/a_2723_115# sky130_asc_res_xhigh_po_2p85_1_29/Rin 0.20fF
C15 porst sky130_asc_cap_mim_m3_1_4/Cout 0.39fF
C16 VSS sky130_asc_nfet_01v8_lvt_1_1/GATE 0.46fF
C17 VDD sky130_asc_pfet_01v8_lvt_6_1/GATE 0.45fF
C18 sky130_asc_res_xhigh_po_2p85_1_9/Rin sky130_asc_res_xhigh_po_2p85_1_19/a_2148_115# 0.23fF
C19 sky130_asc_res_xhigh_po_2p85_1_20/a_2148_115# sky130_asc_res_xhigh_po_2p85_1_18/Rin 0.12fF
C20 sky130_asc_res_xhigh_po_2p85_1_23/Rin vb 0.96fF
C21 sky130_asc_cap_mim_m3_1_4/Cout sky130_asc_res_xhigh_po_2p85_1_29/Rin 1.05fF
C22 VSS sky130_asc_res_xhigh_po_2p85_1_9/Rin 0.25fF
C23 vb sky130_asc_res_xhigh_po_2p85_1_29/Rin 0.04fF
C24 sky130_asc_res_xhigh_po_2p85_1_22/Rin sky130_asc_res_xhigh_po_2p85_1_21/Rin 0.45fF
C25 sky130_asc_res_xhigh_po_2p85_1_14/Rin sky130_asc_res_xhigh_po_2p85_1_13/Rin 0.45fF
C26 VDD sky130_asc_res_xhigh_po_2p85_1_0/Rin 6.93fF
C27 vb sky130_asc_res_xhigh_po_2p85_1_20/a_2148_115# 0.28fF
C28 VDD sky130_asc_res_xhigh_po_2p85_2_0/Rin 1.64fF
C29 VSS sky130_asc_res_xhigh_po_2p85_1_15/Rin 0.68fF
C30 sky130_asc_pfet_01v8_lvt_6_1/GATE sky130_asc_res_xhigh_po_2p85_1_28/Rin 0.03fF
C31 VSS sky130_asc_res_xhigh_po_2p85_1_21/Rin 1.69fF
C32 sky130_asc_res_xhigh_po_2p85_1_20/a_2148_115# sky130_asc_res_xhigh_po_2p85_1_19/Rin 0.08fF
C33 sky130_asc_nfet_01v8_lvt_1_1/GATE va 1.32fF
C34 VSS vbg 0.65fF
C35 sky130_asc_res_xhigh_po_2p85_2_0/Rin sky130_asc_res_xhigh_po_2p85_1_19/Rout 3.52fF
C36 sky130_asc_res_xhigh_po_2p85_2_0/Rin sky130_asc_res_xhigh_po_2p85_1_28/Rin 0.03fF
C37 sky130_asc_res_xhigh_po_2p85_1_12/Rin sky130_asc_res_xhigh_po_2p85_1_13/Rin 0.20fF
C38 sky130_asc_res_xhigh_po_2p85_2_0/Rin sky130_asc_res_xhigh_po_2p85_1_11/Rin 0.05fF
C39 VDD sky130_asc_res_xhigh_po_2p85_1_23/Rin 0.97fF
C40 VDD porst 0.15fF
C41 VSS sky130_asc_pfet_01v8_lvt_6_1/GATE 0.64fF
C42 sky130_asc_res_xhigh_po_2p85_1_10/Rin sky130_asc_res_xhigh_po_2p85_1_18/Rin 1.37fF
C43 VDD sky130_asc_res_xhigh_po_2p85_1_29/Rin 1.38fF
C44 sky130_asc_res_xhigh_po_2p85_1_16/a_2148_115# sky130_asc_res_xhigh_po_2p85_1_24/Rin 0.20fF
C45 sky130_asc_res_xhigh_po_2p85_1_10/Rin sky130_asc_res_xhigh_po_2p85_1_17/Rin 0.03fF
C46 sky130_asc_res_xhigh_po_2p85_1_0/a_2148_115# sky130_asc_res_xhigh_po_2p85_1_0/Rin 0.19fF
C47 sky130_asc_res_xhigh_po_2p85_1_26/Rin sky130_asc_cap_mim_m3_1_4/Cout 1.35fF
C48 sky130_asc_res_xhigh_po_2p85_1_10/Rin vb 0.07fF
C49 sky130_asc_res_xhigh_po_2p85_2_0/Rin sky130_asc_res_xhigh_po_2p85_1_19/a_2148_115# 0.50fF
C50 VSS sky130_asc_res_xhigh_po_2p85_2_0/Rin 3.27fF
C51 sky130_asc_res_xhigh_po_2p85_1_26/Rin vb 0.07fF
C52 VSS sky130_asc_res_xhigh_po_2p85_1_14/a_2148_115# 0.20fF
C53 sky130_asc_res_xhigh_po_2p85_1_29/Rin sky130_asc_res_xhigh_po_2p85_1_28/Rin 1.82fF
C54 sky130_asc_res_xhigh_po_2p85_1_23/Rin sky130_asc_res_xhigh_po_2p85_1_22/Rin 0.45fF
C55 va sky130_asc_pfet_01v8_lvt_6_1/GATE 0.08fF
C56 sky130_asc_res_xhigh_po_2p85_1_10/a_2148_115# sky130_asc_res_xhigh_po_2p85_1_18/Rin 0.05fF
C57 sky130_asc_nfet_01v8_lvt_1_1/DRAIN sky130_asc_cap_mim_m3_1_4/Cout 4.50fF
C58 vb sky130_asc_nfet_01v8_lvt_1_1/DRAIN 0.58fF
C59 sky130_asc_res_xhigh_po_2p85_1_6/a_2148_115# sky130_asc_res_xhigh_po_2p85_1_0/Rin 0.17fF
C60 sky130_asc_res_xhigh_po_2p85_1_10/a_2148_115# vb 0.20fF
C61 sky130_asc_res_xhigh_po_2p85_2_1/Rin sky130_asc_cap_mim_m3_1_4/Cout 1.95fF
C62 sky130_asc_res_xhigh_po_2p85_1_1/Rin sky130_asc_res_xhigh_po_2p85_1_0/Rin 0.48fF
C63 VSS porst 0.42fF
C64 vb sky130_asc_res_xhigh_po_2p85_2_1/Rin 0.04fF
C65 VSS sky130_asc_res_xhigh_po_2p85_1_29/Rin 0.42fF
C66 sky130_asc_res_xhigh_po_2p85_1_30/a_2148_115# sky130_asc_pfet_01v8_lvt_6_1/GATE 0.16fF
C67 VDD sky130_asc_res_xhigh_po_2p85_1_10/Rin 2.79fF
C68 sky130_asc_res_xhigh_po_2p85_1_26/a_2148_115# sky130_asc_res_xhigh_po_2p85_1_25/Rin 0.02fF
C69 VDD sky130_asc_res_xhigh_po_2p85_1_26/Rin 1.26fF
C70 sky130_asc_res_xhigh_po_2p85_1_10/a_2148_115# sky130_asc_res_xhigh_po_2p85_1_19/Rin 0.20fF
C71 VDD sky130_asc_res_xhigh_po_2p85_1_13/Rin 0.11fF
C72 sky130_asc_res_xhigh_po_2p85_1_10/Rin sky130_asc_res_xhigh_po_2p85_1_19/Rout 0.56fF
C73 sky130_asc_res_xhigh_po_2p85_1_23/Rin sky130_asc_res_xhigh_po_2p85_1_24/Rin 0.49fF
C74 va sky130_asc_res_xhigh_po_2p85_1_29/Rin 0.50fF
C75 sky130_asc_res_xhigh_po_2p85_1_10/Rin sky130_asc_res_xhigh_po_2p85_1_11/Rin 0.57fF
C76 sky130_asc_res_xhigh_po_2p85_1_26/Rin sky130_asc_res_xhigh_po_2p85_1_28/Rin 2.81fF
C77 VDD sky130_asc_nfet_01v8_lvt_1_1/DRAIN 1.08fF
C78 vb sky130_asc_res_xhigh_po_2p85_1_18/a_2148_115# 0.28fF
C79 VDD sky130_asc_res_xhigh_po_2p85_1_7/Rin 0.80fF
C80 VDD sky130_asc_res_xhigh_po_2p85_2_1/Rin 0.65fF
C81 sky130_asc_res_xhigh_po_2p85_1_23/Rin sky130_asc_res_xhigh_po_2p85_1_24/a_2148_115# 0.62fF
C82 sky130_asc_res_xhigh_po_2p85_1_11/Rin sky130_asc_res_xhigh_po_2p85_1_13/Rin 0.05fF
C83 sky130_asc_nfet_01v8_lvt_1_1/GATE sky130_asc_res_xhigh_po_2p85_1_21/Rin 0.19fF
C84 VSS sky130_asc_res_xhigh_po_2p85_1_10/Rin 0.36fF
C85 VSS sky130_asc_res_xhigh_po_2p85_1_26/Rin 0.42fF
C86 VDD sky130_asc_res_xhigh_po_2p85_1_27/Rin 1.50fF
C87 sky130_asc_nfet_01v8_lvt_1_1/DRAIN sky130_asc_res_xhigh_po_2p85_1_28/Rin 0.07fF
C88 sky130_asc_res_xhigh_po_2p85_1_25/Rin sky130_asc_cap_mim_m3_1_4/Cout 0.24fF
C89 VSS sky130_asc_res_xhigh_po_2p85_1_13/Rin 0.11fF
C90 sky130_asc_res_xhigh_po_2p85_2_1/Rin sky130_asc_res_xhigh_po_2p85_1_28/Rin 0.52fF
C91 sky130_asc_res_xhigh_po_2p85_1_1/Rin sky130_asc_res_xhigh_po_2p85_1_7/a_2148_115# 0.20fF
C92 sky130_asc_res_xhigh_po_2p85_1_12/a_2148_115# sky130_asc_res_xhigh_po_2p85_1_13/Rin 1.05fF
C93 vb sky130_asc_res_xhigh_po_2p85_1_25/Rin 0.05fF
C94 sky130_asc_res_xhigh_po_2p85_1_8/a_2148_115# sky130_asc_res_xhigh_po_2p85_1_2/Rin 0.20fF
C95 VSS sky130_asc_nfet_01v8_lvt_1_1/DRAIN 0.34fF
C96 sky130_asc_res_xhigh_po_2p85_1_27/Rin sky130_asc_res_xhigh_po_2p85_1_28/Rin 1.14fF
C97 sky130_asc_res_xhigh_po_2p85_2_0/Rin sky130_asc_res_xhigh_po_2p85_1_9/Rin 0.29fF
C98 VSS sky130_asc_res_xhigh_po_2p85_1_7/Rin 0.11fF
C99 VSS sky130_asc_res_xhigh_po_2p85_2_1/Rin 1.88fF
C100 sky130_asc_res_xhigh_po_2p85_1_11/Rin sky130_asc_res_xhigh_po_2p85_1_9/a_2148_115# 0.51fF
C101 va sky130_asc_res_xhigh_po_2p85_1_26/Rin 0.04fF
C102 VDD sky130_asc_res_xhigh_po_2p85_1_14/Rin 0.89fF
C103 vb sky130_asc_res_xhigh_po_2p85_1_18/Rin 1.33fF
C104 sky130_asc_res_xhigh_po_2p85_1_17/Rin vb 0.25fF
C105 vb sky130_asc_cap_mim_m3_1_4/Cout 1.62fF
C106 VDD sky130_asc_res_xhigh_po_2p85_1_25/Rin 1.64fF
C107 va sky130_asc_nfet_01v8_lvt_1_1/DRAIN 0.35fF
C108 sky130_asc_res_xhigh_po_2p85_1_7/Rin sky130_asc_res_xhigh_po_2p85_1_6/a_2148_115# 0.20fF
C109 sky130_asc_res_xhigh_po_2p85_1_15/a_2148_115# sky130_asc_res_xhigh_po_2p85_1_13/Rin 0.20fF
C110 va sky130_asc_res_xhigh_po_2p85_2_1/Rin 0.07fF
C111 vbg sky130_asc_res_xhigh_po_2p85_1_5/a_2148_115# 0.20fF
C112 VSS sky130_asc_res_xhigh_po_2p85_1_18/a_2148_115# 0.16fF
C113 VDD sky130_asc_res_xhigh_po_2p85_1_12/Rin 0.90fF
C114 sky130_asc_res_xhigh_po_2p85_1_16/a_2148_115# sky130_asc_res_xhigh_po_2p85_1_23/Rin 0.20fF
C115 sky130_asc_res_xhigh_po_2p85_1_22/Rin sky130_asc_res_xhigh_po_2p85_1_25/Rin 0.45fF
C116 sky130_asc_res_xhigh_po_2p85_1_13/a_2148_115# sky130_asc_res_xhigh_po_2p85_1_19/Rin 0.21fF
C117 sky130_asc_res_xhigh_po_2p85_1_14/a_2148_115# sky130_asc_res_xhigh_po_2p85_1_0/Rin 0.20fF
C118 VDD sky130_asc_res_xhigh_po_2p85_1_18/Rin 5.98fF
C119 VDD sky130_asc_res_xhigh_po_2p85_1_17/Rin 0.11fF
C120 VDD sky130_asc_cap_mim_m3_1_4/Cout 3.35fF
C121 sky130_asc_res_xhigh_po_2p85_1_12/Rin sky130_asc_res_xhigh_po_2p85_1_11/Rin 0.05fF
C122 VDD vb 8.37fF
C123 VSS sky130_asc_res_xhigh_po_2p85_1_25/Rin 4.85fF
C124 VDD sky130_asc_res_xhigh_po_2p85_1_6/Rin 0.65fF
C125 vb sky130_asc_res_xhigh_po_2p85_1_21/a_2148_115# 1.19fF
C126 sky130_asc_res_xhigh_po_2p85_1_28/a_2148_115# sky130_asc_res_xhigh_po_2p85_1_26/Rin 0.20fF
C127 sky130_asc_res_xhigh_po_2p85_1_17/Rin sky130_asc_res_xhigh_po_2p85_1_19/Rout 0.03fF
C128 sky130_asc_res_xhigh_po_2p85_1_8/a_2148_115# sky130_asc_res_xhigh_po_2p85_1_1/Rin 0.32fF
C129 VDD sky130_asc_res_xhigh_po_2p85_1_19/Rin 2.60fF
C130 sky130_asc_cap_mim_m3_1_4/Cout sky130_asc_res_xhigh_po_2p85_1_28/Rin 1.06fF
C131 sky130_asc_res_xhigh_po_2p85_1_12/Rin sky130_asc_res_xhigh_po_2p85_1_12/a_2148_115# 0.46fF
C132 sky130_asc_res_xhigh_po_2p85_1_29/a_2148_115# sky130_asc_res_xhigh_po_2p85_1_21/Rin 0.20fF
C133 vb sky130_asc_res_xhigh_po_2p85_1_19/Rout 0.55fF
C134 sky130_asc_res_xhigh_po_2p85_1_2/Rin sky130_asc_res_xhigh_po_2p85_1_3/Rin 2.33fF
C135 vb sky130_asc_res_xhigh_po_2p85_1_28/Rin 0.07fF
C136 VDD sky130_asc_res_xhigh_po_2p85_1_2/Rin 0.11fF
C137 sky130_asc_res_xhigh_po_2p85_1_27/Rin sky130_asc_res_xhigh_po_2p85_2_0/a_2723_115# 0.20fF
C138 sky130_asc_res_xhigh_po_2p85_1_24/Rin sky130_asc_res_xhigh_po_2p85_1_25/Rin 0.08fF
C139 VSS sky130_asc_res_xhigh_po_2p85_2_1/a_2723_115# 0.00fF
C140 VSS sky130_asc_res_xhigh_po_2p85_1_18/Rin 0.11fF
C141 sky130_asc_res_xhigh_po_2p85_1_13/a_2148_115# sky130_asc_res_xhigh_po_2p85_1_11/Rin -0.01fF
C142 VSS sky130_asc_res_xhigh_po_2p85_1_17/Rin 0.11fF
C143 sky130_asc_res_xhigh_po_2p85_1_14/Rin sky130_asc_res_xhigh_po_2p85_1_15/a_2148_115# 0.69fF
C144 VDD sky130_asc_res_xhigh_po_2p85_1_3/Rin 0.11fF
C145 sky130_asc_nfet_01v8_lvt_1_1/GATE sky130_asc_nfet_01v8_lvt_1_1/DRAIN 0.19fF
C146 VSS sky130_asc_cap_mim_m3_1_4/Cout 3.66fF
C147 sky130_asc_nfet_01v8_lvt_1_1/GATE sky130_asc_res_xhigh_po_2p85_2_1/Rin 0.04fF
C148 VSS vb 4.68fF
C149 sky130_asc_res_xhigh_po_2p85_1_0/Rin sky130_asc_res_xhigh_po_2p85_1_7/a_2148_115# 0.38fF
C150 sky130_asc_res_xhigh_po_2p85_1_0/a_2148_115# sky130_asc_res_xhigh_po_2p85_1_6/Rin 0.20fF
C151 sky130_asc_res_xhigh_po_2p85_1_28/a_2148_115# sky130_asc_res_xhigh_po_2p85_1_27/Rin 0.49fF
C152 sky130_asc_res_xhigh_po_2p85_1_26/Rin sky130_asc_pfet_01v8_lvt_6_1/GATE 0.03fF
C153 VDD sky130_asc_res_xhigh_po_2p85_1_19/Rout 0.53fF
C154 VSS sky130_asc_res_xhigh_po_2p85_1_19/Rin 1.24fF
C155 va sky130_asc_res_xhigh_po_2p85_2_1/a_2723_115# 0.19fF
C156 VDD sky130_asc_res_xhigh_po_2p85_1_28/Rin 0.58fF
C157 sky130_asc_res_xhigh_po_2p85_2_1/Rin sky130_asc_res_xhigh_po_2p85_1_21/Rin 0.45fF
C158 VSS sky130_asc_res_xhigh_po_2p85_1_2/Rin 0.12fF
C159 sky130_asc_res_xhigh_po_2p85_1_1/a_2148_115# sky130_asc_res_xhigh_po_2p85_1_2/Rin 0.20fF
C160 sky130_asc_res_xhigh_po_2p85_2_0/Rin sky130_asc_res_xhigh_po_2p85_1_10/Rin 0.03fF
C161 VDD sky130_asc_res_xhigh_po_2p85_1_22/Rin 0.21fF
C162 va sky130_asc_cap_mim_m3_1_4/Cout 2.03fF
C163 sky130_asc_res_xhigh_po_2p85_2_0/Rin sky130_asc_res_xhigh_po_2p85_1_26/Rin 0.03fF
C164 va vb 0.04fF
C165 sky130_asc_res_xhigh_po_2p85_1_24/Rin vb 0.03fF
C166 sky130_asc_res_xhigh_po_2p85_1_6/a_2148_115# sky130_asc_res_xhigh_po_2p85_1_6/Rin 0.72fF
C167 VSS sky130_asc_res_xhigh_po_2p85_1_3/Rin 2.54fF
C168 sky130_asc_res_xhigh_po_2p85_1_1/a_2148_115# sky130_asc_res_xhigh_po_2p85_1_3/Rin 0.20fF
C169 sky130_asc_pfet_01v8_lvt_6_1/GATE sky130_asc_nfet_01v8_lvt_1_1/DRAIN 1.64fF
C170 VSS sky130_asc_res_xhigh_po_2p85_1_22/a_2148_115# 0.02fF
C171 VDD VSS 22.87fF
C172 sky130_asc_res_xhigh_po_2p85_1_11/Rin sky130_asc_res_xhigh_po_2p85_1_19/Rout 0.05fF
C173 sky130_asc_res_xhigh_po_2p85_1_7/Rin sky130_asc_res_xhigh_po_2p85_1_0/Rin 2.58fF
C174 VSS sky130_asc_res_xhigh_po_2p85_1_19/Rout 4.18fF
C175 sky130_asc_res_xhigh_po_2p85_1_26/Rin sky130_asc_res_xhigh_po_2p85_1_29/Rin 0.03fF
C176 VSS sky130_asc_res_xhigh_po_2p85_1_28/Rin 0.42fF
C177 sky130_asc_res_xhigh_po_2p85_1_5/Rin sky130_asc_res_xhigh_po_2p85_1_4/Rin 0.17fF
C178 sky130_asc_res_xhigh_po_2p85_1_7/Rin sky130_asc_res_xhigh_po_2p85_1_5/a_2148_115# 0.22fF
C179 sky130_asc_res_xhigh_po_2p85_1_19/a_2148_115# sky130_asc_res_xhigh_po_2p85_1_11/Rin 0.29fF
C180 VSS sky130_asc_res_xhigh_po_2p85_1_11/Rin -0.64fF
C181 VSS sky130_asc_res_xhigh_po_2p85_1_22/Rin 0.21fF
C182 sky130_asc_res_xhigh_po_2p85_1_12/a_2148_115# sky130_asc_res_xhigh_po_2p85_1_11/Rin -0.08fF
C183 sky130_asc_res_xhigh_po_2p85_1_14/Rin sky130_asc_res_xhigh_po_2p85_1_15/Rin 0.03fF
C184 sky130_asc_res_xhigh_po_2p85_1_1/Rin sky130_asc_res_xhigh_po_2p85_1_3/Rin 0.87fF
C185 VDD va 3.39fF
C186 VDD sky130_asc_res_xhigh_po_2p85_1_5/Rin 1.12fF
C187 VDD sky130_asc_res_xhigh_po_2p85_1_24/Rin 0.31fF
C188 VDD sky130_asc_res_xhigh_po_2p85_1_1/Rin 0.11fF
C189 sky130_asc_nfet_01v8_lvt_1_1/DRAIN sky130_asc_res_xhigh_po_2p85_1_29/Rin 0.04fF
C190 sky130_asc_res_xhigh_po_2p85_2_1/Rin sky130_asc_res_xhigh_po_2p85_1_29/Rin 0.03fF
C191 va sky130_asc_res_xhigh_po_2p85_1_28/Rin 1.13fF
C192 sky130_asc_res_xhigh_po_2p85_1_24/Rin sky130_asc_res_xhigh_po_2p85_1_22/Rin 0.45fF
C193 sky130_asc_res_xhigh_po_2p85_1_9/Rin sky130_asc_res_xhigh_po_2p85_1_17/Rin 0.73fF
C194 sky130_asc_nfet_01v8_lvt_1_1/GATE sky130_asc_cap_mim_m3_1_4/Cout 2.12fF
C195 sky130_asc_res_xhigh_po_2p85_1_4/a_2148_115# sky130_asc_res_xhigh_po_2p85_1_4/Rin 0.61fF
C196 sky130_asc_nfet_01v8_lvt_1_1/GATE vb 0.08fF
C197 sky130_asc_res_xhigh_po_2p85_1_4/a_2148_115# sky130_asc_res_xhigh_po_2p85_1_3/Rin 0.04fF
C198 sky130_asc_res_xhigh_po_2p85_1_24/a_2148_115# sky130_asc_res_xhigh_po_2p85_1_22/Rin 0.23fF
C199 VSS va 2.30fF
C200 VSS sky130_asc_res_xhigh_po_2p85_1_5/Rin -0.06fF
C201 VSS sky130_asc_res_xhigh_po_2p85_1_24/Rin 0.63fF
C202 sky130_asc_res_xhigh_po_2p85_1_0/a_2148_115# sky130_asc_res_xhigh_po_2p85_1_5/Rin 0.20fF
C203 VSS sky130_asc_res_xhigh_po_2p85_1_1/Rin 1.78fF
C204 sky130_asc_res_xhigh_po_2p85_1_7/Rin sky130_asc_res_xhigh_po_2p85_1_7/a_2148_115# 0.50fF
C205 sky130_asc_res_xhigh_po_2p85_1_15/Rin sky130_asc_res_xhigh_po_2p85_1_18/Rin 0.45fF
C206 sky130_asc_res_xhigh_po_2p85_1_29/a_2148_115# sky130_asc_res_xhigh_po_2p85_2_1/Rin 0.20fF
C207 sky130_asc_res_xhigh_po_2p85_1_21/Rin sky130_asc_cap_mim_m3_1_4/Cout 2.48fF
C208 sky130_asc_res_xhigh_po_2p85_1_9/Rin sky130_asc_res_xhigh_po_2p85_1_19/Rin 0.03fF
C209 vb sky130_asc_res_xhigh_po_2p85_1_21/Rin 0.04fF
C210 VSS sky130_asc_res_xhigh_po_2p85_1_30/a_2148_115# 0.01fF
C211 vbg sky130_asc_cap_mim_m3_1_4/Cout 0.37fF
C212 sky130_asc_res_xhigh_po_2p85_1_26/Rin sky130_asc_nfet_01v8_lvt_1_1/DRAIN 0.03fF
C213 sky130_asc_res_xhigh_po_2p85_2_0/a_2723_115# sky130_asc_res_xhigh_po_2p85_1_28/Rin 0.19fF
C214 sky130_asc_res_xhigh_po_2p85_1_11/a_2148_115# sky130_asc_res_xhigh_po_2p85_1_17/Rin 0.20fF
C215 sky130_asc_res_xhigh_po_2p85_1_26/Rin sky130_asc_res_xhigh_po_2p85_2_1/Rin 0.03fF
C216 sky130_asc_res_xhigh_po_2p85_1_11/a_2148_115# vb 0.22fF
C217 sky130_asc_pfet_01v8_lvt_6_1/GATE sky130_asc_cap_mim_m3_1_4/Cout 0.95fF
C218 sky130_asc_nfet_01v8_lvt_1_1/GATE sky130_asc_res_xhigh_po_2p85_1_22/a_2148_115# -0.26fF
C219 VDD sky130_asc_nfet_01v8_lvt_1_1/GATE -0.36fF
C220 VDD sky130_asc_res_xhigh_po_2p85_1_9/Rin 0.18fF
C221 vb sky130_asc_pfet_01v8_lvt_6_1/GATE -0.08fF
C222 VSS 0 708.39fF
C223 VDD 0 1018.97fF
C224 vbg 0 13.66fF
C225 sky130_asc_res_xhigh_po_2p85_1_11/Rin 0 5.90fF
C226 sky130_asc_res_xhigh_po_2p85_1_25/Rin 0 3.74fF
C227 sky130_asc_res_xhigh_po_2p85_1_2/Rin 0 2.78fF
C228 sky130_asc_res_xhigh_po_2p85_1_1/Rin 0 3.72fF
C229 sky130_asc_res_xhigh_po_2p85_1_3/Rin 0 4.18fF
C230 sky130_asc_res_xhigh_po_2p85_1_0/Rin 0 7.34fF
C231 sky130_asc_res_xhigh_po_2p85_1_5/Rin 0 3.90fF
C232 sky130_asc_res_xhigh_po_2p85_1_27/Rin 0 3.36fF
C233 sky130_asc_res_xhigh_po_2p85_1_17/Rin 0 4.04fF
C234 sky130_asc_res_xhigh_po_2p85_1_12/Rin 0 3.62fF
C235 sky130_asc_res_xhigh_po_2p85_1_13/Rin 0 2.58fF
C236 sky130_asc_res_xhigh_po_2p85_1_22/Rin 0 2.49fF
C237 sky130_asc_res_xhigh_po_2p85_1_18/Rin 0 4.72fF
C238 sky130_asc_res_xhigh_po_2p85_1_15/Rin 0 3.65fF
C239 sky130_asc_res_xhigh_po_2p85_1_28/Rin 0 5.08fF
C240 sky130_asc_res_xhigh_po_2p85_1_29/Rin 0 4.80fF
C241 sky130_asc_res_xhigh_po_2p85_2_1/Rin 0 7.65fF
C242 sky130_asc_res_xhigh_po_2p85_1_26/Rin 0 5.38fF
C243 porst 0 12.68fF
C244 sky130_asc_nfet_01v8_lvt_1_1/GATE 0 9.98fF
C245 sky130_asc_nfet_01v8_lvt_1_1/DRAIN 0 8.50fF
C246 sky130_asc_res_xhigh_po_2p85_1_6/a_2148_115# 0 2.70fF
C247 sky130_asc_res_xhigh_po_2p85_1_4/Rin 0 3.30fF
C248 sky130_asc_res_xhigh_po_2p85_1_5/a_2148_115# 0 2.70fF
C249 sky130_asc_res_xhigh_po_2p85_1_4/a_2148_115# 0 2.70fF
C250 va 0 68.89fF
C251 sky130_asc_res_xhigh_po_2p85_1_3/a_2148_115# 0 2.70fF
C252 sky130_asc_res_xhigh_po_2p85_1_2/a_2148_115# 0 2.70fF
C253 sky130_asc_res_xhigh_po_2p85_1_1/a_2148_115# 0 2.70fF
C254 sky130_asc_res_xhigh_po_2p85_1_0/a_2148_115# 0 2.70fF
C255 sky130_asc_pfet_01v8_lvt_6_1/GATE 0 11.12fF
C256 sky130_asc_res_xhigh_po_2p85_1_19/Rout 0 54.88fF
C257 sky130_asc_res_xhigh_po_2p85_1_19/Rin 0 4.26fF
C258 sky130_asc_res_xhigh_po_2p85_1_19/a_2148_115# 0 2.70fF
C259 sky130_asc_res_xhigh_po_2p85_1_29/a_2148_115# 0 2.70fF
C260 sky130_asc_res_xhigh_po_2p85_1_18/a_2148_115# 0 2.70fF
C261 sky130_asc_res_xhigh_po_2p85_1_28/a_2148_115# 0 2.70fF
C262 sky130_asc_res_xhigh_po_2p85_1_17/a_2148_115# 0 2.70fF
C263 sky130_asc_res_xhigh_po_2p85_1_27/a_2148_115# 0 2.70fF
C264 sky130_asc_res_xhigh_po_2p85_1_16/a_2148_115# 0 2.70fF
C265 sky130_asc_res_xhigh_po_2p85_1_26/a_2148_115# 0 2.70fF
C266 sky130_asc_res_xhigh_po_2p85_1_14/Rin 0 3.87fF
C267 sky130_asc_res_xhigh_po_2p85_1_15/a_2148_115# 0 2.70fF
C268 sky130_asc_res_xhigh_po_2p85_1_25/a_2148_115# 0 2.70fF
C269 sky130_asc_res_xhigh_po_2p85_1_14/a_2148_115# 0 2.70fF
C270 sky130_asc_res_xhigh_po_2p85_1_23/Rin 0 3.26fF
C271 sky130_asc_res_xhigh_po_2p85_1_24/Rin 0 3.37fF
C272 sky130_asc_res_xhigh_po_2p85_1_24/a_2148_115# 0 2.70fF
C273 sky130_asc_res_xhigh_po_2p85_1_13/a_2148_115# 0 2.70fF
C274 sky130_asc_res_xhigh_po_2p85_1_23/a_2148_115# 0 2.70fF
C275 sky130_asc_res_xhigh_po_2p85_1_12/a_2148_115# 0 2.70fF
C276 sky130_asc_res_xhigh_po_2p85_2_1/a_2723_115# 0 2.70fF
C277 sky130_asc_res_xhigh_po_2p85_1_22/a_2148_115# 0 2.70fF
C278 sky130_asc_res_xhigh_po_2p85_1_11/a_2148_115# 0 2.70fF
C279 sky130_asc_res_xhigh_po_2p85_2_0/a_2723_115# 0 2.70fF
C280 sky130_asc_res_xhigh_po_2p85_1_21/Rin 0 2.99fF
C281 sky130_asc_res_xhigh_po_2p85_1_21/a_2148_115# 0 2.70fF
C282 sky130_asc_res_xhigh_po_2p85_1_10/Rin 0 5.89fF
C283 sky130_asc_res_xhigh_po_2p85_1_10/a_2148_115# 0 2.70fF
C284 vb 0 29.85fF
C285 sky130_asc_res_xhigh_po_2p85_1_20/a_2148_115# 0 2.70fF
C286 sky130_asc_res_xhigh_po_2p85_1_30/a_2148_115# 0 2.70fF
C287 sky130_asc_cap_mim_m3_1_4/Cout 0 128.21fF
C288 sky130_asc_res_xhigh_po_2p85_2_0/Rin 0 5.29fF
C289 sky130_asc_res_xhigh_po_2p85_1_9/Rin 0 8.73fF
C290 sky130_asc_res_xhigh_po_2p85_1_9/a_2148_115# 0 2.70fF
C291 sky130_asc_res_xhigh_po_2p85_1_7/Rin 0 4.15fF
C292 sky130_asc_res_xhigh_po_2p85_1_8/a_2148_115# 0 2.70fF
C293 sky130_asc_res_xhigh_po_2p85_1_6/Rin 0 3.60fF
C294 sky130_asc_res_xhigh_po_2p85_1_7/a_2148_115# 0 2.70fF
.ends

