magic
tech sky130A
magscale 1 2
timestamp 1652146737
<< locali >>
rect 2 1850 172 1910
rect 232 1850 572 1910
rect 632 1850 972 1910
rect 1032 1850 1372 1910
rect 1432 1850 1772 1910
rect 1832 1850 2172 1910
rect 2232 1850 2572 1910
rect 2632 1850 2972 1910
rect 3032 1850 3372 1910
rect 3432 1850 3772 1910
rect 3832 1850 4172 1910
rect 4232 1850 4572 1910
rect 4632 1850 4972 1910
rect 5032 1850 5372 1910
rect 5432 1850 5772 1910
rect 5832 1850 6172 1910
rect 6232 1850 6572 1910
rect 6632 1850 6972 1910
rect 7032 1850 7170 1910
rect 2 -30 172 30
rect 232 -30 572 30
rect 632 -30 972 30
rect 1032 -30 1372 30
rect 1432 -30 1772 30
rect 1832 -30 2172 30
rect 2232 -30 2572 30
rect 2632 -30 2972 30
rect 3032 -30 3372 30
rect 3432 -30 3772 30
rect 3832 -30 4172 30
rect 4232 -30 4572 30
rect 4632 -30 4972 30
rect 5032 -30 5372 30
rect 5432 -30 5772 30
rect 5832 -30 6172 30
rect 6232 -30 6572 30
rect 6632 -30 6972 30
rect 7032 -30 7170 30
<< viali >>
rect 172 1850 232 1910
rect 572 1850 632 1910
rect 972 1850 1032 1910
rect 1372 1850 1432 1910
rect 1772 1850 1832 1910
rect 2172 1850 2232 1910
rect 2572 1850 2632 1910
rect 2972 1850 3032 1910
rect 3372 1850 3432 1910
rect 3772 1850 3832 1910
rect 4172 1850 4232 1910
rect 4572 1850 4632 1910
rect 4972 1850 5032 1910
rect 5372 1850 5432 1910
rect 5772 1850 5832 1910
rect 6172 1850 6232 1910
rect 6572 1850 6632 1910
rect 6972 1850 7032 1910
rect 172 -30 232 30
rect 572 -30 632 30
rect 972 -30 1032 30
rect 1372 -30 1432 30
rect 1772 -30 1832 30
rect 2172 -30 2232 30
rect 2572 -30 2632 30
rect 2972 -30 3032 30
rect 3372 -30 3432 30
rect 3772 -30 3832 30
rect 4172 -30 4232 30
rect 4572 -30 4632 30
rect 4972 -30 5032 30
rect 5372 -30 5432 30
rect 5772 -30 5832 30
rect 6172 -30 6232 30
rect 6572 -30 6632 30
rect 6972 -30 7032 30
<< metal1 >>
rect 2 1910 7170 1940
rect 2 1850 172 1910
rect 232 1850 572 1910
rect 632 1850 972 1910
rect 1032 1850 1372 1910
rect 1432 1850 1772 1910
rect 1832 1850 2172 1910
rect 2232 1850 2572 1910
rect 2632 1850 2972 1910
rect 3032 1850 3372 1910
rect 3432 1850 3772 1910
rect 3832 1850 4172 1910
rect 4232 1850 4572 1910
rect 4632 1850 4972 1910
rect 5032 1850 5372 1910
rect 5432 1850 5772 1910
rect 5832 1850 6172 1910
rect 6232 1850 6572 1910
rect 6632 1850 6972 1910
rect 7032 1850 7170 1910
rect 2 1820 7170 1850
rect 2 30 7170 60
rect 2 -30 172 30
rect 232 -30 572 30
rect 632 -30 972 30
rect 1032 -30 1372 30
rect 1432 -30 1772 30
rect 1832 -30 2172 30
rect 2232 -30 2572 30
rect 2632 -30 2972 30
rect 3032 -30 3372 30
rect 3432 -30 3772 30
rect 3832 -30 4172 30
rect 4232 -30 4572 30
rect 4632 -30 4972 30
rect 5032 -30 5372 30
rect 5432 -30 5772 30
rect 5832 -30 6172 30
rect 6232 -30 6572 30
rect 6632 -30 6972 30
rect 7032 -30 7170 30
rect 2 -60 7170 -30
<< metal3 >>
rect 0 1650 7170 1690
rect 0 1622 7171 1650
rect 0 1078 616 1622
rect 680 1078 1335 1622
rect 1399 1078 2054 1622
rect 2118 1078 2773 1622
rect 2837 1078 3492 1622
rect 3556 1078 4211 1622
rect 4275 1078 4930 1622
rect 4994 1078 5649 1622
rect 5713 1078 6368 1622
rect 6432 1078 7087 1622
rect 7151 1078 7171 1622
rect 0 1050 7171 1078
rect 0 950 7170 1050
rect 0 922 7171 950
rect 0 378 616 922
rect 680 378 1335 922
rect 1399 378 2054 922
rect 2118 378 2773 922
rect 2837 378 3492 922
rect 3556 378 4211 922
rect 4275 378 4930 922
rect 4994 378 5649 922
rect 5713 378 6368 922
rect 6432 378 7087 922
rect 7151 378 7171 922
rect 0 350 7171 378
<< via3 >>
rect 616 1078 680 1622
rect 1335 1078 1399 1622
rect 2054 1078 2118 1622
rect 2773 1078 2837 1622
rect 3492 1078 3556 1622
rect 4211 1078 4275 1622
rect 4930 1078 4994 1622
rect 5649 1078 5713 1622
rect 6368 1078 6432 1622
rect 7087 1078 7151 1622
rect 616 378 680 922
rect 1335 378 1399 922
rect 2054 378 2118 922
rect 2773 378 2837 922
rect 3492 378 3556 922
rect 4211 378 4275 922
rect 4930 378 4994 922
rect 5649 378 5713 922
rect 6368 378 6432 922
rect 7087 378 7151 922
<< mimcap >>
rect 101 1510 501 1550
rect 101 1190 141 1510
rect 461 1190 501 1510
rect 101 1150 501 1190
rect 820 1510 1220 1550
rect 820 1190 860 1510
rect 1180 1190 1220 1510
rect 820 1150 1220 1190
rect 1539 1510 1939 1550
rect 1539 1190 1579 1510
rect 1899 1190 1939 1510
rect 1539 1150 1939 1190
rect 2258 1510 2658 1550
rect 2258 1190 2298 1510
rect 2618 1190 2658 1510
rect 2258 1150 2658 1190
rect 2977 1510 3377 1550
rect 2977 1190 3017 1510
rect 3337 1190 3377 1510
rect 2977 1150 3377 1190
rect 3696 1510 4096 1550
rect 3696 1190 3736 1510
rect 4056 1190 4096 1510
rect 3696 1150 4096 1190
rect 4415 1510 4815 1550
rect 4415 1190 4455 1510
rect 4775 1190 4815 1510
rect 4415 1150 4815 1190
rect 5134 1510 5534 1550
rect 5134 1190 5174 1510
rect 5494 1190 5534 1510
rect 5134 1150 5534 1190
rect 5853 1510 6253 1550
rect 5853 1190 5893 1510
rect 6213 1190 6253 1510
rect 5853 1150 6253 1190
rect 6572 1510 6972 1550
rect 6572 1190 6612 1510
rect 6932 1190 6972 1510
rect 6572 1150 6972 1190
rect 101 810 501 850
rect 101 490 141 810
rect 461 490 501 810
rect 101 450 501 490
rect 820 810 1220 850
rect 820 490 860 810
rect 1180 490 1220 810
rect 820 450 1220 490
rect 1539 810 1939 850
rect 1539 490 1579 810
rect 1899 490 1939 810
rect 1539 450 1939 490
rect 2258 810 2658 850
rect 2258 490 2298 810
rect 2618 490 2658 810
rect 2258 450 2658 490
rect 2977 810 3377 850
rect 2977 490 3017 810
rect 3337 490 3377 810
rect 2977 450 3377 490
rect 3696 810 4096 850
rect 3696 490 3736 810
rect 4056 490 4096 810
rect 3696 450 4096 490
rect 4415 810 4815 850
rect 4415 490 4455 810
rect 4775 490 4815 810
rect 4415 450 4815 490
rect 5134 810 5534 850
rect 5134 490 5174 810
rect 5494 490 5534 810
rect 5134 450 5534 490
rect 5853 810 6253 850
rect 5853 490 5893 810
rect 6213 490 6253 810
rect 5853 450 6253 490
rect 6572 810 6972 850
rect 6572 490 6612 810
rect 6932 490 6972 810
rect 6572 450 6972 490
<< mimcapcontact >>
rect 141 1190 461 1510
rect 860 1190 1180 1510
rect 1579 1190 1899 1510
rect 2298 1190 2618 1510
rect 3017 1190 3337 1510
rect 3736 1190 4056 1510
rect 4455 1190 4775 1510
rect 5174 1190 5494 1510
rect 5893 1190 6213 1510
rect 6612 1190 6932 1510
rect 141 490 461 810
rect 860 490 1180 810
rect 1579 490 1899 810
rect 2298 490 2618 810
rect 3017 490 3337 810
rect 3736 490 4056 810
rect 4455 490 4775 810
rect 5174 490 5494 810
rect 5893 490 6213 810
rect 6612 490 6932 810
<< metal4 >>
rect 600 1622 696 1638
rect 140 1511 460 1530
rect 140 1510 462 1511
rect 140 1190 141 1510
rect 461 1190 462 1510
rect 140 1189 462 1190
rect 140 811 460 1189
rect 600 1078 616 1622
rect 680 1078 696 1622
rect 1319 1622 1415 1638
rect 860 1511 1180 1530
rect 859 1510 1181 1511
rect 859 1190 860 1510
rect 1180 1190 1181 1510
rect 859 1189 1181 1190
rect 600 1062 696 1078
rect 600 922 696 938
rect 140 810 462 811
rect 140 490 141 810
rect 461 490 462 810
rect 140 489 462 490
rect 140 290 460 489
rect 600 378 616 922
rect 680 378 696 922
rect 860 811 1180 1189
rect 1319 1078 1335 1622
rect 1399 1078 1415 1622
rect 2038 1622 2134 1638
rect 1580 1511 1900 1530
rect 1578 1510 1900 1511
rect 1578 1190 1579 1510
rect 1899 1190 1900 1510
rect 1578 1189 1900 1190
rect 1319 1062 1415 1078
rect 1319 922 1415 938
rect 859 810 1181 811
rect 859 490 860 810
rect 1180 490 1181 810
rect 859 489 1181 490
rect 600 362 696 378
rect 860 290 1180 489
rect 1319 378 1335 922
rect 1399 378 1415 922
rect 1580 811 1900 1189
rect 2038 1078 2054 1622
rect 2118 1078 2134 1622
rect 2757 1622 2853 1638
rect 2300 1511 2620 1530
rect 2297 1510 2620 1511
rect 2297 1190 2298 1510
rect 2618 1190 2620 1510
rect 2297 1189 2620 1190
rect 2038 1062 2134 1078
rect 1578 810 1900 811
rect 1578 490 1579 810
rect 1899 490 1900 810
rect 1578 489 1900 490
rect 1319 362 1415 378
rect 1580 290 1900 489
rect 2038 922 2134 938
rect 2038 378 2054 922
rect 2118 378 2134 922
rect 2300 811 2620 1189
rect 2757 1078 2773 1622
rect 2837 1078 2853 1622
rect 3476 1622 3572 1638
rect 3020 1511 3340 1530
rect 3016 1510 3340 1511
rect 3016 1190 3017 1510
rect 3337 1190 3340 1510
rect 3016 1189 3340 1190
rect 2757 1062 2853 1078
rect 2297 810 2620 811
rect 2297 490 2298 810
rect 2618 490 2620 810
rect 2297 489 2620 490
rect 2038 362 2134 378
rect 2300 290 2620 489
rect 2757 922 2853 938
rect 2757 378 2773 922
rect 2837 378 2853 922
rect 3020 811 3340 1189
rect 3476 1078 3492 1622
rect 3556 1078 3572 1622
rect 4195 1622 4291 1638
rect 3740 1511 4060 1530
rect 3735 1510 4060 1511
rect 3735 1190 3736 1510
rect 4056 1190 4060 1510
rect 3735 1189 4060 1190
rect 3476 1062 3572 1078
rect 3016 810 3340 811
rect 3016 490 3017 810
rect 3337 490 3340 810
rect 3016 489 3340 490
rect 2757 362 2853 378
rect 3020 290 3340 489
rect 3476 922 3572 938
rect 3476 378 3492 922
rect 3556 378 3572 922
rect 3740 811 4060 1189
rect 4195 1078 4211 1622
rect 4275 1078 4291 1622
rect 4914 1622 5010 1638
rect 4460 1511 4780 1530
rect 4454 1510 4780 1511
rect 4454 1190 4455 1510
rect 4775 1190 4780 1510
rect 4454 1189 4780 1190
rect 4195 1062 4291 1078
rect 3735 810 4060 811
rect 3735 490 3736 810
rect 4056 490 4060 810
rect 3735 489 4060 490
rect 3476 362 3572 378
rect 3740 290 4060 489
rect 4195 922 4291 938
rect 4195 378 4211 922
rect 4275 378 4291 922
rect 4460 811 4780 1189
rect 4914 1078 4930 1622
rect 4994 1078 5010 1622
rect 5633 1622 5729 1638
rect 5180 1511 5500 1530
rect 5173 1510 5500 1511
rect 5173 1190 5174 1510
rect 5494 1190 5500 1510
rect 5173 1189 5500 1190
rect 4914 1062 5010 1078
rect 4454 810 4780 811
rect 4454 490 4455 810
rect 4775 490 4780 810
rect 4454 489 4780 490
rect 4195 362 4291 378
rect 4460 290 4780 489
rect 4914 922 5010 938
rect 4914 378 4930 922
rect 4994 378 5010 922
rect 5180 811 5500 1189
rect 5633 1078 5649 1622
rect 5713 1078 5729 1622
rect 6352 1622 6448 1638
rect 5900 1511 6220 1530
rect 5892 1510 6220 1511
rect 5892 1190 5893 1510
rect 6213 1190 6220 1510
rect 5892 1189 6220 1190
rect 5633 1062 5729 1078
rect 5173 810 5500 811
rect 5173 490 5174 810
rect 5494 490 5500 810
rect 5173 489 5500 490
rect 4914 362 5010 378
rect 5180 290 5500 489
rect 5633 922 5729 938
rect 5633 378 5649 922
rect 5713 378 5729 922
rect 5900 811 6220 1189
rect 6352 1078 6368 1622
rect 6432 1078 6448 1622
rect 7071 1622 7167 1638
rect 6620 1511 6940 1530
rect 6611 1510 6940 1511
rect 6611 1190 6612 1510
rect 6932 1190 6940 1510
rect 6611 1189 6940 1190
rect 6352 1062 6448 1078
rect 5892 810 6220 811
rect 5892 490 5893 810
rect 6213 490 6220 810
rect 5892 489 6220 490
rect 5633 362 5729 378
rect 5900 290 6220 489
rect 6352 922 6448 938
rect 6352 378 6368 922
rect 6432 378 6448 922
rect 6620 811 6940 1189
rect 7071 1078 7087 1622
rect 7151 1078 7167 1622
rect 7071 1062 7167 1078
rect 6611 810 6940 811
rect 6611 490 6612 810
rect 6932 490 6940 810
rect 6611 489 6940 490
rect 6352 362 6448 378
rect 6620 290 6940 489
rect 7071 922 7167 938
rect 7071 378 7087 922
rect 7151 378 7167 922
rect 7071 362 7167 378
rect 2 190 7170 290
<< labels >>
flabel metal3 0 1630 60 1690 1 FreeSans 800 0 0 0 Cin
port 1 n default bidirectional
flabel metal4 2 210 62 270 1 FreeSans 800 0 0 0 Cout
port 2 n default bidirectional
flabel metal1 2 1850 62 1910 1 FreeSans 800 0 0 0 VPWR
port 3 n power bidirectional
flabel metal1 2 -30 62 30 1 FreeSans 800 0 0 0 VGND
port 4 n ground bidirectional
<< properties >>
string FIXED_BBOX 0 0 7171 1880
string LEFclass CORE
string LEFsite unitasc
<< end >>
