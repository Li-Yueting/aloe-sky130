VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO sky130_asc_pnp_05v5_W3p40L3p40_8
  CLASS CORE ;
  FOREIGN sky130_asc_pnp_05v5_W3p40L3p40_8 ;
  ORIGIN 0.000 0.000 ;
  SIZE 54.500 BY 9.400 ;
  SITE unitasc ;
  PIN Emitter
    DIRECTION INOUT ;
    ANTENNADIFFAREA 92.479996 ;
    PORT
      LAYER li1 ;
        RECT 2.065 2.965 5.535 6.435 ;
        RECT 8.765 2.965 12.235 6.435 ;
        RECT 15.465 2.965 18.935 6.435 ;
        RECT 22.165 2.965 25.635 6.435 ;
        RECT 28.865 2.965 32.335 6.435 ;
        RECT 35.565 2.965 39.035 6.435 ;
        RECT 42.265 2.965 45.735 6.435 ;
        RECT 48.965 2.965 52.435 6.435 ;
      LAYER mcon ;
        RECT 2.430 5.830 2.600 6.000 ;
        RECT 2.930 5.830 3.100 6.000 ;
        RECT 3.430 5.830 3.600 6.000 ;
        RECT 3.930 5.830 4.100 6.000 ;
        RECT 4.430 5.830 4.600 6.000 ;
        RECT 4.930 5.830 5.100 6.000 ;
        RECT 2.430 5.330 2.600 5.500 ;
        RECT 2.930 5.330 3.100 5.500 ;
        RECT 3.430 5.330 3.600 5.500 ;
        RECT 3.930 5.330 4.100 5.500 ;
        RECT 4.430 5.330 4.600 5.500 ;
        RECT 4.930 5.330 5.100 5.500 ;
        RECT 2.430 4.830 2.600 5.000 ;
        RECT 2.930 4.830 3.100 5.000 ;
        RECT 3.430 4.830 3.600 5.000 ;
        RECT 3.930 4.830 4.100 5.000 ;
        RECT 4.430 4.830 4.600 5.000 ;
        RECT 4.930 4.830 5.100 5.000 ;
        RECT 2.430 4.330 2.600 4.500 ;
        RECT 2.930 4.330 3.100 4.500 ;
        RECT 3.430 4.330 3.600 4.500 ;
        RECT 3.930 4.330 4.100 4.500 ;
        RECT 4.430 4.330 4.600 4.500 ;
        RECT 4.930 4.330 5.100 4.500 ;
        RECT 2.430 3.830 2.600 4.000 ;
        RECT 2.930 3.830 3.100 4.000 ;
        RECT 3.430 3.830 3.600 4.000 ;
        RECT 3.930 3.830 4.100 4.000 ;
        RECT 4.430 3.830 4.600 4.000 ;
        RECT 4.930 3.830 5.100 4.000 ;
        RECT 2.430 3.330 2.600 3.500 ;
        RECT 2.930 3.330 3.100 3.500 ;
        RECT 3.430 3.330 3.600 3.500 ;
        RECT 3.930 3.330 4.100 3.500 ;
        RECT 4.430 3.330 4.600 3.500 ;
        RECT 4.930 3.330 5.100 3.500 ;
        RECT 9.130 5.830 9.300 6.000 ;
        RECT 9.630 5.830 9.800 6.000 ;
        RECT 10.130 5.830 10.300 6.000 ;
        RECT 10.630 5.830 10.800 6.000 ;
        RECT 11.130 5.830 11.300 6.000 ;
        RECT 11.630 5.830 11.800 6.000 ;
        RECT 9.130 5.330 9.300 5.500 ;
        RECT 9.630 5.330 9.800 5.500 ;
        RECT 10.130 5.330 10.300 5.500 ;
        RECT 10.630 5.330 10.800 5.500 ;
        RECT 11.130 5.330 11.300 5.500 ;
        RECT 11.630 5.330 11.800 5.500 ;
        RECT 9.130 4.830 9.300 5.000 ;
        RECT 9.630 4.830 9.800 5.000 ;
        RECT 10.130 4.830 10.300 5.000 ;
        RECT 10.630 4.830 10.800 5.000 ;
        RECT 11.130 4.830 11.300 5.000 ;
        RECT 11.630 4.830 11.800 5.000 ;
        RECT 9.130 4.330 9.300 4.500 ;
        RECT 9.630 4.330 9.800 4.500 ;
        RECT 10.130 4.330 10.300 4.500 ;
        RECT 10.630 4.330 10.800 4.500 ;
        RECT 11.130 4.330 11.300 4.500 ;
        RECT 11.630 4.330 11.800 4.500 ;
        RECT 9.130 3.830 9.300 4.000 ;
        RECT 9.630 3.830 9.800 4.000 ;
        RECT 10.130 3.830 10.300 4.000 ;
        RECT 10.630 3.830 10.800 4.000 ;
        RECT 11.130 3.830 11.300 4.000 ;
        RECT 11.630 3.830 11.800 4.000 ;
        RECT 9.130 3.330 9.300 3.500 ;
        RECT 9.630 3.330 9.800 3.500 ;
        RECT 10.130 3.330 10.300 3.500 ;
        RECT 10.630 3.330 10.800 3.500 ;
        RECT 11.130 3.330 11.300 3.500 ;
        RECT 11.630 3.330 11.800 3.500 ;
        RECT 15.830 5.830 16.000 6.000 ;
        RECT 16.330 5.830 16.500 6.000 ;
        RECT 16.830 5.830 17.000 6.000 ;
        RECT 17.330 5.830 17.500 6.000 ;
        RECT 17.830 5.830 18.000 6.000 ;
        RECT 18.330 5.830 18.500 6.000 ;
        RECT 15.830 5.330 16.000 5.500 ;
        RECT 16.330 5.330 16.500 5.500 ;
        RECT 16.830 5.330 17.000 5.500 ;
        RECT 17.330 5.330 17.500 5.500 ;
        RECT 17.830 5.330 18.000 5.500 ;
        RECT 18.330 5.330 18.500 5.500 ;
        RECT 15.830 4.830 16.000 5.000 ;
        RECT 16.330 4.830 16.500 5.000 ;
        RECT 16.830 4.830 17.000 5.000 ;
        RECT 17.330 4.830 17.500 5.000 ;
        RECT 17.830 4.830 18.000 5.000 ;
        RECT 18.330 4.830 18.500 5.000 ;
        RECT 15.830 4.330 16.000 4.500 ;
        RECT 16.330 4.330 16.500 4.500 ;
        RECT 16.830 4.330 17.000 4.500 ;
        RECT 17.330 4.330 17.500 4.500 ;
        RECT 17.830 4.330 18.000 4.500 ;
        RECT 18.330 4.330 18.500 4.500 ;
        RECT 15.830 3.830 16.000 4.000 ;
        RECT 16.330 3.830 16.500 4.000 ;
        RECT 16.830 3.830 17.000 4.000 ;
        RECT 17.330 3.830 17.500 4.000 ;
        RECT 17.830 3.830 18.000 4.000 ;
        RECT 18.330 3.830 18.500 4.000 ;
        RECT 15.830 3.330 16.000 3.500 ;
        RECT 16.330 3.330 16.500 3.500 ;
        RECT 16.830 3.330 17.000 3.500 ;
        RECT 17.330 3.330 17.500 3.500 ;
        RECT 17.830 3.330 18.000 3.500 ;
        RECT 18.330 3.330 18.500 3.500 ;
        RECT 22.530 5.830 22.700 6.000 ;
        RECT 23.030 5.830 23.200 6.000 ;
        RECT 23.530 5.830 23.700 6.000 ;
        RECT 24.030 5.830 24.200 6.000 ;
        RECT 24.530 5.830 24.700 6.000 ;
        RECT 25.030 5.830 25.200 6.000 ;
        RECT 22.530 5.330 22.700 5.500 ;
        RECT 23.030 5.330 23.200 5.500 ;
        RECT 23.530 5.330 23.700 5.500 ;
        RECT 24.030 5.330 24.200 5.500 ;
        RECT 24.530 5.330 24.700 5.500 ;
        RECT 25.030 5.330 25.200 5.500 ;
        RECT 22.530 4.830 22.700 5.000 ;
        RECT 23.030 4.830 23.200 5.000 ;
        RECT 23.530 4.830 23.700 5.000 ;
        RECT 24.030 4.830 24.200 5.000 ;
        RECT 24.530 4.830 24.700 5.000 ;
        RECT 25.030 4.830 25.200 5.000 ;
        RECT 22.530 4.330 22.700 4.500 ;
        RECT 23.030 4.330 23.200 4.500 ;
        RECT 23.530 4.330 23.700 4.500 ;
        RECT 24.030 4.330 24.200 4.500 ;
        RECT 24.530 4.330 24.700 4.500 ;
        RECT 25.030 4.330 25.200 4.500 ;
        RECT 22.530 3.830 22.700 4.000 ;
        RECT 23.030 3.830 23.200 4.000 ;
        RECT 23.530 3.830 23.700 4.000 ;
        RECT 24.030 3.830 24.200 4.000 ;
        RECT 24.530 3.830 24.700 4.000 ;
        RECT 25.030 3.830 25.200 4.000 ;
        RECT 22.530 3.330 22.700 3.500 ;
        RECT 23.030 3.330 23.200 3.500 ;
        RECT 23.530 3.330 23.700 3.500 ;
        RECT 24.030 3.330 24.200 3.500 ;
        RECT 24.530 3.330 24.700 3.500 ;
        RECT 25.030 3.330 25.200 3.500 ;
        RECT 29.230 5.830 29.400 6.000 ;
        RECT 29.730 5.830 29.900 6.000 ;
        RECT 30.230 5.830 30.400 6.000 ;
        RECT 30.730 5.830 30.900 6.000 ;
        RECT 31.230 5.830 31.400 6.000 ;
        RECT 31.730 5.830 31.900 6.000 ;
        RECT 29.230 5.330 29.400 5.500 ;
        RECT 29.730 5.330 29.900 5.500 ;
        RECT 30.230 5.330 30.400 5.500 ;
        RECT 30.730 5.330 30.900 5.500 ;
        RECT 31.230 5.330 31.400 5.500 ;
        RECT 31.730 5.330 31.900 5.500 ;
        RECT 29.230 4.830 29.400 5.000 ;
        RECT 29.730 4.830 29.900 5.000 ;
        RECT 30.230 4.830 30.400 5.000 ;
        RECT 30.730 4.830 30.900 5.000 ;
        RECT 31.230 4.830 31.400 5.000 ;
        RECT 31.730 4.830 31.900 5.000 ;
        RECT 29.230 4.330 29.400 4.500 ;
        RECT 29.730 4.330 29.900 4.500 ;
        RECT 30.230 4.330 30.400 4.500 ;
        RECT 30.730 4.330 30.900 4.500 ;
        RECT 31.230 4.330 31.400 4.500 ;
        RECT 31.730 4.330 31.900 4.500 ;
        RECT 29.230 3.830 29.400 4.000 ;
        RECT 29.730 3.830 29.900 4.000 ;
        RECT 30.230 3.830 30.400 4.000 ;
        RECT 30.730 3.830 30.900 4.000 ;
        RECT 31.230 3.830 31.400 4.000 ;
        RECT 31.730 3.830 31.900 4.000 ;
        RECT 29.230 3.330 29.400 3.500 ;
        RECT 29.730 3.330 29.900 3.500 ;
        RECT 30.230 3.330 30.400 3.500 ;
        RECT 30.730 3.330 30.900 3.500 ;
        RECT 31.230 3.330 31.400 3.500 ;
        RECT 31.730 3.330 31.900 3.500 ;
        RECT 35.930 5.830 36.100 6.000 ;
        RECT 36.430 5.830 36.600 6.000 ;
        RECT 36.930 5.830 37.100 6.000 ;
        RECT 37.430 5.830 37.600 6.000 ;
        RECT 37.930 5.830 38.100 6.000 ;
        RECT 38.430 5.830 38.600 6.000 ;
        RECT 35.930 5.330 36.100 5.500 ;
        RECT 36.430 5.330 36.600 5.500 ;
        RECT 36.930 5.330 37.100 5.500 ;
        RECT 37.430 5.330 37.600 5.500 ;
        RECT 37.930 5.330 38.100 5.500 ;
        RECT 38.430 5.330 38.600 5.500 ;
        RECT 35.930 4.830 36.100 5.000 ;
        RECT 36.430 4.830 36.600 5.000 ;
        RECT 36.930 4.830 37.100 5.000 ;
        RECT 37.430 4.830 37.600 5.000 ;
        RECT 37.930 4.830 38.100 5.000 ;
        RECT 38.430 4.830 38.600 5.000 ;
        RECT 35.930 4.330 36.100 4.500 ;
        RECT 36.430 4.330 36.600 4.500 ;
        RECT 36.930 4.330 37.100 4.500 ;
        RECT 37.430 4.330 37.600 4.500 ;
        RECT 37.930 4.330 38.100 4.500 ;
        RECT 38.430 4.330 38.600 4.500 ;
        RECT 35.930 3.830 36.100 4.000 ;
        RECT 36.430 3.830 36.600 4.000 ;
        RECT 36.930 3.830 37.100 4.000 ;
        RECT 37.430 3.830 37.600 4.000 ;
        RECT 37.930 3.830 38.100 4.000 ;
        RECT 38.430 3.830 38.600 4.000 ;
        RECT 35.930 3.330 36.100 3.500 ;
        RECT 36.430 3.330 36.600 3.500 ;
        RECT 36.930 3.330 37.100 3.500 ;
        RECT 37.430 3.330 37.600 3.500 ;
        RECT 37.930 3.330 38.100 3.500 ;
        RECT 38.430 3.330 38.600 3.500 ;
        RECT 42.630 5.830 42.800 6.000 ;
        RECT 43.130 5.830 43.300 6.000 ;
        RECT 43.630 5.830 43.800 6.000 ;
        RECT 44.130 5.830 44.300 6.000 ;
        RECT 44.630 5.830 44.800 6.000 ;
        RECT 45.130 5.830 45.300 6.000 ;
        RECT 42.630 5.330 42.800 5.500 ;
        RECT 43.130 5.330 43.300 5.500 ;
        RECT 43.630 5.330 43.800 5.500 ;
        RECT 44.130 5.330 44.300 5.500 ;
        RECT 44.630 5.330 44.800 5.500 ;
        RECT 45.130 5.330 45.300 5.500 ;
        RECT 42.630 4.830 42.800 5.000 ;
        RECT 43.130 4.830 43.300 5.000 ;
        RECT 43.630 4.830 43.800 5.000 ;
        RECT 44.130 4.830 44.300 5.000 ;
        RECT 44.630 4.830 44.800 5.000 ;
        RECT 45.130 4.830 45.300 5.000 ;
        RECT 42.630 4.330 42.800 4.500 ;
        RECT 43.130 4.330 43.300 4.500 ;
        RECT 43.630 4.330 43.800 4.500 ;
        RECT 44.130 4.330 44.300 4.500 ;
        RECT 44.630 4.330 44.800 4.500 ;
        RECT 45.130 4.330 45.300 4.500 ;
        RECT 42.630 3.830 42.800 4.000 ;
        RECT 43.130 3.830 43.300 4.000 ;
        RECT 43.630 3.830 43.800 4.000 ;
        RECT 44.130 3.830 44.300 4.000 ;
        RECT 44.630 3.830 44.800 4.000 ;
        RECT 45.130 3.830 45.300 4.000 ;
        RECT 42.630 3.330 42.800 3.500 ;
        RECT 43.130 3.330 43.300 3.500 ;
        RECT 43.630 3.330 43.800 3.500 ;
        RECT 44.130 3.330 44.300 3.500 ;
        RECT 44.630 3.330 44.800 3.500 ;
        RECT 45.130 3.330 45.300 3.500 ;
        RECT 49.330 5.830 49.500 6.000 ;
        RECT 49.830 5.830 50.000 6.000 ;
        RECT 50.330 5.830 50.500 6.000 ;
        RECT 50.830 5.830 51.000 6.000 ;
        RECT 51.330 5.830 51.500 6.000 ;
        RECT 51.830 5.830 52.000 6.000 ;
        RECT 49.330 5.330 49.500 5.500 ;
        RECT 49.830 5.330 50.000 5.500 ;
        RECT 50.330 5.330 50.500 5.500 ;
        RECT 50.830 5.330 51.000 5.500 ;
        RECT 51.330 5.330 51.500 5.500 ;
        RECT 51.830 5.330 52.000 5.500 ;
        RECT 49.330 4.830 49.500 5.000 ;
        RECT 49.830 4.830 50.000 5.000 ;
        RECT 50.330 4.830 50.500 5.000 ;
        RECT 50.830 4.830 51.000 5.000 ;
        RECT 51.330 4.830 51.500 5.000 ;
        RECT 51.830 4.830 52.000 5.000 ;
        RECT 49.330 4.330 49.500 4.500 ;
        RECT 49.830 4.330 50.000 4.500 ;
        RECT 50.330 4.330 50.500 4.500 ;
        RECT 50.830 4.330 51.000 4.500 ;
        RECT 51.330 4.330 51.500 4.500 ;
        RECT 51.830 4.330 52.000 4.500 ;
        RECT 49.330 3.830 49.500 4.000 ;
        RECT 49.830 3.830 50.000 4.000 ;
        RECT 50.330 3.830 50.500 4.000 ;
        RECT 50.830 3.830 51.000 4.000 ;
        RECT 51.330 3.830 51.500 4.000 ;
        RECT 51.830 3.830 52.000 4.000 ;
        RECT 49.330 3.330 49.500 3.500 ;
        RECT 49.830 3.330 50.000 3.500 ;
        RECT 50.330 3.330 50.500 3.500 ;
        RECT 50.830 3.330 51.000 3.500 ;
        RECT 51.330 3.330 51.500 3.500 ;
        RECT 51.830 3.330 52.000 3.500 ;
      LAYER met1 ;
        RECT 2.270 3.170 52.230 6.230 ;
    END
  END Emitter
  PIN Base
    DIRECTION INOUT ;
    ANTENNAGATEAREA 213.831192 ;
    ANTENNADIFFAREA 51.264000 ;
    PORT
      LAYER li1 ;
        RECT 1.395 6.745 6.205 7.105 ;
        RECT 1.395 2.655 1.755 6.745 ;
        RECT 5.845 2.655 6.205 6.745 ;
        RECT 1.395 2.295 6.205 2.655 ;
        RECT 8.095 6.745 12.905 7.105 ;
        RECT 8.095 2.655 8.455 6.745 ;
        RECT 12.545 2.655 12.905 6.745 ;
        RECT 8.095 2.295 12.905 2.655 ;
        RECT 14.795 6.745 19.605 7.105 ;
        RECT 14.795 2.655 15.155 6.745 ;
        RECT 19.245 2.655 19.605 6.745 ;
        RECT 14.795 2.295 19.605 2.655 ;
        RECT 21.495 6.745 26.305 7.105 ;
        RECT 21.495 2.655 21.855 6.745 ;
        RECT 25.945 2.655 26.305 6.745 ;
        RECT 21.495 2.295 26.305 2.655 ;
        RECT 28.195 6.745 33.005 7.105 ;
        RECT 28.195 2.655 28.555 6.745 ;
        RECT 32.645 2.655 33.005 6.745 ;
        RECT 28.195 2.295 33.005 2.655 ;
        RECT 34.895 6.745 39.705 7.105 ;
        RECT 34.895 2.655 35.255 6.745 ;
        RECT 39.345 2.655 39.705 6.745 ;
        RECT 34.895 2.295 39.705 2.655 ;
        RECT 41.595 6.745 46.405 7.105 ;
        RECT 41.595 2.655 41.955 6.745 ;
        RECT 46.045 2.655 46.405 6.745 ;
        RECT 41.595 2.295 46.405 2.655 ;
        RECT 48.295 6.745 53.105 7.105 ;
        RECT 48.295 2.655 48.655 6.745 ;
        RECT 52.745 2.655 53.105 6.745 ;
        RECT 48.295 2.295 53.105 2.655 ;
      LAYER mcon ;
        RECT 1.500 6.850 1.670 7.020 ;
        RECT 1.950 6.850 2.120 7.020 ;
        RECT 2.400 6.850 2.570 7.020 ;
        RECT 2.850 6.850 3.020 7.020 ;
        RECT 3.300 6.850 3.470 7.020 ;
        RECT 3.750 6.850 3.920 7.020 ;
        RECT 4.200 6.850 4.370 7.020 ;
        RECT 4.650 6.850 4.820 7.020 ;
        RECT 5.100 6.850 5.270 7.020 ;
        RECT 5.550 6.850 5.720 7.020 ;
        RECT 6.000 6.850 6.170 7.020 ;
        RECT 8.200 6.850 8.370 7.020 ;
        RECT 8.650 6.850 8.820 7.020 ;
        RECT 9.100 6.850 9.270 7.020 ;
        RECT 9.550 6.850 9.720 7.020 ;
        RECT 10.000 6.850 10.170 7.020 ;
        RECT 10.450 6.850 10.620 7.020 ;
        RECT 10.900 6.850 11.070 7.020 ;
        RECT 11.350 6.850 11.520 7.020 ;
        RECT 11.800 6.850 11.970 7.020 ;
        RECT 12.250 6.850 12.420 7.020 ;
        RECT 12.700 6.850 12.870 7.020 ;
        RECT 14.900 6.850 15.070 7.020 ;
        RECT 15.350 6.850 15.520 7.020 ;
        RECT 15.800 6.850 15.970 7.020 ;
        RECT 16.250 6.850 16.420 7.020 ;
        RECT 16.700 6.850 16.870 7.020 ;
        RECT 17.150 6.850 17.320 7.020 ;
        RECT 17.600 6.850 17.770 7.020 ;
        RECT 18.050 6.850 18.220 7.020 ;
        RECT 18.500 6.850 18.670 7.020 ;
        RECT 18.950 6.850 19.120 7.020 ;
        RECT 19.400 6.850 19.570 7.020 ;
        RECT 21.600 6.850 21.770 7.020 ;
        RECT 22.050 6.850 22.220 7.020 ;
        RECT 22.500 6.850 22.670 7.020 ;
        RECT 22.950 6.850 23.120 7.020 ;
        RECT 23.400 6.850 23.570 7.020 ;
        RECT 23.850 6.850 24.020 7.020 ;
        RECT 24.300 6.850 24.470 7.020 ;
        RECT 24.750 6.850 24.920 7.020 ;
        RECT 25.200 6.850 25.370 7.020 ;
        RECT 25.650 6.850 25.820 7.020 ;
        RECT 26.100 6.850 26.270 7.020 ;
        RECT 28.300 6.850 28.470 7.020 ;
        RECT 28.750 6.850 28.920 7.020 ;
        RECT 29.200 6.850 29.370 7.020 ;
        RECT 29.650 6.850 29.820 7.020 ;
        RECT 30.100 6.850 30.270 7.020 ;
        RECT 30.550 6.850 30.720 7.020 ;
        RECT 31.000 6.850 31.170 7.020 ;
        RECT 31.450 6.850 31.620 7.020 ;
        RECT 31.900 6.850 32.070 7.020 ;
        RECT 32.350 6.850 32.520 7.020 ;
        RECT 32.800 6.850 32.970 7.020 ;
        RECT 35.000 6.850 35.170 7.020 ;
        RECT 35.450 6.850 35.620 7.020 ;
        RECT 35.900 6.850 36.070 7.020 ;
        RECT 36.350 6.850 36.520 7.020 ;
        RECT 36.800 6.850 36.970 7.020 ;
        RECT 37.250 6.850 37.420 7.020 ;
        RECT 37.700 6.850 37.870 7.020 ;
        RECT 38.150 6.850 38.320 7.020 ;
        RECT 38.600 6.850 38.770 7.020 ;
        RECT 39.050 6.850 39.220 7.020 ;
        RECT 39.500 6.850 39.670 7.020 ;
        RECT 41.700 6.850 41.870 7.020 ;
        RECT 42.150 6.850 42.320 7.020 ;
        RECT 42.600 6.850 42.770 7.020 ;
        RECT 43.050 6.850 43.220 7.020 ;
        RECT 43.500 6.850 43.670 7.020 ;
        RECT 43.950 6.850 44.120 7.020 ;
        RECT 44.400 6.850 44.570 7.020 ;
        RECT 44.850 6.850 45.020 7.020 ;
        RECT 45.300 6.850 45.470 7.020 ;
        RECT 45.750 6.850 45.920 7.020 ;
        RECT 46.200 6.850 46.370 7.020 ;
        RECT 48.400 6.850 48.570 7.020 ;
        RECT 48.850 6.850 49.020 7.020 ;
        RECT 49.300 6.850 49.470 7.020 ;
        RECT 49.750 6.850 49.920 7.020 ;
        RECT 50.200 6.850 50.370 7.020 ;
        RECT 50.650 6.850 50.820 7.020 ;
        RECT 51.100 6.850 51.270 7.020 ;
        RECT 51.550 6.850 51.720 7.020 ;
        RECT 52.000 6.850 52.170 7.020 ;
        RECT 52.450 6.850 52.620 7.020 ;
        RECT 52.900 6.850 53.070 7.020 ;
      LAYER met1 ;
        RECT 1.400 6.750 53.100 7.100 ;
    END
  END Base
  PIN Collector
    DIRECTION INOUT ;
    ANTENNADIFFAREA 107.630394 ;
    PORT
      LAYER pwell ;
        RECT 0.450 7.285 54.050 8.050 ;
        RECT 0.450 2.115 1.215 7.285 ;
        RECT 6.385 2.115 7.915 7.285 ;
        RECT 13.085 2.115 14.615 7.285 ;
        RECT 19.785 2.115 21.315 7.285 ;
        RECT 26.485 2.115 28.015 7.285 ;
        RECT 33.185 2.115 34.715 7.285 ;
        RECT 39.885 2.115 41.415 7.285 ;
        RECT 46.585 2.115 48.115 7.285 ;
        RECT 53.285 2.115 54.050 7.285 ;
        RECT 0.450 1.350 54.050 2.115 ;
      LAYER li1 ;
        RECT 0.580 7.425 53.920 7.920 ;
        RECT 0.580 1.975 1.075 7.425 ;
        RECT 6.525 1.975 7.775 7.425 ;
        RECT 13.225 1.975 14.475 7.425 ;
        RECT 19.925 1.975 21.175 7.425 ;
        RECT 26.625 1.975 27.875 7.425 ;
        RECT 33.325 1.975 34.575 7.425 ;
        RECT 40.025 1.975 41.275 7.425 ;
        RECT 46.725 1.975 47.975 7.425 ;
        RECT 53.425 1.975 53.920 7.425 ;
        RECT 0.580 1.480 53.920 1.975 ;
      LAYER mcon ;
        RECT 0.680 7.650 0.850 7.820 ;
        RECT 1.130 7.650 1.300 7.820 ;
        RECT 1.580 7.650 1.750 7.820 ;
        RECT 2.030 7.650 2.200 7.820 ;
        RECT 2.480 7.650 2.650 7.820 ;
        RECT 2.930 7.650 3.100 7.820 ;
        RECT 3.380 7.650 3.550 7.820 ;
        RECT 3.830 7.650 4.000 7.820 ;
        RECT 4.280 7.650 4.450 7.820 ;
        RECT 4.730 7.650 4.900 7.820 ;
        RECT 5.180 7.650 5.350 7.820 ;
        RECT 5.630 7.650 5.800 7.820 ;
        RECT 6.080 7.650 6.250 7.820 ;
        RECT 6.530 7.650 6.700 7.820 ;
        RECT 7.380 7.650 7.550 7.820 ;
        RECT 7.830 7.650 8.000 7.820 ;
        RECT 8.280 7.650 8.450 7.820 ;
        RECT 8.730 7.650 8.900 7.820 ;
        RECT 9.180 7.650 9.350 7.820 ;
        RECT 9.630 7.650 9.800 7.820 ;
        RECT 10.080 7.650 10.250 7.820 ;
        RECT 10.530 7.650 10.700 7.820 ;
        RECT 10.980 7.650 11.150 7.820 ;
        RECT 11.430 7.650 11.600 7.820 ;
        RECT 11.880 7.650 12.050 7.820 ;
        RECT 12.330 7.650 12.500 7.820 ;
        RECT 12.780 7.650 12.950 7.820 ;
        RECT 13.230 7.650 13.400 7.820 ;
        RECT 14.080 7.650 14.250 7.820 ;
        RECT 14.530 7.650 14.700 7.820 ;
        RECT 14.980 7.650 15.150 7.820 ;
        RECT 15.430 7.650 15.600 7.820 ;
        RECT 15.880 7.650 16.050 7.820 ;
        RECT 16.330 7.650 16.500 7.820 ;
        RECT 16.780 7.650 16.950 7.820 ;
        RECT 17.230 7.650 17.400 7.820 ;
        RECT 17.680 7.650 17.850 7.820 ;
        RECT 18.130 7.650 18.300 7.820 ;
        RECT 18.580 7.650 18.750 7.820 ;
        RECT 19.030 7.650 19.200 7.820 ;
        RECT 19.480 7.650 19.650 7.820 ;
        RECT 19.930 7.650 20.100 7.820 ;
        RECT 20.780 7.650 20.950 7.820 ;
        RECT 21.230 7.650 21.400 7.820 ;
        RECT 21.680 7.650 21.850 7.820 ;
        RECT 22.130 7.650 22.300 7.820 ;
        RECT 22.580 7.650 22.750 7.820 ;
        RECT 23.030 7.650 23.200 7.820 ;
        RECT 23.480 7.650 23.650 7.820 ;
        RECT 23.930 7.650 24.100 7.820 ;
        RECT 24.380 7.650 24.550 7.820 ;
        RECT 24.830 7.650 25.000 7.820 ;
        RECT 25.280 7.650 25.450 7.820 ;
        RECT 25.730 7.650 25.900 7.820 ;
        RECT 26.180 7.650 26.350 7.820 ;
        RECT 26.630 7.650 26.800 7.820 ;
        RECT 27.480 7.650 27.650 7.820 ;
        RECT 27.930 7.650 28.100 7.820 ;
        RECT 28.380 7.650 28.550 7.820 ;
        RECT 28.830 7.650 29.000 7.820 ;
        RECT 29.280 7.650 29.450 7.820 ;
        RECT 29.730 7.650 29.900 7.820 ;
        RECT 30.180 7.650 30.350 7.820 ;
        RECT 30.630 7.650 30.800 7.820 ;
        RECT 31.080 7.650 31.250 7.820 ;
        RECT 31.530 7.650 31.700 7.820 ;
        RECT 31.980 7.650 32.150 7.820 ;
        RECT 32.430 7.650 32.600 7.820 ;
        RECT 32.880 7.650 33.050 7.820 ;
        RECT 33.330 7.650 33.500 7.820 ;
        RECT 34.180 7.650 34.350 7.820 ;
        RECT 34.630 7.650 34.800 7.820 ;
        RECT 35.080 7.650 35.250 7.820 ;
        RECT 35.530 7.650 35.700 7.820 ;
        RECT 35.980 7.650 36.150 7.820 ;
        RECT 36.430 7.650 36.600 7.820 ;
        RECT 36.880 7.650 37.050 7.820 ;
        RECT 37.330 7.650 37.500 7.820 ;
        RECT 37.780 7.650 37.950 7.820 ;
        RECT 38.230 7.650 38.400 7.820 ;
        RECT 38.680 7.650 38.850 7.820 ;
        RECT 39.130 7.650 39.300 7.820 ;
        RECT 39.580 7.650 39.750 7.820 ;
        RECT 40.030 7.650 40.200 7.820 ;
        RECT 40.880 7.650 41.050 7.820 ;
        RECT 41.330 7.650 41.500 7.820 ;
        RECT 41.780 7.650 41.950 7.820 ;
        RECT 42.230 7.650 42.400 7.820 ;
        RECT 42.680 7.650 42.850 7.820 ;
        RECT 43.130 7.650 43.300 7.820 ;
        RECT 43.580 7.650 43.750 7.820 ;
        RECT 44.030 7.650 44.200 7.820 ;
        RECT 44.480 7.650 44.650 7.820 ;
        RECT 44.930 7.650 45.100 7.820 ;
        RECT 45.380 7.650 45.550 7.820 ;
        RECT 45.830 7.650 46.000 7.820 ;
        RECT 46.280 7.650 46.450 7.820 ;
        RECT 46.730 7.650 46.900 7.820 ;
        RECT 47.580 7.650 47.750 7.820 ;
        RECT 48.030 7.650 48.200 7.820 ;
        RECT 48.480 7.650 48.650 7.820 ;
        RECT 48.930 7.650 49.100 7.820 ;
        RECT 49.380 7.650 49.550 7.820 ;
        RECT 49.830 7.650 50.000 7.820 ;
        RECT 50.280 7.650 50.450 7.820 ;
        RECT 50.730 7.650 50.900 7.820 ;
        RECT 51.180 7.650 51.350 7.820 ;
        RECT 51.630 7.650 51.800 7.820 ;
        RECT 52.080 7.650 52.250 7.820 ;
        RECT 52.530 7.650 52.700 7.820 ;
        RECT 52.980 7.650 53.150 7.820 ;
        RECT 53.430 7.650 53.600 7.820 ;
      LAYER met1 ;
        RECT 0.580 7.500 53.920 7.850 ;
    END
  END Collector
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER li1 ;
        RECT 0.450 9.250 54.050 9.550 ;
      LAYER mcon ;
        RECT 1.300 9.250 1.600 9.550 ;
        RECT 2.300 9.250 2.600 9.550 ;
        RECT 3.300 9.250 3.600 9.550 ;
        RECT 4.300 9.250 4.600 9.550 ;
        RECT 5.300 9.250 5.600 9.550 ;
        RECT 6.300 9.250 6.600 9.550 ;
        RECT 7.300 9.250 7.600 9.550 ;
        RECT 8.300 9.250 8.600 9.550 ;
        RECT 9.300 9.250 9.600 9.550 ;
        RECT 10.300 9.250 10.600 9.550 ;
        RECT 11.300 9.250 11.600 9.550 ;
        RECT 12.300 9.250 12.600 9.550 ;
        RECT 13.300 9.250 13.600 9.550 ;
        RECT 14.300 9.250 14.600 9.550 ;
        RECT 15.300 9.250 15.600 9.550 ;
        RECT 16.300 9.250 16.600 9.550 ;
        RECT 17.300 9.250 17.600 9.550 ;
        RECT 18.300 9.250 18.600 9.550 ;
        RECT 19.300 9.250 19.600 9.550 ;
        RECT 20.300 9.250 20.600 9.550 ;
        RECT 21.300 9.250 21.600 9.550 ;
        RECT 22.300 9.250 22.600 9.550 ;
        RECT 23.300 9.250 23.600 9.550 ;
        RECT 24.300 9.250 24.600 9.550 ;
        RECT 25.300 9.250 25.600 9.550 ;
        RECT 26.300 9.250 26.600 9.550 ;
        RECT 27.300 9.250 27.600 9.550 ;
        RECT 28.300 9.250 28.600 9.550 ;
        RECT 29.300 9.250 29.600 9.550 ;
        RECT 30.300 9.250 30.600 9.550 ;
        RECT 31.300 9.250 31.600 9.550 ;
        RECT 32.300 9.250 32.600 9.550 ;
        RECT 33.300 9.250 33.600 9.550 ;
        RECT 34.300 9.250 34.600 9.550 ;
        RECT 35.300 9.250 35.600 9.550 ;
        RECT 36.300 9.250 36.600 9.550 ;
        RECT 37.300 9.250 37.600 9.550 ;
        RECT 38.300 9.250 38.600 9.550 ;
        RECT 39.300 9.250 39.600 9.550 ;
        RECT 40.300 9.250 40.600 9.550 ;
        RECT 41.300 9.250 41.600 9.550 ;
        RECT 42.300 9.250 42.600 9.550 ;
        RECT 43.300 9.250 43.600 9.550 ;
        RECT 44.300 9.250 44.600 9.550 ;
        RECT 45.300 9.250 45.600 9.550 ;
        RECT 46.300 9.250 46.600 9.550 ;
        RECT 47.300 9.250 47.600 9.550 ;
        RECT 48.300 9.250 48.600 9.550 ;
        RECT 49.300 9.250 49.600 9.550 ;
        RECT 50.300 9.250 50.600 9.550 ;
        RECT 51.300 9.250 51.600 9.550 ;
        RECT 52.300 9.250 52.600 9.550 ;
        RECT 53.300 9.250 53.600 9.550 ;
      LAYER met1 ;
        RECT 0.450 9.100 54.050 9.700 ;
    END
  END VPWR
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER li1 ;
        RECT 0.450 -0.150 54.050 0.150 ;
      LAYER mcon ;
        RECT 1.300 -0.150 1.600 0.150 ;
        RECT 2.300 -0.150 2.600 0.150 ;
        RECT 3.300 -0.150 3.600 0.150 ;
        RECT 4.300 -0.150 4.600 0.150 ;
        RECT 5.300 -0.150 5.600 0.150 ;
        RECT 6.300 -0.150 6.600 0.150 ;
        RECT 7.300 -0.150 7.600 0.150 ;
        RECT 8.300 -0.150 8.600 0.150 ;
        RECT 9.300 -0.150 9.600 0.150 ;
        RECT 10.300 -0.150 10.600 0.150 ;
        RECT 11.300 -0.150 11.600 0.150 ;
        RECT 12.300 -0.150 12.600 0.150 ;
        RECT 13.300 -0.150 13.600 0.150 ;
        RECT 14.300 -0.150 14.600 0.150 ;
        RECT 15.300 -0.150 15.600 0.150 ;
        RECT 16.300 -0.150 16.600 0.150 ;
        RECT 17.300 -0.150 17.600 0.150 ;
        RECT 18.300 -0.150 18.600 0.150 ;
        RECT 19.300 -0.150 19.600 0.150 ;
        RECT 20.300 -0.150 20.600 0.150 ;
        RECT 21.300 -0.150 21.600 0.150 ;
        RECT 22.300 -0.150 22.600 0.150 ;
        RECT 23.300 -0.150 23.600 0.150 ;
        RECT 24.300 -0.150 24.600 0.150 ;
        RECT 25.300 -0.150 25.600 0.150 ;
        RECT 26.300 -0.150 26.600 0.150 ;
        RECT 27.300 -0.150 27.600 0.150 ;
        RECT 28.300 -0.150 28.600 0.150 ;
        RECT 29.300 -0.150 29.600 0.150 ;
        RECT 30.300 -0.150 30.600 0.150 ;
        RECT 31.300 -0.150 31.600 0.150 ;
        RECT 32.300 -0.150 32.600 0.150 ;
        RECT 33.300 -0.150 33.600 0.150 ;
        RECT 34.300 -0.150 34.600 0.150 ;
        RECT 35.300 -0.150 35.600 0.150 ;
        RECT 36.300 -0.150 36.600 0.150 ;
        RECT 37.300 -0.150 37.600 0.150 ;
        RECT 38.300 -0.150 38.600 0.150 ;
        RECT 39.300 -0.150 39.600 0.150 ;
        RECT 40.300 -0.150 40.600 0.150 ;
        RECT 41.300 -0.150 41.600 0.150 ;
        RECT 42.300 -0.150 42.600 0.150 ;
        RECT 43.300 -0.150 43.600 0.150 ;
        RECT 44.300 -0.150 44.600 0.150 ;
        RECT 45.300 -0.150 45.600 0.150 ;
        RECT 46.300 -0.150 46.600 0.150 ;
        RECT 47.300 -0.150 47.600 0.150 ;
        RECT 48.300 -0.150 48.600 0.150 ;
        RECT 49.300 -0.150 49.600 0.150 ;
        RECT 50.300 -0.150 50.600 0.150 ;
        RECT 51.300 -0.150 51.600 0.150 ;
        RECT 52.300 -0.150 52.600 0.150 ;
        RECT 53.300 -0.150 53.600 0.150 ;
      LAYER met1 ;
        RECT 0.450 -0.300 54.050 0.300 ;
    END
  END VGND
END sky130_asc_pnp_05v5_W3p40L3p40_8
END LIBRARY

