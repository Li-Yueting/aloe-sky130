VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO sky130_asc_pfet_01v8_lvt_60
  CLASS CORE ;
  FOREIGN sky130_asc_pfet_01v8_lvt_60 ;
  ORIGIN 0.000 0.000 ;
  SIZE 139.735 BY 9.400 ;
  SITE unitasc ;
  PIN GATE
    DIRECTION INOUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 774.000000 ;
    PORT
      LAYER li1 ;
        RECT 1.090 0.520 139.130 0.820 ;
    END
  END GATE
  PIN SOURCE
    DIRECTION INOUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 56.114998 ;
    PORT
      LAYER li1 ;
        RECT 1.390 8.450 139.130 8.650 ;
        RECT 3.615 1.755 3.785 8.450 ;
        RECT 8.195 1.755 8.365 8.450 ;
        RECT 12.775 1.755 12.945 8.450 ;
        RECT 17.355 1.755 17.525 8.450 ;
        RECT 21.935 1.755 22.105 8.450 ;
        RECT 26.515 1.755 26.685 8.450 ;
        RECT 31.095 1.755 31.265 8.450 ;
        RECT 35.675 1.755 35.845 8.450 ;
        RECT 40.255 1.755 40.425 8.450 ;
        RECT 44.835 1.755 45.005 8.450 ;
        RECT 49.415 1.755 49.585 8.450 ;
        RECT 53.995 1.755 54.165 8.450 ;
        RECT 58.575 1.755 58.745 8.450 ;
        RECT 63.155 1.755 63.325 8.450 ;
        RECT 67.735 1.755 67.905 8.450 ;
        RECT 72.315 1.755 72.485 8.450 ;
        RECT 76.895 1.755 77.065 8.450 ;
        RECT 81.475 1.755 81.645 8.450 ;
        RECT 86.055 1.755 86.225 8.450 ;
        RECT 90.635 1.755 90.805 8.450 ;
        RECT 95.215 1.755 95.385 8.450 ;
        RECT 99.795 1.755 99.965 8.450 ;
        RECT 104.375 1.755 104.545 8.450 ;
        RECT 108.955 1.755 109.125 8.450 ;
        RECT 113.535 1.755 113.705 8.450 ;
        RECT 118.115 1.755 118.285 8.450 ;
        RECT 122.695 1.755 122.865 8.450 ;
        RECT 127.275 1.755 127.445 8.450 ;
        RECT 131.855 1.755 132.025 8.450 ;
        RECT 136.435 1.755 136.605 8.450 ;
      LAYER mcon ;
        RECT 3.615 1.835 3.785 8.165 ;
        RECT 8.195 1.835 8.365 8.165 ;
        RECT 12.775 1.835 12.945 8.165 ;
        RECT 17.355 1.835 17.525 8.165 ;
        RECT 21.935 1.835 22.105 8.165 ;
        RECT 26.515 1.835 26.685 8.165 ;
        RECT 31.095 1.835 31.265 8.165 ;
        RECT 35.675 1.835 35.845 8.165 ;
        RECT 40.255 1.835 40.425 8.165 ;
        RECT 44.835 1.835 45.005 8.165 ;
        RECT 49.415 1.835 49.585 8.165 ;
        RECT 53.995 1.835 54.165 8.165 ;
        RECT 58.575 1.835 58.745 8.165 ;
        RECT 63.155 1.835 63.325 8.165 ;
        RECT 67.735 1.835 67.905 8.165 ;
        RECT 72.315 1.835 72.485 8.165 ;
        RECT 76.895 1.835 77.065 8.165 ;
        RECT 81.475 1.835 81.645 8.165 ;
        RECT 86.055 1.835 86.225 8.165 ;
        RECT 90.635 1.835 90.805 8.165 ;
        RECT 95.215 1.835 95.385 8.165 ;
        RECT 99.795 1.835 99.965 8.165 ;
        RECT 104.375 1.835 104.545 8.165 ;
        RECT 108.955 1.835 109.125 8.165 ;
        RECT 113.535 1.835 113.705 8.165 ;
        RECT 118.115 1.835 118.285 8.165 ;
        RECT 122.695 1.835 122.865 8.165 ;
        RECT 127.275 1.835 127.445 8.165 ;
        RECT 131.855 1.835 132.025 8.165 ;
        RECT 136.435 1.835 136.605 8.165 ;
      LAYER met1 ;
        RECT 3.585 1.775 3.815 8.225 ;
        RECT 8.165 1.775 8.395 8.225 ;
        RECT 12.745 1.775 12.975 8.225 ;
        RECT 17.325 1.775 17.555 8.225 ;
        RECT 21.905 1.775 22.135 8.225 ;
        RECT 26.485 1.775 26.715 8.225 ;
        RECT 31.065 1.775 31.295 8.225 ;
        RECT 35.645 1.775 35.875 8.225 ;
        RECT 40.225 1.775 40.455 8.225 ;
        RECT 44.805 1.775 45.035 8.225 ;
        RECT 49.385 1.775 49.615 8.225 ;
        RECT 53.965 1.775 54.195 8.225 ;
        RECT 58.545 1.775 58.775 8.225 ;
        RECT 63.125 1.775 63.355 8.225 ;
        RECT 67.705 1.775 67.935 8.225 ;
        RECT 72.285 1.775 72.515 8.225 ;
        RECT 76.865 1.775 77.095 8.225 ;
        RECT 81.445 1.775 81.675 8.225 ;
        RECT 86.025 1.775 86.255 8.225 ;
        RECT 90.605 1.775 90.835 8.225 ;
        RECT 95.185 1.775 95.415 8.225 ;
        RECT 99.765 1.775 99.995 8.225 ;
        RECT 104.345 1.775 104.575 8.225 ;
        RECT 108.925 1.775 109.155 8.225 ;
        RECT 113.505 1.775 113.735 8.225 ;
        RECT 118.085 1.775 118.315 8.225 ;
        RECT 122.665 1.775 122.895 8.225 ;
        RECT 127.245 1.775 127.475 8.225 ;
        RECT 131.825 1.775 132.055 8.225 ;
        RECT 136.405 1.775 136.635 8.225 ;
    END
  END SOURCE
  PIN DRAIN
    DIRECTION INOUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 57.985500 ;
    PORT
      LAYER li1 ;
        RECT 1.325 1.350 1.495 8.245 ;
        RECT 5.905 1.350 6.075 8.245 ;
        RECT 10.485 1.350 10.655 8.245 ;
        RECT 15.065 1.350 15.235 8.245 ;
        RECT 19.645 1.350 19.815 8.245 ;
        RECT 24.225 1.350 24.395 8.245 ;
        RECT 28.805 1.350 28.975 8.245 ;
        RECT 33.385 1.350 33.555 8.245 ;
        RECT 37.965 1.350 38.135 8.245 ;
        RECT 42.545 1.350 42.715 8.245 ;
        RECT 47.125 1.350 47.295 8.245 ;
        RECT 51.705 1.350 51.875 8.245 ;
        RECT 56.285 1.350 56.455 8.245 ;
        RECT 60.865 1.350 61.035 8.245 ;
        RECT 65.445 1.350 65.615 8.245 ;
        RECT 70.025 1.350 70.195 8.245 ;
        RECT 74.605 1.350 74.775 8.245 ;
        RECT 79.185 1.350 79.355 8.245 ;
        RECT 83.765 1.350 83.935 8.245 ;
        RECT 88.345 1.350 88.515 8.245 ;
        RECT 92.925 1.350 93.095 8.245 ;
        RECT 97.505 1.350 97.675 8.245 ;
        RECT 102.085 1.350 102.255 8.245 ;
        RECT 106.665 1.350 106.835 8.245 ;
        RECT 111.245 1.350 111.415 8.245 ;
        RECT 115.825 1.350 115.995 8.245 ;
        RECT 120.405 1.350 120.575 8.245 ;
        RECT 124.985 1.350 125.155 8.245 ;
        RECT 129.565 1.350 129.735 8.245 ;
        RECT 134.145 1.350 134.315 8.245 ;
        RECT 138.725 1.350 138.895 8.245 ;
        RECT 1.090 1.050 139.130 1.350 ;
      LAYER mcon ;
        RECT 1.325 1.835 1.495 8.165 ;
        RECT 5.905 1.835 6.075 8.165 ;
        RECT 10.485 1.835 10.655 8.165 ;
        RECT 15.065 1.835 15.235 8.165 ;
        RECT 19.645 1.835 19.815 8.165 ;
        RECT 24.225 1.835 24.395 8.165 ;
        RECT 28.805 1.835 28.975 8.165 ;
        RECT 33.385 1.835 33.555 8.165 ;
        RECT 37.965 1.835 38.135 8.165 ;
        RECT 42.545 1.835 42.715 8.165 ;
        RECT 47.125 1.835 47.295 8.165 ;
        RECT 51.705 1.835 51.875 8.165 ;
        RECT 56.285 1.835 56.455 8.165 ;
        RECT 60.865 1.835 61.035 8.165 ;
        RECT 65.445 1.835 65.615 8.165 ;
        RECT 70.025 1.835 70.195 8.165 ;
        RECT 74.605 1.835 74.775 8.165 ;
        RECT 79.185 1.835 79.355 8.165 ;
        RECT 83.765 1.835 83.935 8.165 ;
        RECT 88.345 1.835 88.515 8.165 ;
        RECT 92.925 1.835 93.095 8.165 ;
        RECT 97.505 1.835 97.675 8.165 ;
        RECT 102.085 1.835 102.255 8.165 ;
        RECT 106.665 1.835 106.835 8.165 ;
        RECT 111.245 1.835 111.415 8.165 ;
        RECT 115.825 1.835 115.995 8.165 ;
        RECT 120.405 1.835 120.575 8.165 ;
        RECT 124.985 1.835 125.155 8.165 ;
        RECT 129.565 1.835 129.735 8.165 ;
        RECT 134.145 1.835 134.315 8.165 ;
        RECT 138.725 1.835 138.895 8.165 ;
      LAYER met1 ;
        RECT 1.295 1.775 1.525 8.225 ;
        RECT 5.875 1.775 6.105 8.225 ;
        RECT 10.455 1.775 10.685 8.225 ;
        RECT 15.035 1.775 15.265 8.225 ;
        RECT 19.615 1.775 19.845 8.225 ;
        RECT 24.195 1.775 24.425 8.225 ;
        RECT 28.775 1.775 29.005 8.225 ;
        RECT 33.355 1.775 33.585 8.225 ;
        RECT 37.935 1.775 38.165 8.225 ;
        RECT 42.515 1.775 42.745 8.225 ;
        RECT 47.095 1.775 47.325 8.225 ;
        RECT 51.675 1.775 51.905 8.225 ;
        RECT 56.255 1.775 56.485 8.225 ;
        RECT 60.835 1.775 61.065 8.225 ;
        RECT 65.415 1.775 65.645 8.225 ;
        RECT 69.995 1.775 70.225 8.225 ;
        RECT 74.575 1.775 74.805 8.225 ;
        RECT 79.155 1.775 79.385 8.225 ;
        RECT 83.735 1.775 83.965 8.225 ;
        RECT 88.315 1.775 88.545 8.225 ;
        RECT 92.895 1.775 93.125 8.225 ;
        RECT 97.475 1.775 97.705 8.225 ;
        RECT 102.055 1.775 102.285 8.225 ;
        RECT 106.635 1.775 106.865 8.225 ;
        RECT 111.215 1.775 111.445 8.225 ;
        RECT 115.795 1.775 116.025 8.225 ;
        RECT 120.375 1.775 120.605 8.225 ;
        RECT 124.955 1.775 125.185 8.225 ;
        RECT 129.535 1.775 129.765 8.225 ;
        RECT 134.115 1.775 134.345 8.225 ;
        RECT 138.695 1.775 138.925 8.225 ;
    END
  END DRAIN
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT 0.600 8.535 139.130 9.700 ;
        RECT 0.600 1.470 139.135 8.535 ;
        RECT 1.085 1.465 139.135 1.470 ;
      LAYER li1 ;
        RECT 0.600 9.250 139.130 9.550 ;
        RECT 0.740 8.200 1.040 9.250 ;
        RECT 5.980 8.850 6.780 9.250 ;
        RECT 12.480 8.850 13.280 9.250 ;
        RECT 18.980 8.850 19.780 9.250 ;
        RECT 25.480 8.850 26.280 9.250 ;
        RECT 31.980 8.850 32.780 9.250 ;
        RECT 38.480 8.850 39.280 9.250 ;
        RECT 44.980 8.850 45.780 9.250 ;
        RECT 51.480 8.850 52.280 9.250 ;
        RECT 57.980 8.850 58.780 9.250 ;
        RECT 64.480 8.850 65.280 9.250 ;
        RECT 70.980 8.850 71.780 9.250 ;
        RECT 77.480 8.850 78.280 9.250 ;
        RECT 83.980 8.850 84.780 9.250 ;
        RECT 90.480 8.850 91.280 9.250 ;
        RECT 96.980 8.850 97.780 9.250 ;
        RECT 103.480 8.850 104.280 9.250 ;
        RECT 109.980 8.850 110.780 9.250 ;
        RECT 116.480 8.850 117.280 9.250 ;
        RECT 122.980 8.850 123.780 9.250 ;
        RECT 129.480 8.850 130.280 9.250 ;
      LAYER mcon ;
        RECT 1.940 9.250 2.240 9.550 ;
        RECT 3.940 9.250 4.240 9.550 ;
        RECT 5.940 9.250 6.240 9.550 ;
        RECT 7.940 9.250 8.240 9.550 ;
        RECT 9.940 9.250 10.240 9.550 ;
        RECT 11.940 9.250 12.240 9.550 ;
        RECT 13.940 9.250 14.240 9.550 ;
        RECT 15.940 9.250 16.240 9.550 ;
        RECT 17.940 9.250 18.240 9.550 ;
        RECT 19.940 9.250 20.240 9.550 ;
        RECT 21.940 9.250 22.240 9.550 ;
        RECT 23.940 9.250 24.240 9.550 ;
        RECT 25.940 9.250 26.240 9.550 ;
        RECT 27.940 9.250 28.240 9.550 ;
        RECT 29.940 9.250 30.240 9.550 ;
        RECT 31.940 9.250 32.240 9.550 ;
        RECT 33.940 9.250 34.240 9.550 ;
        RECT 35.940 9.250 36.240 9.550 ;
        RECT 37.940 9.250 38.240 9.550 ;
        RECT 39.940 9.250 40.240 9.550 ;
        RECT 41.940 9.250 42.240 9.550 ;
        RECT 43.940 9.250 44.240 9.550 ;
        RECT 45.940 9.250 46.240 9.550 ;
        RECT 47.940 9.250 48.240 9.550 ;
        RECT 49.940 9.250 50.240 9.550 ;
        RECT 51.940 9.250 52.240 9.550 ;
        RECT 53.940 9.250 54.240 9.550 ;
        RECT 55.940 9.250 56.240 9.550 ;
        RECT 57.940 9.250 58.240 9.550 ;
        RECT 59.940 9.250 60.240 9.550 ;
        RECT 61.940 9.250 62.240 9.550 ;
        RECT 63.940 9.250 64.240 9.550 ;
        RECT 65.940 9.250 66.240 9.550 ;
        RECT 67.940 9.250 68.240 9.550 ;
        RECT 69.940 9.250 70.240 9.550 ;
        RECT 71.940 9.250 72.240 9.550 ;
        RECT 73.940 9.250 74.240 9.550 ;
        RECT 75.940 9.250 76.240 9.550 ;
        RECT 77.940 9.250 78.240 9.550 ;
        RECT 79.940 9.250 80.240 9.550 ;
        RECT 81.940 9.250 82.240 9.550 ;
        RECT 83.940 9.250 84.240 9.550 ;
        RECT 85.940 9.250 86.240 9.550 ;
        RECT 87.940 9.250 88.240 9.550 ;
        RECT 89.940 9.250 90.240 9.550 ;
        RECT 91.940 9.250 92.240 9.550 ;
        RECT 93.940 9.250 94.240 9.550 ;
        RECT 95.940 9.250 96.240 9.550 ;
        RECT 97.940 9.250 98.240 9.550 ;
        RECT 99.940 9.250 100.240 9.550 ;
        RECT 101.940 9.250 102.240 9.550 ;
        RECT 103.940 9.250 104.240 9.550 ;
        RECT 105.940 9.250 106.240 9.550 ;
        RECT 107.940 9.250 108.240 9.550 ;
        RECT 109.940 9.250 110.240 9.550 ;
        RECT 111.940 9.250 112.240 9.550 ;
        RECT 113.940 9.250 114.240 9.550 ;
        RECT 115.940 9.250 116.240 9.550 ;
        RECT 117.940 9.250 118.240 9.550 ;
        RECT 119.940 9.250 120.240 9.550 ;
        RECT 121.940 9.250 122.240 9.550 ;
        RECT 123.940 9.250 124.240 9.550 ;
        RECT 125.940 9.250 126.240 9.550 ;
        RECT 127.940 9.250 128.240 9.550 ;
        RECT 129.940 9.250 130.240 9.550 ;
        RECT 131.940 9.250 132.240 9.550 ;
        RECT 133.940 9.250 134.240 9.550 ;
        RECT 135.940 9.250 136.240 9.550 ;
        RECT 137.940 9.250 138.240 9.550 ;
      LAYER met1 ;
        RECT 0.600 9.100 139.130 9.700 ;
    END
  END VPWR
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER li1 ;
        RECT 0.600 -0.150 139.130 0.150 ;
      LAYER mcon ;
        RECT 1.940 -0.150 2.240 0.150 ;
        RECT 3.940 -0.150 4.240 0.150 ;
        RECT 5.940 -0.150 6.240 0.150 ;
        RECT 7.940 -0.150 8.240 0.150 ;
        RECT 9.940 -0.150 10.240 0.150 ;
        RECT 11.940 -0.150 12.240 0.150 ;
        RECT 13.940 -0.150 14.240 0.150 ;
        RECT 15.940 -0.150 16.240 0.150 ;
        RECT 17.940 -0.150 18.240 0.150 ;
        RECT 19.940 -0.150 20.240 0.150 ;
        RECT 21.940 -0.150 22.240 0.150 ;
        RECT 23.940 -0.150 24.240 0.150 ;
        RECT 25.940 -0.150 26.240 0.150 ;
        RECT 27.940 -0.150 28.240 0.150 ;
        RECT 29.940 -0.150 30.240 0.150 ;
        RECT 31.940 -0.150 32.240 0.150 ;
        RECT 33.940 -0.150 34.240 0.150 ;
        RECT 35.940 -0.150 36.240 0.150 ;
        RECT 37.940 -0.150 38.240 0.150 ;
        RECT 39.940 -0.150 40.240 0.150 ;
        RECT 41.940 -0.150 42.240 0.150 ;
        RECT 43.940 -0.150 44.240 0.150 ;
        RECT 45.940 -0.150 46.240 0.150 ;
        RECT 47.940 -0.150 48.240 0.150 ;
        RECT 49.940 -0.150 50.240 0.150 ;
        RECT 51.940 -0.150 52.240 0.150 ;
        RECT 53.940 -0.150 54.240 0.150 ;
        RECT 55.940 -0.150 56.240 0.150 ;
        RECT 57.940 -0.150 58.240 0.150 ;
        RECT 59.940 -0.150 60.240 0.150 ;
        RECT 61.940 -0.150 62.240 0.150 ;
        RECT 63.940 -0.150 64.240 0.150 ;
        RECT 65.940 -0.150 66.240 0.150 ;
        RECT 67.940 -0.150 68.240 0.150 ;
        RECT 69.940 -0.150 70.240 0.150 ;
        RECT 71.940 -0.150 72.240 0.150 ;
        RECT 73.940 -0.150 74.240 0.150 ;
        RECT 75.940 -0.150 76.240 0.150 ;
        RECT 77.940 -0.150 78.240 0.150 ;
        RECT 79.940 -0.150 80.240 0.150 ;
        RECT 81.940 -0.150 82.240 0.150 ;
        RECT 83.940 -0.150 84.240 0.150 ;
        RECT 85.940 -0.150 86.240 0.150 ;
        RECT 87.940 -0.150 88.240 0.150 ;
        RECT 89.940 -0.150 90.240 0.150 ;
        RECT 91.940 -0.150 92.240 0.150 ;
        RECT 93.940 -0.150 94.240 0.150 ;
        RECT 95.940 -0.150 96.240 0.150 ;
        RECT 97.940 -0.150 98.240 0.150 ;
        RECT 99.940 -0.150 100.240 0.150 ;
        RECT 101.940 -0.150 102.240 0.150 ;
        RECT 103.940 -0.150 104.240 0.150 ;
        RECT 105.940 -0.150 106.240 0.150 ;
        RECT 107.940 -0.150 108.240 0.150 ;
        RECT 109.940 -0.150 110.240 0.150 ;
        RECT 111.940 -0.150 112.240 0.150 ;
        RECT 113.940 -0.150 114.240 0.150 ;
        RECT 115.940 -0.150 116.240 0.150 ;
        RECT 117.940 -0.150 118.240 0.150 ;
        RECT 119.940 -0.150 120.240 0.150 ;
        RECT 121.940 -0.150 122.240 0.150 ;
        RECT 123.940 -0.150 124.240 0.150 ;
        RECT 125.940 -0.150 126.240 0.150 ;
        RECT 127.940 -0.150 128.240 0.150 ;
        RECT 129.940 -0.150 130.240 0.150 ;
        RECT 131.940 -0.150 132.240 0.150 ;
        RECT 133.940 -0.150 134.240 0.150 ;
        RECT 135.940 -0.150 136.240 0.150 ;
        RECT 137.940 -0.150 138.240 0.150 ;
      LAYER met1 ;
        RECT 0.600 -0.300 139.130 0.300 ;
    END
  END VGND
END sky130_asc_pfet_01v8_lvt_60
END LIBRARY

