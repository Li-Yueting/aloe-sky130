.subckt sky130_fd_sc_hd__pfet GATE SOURCE DRAIN VPB VPWR VGND
X0 SOURCE GATE DRAIN VPB sky130_fd_pr__pfet_01v8_lvt w=6450000u l=2000000u
.ends

.subckt sky130_fd_sc_hd__nfet GATE SOURCE DRAIN VNB VPWR VGND
X0 SOURCE GATE DRAIN VNB sky130_fd_pr__nfet_01v8_lvt w=4000000u l=2000000u
.ends