magic
tech sky130A
magscale 1 2
timestamp 1652221618
<< nwell >>
rect 0 294 4350 1940
rect 98 293 4350 294
<< pmoslvt >>
rect 192 355 592 1645
rect 650 355 1050 1645
rect 1108 355 1508 1645
rect 1566 355 1966 1645
rect 2024 355 2424 1645
rect 2482 355 2882 1645
rect 2940 355 3340 1645
rect 3398 355 3798 1645
rect 3856 355 4256 1645
<< pdiff >>
rect 134 1633 192 1645
rect 134 367 146 1633
rect 180 367 192 1633
rect 134 355 192 367
rect 592 1633 650 1645
rect 592 367 604 1633
rect 638 367 650 1633
rect 592 355 650 367
rect 1050 1633 1108 1645
rect 1050 367 1062 1633
rect 1096 367 1108 1633
rect 1050 355 1108 367
rect 1508 1633 1566 1645
rect 1508 367 1520 1633
rect 1554 367 1566 1633
rect 1508 355 1566 367
rect 1966 1633 2024 1645
rect 1966 367 1978 1633
rect 2012 367 2024 1633
rect 1966 355 2024 367
rect 2424 1633 2482 1645
rect 2424 367 2436 1633
rect 2470 367 2482 1633
rect 2424 355 2482 367
rect 2882 1633 2940 1645
rect 2882 367 2894 1633
rect 2928 367 2940 1633
rect 2882 355 2940 367
rect 3340 1633 3398 1645
rect 3340 367 3352 1633
rect 3386 367 3398 1633
rect 3340 355 3398 367
rect 3798 1633 3856 1645
rect 3798 367 3810 1633
rect 3844 367 3856 1633
rect 3798 355 3856 367
rect 4256 1633 4314 1645
rect 4256 367 4268 1633
rect 4302 367 4314 1633
rect 4256 355 4314 367
<< pdiffc >>
rect 146 367 180 1633
rect 604 367 638 1633
rect 1062 367 1096 1633
rect 1520 367 1554 1633
rect 1978 367 2012 1633
rect 2436 367 2470 1633
rect 2894 367 2928 1633
rect 3352 367 3386 1633
rect 3810 367 3844 1633
rect 4268 367 4302 1633
<< nsubdiff >>
rect 38 1760 78 1800
rect 38 1680 78 1720
<< nsubdiffcont >>
rect 38 1720 78 1760
<< poly >>
rect 192 1645 592 1671
rect 650 1645 1050 1671
rect 1108 1645 1508 1671
rect 1566 1645 1966 1671
rect 2024 1645 2424 1671
rect 2482 1645 2882 1671
rect 2940 1645 3340 1671
rect 3398 1645 3798 1671
rect 3856 1645 4256 1671
rect 192 329 592 355
rect 650 329 1050 355
rect 1108 329 1508 355
rect 1566 329 1966 355
rect 2024 329 2424 355
rect 2482 329 2882 355
rect 2940 329 3340 355
rect 3398 329 3798 355
rect 3856 329 4256 355
rect 338 184 458 329
rect 794 184 914 329
rect 1250 184 1370 329
rect 1706 184 1826 329
rect 2162 184 2282 329
rect 2618 184 2738 329
rect 3074 184 3194 329
rect 3530 184 3650 329
rect 3986 184 4106 329
rect 98 164 4350 184
rect 98 104 268 164
rect 328 104 668 164
rect 728 104 1068 164
rect 1128 104 1468 164
rect 1528 104 1868 164
rect 1928 104 2268 164
rect 2328 104 2668 164
rect 2728 104 3068 164
rect 3128 104 3468 164
rect 3528 104 3868 164
rect 3928 104 4350 164
rect 98 84 4350 104
<< polycont >>
rect 268 104 328 164
rect 668 104 728 164
rect 1068 104 1128 164
rect 1468 104 1528 164
rect 1868 104 1928 164
rect 2268 104 2328 164
rect 2668 104 2728 164
rect 3068 104 3128 164
rect 3468 104 3528 164
rect 3868 104 3928 164
<< locali >>
rect 0 1850 268 1910
rect 328 1850 668 1910
rect 728 1850 1068 1910
rect 1128 1850 1468 1910
rect 1528 1850 1868 1910
rect 1928 1850 2268 1910
rect 2328 1850 2668 1910
rect 2728 1850 3068 1910
rect 3128 1850 3468 1910
rect 3528 1850 3868 1910
rect 3928 1850 4350 1910
rect 28 1760 88 1850
rect 28 1720 38 1760
rect 78 1720 88 1760
rect 158 1730 4350 1790
rect 28 1640 88 1720
rect 603 1649 637 1730
rect 1519 1649 1553 1730
rect 2435 1649 2469 1730
rect 3351 1649 3385 1730
rect 4267 1649 4301 1730
rect 146 1633 180 1649
rect 145 367 146 374
rect 603 1633 638 1649
rect 603 1626 604 1633
rect 145 351 180 367
rect 1062 1633 1096 1649
rect 604 351 638 367
rect 1061 367 1062 374
rect 1519 1633 1554 1649
rect 1519 1626 1520 1633
rect 1061 351 1096 367
rect 1978 1633 2012 1649
rect 1520 351 1554 367
rect 1977 367 1978 374
rect 2435 1633 2470 1649
rect 2435 1626 2436 1633
rect 1977 351 2012 367
rect 2894 1633 2928 1649
rect 2436 351 2470 367
rect 2893 367 2894 374
rect 3351 1633 3386 1649
rect 3351 1626 3352 1633
rect 2893 351 2928 367
rect 3810 1633 3844 1649
rect 3352 351 3386 367
rect 3809 367 3810 374
rect 4267 1633 4302 1649
rect 4267 1626 4268 1633
rect 3809 351 3844 367
rect 4268 351 4302 367
rect 145 270 179 351
rect 1061 270 1095 351
rect 1977 270 2011 351
rect 2893 270 2927 351
rect 3809 270 3843 351
rect 98 210 4350 270
rect 98 104 268 164
rect 328 104 668 164
rect 728 104 1068 164
rect 1128 104 1468 164
rect 1528 104 1868 164
rect 1928 104 2268 164
rect 2328 104 2668 164
rect 2728 104 3068 164
rect 3128 104 3468 164
rect 3528 104 3868 164
rect 3928 104 4350 164
rect 0 -30 268 30
rect 328 -30 668 30
rect 728 -30 1068 30
rect 1128 -30 1468 30
rect 1528 -30 1868 30
rect 1928 -30 2268 30
rect 2328 -30 2668 30
rect 2728 -30 3068 30
rect 3128 -30 3468 30
rect 3528 -30 3868 30
rect 3928 -30 4350 30
<< viali >>
rect 268 1850 328 1910
rect 668 1850 728 1910
rect 1068 1850 1128 1910
rect 1468 1850 1528 1910
rect 1868 1850 1928 1910
rect 2268 1850 2328 1910
rect 2668 1850 2728 1910
rect 3068 1850 3128 1910
rect 3468 1850 3528 1910
rect 3868 1850 3928 1910
rect 146 367 180 1633
rect 604 367 638 1633
rect 1062 367 1096 1633
rect 1520 367 1554 1633
rect 1978 367 2012 1633
rect 2436 367 2470 1633
rect 2894 367 2928 1633
rect 3352 367 3386 1633
rect 3810 367 3844 1633
rect 4268 367 4302 1633
rect 268 -30 328 30
rect 668 -30 728 30
rect 1068 -30 1128 30
rect 1468 -30 1528 30
rect 1868 -30 1928 30
rect 2268 -30 2328 30
rect 2668 -30 2728 30
rect 3068 -30 3128 30
rect 3468 -30 3528 30
rect 3868 -30 3928 30
<< metal1 >>
rect 0 1910 4350 1940
rect 0 1850 268 1910
rect 328 1850 668 1910
rect 728 1850 1068 1910
rect 1128 1850 1468 1910
rect 1528 1850 1868 1910
rect 1928 1850 2268 1910
rect 2328 1850 2668 1910
rect 2728 1850 3068 1910
rect 3128 1850 3468 1910
rect 3528 1850 3868 1910
rect 3928 1850 4350 1910
rect 0 1820 4350 1850
rect 140 1633 186 1645
rect 140 367 146 1633
rect 180 367 186 1633
rect 140 355 186 367
rect 598 1633 644 1645
rect 598 367 604 1633
rect 638 367 644 1633
rect 598 355 644 367
rect 1056 1633 1102 1645
rect 1056 367 1062 1633
rect 1096 367 1102 1633
rect 1056 355 1102 367
rect 1514 1633 1560 1645
rect 1514 367 1520 1633
rect 1554 367 1560 1633
rect 1514 355 1560 367
rect 1972 1633 2018 1645
rect 1972 367 1978 1633
rect 2012 367 2018 1633
rect 1972 355 2018 367
rect 2430 1633 2476 1645
rect 2430 367 2436 1633
rect 2470 367 2476 1633
rect 2430 355 2476 367
rect 2888 1633 2934 1645
rect 2888 367 2894 1633
rect 2928 367 2934 1633
rect 2888 355 2934 367
rect 3346 1633 3392 1645
rect 3346 367 3352 1633
rect 3386 367 3392 1633
rect 3346 355 3392 367
rect 3804 1633 3850 1645
rect 3804 367 3810 1633
rect 3844 367 3850 1633
rect 3804 355 3850 367
rect 4262 1633 4308 1645
rect 4262 367 4268 1633
rect 4302 367 4308 1633
rect 4262 355 4308 367
rect 0 30 4350 60
rect 0 -30 268 30
rect 328 -30 668 30
rect 728 -30 1068 30
rect 1128 -30 1468 30
rect 1528 -30 1868 30
rect 1928 -30 2268 30
rect 2328 -30 2668 30
rect 2728 -30 3068 30
rect 3128 -30 3468 30
rect 3528 -30 3868 30
rect 3928 -30 4350 30
rect 0 -60 4350 -30
<< labels >>
flabel nwell 0 1850 60 1910 1 FreeSans 800 0 0 0 VPWR
port 4 n power bidirectional
flabel metal1 0 -30 158 30 1 FreeSans 800 0 0 0 VGND
port 5 n ground bidirectional
flabel locali 4290 1730 4350 1790 1 FreeSans 800 0 0 0 SOURCE
port 2 n signal bidirectional
flabel locali 4290 210 4350 270 1 FreeSans 800 0 0 0 DRAIN
port 3 n signal bidirectional
flabel locali 4290 104 4350 164 1 FreeSans 800 0 0 0 GATE
port 1 n signal bidirectional
<< properties >>
string FIXED_BBOX 0 0 4350 1880
string LEFclass CORE
string LEFsite unitasc
<< end >>
