VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO sky130_asc_pfet_01v8_lvt_12
  CLASS CORE ;
  FOREIGN sky130_asc_pfet_01v8_lvt_12 ;
  ORIGIN 0.000 0.000 ;
  SIZE 29.815 BY 9.400 ;
  SITE unitasc ;
  PIN GATE
    DIRECTION INOUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 154.800003 ;
    PORT
      LAYER li1 ;
        RECT 1.090 0.520 29.210 0.820 ;
    END
  END GATE
  PIN SOURCE
    DIRECTION INOUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 11.223000 ;
    PORT
      LAYER li1 ;
        RECT 1.390 8.450 29.210 8.650 ;
        RECT 3.615 1.755 3.785 8.450 ;
        RECT 8.195 1.755 8.365 8.450 ;
        RECT 12.775 1.755 12.945 8.450 ;
        RECT 17.355 1.755 17.525 8.450 ;
        RECT 21.935 1.755 22.105 8.450 ;
        RECT 26.515 1.755 26.685 8.450 ;
      LAYER mcon ;
        RECT 3.615 1.835 3.785 8.165 ;
        RECT 8.195 1.835 8.365 8.165 ;
        RECT 12.775 1.835 12.945 8.165 ;
        RECT 17.355 1.835 17.525 8.165 ;
        RECT 21.935 1.835 22.105 8.165 ;
        RECT 26.515 1.835 26.685 8.165 ;
      LAYER met1 ;
        RECT 3.585 1.775 3.815 8.225 ;
        RECT 8.165 1.775 8.395 8.225 ;
        RECT 12.745 1.775 12.975 8.225 ;
        RECT 17.325 1.775 17.555 8.225 ;
        RECT 21.905 1.775 22.135 8.225 ;
        RECT 26.485 1.775 26.715 8.225 ;
    END
  END SOURCE
  PIN DRAIN
    DIRECTION INOUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 13.093500 ;
    PORT
      LAYER li1 ;
        RECT 1.325 1.350 1.495 8.245 ;
        RECT 5.905 1.350 6.075 8.245 ;
        RECT 10.485 1.350 10.655 8.245 ;
        RECT 15.065 1.350 15.235 8.245 ;
        RECT 19.645 1.350 19.815 8.245 ;
        RECT 24.225 1.350 24.395 8.245 ;
        RECT 28.805 1.350 28.975 8.245 ;
        RECT 1.090 1.050 29.210 1.350 ;
      LAYER mcon ;
        RECT 1.325 1.835 1.495 8.165 ;
        RECT 5.905 1.835 6.075 8.165 ;
        RECT 10.485 1.835 10.655 8.165 ;
        RECT 15.065 1.835 15.235 8.165 ;
        RECT 19.645 1.835 19.815 8.165 ;
        RECT 24.225 1.835 24.395 8.165 ;
        RECT 28.805 1.835 28.975 8.165 ;
      LAYER met1 ;
        RECT 1.295 1.775 1.525 8.225 ;
        RECT 5.875 1.775 6.105 8.225 ;
        RECT 10.455 1.775 10.685 8.225 ;
        RECT 15.035 1.775 15.265 8.225 ;
        RECT 19.615 1.775 19.845 8.225 ;
        RECT 24.195 1.775 24.425 8.225 ;
        RECT 28.775 1.775 29.005 8.225 ;
    END
  END DRAIN
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT 0.600 8.535 29.210 9.700 ;
        RECT 0.600 1.470 29.215 8.535 ;
        RECT 1.085 1.465 29.215 1.470 ;
      LAYER li1 ;
        RECT 0.600 9.250 29.210 9.550 ;
        RECT 0.740 8.200 1.040 9.250 ;
        RECT 5.980 8.850 6.780 9.250 ;
        RECT 12.480 8.850 13.280 9.250 ;
        RECT 18.980 8.850 19.780 9.250 ;
      LAYER mcon ;
        RECT 1.940 9.250 2.240 9.550 ;
        RECT 3.940 9.250 4.240 9.550 ;
        RECT 5.940 9.250 6.240 9.550 ;
        RECT 7.940 9.250 8.240 9.550 ;
        RECT 9.940 9.250 10.240 9.550 ;
        RECT 11.940 9.250 12.240 9.550 ;
        RECT 13.940 9.250 14.240 9.550 ;
        RECT 15.940 9.250 16.240 9.550 ;
        RECT 17.940 9.250 18.240 9.550 ;
        RECT 19.940 9.250 20.240 9.550 ;
        RECT 21.940 9.250 22.240 9.550 ;
        RECT 23.940 9.250 24.240 9.550 ;
        RECT 25.940 9.250 26.240 9.550 ;
        RECT 27.940 9.250 28.240 9.550 ;
      LAYER met1 ;
        RECT 0.600 9.100 29.210 9.700 ;
    END
  END VPWR
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER li1 ;
        RECT 0.600 -0.150 29.210 0.150 ;
      LAYER mcon ;
        RECT 1.940 -0.150 2.240 0.150 ;
        RECT 3.940 -0.150 4.240 0.150 ;
        RECT 5.940 -0.150 6.240 0.150 ;
        RECT 7.940 -0.150 8.240 0.150 ;
        RECT 9.940 -0.150 10.240 0.150 ;
        RECT 11.940 -0.150 12.240 0.150 ;
        RECT 13.940 -0.150 14.240 0.150 ;
        RECT 15.940 -0.150 16.240 0.150 ;
        RECT 17.940 -0.150 18.240 0.150 ;
        RECT 19.940 -0.150 20.240 0.150 ;
        RECT 21.940 -0.150 22.240 0.150 ;
        RECT 23.940 -0.150 24.240 0.150 ;
        RECT 25.940 -0.150 26.240 0.150 ;
        RECT 27.940 -0.150 28.240 0.150 ;
      LAYER met1 ;
        RECT 0.600 -0.300 29.210 0.300 ;
    END
  END VGND
END sky130_asc_pfet_01v8_lvt_12
END LIBRARY

