magic
tech sky130A
magscale 1 2
timestamp 1652753088
<< pwell >>
rect 90 1457 9470 1610
rect 90 423 243 1457
rect 1277 423 1583 1457
rect 2617 423 2923 1457
rect 3957 423 4263 1457
rect 5297 423 5603 1457
rect 6637 423 6943 1457
rect 7977 423 8283 1457
rect 9317 423 9470 1457
rect 90 270 9470 423
<< nbase >>
rect 243 423 1277 1457
rect 1583 423 2617 1457
rect 2923 423 3957 1457
rect 4263 423 5297 1457
rect 5603 423 6637 1457
rect 6943 423 7977 1457
rect 8283 423 9317 1457
<< pdiff >>
rect 420 1228 1100 1280
rect 420 1194 474 1228
rect 508 1194 564 1228
rect 598 1194 654 1228
rect 688 1194 744 1228
rect 778 1194 834 1228
rect 868 1194 924 1228
rect 958 1194 1014 1228
rect 1048 1194 1100 1228
rect 420 1138 1100 1194
rect 420 1104 474 1138
rect 508 1104 564 1138
rect 598 1104 654 1138
rect 688 1104 744 1138
rect 778 1104 834 1138
rect 868 1104 924 1138
rect 958 1104 1014 1138
rect 1048 1104 1100 1138
rect 420 1048 1100 1104
rect 420 1014 474 1048
rect 508 1014 564 1048
rect 598 1014 654 1048
rect 688 1014 744 1048
rect 778 1014 834 1048
rect 868 1014 924 1048
rect 958 1014 1014 1048
rect 1048 1014 1100 1048
rect 420 958 1100 1014
rect 420 924 474 958
rect 508 924 564 958
rect 598 924 654 958
rect 688 924 744 958
rect 778 924 834 958
rect 868 924 924 958
rect 958 924 1014 958
rect 1048 924 1100 958
rect 420 868 1100 924
rect 420 834 474 868
rect 508 834 564 868
rect 598 834 654 868
rect 688 834 744 868
rect 778 834 834 868
rect 868 834 924 868
rect 958 834 1014 868
rect 1048 834 1100 868
rect 420 778 1100 834
rect 420 744 474 778
rect 508 744 564 778
rect 598 744 654 778
rect 688 744 744 778
rect 778 744 834 778
rect 868 744 924 778
rect 958 744 1014 778
rect 1048 744 1100 778
rect 420 688 1100 744
rect 420 654 474 688
rect 508 654 564 688
rect 598 654 654 688
rect 688 654 744 688
rect 778 654 834 688
rect 868 654 924 688
rect 958 654 1014 688
rect 1048 654 1100 688
rect 420 600 1100 654
rect 1760 1228 2440 1280
rect 1760 1194 1814 1228
rect 1848 1194 1904 1228
rect 1938 1194 1994 1228
rect 2028 1194 2084 1228
rect 2118 1194 2174 1228
rect 2208 1194 2264 1228
rect 2298 1194 2354 1228
rect 2388 1194 2440 1228
rect 1760 1138 2440 1194
rect 1760 1104 1814 1138
rect 1848 1104 1904 1138
rect 1938 1104 1994 1138
rect 2028 1104 2084 1138
rect 2118 1104 2174 1138
rect 2208 1104 2264 1138
rect 2298 1104 2354 1138
rect 2388 1104 2440 1138
rect 1760 1048 2440 1104
rect 1760 1014 1814 1048
rect 1848 1014 1904 1048
rect 1938 1014 1994 1048
rect 2028 1014 2084 1048
rect 2118 1014 2174 1048
rect 2208 1014 2264 1048
rect 2298 1014 2354 1048
rect 2388 1014 2440 1048
rect 1760 958 2440 1014
rect 1760 924 1814 958
rect 1848 924 1904 958
rect 1938 924 1994 958
rect 2028 924 2084 958
rect 2118 924 2174 958
rect 2208 924 2264 958
rect 2298 924 2354 958
rect 2388 924 2440 958
rect 1760 868 2440 924
rect 1760 834 1814 868
rect 1848 834 1904 868
rect 1938 834 1994 868
rect 2028 834 2084 868
rect 2118 834 2174 868
rect 2208 834 2264 868
rect 2298 834 2354 868
rect 2388 834 2440 868
rect 1760 778 2440 834
rect 1760 744 1814 778
rect 1848 744 1904 778
rect 1938 744 1994 778
rect 2028 744 2084 778
rect 2118 744 2174 778
rect 2208 744 2264 778
rect 2298 744 2354 778
rect 2388 744 2440 778
rect 1760 688 2440 744
rect 1760 654 1814 688
rect 1848 654 1904 688
rect 1938 654 1994 688
rect 2028 654 2084 688
rect 2118 654 2174 688
rect 2208 654 2264 688
rect 2298 654 2354 688
rect 2388 654 2440 688
rect 1760 600 2440 654
rect 3100 1228 3780 1280
rect 3100 1194 3154 1228
rect 3188 1194 3244 1228
rect 3278 1194 3334 1228
rect 3368 1194 3424 1228
rect 3458 1194 3514 1228
rect 3548 1194 3604 1228
rect 3638 1194 3694 1228
rect 3728 1194 3780 1228
rect 3100 1138 3780 1194
rect 3100 1104 3154 1138
rect 3188 1104 3244 1138
rect 3278 1104 3334 1138
rect 3368 1104 3424 1138
rect 3458 1104 3514 1138
rect 3548 1104 3604 1138
rect 3638 1104 3694 1138
rect 3728 1104 3780 1138
rect 3100 1048 3780 1104
rect 3100 1014 3154 1048
rect 3188 1014 3244 1048
rect 3278 1014 3334 1048
rect 3368 1014 3424 1048
rect 3458 1014 3514 1048
rect 3548 1014 3604 1048
rect 3638 1014 3694 1048
rect 3728 1014 3780 1048
rect 3100 958 3780 1014
rect 3100 924 3154 958
rect 3188 924 3244 958
rect 3278 924 3334 958
rect 3368 924 3424 958
rect 3458 924 3514 958
rect 3548 924 3604 958
rect 3638 924 3694 958
rect 3728 924 3780 958
rect 3100 868 3780 924
rect 3100 834 3154 868
rect 3188 834 3244 868
rect 3278 834 3334 868
rect 3368 834 3424 868
rect 3458 834 3514 868
rect 3548 834 3604 868
rect 3638 834 3694 868
rect 3728 834 3780 868
rect 3100 778 3780 834
rect 3100 744 3154 778
rect 3188 744 3244 778
rect 3278 744 3334 778
rect 3368 744 3424 778
rect 3458 744 3514 778
rect 3548 744 3604 778
rect 3638 744 3694 778
rect 3728 744 3780 778
rect 3100 688 3780 744
rect 3100 654 3154 688
rect 3188 654 3244 688
rect 3278 654 3334 688
rect 3368 654 3424 688
rect 3458 654 3514 688
rect 3548 654 3604 688
rect 3638 654 3694 688
rect 3728 654 3780 688
rect 3100 600 3780 654
rect 4440 1228 5120 1280
rect 4440 1194 4494 1228
rect 4528 1194 4584 1228
rect 4618 1194 4674 1228
rect 4708 1194 4764 1228
rect 4798 1194 4854 1228
rect 4888 1194 4944 1228
rect 4978 1194 5034 1228
rect 5068 1194 5120 1228
rect 4440 1138 5120 1194
rect 4440 1104 4494 1138
rect 4528 1104 4584 1138
rect 4618 1104 4674 1138
rect 4708 1104 4764 1138
rect 4798 1104 4854 1138
rect 4888 1104 4944 1138
rect 4978 1104 5034 1138
rect 5068 1104 5120 1138
rect 4440 1048 5120 1104
rect 4440 1014 4494 1048
rect 4528 1014 4584 1048
rect 4618 1014 4674 1048
rect 4708 1014 4764 1048
rect 4798 1014 4854 1048
rect 4888 1014 4944 1048
rect 4978 1014 5034 1048
rect 5068 1014 5120 1048
rect 4440 958 5120 1014
rect 4440 924 4494 958
rect 4528 924 4584 958
rect 4618 924 4674 958
rect 4708 924 4764 958
rect 4798 924 4854 958
rect 4888 924 4944 958
rect 4978 924 5034 958
rect 5068 924 5120 958
rect 4440 868 5120 924
rect 4440 834 4494 868
rect 4528 834 4584 868
rect 4618 834 4674 868
rect 4708 834 4764 868
rect 4798 834 4854 868
rect 4888 834 4944 868
rect 4978 834 5034 868
rect 5068 834 5120 868
rect 4440 778 5120 834
rect 4440 744 4494 778
rect 4528 744 4584 778
rect 4618 744 4674 778
rect 4708 744 4764 778
rect 4798 744 4854 778
rect 4888 744 4944 778
rect 4978 744 5034 778
rect 5068 744 5120 778
rect 4440 688 5120 744
rect 4440 654 4494 688
rect 4528 654 4584 688
rect 4618 654 4674 688
rect 4708 654 4764 688
rect 4798 654 4854 688
rect 4888 654 4944 688
rect 4978 654 5034 688
rect 5068 654 5120 688
rect 4440 600 5120 654
rect 5780 1228 6460 1280
rect 5780 1194 5834 1228
rect 5868 1194 5924 1228
rect 5958 1194 6014 1228
rect 6048 1194 6104 1228
rect 6138 1194 6194 1228
rect 6228 1194 6284 1228
rect 6318 1194 6374 1228
rect 6408 1194 6460 1228
rect 5780 1138 6460 1194
rect 5780 1104 5834 1138
rect 5868 1104 5924 1138
rect 5958 1104 6014 1138
rect 6048 1104 6104 1138
rect 6138 1104 6194 1138
rect 6228 1104 6284 1138
rect 6318 1104 6374 1138
rect 6408 1104 6460 1138
rect 5780 1048 6460 1104
rect 5780 1014 5834 1048
rect 5868 1014 5924 1048
rect 5958 1014 6014 1048
rect 6048 1014 6104 1048
rect 6138 1014 6194 1048
rect 6228 1014 6284 1048
rect 6318 1014 6374 1048
rect 6408 1014 6460 1048
rect 5780 958 6460 1014
rect 5780 924 5834 958
rect 5868 924 5924 958
rect 5958 924 6014 958
rect 6048 924 6104 958
rect 6138 924 6194 958
rect 6228 924 6284 958
rect 6318 924 6374 958
rect 6408 924 6460 958
rect 5780 868 6460 924
rect 5780 834 5834 868
rect 5868 834 5924 868
rect 5958 834 6014 868
rect 6048 834 6104 868
rect 6138 834 6194 868
rect 6228 834 6284 868
rect 6318 834 6374 868
rect 6408 834 6460 868
rect 5780 778 6460 834
rect 5780 744 5834 778
rect 5868 744 5924 778
rect 5958 744 6014 778
rect 6048 744 6104 778
rect 6138 744 6194 778
rect 6228 744 6284 778
rect 6318 744 6374 778
rect 6408 744 6460 778
rect 5780 688 6460 744
rect 5780 654 5834 688
rect 5868 654 5924 688
rect 5958 654 6014 688
rect 6048 654 6104 688
rect 6138 654 6194 688
rect 6228 654 6284 688
rect 6318 654 6374 688
rect 6408 654 6460 688
rect 5780 600 6460 654
rect 7120 1228 7800 1280
rect 7120 1194 7174 1228
rect 7208 1194 7264 1228
rect 7298 1194 7354 1228
rect 7388 1194 7444 1228
rect 7478 1194 7534 1228
rect 7568 1194 7624 1228
rect 7658 1194 7714 1228
rect 7748 1194 7800 1228
rect 7120 1138 7800 1194
rect 7120 1104 7174 1138
rect 7208 1104 7264 1138
rect 7298 1104 7354 1138
rect 7388 1104 7444 1138
rect 7478 1104 7534 1138
rect 7568 1104 7624 1138
rect 7658 1104 7714 1138
rect 7748 1104 7800 1138
rect 7120 1048 7800 1104
rect 7120 1014 7174 1048
rect 7208 1014 7264 1048
rect 7298 1014 7354 1048
rect 7388 1014 7444 1048
rect 7478 1014 7534 1048
rect 7568 1014 7624 1048
rect 7658 1014 7714 1048
rect 7748 1014 7800 1048
rect 7120 958 7800 1014
rect 7120 924 7174 958
rect 7208 924 7264 958
rect 7298 924 7354 958
rect 7388 924 7444 958
rect 7478 924 7534 958
rect 7568 924 7624 958
rect 7658 924 7714 958
rect 7748 924 7800 958
rect 7120 868 7800 924
rect 7120 834 7174 868
rect 7208 834 7264 868
rect 7298 834 7354 868
rect 7388 834 7444 868
rect 7478 834 7534 868
rect 7568 834 7624 868
rect 7658 834 7714 868
rect 7748 834 7800 868
rect 7120 778 7800 834
rect 7120 744 7174 778
rect 7208 744 7264 778
rect 7298 744 7354 778
rect 7388 744 7444 778
rect 7478 744 7534 778
rect 7568 744 7624 778
rect 7658 744 7714 778
rect 7748 744 7800 778
rect 7120 688 7800 744
rect 7120 654 7174 688
rect 7208 654 7264 688
rect 7298 654 7354 688
rect 7388 654 7444 688
rect 7478 654 7534 688
rect 7568 654 7624 688
rect 7658 654 7714 688
rect 7748 654 7800 688
rect 7120 600 7800 654
rect 8460 1228 9140 1280
rect 8460 1194 8514 1228
rect 8548 1194 8604 1228
rect 8638 1194 8694 1228
rect 8728 1194 8784 1228
rect 8818 1194 8874 1228
rect 8908 1194 8964 1228
rect 8998 1194 9054 1228
rect 9088 1194 9140 1228
rect 8460 1138 9140 1194
rect 8460 1104 8514 1138
rect 8548 1104 8604 1138
rect 8638 1104 8694 1138
rect 8728 1104 8784 1138
rect 8818 1104 8874 1138
rect 8908 1104 8964 1138
rect 8998 1104 9054 1138
rect 9088 1104 9140 1138
rect 8460 1048 9140 1104
rect 8460 1014 8514 1048
rect 8548 1014 8604 1048
rect 8638 1014 8694 1048
rect 8728 1014 8784 1048
rect 8818 1014 8874 1048
rect 8908 1014 8964 1048
rect 8998 1014 9054 1048
rect 9088 1014 9140 1048
rect 8460 958 9140 1014
rect 8460 924 8514 958
rect 8548 924 8604 958
rect 8638 924 8694 958
rect 8728 924 8784 958
rect 8818 924 8874 958
rect 8908 924 8964 958
rect 8998 924 9054 958
rect 9088 924 9140 958
rect 8460 868 9140 924
rect 8460 834 8514 868
rect 8548 834 8604 868
rect 8638 834 8694 868
rect 8728 834 8784 868
rect 8818 834 8874 868
rect 8908 834 8964 868
rect 8998 834 9054 868
rect 9088 834 9140 868
rect 8460 778 9140 834
rect 8460 744 8514 778
rect 8548 744 8604 778
rect 8638 744 8694 778
rect 8728 744 8784 778
rect 8818 744 8874 778
rect 8908 744 8964 778
rect 8998 744 9054 778
rect 9088 744 9140 778
rect 8460 688 9140 744
rect 8460 654 8514 688
rect 8548 654 8604 688
rect 8638 654 8694 688
rect 8728 654 8784 688
rect 8818 654 8874 688
rect 8908 654 8964 688
rect 8998 654 9054 688
rect 9088 654 9140 688
rect 8460 600 9140 654
<< pdiffc >>
rect 474 1194 508 1228
rect 564 1194 598 1228
rect 654 1194 688 1228
rect 744 1194 778 1228
rect 834 1194 868 1228
rect 924 1194 958 1228
rect 1014 1194 1048 1228
rect 474 1104 508 1138
rect 564 1104 598 1138
rect 654 1104 688 1138
rect 744 1104 778 1138
rect 834 1104 868 1138
rect 924 1104 958 1138
rect 1014 1104 1048 1138
rect 474 1014 508 1048
rect 564 1014 598 1048
rect 654 1014 688 1048
rect 744 1014 778 1048
rect 834 1014 868 1048
rect 924 1014 958 1048
rect 1014 1014 1048 1048
rect 474 924 508 958
rect 564 924 598 958
rect 654 924 688 958
rect 744 924 778 958
rect 834 924 868 958
rect 924 924 958 958
rect 1014 924 1048 958
rect 474 834 508 868
rect 564 834 598 868
rect 654 834 688 868
rect 744 834 778 868
rect 834 834 868 868
rect 924 834 958 868
rect 1014 834 1048 868
rect 474 744 508 778
rect 564 744 598 778
rect 654 744 688 778
rect 744 744 778 778
rect 834 744 868 778
rect 924 744 958 778
rect 1014 744 1048 778
rect 474 654 508 688
rect 564 654 598 688
rect 654 654 688 688
rect 744 654 778 688
rect 834 654 868 688
rect 924 654 958 688
rect 1014 654 1048 688
rect 1814 1194 1848 1228
rect 1904 1194 1938 1228
rect 1994 1194 2028 1228
rect 2084 1194 2118 1228
rect 2174 1194 2208 1228
rect 2264 1194 2298 1228
rect 2354 1194 2388 1228
rect 1814 1104 1848 1138
rect 1904 1104 1938 1138
rect 1994 1104 2028 1138
rect 2084 1104 2118 1138
rect 2174 1104 2208 1138
rect 2264 1104 2298 1138
rect 2354 1104 2388 1138
rect 1814 1014 1848 1048
rect 1904 1014 1938 1048
rect 1994 1014 2028 1048
rect 2084 1014 2118 1048
rect 2174 1014 2208 1048
rect 2264 1014 2298 1048
rect 2354 1014 2388 1048
rect 1814 924 1848 958
rect 1904 924 1938 958
rect 1994 924 2028 958
rect 2084 924 2118 958
rect 2174 924 2208 958
rect 2264 924 2298 958
rect 2354 924 2388 958
rect 1814 834 1848 868
rect 1904 834 1938 868
rect 1994 834 2028 868
rect 2084 834 2118 868
rect 2174 834 2208 868
rect 2264 834 2298 868
rect 2354 834 2388 868
rect 1814 744 1848 778
rect 1904 744 1938 778
rect 1994 744 2028 778
rect 2084 744 2118 778
rect 2174 744 2208 778
rect 2264 744 2298 778
rect 2354 744 2388 778
rect 1814 654 1848 688
rect 1904 654 1938 688
rect 1994 654 2028 688
rect 2084 654 2118 688
rect 2174 654 2208 688
rect 2264 654 2298 688
rect 2354 654 2388 688
rect 3154 1194 3188 1228
rect 3244 1194 3278 1228
rect 3334 1194 3368 1228
rect 3424 1194 3458 1228
rect 3514 1194 3548 1228
rect 3604 1194 3638 1228
rect 3694 1194 3728 1228
rect 3154 1104 3188 1138
rect 3244 1104 3278 1138
rect 3334 1104 3368 1138
rect 3424 1104 3458 1138
rect 3514 1104 3548 1138
rect 3604 1104 3638 1138
rect 3694 1104 3728 1138
rect 3154 1014 3188 1048
rect 3244 1014 3278 1048
rect 3334 1014 3368 1048
rect 3424 1014 3458 1048
rect 3514 1014 3548 1048
rect 3604 1014 3638 1048
rect 3694 1014 3728 1048
rect 3154 924 3188 958
rect 3244 924 3278 958
rect 3334 924 3368 958
rect 3424 924 3458 958
rect 3514 924 3548 958
rect 3604 924 3638 958
rect 3694 924 3728 958
rect 3154 834 3188 868
rect 3244 834 3278 868
rect 3334 834 3368 868
rect 3424 834 3458 868
rect 3514 834 3548 868
rect 3604 834 3638 868
rect 3694 834 3728 868
rect 3154 744 3188 778
rect 3244 744 3278 778
rect 3334 744 3368 778
rect 3424 744 3458 778
rect 3514 744 3548 778
rect 3604 744 3638 778
rect 3694 744 3728 778
rect 3154 654 3188 688
rect 3244 654 3278 688
rect 3334 654 3368 688
rect 3424 654 3458 688
rect 3514 654 3548 688
rect 3604 654 3638 688
rect 3694 654 3728 688
rect 4494 1194 4528 1228
rect 4584 1194 4618 1228
rect 4674 1194 4708 1228
rect 4764 1194 4798 1228
rect 4854 1194 4888 1228
rect 4944 1194 4978 1228
rect 5034 1194 5068 1228
rect 4494 1104 4528 1138
rect 4584 1104 4618 1138
rect 4674 1104 4708 1138
rect 4764 1104 4798 1138
rect 4854 1104 4888 1138
rect 4944 1104 4978 1138
rect 5034 1104 5068 1138
rect 4494 1014 4528 1048
rect 4584 1014 4618 1048
rect 4674 1014 4708 1048
rect 4764 1014 4798 1048
rect 4854 1014 4888 1048
rect 4944 1014 4978 1048
rect 5034 1014 5068 1048
rect 4494 924 4528 958
rect 4584 924 4618 958
rect 4674 924 4708 958
rect 4764 924 4798 958
rect 4854 924 4888 958
rect 4944 924 4978 958
rect 5034 924 5068 958
rect 4494 834 4528 868
rect 4584 834 4618 868
rect 4674 834 4708 868
rect 4764 834 4798 868
rect 4854 834 4888 868
rect 4944 834 4978 868
rect 5034 834 5068 868
rect 4494 744 4528 778
rect 4584 744 4618 778
rect 4674 744 4708 778
rect 4764 744 4798 778
rect 4854 744 4888 778
rect 4944 744 4978 778
rect 5034 744 5068 778
rect 4494 654 4528 688
rect 4584 654 4618 688
rect 4674 654 4708 688
rect 4764 654 4798 688
rect 4854 654 4888 688
rect 4944 654 4978 688
rect 5034 654 5068 688
rect 5834 1194 5868 1228
rect 5924 1194 5958 1228
rect 6014 1194 6048 1228
rect 6104 1194 6138 1228
rect 6194 1194 6228 1228
rect 6284 1194 6318 1228
rect 6374 1194 6408 1228
rect 5834 1104 5868 1138
rect 5924 1104 5958 1138
rect 6014 1104 6048 1138
rect 6104 1104 6138 1138
rect 6194 1104 6228 1138
rect 6284 1104 6318 1138
rect 6374 1104 6408 1138
rect 5834 1014 5868 1048
rect 5924 1014 5958 1048
rect 6014 1014 6048 1048
rect 6104 1014 6138 1048
rect 6194 1014 6228 1048
rect 6284 1014 6318 1048
rect 6374 1014 6408 1048
rect 5834 924 5868 958
rect 5924 924 5958 958
rect 6014 924 6048 958
rect 6104 924 6138 958
rect 6194 924 6228 958
rect 6284 924 6318 958
rect 6374 924 6408 958
rect 5834 834 5868 868
rect 5924 834 5958 868
rect 6014 834 6048 868
rect 6104 834 6138 868
rect 6194 834 6228 868
rect 6284 834 6318 868
rect 6374 834 6408 868
rect 5834 744 5868 778
rect 5924 744 5958 778
rect 6014 744 6048 778
rect 6104 744 6138 778
rect 6194 744 6228 778
rect 6284 744 6318 778
rect 6374 744 6408 778
rect 5834 654 5868 688
rect 5924 654 5958 688
rect 6014 654 6048 688
rect 6104 654 6138 688
rect 6194 654 6228 688
rect 6284 654 6318 688
rect 6374 654 6408 688
rect 7174 1194 7208 1228
rect 7264 1194 7298 1228
rect 7354 1194 7388 1228
rect 7444 1194 7478 1228
rect 7534 1194 7568 1228
rect 7624 1194 7658 1228
rect 7714 1194 7748 1228
rect 7174 1104 7208 1138
rect 7264 1104 7298 1138
rect 7354 1104 7388 1138
rect 7444 1104 7478 1138
rect 7534 1104 7568 1138
rect 7624 1104 7658 1138
rect 7714 1104 7748 1138
rect 7174 1014 7208 1048
rect 7264 1014 7298 1048
rect 7354 1014 7388 1048
rect 7444 1014 7478 1048
rect 7534 1014 7568 1048
rect 7624 1014 7658 1048
rect 7714 1014 7748 1048
rect 7174 924 7208 958
rect 7264 924 7298 958
rect 7354 924 7388 958
rect 7444 924 7478 958
rect 7534 924 7568 958
rect 7624 924 7658 958
rect 7714 924 7748 958
rect 7174 834 7208 868
rect 7264 834 7298 868
rect 7354 834 7388 868
rect 7444 834 7478 868
rect 7534 834 7568 868
rect 7624 834 7658 868
rect 7714 834 7748 868
rect 7174 744 7208 778
rect 7264 744 7298 778
rect 7354 744 7388 778
rect 7444 744 7478 778
rect 7534 744 7568 778
rect 7624 744 7658 778
rect 7714 744 7748 778
rect 7174 654 7208 688
rect 7264 654 7298 688
rect 7354 654 7388 688
rect 7444 654 7478 688
rect 7534 654 7568 688
rect 7624 654 7658 688
rect 7714 654 7748 688
rect 8514 1194 8548 1228
rect 8604 1194 8638 1228
rect 8694 1194 8728 1228
rect 8784 1194 8818 1228
rect 8874 1194 8908 1228
rect 8964 1194 8998 1228
rect 9054 1194 9088 1228
rect 8514 1104 8548 1138
rect 8604 1104 8638 1138
rect 8694 1104 8728 1138
rect 8784 1104 8818 1138
rect 8874 1104 8908 1138
rect 8964 1104 8998 1138
rect 9054 1104 9088 1138
rect 8514 1014 8548 1048
rect 8604 1014 8638 1048
rect 8694 1014 8728 1048
rect 8784 1014 8818 1048
rect 8874 1014 8908 1048
rect 8964 1014 8998 1048
rect 9054 1014 9088 1048
rect 8514 924 8548 958
rect 8604 924 8638 958
rect 8694 924 8728 958
rect 8784 924 8818 958
rect 8874 924 8908 958
rect 8964 924 8998 958
rect 9054 924 9088 958
rect 8514 834 8548 868
rect 8604 834 8638 868
rect 8694 834 8728 868
rect 8784 834 8818 868
rect 8874 834 8908 868
rect 8964 834 8998 868
rect 9054 834 9088 868
rect 8514 744 8548 778
rect 8604 744 8638 778
rect 8694 744 8728 778
rect 8784 744 8818 778
rect 8874 744 8908 778
rect 8964 744 8998 778
rect 9054 744 9088 778
rect 8514 654 8548 688
rect 8604 654 8638 688
rect 8694 654 8728 688
rect 8784 654 8818 688
rect 8874 654 8908 688
rect 8964 654 8998 688
rect 9054 654 9088 688
<< psubdiff >>
rect 116 1549 9444 1584
rect 116 1526 246 1549
rect 116 1492 150 1526
rect 184 1515 246 1526
rect 280 1515 336 1549
rect 370 1515 426 1549
rect 460 1515 516 1549
rect 550 1515 606 1549
rect 640 1515 696 1549
rect 730 1515 786 1549
rect 820 1515 876 1549
rect 910 1515 966 1549
rect 1000 1515 1056 1549
rect 1090 1515 1146 1549
rect 1180 1515 1236 1549
rect 1270 1526 1586 1549
rect 1270 1515 1337 1526
rect 184 1492 1337 1515
rect 1371 1492 1490 1526
rect 1524 1515 1586 1526
rect 1620 1515 1676 1549
rect 1710 1515 1766 1549
rect 1800 1515 1856 1549
rect 1890 1515 1946 1549
rect 1980 1515 2036 1549
rect 2070 1515 2126 1549
rect 2160 1515 2216 1549
rect 2250 1515 2306 1549
rect 2340 1515 2396 1549
rect 2430 1515 2486 1549
rect 2520 1515 2576 1549
rect 2610 1526 2926 1549
rect 2610 1515 2677 1526
rect 1524 1492 2677 1515
rect 2711 1492 2830 1526
rect 2864 1515 2926 1526
rect 2960 1515 3016 1549
rect 3050 1515 3106 1549
rect 3140 1515 3196 1549
rect 3230 1515 3286 1549
rect 3320 1515 3376 1549
rect 3410 1515 3466 1549
rect 3500 1515 3556 1549
rect 3590 1515 3646 1549
rect 3680 1515 3736 1549
rect 3770 1515 3826 1549
rect 3860 1515 3916 1549
rect 3950 1526 4266 1549
rect 3950 1515 4017 1526
rect 2864 1492 4017 1515
rect 4051 1492 4170 1526
rect 4204 1515 4266 1526
rect 4300 1515 4356 1549
rect 4390 1515 4446 1549
rect 4480 1515 4536 1549
rect 4570 1515 4626 1549
rect 4660 1515 4716 1549
rect 4750 1515 4806 1549
rect 4840 1515 4896 1549
rect 4930 1515 4986 1549
rect 5020 1515 5076 1549
rect 5110 1515 5166 1549
rect 5200 1515 5256 1549
rect 5290 1526 5606 1549
rect 5290 1515 5357 1526
rect 4204 1492 5357 1515
rect 5391 1492 5510 1526
rect 5544 1515 5606 1526
rect 5640 1515 5696 1549
rect 5730 1515 5786 1549
rect 5820 1515 5876 1549
rect 5910 1515 5966 1549
rect 6000 1515 6056 1549
rect 6090 1515 6146 1549
rect 6180 1515 6236 1549
rect 6270 1515 6326 1549
rect 6360 1515 6416 1549
rect 6450 1515 6506 1549
rect 6540 1515 6596 1549
rect 6630 1526 6946 1549
rect 6630 1515 6697 1526
rect 5544 1492 6697 1515
rect 6731 1492 6850 1526
rect 6884 1515 6946 1526
rect 6980 1515 7036 1549
rect 7070 1515 7126 1549
rect 7160 1515 7216 1549
rect 7250 1515 7306 1549
rect 7340 1515 7396 1549
rect 7430 1515 7486 1549
rect 7520 1515 7576 1549
rect 7610 1515 7666 1549
rect 7700 1515 7756 1549
rect 7790 1515 7846 1549
rect 7880 1515 7936 1549
rect 7970 1526 8286 1549
rect 7970 1515 8037 1526
rect 6884 1492 8037 1515
rect 8071 1492 8190 1526
rect 8224 1515 8286 1526
rect 8320 1515 8376 1549
rect 8410 1515 8466 1549
rect 8500 1515 8556 1549
rect 8590 1515 8646 1549
rect 8680 1515 8736 1549
rect 8770 1515 8826 1549
rect 8860 1515 8916 1549
rect 8950 1515 9006 1549
rect 9040 1515 9096 1549
rect 9130 1515 9186 1549
rect 9220 1515 9276 1549
rect 9310 1526 9444 1549
rect 9310 1515 9377 1526
rect 8224 1492 9377 1515
rect 9411 1492 9444 1526
rect 116 1483 9444 1492
rect 116 1436 217 1483
rect 116 1402 150 1436
rect 184 1402 217 1436
rect 1303 1436 1557 1483
rect 116 1346 217 1402
rect 116 1312 150 1346
rect 184 1312 217 1346
rect 116 1256 217 1312
rect 116 1222 150 1256
rect 184 1222 217 1256
rect 116 1166 217 1222
rect 116 1132 150 1166
rect 184 1132 217 1166
rect 116 1076 217 1132
rect 116 1042 150 1076
rect 184 1042 217 1076
rect 116 986 217 1042
rect 116 952 150 986
rect 184 952 217 986
rect 116 896 217 952
rect 116 862 150 896
rect 184 862 217 896
rect 116 806 217 862
rect 116 772 150 806
rect 184 772 217 806
rect 116 716 217 772
rect 116 682 150 716
rect 184 682 217 716
rect 116 626 217 682
rect 116 592 150 626
rect 184 592 217 626
rect 116 536 217 592
rect 116 502 150 536
rect 184 502 217 536
rect 116 446 217 502
rect 1303 1402 1337 1436
rect 1371 1402 1490 1436
rect 1524 1402 1557 1436
rect 2643 1436 2897 1483
rect 1303 1346 1557 1402
rect 1303 1312 1337 1346
rect 1371 1312 1490 1346
rect 1524 1312 1557 1346
rect 1303 1256 1557 1312
rect 1303 1222 1337 1256
rect 1371 1222 1490 1256
rect 1524 1222 1557 1256
rect 1303 1166 1557 1222
rect 1303 1132 1337 1166
rect 1371 1132 1490 1166
rect 1524 1132 1557 1166
rect 1303 1076 1557 1132
rect 1303 1042 1337 1076
rect 1371 1042 1490 1076
rect 1524 1042 1557 1076
rect 1303 986 1557 1042
rect 1303 952 1337 986
rect 1371 952 1490 986
rect 1524 952 1557 986
rect 1303 896 1557 952
rect 1303 862 1337 896
rect 1371 862 1490 896
rect 1524 862 1557 896
rect 1303 806 1557 862
rect 1303 772 1337 806
rect 1371 772 1490 806
rect 1524 772 1557 806
rect 1303 716 1557 772
rect 1303 682 1337 716
rect 1371 682 1490 716
rect 1524 682 1557 716
rect 1303 626 1557 682
rect 1303 592 1337 626
rect 1371 592 1490 626
rect 1524 592 1557 626
rect 1303 536 1557 592
rect 1303 502 1337 536
rect 1371 502 1490 536
rect 1524 502 1557 536
rect 116 412 150 446
rect 184 412 217 446
rect 116 397 217 412
rect 1303 446 1557 502
rect 2643 1402 2677 1436
rect 2711 1402 2830 1436
rect 2864 1402 2897 1436
rect 3983 1436 4237 1483
rect 2643 1346 2897 1402
rect 2643 1312 2677 1346
rect 2711 1312 2830 1346
rect 2864 1312 2897 1346
rect 2643 1256 2897 1312
rect 2643 1222 2677 1256
rect 2711 1222 2830 1256
rect 2864 1222 2897 1256
rect 2643 1166 2897 1222
rect 2643 1132 2677 1166
rect 2711 1132 2830 1166
rect 2864 1132 2897 1166
rect 2643 1076 2897 1132
rect 2643 1042 2677 1076
rect 2711 1042 2830 1076
rect 2864 1042 2897 1076
rect 2643 986 2897 1042
rect 2643 952 2677 986
rect 2711 952 2830 986
rect 2864 952 2897 986
rect 2643 896 2897 952
rect 2643 862 2677 896
rect 2711 862 2830 896
rect 2864 862 2897 896
rect 2643 806 2897 862
rect 2643 772 2677 806
rect 2711 772 2830 806
rect 2864 772 2897 806
rect 2643 716 2897 772
rect 2643 682 2677 716
rect 2711 682 2830 716
rect 2864 682 2897 716
rect 2643 626 2897 682
rect 2643 592 2677 626
rect 2711 592 2830 626
rect 2864 592 2897 626
rect 2643 536 2897 592
rect 2643 502 2677 536
rect 2711 502 2830 536
rect 2864 502 2897 536
rect 1303 412 1337 446
rect 1371 412 1490 446
rect 1524 412 1557 446
rect 1303 397 1557 412
rect 2643 446 2897 502
rect 3983 1402 4017 1436
rect 4051 1402 4170 1436
rect 4204 1402 4237 1436
rect 5323 1436 5577 1483
rect 3983 1346 4237 1402
rect 3983 1312 4017 1346
rect 4051 1312 4170 1346
rect 4204 1312 4237 1346
rect 3983 1256 4237 1312
rect 3983 1222 4017 1256
rect 4051 1222 4170 1256
rect 4204 1222 4237 1256
rect 3983 1166 4237 1222
rect 3983 1132 4017 1166
rect 4051 1132 4170 1166
rect 4204 1132 4237 1166
rect 3983 1076 4237 1132
rect 3983 1042 4017 1076
rect 4051 1042 4170 1076
rect 4204 1042 4237 1076
rect 3983 986 4237 1042
rect 3983 952 4017 986
rect 4051 952 4170 986
rect 4204 952 4237 986
rect 3983 896 4237 952
rect 3983 862 4017 896
rect 4051 862 4170 896
rect 4204 862 4237 896
rect 3983 806 4237 862
rect 3983 772 4017 806
rect 4051 772 4170 806
rect 4204 772 4237 806
rect 3983 716 4237 772
rect 3983 682 4017 716
rect 4051 682 4170 716
rect 4204 682 4237 716
rect 3983 626 4237 682
rect 3983 592 4017 626
rect 4051 592 4170 626
rect 4204 592 4237 626
rect 3983 536 4237 592
rect 3983 502 4017 536
rect 4051 502 4170 536
rect 4204 502 4237 536
rect 2643 412 2677 446
rect 2711 412 2830 446
rect 2864 412 2897 446
rect 2643 397 2897 412
rect 3983 446 4237 502
rect 5323 1402 5357 1436
rect 5391 1402 5510 1436
rect 5544 1402 5577 1436
rect 6663 1436 6917 1483
rect 5323 1346 5577 1402
rect 5323 1312 5357 1346
rect 5391 1312 5510 1346
rect 5544 1312 5577 1346
rect 5323 1256 5577 1312
rect 5323 1222 5357 1256
rect 5391 1222 5510 1256
rect 5544 1222 5577 1256
rect 5323 1166 5577 1222
rect 5323 1132 5357 1166
rect 5391 1132 5510 1166
rect 5544 1132 5577 1166
rect 5323 1076 5577 1132
rect 5323 1042 5357 1076
rect 5391 1042 5510 1076
rect 5544 1042 5577 1076
rect 5323 986 5577 1042
rect 5323 952 5357 986
rect 5391 952 5510 986
rect 5544 952 5577 986
rect 5323 896 5577 952
rect 5323 862 5357 896
rect 5391 862 5510 896
rect 5544 862 5577 896
rect 5323 806 5577 862
rect 5323 772 5357 806
rect 5391 772 5510 806
rect 5544 772 5577 806
rect 5323 716 5577 772
rect 5323 682 5357 716
rect 5391 682 5510 716
rect 5544 682 5577 716
rect 5323 626 5577 682
rect 5323 592 5357 626
rect 5391 592 5510 626
rect 5544 592 5577 626
rect 5323 536 5577 592
rect 5323 502 5357 536
rect 5391 502 5510 536
rect 5544 502 5577 536
rect 3983 412 4017 446
rect 4051 412 4170 446
rect 4204 412 4237 446
rect 3983 397 4237 412
rect 5323 446 5577 502
rect 6663 1402 6697 1436
rect 6731 1402 6850 1436
rect 6884 1402 6917 1436
rect 8003 1436 8257 1483
rect 6663 1346 6917 1402
rect 6663 1312 6697 1346
rect 6731 1312 6850 1346
rect 6884 1312 6917 1346
rect 6663 1256 6917 1312
rect 6663 1222 6697 1256
rect 6731 1222 6850 1256
rect 6884 1222 6917 1256
rect 6663 1166 6917 1222
rect 6663 1132 6697 1166
rect 6731 1132 6850 1166
rect 6884 1132 6917 1166
rect 6663 1076 6917 1132
rect 6663 1042 6697 1076
rect 6731 1042 6850 1076
rect 6884 1042 6917 1076
rect 6663 986 6917 1042
rect 6663 952 6697 986
rect 6731 952 6850 986
rect 6884 952 6917 986
rect 6663 896 6917 952
rect 6663 862 6697 896
rect 6731 862 6850 896
rect 6884 862 6917 896
rect 6663 806 6917 862
rect 6663 772 6697 806
rect 6731 772 6850 806
rect 6884 772 6917 806
rect 6663 716 6917 772
rect 6663 682 6697 716
rect 6731 682 6850 716
rect 6884 682 6917 716
rect 6663 626 6917 682
rect 6663 592 6697 626
rect 6731 592 6850 626
rect 6884 592 6917 626
rect 6663 536 6917 592
rect 6663 502 6697 536
rect 6731 502 6850 536
rect 6884 502 6917 536
rect 5323 412 5357 446
rect 5391 412 5510 446
rect 5544 412 5577 446
rect 5323 397 5577 412
rect 6663 446 6917 502
rect 8003 1402 8037 1436
rect 8071 1402 8190 1436
rect 8224 1402 8257 1436
rect 9343 1436 9444 1483
rect 8003 1346 8257 1402
rect 8003 1312 8037 1346
rect 8071 1312 8190 1346
rect 8224 1312 8257 1346
rect 8003 1256 8257 1312
rect 8003 1222 8037 1256
rect 8071 1222 8190 1256
rect 8224 1222 8257 1256
rect 8003 1166 8257 1222
rect 8003 1132 8037 1166
rect 8071 1132 8190 1166
rect 8224 1132 8257 1166
rect 8003 1076 8257 1132
rect 8003 1042 8037 1076
rect 8071 1042 8190 1076
rect 8224 1042 8257 1076
rect 8003 986 8257 1042
rect 8003 952 8037 986
rect 8071 952 8190 986
rect 8224 952 8257 986
rect 8003 896 8257 952
rect 8003 862 8037 896
rect 8071 862 8190 896
rect 8224 862 8257 896
rect 8003 806 8257 862
rect 8003 772 8037 806
rect 8071 772 8190 806
rect 8224 772 8257 806
rect 8003 716 8257 772
rect 8003 682 8037 716
rect 8071 682 8190 716
rect 8224 682 8257 716
rect 8003 626 8257 682
rect 8003 592 8037 626
rect 8071 592 8190 626
rect 8224 592 8257 626
rect 8003 536 8257 592
rect 8003 502 8037 536
rect 8071 502 8190 536
rect 8224 502 8257 536
rect 6663 412 6697 446
rect 6731 412 6850 446
rect 6884 412 6917 446
rect 6663 397 6917 412
rect 8003 446 8257 502
rect 9343 1402 9377 1436
rect 9411 1402 9444 1436
rect 9343 1346 9444 1402
rect 9343 1312 9377 1346
rect 9411 1312 9444 1346
rect 9343 1256 9444 1312
rect 9343 1222 9377 1256
rect 9411 1222 9444 1256
rect 9343 1166 9444 1222
rect 9343 1132 9377 1166
rect 9411 1132 9444 1166
rect 9343 1076 9444 1132
rect 9343 1042 9377 1076
rect 9411 1042 9444 1076
rect 9343 986 9444 1042
rect 9343 952 9377 986
rect 9411 952 9444 986
rect 9343 896 9444 952
rect 9343 862 9377 896
rect 9411 862 9444 896
rect 9343 806 9444 862
rect 9343 772 9377 806
rect 9411 772 9444 806
rect 9343 716 9444 772
rect 9343 682 9377 716
rect 9411 682 9444 716
rect 9343 626 9444 682
rect 9343 592 9377 626
rect 9411 592 9444 626
rect 9343 536 9444 592
rect 9343 502 9377 536
rect 9411 502 9444 536
rect 8003 412 8037 446
rect 8071 412 8190 446
rect 8224 412 8257 446
rect 8003 397 8257 412
rect 9343 446 9444 502
rect 9343 412 9377 446
rect 9411 412 9444 446
rect 9343 397 9444 412
rect 116 362 9444 397
rect 116 328 246 362
rect 280 328 336 362
rect 370 328 426 362
rect 460 328 516 362
rect 550 328 606 362
rect 640 328 696 362
rect 730 328 786 362
rect 820 328 876 362
rect 910 328 966 362
rect 1000 328 1056 362
rect 1090 328 1146 362
rect 1180 328 1236 362
rect 1270 328 1586 362
rect 1620 328 1676 362
rect 1710 328 1766 362
rect 1800 328 1856 362
rect 1890 328 1946 362
rect 1980 328 2036 362
rect 2070 328 2126 362
rect 2160 328 2216 362
rect 2250 328 2306 362
rect 2340 328 2396 362
rect 2430 328 2486 362
rect 2520 328 2576 362
rect 2610 328 2926 362
rect 2960 328 3016 362
rect 3050 328 3106 362
rect 3140 328 3196 362
rect 3230 328 3286 362
rect 3320 328 3376 362
rect 3410 328 3466 362
rect 3500 328 3556 362
rect 3590 328 3646 362
rect 3680 328 3736 362
rect 3770 328 3826 362
rect 3860 328 3916 362
rect 3950 328 4266 362
rect 4300 328 4356 362
rect 4390 328 4446 362
rect 4480 328 4536 362
rect 4570 328 4626 362
rect 4660 328 4716 362
rect 4750 328 4806 362
rect 4840 328 4896 362
rect 4930 328 4986 362
rect 5020 328 5076 362
rect 5110 328 5166 362
rect 5200 328 5256 362
rect 5290 328 5606 362
rect 5640 328 5696 362
rect 5730 328 5786 362
rect 5820 328 5876 362
rect 5910 328 5966 362
rect 6000 328 6056 362
rect 6090 328 6146 362
rect 6180 328 6236 362
rect 6270 328 6326 362
rect 6360 328 6416 362
rect 6450 328 6506 362
rect 6540 328 6596 362
rect 6630 328 6946 362
rect 6980 328 7036 362
rect 7070 328 7126 362
rect 7160 328 7216 362
rect 7250 328 7306 362
rect 7340 328 7396 362
rect 7430 328 7486 362
rect 7520 328 7576 362
rect 7610 328 7666 362
rect 7700 328 7756 362
rect 7790 328 7846 362
rect 7880 328 7936 362
rect 7970 328 8286 362
rect 8320 328 8376 362
rect 8410 328 8466 362
rect 8500 328 8556 362
rect 8590 328 8646 362
rect 8680 328 8736 362
rect 8770 328 8826 362
rect 8860 328 8916 362
rect 8950 328 9006 362
rect 9040 328 9096 362
rect 9130 328 9186 362
rect 9220 328 9276 362
rect 9310 328 9444 362
rect 116 296 9444 328
<< nsubdiff >>
rect 279 1402 1241 1421
rect 279 1368 410 1402
rect 444 1368 500 1402
rect 534 1368 590 1402
rect 624 1368 680 1402
rect 714 1368 770 1402
rect 804 1368 860 1402
rect 894 1368 950 1402
rect 984 1368 1040 1402
rect 1074 1368 1130 1402
rect 1164 1368 1241 1402
rect 279 1349 1241 1368
rect 279 1345 351 1349
rect 279 1311 298 1345
rect 332 1311 351 1345
rect 279 1255 351 1311
rect 1169 1326 1241 1349
rect 1169 1292 1188 1326
rect 1222 1292 1241 1326
rect 279 1221 298 1255
rect 332 1221 351 1255
rect 279 1165 351 1221
rect 279 1131 298 1165
rect 332 1131 351 1165
rect 279 1075 351 1131
rect 279 1041 298 1075
rect 332 1041 351 1075
rect 279 985 351 1041
rect 279 951 298 985
rect 332 951 351 985
rect 279 895 351 951
rect 279 861 298 895
rect 332 861 351 895
rect 279 805 351 861
rect 279 771 298 805
rect 332 771 351 805
rect 279 715 351 771
rect 279 681 298 715
rect 332 681 351 715
rect 279 625 351 681
rect 279 591 298 625
rect 332 591 351 625
rect 1169 1236 1241 1292
rect 1169 1202 1188 1236
rect 1222 1202 1241 1236
rect 1169 1146 1241 1202
rect 1169 1112 1188 1146
rect 1222 1112 1241 1146
rect 1169 1056 1241 1112
rect 1169 1022 1188 1056
rect 1222 1022 1241 1056
rect 1169 966 1241 1022
rect 1169 932 1188 966
rect 1222 932 1241 966
rect 1169 876 1241 932
rect 1169 842 1188 876
rect 1222 842 1241 876
rect 1169 786 1241 842
rect 1169 752 1188 786
rect 1222 752 1241 786
rect 1169 696 1241 752
rect 1169 662 1188 696
rect 1222 662 1241 696
rect 1169 606 1241 662
rect 279 531 351 591
rect 1169 572 1188 606
rect 1222 572 1241 606
rect 1169 531 1241 572
rect 279 512 1241 531
rect 279 478 376 512
rect 410 478 466 512
rect 500 478 556 512
rect 590 478 646 512
rect 680 478 736 512
rect 770 478 826 512
rect 860 478 916 512
rect 950 478 1006 512
rect 1040 478 1096 512
rect 1130 478 1241 512
rect 279 459 1241 478
rect 1619 1402 2581 1421
rect 1619 1368 1750 1402
rect 1784 1368 1840 1402
rect 1874 1368 1930 1402
rect 1964 1368 2020 1402
rect 2054 1368 2110 1402
rect 2144 1368 2200 1402
rect 2234 1368 2290 1402
rect 2324 1368 2380 1402
rect 2414 1368 2470 1402
rect 2504 1368 2581 1402
rect 1619 1349 2581 1368
rect 1619 1345 1691 1349
rect 1619 1311 1638 1345
rect 1672 1311 1691 1345
rect 1619 1255 1691 1311
rect 2509 1326 2581 1349
rect 2509 1292 2528 1326
rect 2562 1292 2581 1326
rect 1619 1221 1638 1255
rect 1672 1221 1691 1255
rect 1619 1165 1691 1221
rect 1619 1131 1638 1165
rect 1672 1131 1691 1165
rect 1619 1075 1691 1131
rect 1619 1041 1638 1075
rect 1672 1041 1691 1075
rect 1619 985 1691 1041
rect 1619 951 1638 985
rect 1672 951 1691 985
rect 1619 895 1691 951
rect 1619 861 1638 895
rect 1672 861 1691 895
rect 1619 805 1691 861
rect 1619 771 1638 805
rect 1672 771 1691 805
rect 1619 715 1691 771
rect 1619 681 1638 715
rect 1672 681 1691 715
rect 1619 625 1691 681
rect 1619 591 1638 625
rect 1672 591 1691 625
rect 2509 1236 2581 1292
rect 2509 1202 2528 1236
rect 2562 1202 2581 1236
rect 2509 1146 2581 1202
rect 2509 1112 2528 1146
rect 2562 1112 2581 1146
rect 2509 1056 2581 1112
rect 2509 1022 2528 1056
rect 2562 1022 2581 1056
rect 2509 966 2581 1022
rect 2509 932 2528 966
rect 2562 932 2581 966
rect 2509 876 2581 932
rect 2509 842 2528 876
rect 2562 842 2581 876
rect 2509 786 2581 842
rect 2509 752 2528 786
rect 2562 752 2581 786
rect 2509 696 2581 752
rect 2509 662 2528 696
rect 2562 662 2581 696
rect 2509 606 2581 662
rect 1619 531 1691 591
rect 2509 572 2528 606
rect 2562 572 2581 606
rect 2509 531 2581 572
rect 1619 512 2581 531
rect 1619 478 1716 512
rect 1750 478 1806 512
rect 1840 478 1896 512
rect 1930 478 1986 512
rect 2020 478 2076 512
rect 2110 478 2166 512
rect 2200 478 2256 512
rect 2290 478 2346 512
rect 2380 478 2436 512
rect 2470 478 2581 512
rect 1619 459 2581 478
rect 2959 1402 3921 1421
rect 2959 1368 3090 1402
rect 3124 1368 3180 1402
rect 3214 1368 3270 1402
rect 3304 1368 3360 1402
rect 3394 1368 3450 1402
rect 3484 1368 3540 1402
rect 3574 1368 3630 1402
rect 3664 1368 3720 1402
rect 3754 1368 3810 1402
rect 3844 1368 3921 1402
rect 2959 1349 3921 1368
rect 2959 1345 3031 1349
rect 2959 1311 2978 1345
rect 3012 1311 3031 1345
rect 2959 1255 3031 1311
rect 3849 1326 3921 1349
rect 3849 1292 3868 1326
rect 3902 1292 3921 1326
rect 2959 1221 2978 1255
rect 3012 1221 3031 1255
rect 2959 1165 3031 1221
rect 2959 1131 2978 1165
rect 3012 1131 3031 1165
rect 2959 1075 3031 1131
rect 2959 1041 2978 1075
rect 3012 1041 3031 1075
rect 2959 985 3031 1041
rect 2959 951 2978 985
rect 3012 951 3031 985
rect 2959 895 3031 951
rect 2959 861 2978 895
rect 3012 861 3031 895
rect 2959 805 3031 861
rect 2959 771 2978 805
rect 3012 771 3031 805
rect 2959 715 3031 771
rect 2959 681 2978 715
rect 3012 681 3031 715
rect 2959 625 3031 681
rect 2959 591 2978 625
rect 3012 591 3031 625
rect 3849 1236 3921 1292
rect 3849 1202 3868 1236
rect 3902 1202 3921 1236
rect 3849 1146 3921 1202
rect 3849 1112 3868 1146
rect 3902 1112 3921 1146
rect 3849 1056 3921 1112
rect 3849 1022 3868 1056
rect 3902 1022 3921 1056
rect 3849 966 3921 1022
rect 3849 932 3868 966
rect 3902 932 3921 966
rect 3849 876 3921 932
rect 3849 842 3868 876
rect 3902 842 3921 876
rect 3849 786 3921 842
rect 3849 752 3868 786
rect 3902 752 3921 786
rect 3849 696 3921 752
rect 3849 662 3868 696
rect 3902 662 3921 696
rect 3849 606 3921 662
rect 2959 531 3031 591
rect 3849 572 3868 606
rect 3902 572 3921 606
rect 3849 531 3921 572
rect 2959 512 3921 531
rect 2959 478 3056 512
rect 3090 478 3146 512
rect 3180 478 3236 512
rect 3270 478 3326 512
rect 3360 478 3416 512
rect 3450 478 3506 512
rect 3540 478 3596 512
rect 3630 478 3686 512
rect 3720 478 3776 512
rect 3810 478 3921 512
rect 2959 459 3921 478
rect 4299 1402 5261 1421
rect 4299 1368 4430 1402
rect 4464 1368 4520 1402
rect 4554 1368 4610 1402
rect 4644 1368 4700 1402
rect 4734 1368 4790 1402
rect 4824 1368 4880 1402
rect 4914 1368 4970 1402
rect 5004 1368 5060 1402
rect 5094 1368 5150 1402
rect 5184 1368 5261 1402
rect 4299 1349 5261 1368
rect 4299 1345 4371 1349
rect 4299 1311 4318 1345
rect 4352 1311 4371 1345
rect 4299 1255 4371 1311
rect 5189 1326 5261 1349
rect 5189 1292 5208 1326
rect 5242 1292 5261 1326
rect 4299 1221 4318 1255
rect 4352 1221 4371 1255
rect 4299 1165 4371 1221
rect 4299 1131 4318 1165
rect 4352 1131 4371 1165
rect 4299 1075 4371 1131
rect 4299 1041 4318 1075
rect 4352 1041 4371 1075
rect 4299 985 4371 1041
rect 4299 951 4318 985
rect 4352 951 4371 985
rect 4299 895 4371 951
rect 4299 861 4318 895
rect 4352 861 4371 895
rect 4299 805 4371 861
rect 4299 771 4318 805
rect 4352 771 4371 805
rect 4299 715 4371 771
rect 4299 681 4318 715
rect 4352 681 4371 715
rect 4299 625 4371 681
rect 4299 591 4318 625
rect 4352 591 4371 625
rect 5189 1236 5261 1292
rect 5189 1202 5208 1236
rect 5242 1202 5261 1236
rect 5189 1146 5261 1202
rect 5189 1112 5208 1146
rect 5242 1112 5261 1146
rect 5189 1056 5261 1112
rect 5189 1022 5208 1056
rect 5242 1022 5261 1056
rect 5189 966 5261 1022
rect 5189 932 5208 966
rect 5242 932 5261 966
rect 5189 876 5261 932
rect 5189 842 5208 876
rect 5242 842 5261 876
rect 5189 786 5261 842
rect 5189 752 5208 786
rect 5242 752 5261 786
rect 5189 696 5261 752
rect 5189 662 5208 696
rect 5242 662 5261 696
rect 5189 606 5261 662
rect 4299 531 4371 591
rect 5189 572 5208 606
rect 5242 572 5261 606
rect 5189 531 5261 572
rect 4299 512 5261 531
rect 4299 478 4396 512
rect 4430 478 4486 512
rect 4520 478 4576 512
rect 4610 478 4666 512
rect 4700 478 4756 512
rect 4790 478 4846 512
rect 4880 478 4936 512
rect 4970 478 5026 512
rect 5060 478 5116 512
rect 5150 478 5261 512
rect 4299 459 5261 478
rect 5639 1402 6601 1421
rect 5639 1368 5770 1402
rect 5804 1368 5860 1402
rect 5894 1368 5950 1402
rect 5984 1368 6040 1402
rect 6074 1368 6130 1402
rect 6164 1368 6220 1402
rect 6254 1368 6310 1402
rect 6344 1368 6400 1402
rect 6434 1368 6490 1402
rect 6524 1368 6601 1402
rect 5639 1349 6601 1368
rect 5639 1345 5711 1349
rect 5639 1311 5658 1345
rect 5692 1311 5711 1345
rect 5639 1255 5711 1311
rect 6529 1326 6601 1349
rect 6529 1292 6548 1326
rect 6582 1292 6601 1326
rect 5639 1221 5658 1255
rect 5692 1221 5711 1255
rect 5639 1165 5711 1221
rect 5639 1131 5658 1165
rect 5692 1131 5711 1165
rect 5639 1075 5711 1131
rect 5639 1041 5658 1075
rect 5692 1041 5711 1075
rect 5639 985 5711 1041
rect 5639 951 5658 985
rect 5692 951 5711 985
rect 5639 895 5711 951
rect 5639 861 5658 895
rect 5692 861 5711 895
rect 5639 805 5711 861
rect 5639 771 5658 805
rect 5692 771 5711 805
rect 5639 715 5711 771
rect 5639 681 5658 715
rect 5692 681 5711 715
rect 5639 625 5711 681
rect 5639 591 5658 625
rect 5692 591 5711 625
rect 6529 1236 6601 1292
rect 6529 1202 6548 1236
rect 6582 1202 6601 1236
rect 6529 1146 6601 1202
rect 6529 1112 6548 1146
rect 6582 1112 6601 1146
rect 6529 1056 6601 1112
rect 6529 1022 6548 1056
rect 6582 1022 6601 1056
rect 6529 966 6601 1022
rect 6529 932 6548 966
rect 6582 932 6601 966
rect 6529 876 6601 932
rect 6529 842 6548 876
rect 6582 842 6601 876
rect 6529 786 6601 842
rect 6529 752 6548 786
rect 6582 752 6601 786
rect 6529 696 6601 752
rect 6529 662 6548 696
rect 6582 662 6601 696
rect 6529 606 6601 662
rect 5639 531 5711 591
rect 6529 572 6548 606
rect 6582 572 6601 606
rect 6529 531 6601 572
rect 5639 512 6601 531
rect 5639 478 5736 512
rect 5770 478 5826 512
rect 5860 478 5916 512
rect 5950 478 6006 512
rect 6040 478 6096 512
rect 6130 478 6186 512
rect 6220 478 6276 512
rect 6310 478 6366 512
rect 6400 478 6456 512
rect 6490 478 6601 512
rect 5639 459 6601 478
rect 6979 1402 7941 1421
rect 6979 1368 7110 1402
rect 7144 1368 7200 1402
rect 7234 1368 7290 1402
rect 7324 1368 7380 1402
rect 7414 1368 7470 1402
rect 7504 1368 7560 1402
rect 7594 1368 7650 1402
rect 7684 1368 7740 1402
rect 7774 1368 7830 1402
rect 7864 1368 7941 1402
rect 6979 1349 7941 1368
rect 6979 1345 7051 1349
rect 6979 1311 6998 1345
rect 7032 1311 7051 1345
rect 6979 1255 7051 1311
rect 7869 1326 7941 1349
rect 7869 1292 7888 1326
rect 7922 1292 7941 1326
rect 6979 1221 6998 1255
rect 7032 1221 7051 1255
rect 6979 1165 7051 1221
rect 6979 1131 6998 1165
rect 7032 1131 7051 1165
rect 6979 1075 7051 1131
rect 6979 1041 6998 1075
rect 7032 1041 7051 1075
rect 6979 985 7051 1041
rect 6979 951 6998 985
rect 7032 951 7051 985
rect 6979 895 7051 951
rect 6979 861 6998 895
rect 7032 861 7051 895
rect 6979 805 7051 861
rect 6979 771 6998 805
rect 7032 771 7051 805
rect 6979 715 7051 771
rect 6979 681 6998 715
rect 7032 681 7051 715
rect 6979 625 7051 681
rect 6979 591 6998 625
rect 7032 591 7051 625
rect 7869 1236 7941 1292
rect 7869 1202 7888 1236
rect 7922 1202 7941 1236
rect 7869 1146 7941 1202
rect 7869 1112 7888 1146
rect 7922 1112 7941 1146
rect 7869 1056 7941 1112
rect 7869 1022 7888 1056
rect 7922 1022 7941 1056
rect 7869 966 7941 1022
rect 7869 932 7888 966
rect 7922 932 7941 966
rect 7869 876 7941 932
rect 7869 842 7888 876
rect 7922 842 7941 876
rect 7869 786 7941 842
rect 7869 752 7888 786
rect 7922 752 7941 786
rect 7869 696 7941 752
rect 7869 662 7888 696
rect 7922 662 7941 696
rect 7869 606 7941 662
rect 6979 531 7051 591
rect 7869 572 7888 606
rect 7922 572 7941 606
rect 7869 531 7941 572
rect 6979 512 7941 531
rect 6979 478 7076 512
rect 7110 478 7166 512
rect 7200 478 7256 512
rect 7290 478 7346 512
rect 7380 478 7436 512
rect 7470 478 7526 512
rect 7560 478 7616 512
rect 7650 478 7706 512
rect 7740 478 7796 512
rect 7830 478 7941 512
rect 6979 459 7941 478
rect 8319 1402 9281 1421
rect 8319 1368 8450 1402
rect 8484 1368 8540 1402
rect 8574 1368 8630 1402
rect 8664 1368 8720 1402
rect 8754 1368 8810 1402
rect 8844 1368 8900 1402
rect 8934 1368 8990 1402
rect 9024 1368 9080 1402
rect 9114 1368 9170 1402
rect 9204 1368 9281 1402
rect 8319 1349 9281 1368
rect 8319 1345 8391 1349
rect 8319 1311 8338 1345
rect 8372 1311 8391 1345
rect 8319 1255 8391 1311
rect 9209 1326 9281 1349
rect 9209 1292 9228 1326
rect 9262 1292 9281 1326
rect 8319 1221 8338 1255
rect 8372 1221 8391 1255
rect 8319 1165 8391 1221
rect 8319 1131 8338 1165
rect 8372 1131 8391 1165
rect 8319 1075 8391 1131
rect 8319 1041 8338 1075
rect 8372 1041 8391 1075
rect 8319 985 8391 1041
rect 8319 951 8338 985
rect 8372 951 8391 985
rect 8319 895 8391 951
rect 8319 861 8338 895
rect 8372 861 8391 895
rect 8319 805 8391 861
rect 8319 771 8338 805
rect 8372 771 8391 805
rect 8319 715 8391 771
rect 8319 681 8338 715
rect 8372 681 8391 715
rect 8319 625 8391 681
rect 8319 591 8338 625
rect 8372 591 8391 625
rect 9209 1236 9281 1292
rect 9209 1202 9228 1236
rect 9262 1202 9281 1236
rect 9209 1146 9281 1202
rect 9209 1112 9228 1146
rect 9262 1112 9281 1146
rect 9209 1056 9281 1112
rect 9209 1022 9228 1056
rect 9262 1022 9281 1056
rect 9209 966 9281 1022
rect 9209 932 9228 966
rect 9262 932 9281 966
rect 9209 876 9281 932
rect 9209 842 9228 876
rect 9262 842 9281 876
rect 9209 786 9281 842
rect 9209 752 9228 786
rect 9262 752 9281 786
rect 9209 696 9281 752
rect 9209 662 9228 696
rect 9262 662 9281 696
rect 9209 606 9281 662
rect 8319 531 8391 591
rect 9209 572 9228 606
rect 9262 572 9281 606
rect 9209 531 9281 572
rect 8319 512 9281 531
rect 8319 478 8416 512
rect 8450 478 8506 512
rect 8540 478 8596 512
rect 8630 478 8686 512
rect 8720 478 8776 512
rect 8810 478 8866 512
rect 8900 478 8956 512
rect 8990 478 9046 512
rect 9080 478 9136 512
rect 9170 478 9281 512
rect 8319 459 9281 478
<< psubdiffcont >>
rect 150 1492 184 1526
rect 246 1515 280 1549
rect 336 1515 370 1549
rect 426 1515 460 1549
rect 516 1515 550 1549
rect 606 1515 640 1549
rect 696 1515 730 1549
rect 786 1515 820 1549
rect 876 1515 910 1549
rect 966 1515 1000 1549
rect 1056 1515 1090 1549
rect 1146 1515 1180 1549
rect 1236 1515 1270 1549
rect 1337 1492 1371 1526
rect 1490 1492 1524 1526
rect 1586 1515 1620 1549
rect 1676 1515 1710 1549
rect 1766 1515 1800 1549
rect 1856 1515 1890 1549
rect 1946 1515 1980 1549
rect 2036 1515 2070 1549
rect 2126 1515 2160 1549
rect 2216 1515 2250 1549
rect 2306 1515 2340 1549
rect 2396 1515 2430 1549
rect 2486 1515 2520 1549
rect 2576 1515 2610 1549
rect 2677 1492 2711 1526
rect 2830 1492 2864 1526
rect 2926 1515 2960 1549
rect 3016 1515 3050 1549
rect 3106 1515 3140 1549
rect 3196 1515 3230 1549
rect 3286 1515 3320 1549
rect 3376 1515 3410 1549
rect 3466 1515 3500 1549
rect 3556 1515 3590 1549
rect 3646 1515 3680 1549
rect 3736 1515 3770 1549
rect 3826 1515 3860 1549
rect 3916 1515 3950 1549
rect 4017 1492 4051 1526
rect 4170 1492 4204 1526
rect 4266 1515 4300 1549
rect 4356 1515 4390 1549
rect 4446 1515 4480 1549
rect 4536 1515 4570 1549
rect 4626 1515 4660 1549
rect 4716 1515 4750 1549
rect 4806 1515 4840 1549
rect 4896 1515 4930 1549
rect 4986 1515 5020 1549
rect 5076 1515 5110 1549
rect 5166 1515 5200 1549
rect 5256 1515 5290 1549
rect 5357 1492 5391 1526
rect 5510 1492 5544 1526
rect 5606 1515 5640 1549
rect 5696 1515 5730 1549
rect 5786 1515 5820 1549
rect 5876 1515 5910 1549
rect 5966 1515 6000 1549
rect 6056 1515 6090 1549
rect 6146 1515 6180 1549
rect 6236 1515 6270 1549
rect 6326 1515 6360 1549
rect 6416 1515 6450 1549
rect 6506 1515 6540 1549
rect 6596 1515 6630 1549
rect 6697 1492 6731 1526
rect 6850 1492 6884 1526
rect 6946 1515 6980 1549
rect 7036 1515 7070 1549
rect 7126 1515 7160 1549
rect 7216 1515 7250 1549
rect 7306 1515 7340 1549
rect 7396 1515 7430 1549
rect 7486 1515 7520 1549
rect 7576 1515 7610 1549
rect 7666 1515 7700 1549
rect 7756 1515 7790 1549
rect 7846 1515 7880 1549
rect 7936 1515 7970 1549
rect 8037 1492 8071 1526
rect 8190 1492 8224 1526
rect 8286 1515 8320 1549
rect 8376 1515 8410 1549
rect 8466 1515 8500 1549
rect 8556 1515 8590 1549
rect 8646 1515 8680 1549
rect 8736 1515 8770 1549
rect 8826 1515 8860 1549
rect 8916 1515 8950 1549
rect 9006 1515 9040 1549
rect 9096 1515 9130 1549
rect 9186 1515 9220 1549
rect 9276 1515 9310 1549
rect 9377 1492 9411 1526
rect 150 1402 184 1436
rect 150 1312 184 1346
rect 150 1222 184 1256
rect 150 1132 184 1166
rect 150 1042 184 1076
rect 150 952 184 986
rect 150 862 184 896
rect 150 772 184 806
rect 150 682 184 716
rect 150 592 184 626
rect 150 502 184 536
rect 1337 1402 1371 1436
rect 1490 1402 1524 1436
rect 1337 1312 1371 1346
rect 1490 1312 1524 1346
rect 1337 1222 1371 1256
rect 1490 1222 1524 1256
rect 1337 1132 1371 1166
rect 1490 1132 1524 1166
rect 1337 1042 1371 1076
rect 1490 1042 1524 1076
rect 1337 952 1371 986
rect 1490 952 1524 986
rect 1337 862 1371 896
rect 1490 862 1524 896
rect 1337 772 1371 806
rect 1490 772 1524 806
rect 1337 682 1371 716
rect 1490 682 1524 716
rect 1337 592 1371 626
rect 1490 592 1524 626
rect 1337 502 1371 536
rect 1490 502 1524 536
rect 150 412 184 446
rect 2677 1402 2711 1436
rect 2830 1402 2864 1436
rect 2677 1312 2711 1346
rect 2830 1312 2864 1346
rect 2677 1222 2711 1256
rect 2830 1222 2864 1256
rect 2677 1132 2711 1166
rect 2830 1132 2864 1166
rect 2677 1042 2711 1076
rect 2830 1042 2864 1076
rect 2677 952 2711 986
rect 2830 952 2864 986
rect 2677 862 2711 896
rect 2830 862 2864 896
rect 2677 772 2711 806
rect 2830 772 2864 806
rect 2677 682 2711 716
rect 2830 682 2864 716
rect 2677 592 2711 626
rect 2830 592 2864 626
rect 2677 502 2711 536
rect 2830 502 2864 536
rect 1337 412 1371 446
rect 1490 412 1524 446
rect 4017 1402 4051 1436
rect 4170 1402 4204 1436
rect 4017 1312 4051 1346
rect 4170 1312 4204 1346
rect 4017 1222 4051 1256
rect 4170 1222 4204 1256
rect 4017 1132 4051 1166
rect 4170 1132 4204 1166
rect 4017 1042 4051 1076
rect 4170 1042 4204 1076
rect 4017 952 4051 986
rect 4170 952 4204 986
rect 4017 862 4051 896
rect 4170 862 4204 896
rect 4017 772 4051 806
rect 4170 772 4204 806
rect 4017 682 4051 716
rect 4170 682 4204 716
rect 4017 592 4051 626
rect 4170 592 4204 626
rect 4017 502 4051 536
rect 4170 502 4204 536
rect 2677 412 2711 446
rect 2830 412 2864 446
rect 5357 1402 5391 1436
rect 5510 1402 5544 1436
rect 5357 1312 5391 1346
rect 5510 1312 5544 1346
rect 5357 1222 5391 1256
rect 5510 1222 5544 1256
rect 5357 1132 5391 1166
rect 5510 1132 5544 1166
rect 5357 1042 5391 1076
rect 5510 1042 5544 1076
rect 5357 952 5391 986
rect 5510 952 5544 986
rect 5357 862 5391 896
rect 5510 862 5544 896
rect 5357 772 5391 806
rect 5510 772 5544 806
rect 5357 682 5391 716
rect 5510 682 5544 716
rect 5357 592 5391 626
rect 5510 592 5544 626
rect 5357 502 5391 536
rect 5510 502 5544 536
rect 4017 412 4051 446
rect 4170 412 4204 446
rect 6697 1402 6731 1436
rect 6850 1402 6884 1436
rect 6697 1312 6731 1346
rect 6850 1312 6884 1346
rect 6697 1222 6731 1256
rect 6850 1222 6884 1256
rect 6697 1132 6731 1166
rect 6850 1132 6884 1166
rect 6697 1042 6731 1076
rect 6850 1042 6884 1076
rect 6697 952 6731 986
rect 6850 952 6884 986
rect 6697 862 6731 896
rect 6850 862 6884 896
rect 6697 772 6731 806
rect 6850 772 6884 806
rect 6697 682 6731 716
rect 6850 682 6884 716
rect 6697 592 6731 626
rect 6850 592 6884 626
rect 6697 502 6731 536
rect 6850 502 6884 536
rect 5357 412 5391 446
rect 5510 412 5544 446
rect 8037 1402 8071 1436
rect 8190 1402 8224 1436
rect 8037 1312 8071 1346
rect 8190 1312 8224 1346
rect 8037 1222 8071 1256
rect 8190 1222 8224 1256
rect 8037 1132 8071 1166
rect 8190 1132 8224 1166
rect 8037 1042 8071 1076
rect 8190 1042 8224 1076
rect 8037 952 8071 986
rect 8190 952 8224 986
rect 8037 862 8071 896
rect 8190 862 8224 896
rect 8037 772 8071 806
rect 8190 772 8224 806
rect 8037 682 8071 716
rect 8190 682 8224 716
rect 8037 592 8071 626
rect 8190 592 8224 626
rect 8037 502 8071 536
rect 8190 502 8224 536
rect 6697 412 6731 446
rect 6850 412 6884 446
rect 9377 1402 9411 1436
rect 9377 1312 9411 1346
rect 9377 1222 9411 1256
rect 9377 1132 9411 1166
rect 9377 1042 9411 1076
rect 9377 952 9411 986
rect 9377 862 9411 896
rect 9377 772 9411 806
rect 9377 682 9411 716
rect 9377 592 9411 626
rect 9377 502 9411 536
rect 8037 412 8071 446
rect 8190 412 8224 446
rect 9377 412 9411 446
rect 246 328 280 362
rect 336 328 370 362
rect 426 328 460 362
rect 516 328 550 362
rect 606 328 640 362
rect 696 328 730 362
rect 786 328 820 362
rect 876 328 910 362
rect 966 328 1000 362
rect 1056 328 1090 362
rect 1146 328 1180 362
rect 1236 328 1270 362
rect 1586 328 1620 362
rect 1676 328 1710 362
rect 1766 328 1800 362
rect 1856 328 1890 362
rect 1946 328 1980 362
rect 2036 328 2070 362
rect 2126 328 2160 362
rect 2216 328 2250 362
rect 2306 328 2340 362
rect 2396 328 2430 362
rect 2486 328 2520 362
rect 2576 328 2610 362
rect 2926 328 2960 362
rect 3016 328 3050 362
rect 3106 328 3140 362
rect 3196 328 3230 362
rect 3286 328 3320 362
rect 3376 328 3410 362
rect 3466 328 3500 362
rect 3556 328 3590 362
rect 3646 328 3680 362
rect 3736 328 3770 362
rect 3826 328 3860 362
rect 3916 328 3950 362
rect 4266 328 4300 362
rect 4356 328 4390 362
rect 4446 328 4480 362
rect 4536 328 4570 362
rect 4626 328 4660 362
rect 4716 328 4750 362
rect 4806 328 4840 362
rect 4896 328 4930 362
rect 4986 328 5020 362
rect 5076 328 5110 362
rect 5166 328 5200 362
rect 5256 328 5290 362
rect 5606 328 5640 362
rect 5696 328 5730 362
rect 5786 328 5820 362
rect 5876 328 5910 362
rect 5966 328 6000 362
rect 6056 328 6090 362
rect 6146 328 6180 362
rect 6236 328 6270 362
rect 6326 328 6360 362
rect 6416 328 6450 362
rect 6506 328 6540 362
rect 6596 328 6630 362
rect 6946 328 6980 362
rect 7036 328 7070 362
rect 7126 328 7160 362
rect 7216 328 7250 362
rect 7306 328 7340 362
rect 7396 328 7430 362
rect 7486 328 7520 362
rect 7576 328 7610 362
rect 7666 328 7700 362
rect 7756 328 7790 362
rect 7846 328 7880 362
rect 7936 328 7970 362
rect 8286 328 8320 362
rect 8376 328 8410 362
rect 8466 328 8500 362
rect 8556 328 8590 362
rect 8646 328 8680 362
rect 8736 328 8770 362
rect 8826 328 8860 362
rect 8916 328 8950 362
rect 9006 328 9040 362
rect 9096 328 9130 362
rect 9186 328 9220 362
rect 9276 328 9310 362
<< nsubdiffcont >>
rect 410 1368 444 1402
rect 500 1368 534 1402
rect 590 1368 624 1402
rect 680 1368 714 1402
rect 770 1368 804 1402
rect 860 1368 894 1402
rect 950 1368 984 1402
rect 1040 1368 1074 1402
rect 1130 1368 1164 1402
rect 298 1311 332 1345
rect 1188 1292 1222 1326
rect 298 1221 332 1255
rect 298 1131 332 1165
rect 298 1041 332 1075
rect 298 951 332 985
rect 298 861 332 895
rect 298 771 332 805
rect 298 681 332 715
rect 298 591 332 625
rect 1188 1202 1222 1236
rect 1188 1112 1222 1146
rect 1188 1022 1222 1056
rect 1188 932 1222 966
rect 1188 842 1222 876
rect 1188 752 1222 786
rect 1188 662 1222 696
rect 1188 572 1222 606
rect 376 478 410 512
rect 466 478 500 512
rect 556 478 590 512
rect 646 478 680 512
rect 736 478 770 512
rect 826 478 860 512
rect 916 478 950 512
rect 1006 478 1040 512
rect 1096 478 1130 512
rect 1750 1368 1784 1402
rect 1840 1368 1874 1402
rect 1930 1368 1964 1402
rect 2020 1368 2054 1402
rect 2110 1368 2144 1402
rect 2200 1368 2234 1402
rect 2290 1368 2324 1402
rect 2380 1368 2414 1402
rect 2470 1368 2504 1402
rect 1638 1311 1672 1345
rect 2528 1292 2562 1326
rect 1638 1221 1672 1255
rect 1638 1131 1672 1165
rect 1638 1041 1672 1075
rect 1638 951 1672 985
rect 1638 861 1672 895
rect 1638 771 1672 805
rect 1638 681 1672 715
rect 1638 591 1672 625
rect 2528 1202 2562 1236
rect 2528 1112 2562 1146
rect 2528 1022 2562 1056
rect 2528 932 2562 966
rect 2528 842 2562 876
rect 2528 752 2562 786
rect 2528 662 2562 696
rect 2528 572 2562 606
rect 1716 478 1750 512
rect 1806 478 1840 512
rect 1896 478 1930 512
rect 1986 478 2020 512
rect 2076 478 2110 512
rect 2166 478 2200 512
rect 2256 478 2290 512
rect 2346 478 2380 512
rect 2436 478 2470 512
rect 3090 1368 3124 1402
rect 3180 1368 3214 1402
rect 3270 1368 3304 1402
rect 3360 1368 3394 1402
rect 3450 1368 3484 1402
rect 3540 1368 3574 1402
rect 3630 1368 3664 1402
rect 3720 1368 3754 1402
rect 3810 1368 3844 1402
rect 2978 1311 3012 1345
rect 3868 1292 3902 1326
rect 2978 1221 3012 1255
rect 2978 1131 3012 1165
rect 2978 1041 3012 1075
rect 2978 951 3012 985
rect 2978 861 3012 895
rect 2978 771 3012 805
rect 2978 681 3012 715
rect 2978 591 3012 625
rect 3868 1202 3902 1236
rect 3868 1112 3902 1146
rect 3868 1022 3902 1056
rect 3868 932 3902 966
rect 3868 842 3902 876
rect 3868 752 3902 786
rect 3868 662 3902 696
rect 3868 572 3902 606
rect 3056 478 3090 512
rect 3146 478 3180 512
rect 3236 478 3270 512
rect 3326 478 3360 512
rect 3416 478 3450 512
rect 3506 478 3540 512
rect 3596 478 3630 512
rect 3686 478 3720 512
rect 3776 478 3810 512
rect 4430 1368 4464 1402
rect 4520 1368 4554 1402
rect 4610 1368 4644 1402
rect 4700 1368 4734 1402
rect 4790 1368 4824 1402
rect 4880 1368 4914 1402
rect 4970 1368 5004 1402
rect 5060 1368 5094 1402
rect 5150 1368 5184 1402
rect 4318 1311 4352 1345
rect 5208 1292 5242 1326
rect 4318 1221 4352 1255
rect 4318 1131 4352 1165
rect 4318 1041 4352 1075
rect 4318 951 4352 985
rect 4318 861 4352 895
rect 4318 771 4352 805
rect 4318 681 4352 715
rect 4318 591 4352 625
rect 5208 1202 5242 1236
rect 5208 1112 5242 1146
rect 5208 1022 5242 1056
rect 5208 932 5242 966
rect 5208 842 5242 876
rect 5208 752 5242 786
rect 5208 662 5242 696
rect 5208 572 5242 606
rect 4396 478 4430 512
rect 4486 478 4520 512
rect 4576 478 4610 512
rect 4666 478 4700 512
rect 4756 478 4790 512
rect 4846 478 4880 512
rect 4936 478 4970 512
rect 5026 478 5060 512
rect 5116 478 5150 512
rect 5770 1368 5804 1402
rect 5860 1368 5894 1402
rect 5950 1368 5984 1402
rect 6040 1368 6074 1402
rect 6130 1368 6164 1402
rect 6220 1368 6254 1402
rect 6310 1368 6344 1402
rect 6400 1368 6434 1402
rect 6490 1368 6524 1402
rect 5658 1311 5692 1345
rect 6548 1292 6582 1326
rect 5658 1221 5692 1255
rect 5658 1131 5692 1165
rect 5658 1041 5692 1075
rect 5658 951 5692 985
rect 5658 861 5692 895
rect 5658 771 5692 805
rect 5658 681 5692 715
rect 5658 591 5692 625
rect 6548 1202 6582 1236
rect 6548 1112 6582 1146
rect 6548 1022 6582 1056
rect 6548 932 6582 966
rect 6548 842 6582 876
rect 6548 752 6582 786
rect 6548 662 6582 696
rect 6548 572 6582 606
rect 5736 478 5770 512
rect 5826 478 5860 512
rect 5916 478 5950 512
rect 6006 478 6040 512
rect 6096 478 6130 512
rect 6186 478 6220 512
rect 6276 478 6310 512
rect 6366 478 6400 512
rect 6456 478 6490 512
rect 7110 1368 7144 1402
rect 7200 1368 7234 1402
rect 7290 1368 7324 1402
rect 7380 1368 7414 1402
rect 7470 1368 7504 1402
rect 7560 1368 7594 1402
rect 7650 1368 7684 1402
rect 7740 1368 7774 1402
rect 7830 1368 7864 1402
rect 6998 1311 7032 1345
rect 7888 1292 7922 1326
rect 6998 1221 7032 1255
rect 6998 1131 7032 1165
rect 6998 1041 7032 1075
rect 6998 951 7032 985
rect 6998 861 7032 895
rect 6998 771 7032 805
rect 6998 681 7032 715
rect 6998 591 7032 625
rect 7888 1202 7922 1236
rect 7888 1112 7922 1146
rect 7888 1022 7922 1056
rect 7888 932 7922 966
rect 7888 842 7922 876
rect 7888 752 7922 786
rect 7888 662 7922 696
rect 7888 572 7922 606
rect 7076 478 7110 512
rect 7166 478 7200 512
rect 7256 478 7290 512
rect 7346 478 7380 512
rect 7436 478 7470 512
rect 7526 478 7560 512
rect 7616 478 7650 512
rect 7706 478 7740 512
rect 7796 478 7830 512
rect 8450 1368 8484 1402
rect 8540 1368 8574 1402
rect 8630 1368 8664 1402
rect 8720 1368 8754 1402
rect 8810 1368 8844 1402
rect 8900 1368 8934 1402
rect 8990 1368 9024 1402
rect 9080 1368 9114 1402
rect 9170 1368 9204 1402
rect 8338 1311 8372 1345
rect 9228 1292 9262 1326
rect 8338 1221 8372 1255
rect 8338 1131 8372 1165
rect 8338 1041 8372 1075
rect 8338 951 8372 985
rect 8338 861 8372 895
rect 8338 771 8372 805
rect 8338 681 8372 715
rect 8338 591 8372 625
rect 9228 1202 9262 1236
rect 9228 1112 9262 1146
rect 9228 1022 9262 1056
rect 9228 932 9262 966
rect 9228 842 9262 876
rect 9228 752 9262 786
rect 9228 662 9262 696
rect 9228 572 9262 606
rect 8416 478 8450 512
rect 8506 478 8540 512
rect 8596 478 8630 512
rect 8686 478 8720 512
rect 8776 478 8810 512
rect 8866 478 8900 512
rect 8956 478 8990 512
rect 9046 478 9080 512
rect 9136 478 9170 512
<< locali >>
rect 90 1850 260 1910
rect 320 1850 460 1910
rect 520 1850 660 1910
rect 720 1850 860 1910
rect 920 1850 1060 1910
rect 1120 1850 1260 1910
rect 1320 1850 1460 1910
rect 1520 1850 1660 1910
rect 1720 1850 1860 1910
rect 1920 1850 2060 1910
rect 2120 1850 2260 1910
rect 2320 1850 2460 1910
rect 2520 1850 2660 1910
rect 2720 1850 2860 1910
rect 2920 1850 3060 1910
rect 3120 1850 3260 1910
rect 3320 1850 3460 1910
rect 3520 1850 3660 1910
rect 3720 1850 3860 1910
rect 3920 1850 4060 1910
rect 4120 1850 4260 1910
rect 4320 1850 4460 1910
rect 4520 1850 4660 1910
rect 4720 1850 4860 1910
rect 4920 1850 5060 1910
rect 5120 1850 5260 1910
rect 5320 1850 5460 1910
rect 5520 1850 5660 1910
rect 5720 1850 5860 1910
rect 5920 1850 6060 1910
rect 6120 1850 6260 1910
rect 6320 1850 6460 1910
rect 6520 1850 6660 1910
rect 6720 1850 6860 1910
rect 6920 1850 7060 1910
rect 7120 1850 7260 1910
rect 7320 1850 7460 1910
rect 7520 1850 7660 1910
rect 7720 1850 7860 1910
rect 7920 1850 8060 1910
rect 8120 1850 8260 1910
rect 8320 1850 8460 1910
rect 8520 1850 8660 1910
rect 8720 1850 8860 1910
rect 8920 1850 9060 1910
rect 9120 1850 9260 1910
rect 9320 1850 9470 1910
rect 116 1564 9444 1584
rect 116 1530 136 1564
rect 170 1530 226 1564
rect 260 1549 316 1564
rect 350 1549 406 1564
rect 440 1549 496 1564
rect 530 1549 586 1564
rect 620 1549 676 1564
rect 710 1549 766 1564
rect 800 1549 856 1564
rect 890 1549 946 1564
rect 980 1549 1036 1564
rect 1070 1549 1126 1564
rect 1160 1549 1216 1564
rect 1250 1549 1306 1564
rect 280 1530 316 1549
rect 370 1530 406 1549
rect 460 1530 496 1549
rect 550 1530 586 1549
rect 640 1530 676 1549
rect 730 1530 766 1549
rect 820 1530 856 1549
rect 910 1530 946 1549
rect 1000 1530 1036 1549
rect 1090 1530 1126 1549
rect 1180 1530 1216 1549
rect 1270 1530 1306 1549
rect 1340 1530 1476 1564
rect 1510 1530 1566 1564
rect 1600 1549 1656 1564
rect 1690 1549 1746 1564
rect 1780 1549 1836 1564
rect 1870 1549 1926 1564
rect 1960 1549 2016 1564
rect 2050 1549 2106 1564
rect 2140 1549 2196 1564
rect 2230 1549 2286 1564
rect 2320 1549 2376 1564
rect 2410 1549 2466 1564
rect 2500 1549 2556 1564
rect 2590 1549 2646 1564
rect 1620 1530 1656 1549
rect 1710 1530 1746 1549
rect 1800 1530 1836 1549
rect 1890 1530 1926 1549
rect 1980 1530 2016 1549
rect 2070 1530 2106 1549
rect 2160 1530 2196 1549
rect 2250 1530 2286 1549
rect 2340 1530 2376 1549
rect 2430 1530 2466 1549
rect 2520 1530 2556 1549
rect 2610 1530 2646 1549
rect 2680 1530 2816 1564
rect 2850 1530 2906 1564
rect 2940 1549 2996 1564
rect 3030 1549 3086 1564
rect 3120 1549 3176 1564
rect 3210 1549 3266 1564
rect 3300 1549 3356 1564
rect 3390 1549 3446 1564
rect 3480 1549 3536 1564
rect 3570 1549 3626 1564
rect 3660 1549 3716 1564
rect 3750 1549 3806 1564
rect 3840 1549 3896 1564
rect 3930 1549 3986 1564
rect 2960 1530 2996 1549
rect 3050 1530 3086 1549
rect 3140 1530 3176 1549
rect 3230 1530 3266 1549
rect 3320 1530 3356 1549
rect 3410 1530 3446 1549
rect 3500 1530 3536 1549
rect 3590 1530 3626 1549
rect 3680 1530 3716 1549
rect 3770 1530 3806 1549
rect 3860 1530 3896 1549
rect 3950 1530 3986 1549
rect 4020 1530 4156 1564
rect 4190 1530 4246 1564
rect 4280 1549 4336 1564
rect 4370 1549 4426 1564
rect 4460 1549 4516 1564
rect 4550 1549 4606 1564
rect 4640 1549 4696 1564
rect 4730 1549 4786 1564
rect 4820 1549 4876 1564
rect 4910 1549 4966 1564
rect 5000 1549 5056 1564
rect 5090 1549 5146 1564
rect 5180 1549 5236 1564
rect 5270 1549 5326 1564
rect 4300 1530 4336 1549
rect 4390 1530 4426 1549
rect 4480 1530 4516 1549
rect 4570 1530 4606 1549
rect 4660 1530 4696 1549
rect 4750 1530 4786 1549
rect 4840 1530 4876 1549
rect 4930 1530 4966 1549
rect 5020 1530 5056 1549
rect 5110 1530 5146 1549
rect 5200 1530 5236 1549
rect 5290 1530 5326 1549
rect 5360 1530 5496 1564
rect 5530 1530 5586 1564
rect 5620 1549 5676 1564
rect 5710 1549 5766 1564
rect 5800 1549 5856 1564
rect 5890 1549 5946 1564
rect 5980 1549 6036 1564
rect 6070 1549 6126 1564
rect 6160 1549 6216 1564
rect 6250 1549 6306 1564
rect 6340 1549 6396 1564
rect 6430 1549 6486 1564
rect 6520 1549 6576 1564
rect 6610 1549 6666 1564
rect 5640 1530 5676 1549
rect 5730 1530 5766 1549
rect 5820 1530 5856 1549
rect 5910 1530 5946 1549
rect 6000 1530 6036 1549
rect 6090 1530 6126 1549
rect 6180 1530 6216 1549
rect 6270 1530 6306 1549
rect 6360 1530 6396 1549
rect 6450 1530 6486 1549
rect 6540 1530 6576 1549
rect 6630 1530 6666 1549
rect 6700 1530 6836 1564
rect 6870 1530 6926 1564
rect 6960 1549 7016 1564
rect 7050 1549 7106 1564
rect 7140 1549 7196 1564
rect 7230 1549 7286 1564
rect 7320 1549 7376 1564
rect 7410 1549 7466 1564
rect 7500 1549 7556 1564
rect 7590 1549 7646 1564
rect 7680 1549 7736 1564
rect 7770 1549 7826 1564
rect 7860 1549 7916 1564
rect 7950 1549 8006 1564
rect 6980 1530 7016 1549
rect 7070 1530 7106 1549
rect 7160 1530 7196 1549
rect 7250 1530 7286 1549
rect 7340 1530 7376 1549
rect 7430 1530 7466 1549
rect 7520 1530 7556 1549
rect 7610 1530 7646 1549
rect 7700 1530 7736 1549
rect 7790 1530 7826 1549
rect 7880 1530 7916 1549
rect 7970 1530 8006 1549
rect 8040 1530 8176 1564
rect 8210 1530 8266 1564
rect 8300 1549 8356 1564
rect 8390 1549 8446 1564
rect 8480 1549 8536 1564
rect 8570 1549 8626 1564
rect 8660 1549 8716 1564
rect 8750 1549 8806 1564
rect 8840 1549 8896 1564
rect 8930 1549 8986 1564
rect 9020 1549 9076 1564
rect 9110 1549 9166 1564
rect 9200 1549 9256 1564
rect 9290 1549 9346 1564
rect 8320 1530 8356 1549
rect 8410 1530 8446 1549
rect 8500 1530 8536 1549
rect 8590 1530 8626 1549
rect 8680 1530 8716 1549
rect 8770 1530 8806 1549
rect 8860 1530 8896 1549
rect 8950 1530 8986 1549
rect 9040 1530 9076 1549
rect 9130 1530 9166 1549
rect 9220 1530 9256 1549
rect 9310 1530 9346 1549
rect 9380 1530 9444 1564
rect 116 1526 246 1530
rect 116 1492 150 1526
rect 184 1515 246 1526
rect 280 1515 336 1530
rect 370 1515 426 1530
rect 460 1515 516 1530
rect 550 1515 606 1530
rect 640 1515 696 1530
rect 730 1515 786 1530
rect 820 1515 876 1530
rect 910 1515 966 1530
rect 1000 1515 1056 1530
rect 1090 1515 1146 1530
rect 1180 1515 1236 1530
rect 1270 1526 1586 1530
rect 1270 1515 1337 1526
rect 184 1492 1337 1515
rect 1371 1492 1490 1526
rect 1524 1515 1586 1526
rect 1620 1515 1676 1530
rect 1710 1515 1766 1530
rect 1800 1515 1856 1530
rect 1890 1515 1946 1530
rect 1980 1515 2036 1530
rect 2070 1515 2126 1530
rect 2160 1515 2216 1530
rect 2250 1515 2306 1530
rect 2340 1515 2396 1530
rect 2430 1515 2486 1530
rect 2520 1515 2576 1530
rect 2610 1526 2926 1530
rect 2610 1515 2677 1526
rect 1524 1492 2677 1515
rect 2711 1492 2830 1526
rect 2864 1515 2926 1526
rect 2960 1515 3016 1530
rect 3050 1515 3106 1530
rect 3140 1515 3196 1530
rect 3230 1515 3286 1530
rect 3320 1515 3376 1530
rect 3410 1515 3466 1530
rect 3500 1515 3556 1530
rect 3590 1515 3646 1530
rect 3680 1515 3736 1530
rect 3770 1515 3826 1530
rect 3860 1515 3916 1530
rect 3950 1526 4266 1530
rect 3950 1515 4017 1526
rect 2864 1492 4017 1515
rect 4051 1492 4170 1526
rect 4204 1515 4266 1526
rect 4300 1515 4356 1530
rect 4390 1515 4446 1530
rect 4480 1515 4536 1530
rect 4570 1515 4626 1530
rect 4660 1515 4716 1530
rect 4750 1515 4806 1530
rect 4840 1515 4896 1530
rect 4930 1515 4986 1530
rect 5020 1515 5076 1530
rect 5110 1515 5166 1530
rect 5200 1515 5256 1530
rect 5290 1526 5606 1530
rect 5290 1515 5357 1526
rect 4204 1492 5357 1515
rect 5391 1492 5510 1526
rect 5544 1515 5606 1526
rect 5640 1515 5696 1530
rect 5730 1515 5786 1530
rect 5820 1515 5876 1530
rect 5910 1515 5966 1530
rect 6000 1515 6056 1530
rect 6090 1515 6146 1530
rect 6180 1515 6236 1530
rect 6270 1515 6326 1530
rect 6360 1515 6416 1530
rect 6450 1515 6506 1530
rect 6540 1515 6596 1530
rect 6630 1526 6946 1530
rect 6630 1515 6697 1526
rect 5544 1492 6697 1515
rect 6731 1492 6850 1526
rect 6884 1515 6946 1526
rect 6980 1515 7036 1530
rect 7070 1515 7126 1530
rect 7160 1515 7216 1530
rect 7250 1515 7306 1530
rect 7340 1515 7396 1530
rect 7430 1515 7486 1530
rect 7520 1515 7576 1530
rect 7610 1515 7666 1530
rect 7700 1515 7756 1530
rect 7790 1515 7846 1530
rect 7880 1515 7936 1530
rect 7970 1526 8286 1530
rect 7970 1515 8037 1526
rect 6884 1492 8037 1515
rect 8071 1492 8190 1526
rect 8224 1515 8286 1526
rect 8320 1515 8376 1530
rect 8410 1515 8466 1530
rect 8500 1515 8556 1530
rect 8590 1515 8646 1530
rect 8680 1515 8736 1530
rect 8770 1515 8826 1530
rect 8860 1515 8916 1530
rect 8950 1515 9006 1530
rect 9040 1515 9096 1530
rect 9130 1515 9186 1530
rect 9220 1515 9276 1530
rect 9310 1526 9444 1530
rect 9310 1515 9377 1526
rect 8224 1492 9377 1515
rect 9411 1492 9444 1526
rect 116 1485 9444 1492
rect 116 1436 215 1485
rect 116 1402 150 1436
rect 184 1402 215 1436
rect 1305 1436 1555 1485
rect 116 1346 215 1402
rect 116 1312 150 1346
rect 184 1312 215 1346
rect 116 1256 215 1312
rect 116 1222 150 1256
rect 184 1222 215 1256
rect 116 1166 215 1222
rect 116 1132 150 1166
rect 184 1132 215 1166
rect 116 1076 215 1132
rect 116 1042 150 1076
rect 184 1042 215 1076
rect 116 986 215 1042
rect 116 952 150 986
rect 184 952 215 986
rect 116 896 215 952
rect 116 862 150 896
rect 184 862 215 896
rect 116 806 215 862
rect 116 772 150 806
rect 184 772 215 806
rect 116 716 215 772
rect 116 682 150 716
rect 184 682 215 716
rect 116 626 215 682
rect 116 592 150 626
rect 184 592 215 626
rect 116 536 215 592
rect 116 502 150 536
rect 184 502 215 536
rect 116 446 215 502
rect 279 1404 1241 1421
rect 279 1370 300 1404
rect 334 1370 390 1404
rect 424 1402 480 1404
rect 514 1402 570 1404
rect 604 1402 660 1404
rect 694 1402 750 1404
rect 784 1402 840 1404
rect 874 1402 930 1404
rect 964 1402 1020 1404
rect 1054 1402 1110 1404
rect 1144 1402 1200 1404
rect 444 1370 480 1402
rect 534 1370 570 1402
rect 624 1370 660 1402
rect 714 1370 750 1402
rect 804 1370 840 1402
rect 894 1370 930 1402
rect 984 1370 1020 1402
rect 1074 1370 1110 1402
rect 1164 1370 1200 1402
rect 1234 1370 1241 1404
rect 279 1368 410 1370
rect 444 1368 500 1370
rect 534 1368 590 1370
rect 624 1368 680 1370
rect 714 1368 770 1370
rect 804 1368 860 1370
rect 894 1368 950 1370
rect 984 1368 1040 1370
rect 1074 1368 1130 1370
rect 1164 1368 1241 1370
rect 279 1349 1241 1368
rect 279 1345 351 1349
rect 279 1311 298 1345
rect 332 1311 351 1345
rect 279 1255 351 1311
rect 1169 1326 1241 1349
rect 1169 1292 1188 1326
rect 1222 1292 1241 1326
rect 279 1221 298 1255
rect 332 1221 351 1255
rect 279 1165 351 1221
rect 279 1131 298 1165
rect 332 1131 351 1165
rect 279 1075 351 1131
rect 279 1041 298 1075
rect 332 1041 351 1075
rect 279 985 351 1041
rect 279 951 298 985
rect 332 951 351 985
rect 279 895 351 951
rect 279 861 298 895
rect 332 861 351 895
rect 279 805 351 861
rect 279 771 298 805
rect 332 771 351 805
rect 279 715 351 771
rect 279 681 298 715
rect 332 681 351 715
rect 279 625 351 681
rect 279 591 298 625
rect 332 591 351 625
rect 413 1228 1107 1287
rect 413 1194 474 1228
rect 508 1200 564 1228
rect 598 1200 654 1228
rect 688 1200 744 1228
rect 520 1194 564 1200
rect 620 1194 654 1200
rect 720 1194 744 1200
rect 778 1200 834 1228
rect 778 1194 786 1200
rect 413 1166 486 1194
rect 520 1166 586 1194
rect 620 1166 686 1194
rect 720 1166 786 1194
rect 820 1194 834 1200
rect 868 1200 924 1228
rect 868 1194 886 1200
rect 820 1166 886 1194
rect 920 1194 924 1200
rect 958 1200 1014 1228
rect 958 1194 986 1200
rect 1048 1194 1107 1228
rect 920 1166 986 1194
rect 1020 1166 1107 1194
rect 413 1138 1107 1166
rect 413 1104 474 1138
rect 508 1104 564 1138
rect 598 1104 654 1138
rect 688 1104 744 1138
rect 778 1104 834 1138
rect 868 1104 924 1138
rect 958 1104 1014 1138
rect 1048 1104 1107 1138
rect 413 1100 1107 1104
rect 413 1066 486 1100
rect 520 1066 586 1100
rect 620 1066 686 1100
rect 720 1066 786 1100
rect 820 1066 886 1100
rect 920 1066 986 1100
rect 1020 1066 1107 1100
rect 413 1048 1107 1066
rect 413 1014 474 1048
rect 508 1014 564 1048
rect 598 1014 654 1048
rect 688 1014 744 1048
rect 778 1014 834 1048
rect 868 1014 924 1048
rect 958 1014 1014 1048
rect 1048 1014 1107 1048
rect 413 1000 1107 1014
rect 413 966 486 1000
rect 520 966 586 1000
rect 620 966 686 1000
rect 720 966 786 1000
rect 820 966 886 1000
rect 920 966 986 1000
rect 1020 966 1107 1000
rect 413 958 1107 966
rect 413 924 474 958
rect 508 924 564 958
rect 598 924 654 958
rect 688 924 744 958
rect 778 924 834 958
rect 868 924 924 958
rect 958 924 1014 958
rect 1048 924 1107 958
rect 413 900 1107 924
rect 413 868 486 900
rect 520 868 586 900
rect 620 868 686 900
rect 720 868 786 900
rect 413 834 474 868
rect 520 866 564 868
rect 620 866 654 868
rect 720 866 744 868
rect 508 834 564 866
rect 598 834 654 866
rect 688 834 744 866
rect 778 866 786 868
rect 820 868 886 900
rect 820 866 834 868
rect 778 834 834 866
rect 868 866 886 868
rect 920 868 986 900
rect 1020 868 1107 900
rect 920 866 924 868
rect 868 834 924 866
rect 958 866 986 868
rect 958 834 1014 866
rect 1048 834 1107 868
rect 413 800 1107 834
rect 413 778 486 800
rect 520 778 586 800
rect 620 778 686 800
rect 720 778 786 800
rect 413 744 474 778
rect 520 766 564 778
rect 620 766 654 778
rect 720 766 744 778
rect 508 744 564 766
rect 598 744 654 766
rect 688 744 744 766
rect 778 766 786 778
rect 820 778 886 800
rect 820 766 834 778
rect 778 744 834 766
rect 868 766 886 778
rect 920 778 986 800
rect 1020 778 1107 800
rect 920 766 924 778
rect 868 744 924 766
rect 958 766 986 778
rect 958 744 1014 766
rect 1048 744 1107 778
rect 413 700 1107 744
rect 413 688 486 700
rect 520 688 586 700
rect 620 688 686 700
rect 720 688 786 700
rect 413 654 474 688
rect 520 666 564 688
rect 620 666 654 688
rect 720 666 744 688
rect 508 654 564 666
rect 598 654 654 666
rect 688 654 744 666
rect 778 666 786 688
rect 820 688 886 700
rect 820 666 834 688
rect 778 654 834 666
rect 868 666 886 688
rect 920 688 986 700
rect 1020 688 1107 700
rect 920 666 924 688
rect 868 654 924 666
rect 958 666 986 688
rect 958 654 1014 666
rect 1048 654 1107 688
rect 413 593 1107 654
rect 1169 1236 1241 1292
rect 1169 1202 1188 1236
rect 1222 1202 1241 1236
rect 1169 1146 1241 1202
rect 1169 1112 1188 1146
rect 1222 1112 1241 1146
rect 1169 1056 1241 1112
rect 1169 1022 1188 1056
rect 1222 1022 1241 1056
rect 1169 966 1241 1022
rect 1169 932 1188 966
rect 1222 932 1241 966
rect 1169 876 1241 932
rect 1169 842 1188 876
rect 1222 842 1241 876
rect 1169 786 1241 842
rect 1169 752 1188 786
rect 1222 752 1241 786
rect 1169 696 1241 752
rect 1169 662 1188 696
rect 1222 662 1241 696
rect 1169 606 1241 662
rect 279 531 351 591
rect 1169 572 1188 606
rect 1222 572 1241 606
rect 1169 531 1241 572
rect 279 512 1241 531
rect 279 478 376 512
rect 410 478 466 512
rect 500 478 556 512
rect 590 478 646 512
rect 680 478 736 512
rect 770 478 826 512
rect 860 478 916 512
rect 950 478 1006 512
rect 1040 478 1096 512
rect 1130 478 1241 512
rect 279 459 1241 478
rect 1305 1402 1337 1436
rect 1371 1402 1490 1436
rect 1524 1402 1555 1436
rect 2645 1436 2895 1485
rect 1305 1346 1555 1402
rect 1305 1312 1337 1346
rect 1371 1312 1490 1346
rect 1524 1312 1555 1346
rect 1305 1256 1555 1312
rect 1305 1222 1337 1256
rect 1371 1222 1490 1256
rect 1524 1222 1555 1256
rect 1305 1166 1555 1222
rect 1305 1132 1337 1166
rect 1371 1132 1490 1166
rect 1524 1132 1555 1166
rect 1305 1076 1555 1132
rect 1305 1042 1337 1076
rect 1371 1042 1490 1076
rect 1524 1042 1555 1076
rect 1305 986 1555 1042
rect 1305 952 1337 986
rect 1371 952 1490 986
rect 1524 952 1555 986
rect 1305 896 1555 952
rect 1305 862 1337 896
rect 1371 862 1490 896
rect 1524 862 1555 896
rect 1305 806 1555 862
rect 1305 772 1337 806
rect 1371 772 1490 806
rect 1524 772 1555 806
rect 1305 716 1555 772
rect 1305 682 1337 716
rect 1371 682 1490 716
rect 1524 682 1555 716
rect 1305 626 1555 682
rect 1305 592 1337 626
rect 1371 592 1490 626
rect 1524 592 1555 626
rect 1305 536 1555 592
rect 1305 502 1337 536
rect 1371 502 1490 536
rect 1524 502 1555 536
rect 116 412 150 446
rect 184 412 215 446
rect 116 395 215 412
rect 1305 446 1555 502
rect 1619 1404 2581 1421
rect 1619 1370 1640 1404
rect 1674 1370 1730 1404
rect 1764 1402 1820 1404
rect 1854 1402 1910 1404
rect 1944 1402 2000 1404
rect 2034 1402 2090 1404
rect 2124 1402 2180 1404
rect 2214 1402 2270 1404
rect 2304 1402 2360 1404
rect 2394 1402 2450 1404
rect 2484 1402 2540 1404
rect 1784 1370 1820 1402
rect 1874 1370 1910 1402
rect 1964 1370 2000 1402
rect 2054 1370 2090 1402
rect 2144 1370 2180 1402
rect 2234 1370 2270 1402
rect 2324 1370 2360 1402
rect 2414 1370 2450 1402
rect 2504 1370 2540 1402
rect 2574 1370 2581 1404
rect 1619 1368 1750 1370
rect 1784 1368 1840 1370
rect 1874 1368 1930 1370
rect 1964 1368 2020 1370
rect 2054 1368 2110 1370
rect 2144 1368 2200 1370
rect 2234 1368 2290 1370
rect 2324 1368 2380 1370
rect 2414 1368 2470 1370
rect 2504 1368 2581 1370
rect 1619 1349 2581 1368
rect 1619 1345 1691 1349
rect 1619 1311 1638 1345
rect 1672 1311 1691 1345
rect 1619 1255 1691 1311
rect 2509 1326 2581 1349
rect 2509 1292 2528 1326
rect 2562 1292 2581 1326
rect 1619 1221 1638 1255
rect 1672 1221 1691 1255
rect 1619 1165 1691 1221
rect 1619 1131 1638 1165
rect 1672 1131 1691 1165
rect 1619 1075 1691 1131
rect 1619 1041 1638 1075
rect 1672 1041 1691 1075
rect 1619 985 1691 1041
rect 1619 951 1638 985
rect 1672 951 1691 985
rect 1619 895 1691 951
rect 1619 861 1638 895
rect 1672 861 1691 895
rect 1619 805 1691 861
rect 1619 771 1638 805
rect 1672 771 1691 805
rect 1619 715 1691 771
rect 1619 681 1638 715
rect 1672 681 1691 715
rect 1619 625 1691 681
rect 1619 591 1638 625
rect 1672 591 1691 625
rect 1753 1228 2447 1287
rect 1753 1194 1814 1228
rect 1848 1200 1904 1228
rect 1938 1200 1994 1228
rect 2028 1200 2084 1228
rect 1860 1194 1904 1200
rect 1960 1194 1994 1200
rect 2060 1194 2084 1200
rect 2118 1200 2174 1228
rect 2118 1194 2126 1200
rect 1753 1166 1826 1194
rect 1860 1166 1926 1194
rect 1960 1166 2026 1194
rect 2060 1166 2126 1194
rect 2160 1194 2174 1200
rect 2208 1200 2264 1228
rect 2208 1194 2226 1200
rect 2160 1166 2226 1194
rect 2260 1194 2264 1200
rect 2298 1200 2354 1228
rect 2298 1194 2326 1200
rect 2388 1194 2447 1228
rect 2260 1166 2326 1194
rect 2360 1166 2447 1194
rect 1753 1138 2447 1166
rect 1753 1104 1814 1138
rect 1848 1104 1904 1138
rect 1938 1104 1994 1138
rect 2028 1104 2084 1138
rect 2118 1104 2174 1138
rect 2208 1104 2264 1138
rect 2298 1104 2354 1138
rect 2388 1104 2447 1138
rect 1753 1100 2447 1104
rect 1753 1066 1826 1100
rect 1860 1066 1926 1100
rect 1960 1066 2026 1100
rect 2060 1066 2126 1100
rect 2160 1066 2226 1100
rect 2260 1066 2326 1100
rect 2360 1066 2447 1100
rect 1753 1048 2447 1066
rect 1753 1014 1814 1048
rect 1848 1014 1904 1048
rect 1938 1014 1994 1048
rect 2028 1014 2084 1048
rect 2118 1014 2174 1048
rect 2208 1014 2264 1048
rect 2298 1014 2354 1048
rect 2388 1014 2447 1048
rect 1753 1000 2447 1014
rect 1753 966 1826 1000
rect 1860 966 1926 1000
rect 1960 966 2026 1000
rect 2060 966 2126 1000
rect 2160 966 2226 1000
rect 2260 966 2326 1000
rect 2360 966 2447 1000
rect 1753 958 2447 966
rect 1753 924 1814 958
rect 1848 924 1904 958
rect 1938 924 1994 958
rect 2028 924 2084 958
rect 2118 924 2174 958
rect 2208 924 2264 958
rect 2298 924 2354 958
rect 2388 924 2447 958
rect 1753 900 2447 924
rect 1753 868 1826 900
rect 1860 868 1926 900
rect 1960 868 2026 900
rect 2060 868 2126 900
rect 1753 834 1814 868
rect 1860 866 1904 868
rect 1960 866 1994 868
rect 2060 866 2084 868
rect 1848 834 1904 866
rect 1938 834 1994 866
rect 2028 834 2084 866
rect 2118 866 2126 868
rect 2160 868 2226 900
rect 2160 866 2174 868
rect 2118 834 2174 866
rect 2208 866 2226 868
rect 2260 868 2326 900
rect 2360 868 2447 900
rect 2260 866 2264 868
rect 2208 834 2264 866
rect 2298 866 2326 868
rect 2298 834 2354 866
rect 2388 834 2447 868
rect 1753 800 2447 834
rect 1753 778 1826 800
rect 1860 778 1926 800
rect 1960 778 2026 800
rect 2060 778 2126 800
rect 1753 744 1814 778
rect 1860 766 1904 778
rect 1960 766 1994 778
rect 2060 766 2084 778
rect 1848 744 1904 766
rect 1938 744 1994 766
rect 2028 744 2084 766
rect 2118 766 2126 778
rect 2160 778 2226 800
rect 2160 766 2174 778
rect 2118 744 2174 766
rect 2208 766 2226 778
rect 2260 778 2326 800
rect 2360 778 2447 800
rect 2260 766 2264 778
rect 2208 744 2264 766
rect 2298 766 2326 778
rect 2298 744 2354 766
rect 2388 744 2447 778
rect 1753 700 2447 744
rect 1753 688 1826 700
rect 1860 688 1926 700
rect 1960 688 2026 700
rect 2060 688 2126 700
rect 1753 654 1814 688
rect 1860 666 1904 688
rect 1960 666 1994 688
rect 2060 666 2084 688
rect 1848 654 1904 666
rect 1938 654 1994 666
rect 2028 654 2084 666
rect 2118 666 2126 688
rect 2160 688 2226 700
rect 2160 666 2174 688
rect 2118 654 2174 666
rect 2208 666 2226 688
rect 2260 688 2326 700
rect 2360 688 2447 700
rect 2260 666 2264 688
rect 2208 654 2264 666
rect 2298 666 2326 688
rect 2298 654 2354 666
rect 2388 654 2447 688
rect 1753 593 2447 654
rect 2509 1236 2581 1292
rect 2509 1202 2528 1236
rect 2562 1202 2581 1236
rect 2509 1146 2581 1202
rect 2509 1112 2528 1146
rect 2562 1112 2581 1146
rect 2509 1056 2581 1112
rect 2509 1022 2528 1056
rect 2562 1022 2581 1056
rect 2509 966 2581 1022
rect 2509 932 2528 966
rect 2562 932 2581 966
rect 2509 876 2581 932
rect 2509 842 2528 876
rect 2562 842 2581 876
rect 2509 786 2581 842
rect 2509 752 2528 786
rect 2562 752 2581 786
rect 2509 696 2581 752
rect 2509 662 2528 696
rect 2562 662 2581 696
rect 2509 606 2581 662
rect 1619 531 1691 591
rect 2509 572 2528 606
rect 2562 572 2581 606
rect 2509 531 2581 572
rect 1619 512 2581 531
rect 1619 478 1716 512
rect 1750 478 1806 512
rect 1840 478 1896 512
rect 1930 478 1986 512
rect 2020 478 2076 512
rect 2110 478 2166 512
rect 2200 478 2256 512
rect 2290 478 2346 512
rect 2380 478 2436 512
rect 2470 478 2581 512
rect 1619 459 2581 478
rect 2645 1402 2677 1436
rect 2711 1402 2830 1436
rect 2864 1402 2895 1436
rect 3985 1436 4235 1485
rect 2645 1346 2895 1402
rect 2645 1312 2677 1346
rect 2711 1312 2830 1346
rect 2864 1312 2895 1346
rect 2645 1256 2895 1312
rect 2645 1222 2677 1256
rect 2711 1222 2830 1256
rect 2864 1222 2895 1256
rect 2645 1166 2895 1222
rect 2645 1132 2677 1166
rect 2711 1132 2830 1166
rect 2864 1132 2895 1166
rect 2645 1076 2895 1132
rect 2645 1042 2677 1076
rect 2711 1042 2830 1076
rect 2864 1042 2895 1076
rect 2645 986 2895 1042
rect 2645 952 2677 986
rect 2711 952 2830 986
rect 2864 952 2895 986
rect 2645 896 2895 952
rect 2645 862 2677 896
rect 2711 862 2830 896
rect 2864 862 2895 896
rect 2645 806 2895 862
rect 2645 772 2677 806
rect 2711 772 2830 806
rect 2864 772 2895 806
rect 2645 716 2895 772
rect 2645 682 2677 716
rect 2711 682 2830 716
rect 2864 682 2895 716
rect 2645 626 2895 682
rect 2645 592 2677 626
rect 2711 592 2830 626
rect 2864 592 2895 626
rect 2645 536 2895 592
rect 2645 502 2677 536
rect 2711 502 2830 536
rect 2864 502 2895 536
rect 1305 412 1337 446
rect 1371 412 1490 446
rect 1524 412 1555 446
rect 1305 395 1555 412
rect 2645 446 2895 502
rect 2959 1404 3921 1421
rect 2959 1370 2980 1404
rect 3014 1370 3070 1404
rect 3104 1402 3160 1404
rect 3194 1402 3250 1404
rect 3284 1402 3340 1404
rect 3374 1402 3430 1404
rect 3464 1402 3520 1404
rect 3554 1402 3610 1404
rect 3644 1402 3700 1404
rect 3734 1402 3790 1404
rect 3824 1402 3880 1404
rect 3124 1370 3160 1402
rect 3214 1370 3250 1402
rect 3304 1370 3340 1402
rect 3394 1370 3430 1402
rect 3484 1370 3520 1402
rect 3574 1370 3610 1402
rect 3664 1370 3700 1402
rect 3754 1370 3790 1402
rect 3844 1370 3880 1402
rect 3914 1370 3921 1404
rect 2959 1368 3090 1370
rect 3124 1368 3180 1370
rect 3214 1368 3270 1370
rect 3304 1368 3360 1370
rect 3394 1368 3450 1370
rect 3484 1368 3540 1370
rect 3574 1368 3630 1370
rect 3664 1368 3720 1370
rect 3754 1368 3810 1370
rect 3844 1368 3921 1370
rect 2959 1349 3921 1368
rect 2959 1345 3031 1349
rect 2959 1311 2978 1345
rect 3012 1311 3031 1345
rect 2959 1255 3031 1311
rect 3849 1326 3921 1349
rect 3849 1292 3868 1326
rect 3902 1292 3921 1326
rect 2959 1221 2978 1255
rect 3012 1221 3031 1255
rect 2959 1165 3031 1221
rect 2959 1131 2978 1165
rect 3012 1131 3031 1165
rect 2959 1075 3031 1131
rect 2959 1041 2978 1075
rect 3012 1041 3031 1075
rect 2959 985 3031 1041
rect 2959 951 2978 985
rect 3012 951 3031 985
rect 2959 895 3031 951
rect 2959 861 2978 895
rect 3012 861 3031 895
rect 2959 805 3031 861
rect 2959 771 2978 805
rect 3012 771 3031 805
rect 2959 715 3031 771
rect 2959 681 2978 715
rect 3012 681 3031 715
rect 2959 625 3031 681
rect 2959 591 2978 625
rect 3012 591 3031 625
rect 3093 1228 3787 1287
rect 3093 1194 3154 1228
rect 3188 1200 3244 1228
rect 3278 1200 3334 1228
rect 3368 1200 3424 1228
rect 3200 1194 3244 1200
rect 3300 1194 3334 1200
rect 3400 1194 3424 1200
rect 3458 1200 3514 1228
rect 3458 1194 3466 1200
rect 3093 1166 3166 1194
rect 3200 1166 3266 1194
rect 3300 1166 3366 1194
rect 3400 1166 3466 1194
rect 3500 1194 3514 1200
rect 3548 1200 3604 1228
rect 3548 1194 3566 1200
rect 3500 1166 3566 1194
rect 3600 1194 3604 1200
rect 3638 1200 3694 1228
rect 3638 1194 3666 1200
rect 3728 1194 3787 1228
rect 3600 1166 3666 1194
rect 3700 1166 3787 1194
rect 3093 1138 3787 1166
rect 3093 1104 3154 1138
rect 3188 1104 3244 1138
rect 3278 1104 3334 1138
rect 3368 1104 3424 1138
rect 3458 1104 3514 1138
rect 3548 1104 3604 1138
rect 3638 1104 3694 1138
rect 3728 1104 3787 1138
rect 3093 1100 3787 1104
rect 3093 1066 3166 1100
rect 3200 1066 3266 1100
rect 3300 1066 3366 1100
rect 3400 1066 3466 1100
rect 3500 1066 3566 1100
rect 3600 1066 3666 1100
rect 3700 1066 3787 1100
rect 3093 1048 3787 1066
rect 3093 1014 3154 1048
rect 3188 1014 3244 1048
rect 3278 1014 3334 1048
rect 3368 1014 3424 1048
rect 3458 1014 3514 1048
rect 3548 1014 3604 1048
rect 3638 1014 3694 1048
rect 3728 1014 3787 1048
rect 3093 1000 3787 1014
rect 3093 966 3166 1000
rect 3200 966 3266 1000
rect 3300 966 3366 1000
rect 3400 966 3466 1000
rect 3500 966 3566 1000
rect 3600 966 3666 1000
rect 3700 966 3787 1000
rect 3093 958 3787 966
rect 3093 924 3154 958
rect 3188 924 3244 958
rect 3278 924 3334 958
rect 3368 924 3424 958
rect 3458 924 3514 958
rect 3548 924 3604 958
rect 3638 924 3694 958
rect 3728 924 3787 958
rect 3093 900 3787 924
rect 3093 868 3166 900
rect 3200 868 3266 900
rect 3300 868 3366 900
rect 3400 868 3466 900
rect 3093 834 3154 868
rect 3200 866 3244 868
rect 3300 866 3334 868
rect 3400 866 3424 868
rect 3188 834 3244 866
rect 3278 834 3334 866
rect 3368 834 3424 866
rect 3458 866 3466 868
rect 3500 868 3566 900
rect 3500 866 3514 868
rect 3458 834 3514 866
rect 3548 866 3566 868
rect 3600 868 3666 900
rect 3700 868 3787 900
rect 3600 866 3604 868
rect 3548 834 3604 866
rect 3638 866 3666 868
rect 3638 834 3694 866
rect 3728 834 3787 868
rect 3093 800 3787 834
rect 3093 778 3166 800
rect 3200 778 3266 800
rect 3300 778 3366 800
rect 3400 778 3466 800
rect 3093 744 3154 778
rect 3200 766 3244 778
rect 3300 766 3334 778
rect 3400 766 3424 778
rect 3188 744 3244 766
rect 3278 744 3334 766
rect 3368 744 3424 766
rect 3458 766 3466 778
rect 3500 778 3566 800
rect 3500 766 3514 778
rect 3458 744 3514 766
rect 3548 766 3566 778
rect 3600 778 3666 800
rect 3700 778 3787 800
rect 3600 766 3604 778
rect 3548 744 3604 766
rect 3638 766 3666 778
rect 3638 744 3694 766
rect 3728 744 3787 778
rect 3093 700 3787 744
rect 3093 688 3166 700
rect 3200 688 3266 700
rect 3300 688 3366 700
rect 3400 688 3466 700
rect 3093 654 3154 688
rect 3200 666 3244 688
rect 3300 666 3334 688
rect 3400 666 3424 688
rect 3188 654 3244 666
rect 3278 654 3334 666
rect 3368 654 3424 666
rect 3458 666 3466 688
rect 3500 688 3566 700
rect 3500 666 3514 688
rect 3458 654 3514 666
rect 3548 666 3566 688
rect 3600 688 3666 700
rect 3700 688 3787 700
rect 3600 666 3604 688
rect 3548 654 3604 666
rect 3638 666 3666 688
rect 3638 654 3694 666
rect 3728 654 3787 688
rect 3093 593 3787 654
rect 3849 1236 3921 1292
rect 3849 1202 3868 1236
rect 3902 1202 3921 1236
rect 3849 1146 3921 1202
rect 3849 1112 3868 1146
rect 3902 1112 3921 1146
rect 3849 1056 3921 1112
rect 3849 1022 3868 1056
rect 3902 1022 3921 1056
rect 3849 966 3921 1022
rect 3849 932 3868 966
rect 3902 932 3921 966
rect 3849 876 3921 932
rect 3849 842 3868 876
rect 3902 842 3921 876
rect 3849 786 3921 842
rect 3849 752 3868 786
rect 3902 752 3921 786
rect 3849 696 3921 752
rect 3849 662 3868 696
rect 3902 662 3921 696
rect 3849 606 3921 662
rect 2959 531 3031 591
rect 3849 572 3868 606
rect 3902 572 3921 606
rect 3849 531 3921 572
rect 2959 512 3921 531
rect 2959 478 3056 512
rect 3090 478 3146 512
rect 3180 478 3236 512
rect 3270 478 3326 512
rect 3360 478 3416 512
rect 3450 478 3506 512
rect 3540 478 3596 512
rect 3630 478 3686 512
rect 3720 478 3776 512
rect 3810 478 3921 512
rect 2959 459 3921 478
rect 3985 1402 4017 1436
rect 4051 1402 4170 1436
rect 4204 1402 4235 1436
rect 5325 1436 5575 1485
rect 3985 1346 4235 1402
rect 3985 1312 4017 1346
rect 4051 1312 4170 1346
rect 4204 1312 4235 1346
rect 3985 1256 4235 1312
rect 3985 1222 4017 1256
rect 4051 1222 4170 1256
rect 4204 1222 4235 1256
rect 3985 1166 4235 1222
rect 3985 1132 4017 1166
rect 4051 1132 4170 1166
rect 4204 1132 4235 1166
rect 3985 1076 4235 1132
rect 3985 1042 4017 1076
rect 4051 1042 4170 1076
rect 4204 1042 4235 1076
rect 3985 986 4235 1042
rect 3985 952 4017 986
rect 4051 952 4170 986
rect 4204 952 4235 986
rect 3985 896 4235 952
rect 3985 862 4017 896
rect 4051 862 4170 896
rect 4204 862 4235 896
rect 3985 806 4235 862
rect 3985 772 4017 806
rect 4051 772 4170 806
rect 4204 772 4235 806
rect 3985 716 4235 772
rect 3985 682 4017 716
rect 4051 682 4170 716
rect 4204 682 4235 716
rect 3985 626 4235 682
rect 3985 592 4017 626
rect 4051 592 4170 626
rect 4204 592 4235 626
rect 3985 536 4235 592
rect 3985 502 4017 536
rect 4051 502 4170 536
rect 4204 502 4235 536
rect 2645 412 2677 446
rect 2711 412 2830 446
rect 2864 412 2895 446
rect 2645 395 2895 412
rect 3985 446 4235 502
rect 4299 1404 5261 1421
rect 4299 1370 4320 1404
rect 4354 1370 4410 1404
rect 4444 1402 4500 1404
rect 4534 1402 4590 1404
rect 4624 1402 4680 1404
rect 4714 1402 4770 1404
rect 4804 1402 4860 1404
rect 4894 1402 4950 1404
rect 4984 1402 5040 1404
rect 5074 1402 5130 1404
rect 5164 1402 5220 1404
rect 4464 1370 4500 1402
rect 4554 1370 4590 1402
rect 4644 1370 4680 1402
rect 4734 1370 4770 1402
rect 4824 1370 4860 1402
rect 4914 1370 4950 1402
rect 5004 1370 5040 1402
rect 5094 1370 5130 1402
rect 5184 1370 5220 1402
rect 5254 1370 5261 1404
rect 4299 1368 4430 1370
rect 4464 1368 4520 1370
rect 4554 1368 4610 1370
rect 4644 1368 4700 1370
rect 4734 1368 4790 1370
rect 4824 1368 4880 1370
rect 4914 1368 4970 1370
rect 5004 1368 5060 1370
rect 5094 1368 5150 1370
rect 5184 1368 5261 1370
rect 4299 1349 5261 1368
rect 4299 1345 4371 1349
rect 4299 1311 4318 1345
rect 4352 1311 4371 1345
rect 4299 1255 4371 1311
rect 5189 1326 5261 1349
rect 5189 1292 5208 1326
rect 5242 1292 5261 1326
rect 4299 1221 4318 1255
rect 4352 1221 4371 1255
rect 4299 1165 4371 1221
rect 4299 1131 4318 1165
rect 4352 1131 4371 1165
rect 4299 1075 4371 1131
rect 4299 1041 4318 1075
rect 4352 1041 4371 1075
rect 4299 985 4371 1041
rect 4299 951 4318 985
rect 4352 951 4371 985
rect 4299 895 4371 951
rect 4299 861 4318 895
rect 4352 861 4371 895
rect 4299 805 4371 861
rect 4299 771 4318 805
rect 4352 771 4371 805
rect 4299 715 4371 771
rect 4299 681 4318 715
rect 4352 681 4371 715
rect 4299 625 4371 681
rect 4299 591 4318 625
rect 4352 591 4371 625
rect 4433 1228 5127 1287
rect 4433 1194 4494 1228
rect 4528 1200 4584 1228
rect 4618 1200 4674 1228
rect 4708 1200 4764 1228
rect 4540 1194 4584 1200
rect 4640 1194 4674 1200
rect 4740 1194 4764 1200
rect 4798 1200 4854 1228
rect 4798 1194 4806 1200
rect 4433 1166 4506 1194
rect 4540 1166 4606 1194
rect 4640 1166 4706 1194
rect 4740 1166 4806 1194
rect 4840 1194 4854 1200
rect 4888 1200 4944 1228
rect 4888 1194 4906 1200
rect 4840 1166 4906 1194
rect 4940 1194 4944 1200
rect 4978 1200 5034 1228
rect 4978 1194 5006 1200
rect 5068 1194 5127 1228
rect 4940 1166 5006 1194
rect 5040 1166 5127 1194
rect 4433 1138 5127 1166
rect 4433 1104 4494 1138
rect 4528 1104 4584 1138
rect 4618 1104 4674 1138
rect 4708 1104 4764 1138
rect 4798 1104 4854 1138
rect 4888 1104 4944 1138
rect 4978 1104 5034 1138
rect 5068 1104 5127 1138
rect 4433 1100 5127 1104
rect 4433 1066 4506 1100
rect 4540 1066 4606 1100
rect 4640 1066 4706 1100
rect 4740 1066 4806 1100
rect 4840 1066 4906 1100
rect 4940 1066 5006 1100
rect 5040 1066 5127 1100
rect 4433 1048 5127 1066
rect 4433 1014 4494 1048
rect 4528 1014 4584 1048
rect 4618 1014 4674 1048
rect 4708 1014 4764 1048
rect 4798 1014 4854 1048
rect 4888 1014 4944 1048
rect 4978 1014 5034 1048
rect 5068 1014 5127 1048
rect 4433 1000 5127 1014
rect 4433 966 4506 1000
rect 4540 966 4606 1000
rect 4640 966 4706 1000
rect 4740 966 4806 1000
rect 4840 966 4906 1000
rect 4940 966 5006 1000
rect 5040 966 5127 1000
rect 4433 958 5127 966
rect 4433 924 4494 958
rect 4528 924 4584 958
rect 4618 924 4674 958
rect 4708 924 4764 958
rect 4798 924 4854 958
rect 4888 924 4944 958
rect 4978 924 5034 958
rect 5068 924 5127 958
rect 4433 900 5127 924
rect 4433 868 4506 900
rect 4540 868 4606 900
rect 4640 868 4706 900
rect 4740 868 4806 900
rect 4433 834 4494 868
rect 4540 866 4584 868
rect 4640 866 4674 868
rect 4740 866 4764 868
rect 4528 834 4584 866
rect 4618 834 4674 866
rect 4708 834 4764 866
rect 4798 866 4806 868
rect 4840 868 4906 900
rect 4840 866 4854 868
rect 4798 834 4854 866
rect 4888 866 4906 868
rect 4940 868 5006 900
rect 5040 868 5127 900
rect 4940 866 4944 868
rect 4888 834 4944 866
rect 4978 866 5006 868
rect 4978 834 5034 866
rect 5068 834 5127 868
rect 4433 800 5127 834
rect 4433 778 4506 800
rect 4540 778 4606 800
rect 4640 778 4706 800
rect 4740 778 4806 800
rect 4433 744 4494 778
rect 4540 766 4584 778
rect 4640 766 4674 778
rect 4740 766 4764 778
rect 4528 744 4584 766
rect 4618 744 4674 766
rect 4708 744 4764 766
rect 4798 766 4806 778
rect 4840 778 4906 800
rect 4840 766 4854 778
rect 4798 744 4854 766
rect 4888 766 4906 778
rect 4940 778 5006 800
rect 5040 778 5127 800
rect 4940 766 4944 778
rect 4888 744 4944 766
rect 4978 766 5006 778
rect 4978 744 5034 766
rect 5068 744 5127 778
rect 4433 700 5127 744
rect 4433 688 4506 700
rect 4540 688 4606 700
rect 4640 688 4706 700
rect 4740 688 4806 700
rect 4433 654 4494 688
rect 4540 666 4584 688
rect 4640 666 4674 688
rect 4740 666 4764 688
rect 4528 654 4584 666
rect 4618 654 4674 666
rect 4708 654 4764 666
rect 4798 666 4806 688
rect 4840 688 4906 700
rect 4840 666 4854 688
rect 4798 654 4854 666
rect 4888 666 4906 688
rect 4940 688 5006 700
rect 5040 688 5127 700
rect 4940 666 4944 688
rect 4888 654 4944 666
rect 4978 666 5006 688
rect 4978 654 5034 666
rect 5068 654 5127 688
rect 4433 593 5127 654
rect 5189 1236 5261 1292
rect 5189 1202 5208 1236
rect 5242 1202 5261 1236
rect 5189 1146 5261 1202
rect 5189 1112 5208 1146
rect 5242 1112 5261 1146
rect 5189 1056 5261 1112
rect 5189 1022 5208 1056
rect 5242 1022 5261 1056
rect 5189 966 5261 1022
rect 5189 932 5208 966
rect 5242 932 5261 966
rect 5189 876 5261 932
rect 5189 842 5208 876
rect 5242 842 5261 876
rect 5189 786 5261 842
rect 5189 752 5208 786
rect 5242 752 5261 786
rect 5189 696 5261 752
rect 5189 662 5208 696
rect 5242 662 5261 696
rect 5189 606 5261 662
rect 4299 531 4371 591
rect 5189 572 5208 606
rect 5242 572 5261 606
rect 5189 531 5261 572
rect 4299 512 5261 531
rect 4299 478 4396 512
rect 4430 478 4486 512
rect 4520 478 4576 512
rect 4610 478 4666 512
rect 4700 478 4756 512
rect 4790 478 4846 512
rect 4880 478 4936 512
rect 4970 478 5026 512
rect 5060 478 5116 512
rect 5150 478 5261 512
rect 4299 459 5261 478
rect 5325 1402 5357 1436
rect 5391 1402 5510 1436
rect 5544 1402 5575 1436
rect 6665 1436 6915 1485
rect 5325 1346 5575 1402
rect 5325 1312 5357 1346
rect 5391 1312 5510 1346
rect 5544 1312 5575 1346
rect 5325 1256 5575 1312
rect 5325 1222 5357 1256
rect 5391 1222 5510 1256
rect 5544 1222 5575 1256
rect 5325 1166 5575 1222
rect 5325 1132 5357 1166
rect 5391 1132 5510 1166
rect 5544 1132 5575 1166
rect 5325 1076 5575 1132
rect 5325 1042 5357 1076
rect 5391 1042 5510 1076
rect 5544 1042 5575 1076
rect 5325 986 5575 1042
rect 5325 952 5357 986
rect 5391 952 5510 986
rect 5544 952 5575 986
rect 5325 896 5575 952
rect 5325 862 5357 896
rect 5391 862 5510 896
rect 5544 862 5575 896
rect 5325 806 5575 862
rect 5325 772 5357 806
rect 5391 772 5510 806
rect 5544 772 5575 806
rect 5325 716 5575 772
rect 5325 682 5357 716
rect 5391 682 5510 716
rect 5544 682 5575 716
rect 5325 626 5575 682
rect 5325 592 5357 626
rect 5391 592 5510 626
rect 5544 592 5575 626
rect 5325 536 5575 592
rect 5325 502 5357 536
rect 5391 502 5510 536
rect 5544 502 5575 536
rect 3985 412 4017 446
rect 4051 412 4170 446
rect 4204 412 4235 446
rect 3985 395 4235 412
rect 5325 446 5575 502
rect 5639 1404 6601 1421
rect 5639 1370 5660 1404
rect 5694 1370 5750 1404
rect 5784 1402 5840 1404
rect 5874 1402 5930 1404
rect 5964 1402 6020 1404
rect 6054 1402 6110 1404
rect 6144 1402 6200 1404
rect 6234 1402 6290 1404
rect 6324 1402 6380 1404
rect 6414 1402 6470 1404
rect 6504 1402 6560 1404
rect 5804 1370 5840 1402
rect 5894 1370 5930 1402
rect 5984 1370 6020 1402
rect 6074 1370 6110 1402
rect 6164 1370 6200 1402
rect 6254 1370 6290 1402
rect 6344 1370 6380 1402
rect 6434 1370 6470 1402
rect 6524 1370 6560 1402
rect 6594 1370 6601 1404
rect 5639 1368 5770 1370
rect 5804 1368 5860 1370
rect 5894 1368 5950 1370
rect 5984 1368 6040 1370
rect 6074 1368 6130 1370
rect 6164 1368 6220 1370
rect 6254 1368 6310 1370
rect 6344 1368 6400 1370
rect 6434 1368 6490 1370
rect 6524 1368 6601 1370
rect 5639 1349 6601 1368
rect 5639 1345 5711 1349
rect 5639 1311 5658 1345
rect 5692 1311 5711 1345
rect 5639 1255 5711 1311
rect 6529 1326 6601 1349
rect 6529 1292 6548 1326
rect 6582 1292 6601 1326
rect 5639 1221 5658 1255
rect 5692 1221 5711 1255
rect 5639 1165 5711 1221
rect 5639 1131 5658 1165
rect 5692 1131 5711 1165
rect 5639 1075 5711 1131
rect 5639 1041 5658 1075
rect 5692 1041 5711 1075
rect 5639 985 5711 1041
rect 5639 951 5658 985
rect 5692 951 5711 985
rect 5639 895 5711 951
rect 5639 861 5658 895
rect 5692 861 5711 895
rect 5639 805 5711 861
rect 5639 771 5658 805
rect 5692 771 5711 805
rect 5639 715 5711 771
rect 5639 681 5658 715
rect 5692 681 5711 715
rect 5639 625 5711 681
rect 5639 591 5658 625
rect 5692 591 5711 625
rect 5773 1228 6467 1287
rect 5773 1194 5834 1228
rect 5868 1200 5924 1228
rect 5958 1200 6014 1228
rect 6048 1200 6104 1228
rect 5880 1194 5924 1200
rect 5980 1194 6014 1200
rect 6080 1194 6104 1200
rect 6138 1200 6194 1228
rect 6138 1194 6146 1200
rect 5773 1166 5846 1194
rect 5880 1166 5946 1194
rect 5980 1166 6046 1194
rect 6080 1166 6146 1194
rect 6180 1194 6194 1200
rect 6228 1200 6284 1228
rect 6228 1194 6246 1200
rect 6180 1166 6246 1194
rect 6280 1194 6284 1200
rect 6318 1200 6374 1228
rect 6318 1194 6346 1200
rect 6408 1194 6467 1228
rect 6280 1166 6346 1194
rect 6380 1166 6467 1194
rect 5773 1138 6467 1166
rect 5773 1104 5834 1138
rect 5868 1104 5924 1138
rect 5958 1104 6014 1138
rect 6048 1104 6104 1138
rect 6138 1104 6194 1138
rect 6228 1104 6284 1138
rect 6318 1104 6374 1138
rect 6408 1104 6467 1138
rect 5773 1100 6467 1104
rect 5773 1066 5846 1100
rect 5880 1066 5946 1100
rect 5980 1066 6046 1100
rect 6080 1066 6146 1100
rect 6180 1066 6246 1100
rect 6280 1066 6346 1100
rect 6380 1066 6467 1100
rect 5773 1048 6467 1066
rect 5773 1014 5834 1048
rect 5868 1014 5924 1048
rect 5958 1014 6014 1048
rect 6048 1014 6104 1048
rect 6138 1014 6194 1048
rect 6228 1014 6284 1048
rect 6318 1014 6374 1048
rect 6408 1014 6467 1048
rect 5773 1000 6467 1014
rect 5773 966 5846 1000
rect 5880 966 5946 1000
rect 5980 966 6046 1000
rect 6080 966 6146 1000
rect 6180 966 6246 1000
rect 6280 966 6346 1000
rect 6380 966 6467 1000
rect 5773 958 6467 966
rect 5773 924 5834 958
rect 5868 924 5924 958
rect 5958 924 6014 958
rect 6048 924 6104 958
rect 6138 924 6194 958
rect 6228 924 6284 958
rect 6318 924 6374 958
rect 6408 924 6467 958
rect 5773 900 6467 924
rect 5773 868 5846 900
rect 5880 868 5946 900
rect 5980 868 6046 900
rect 6080 868 6146 900
rect 5773 834 5834 868
rect 5880 866 5924 868
rect 5980 866 6014 868
rect 6080 866 6104 868
rect 5868 834 5924 866
rect 5958 834 6014 866
rect 6048 834 6104 866
rect 6138 866 6146 868
rect 6180 868 6246 900
rect 6180 866 6194 868
rect 6138 834 6194 866
rect 6228 866 6246 868
rect 6280 868 6346 900
rect 6380 868 6467 900
rect 6280 866 6284 868
rect 6228 834 6284 866
rect 6318 866 6346 868
rect 6318 834 6374 866
rect 6408 834 6467 868
rect 5773 800 6467 834
rect 5773 778 5846 800
rect 5880 778 5946 800
rect 5980 778 6046 800
rect 6080 778 6146 800
rect 5773 744 5834 778
rect 5880 766 5924 778
rect 5980 766 6014 778
rect 6080 766 6104 778
rect 5868 744 5924 766
rect 5958 744 6014 766
rect 6048 744 6104 766
rect 6138 766 6146 778
rect 6180 778 6246 800
rect 6180 766 6194 778
rect 6138 744 6194 766
rect 6228 766 6246 778
rect 6280 778 6346 800
rect 6380 778 6467 800
rect 6280 766 6284 778
rect 6228 744 6284 766
rect 6318 766 6346 778
rect 6318 744 6374 766
rect 6408 744 6467 778
rect 5773 700 6467 744
rect 5773 688 5846 700
rect 5880 688 5946 700
rect 5980 688 6046 700
rect 6080 688 6146 700
rect 5773 654 5834 688
rect 5880 666 5924 688
rect 5980 666 6014 688
rect 6080 666 6104 688
rect 5868 654 5924 666
rect 5958 654 6014 666
rect 6048 654 6104 666
rect 6138 666 6146 688
rect 6180 688 6246 700
rect 6180 666 6194 688
rect 6138 654 6194 666
rect 6228 666 6246 688
rect 6280 688 6346 700
rect 6380 688 6467 700
rect 6280 666 6284 688
rect 6228 654 6284 666
rect 6318 666 6346 688
rect 6318 654 6374 666
rect 6408 654 6467 688
rect 5773 593 6467 654
rect 6529 1236 6601 1292
rect 6529 1202 6548 1236
rect 6582 1202 6601 1236
rect 6529 1146 6601 1202
rect 6529 1112 6548 1146
rect 6582 1112 6601 1146
rect 6529 1056 6601 1112
rect 6529 1022 6548 1056
rect 6582 1022 6601 1056
rect 6529 966 6601 1022
rect 6529 932 6548 966
rect 6582 932 6601 966
rect 6529 876 6601 932
rect 6529 842 6548 876
rect 6582 842 6601 876
rect 6529 786 6601 842
rect 6529 752 6548 786
rect 6582 752 6601 786
rect 6529 696 6601 752
rect 6529 662 6548 696
rect 6582 662 6601 696
rect 6529 606 6601 662
rect 5639 531 5711 591
rect 6529 572 6548 606
rect 6582 572 6601 606
rect 6529 531 6601 572
rect 5639 512 6601 531
rect 5639 478 5736 512
rect 5770 478 5826 512
rect 5860 478 5916 512
rect 5950 478 6006 512
rect 6040 478 6096 512
rect 6130 478 6186 512
rect 6220 478 6276 512
rect 6310 478 6366 512
rect 6400 478 6456 512
rect 6490 478 6601 512
rect 5639 459 6601 478
rect 6665 1402 6697 1436
rect 6731 1402 6850 1436
rect 6884 1402 6915 1436
rect 8005 1436 8255 1485
rect 6665 1346 6915 1402
rect 6665 1312 6697 1346
rect 6731 1312 6850 1346
rect 6884 1312 6915 1346
rect 6665 1256 6915 1312
rect 6665 1222 6697 1256
rect 6731 1222 6850 1256
rect 6884 1222 6915 1256
rect 6665 1166 6915 1222
rect 6665 1132 6697 1166
rect 6731 1132 6850 1166
rect 6884 1132 6915 1166
rect 6665 1076 6915 1132
rect 6665 1042 6697 1076
rect 6731 1042 6850 1076
rect 6884 1042 6915 1076
rect 6665 986 6915 1042
rect 6665 952 6697 986
rect 6731 952 6850 986
rect 6884 952 6915 986
rect 6665 896 6915 952
rect 6665 862 6697 896
rect 6731 862 6850 896
rect 6884 862 6915 896
rect 6665 806 6915 862
rect 6665 772 6697 806
rect 6731 772 6850 806
rect 6884 772 6915 806
rect 6665 716 6915 772
rect 6665 682 6697 716
rect 6731 682 6850 716
rect 6884 682 6915 716
rect 6665 626 6915 682
rect 6665 592 6697 626
rect 6731 592 6850 626
rect 6884 592 6915 626
rect 6665 536 6915 592
rect 6665 502 6697 536
rect 6731 502 6850 536
rect 6884 502 6915 536
rect 5325 412 5357 446
rect 5391 412 5510 446
rect 5544 412 5575 446
rect 5325 395 5575 412
rect 6665 446 6915 502
rect 6979 1404 7941 1421
rect 6979 1370 7000 1404
rect 7034 1370 7090 1404
rect 7124 1402 7180 1404
rect 7214 1402 7270 1404
rect 7304 1402 7360 1404
rect 7394 1402 7450 1404
rect 7484 1402 7540 1404
rect 7574 1402 7630 1404
rect 7664 1402 7720 1404
rect 7754 1402 7810 1404
rect 7844 1402 7900 1404
rect 7144 1370 7180 1402
rect 7234 1370 7270 1402
rect 7324 1370 7360 1402
rect 7414 1370 7450 1402
rect 7504 1370 7540 1402
rect 7594 1370 7630 1402
rect 7684 1370 7720 1402
rect 7774 1370 7810 1402
rect 7864 1370 7900 1402
rect 7934 1370 7941 1404
rect 6979 1368 7110 1370
rect 7144 1368 7200 1370
rect 7234 1368 7290 1370
rect 7324 1368 7380 1370
rect 7414 1368 7470 1370
rect 7504 1368 7560 1370
rect 7594 1368 7650 1370
rect 7684 1368 7740 1370
rect 7774 1368 7830 1370
rect 7864 1368 7941 1370
rect 6979 1349 7941 1368
rect 6979 1345 7051 1349
rect 6979 1311 6998 1345
rect 7032 1311 7051 1345
rect 6979 1255 7051 1311
rect 7869 1326 7941 1349
rect 7869 1292 7888 1326
rect 7922 1292 7941 1326
rect 6979 1221 6998 1255
rect 7032 1221 7051 1255
rect 6979 1165 7051 1221
rect 6979 1131 6998 1165
rect 7032 1131 7051 1165
rect 6979 1075 7051 1131
rect 6979 1041 6998 1075
rect 7032 1041 7051 1075
rect 6979 985 7051 1041
rect 6979 951 6998 985
rect 7032 951 7051 985
rect 6979 895 7051 951
rect 6979 861 6998 895
rect 7032 861 7051 895
rect 6979 805 7051 861
rect 6979 771 6998 805
rect 7032 771 7051 805
rect 6979 715 7051 771
rect 6979 681 6998 715
rect 7032 681 7051 715
rect 6979 625 7051 681
rect 6979 591 6998 625
rect 7032 591 7051 625
rect 7113 1228 7807 1287
rect 7113 1194 7174 1228
rect 7208 1200 7264 1228
rect 7298 1200 7354 1228
rect 7388 1200 7444 1228
rect 7220 1194 7264 1200
rect 7320 1194 7354 1200
rect 7420 1194 7444 1200
rect 7478 1200 7534 1228
rect 7478 1194 7486 1200
rect 7113 1166 7186 1194
rect 7220 1166 7286 1194
rect 7320 1166 7386 1194
rect 7420 1166 7486 1194
rect 7520 1194 7534 1200
rect 7568 1200 7624 1228
rect 7568 1194 7586 1200
rect 7520 1166 7586 1194
rect 7620 1194 7624 1200
rect 7658 1200 7714 1228
rect 7658 1194 7686 1200
rect 7748 1194 7807 1228
rect 7620 1166 7686 1194
rect 7720 1166 7807 1194
rect 7113 1138 7807 1166
rect 7113 1104 7174 1138
rect 7208 1104 7264 1138
rect 7298 1104 7354 1138
rect 7388 1104 7444 1138
rect 7478 1104 7534 1138
rect 7568 1104 7624 1138
rect 7658 1104 7714 1138
rect 7748 1104 7807 1138
rect 7113 1100 7807 1104
rect 7113 1066 7186 1100
rect 7220 1066 7286 1100
rect 7320 1066 7386 1100
rect 7420 1066 7486 1100
rect 7520 1066 7586 1100
rect 7620 1066 7686 1100
rect 7720 1066 7807 1100
rect 7113 1048 7807 1066
rect 7113 1014 7174 1048
rect 7208 1014 7264 1048
rect 7298 1014 7354 1048
rect 7388 1014 7444 1048
rect 7478 1014 7534 1048
rect 7568 1014 7624 1048
rect 7658 1014 7714 1048
rect 7748 1014 7807 1048
rect 7113 1000 7807 1014
rect 7113 966 7186 1000
rect 7220 966 7286 1000
rect 7320 966 7386 1000
rect 7420 966 7486 1000
rect 7520 966 7586 1000
rect 7620 966 7686 1000
rect 7720 966 7807 1000
rect 7113 958 7807 966
rect 7113 924 7174 958
rect 7208 924 7264 958
rect 7298 924 7354 958
rect 7388 924 7444 958
rect 7478 924 7534 958
rect 7568 924 7624 958
rect 7658 924 7714 958
rect 7748 924 7807 958
rect 7113 900 7807 924
rect 7113 868 7186 900
rect 7220 868 7286 900
rect 7320 868 7386 900
rect 7420 868 7486 900
rect 7113 834 7174 868
rect 7220 866 7264 868
rect 7320 866 7354 868
rect 7420 866 7444 868
rect 7208 834 7264 866
rect 7298 834 7354 866
rect 7388 834 7444 866
rect 7478 866 7486 868
rect 7520 868 7586 900
rect 7520 866 7534 868
rect 7478 834 7534 866
rect 7568 866 7586 868
rect 7620 868 7686 900
rect 7720 868 7807 900
rect 7620 866 7624 868
rect 7568 834 7624 866
rect 7658 866 7686 868
rect 7658 834 7714 866
rect 7748 834 7807 868
rect 7113 800 7807 834
rect 7113 778 7186 800
rect 7220 778 7286 800
rect 7320 778 7386 800
rect 7420 778 7486 800
rect 7113 744 7174 778
rect 7220 766 7264 778
rect 7320 766 7354 778
rect 7420 766 7444 778
rect 7208 744 7264 766
rect 7298 744 7354 766
rect 7388 744 7444 766
rect 7478 766 7486 778
rect 7520 778 7586 800
rect 7520 766 7534 778
rect 7478 744 7534 766
rect 7568 766 7586 778
rect 7620 778 7686 800
rect 7720 778 7807 800
rect 7620 766 7624 778
rect 7568 744 7624 766
rect 7658 766 7686 778
rect 7658 744 7714 766
rect 7748 744 7807 778
rect 7113 700 7807 744
rect 7113 688 7186 700
rect 7220 688 7286 700
rect 7320 688 7386 700
rect 7420 688 7486 700
rect 7113 654 7174 688
rect 7220 666 7264 688
rect 7320 666 7354 688
rect 7420 666 7444 688
rect 7208 654 7264 666
rect 7298 654 7354 666
rect 7388 654 7444 666
rect 7478 666 7486 688
rect 7520 688 7586 700
rect 7520 666 7534 688
rect 7478 654 7534 666
rect 7568 666 7586 688
rect 7620 688 7686 700
rect 7720 688 7807 700
rect 7620 666 7624 688
rect 7568 654 7624 666
rect 7658 666 7686 688
rect 7658 654 7714 666
rect 7748 654 7807 688
rect 7113 593 7807 654
rect 7869 1236 7941 1292
rect 7869 1202 7888 1236
rect 7922 1202 7941 1236
rect 7869 1146 7941 1202
rect 7869 1112 7888 1146
rect 7922 1112 7941 1146
rect 7869 1056 7941 1112
rect 7869 1022 7888 1056
rect 7922 1022 7941 1056
rect 7869 966 7941 1022
rect 7869 932 7888 966
rect 7922 932 7941 966
rect 7869 876 7941 932
rect 7869 842 7888 876
rect 7922 842 7941 876
rect 7869 786 7941 842
rect 7869 752 7888 786
rect 7922 752 7941 786
rect 7869 696 7941 752
rect 7869 662 7888 696
rect 7922 662 7941 696
rect 7869 606 7941 662
rect 6979 531 7051 591
rect 7869 572 7888 606
rect 7922 572 7941 606
rect 7869 531 7941 572
rect 6979 512 7941 531
rect 6979 478 7076 512
rect 7110 478 7166 512
rect 7200 478 7256 512
rect 7290 478 7346 512
rect 7380 478 7436 512
rect 7470 478 7526 512
rect 7560 478 7616 512
rect 7650 478 7706 512
rect 7740 478 7796 512
rect 7830 478 7941 512
rect 6979 459 7941 478
rect 8005 1402 8037 1436
rect 8071 1402 8190 1436
rect 8224 1402 8255 1436
rect 9345 1436 9444 1485
rect 8005 1346 8255 1402
rect 8005 1312 8037 1346
rect 8071 1312 8190 1346
rect 8224 1312 8255 1346
rect 8005 1256 8255 1312
rect 8005 1222 8037 1256
rect 8071 1222 8190 1256
rect 8224 1222 8255 1256
rect 8005 1166 8255 1222
rect 8005 1132 8037 1166
rect 8071 1132 8190 1166
rect 8224 1132 8255 1166
rect 8005 1076 8255 1132
rect 8005 1042 8037 1076
rect 8071 1042 8190 1076
rect 8224 1042 8255 1076
rect 8005 986 8255 1042
rect 8005 952 8037 986
rect 8071 952 8190 986
rect 8224 952 8255 986
rect 8005 896 8255 952
rect 8005 862 8037 896
rect 8071 862 8190 896
rect 8224 862 8255 896
rect 8005 806 8255 862
rect 8005 772 8037 806
rect 8071 772 8190 806
rect 8224 772 8255 806
rect 8005 716 8255 772
rect 8005 682 8037 716
rect 8071 682 8190 716
rect 8224 682 8255 716
rect 8005 626 8255 682
rect 8005 592 8037 626
rect 8071 592 8190 626
rect 8224 592 8255 626
rect 8005 536 8255 592
rect 8005 502 8037 536
rect 8071 502 8190 536
rect 8224 502 8255 536
rect 6665 412 6697 446
rect 6731 412 6850 446
rect 6884 412 6915 446
rect 6665 395 6915 412
rect 8005 446 8255 502
rect 8319 1404 9281 1421
rect 8319 1370 8340 1404
rect 8374 1370 8430 1404
rect 8464 1402 8520 1404
rect 8554 1402 8610 1404
rect 8644 1402 8700 1404
rect 8734 1402 8790 1404
rect 8824 1402 8880 1404
rect 8914 1402 8970 1404
rect 9004 1402 9060 1404
rect 9094 1402 9150 1404
rect 9184 1402 9240 1404
rect 8484 1370 8520 1402
rect 8574 1370 8610 1402
rect 8664 1370 8700 1402
rect 8754 1370 8790 1402
rect 8844 1370 8880 1402
rect 8934 1370 8970 1402
rect 9024 1370 9060 1402
rect 9114 1370 9150 1402
rect 9204 1370 9240 1402
rect 9274 1370 9281 1404
rect 8319 1368 8450 1370
rect 8484 1368 8540 1370
rect 8574 1368 8630 1370
rect 8664 1368 8720 1370
rect 8754 1368 8810 1370
rect 8844 1368 8900 1370
rect 8934 1368 8990 1370
rect 9024 1368 9080 1370
rect 9114 1368 9170 1370
rect 9204 1368 9281 1370
rect 8319 1349 9281 1368
rect 8319 1345 8391 1349
rect 8319 1311 8338 1345
rect 8372 1311 8391 1345
rect 8319 1255 8391 1311
rect 9209 1326 9281 1349
rect 9209 1292 9228 1326
rect 9262 1292 9281 1326
rect 8319 1221 8338 1255
rect 8372 1221 8391 1255
rect 8319 1165 8391 1221
rect 8319 1131 8338 1165
rect 8372 1131 8391 1165
rect 8319 1075 8391 1131
rect 8319 1041 8338 1075
rect 8372 1041 8391 1075
rect 8319 985 8391 1041
rect 8319 951 8338 985
rect 8372 951 8391 985
rect 8319 895 8391 951
rect 8319 861 8338 895
rect 8372 861 8391 895
rect 8319 805 8391 861
rect 8319 771 8338 805
rect 8372 771 8391 805
rect 8319 715 8391 771
rect 8319 681 8338 715
rect 8372 681 8391 715
rect 8319 625 8391 681
rect 8319 591 8338 625
rect 8372 591 8391 625
rect 8453 1228 9147 1287
rect 8453 1194 8514 1228
rect 8548 1200 8604 1228
rect 8638 1200 8694 1228
rect 8728 1200 8784 1228
rect 8560 1194 8604 1200
rect 8660 1194 8694 1200
rect 8760 1194 8784 1200
rect 8818 1200 8874 1228
rect 8818 1194 8826 1200
rect 8453 1166 8526 1194
rect 8560 1166 8626 1194
rect 8660 1166 8726 1194
rect 8760 1166 8826 1194
rect 8860 1194 8874 1200
rect 8908 1200 8964 1228
rect 8908 1194 8926 1200
rect 8860 1166 8926 1194
rect 8960 1194 8964 1200
rect 8998 1200 9054 1228
rect 8998 1194 9026 1200
rect 9088 1194 9147 1228
rect 8960 1166 9026 1194
rect 9060 1166 9147 1194
rect 8453 1138 9147 1166
rect 8453 1104 8514 1138
rect 8548 1104 8604 1138
rect 8638 1104 8694 1138
rect 8728 1104 8784 1138
rect 8818 1104 8874 1138
rect 8908 1104 8964 1138
rect 8998 1104 9054 1138
rect 9088 1104 9147 1138
rect 8453 1100 9147 1104
rect 8453 1066 8526 1100
rect 8560 1066 8626 1100
rect 8660 1066 8726 1100
rect 8760 1066 8826 1100
rect 8860 1066 8926 1100
rect 8960 1066 9026 1100
rect 9060 1066 9147 1100
rect 8453 1048 9147 1066
rect 8453 1014 8514 1048
rect 8548 1014 8604 1048
rect 8638 1014 8694 1048
rect 8728 1014 8784 1048
rect 8818 1014 8874 1048
rect 8908 1014 8964 1048
rect 8998 1014 9054 1048
rect 9088 1014 9147 1048
rect 8453 1000 9147 1014
rect 8453 966 8526 1000
rect 8560 966 8626 1000
rect 8660 966 8726 1000
rect 8760 966 8826 1000
rect 8860 966 8926 1000
rect 8960 966 9026 1000
rect 9060 966 9147 1000
rect 8453 958 9147 966
rect 8453 924 8514 958
rect 8548 924 8604 958
rect 8638 924 8694 958
rect 8728 924 8784 958
rect 8818 924 8874 958
rect 8908 924 8964 958
rect 8998 924 9054 958
rect 9088 924 9147 958
rect 8453 900 9147 924
rect 8453 868 8526 900
rect 8560 868 8626 900
rect 8660 868 8726 900
rect 8760 868 8826 900
rect 8453 834 8514 868
rect 8560 866 8604 868
rect 8660 866 8694 868
rect 8760 866 8784 868
rect 8548 834 8604 866
rect 8638 834 8694 866
rect 8728 834 8784 866
rect 8818 866 8826 868
rect 8860 868 8926 900
rect 8860 866 8874 868
rect 8818 834 8874 866
rect 8908 866 8926 868
rect 8960 868 9026 900
rect 9060 868 9147 900
rect 8960 866 8964 868
rect 8908 834 8964 866
rect 8998 866 9026 868
rect 8998 834 9054 866
rect 9088 834 9147 868
rect 8453 800 9147 834
rect 8453 778 8526 800
rect 8560 778 8626 800
rect 8660 778 8726 800
rect 8760 778 8826 800
rect 8453 744 8514 778
rect 8560 766 8604 778
rect 8660 766 8694 778
rect 8760 766 8784 778
rect 8548 744 8604 766
rect 8638 744 8694 766
rect 8728 744 8784 766
rect 8818 766 8826 778
rect 8860 778 8926 800
rect 8860 766 8874 778
rect 8818 744 8874 766
rect 8908 766 8926 778
rect 8960 778 9026 800
rect 9060 778 9147 800
rect 8960 766 8964 778
rect 8908 744 8964 766
rect 8998 766 9026 778
rect 8998 744 9054 766
rect 9088 744 9147 778
rect 8453 700 9147 744
rect 8453 688 8526 700
rect 8560 688 8626 700
rect 8660 688 8726 700
rect 8760 688 8826 700
rect 8453 654 8514 688
rect 8560 666 8604 688
rect 8660 666 8694 688
rect 8760 666 8784 688
rect 8548 654 8604 666
rect 8638 654 8694 666
rect 8728 654 8784 666
rect 8818 666 8826 688
rect 8860 688 8926 700
rect 8860 666 8874 688
rect 8818 654 8874 666
rect 8908 666 8926 688
rect 8960 688 9026 700
rect 9060 688 9147 700
rect 8960 666 8964 688
rect 8908 654 8964 666
rect 8998 666 9026 688
rect 8998 654 9054 666
rect 9088 654 9147 688
rect 8453 593 9147 654
rect 9209 1236 9281 1292
rect 9209 1202 9228 1236
rect 9262 1202 9281 1236
rect 9209 1146 9281 1202
rect 9209 1112 9228 1146
rect 9262 1112 9281 1146
rect 9209 1056 9281 1112
rect 9209 1022 9228 1056
rect 9262 1022 9281 1056
rect 9209 966 9281 1022
rect 9209 932 9228 966
rect 9262 932 9281 966
rect 9209 876 9281 932
rect 9209 842 9228 876
rect 9262 842 9281 876
rect 9209 786 9281 842
rect 9209 752 9228 786
rect 9262 752 9281 786
rect 9209 696 9281 752
rect 9209 662 9228 696
rect 9262 662 9281 696
rect 9209 606 9281 662
rect 8319 531 8391 591
rect 9209 572 9228 606
rect 9262 572 9281 606
rect 9209 531 9281 572
rect 8319 512 9281 531
rect 8319 478 8416 512
rect 8450 478 8506 512
rect 8540 478 8596 512
rect 8630 478 8686 512
rect 8720 478 8776 512
rect 8810 478 8866 512
rect 8900 478 8956 512
rect 8990 478 9046 512
rect 9080 478 9136 512
rect 9170 478 9281 512
rect 8319 459 9281 478
rect 9345 1402 9377 1436
rect 9411 1402 9444 1436
rect 9345 1346 9444 1402
rect 9345 1312 9377 1346
rect 9411 1312 9444 1346
rect 9345 1256 9444 1312
rect 9345 1222 9377 1256
rect 9411 1222 9444 1256
rect 9345 1166 9444 1222
rect 9345 1132 9377 1166
rect 9411 1132 9444 1166
rect 9345 1076 9444 1132
rect 9345 1042 9377 1076
rect 9411 1042 9444 1076
rect 9345 986 9444 1042
rect 9345 952 9377 986
rect 9411 952 9444 986
rect 9345 896 9444 952
rect 9345 862 9377 896
rect 9411 862 9444 896
rect 9345 806 9444 862
rect 9345 772 9377 806
rect 9411 772 9444 806
rect 9345 716 9444 772
rect 9345 682 9377 716
rect 9411 682 9444 716
rect 9345 626 9444 682
rect 9345 592 9377 626
rect 9411 592 9444 626
rect 9345 536 9444 592
rect 9345 502 9377 536
rect 9411 502 9444 536
rect 8005 412 8037 446
rect 8071 412 8190 446
rect 8224 412 8255 446
rect 8005 395 8255 412
rect 9345 446 9444 502
rect 9345 412 9377 446
rect 9411 412 9444 446
rect 9345 395 9444 412
rect 116 362 9444 395
rect 116 328 246 362
rect 280 328 336 362
rect 370 328 426 362
rect 460 328 516 362
rect 550 328 606 362
rect 640 328 696 362
rect 730 328 786 362
rect 820 328 876 362
rect 910 328 966 362
rect 1000 328 1056 362
rect 1090 328 1146 362
rect 1180 328 1236 362
rect 1270 328 1586 362
rect 1620 328 1676 362
rect 1710 328 1766 362
rect 1800 328 1856 362
rect 1890 328 1946 362
rect 1980 328 2036 362
rect 2070 328 2126 362
rect 2160 328 2216 362
rect 2250 328 2306 362
rect 2340 328 2396 362
rect 2430 328 2486 362
rect 2520 328 2576 362
rect 2610 328 2926 362
rect 2960 328 3016 362
rect 3050 328 3106 362
rect 3140 328 3196 362
rect 3230 328 3286 362
rect 3320 328 3376 362
rect 3410 328 3466 362
rect 3500 328 3556 362
rect 3590 328 3646 362
rect 3680 328 3736 362
rect 3770 328 3826 362
rect 3860 328 3916 362
rect 3950 328 4266 362
rect 4300 328 4356 362
rect 4390 328 4446 362
rect 4480 328 4536 362
rect 4570 328 4626 362
rect 4660 328 4716 362
rect 4750 328 4806 362
rect 4840 328 4896 362
rect 4930 328 4986 362
rect 5020 328 5076 362
rect 5110 328 5166 362
rect 5200 328 5256 362
rect 5290 328 5606 362
rect 5640 328 5696 362
rect 5730 328 5786 362
rect 5820 328 5876 362
rect 5910 328 5966 362
rect 6000 328 6056 362
rect 6090 328 6146 362
rect 6180 328 6236 362
rect 6270 328 6326 362
rect 6360 328 6416 362
rect 6450 328 6506 362
rect 6540 328 6596 362
rect 6630 328 6946 362
rect 6980 328 7036 362
rect 7070 328 7126 362
rect 7160 328 7216 362
rect 7250 328 7306 362
rect 7340 328 7396 362
rect 7430 328 7486 362
rect 7520 328 7576 362
rect 7610 328 7666 362
rect 7700 328 7756 362
rect 7790 328 7846 362
rect 7880 328 7936 362
rect 7970 328 8286 362
rect 8320 328 8376 362
rect 8410 328 8466 362
rect 8500 328 8556 362
rect 8590 328 8646 362
rect 8680 328 8736 362
rect 8770 328 8826 362
rect 8860 328 8916 362
rect 8950 328 9006 362
rect 9040 328 9096 362
rect 9130 328 9186 362
rect 9220 328 9276 362
rect 9310 328 9444 362
rect 116 296 9444 328
rect 90 -30 260 30
rect 320 -30 460 30
rect 520 -30 660 30
rect 720 -30 860 30
rect 920 -30 1060 30
rect 1120 -30 1260 30
rect 1320 -30 1460 30
rect 1520 -30 1660 30
rect 1720 -30 1860 30
rect 1920 -30 2060 30
rect 2120 -30 2260 30
rect 2320 -30 2460 30
rect 2520 -30 2660 30
rect 2720 -30 2860 30
rect 2920 -30 3060 30
rect 3120 -30 3260 30
rect 3320 -30 3460 30
rect 3520 -30 3660 30
rect 3720 -30 3860 30
rect 3920 -30 4060 30
rect 4120 -30 4260 30
rect 4320 -30 4460 30
rect 4520 -30 4660 30
rect 4720 -30 4860 30
rect 4920 -30 5060 30
rect 5120 -30 5260 30
rect 5320 -30 5460 30
rect 5520 -30 5660 30
rect 5720 -30 5860 30
rect 5920 -30 6060 30
rect 6120 -30 6260 30
rect 6320 -30 6460 30
rect 6520 -30 6660 30
rect 6720 -30 6860 30
rect 6920 -30 7060 30
rect 7120 -30 7260 30
rect 7320 -30 7460 30
rect 7520 -30 7660 30
rect 7720 -30 7860 30
rect 7920 -30 8060 30
rect 8120 -30 8260 30
rect 8320 -30 8460 30
rect 8520 -30 8660 30
rect 8720 -30 8860 30
rect 8920 -30 9060 30
rect 9120 -30 9260 30
rect 9320 -30 9470 30
<< viali >>
rect 260 1850 320 1910
rect 460 1850 520 1910
rect 660 1850 720 1910
rect 860 1850 920 1910
rect 1060 1850 1120 1910
rect 1260 1850 1320 1910
rect 1460 1850 1520 1910
rect 1660 1850 1720 1910
rect 1860 1850 1920 1910
rect 2060 1850 2120 1910
rect 2260 1850 2320 1910
rect 2460 1850 2520 1910
rect 2660 1850 2720 1910
rect 2860 1850 2920 1910
rect 3060 1850 3120 1910
rect 3260 1850 3320 1910
rect 3460 1850 3520 1910
rect 3660 1850 3720 1910
rect 3860 1850 3920 1910
rect 4060 1850 4120 1910
rect 4260 1850 4320 1910
rect 4460 1850 4520 1910
rect 4660 1850 4720 1910
rect 4860 1850 4920 1910
rect 5060 1850 5120 1910
rect 5260 1850 5320 1910
rect 5460 1850 5520 1910
rect 5660 1850 5720 1910
rect 5860 1850 5920 1910
rect 6060 1850 6120 1910
rect 6260 1850 6320 1910
rect 6460 1850 6520 1910
rect 6660 1850 6720 1910
rect 6860 1850 6920 1910
rect 7060 1850 7120 1910
rect 7260 1850 7320 1910
rect 7460 1850 7520 1910
rect 7660 1850 7720 1910
rect 7860 1850 7920 1910
rect 8060 1850 8120 1910
rect 8260 1850 8320 1910
rect 8460 1850 8520 1910
rect 8660 1850 8720 1910
rect 8860 1850 8920 1910
rect 9060 1850 9120 1910
rect 9260 1850 9320 1910
rect 136 1530 170 1564
rect 226 1549 260 1564
rect 316 1549 350 1564
rect 406 1549 440 1564
rect 496 1549 530 1564
rect 586 1549 620 1564
rect 676 1549 710 1564
rect 766 1549 800 1564
rect 856 1549 890 1564
rect 946 1549 980 1564
rect 1036 1549 1070 1564
rect 1126 1549 1160 1564
rect 1216 1549 1250 1564
rect 226 1530 246 1549
rect 246 1530 260 1549
rect 316 1530 336 1549
rect 336 1530 350 1549
rect 406 1530 426 1549
rect 426 1530 440 1549
rect 496 1530 516 1549
rect 516 1530 530 1549
rect 586 1530 606 1549
rect 606 1530 620 1549
rect 676 1530 696 1549
rect 696 1530 710 1549
rect 766 1530 786 1549
rect 786 1530 800 1549
rect 856 1530 876 1549
rect 876 1530 890 1549
rect 946 1530 966 1549
rect 966 1530 980 1549
rect 1036 1530 1056 1549
rect 1056 1530 1070 1549
rect 1126 1530 1146 1549
rect 1146 1530 1160 1549
rect 1216 1530 1236 1549
rect 1236 1530 1250 1549
rect 1306 1530 1340 1564
rect 1476 1530 1510 1564
rect 1566 1549 1600 1564
rect 1656 1549 1690 1564
rect 1746 1549 1780 1564
rect 1836 1549 1870 1564
rect 1926 1549 1960 1564
rect 2016 1549 2050 1564
rect 2106 1549 2140 1564
rect 2196 1549 2230 1564
rect 2286 1549 2320 1564
rect 2376 1549 2410 1564
rect 2466 1549 2500 1564
rect 2556 1549 2590 1564
rect 1566 1530 1586 1549
rect 1586 1530 1600 1549
rect 1656 1530 1676 1549
rect 1676 1530 1690 1549
rect 1746 1530 1766 1549
rect 1766 1530 1780 1549
rect 1836 1530 1856 1549
rect 1856 1530 1870 1549
rect 1926 1530 1946 1549
rect 1946 1530 1960 1549
rect 2016 1530 2036 1549
rect 2036 1530 2050 1549
rect 2106 1530 2126 1549
rect 2126 1530 2140 1549
rect 2196 1530 2216 1549
rect 2216 1530 2230 1549
rect 2286 1530 2306 1549
rect 2306 1530 2320 1549
rect 2376 1530 2396 1549
rect 2396 1530 2410 1549
rect 2466 1530 2486 1549
rect 2486 1530 2500 1549
rect 2556 1530 2576 1549
rect 2576 1530 2590 1549
rect 2646 1530 2680 1564
rect 2816 1530 2850 1564
rect 2906 1549 2940 1564
rect 2996 1549 3030 1564
rect 3086 1549 3120 1564
rect 3176 1549 3210 1564
rect 3266 1549 3300 1564
rect 3356 1549 3390 1564
rect 3446 1549 3480 1564
rect 3536 1549 3570 1564
rect 3626 1549 3660 1564
rect 3716 1549 3750 1564
rect 3806 1549 3840 1564
rect 3896 1549 3930 1564
rect 2906 1530 2926 1549
rect 2926 1530 2940 1549
rect 2996 1530 3016 1549
rect 3016 1530 3030 1549
rect 3086 1530 3106 1549
rect 3106 1530 3120 1549
rect 3176 1530 3196 1549
rect 3196 1530 3210 1549
rect 3266 1530 3286 1549
rect 3286 1530 3300 1549
rect 3356 1530 3376 1549
rect 3376 1530 3390 1549
rect 3446 1530 3466 1549
rect 3466 1530 3480 1549
rect 3536 1530 3556 1549
rect 3556 1530 3570 1549
rect 3626 1530 3646 1549
rect 3646 1530 3660 1549
rect 3716 1530 3736 1549
rect 3736 1530 3750 1549
rect 3806 1530 3826 1549
rect 3826 1530 3840 1549
rect 3896 1530 3916 1549
rect 3916 1530 3930 1549
rect 3986 1530 4020 1564
rect 4156 1530 4190 1564
rect 4246 1549 4280 1564
rect 4336 1549 4370 1564
rect 4426 1549 4460 1564
rect 4516 1549 4550 1564
rect 4606 1549 4640 1564
rect 4696 1549 4730 1564
rect 4786 1549 4820 1564
rect 4876 1549 4910 1564
rect 4966 1549 5000 1564
rect 5056 1549 5090 1564
rect 5146 1549 5180 1564
rect 5236 1549 5270 1564
rect 4246 1530 4266 1549
rect 4266 1530 4280 1549
rect 4336 1530 4356 1549
rect 4356 1530 4370 1549
rect 4426 1530 4446 1549
rect 4446 1530 4460 1549
rect 4516 1530 4536 1549
rect 4536 1530 4550 1549
rect 4606 1530 4626 1549
rect 4626 1530 4640 1549
rect 4696 1530 4716 1549
rect 4716 1530 4730 1549
rect 4786 1530 4806 1549
rect 4806 1530 4820 1549
rect 4876 1530 4896 1549
rect 4896 1530 4910 1549
rect 4966 1530 4986 1549
rect 4986 1530 5000 1549
rect 5056 1530 5076 1549
rect 5076 1530 5090 1549
rect 5146 1530 5166 1549
rect 5166 1530 5180 1549
rect 5236 1530 5256 1549
rect 5256 1530 5270 1549
rect 5326 1530 5360 1564
rect 5496 1530 5530 1564
rect 5586 1549 5620 1564
rect 5676 1549 5710 1564
rect 5766 1549 5800 1564
rect 5856 1549 5890 1564
rect 5946 1549 5980 1564
rect 6036 1549 6070 1564
rect 6126 1549 6160 1564
rect 6216 1549 6250 1564
rect 6306 1549 6340 1564
rect 6396 1549 6430 1564
rect 6486 1549 6520 1564
rect 6576 1549 6610 1564
rect 5586 1530 5606 1549
rect 5606 1530 5620 1549
rect 5676 1530 5696 1549
rect 5696 1530 5710 1549
rect 5766 1530 5786 1549
rect 5786 1530 5800 1549
rect 5856 1530 5876 1549
rect 5876 1530 5890 1549
rect 5946 1530 5966 1549
rect 5966 1530 5980 1549
rect 6036 1530 6056 1549
rect 6056 1530 6070 1549
rect 6126 1530 6146 1549
rect 6146 1530 6160 1549
rect 6216 1530 6236 1549
rect 6236 1530 6250 1549
rect 6306 1530 6326 1549
rect 6326 1530 6340 1549
rect 6396 1530 6416 1549
rect 6416 1530 6430 1549
rect 6486 1530 6506 1549
rect 6506 1530 6520 1549
rect 6576 1530 6596 1549
rect 6596 1530 6610 1549
rect 6666 1530 6700 1564
rect 6836 1530 6870 1564
rect 6926 1549 6960 1564
rect 7016 1549 7050 1564
rect 7106 1549 7140 1564
rect 7196 1549 7230 1564
rect 7286 1549 7320 1564
rect 7376 1549 7410 1564
rect 7466 1549 7500 1564
rect 7556 1549 7590 1564
rect 7646 1549 7680 1564
rect 7736 1549 7770 1564
rect 7826 1549 7860 1564
rect 7916 1549 7950 1564
rect 6926 1530 6946 1549
rect 6946 1530 6960 1549
rect 7016 1530 7036 1549
rect 7036 1530 7050 1549
rect 7106 1530 7126 1549
rect 7126 1530 7140 1549
rect 7196 1530 7216 1549
rect 7216 1530 7230 1549
rect 7286 1530 7306 1549
rect 7306 1530 7320 1549
rect 7376 1530 7396 1549
rect 7396 1530 7410 1549
rect 7466 1530 7486 1549
rect 7486 1530 7500 1549
rect 7556 1530 7576 1549
rect 7576 1530 7590 1549
rect 7646 1530 7666 1549
rect 7666 1530 7680 1549
rect 7736 1530 7756 1549
rect 7756 1530 7770 1549
rect 7826 1530 7846 1549
rect 7846 1530 7860 1549
rect 7916 1530 7936 1549
rect 7936 1530 7950 1549
rect 8006 1530 8040 1564
rect 8176 1530 8210 1564
rect 8266 1549 8300 1564
rect 8356 1549 8390 1564
rect 8446 1549 8480 1564
rect 8536 1549 8570 1564
rect 8626 1549 8660 1564
rect 8716 1549 8750 1564
rect 8806 1549 8840 1564
rect 8896 1549 8930 1564
rect 8986 1549 9020 1564
rect 9076 1549 9110 1564
rect 9166 1549 9200 1564
rect 9256 1549 9290 1564
rect 8266 1530 8286 1549
rect 8286 1530 8300 1549
rect 8356 1530 8376 1549
rect 8376 1530 8390 1549
rect 8446 1530 8466 1549
rect 8466 1530 8480 1549
rect 8536 1530 8556 1549
rect 8556 1530 8570 1549
rect 8626 1530 8646 1549
rect 8646 1530 8660 1549
rect 8716 1530 8736 1549
rect 8736 1530 8750 1549
rect 8806 1530 8826 1549
rect 8826 1530 8840 1549
rect 8896 1530 8916 1549
rect 8916 1530 8930 1549
rect 8986 1530 9006 1549
rect 9006 1530 9020 1549
rect 9076 1530 9096 1549
rect 9096 1530 9110 1549
rect 9166 1530 9186 1549
rect 9186 1530 9200 1549
rect 9256 1530 9276 1549
rect 9276 1530 9290 1549
rect 9346 1530 9380 1564
rect 300 1370 334 1404
rect 390 1402 424 1404
rect 480 1402 514 1404
rect 570 1402 604 1404
rect 660 1402 694 1404
rect 750 1402 784 1404
rect 840 1402 874 1404
rect 930 1402 964 1404
rect 1020 1402 1054 1404
rect 1110 1402 1144 1404
rect 390 1370 410 1402
rect 410 1370 424 1402
rect 480 1370 500 1402
rect 500 1370 514 1402
rect 570 1370 590 1402
rect 590 1370 604 1402
rect 660 1370 680 1402
rect 680 1370 694 1402
rect 750 1370 770 1402
rect 770 1370 784 1402
rect 840 1370 860 1402
rect 860 1370 874 1402
rect 930 1370 950 1402
rect 950 1370 964 1402
rect 1020 1370 1040 1402
rect 1040 1370 1054 1402
rect 1110 1370 1130 1402
rect 1130 1370 1144 1402
rect 1200 1370 1234 1404
rect 486 1194 508 1200
rect 508 1194 520 1200
rect 586 1194 598 1200
rect 598 1194 620 1200
rect 686 1194 688 1200
rect 688 1194 720 1200
rect 486 1166 520 1194
rect 586 1166 620 1194
rect 686 1166 720 1194
rect 786 1166 820 1200
rect 886 1166 920 1200
rect 986 1194 1014 1200
rect 1014 1194 1020 1200
rect 986 1166 1020 1194
rect 486 1066 520 1100
rect 586 1066 620 1100
rect 686 1066 720 1100
rect 786 1066 820 1100
rect 886 1066 920 1100
rect 986 1066 1020 1100
rect 486 966 520 1000
rect 586 966 620 1000
rect 686 966 720 1000
rect 786 966 820 1000
rect 886 966 920 1000
rect 986 966 1020 1000
rect 486 868 520 900
rect 586 868 620 900
rect 686 868 720 900
rect 486 866 508 868
rect 508 866 520 868
rect 586 866 598 868
rect 598 866 620 868
rect 686 866 688 868
rect 688 866 720 868
rect 786 866 820 900
rect 886 866 920 900
rect 986 868 1020 900
rect 986 866 1014 868
rect 1014 866 1020 868
rect 486 778 520 800
rect 586 778 620 800
rect 686 778 720 800
rect 486 766 508 778
rect 508 766 520 778
rect 586 766 598 778
rect 598 766 620 778
rect 686 766 688 778
rect 688 766 720 778
rect 786 766 820 800
rect 886 766 920 800
rect 986 778 1020 800
rect 986 766 1014 778
rect 1014 766 1020 778
rect 486 688 520 700
rect 586 688 620 700
rect 686 688 720 700
rect 486 666 508 688
rect 508 666 520 688
rect 586 666 598 688
rect 598 666 620 688
rect 686 666 688 688
rect 688 666 720 688
rect 786 666 820 700
rect 886 666 920 700
rect 986 688 1020 700
rect 986 666 1014 688
rect 1014 666 1020 688
rect 1640 1370 1674 1404
rect 1730 1402 1764 1404
rect 1820 1402 1854 1404
rect 1910 1402 1944 1404
rect 2000 1402 2034 1404
rect 2090 1402 2124 1404
rect 2180 1402 2214 1404
rect 2270 1402 2304 1404
rect 2360 1402 2394 1404
rect 2450 1402 2484 1404
rect 1730 1370 1750 1402
rect 1750 1370 1764 1402
rect 1820 1370 1840 1402
rect 1840 1370 1854 1402
rect 1910 1370 1930 1402
rect 1930 1370 1944 1402
rect 2000 1370 2020 1402
rect 2020 1370 2034 1402
rect 2090 1370 2110 1402
rect 2110 1370 2124 1402
rect 2180 1370 2200 1402
rect 2200 1370 2214 1402
rect 2270 1370 2290 1402
rect 2290 1370 2304 1402
rect 2360 1370 2380 1402
rect 2380 1370 2394 1402
rect 2450 1370 2470 1402
rect 2470 1370 2484 1402
rect 2540 1370 2574 1404
rect 1826 1194 1848 1200
rect 1848 1194 1860 1200
rect 1926 1194 1938 1200
rect 1938 1194 1960 1200
rect 2026 1194 2028 1200
rect 2028 1194 2060 1200
rect 1826 1166 1860 1194
rect 1926 1166 1960 1194
rect 2026 1166 2060 1194
rect 2126 1166 2160 1200
rect 2226 1166 2260 1200
rect 2326 1194 2354 1200
rect 2354 1194 2360 1200
rect 2326 1166 2360 1194
rect 1826 1066 1860 1100
rect 1926 1066 1960 1100
rect 2026 1066 2060 1100
rect 2126 1066 2160 1100
rect 2226 1066 2260 1100
rect 2326 1066 2360 1100
rect 1826 966 1860 1000
rect 1926 966 1960 1000
rect 2026 966 2060 1000
rect 2126 966 2160 1000
rect 2226 966 2260 1000
rect 2326 966 2360 1000
rect 1826 868 1860 900
rect 1926 868 1960 900
rect 2026 868 2060 900
rect 1826 866 1848 868
rect 1848 866 1860 868
rect 1926 866 1938 868
rect 1938 866 1960 868
rect 2026 866 2028 868
rect 2028 866 2060 868
rect 2126 866 2160 900
rect 2226 866 2260 900
rect 2326 868 2360 900
rect 2326 866 2354 868
rect 2354 866 2360 868
rect 1826 778 1860 800
rect 1926 778 1960 800
rect 2026 778 2060 800
rect 1826 766 1848 778
rect 1848 766 1860 778
rect 1926 766 1938 778
rect 1938 766 1960 778
rect 2026 766 2028 778
rect 2028 766 2060 778
rect 2126 766 2160 800
rect 2226 766 2260 800
rect 2326 778 2360 800
rect 2326 766 2354 778
rect 2354 766 2360 778
rect 1826 688 1860 700
rect 1926 688 1960 700
rect 2026 688 2060 700
rect 1826 666 1848 688
rect 1848 666 1860 688
rect 1926 666 1938 688
rect 1938 666 1960 688
rect 2026 666 2028 688
rect 2028 666 2060 688
rect 2126 666 2160 700
rect 2226 666 2260 700
rect 2326 688 2360 700
rect 2326 666 2354 688
rect 2354 666 2360 688
rect 2980 1370 3014 1404
rect 3070 1402 3104 1404
rect 3160 1402 3194 1404
rect 3250 1402 3284 1404
rect 3340 1402 3374 1404
rect 3430 1402 3464 1404
rect 3520 1402 3554 1404
rect 3610 1402 3644 1404
rect 3700 1402 3734 1404
rect 3790 1402 3824 1404
rect 3070 1370 3090 1402
rect 3090 1370 3104 1402
rect 3160 1370 3180 1402
rect 3180 1370 3194 1402
rect 3250 1370 3270 1402
rect 3270 1370 3284 1402
rect 3340 1370 3360 1402
rect 3360 1370 3374 1402
rect 3430 1370 3450 1402
rect 3450 1370 3464 1402
rect 3520 1370 3540 1402
rect 3540 1370 3554 1402
rect 3610 1370 3630 1402
rect 3630 1370 3644 1402
rect 3700 1370 3720 1402
rect 3720 1370 3734 1402
rect 3790 1370 3810 1402
rect 3810 1370 3824 1402
rect 3880 1370 3914 1404
rect 3166 1194 3188 1200
rect 3188 1194 3200 1200
rect 3266 1194 3278 1200
rect 3278 1194 3300 1200
rect 3366 1194 3368 1200
rect 3368 1194 3400 1200
rect 3166 1166 3200 1194
rect 3266 1166 3300 1194
rect 3366 1166 3400 1194
rect 3466 1166 3500 1200
rect 3566 1166 3600 1200
rect 3666 1194 3694 1200
rect 3694 1194 3700 1200
rect 3666 1166 3700 1194
rect 3166 1066 3200 1100
rect 3266 1066 3300 1100
rect 3366 1066 3400 1100
rect 3466 1066 3500 1100
rect 3566 1066 3600 1100
rect 3666 1066 3700 1100
rect 3166 966 3200 1000
rect 3266 966 3300 1000
rect 3366 966 3400 1000
rect 3466 966 3500 1000
rect 3566 966 3600 1000
rect 3666 966 3700 1000
rect 3166 868 3200 900
rect 3266 868 3300 900
rect 3366 868 3400 900
rect 3166 866 3188 868
rect 3188 866 3200 868
rect 3266 866 3278 868
rect 3278 866 3300 868
rect 3366 866 3368 868
rect 3368 866 3400 868
rect 3466 866 3500 900
rect 3566 866 3600 900
rect 3666 868 3700 900
rect 3666 866 3694 868
rect 3694 866 3700 868
rect 3166 778 3200 800
rect 3266 778 3300 800
rect 3366 778 3400 800
rect 3166 766 3188 778
rect 3188 766 3200 778
rect 3266 766 3278 778
rect 3278 766 3300 778
rect 3366 766 3368 778
rect 3368 766 3400 778
rect 3466 766 3500 800
rect 3566 766 3600 800
rect 3666 778 3700 800
rect 3666 766 3694 778
rect 3694 766 3700 778
rect 3166 688 3200 700
rect 3266 688 3300 700
rect 3366 688 3400 700
rect 3166 666 3188 688
rect 3188 666 3200 688
rect 3266 666 3278 688
rect 3278 666 3300 688
rect 3366 666 3368 688
rect 3368 666 3400 688
rect 3466 666 3500 700
rect 3566 666 3600 700
rect 3666 688 3700 700
rect 3666 666 3694 688
rect 3694 666 3700 688
rect 4320 1370 4354 1404
rect 4410 1402 4444 1404
rect 4500 1402 4534 1404
rect 4590 1402 4624 1404
rect 4680 1402 4714 1404
rect 4770 1402 4804 1404
rect 4860 1402 4894 1404
rect 4950 1402 4984 1404
rect 5040 1402 5074 1404
rect 5130 1402 5164 1404
rect 4410 1370 4430 1402
rect 4430 1370 4444 1402
rect 4500 1370 4520 1402
rect 4520 1370 4534 1402
rect 4590 1370 4610 1402
rect 4610 1370 4624 1402
rect 4680 1370 4700 1402
rect 4700 1370 4714 1402
rect 4770 1370 4790 1402
rect 4790 1370 4804 1402
rect 4860 1370 4880 1402
rect 4880 1370 4894 1402
rect 4950 1370 4970 1402
rect 4970 1370 4984 1402
rect 5040 1370 5060 1402
rect 5060 1370 5074 1402
rect 5130 1370 5150 1402
rect 5150 1370 5164 1402
rect 5220 1370 5254 1404
rect 4506 1194 4528 1200
rect 4528 1194 4540 1200
rect 4606 1194 4618 1200
rect 4618 1194 4640 1200
rect 4706 1194 4708 1200
rect 4708 1194 4740 1200
rect 4506 1166 4540 1194
rect 4606 1166 4640 1194
rect 4706 1166 4740 1194
rect 4806 1166 4840 1200
rect 4906 1166 4940 1200
rect 5006 1194 5034 1200
rect 5034 1194 5040 1200
rect 5006 1166 5040 1194
rect 4506 1066 4540 1100
rect 4606 1066 4640 1100
rect 4706 1066 4740 1100
rect 4806 1066 4840 1100
rect 4906 1066 4940 1100
rect 5006 1066 5040 1100
rect 4506 966 4540 1000
rect 4606 966 4640 1000
rect 4706 966 4740 1000
rect 4806 966 4840 1000
rect 4906 966 4940 1000
rect 5006 966 5040 1000
rect 4506 868 4540 900
rect 4606 868 4640 900
rect 4706 868 4740 900
rect 4506 866 4528 868
rect 4528 866 4540 868
rect 4606 866 4618 868
rect 4618 866 4640 868
rect 4706 866 4708 868
rect 4708 866 4740 868
rect 4806 866 4840 900
rect 4906 866 4940 900
rect 5006 868 5040 900
rect 5006 866 5034 868
rect 5034 866 5040 868
rect 4506 778 4540 800
rect 4606 778 4640 800
rect 4706 778 4740 800
rect 4506 766 4528 778
rect 4528 766 4540 778
rect 4606 766 4618 778
rect 4618 766 4640 778
rect 4706 766 4708 778
rect 4708 766 4740 778
rect 4806 766 4840 800
rect 4906 766 4940 800
rect 5006 778 5040 800
rect 5006 766 5034 778
rect 5034 766 5040 778
rect 4506 688 4540 700
rect 4606 688 4640 700
rect 4706 688 4740 700
rect 4506 666 4528 688
rect 4528 666 4540 688
rect 4606 666 4618 688
rect 4618 666 4640 688
rect 4706 666 4708 688
rect 4708 666 4740 688
rect 4806 666 4840 700
rect 4906 666 4940 700
rect 5006 688 5040 700
rect 5006 666 5034 688
rect 5034 666 5040 688
rect 5660 1370 5694 1404
rect 5750 1402 5784 1404
rect 5840 1402 5874 1404
rect 5930 1402 5964 1404
rect 6020 1402 6054 1404
rect 6110 1402 6144 1404
rect 6200 1402 6234 1404
rect 6290 1402 6324 1404
rect 6380 1402 6414 1404
rect 6470 1402 6504 1404
rect 5750 1370 5770 1402
rect 5770 1370 5784 1402
rect 5840 1370 5860 1402
rect 5860 1370 5874 1402
rect 5930 1370 5950 1402
rect 5950 1370 5964 1402
rect 6020 1370 6040 1402
rect 6040 1370 6054 1402
rect 6110 1370 6130 1402
rect 6130 1370 6144 1402
rect 6200 1370 6220 1402
rect 6220 1370 6234 1402
rect 6290 1370 6310 1402
rect 6310 1370 6324 1402
rect 6380 1370 6400 1402
rect 6400 1370 6414 1402
rect 6470 1370 6490 1402
rect 6490 1370 6504 1402
rect 6560 1370 6594 1404
rect 5846 1194 5868 1200
rect 5868 1194 5880 1200
rect 5946 1194 5958 1200
rect 5958 1194 5980 1200
rect 6046 1194 6048 1200
rect 6048 1194 6080 1200
rect 5846 1166 5880 1194
rect 5946 1166 5980 1194
rect 6046 1166 6080 1194
rect 6146 1166 6180 1200
rect 6246 1166 6280 1200
rect 6346 1194 6374 1200
rect 6374 1194 6380 1200
rect 6346 1166 6380 1194
rect 5846 1066 5880 1100
rect 5946 1066 5980 1100
rect 6046 1066 6080 1100
rect 6146 1066 6180 1100
rect 6246 1066 6280 1100
rect 6346 1066 6380 1100
rect 5846 966 5880 1000
rect 5946 966 5980 1000
rect 6046 966 6080 1000
rect 6146 966 6180 1000
rect 6246 966 6280 1000
rect 6346 966 6380 1000
rect 5846 868 5880 900
rect 5946 868 5980 900
rect 6046 868 6080 900
rect 5846 866 5868 868
rect 5868 866 5880 868
rect 5946 866 5958 868
rect 5958 866 5980 868
rect 6046 866 6048 868
rect 6048 866 6080 868
rect 6146 866 6180 900
rect 6246 866 6280 900
rect 6346 868 6380 900
rect 6346 866 6374 868
rect 6374 866 6380 868
rect 5846 778 5880 800
rect 5946 778 5980 800
rect 6046 778 6080 800
rect 5846 766 5868 778
rect 5868 766 5880 778
rect 5946 766 5958 778
rect 5958 766 5980 778
rect 6046 766 6048 778
rect 6048 766 6080 778
rect 6146 766 6180 800
rect 6246 766 6280 800
rect 6346 778 6380 800
rect 6346 766 6374 778
rect 6374 766 6380 778
rect 5846 688 5880 700
rect 5946 688 5980 700
rect 6046 688 6080 700
rect 5846 666 5868 688
rect 5868 666 5880 688
rect 5946 666 5958 688
rect 5958 666 5980 688
rect 6046 666 6048 688
rect 6048 666 6080 688
rect 6146 666 6180 700
rect 6246 666 6280 700
rect 6346 688 6380 700
rect 6346 666 6374 688
rect 6374 666 6380 688
rect 7000 1370 7034 1404
rect 7090 1402 7124 1404
rect 7180 1402 7214 1404
rect 7270 1402 7304 1404
rect 7360 1402 7394 1404
rect 7450 1402 7484 1404
rect 7540 1402 7574 1404
rect 7630 1402 7664 1404
rect 7720 1402 7754 1404
rect 7810 1402 7844 1404
rect 7090 1370 7110 1402
rect 7110 1370 7124 1402
rect 7180 1370 7200 1402
rect 7200 1370 7214 1402
rect 7270 1370 7290 1402
rect 7290 1370 7304 1402
rect 7360 1370 7380 1402
rect 7380 1370 7394 1402
rect 7450 1370 7470 1402
rect 7470 1370 7484 1402
rect 7540 1370 7560 1402
rect 7560 1370 7574 1402
rect 7630 1370 7650 1402
rect 7650 1370 7664 1402
rect 7720 1370 7740 1402
rect 7740 1370 7754 1402
rect 7810 1370 7830 1402
rect 7830 1370 7844 1402
rect 7900 1370 7934 1404
rect 7186 1194 7208 1200
rect 7208 1194 7220 1200
rect 7286 1194 7298 1200
rect 7298 1194 7320 1200
rect 7386 1194 7388 1200
rect 7388 1194 7420 1200
rect 7186 1166 7220 1194
rect 7286 1166 7320 1194
rect 7386 1166 7420 1194
rect 7486 1166 7520 1200
rect 7586 1166 7620 1200
rect 7686 1194 7714 1200
rect 7714 1194 7720 1200
rect 7686 1166 7720 1194
rect 7186 1066 7220 1100
rect 7286 1066 7320 1100
rect 7386 1066 7420 1100
rect 7486 1066 7520 1100
rect 7586 1066 7620 1100
rect 7686 1066 7720 1100
rect 7186 966 7220 1000
rect 7286 966 7320 1000
rect 7386 966 7420 1000
rect 7486 966 7520 1000
rect 7586 966 7620 1000
rect 7686 966 7720 1000
rect 7186 868 7220 900
rect 7286 868 7320 900
rect 7386 868 7420 900
rect 7186 866 7208 868
rect 7208 866 7220 868
rect 7286 866 7298 868
rect 7298 866 7320 868
rect 7386 866 7388 868
rect 7388 866 7420 868
rect 7486 866 7520 900
rect 7586 866 7620 900
rect 7686 868 7720 900
rect 7686 866 7714 868
rect 7714 866 7720 868
rect 7186 778 7220 800
rect 7286 778 7320 800
rect 7386 778 7420 800
rect 7186 766 7208 778
rect 7208 766 7220 778
rect 7286 766 7298 778
rect 7298 766 7320 778
rect 7386 766 7388 778
rect 7388 766 7420 778
rect 7486 766 7520 800
rect 7586 766 7620 800
rect 7686 778 7720 800
rect 7686 766 7714 778
rect 7714 766 7720 778
rect 7186 688 7220 700
rect 7286 688 7320 700
rect 7386 688 7420 700
rect 7186 666 7208 688
rect 7208 666 7220 688
rect 7286 666 7298 688
rect 7298 666 7320 688
rect 7386 666 7388 688
rect 7388 666 7420 688
rect 7486 666 7520 700
rect 7586 666 7620 700
rect 7686 688 7720 700
rect 7686 666 7714 688
rect 7714 666 7720 688
rect 8340 1370 8374 1404
rect 8430 1402 8464 1404
rect 8520 1402 8554 1404
rect 8610 1402 8644 1404
rect 8700 1402 8734 1404
rect 8790 1402 8824 1404
rect 8880 1402 8914 1404
rect 8970 1402 9004 1404
rect 9060 1402 9094 1404
rect 9150 1402 9184 1404
rect 8430 1370 8450 1402
rect 8450 1370 8464 1402
rect 8520 1370 8540 1402
rect 8540 1370 8554 1402
rect 8610 1370 8630 1402
rect 8630 1370 8644 1402
rect 8700 1370 8720 1402
rect 8720 1370 8734 1402
rect 8790 1370 8810 1402
rect 8810 1370 8824 1402
rect 8880 1370 8900 1402
rect 8900 1370 8914 1402
rect 8970 1370 8990 1402
rect 8990 1370 9004 1402
rect 9060 1370 9080 1402
rect 9080 1370 9094 1402
rect 9150 1370 9170 1402
rect 9170 1370 9184 1402
rect 9240 1370 9274 1404
rect 8526 1194 8548 1200
rect 8548 1194 8560 1200
rect 8626 1194 8638 1200
rect 8638 1194 8660 1200
rect 8726 1194 8728 1200
rect 8728 1194 8760 1200
rect 8526 1166 8560 1194
rect 8626 1166 8660 1194
rect 8726 1166 8760 1194
rect 8826 1166 8860 1200
rect 8926 1166 8960 1200
rect 9026 1194 9054 1200
rect 9054 1194 9060 1200
rect 9026 1166 9060 1194
rect 8526 1066 8560 1100
rect 8626 1066 8660 1100
rect 8726 1066 8760 1100
rect 8826 1066 8860 1100
rect 8926 1066 8960 1100
rect 9026 1066 9060 1100
rect 8526 966 8560 1000
rect 8626 966 8660 1000
rect 8726 966 8760 1000
rect 8826 966 8860 1000
rect 8926 966 8960 1000
rect 9026 966 9060 1000
rect 8526 868 8560 900
rect 8626 868 8660 900
rect 8726 868 8760 900
rect 8526 866 8548 868
rect 8548 866 8560 868
rect 8626 866 8638 868
rect 8638 866 8660 868
rect 8726 866 8728 868
rect 8728 866 8760 868
rect 8826 866 8860 900
rect 8926 866 8960 900
rect 9026 868 9060 900
rect 9026 866 9054 868
rect 9054 866 9060 868
rect 8526 778 8560 800
rect 8626 778 8660 800
rect 8726 778 8760 800
rect 8526 766 8548 778
rect 8548 766 8560 778
rect 8626 766 8638 778
rect 8638 766 8660 778
rect 8726 766 8728 778
rect 8728 766 8760 778
rect 8826 766 8860 800
rect 8926 766 8960 800
rect 9026 778 9060 800
rect 9026 766 9054 778
rect 9054 766 9060 778
rect 8526 688 8560 700
rect 8626 688 8660 700
rect 8726 688 8760 700
rect 8526 666 8548 688
rect 8548 666 8560 688
rect 8626 666 8638 688
rect 8638 666 8660 688
rect 8726 666 8728 688
rect 8728 666 8760 688
rect 8826 666 8860 700
rect 8926 666 8960 700
rect 9026 688 9060 700
rect 9026 666 9054 688
rect 9054 666 9060 688
rect 260 -30 320 30
rect 460 -30 520 30
rect 660 -30 720 30
rect 860 -30 920 30
rect 1060 -30 1120 30
rect 1260 -30 1320 30
rect 1460 -30 1520 30
rect 1660 -30 1720 30
rect 1860 -30 1920 30
rect 2060 -30 2120 30
rect 2260 -30 2320 30
rect 2460 -30 2520 30
rect 2660 -30 2720 30
rect 2860 -30 2920 30
rect 3060 -30 3120 30
rect 3260 -30 3320 30
rect 3460 -30 3520 30
rect 3660 -30 3720 30
rect 3860 -30 3920 30
rect 4060 -30 4120 30
rect 4260 -30 4320 30
rect 4460 -30 4520 30
rect 4660 -30 4720 30
rect 4860 -30 4920 30
rect 5060 -30 5120 30
rect 5260 -30 5320 30
rect 5460 -30 5520 30
rect 5660 -30 5720 30
rect 5860 -30 5920 30
rect 6060 -30 6120 30
rect 6260 -30 6320 30
rect 6460 -30 6520 30
rect 6660 -30 6720 30
rect 6860 -30 6920 30
rect 7060 -30 7120 30
rect 7260 -30 7320 30
rect 7460 -30 7520 30
rect 7660 -30 7720 30
rect 7860 -30 7920 30
rect 8060 -30 8120 30
rect 8260 -30 8320 30
rect 8460 -30 8520 30
rect 8660 -30 8720 30
rect 8860 -30 8920 30
rect 9060 -30 9120 30
rect 9260 -30 9320 30
<< metal1 >>
rect 90 1910 9470 1940
rect 90 1850 260 1910
rect 320 1850 460 1910
rect 520 1850 660 1910
rect 720 1850 860 1910
rect 920 1850 1060 1910
rect 1120 1850 1260 1910
rect 1320 1850 1460 1910
rect 1520 1850 1660 1910
rect 1720 1850 1860 1910
rect 1920 1850 2060 1910
rect 2120 1850 2260 1910
rect 2320 1850 2460 1910
rect 2520 1850 2660 1910
rect 2720 1850 2860 1910
rect 2920 1850 3060 1910
rect 3120 1850 3260 1910
rect 3320 1850 3460 1910
rect 3520 1850 3660 1910
rect 3720 1850 3860 1910
rect 3920 1850 4060 1910
rect 4120 1850 4260 1910
rect 4320 1850 4460 1910
rect 4520 1850 4660 1910
rect 4720 1850 4860 1910
rect 4920 1850 5060 1910
rect 5120 1850 5260 1910
rect 5320 1850 5460 1910
rect 5520 1850 5660 1910
rect 5720 1850 5860 1910
rect 5920 1850 6060 1910
rect 6120 1850 6260 1910
rect 6320 1850 6460 1910
rect 6520 1850 6660 1910
rect 6720 1850 6860 1910
rect 6920 1850 7060 1910
rect 7120 1850 7260 1910
rect 7320 1850 7460 1910
rect 7520 1850 7660 1910
rect 7720 1850 7860 1910
rect 7920 1850 8060 1910
rect 8120 1850 8260 1910
rect 8320 1850 8460 1910
rect 8520 1850 8660 1910
rect 8720 1850 8860 1910
rect 8920 1850 9060 1910
rect 9120 1850 9260 1910
rect 9320 1850 9470 1910
rect 90 1820 9470 1850
rect 116 1564 9444 1570
rect 116 1530 136 1564
rect 170 1530 226 1564
rect 260 1530 316 1564
rect 350 1530 406 1564
rect 440 1530 496 1564
rect 530 1530 586 1564
rect 620 1530 676 1564
rect 710 1530 766 1564
rect 800 1530 856 1564
rect 890 1530 946 1564
rect 980 1530 1036 1564
rect 1070 1530 1126 1564
rect 1160 1530 1216 1564
rect 1250 1530 1306 1564
rect 1340 1530 1476 1564
rect 1510 1530 1566 1564
rect 1600 1530 1656 1564
rect 1690 1530 1746 1564
rect 1780 1530 1836 1564
rect 1870 1530 1926 1564
rect 1960 1530 2016 1564
rect 2050 1530 2106 1564
rect 2140 1530 2196 1564
rect 2230 1530 2286 1564
rect 2320 1530 2376 1564
rect 2410 1530 2466 1564
rect 2500 1530 2556 1564
rect 2590 1530 2646 1564
rect 2680 1530 2816 1564
rect 2850 1530 2906 1564
rect 2940 1530 2996 1564
rect 3030 1530 3086 1564
rect 3120 1530 3176 1564
rect 3210 1530 3266 1564
rect 3300 1530 3356 1564
rect 3390 1530 3446 1564
rect 3480 1530 3536 1564
rect 3570 1530 3626 1564
rect 3660 1530 3716 1564
rect 3750 1530 3806 1564
rect 3840 1530 3896 1564
rect 3930 1530 3986 1564
rect 4020 1530 4156 1564
rect 4190 1530 4246 1564
rect 4280 1530 4336 1564
rect 4370 1530 4426 1564
rect 4460 1530 4516 1564
rect 4550 1530 4606 1564
rect 4640 1530 4696 1564
rect 4730 1530 4786 1564
rect 4820 1530 4876 1564
rect 4910 1530 4966 1564
rect 5000 1530 5056 1564
rect 5090 1530 5146 1564
rect 5180 1530 5236 1564
rect 5270 1530 5326 1564
rect 5360 1530 5496 1564
rect 5530 1530 5586 1564
rect 5620 1530 5676 1564
rect 5710 1530 5766 1564
rect 5800 1530 5856 1564
rect 5890 1530 5946 1564
rect 5980 1530 6036 1564
rect 6070 1530 6126 1564
rect 6160 1530 6216 1564
rect 6250 1530 6306 1564
rect 6340 1530 6396 1564
rect 6430 1530 6486 1564
rect 6520 1530 6576 1564
rect 6610 1530 6666 1564
rect 6700 1530 6836 1564
rect 6870 1530 6926 1564
rect 6960 1530 7016 1564
rect 7050 1530 7106 1564
rect 7140 1530 7196 1564
rect 7230 1530 7286 1564
rect 7320 1530 7376 1564
rect 7410 1530 7466 1564
rect 7500 1530 7556 1564
rect 7590 1530 7646 1564
rect 7680 1530 7736 1564
rect 7770 1530 7826 1564
rect 7860 1530 7916 1564
rect 7950 1530 8006 1564
rect 8040 1530 8176 1564
rect 8210 1530 8266 1564
rect 8300 1530 8356 1564
rect 8390 1530 8446 1564
rect 8480 1530 8536 1564
rect 8570 1530 8626 1564
rect 8660 1530 8716 1564
rect 8750 1530 8806 1564
rect 8840 1530 8896 1564
rect 8930 1530 8986 1564
rect 9020 1530 9076 1564
rect 9110 1530 9166 1564
rect 9200 1530 9256 1564
rect 9290 1530 9346 1564
rect 9380 1530 9444 1564
rect 116 1500 9444 1530
rect 280 1404 9280 1420
rect 280 1370 300 1404
rect 334 1370 390 1404
rect 424 1370 480 1404
rect 514 1370 570 1404
rect 604 1370 660 1404
rect 694 1370 750 1404
rect 784 1370 840 1404
rect 874 1370 930 1404
rect 964 1370 1020 1404
rect 1054 1370 1110 1404
rect 1144 1370 1200 1404
rect 1234 1370 1640 1404
rect 1674 1370 1730 1404
rect 1764 1370 1820 1404
rect 1854 1370 1910 1404
rect 1944 1370 2000 1404
rect 2034 1370 2090 1404
rect 2124 1370 2180 1404
rect 2214 1370 2270 1404
rect 2304 1370 2360 1404
rect 2394 1370 2450 1404
rect 2484 1370 2540 1404
rect 2574 1370 2980 1404
rect 3014 1370 3070 1404
rect 3104 1370 3160 1404
rect 3194 1370 3250 1404
rect 3284 1370 3340 1404
rect 3374 1370 3430 1404
rect 3464 1370 3520 1404
rect 3554 1370 3610 1404
rect 3644 1370 3700 1404
rect 3734 1370 3790 1404
rect 3824 1370 3880 1404
rect 3914 1370 4320 1404
rect 4354 1370 4410 1404
rect 4444 1370 4500 1404
rect 4534 1370 4590 1404
rect 4624 1370 4680 1404
rect 4714 1370 4770 1404
rect 4804 1370 4860 1404
rect 4894 1370 4950 1404
rect 4984 1370 5040 1404
rect 5074 1370 5130 1404
rect 5164 1370 5220 1404
rect 5254 1370 5660 1404
rect 5694 1370 5750 1404
rect 5784 1370 5840 1404
rect 5874 1370 5930 1404
rect 5964 1370 6020 1404
rect 6054 1370 6110 1404
rect 6144 1370 6200 1404
rect 6234 1370 6290 1404
rect 6324 1370 6380 1404
rect 6414 1370 6470 1404
rect 6504 1370 6560 1404
rect 6594 1370 7000 1404
rect 7034 1370 7090 1404
rect 7124 1370 7180 1404
rect 7214 1370 7270 1404
rect 7304 1370 7360 1404
rect 7394 1370 7450 1404
rect 7484 1370 7540 1404
rect 7574 1370 7630 1404
rect 7664 1370 7720 1404
rect 7754 1370 7810 1404
rect 7844 1370 7900 1404
rect 7934 1370 8340 1404
rect 8374 1370 8430 1404
rect 8464 1370 8520 1404
rect 8554 1370 8610 1404
rect 8644 1370 8700 1404
rect 8734 1370 8790 1404
rect 8824 1370 8880 1404
rect 8914 1370 8970 1404
rect 9004 1370 9060 1404
rect 9094 1370 9150 1404
rect 9184 1370 9240 1404
rect 9274 1370 9280 1404
rect 280 1350 9280 1370
rect 454 1200 9106 1246
rect 454 1166 486 1200
rect 520 1166 586 1200
rect 620 1166 686 1200
rect 720 1166 786 1200
rect 820 1166 886 1200
rect 920 1166 986 1200
rect 1020 1166 1826 1200
rect 1860 1166 1926 1200
rect 1960 1166 2026 1200
rect 2060 1166 2126 1200
rect 2160 1166 2226 1200
rect 2260 1166 2326 1200
rect 2360 1166 3166 1200
rect 3200 1166 3266 1200
rect 3300 1166 3366 1200
rect 3400 1166 3466 1200
rect 3500 1166 3566 1200
rect 3600 1166 3666 1200
rect 3700 1166 4506 1200
rect 4540 1166 4606 1200
rect 4640 1166 4706 1200
rect 4740 1166 4806 1200
rect 4840 1166 4906 1200
rect 4940 1166 5006 1200
rect 5040 1166 5846 1200
rect 5880 1166 5946 1200
rect 5980 1166 6046 1200
rect 6080 1166 6146 1200
rect 6180 1166 6246 1200
rect 6280 1166 6346 1200
rect 6380 1166 7186 1200
rect 7220 1166 7286 1200
rect 7320 1166 7386 1200
rect 7420 1166 7486 1200
rect 7520 1166 7586 1200
rect 7620 1166 7686 1200
rect 7720 1166 8526 1200
rect 8560 1166 8626 1200
rect 8660 1166 8726 1200
rect 8760 1166 8826 1200
rect 8860 1166 8926 1200
rect 8960 1166 9026 1200
rect 9060 1166 9106 1200
rect 454 1100 9106 1166
rect 454 1066 486 1100
rect 520 1066 586 1100
rect 620 1066 686 1100
rect 720 1066 786 1100
rect 820 1066 886 1100
rect 920 1066 986 1100
rect 1020 1066 1826 1100
rect 1860 1066 1926 1100
rect 1960 1066 2026 1100
rect 2060 1066 2126 1100
rect 2160 1066 2226 1100
rect 2260 1066 2326 1100
rect 2360 1066 3166 1100
rect 3200 1066 3266 1100
rect 3300 1066 3366 1100
rect 3400 1066 3466 1100
rect 3500 1066 3566 1100
rect 3600 1066 3666 1100
rect 3700 1066 4506 1100
rect 4540 1066 4606 1100
rect 4640 1066 4706 1100
rect 4740 1066 4806 1100
rect 4840 1066 4906 1100
rect 4940 1066 5006 1100
rect 5040 1066 5846 1100
rect 5880 1066 5946 1100
rect 5980 1066 6046 1100
rect 6080 1066 6146 1100
rect 6180 1066 6246 1100
rect 6280 1066 6346 1100
rect 6380 1066 7186 1100
rect 7220 1066 7286 1100
rect 7320 1066 7386 1100
rect 7420 1066 7486 1100
rect 7520 1066 7586 1100
rect 7620 1066 7686 1100
rect 7720 1066 8526 1100
rect 8560 1066 8626 1100
rect 8660 1066 8726 1100
rect 8760 1066 8826 1100
rect 8860 1066 8926 1100
rect 8960 1066 9026 1100
rect 9060 1066 9106 1100
rect 454 1000 9106 1066
rect 454 966 486 1000
rect 520 966 586 1000
rect 620 966 686 1000
rect 720 966 786 1000
rect 820 966 886 1000
rect 920 966 986 1000
rect 1020 966 1826 1000
rect 1860 966 1926 1000
rect 1960 966 2026 1000
rect 2060 966 2126 1000
rect 2160 966 2226 1000
rect 2260 966 2326 1000
rect 2360 966 3166 1000
rect 3200 966 3266 1000
rect 3300 966 3366 1000
rect 3400 966 3466 1000
rect 3500 966 3566 1000
rect 3600 966 3666 1000
rect 3700 966 4506 1000
rect 4540 966 4606 1000
rect 4640 966 4706 1000
rect 4740 966 4806 1000
rect 4840 966 4906 1000
rect 4940 966 5006 1000
rect 5040 966 5846 1000
rect 5880 966 5946 1000
rect 5980 966 6046 1000
rect 6080 966 6146 1000
rect 6180 966 6246 1000
rect 6280 966 6346 1000
rect 6380 966 7186 1000
rect 7220 966 7286 1000
rect 7320 966 7386 1000
rect 7420 966 7486 1000
rect 7520 966 7586 1000
rect 7620 966 7686 1000
rect 7720 966 8526 1000
rect 8560 966 8626 1000
rect 8660 966 8726 1000
rect 8760 966 8826 1000
rect 8860 966 8926 1000
rect 8960 966 9026 1000
rect 9060 966 9106 1000
rect 454 900 9106 966
rect 454 866 486 900
rect 520 866 586 900
rect 620 866 686 900
rect 720 866 786 900
rect 820 866 886 900
rect 920 866 986 900
rect 1020 866 1826 900
rect 1860 866 1926 900
rect 1960 866 2026 900
rect 2060 866 2126 900
rect 2160 866 2226 900
rect 2260 866 2326 900
rect 2360 866 3166 900
rect 3200 866 3266 900
rect 3300 866 3366 900
rect 3400 866 3466 900
rect 3500 866 3566 900
rect 3600 866 3666 900
rect 3700 866 4506 900
rect 4540 866 4606 900
rect 4640 866 4706 900
rect 4740 866 4806 900
rect 4840 866 4906 900
rect 4940 866 5006 900
rect 5040 866 5846 900
rect 5880 866 5946 900
rect 5980 866 6046 900
rect 6080 866 6146 900
rect 6180 866 6246 900
rect 6280 866 6346 900
rect 6380 866 7186 900
rect 7220 866 7286 900
rect 7320 866 7386 900
rect 7420 866 7486 900
rect 7520 866 7586 900
rect 7620 866 7686 900
rect 7720 866 8526 900
rect 8560 866 8626 900
rect 8660 866 8726 900
rect 8760 866 8826 900
rect 8860 866 8926 900
rect 8960 866 9026 900
rect 9060 866 9106 900
rect 454 800 9106 866
rect 454 766 486 800
rect 520 766 586 800
rect 620 766 686 800
rect 720 766 786 800
rect 820 766 886 800
rect 920 766 986 800
rect 1020 766 1826 800
rect 1860 766 1926 800
rect 1960 766 2026 800
rect 2060 766 2126 800
rect 2160 766 2226 800
rect 2260 766 2326 800
rect 2360 766 3166 800
rect 3200 766 3266 800
rect 3300 766 3366 800
rect 3400 766 3466 800
rect 3500 766 3566 800
rect 3600 766 3666 800
rect 3700 766 4506 800
rect 4540 766 4606 800
rect 4640 766 4706 800
rect 4740 766 4806 800
rect 4840 766 4906 800
rect 4940 766 5006 800
rect 5040 766 5846 800
rect 5880 766 5946 800
rect 5980 766 6046 800
rect 6080 766 6146 800
rect 6180 766 6246 800
rect 6280 766 6346 800
rect 6380 766 7186 800
rect 7220 766 7286 800
rect 7320 766 7386 800
rect 7420 766 7486 800
rect 7520 766 7586 800
rect 7620 766 7686 800
rect 7720 766 8526 800
rect 8560 766 8626 800
rect 8660 766 8726 800
rect 8760 766 8826 800
rect 8860 766 8926 800
rect 8960 766 9026 800
rect 9060 766 9106 800
rect 454 700 9106 766
rect 454 666 486 700
rect 520 666 586 700
rect 620 666 686 700
rect 720 666 786 700
rect 820 666 886 700
rect 920 666 986 700
rect 1020 666 1826 700
rect 1860 666 1926 700
rect 1960 666 2026 700
rect 2060 666 2126 700
rect 2160 666 2226 700
rect 2260 666 2326 700
rect 2360 666 3166 700
rect 3200 666 3266 700
rect 3300 666 3366 700
rect 3400 666 3466 700
rect 3500 666 3566 700
rect 3600 666 3666 700
rect 3700 666 4506 700
rect 4540 666 4606 700
rect 4640 666 4706 700
rect 4740 666 4806 700
rect 4840 666 4906 700
rect 4940 666 5006 700
rect 5040 666 5846 700
rect 5880 666 5946 700
rect 5980 666 6046 700
rect 6080 666 6146 700
rect 6180 666 6246 700
rect 6280 666 6346 700
rect 6380 666 7186 700
rect 7220 666 7286 700
rect 7320 666 7386 700
rect 7420 666 7486 700
rect 7520 666 7586 700
rect 7620 666 7686 700
rect 7720 666 8526 700
rect 8560 666 8626 700
rect 8660 666 8726 700
rect 8760 666 8826 700
rect 8860 666 8926 700
rect 8960 666 9026 700
rect 9060 666 9106 700
rect 454 634 9106 666
rect 90 30 9470 60
rect 90 -30 260 30
rect 320 -30 460 30
rect 520 -30 660 30
rect 720 -30 860 30
rect 920 -30 1060 30
rect 1120 -30 1260 30
rect 1320 -30 1460 30
rect 1520 -30 1660 30
rect 1720 -30 1860 30
rect 1920 -30 2060 30
rect 2120 -30 2260 30
rect 2320 -30 2460 30
rect 2520 -30 2660 30
rect 2720 -30 2860 30
rect 2920 -30 3060 30
rect 3120 -30 3260 30
rect 3320 -30 3460 30
rect 3520 -30 3660 30
rect 3720 -30 3860 30
rect 3920 -30 4060 30
rect 4120 -30 4260 30
rect 4320 -30 4460 30
rect 4520 -30 4660 30
rect 4720 -30 4860 30
rect 4920 -30 5060 30
rect 5120 -30 5260 30
rect 5320 -30 5460 30
rect 5520 -30 5660 30
rect 5720 -30 5860 30
rect 5920 -30 6060 30
rect 6120 -30 6260 30
rect 6320 -30 6460 30
rect 6520 -30 6660 30
rect 6720 -30 6860 30
rect 6920 -30 7060 30
rect 7120 -30 7260 30
rect 7320 -30 7460 30
rect 7520 -30 7660 30
rect 7720 -30 7860 30
rect 7920 -30 8060 30
rect 8120 -30 8260 30
rect 8320 -30 8460 30
rect 8520 -30 8660 30
rect 8720 -30 8860 30
rect 8920 -30 9060 30
rect 9120 -30 9260 30
rect 9320 -30 9470 30
rect 90 -60 9470 -30
<< pnp3p40 >>
rect 243 423 1277 1457
rect 1583 423 2617 1457
rect 2923 423 3957 1457
rect 4263 423 5297 1457
rect 5603 423 6637 1457
rect 6943 423 7977 1457
rect 8283 423 9317 1457
<< labels >>
flabel metal1 116 1524 356 1564 1 FreeSans 480 0 0 0 Collector
port 3 n default bidirectional
flabel metal1 280 1372 520 1412 1 FreeSans 480 0 0 0 Base
port 2 n default bidirectional
flabel metal1 630 1010 870 1140 1 FreeSans 480 0 0 0 Emitter
port 1 n default bidirectional
flabel metal1 90 1850 150 1910 1 FreeSans 800 0 0 0 VPWR
port 4 n power bidirectional
flabel metal1 90 -30 150 30 1 FreeSans 800 0 0 0 VGND
port 5 n ground bidirectional
flabel locali 8684 896 8932 1000 0 FreeSans 400 0 0 0 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_5/Emitter
flabel locali 8743 1522 8844 1571 0 FreeSans 400 0 0 0 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_5/Collector
flabel locali 8720 1372 8838 1412 0 FreeSans 400 0 0 0 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_5/Base
flabel locali 7344 896 7592 1000 0 FreeSans 400 0 0 0 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_4/Emitter
flabel locali 7403 1522 7504 1571 0 FreeSans 400 0 0 0 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_4/Collector
flabel locali 7380 1372 7498 1412 0 FreeSans 400 0 0 0 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_4/Base
flabel locali 6004 896 6252 1000 0 FreeSans 400 0 0 0 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_3/Emitter
flabel locali 6063 1522 6164 1571 0 FreeSans 400 0 0 0 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_3/Collector
flabel locali 6040 1372 6158 1412 0 FreeSans 400 0 0 0 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_3/Base
flabel locali 4664 896 4912 1000 0 FreeSans 400 0 0 0 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_2/Emitter
flabel locali 4723 1522 4824 1571 0 FreeSans 400 0 0 0 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_2/Collector
flabel locali 4700 1372 4818 1412 0 FreeSans 400 0 0 0 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_2/Base
flabel locali 3324 896 3572 1000 0 FreeSans 400 0 0 0 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_1/Emitter
flabel locali 3383 1522 3484 1571 0 FreeSans 400 0 0 0 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_1/Collector
flabel locali 3360 1372 3478 1412 0 FreeSans 400 0 0 0 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_1/Base
flabel locali 1984 896 2232 1000 0 FreeSans 400 0 0 0 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0/Emitter
flabel locali 2043 1522 2144 1571 0 FreeSans 400 0 0 0 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0/Collector
flabel locali 2020 1372 2138 1412 0 FreeSans 400 0 0 0 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0/Base
flabel locali 644 896 892 1000 0 FreeSans 400 0 0 0 xm1/Emitter
flabel locali 703 1522 804 1571 0 FreeSans 400 0 0 0 xm1/Collector
flabel locali 680 1372 798 1412 0 FreeSans 400 0 0 0 xm1/Base
<< properties >>
string FIXED_BBOX 0 0 9560 1880
string LEFclass CORE
string LEFsite unitasc
<< end >>
