magic
tech sky130A
magscale 1 2
timestamp 1658609783
<< nwell >>
rect 130 1707 3008 1940
rect 130 1000 3009 1707
rect 131 293 3009 1000
<< pmoslvt >>
rect 225 355 625 1645
rect 683 355 1083 1645
rect 1141 355 1541 1645
rect 1599 355 1999 1645
rect 2057 355 2457 1645
rect 2515 355 2915 1645
<< pdiff >>
rect 167 1633 225 1645
rect 167 367 179 1633
rect 213 367 225 1633
rect 167 355 225 367
rect 625 1633 683 1645
rect 625 367 637 1633
rect 671 367 683 1633
rect 625 355 683 367
rect 1083 1633 1141 1645
rect 1083 367 1095 1633
rect 1129 367 1141 1633
rect 1083 355 1141 367
rect 1541 1633 1599 1645
rect 1541 367 1553 1633
rect 1587 367 1599 1633
rect 1541 355 1599 367
rect 1999 1633 2057 1645
rect 1999 367 2011 1633
rect 2045 367 2057 1633
rect 1999 355 2057 367
rect 2457 1633 2515 1645
rect 2457 367 2469 1633
rect 2503 367 2515 1633
rect 2457 355 2515 367
rect 2915 1633 2973 1645
rect 2915 367 2927 1633
rect 2961 367 2973 1633
rect 2915 355 2973 367
<< pdiffc >>
rect 179 367 213 1633
rect 637 367 671 1633
rect 1095 367 1129 1633
rect 1553 367 1587 1633
rect 2011 367 2045 1633
rect 2469 367 2503 1633
rect 2927 367 2961 1633
<< poly >>
rect 225 1645 625 1671
rect 683 1645 1083 1671
rect 1141 1645 1541 1671
rect 1599 1645 1999 1671
rect 2057 1645 2457 1671
rect 2515 1645 2915 1671
rect 225 329 625 355
rect 683 329 1083 355
rect 1141 329 1541 355
rect 1599 329 1999 355
rect 2057 329 2457 355
rect 2515 329 2915 355
rect 370 182 490 329
rect 826 182 946 329
rect 1282 182 1402 329
rect 1738 182 1858 329
rect 2194 182 2314 329
rect 2650 182 2770 329
rect 130 162 3008 182
rect 130 102 300 162
rect 360 102 700 162
rect 760 102 1100 162
rect 1160 102 1500 162
rect 1560 102 1900 162
rect 1960 102 2300 162
rect 2360 102 2700 162
rect 2760 102 3008 162
rect 130 82 3008 102
<< polycont >>
rect 300 102 360 162
rect 700 102 760 162
rect 1100 102 1160 162
rect 1500 102 1560 162
rect 1900 102 1960 162
rect 2300 102 2360 162
rect 2700 102 2760 162
<< locali >>
rect 130 1850 300 1910
rect 360 1850 700 1910
rect 760 1850 1100 1910
rect 1160 1850 1500 1910
rect 1560 1850 1900 1910
rect 1960 1850 2300 1910
rect 2360 1850 2700 1910
rect 2760 1850 3008 1910
rect 130 1730 3008 1790
rect 635 1649 669 1730
rect 1551 1649 1585 1730
rect 2467 1649 2501 1730
rect 179 1633 213 1649
rect 177 367 179 372
rect 635 1633 671 1649
rect 635 1626 637 1633
rect 177 351 213 367
rect 1095 1633 1129 1649
rect 637 351 671 367
rect 1093 367 1095 372
rect 1551 1633 1587 1649
rect 1551 1626 1553 1633
rect 1093 351 1129 367
rect 2011 1633 2045 1649
rect 1553 351 1587 367
rect 2009 367 2011 372
rect 2467 1633 2503 1649
rect 2467 1626 2469 1633
rect 2009 351 2045 367
rect 2927 1633 2961 1649
rect 2469 351 2503 367
rect 2925 367 2927 372
rect 2925 351 2961 367
rect 177 270 211 351
rect 1093 270 1127 351
rect 2009 270 2043 351
rect 2925 270 2959 351
rect 130 210 3008 270
rect 130 102 300 162
rect 360 102 700 162
rect 760 102 1100 162
rect 1160 102 1500 162
rect 1560 102 1900 162
rect 1960 102 2300 162
rect 2360 102 2700 162
rect 2760 102 3008 162
rect 130 -30 300 30
rect 360 -30 700 30
rect 760 -30 1100 30
rect 1160 -30 1500 30
rect 1560 -30 1900 30
rect 1960 -30 2300 30
rect 2360 -30 2700 30
rect 2760 -30 3008 30
<< viali >>
rect 300 1850 360 1910
rect 700 1850 760 1910
rect 1100 1850 1160 1910
rect 1500 1850 1560 1910
rect 1900 1850 1960 1910
rect 2300 1850 2360 1910
rect 2700 1850 2760 1910
rect 179 367 213 1633
rect 637 367 671 1633
rect 1095 367 1129 1633
rect 1553 367 1587 1633
rect 2011 367 2045 1633
rect 2469 367 2503 1633
rect 2927 367 2961 1633
rect 300 -30 360 30
rect 700 -30 760 30
rect 1100 -30 1160 30
rect 1500 -30 1560 30
rect 1900 -30 1960 30
rect 2300 -30 2360 30
rect 2700 -30 2760 30
<< metal1 >>
rect 130 1910 3008 1940
rect 130 1850 300 1910
rect 360 1850 700 1910
rect 760 1850 1100 1910
rect 1160 1850 1500 1910
rect 1560 1850 1900 1910
rect 1960 1850 2300 1910
rect 2360 1850 2700 1910
rect 2760 1850 3008 1910
rect 130 1820 3008 1850
rect 173 1633 219 1645
rect 173 367 179 1633
rect 213 367 219 1633
rect 173 355 219 367
rect 631 1633 677 1645
rect 631 367 637 1633
rect 671 367 677 1633
rect 631 355 677 367
rect 1089 1633 1135 1645
rect 1089 367 1095 1633
rect 1129 367 1135 1633
rect 1089 355 1135 367
rect 1547 1633 1593 1645
rect 1547 367 1553 1633
rect 1587 367 1593 1633
rect 1547 355 1593 367
rect 2005 1633 2051 1645
rect 2005 367 2011 1633
rect 2045 367 2051 1633
rect 2005 355 2051 367
rect 2463 1633 2509 1645
rect 2463 367 2469 1633
rect 2503 367 2509 1633
rect 2463 355 2509 367
rect 2921 1633 2967 1645
rect 2921 367 2927 1633
rect 2961 367 2967 1633
rect 2921 355 2967 367
rect 130 30 3008 60
rect 130 -30 300 30
rect 360 -30 700 30
rect 760 -30 1100 30
rect 1160 -30 1500 30
rect 1560 -30 1900 30
rect 1960 -30 2300 30
rect 2360 -30 2700 30
rect 2760 -30 3008 30
rect 130 -60 3008 -30
<< labels >>
flabel metal1 130 1850 190 1910 1 FreeSans 480 0 0 0 VPWR
port 4 n power bidirectional
flabel space 120 1850 180 1910 1 FreeSans 480 0 0 0 VPB
flabel metal1 130 -30 190 30 1 FreeSans 480 0 0 0 VGND
port 5 n ground bidirectional
flabel locali 2948 1730 3008 1790 1 FreeSans 480 0 0 0 SOURCE
port 2 n signal bidirectional
flabel locali 2948 210 3008 270 1 FreeSans 480 0 0 0 DRAIN
port 3 n signal bidirectional
flabel locali 2948 102 3008 162 1 FreeSans 480 0 0 0 GATE
port 1 n signal bidirectional
<< properties >>
string FIXED_BBOX 0 0 3395 1880
string LEFclass CORE
string LEFsite unitasc
<< end >>
