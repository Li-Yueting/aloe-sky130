VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO switch
  CLASS BLOCK ;
  FOREIGN switch ;
  ORIGIN 0.000 0.000 ;
  SIZE 29.230 BY 207.160 ;
  PIN out
    DIRECTION INOUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 116.710396 ;
    PORT
      LAYER li1 ;
        RECT 19.935 203.420 20.105 204.820 ;
        RECT 20.895 203.420 21.065 204.820 ;
        RECT 21.855 203.420 22.025 204.820 ;
        RECT 22.815 203.420 22.985 204.820 ;
        RECT 23.775 203.420 23.945 204.820 ;
        RECT 24.735 203.420 24.905 204.820 ;
        RECT 19.935 201.360 20.105 201.920 ;
        RECT 20.895 201.360 21.065 201.920 ;
        RECT 21.855 201.360 22.025 201.920 ;
        RECT 22.815 201.360 22.985 201.920 ;
        RECT 23.775 201.360 23.945 201.920 ;
        RECT 24.735 201.360 24.905 201.920 ;
        RECT 19.935 196.985 20.105 198.385 ;
        RECT 20.895 196.985 21.065 198.385 ;
        RECT 21.855 196.985 22.025 198.385 ;
        RECT 22.815 196.985 22.985 198.385 ;
        RECT 23.775 196.985 23.945 198.385 ;
        RECT 24.735 196.985 24.905 198.385 ;
        RECT 19.935 194.925 20.105 195.485 ;
        RECT 20.895 194.925 21.065 195.485 ;
        RECT 21.855 194.925 22.025 195.485 ;
        RECT 22.815 194.925 22.985 195.485 ;
        RECT 23.775 194.925 23.945 195.485 ;
        RECT 24.735 194.925 24.905 195.485 ;
        RECT 19.935 190.550 20.105 191.950 ;
        RECT 20.895 190.550 21.065 191.950 ;
        RECT 21.855 190.550 22.025 191.950 ;
        RECT 22.815 190.550 22.985 191.950 ;
        RECT 23.775 190.550 23.945 191.950 ;
        RECT 24.735 190.550 24.905 191.950 ;
        RECT 19.935 188.490 20.105 189.050 ;
        RECT 20.895 188.490 21.065 189.050 ;
        RECT 21.855 188.490 22.025 189.050 ;
        RECT 22.815 188.490 22.985 189.050 ;
        RECT 23.775 188.490 23.945 189.050 ;
        RECT 24.735 188.490 24.905 189.050 ;
        RECT 19.935 184.115 20.105 185.515 ;
        RECT 20.895 184.115 21.065 185.515 ;
        RECT 21.855 184.115 22.025 185.515 ;
        RECT 22.815 184.115 22.985 185.515 ;
        RECT 23.775 184.115 23.945 185.515 ;
        RECT 24.735 184.115 24.905 185.515 ;
        RECT 19.935 182.055 20.105 182.615 ;
        RECT 20.895 182.055 21.065 182.615 ;
        RECT 21.855 182.055 22.025 182.615 ;
        RECT 22.815 182.055 22.985 182.615 ;
        RECT 23.775 182.055 23.945 182.615 ;
        RECT 24.735 182.055 24.905 182.615 ;
        RECT 19.935 177.680 20.105 179.080 ;
        RECT 20.895 177.680 21.065 179.080 ;
        RECT 21.855 177.680 22.025 179.080 ;
        RECT 22.815 177.680 22.985 179.080 ;
        RECT 23.775 177.680 23.945 179.080 ;
        RECT 24.735 177.680 24.905 179.080 ;
        RECT 19.935 175.620 20.105 176.180 ;
        RECT 20.895 175.620 21.065 176.180 ;
        RECT 21.855 175.620 22.025 176.180 ;
        RECT 22.815 175.620 22.985 176.180 ;
        RECT 23.775 175.620 23.945 176.180 ;
        RECT 24.735 175.620 24.905 176.180 ;
        RECT 19.935 171.245 20.105 172.645 ;
        RECT 20.895 171.245 21.065 172.645 ;
        RECT 21.855 171.245 22.025 172.645 ;
        RECT 22.815 171.245 22.985 172.645 ;
        RECT 23.775 171.245 23.945 172.645 ;
        RECT 24.735 171.245 24.905 172.645 ;
        RECT 19.935 169.185 20.105 169.745 ;
        RECT 20.895 169.185 21.065 169.745 ;
        RECT 21.855 169.185 22.025 169.745 ;
        RECT 22.815 169.185 22.985 169.745 ;
        RECT 23.775 169.185 23.945 169.745 ;
        RECT 24.735 169.185 24.905 169.745 ;
        RECT 19.935 164.810 20.105 166.210 ;
        RECT 20.895 164.810 21.065 166.210 ;
        RECT 21.855 164.810 22.025 166.210 ;
        RECT 22.815 164.810 22.985 166.210 ;
        RECT 23.775 164.810 23.945 166.210 ;
        RECT 24.735 164.810 24.905 166.210 ;
        RECT 19.935 162.750 20.105 163.310 ;
        RECT 20.895 162.750 21.065 163.310 ;
        RECT 21.855 162.750 22.025 163.310 ;
        RECT 22.815 162.750 22.985 163.310 ;
        RECT 23.775 162.750 23.945 163.310 ;
        RECT 24.735 162.750 24.905 163.310 ;
        RECT 19.935 158.375 20.105 159.775 ;
        RECT 20.895 158.375 21.065 159.775 ;
        RECT 21.855 158.375 22.025 159.775 ;
        RECT 22.815 158.375 22.985 159.775 ;
        RECT 23.775 158.375 23.945 159.775 ;
        RECT 24.735 158.375 24.905 159.775 ;
        RECT 19.935 156.315 20.105 156.875 ;
        RECT 20.895 156.315 21.065 156.875 ;
        RECT 21.855 156.315 22.025 156.875 ;
        RECT 22.815 156.315 22.985 156.875 ;
        RECT 23.775 156.315 23.945 156.875 ;
        RECT 24.735 156.315 24.905 156.875 ;
        RECT 19.935 151.940 20.105 153.340 ;
        RECT 20.895 151.940 21.065 153.340 ;
        RECT 21.855 151.940 22.025 153.340 ;
        RECT 22.815 151.940 22.985 153.340 ;
        RECT 23.775 151.940 23.945 153.340 ;
        RECT 24.735 151.940 24.905 153.340 ;
        RECT 19.935 149.880 20.105 150.440 ;
        RECT 20.895 149.880 21.065 150.440 ;
        RECT 21.855 149.880 22.025 150.440 ;
        RECT 22.815 149.880 22.985 150.440 ;
        RECT 23.775 149.880 23.945 150.440 ;
        RECT 24.735 149.880 24.905 150.440 ;
        RECT 19.935 145.505 20.105 146.905 ;
        RECT 20.895 145.505 21.065 146.905 ;
        RECT 21.855 145.505 22.025 146.905 ;
        RECT 22.815 145.505 22.985 146.905 ;
        RECT 23.775 145.505 23.945 146.905 ;
        RECT 24.735 145.505 24.905 146.905 ;
        RECT 19.935 143.445 20.105 144.005 ;
        RECT 20.895 143.445 21.065 144.005 ;
        RECT 21.855 143.445 22.025 144.005 ;
        RECT 22.815 143.445 22.985 144.005 ;
        RECT 23.775 143.445 23.945 144.005 ;
        RECT 24.735 143.445 24.905 144.005 ;
        RECT 19.935 139.070 20.105 140.470 ;
        RECT 20.895 139.070 21.065 140.470 ;
        RECT 21.855 139.070 22.025 140.470 ;
        RECT 22.815 139.070 22.985 140.470 ;
        RECT 23.775 139.070 23.945 140.470 ;
        RECT 24.735 139.070 24.905 140.470 ;
        RECT 19.935 137.010 20.105 137.570 ;
        RECT 20.895 137.010 21.065 137.570 ;
        RECT 21.855 137.010 22.025 137.570 ;
        RECT 22.815 137.010 22.985 137.570 ;
        RECT 23.775 137.010 23.945 137.570 ;
        RECT 24.735 137.010 24.905 137.570 ;
        RECT 19.935 132.635 20.105 134.035 ;
        RECT 20.895 132.635 21.065 134.035 ;
        RECT 21.855 132.635 22.025 134.035 ;
        RECT 22.815 132.635 22.985 134.035 ;
        RECT 23.775 132.635 23.945 134.035 ;
        RECT 24.735 132.635 24.905 134.035 ;
        RECT 19.935 130.575 20.105 131.135 ;
        RECT 20.895 130.575 21.065 131.135 ;
        RECT 21.855 130.575 22.025 131.135 ;
        RECT 22.815 130.575 22.985 131.135 ;
        RECT 23.775 130.575 23.945 131.135 ;
        RECT 24.735 130.575 24.905 131.135 ;
        RECT 19.935 126.200 20.105 127.600 ;
        RECT 20.895 126.200 21.065 127.600 ;
        RECT 21.855 126.200 22.025 127.600 ;
        RECT 22.815 126.200 22.985 127.600 ;
        RECT 23.775 126.200 23.945 127.600 ;
        RECT 24.735 126.200 24.905 127.600 ;
        RECT 19.935 124.140 20.105 124.700 ;
        RECT 20.895 124.140 21.065 124.700 ;
        RECT 21.855 124.140 22.025 124.700 ;
        RECT 22.815 124.140 22.985 124.700 ;
        RECT 23.775 124.140 23.945 124.700 ;
        RECT 24.735 124.140 24.905 124.700 ;
        RECT 19.935 119.765 20.105 121.165 ;
        RECT 20.895 119.765 21.065 121.165 ;
        RECT 21.855 119.765 22.025 121.165 ;
        RECT 22.815 119.765 22.985 121.165 ;
        RECT 23.775 119.765 23.945 121.165 ;
        RECT 24.735 119.765 24.905 121.165 ;
        RECT 19.935 117.705 20.105 118.265 ;
        RECT 20.895 117.705 21.065 118.265 ;
        RECT 21.855 117.705 22.025 118.265 ;
        RECT 22.815 117.705 22.985 118.265 ;
        RECT 23.775 117.705 23.945 118.265 ;
        RECT 24.735 117.705 24.905 118.265 ;
        RECT 19.935 113.330 20.105 114.730 ;
        RECT 20.895 113.330 21.065 114.730 ;
        RECT 21.855 113.330 22.025 114.730 ;
        RECT 22.815 113.330 22.985 114.730 ;
        RECT 23.775 113.330 23.945 114.730 ;
        RECT 24.735 113.330 24.905 114.730 ;
        RECT 19.935 111.270 20.105 111.830 ;
        RECT 20.895 111.270 21.065 111.830 ;
        RECT 21.855 111.270 22.025 111.830 ;
        RECT 22.815 111.270 22.985 111.830 ;
        RECT 23.775 111.270 23.945 111.830 ;
        RECT 24.735 111.270 24.905 111.830 ;
        RECT 19.935 106.895 20.105 108.295 ;
        RECT 20.895 106.895 21.065 108.295 ;
        RECT 21.855 106.895 22.025 108.295 ;
        RECT 22.815 106.895 22.985 108.295 ;
        RECT 23.775 106.895 23.945 108.295 ;
        RECT 24.735 106.895 24.905 108.295 ;
        RECT 19.935 104.835 20.105 105.395 ;
        RECT 20.895 104.835 21.065 105.395 ;
        RECT 21.855 104.835 22.025 105.395 ;
        RECT 22.815 104.835 22.985 105.395 ;
        RECT 23.775 104.835 23.945 105.395 ;
        RECT 24.735 104.835 24.905 105.395 ;
        RECT 19.935 100.460 20.105 101.860 ;
        RECT 20.895 100.460 21.065 101.860 ;
        RECT 21.855 100.460 22.025 101.860 ;
        RECT 22.815 100.460 22.985 101.860 ;
        RECT 23.775 100.460 23.945 101.860 ;
        RECT 24.735 100.460 24.905 101.860 ;
        RECT 19.935 98.400 20.105 98.960 ;
        RECT 20.895 98.400 21.065 98.960 ;
        RECT 21.855 98.400 22.025 98.960 ;
        RECT 22.815 98.400 22.985 98.960 ;
        RECT 23.775 98.400 23.945 98.960 ;
        RECT 24.735 98.400 24.905 98.960 ;
        RECT 19.935 94.025 20.105 95.425 ;
        RECT 20.895 94.025 21.065 95.425 ;
        RECT 21.855 94.025 22.025 95.425 ;
        RECT 22.815 94.025 22.985 95.425 ;
        RECT 23.775 94.025 23.945 95.425 ;
        RECT 24.735 94.025 24.905 95.425 ;
        RECT 19.935 91.965 20.105 92.525 ;
        RECT 20.895 91.965 21.065 92.525 ;
        RECT 21.855 91.965 22.025 92.525 ;
        RECT 22.815 91.965 22.985 92.525 ;
        RECT 23.775 91.965 23.945 92.525 ;
        RECT 24.735 91.965 24.905 92.525 ;
        RECT 19.935 87.590 20.105 88.990 ;
        RECT 20.895 87.590 21.065 88.990 ;
        RECT 21.855 87.590 22.025 88.990 ;
        RECT 22.815 87.590 22.985 88.990 ;
        RECT 23.775 87.590 23.945 88.990 ;
        RECT 24.735 87.590 24.905 88.990 ;
        RECT 19.935 85.530 20.105 86.090 ;
        RECT 20.895 85.530 21.065 86.090 ;
        RECT 21.855 85.530 22.025 86.090 ;
        RECT 22.815 85.530 22.985 86.090 ;
        RECT 23.775 85.530 23.945 86.090 ;
        RECT 24.735 85.530 24.905 86.090 ;
        RECT 19.935 81.155 20.105 82.555 ;
        RECT 20.895 81.155 21.065 82.555 ;
        RECT 21.855 81.155 22.025 82.555 ;
        RECT 22.815 81.155 22.985 82.555 ;
        RECT 23.775 81.155 23.945 82.555 ;
        RECT 24.735 81.155 24.905 82.555 ;
        RECT 19.935 79.095 20.105 79.655 ;
        RECT 20.895 79.095 21.065 79.655 ;
        RECT 21.855 79.095 22.025 79.655 ;
        RECT 22.815 79.095 22.985 79.655 ;
        RECT 23.775 79.095 23.945 79.655 ;
        RECT 24.735 79.095 24.905 79.655 ;
        RECT 19.935 74.720 20.105 76.120 ;
        RECT 20.895 74.720 21.065 76.120 ;
        RECT 21.855 74.720 22.025 76.120 ;
        RECT 22.815 74.720 22.985 76.120 ;
        RECT 23.775 74.720 23.945 76.120 ;
        RECT 24.735 74.720 24.905 76.120 ;
        RECT 19.935 72.660 20.105 73.220 ;
        RECT 20.895 72.660 21.065 73.220 ;
        RECT 21.855 72.660 22.025 73.220 ;
        RECT 22.815 72.660 22.985 73.220 ;
        RECT 23.775 72.660 23.945 73.220 ;
        RECT 24.735 72.660 24.905 73.220 ;
        RECT 19.935 68.285 20.105 69.685 ;
        RECT 20.895 68.285 21.065 69.685 ;
        RECT 21.855 68.285 22.025 69.685 ;
        RECT 22.815 68.285 22.985 69.685 ;
        RECT 23.775 68.285 23.945 69.685 ;
        RECT 24.735 68.285 24.905 69.685 ;
        RECT 19.935 66.225 20.105 66.785 ;
        RECT 20.895 66.225 21.065 66.785 ;
        RECT 21.855 66.225 22.025 66.785 ;
        RECT 22.815 66.225 22.985 66.785 ;
        RECT 23.775 66.225 23.945 66.785 ;
        RECT 24.735 66.225 24.905 66.785 ;
        RECT 19.935 61.850 20.105 63.250 ;
        RECT 20.895 61.850 21.065 63.250 ;
        RECT 21.855 61.850 22.025 63.250 ;
        RECT 22.815 61.850 22.985 63.250 ;
        RECT 23.775 61.850 23.945 63.250 ;
        RECT 24.735 61.850 24.905 63.250 ;
        RECT 19.935 59.790 20.105 60.350 ;
        RECT 20.895 59.790 21.065 60.350 ;
        RECT 21.855 59.790 22.025 60.350 ;
        RECT 22.815 59.790 22.985 60.350 ;
        RECT 23.775 59.790 23.945 60.350 ;
        RECT 24.735 59.790 24.905 60.350 ;
        RECT 19.935 55.415 20.105 56.815 ;
        RECT 20.895 55.415 21.065 56.815 ;
        RECT 21.855 55.415 22.025 56.815 ;
        RECT 22.815 55.415 22.985 56.815 ;
        RECT 23.775 55.415 23.945 56.815 ;
        RECT 24.735 55.415 24.905 56.815 ;
        RECT 19.935 53.355 20.105 53.915 ;
        RECT 20.895 53.355 21.065 53.915 ;
        RECT 21.855 53.355 22.025 53.915 ;
        RECT 22.815 53.355 22.985 53.915 ;
        RECT 23.775 53.355 23.945 53.915 ;
        RECT 24.735 53.355 24.905 53.915 ;
        RECT 19.935 48.980 20.105 50.380 ;
        RECT 20.895 48.980 21.065 50.380 ;
        RECT 21.855 48.980 22.025 50.380 ;
        RECT 22.815 48.980 22.985 50.380 ;
        RECT 23.775 48.980 23.945 50.380 ;
        RECT 24.735 48.980 24.905 50.380 ;
        RECT 19.935 46.920 20.105 47.480 ;
        RECT 20.895 46.920 21.065 47.480 ;
        RECT 21.855 46.920 22.025 47.480 ;
        RECT 22.815 46.920 22.985 47.480 ;
        RECT 23.775 46.920 23.945 47.480 ;
        RECT 24.735 46.920 24.905 47.480 ;
        RECT 19.935 42.545 20.105 43.945 ;
        RECT 20.895 42.545 21.065 43.945 ;
        RECT 21.855 42.545 22.025 43.945 ;
        RECT 22.815 42.545 22.985 43.945 ;
        RECT 23.775 42.545 23.945 43.945 ;
        RECT 24.735 42.545 24.905 43.945 ;
        RECT 19.935 40.485 20.105 41.045 ;
        RECT 20.895 40.485 21.065 41.045 ;
        RECT 21.855 40.485 22.025 41.045 ;
        RECT 22.815 40.485 22.985 41.045 ;
        RECT 23.775 40.485 23.945 41.045 ;
        RECT 24.735 40.485 24.905 41.045 ;
        RECT 19.935 36.110 20.105 37.510 ;
        RECT 20.895 36.110 21.065 37.510 ;
        RECT 21.855 36.110 22.025 37.510 ;
        RECT 22.815 36.110 22.985 37.510 ;
        RECT 23.775 36.110 23.945 37.510 ;
        RECT 24.735 36.110 24.905 37.510 ;
        RECT 19.935 34.050 20.105 34.610 ;
        RECT 20.895 34.050 21.065 34.610 ;
        RECT 21.855 34.050 22.025 34.610 ;
        RECT 22.815 34.050 22.985 34.610 ;
        RECT 23.775 34.050 23.945 34.610 ;
        RECT 24.735 34.050 24.905 34.610 ;
        RECT 19.935 29.675 20.105 31.075 ;
        RECT 20.895 29.675 21.065 31.075 ;
        RECT 21.855 29.675 22.025 31.075 ;
        RECT 22.815 29.675 22.985 31.075 ;
        RECT 23.775 29.675 23.945 31.075 ;
        RECT 24.735 29.675 24.905 31.075 ;
        RECT 19.935 27.615 20.105 28.175 ;
        RECT 20.895 27.615 21.065 28.175 ;
        RECT 21.855 27.615 22.025 28.175 ;
        RECT 22.815 27.615 22.985 28.175 ;
        RECT 23.775 27.615 23.945 28.175 ;
        RECT 24.735 27.615 24.905 28.175 ;
        RECT 19.935 23.240 20.105 24.640 ;
        RECT 20.895 23.240 21.065 24.640 ;
        RECT 21.855 23.240 22.025 24.640 ;
        RECT 22.815 23.240 22.985 24.640 ;
        RECT 23.775 23.240 23.945 24.640 ;
        RECT 24.735 23.240 24.905 24.640 ;
        RECT 19.935 21.180 20.105 21.740 ;
        RECT 20.895 21.180 21.065 21.740 ;
        RECT 21.855 21.180 22.025 21.740 ;
        RECT 22.815 21.180 22.985 21.740 ;
        RECT 23.775 21.180 23.945 21.740 ;
        RECT 24.735 21.180 24.905 21.740 ;
        RECT 19.935 16.805 20.105 18.205 ;
        RECT 20.895 16.805 21.065 18.205 ;
        RECT 21.855 16.805 22.025 18.205 ;
        RECT 22.815 16.805 22.985 18.205 ;
        RECT 23.775 16.805 23.945 18.205 ;
        RECT 24.735 16.805 24.905 18.205 ;
        RECT 19.935 14.745 20.105 15.305 ;
        RECT 20.895 14.745 21.065 15.305 ;
        RECT 21.855 14.745 22.025 15.305 ;
        RECT 22.815 14.745 22.985 15.305 ;
        RECT 23.775 14.745 23.945 15.305 ;
        RECT 24.735 14.745 24.905 15.305 ;
        RECT 19.935 10.370 20.105 11.770 ;
        RECT 20.895 10.370 21.065 11.770 ;
        RECT 21.855 10.370 22.025 11.770 ;
        RECT 22.815 10.370 22.985 11.770 ;
        RECT 23.775 10.370 23.945 11.770 ;
        RECT 24.735 10.370 24.905 11.770 ;
        RECT 19.935 8.310 20.105 8.870 ;
        RECT 20.895 8.310 21.065 8.870 ;
        RECT 21.855 8.310 22.025 8.870 ;
        RECT 22.815 8.310 22.985 8.870 ;
        RECT 23.775 8.310 23.945 8.870 ;
        RECT 24.735 8.310 24.905 8.870 ;
        RECT 19.935 3.935 20.105 5.335 ;
        RECT 20.895 3.935 21.065 5.335 ;
        RECT 21.855 3.935 22.025 5.335 ;
        RECT 22.815 3.935 22.985 5.335 ;
        RECT 23.775 3.935 23.945 5.335 ;
        RECT 24.735 3.935 24.905 5.335 ;
        RECT 19.935 1.875 20.105 2.435 ;
        RECT 20.895 1.875 21.065 2.435 ;
        RECT 21.855 1.875 22.025 2.435 ;
        RECT 22.815 1.875 22.985 2.435 ;
        RECT 23.775 1.875 23.945 2.435 ;
        RECT 24.735 1.875 24.905 2.435 ;
      LAYER mcon ;
        RECT 19.935 204.395 20.105 204.565 ;
        RECT 19.935 204.035 20.105 204.205 ;
        RECT 19.935 203.675 20.105 203.845 ;
        RECT 20.895 204.395 21.065 204.565 ;
        RECT 20.895 204.035 21.065 204.205 ;
        RECT 20.895 203.675 21.065 203.845 ;
        RECT 21.855 204.395 22.025 204.565 ;
        RECT 21.855 204.035 22.025 204.205 ;
        RECT 21.855 203.675 22.025 203.845 ;
        RECT 22.815 204.395 22.985 204.565 ;
        RECT 22.815 204.035 22.985 204.205 ;
        RECT 22.815 203.675 22.985 203.845 ;
        RECT 23.775 204.395 23.945 204.565 ;
        RECT 23.775 204.035 23.945 204.205 ;
        RECT 23.775 203.675 23.945 203.845 ;
        RECT 24.735 204.395 24.905 204.565 ;
        RECT 24.735 204.035 24.905 204.205 ;
        RECT 24.735 203.675 24.905 203.845 ;
        RECT 19.935 201.555 20.105 201.725 ;
        RECT 20.895 201.555 21.065 201.725 ;
        RECT 21.855 201.555 22.025 201.725 ;
        RECT 22.815 201.555 22.985 201.725 ;
        RECT 23.775 201.555 23.945 201.725 ;
        RECT 24.735 201.555 24.905 201.725 ;
        RECT 19.935 197.960 20.105 198.130 ;
        RECT 19.935 197.600 20.105 197.770 ;
        RECT 19.935 197.240 20.105 197.410 ;
        RECT 20.895 197.960 21.065 198.130 ;
        RECT 20.895 197.600 21.065 197.770 ;
        RECT 20.895 197.240 21.065 197.410 ;
        RECT 21.855 197.960 22.025 198.130 ;
        RECT 21.855 197.600 22.025 197.770 ;
        RECT 21.855 197.240 22.025 197.410 ;
        RECT 22.815 197.960 22.985 198.130 ;
        RECT 22.815 197.600 22.985 197.770 ;
        RECT 22.815 197.240 22.985 197.410 ;
        RECT 23.775 197.960 23.945 198.130 ;
        RECT 23.775 197.600 23.945 197.770 ;
        RECT 23.775 197.240 23.945 197.410 ;
        RECT 24.735 197.960 24.905 198.130 ;
        RECT 24.735 197.600 24.905 197.770 ;
        RECT 24.735 197.240 24.905 197.410 ;
        RECT 19.935 195.120 20.105 195.290 ;
        RECT 20.895 195.120 21.065 195.290 ;
        RECT 21.855 195.120 22.025 195.290 ;
        RECT 22.815 195.120 22.985 195.290 ;
        RECT 23.775 195.120 23.945 195.290 ;
        RECT 24.735 195.120 24.905 195.290 ;
        RECT 19.935 191.525 20.105 191.695 ;
        RECT 19.935 191.165 20.105 191.335 ;
        RECT 19.935 190.805 20.105 190.975 ;
        RECT 20.895 191.525 21.065 191.695 ;
        RECT 20.895 191.165 21.065 191.335 ;
        RECT 20.895 190.805 21.065 190.975 ;
        RECT 21.855 191.525 22.025 191.695 ;
        RECT 21.855 191.165 22.025 191.335 ;
        RECT 21.855 190.805 22.025 190.975 ;
        RECT 22.815 191.525 22.985 191.695 ;
        RECT 22.815 191.165 22.985 191.335 ;
        RECT 22.815 190.805 22.985 190.975 ;
        RECT 23.775 191.525 23.945 191.695 ;
        RECT 23.775 191.165 23.945 191.335 ;
        RECT 23.775 190.805 23.945 190.975 ;
        RECT 24.735 191.525 24.905 191.695 ;
        RECT 24.735 191.165 24.905 191.335 ;
        RECT 24.735 190.805 24.905 190.975 ;
        RECT 19.935 188.685 20.105 188.855 ;
        RECT 20.895 188.685 21.065 188.855 ;
        RECT 21.855 188.685 22.025 188.855 ;
        RECT 22.815 188.685 22.985 188.855 ;
        RECT 23.775 188.685 23.945 188.855 ;
        RECT 24.735 188.685 24.905 188.855 ;
        RECT 19.935 185.090 20.105 185.260 ;
        RECT 19.935 184.730 20.105 184.900 ;
        RECT 19.935 184.370 20.105 184.540 ;
        RECT 20.895 185.090 21.065 185.260 ;
        RECT 20.895 184.730 21.065 184.900 ;
        RECT 20.895 184.370 21.065 184.540 ;
        RECT 21.855 185.090 22.025 185.260 ;
        RECT 21.855 184.730 22.025 184.900 ;
        RECT 21.855 184.370 22.025 184.540 ;
        RECT 22.815 185.090 22.985 185.260 ;
        RECT 22.815 184.730 22.985 184.900 ;
        RECT 22.815 184.370 22.985 184.540 ;
        RECT 23.775 185.090 23.945 185.260 ;
        RECT 23.775 184.730 23.945 184.900 ;
        RECT 23.775 184.370 23.945 184.540 ;
        RECT 24.735 185.090 24.905 185.260 ;
        RECT 24.735 184.730 24.905 184.900 ;
        RECT 24.735 184.370 24.905 184.540 ;
        RECT 19.935 182.250 20.105 182.420 ;
        RECT 20.895 182.250 21.065 182.420 ;
        RECT 21.855 182.250 22.025 182.420 ;
        RECT 22.815 182.250 22.985 182.420 ;
        RECT 23.775 182.250 23.945 182.420 ;
        RECT 24.735 182.250 24.905 182.420 ;
        RECT 19.935 178.655 20.105 178.825 ;
        RECT 19.935 178.295 20.105 178.465 ;
        RECT 19.935 177.935 20.105 178.105 ;
        RECT 20.895 178.655 21.065 178.825 ;
        RECT 20.895 178.295 21.065 178.465 ;
        RECT 20.895 177.935 21.065 178.105 ;
        RECT 21.855 178.655 22.025 178.825 ;
        RECT 21.855 178.295 22.025 178.465 ;
        RECT 21.855 177.935 22.025 178.105 ;
        RECT 22.815 178.655 22.985 178.825 ;
        RECT 22.815 178.295 22.985 178.465 ;
        RECT 22.815 177.935 22.985 178.105 ;
        RECT 23.775 178.655 23.945 178.825 ;
        RECT 23.775 178.295 23.945 178.465 ;
        RECT 23.775 177.935 23.945 178.105 ;
        RECT 24.735 178.655 24.905 178.825 ;
        RECT 24.735 178.295 24.905 178.465 ;
        RECT 24.735 177.935 24.905 178.105 ;
        RECT 19.935 175.815 20.105 175.985 ;
        RECT 20.895 175.815 21.065 175.985 ;
        RECT 21.855 175.815 22.025 175.985 ;
        RECT 22.815 175.815 22.985 175.985 ;
        RECT 23.775 175.815 23.945 175.985 ;
        RECT 24.735 175.815 24.905 175.985 ;
        RECT 19.935 172.220 20.105 172.390 ;
        RECT 19.935 171.860 20.105 172.030 ;
        RECT 19.935 171.500 20.105 171.670 ;
        RECT 20.895 172.220 21.065 172.390 ;
        RECT 20.895 171.860 21.065 172.030 ;
        RECT 20.895 171.500 21.065 171.670 ;
        RECT 21.855 172.220 22.025 172.390 ;
        RECT 21.855 171.860 22.025 172.030 ;
        RECT 21.855 171.500 22.025 171.670 ;
        RECT 22.815 172.220 22.985 172.390 ;
        RECT 22.815 171.860 22.985 172.030 ;
        RECT 22.815 171.500 22.985 171.670 ;
        RECT 23.775 172.220 23.945 172.390 ;
        RECT 23.775 171.860 23.945 172.030 ;
        RECT 23.775 171.500 23.945 171.670 ;
        RECT 24.735 172.220 24.905 172.390 ;
        RECT 24.735 171.860 24.905 172.030 ;
        RECT 24.735 171.500 24.905 171.670 ;
        RECT 19.935 169.380 20.105 169.550 ;
        RECT 20.895 169.380 21.065 169.550 ;
        RECT 21.855 169.380 22.025 169.550 ;
        RECT 22.815 169.380 22.985 169.550 ;
        RECT 23.775 169.380 23.945 169.550 ;
        RECT 24.735 169.380 24.905 169.550 ;
        RECT 19.935 165.785 20.105 165.955 ;
        RECT 19.935 165.425 20.105 165.595 ;
        RECT 19.935 165.065 20.105 165.235 ;
        RECT 20.895 165.785 21.065 165.955 ;
        RECT 20.895 165.425 21.065 165.595 ;
        RECT 20.895 165.065 21.065 165.235 ;
        RECT 21.855 165.785 22.025 165.955 ;
        RECT 21.855 165.425 22.025 165.595 ;
        RECT 21.855 165.065 22.025 165.235 ;
        RECT 22.815 165.785 22.985 165.955 ;
        RECT 22.815 165.425 22.985 165.595 ;
        RECT 22.815 165.065 22.985 165.235 ;
        RECT 23.775 165.785 23.945 165.955 ;
        RECT 23.775 165.425 23.945 165.595 ;
        RECT 23.775 165.065 23.945 165.235 ;
        RECT 24.735 165.785 24.905 165.955 ;
        RECT 24.735 165.425 24.905 165.595 ;
        RECT 24.735 165.065 24.905 165.235 ;
        RECT 19.935 162.945 20.105 163.115 ;
        RECT 20.895 162.945 21.065 163.115 ;
        RECT 21.855 162.945 22.025 163.115 ;
        RECT 22.815 162.945 22.985 163.115 ;
        RECT 23.775 162.945 23.945 163.115 ;
        RECT 24.735 162.945 24.905 163.115 ;
        RECT 19.935 159.350 20.105 159.520 ;
        RECT 19.935 158.990 20.105 159.160 ;
        RECT 19.935 158.630 20.105 158.800 ;
        RECT 20.895 159.350 21.065 159.520 ;
        RECT 20.895 158.990 21.065 159.160 ;
        RECT 20.895 158.630 21.065 158.800 ;
        RECT 21.855 159.350 22.025 159.520 ;
        RECT 21.855 158.990 22.025 159.160 ;
        RECT 21.855 158.630 22.025 158.800 ;
        RECT 22.815 159.350 22.985 159.520 ;
        RECT 22.815 158.990 22.985 159.160 ;
        RECT 22.815 158.630 22.985 158.800 ;
        RECT 23.775 159.350 23.945 159.520 ;
        RECT 23.775 158.990 23.945 159.160 ;
        RECT 23.775 158.630 23.945 158.800 ;
        RECT 24.735 159.350 24.905 159.520 ;
        RECT 24.735 158.990 24.905 159.160 ;
        RECT 24.735 158.630 24.905 158.800 ;
        RECT 19.935 156.510 20.105 156.680 ;
        RECT 20.895 156.510 21.065 156.680 ;
        RECT 21.855 156.510 22.025 156.680 ;
        RECT 22.815 156.510 22.985 156.680 ;
        RECT 23.775 156.510 23.945 156.680 ;
        RECT 24.735 156.510 24.905 156.680 ;
        RECT 19.935 152.915 20.105 153.085 ;
        RECT 19.935 152.555 20.105 152.725 ;
        RECT 19.935 152.195 20.105 152.365 ;
        RECT 20.895 152.915 21.065 153.085 ;
        RECT 20.895 152.555 21.065 152.725 ;
        RECT 20.895 152.195 21.065 152.365 ;
        RECT 21.855 152.915 22.025 153.085 ;
        RECT 21.855 152.555 22.025 152.725 ;
        RECT 21.855 152.195 22.025 152.365 ;
        RECT 22.815 152.915 22.985 153.085 ;
        RECT 22.815 152.555 22.985 152.725 ;
        RECT 22.815 152.195 22.985 152.365 ;
        RECT 23.775 152.915 23.945 153.085 ;
        RECT 23.775 152.555 23.945 152.725 ;
        RECT 23.775 152.195 23.945 152.365 ;
        RECT 24.735 152.915 24.905 153.085 ;
        RECT 24.735 152.555 24.905 152.725 ;
        RECT 24.735 152.195 24.905 152.365 ;
        RECT 19.935 150.075 20.105 150.245 ;
        RECT 20.895 150.075 21.065 150.245 ;
        RECT 21.855 150.075 22.025 150.245 ;
        RECT 22.815 150.075 22.985 150.245 ;
        RECT 23.775 150.075 23.945 150.245 ;
        RECT 24.735 150.075 24.905 150.245 ;
        RECT 19.935 146.480 20.105 146.650 ;
        RECT 19.935 146.120 20.105 146.290 ;
        RECT 19.935 145.760 20.105 145.930 ;
        RECT 20.895 146.480 21.065 146.650 ;
        RECT 20.895 146.120 21.065 146.290 ;
        RECT 20.895 145.760 21.065 145.930 ;
        RECT 21.855 146.480 22.025 146.650 ;
        RECT 21.855 146.120 22.025 146.290 ;
        RECT 21.855 145.760 22.025 145.930 ;
        RECT 22.815 146.480 22.985 146.650 ;
        RECT 22.815 146.120 22.985 146.290 ;
        RECT 22.815 145.760 22.985 145.930 ;
        RECT 23.775 146.480 23.945 146.650 ;
        RECT 23.775 146.120 23.945 146.290 ;
        RECT 23.775 145.760 23.945 145.930 ;
        RECT 24.735 146.480 24.905 146.650 ;
        RECT 24.735 146.120 24.905 146.290 ;
        RECT 24.735 145.760 24.905 145.930 ;
        RECT 19.935 143.640 20.105 143.810 ;
        RECT 20.895 143.640 21.065 143.810 ;
        RECT 21.855 143.640 22.025 143.810 ;
        RECT 22.815 143.640 22.985 143.810 ;
        RECT 23.775 143.640 23.945 143.810 ;
        RECT 24.735 143.640 24.905 143.810 ;
        RECT 19.935 140.045 20.105 140.215 ;
        RECT 19.935 139.685 20.105 139.855 ;
        RECT 19.935 139.325 20.105 139.495 ;
        RECT 20.895 140.045 21.065 140.215 ;
        RECT 20.895 139.685 21.065 139.855 ;
        RECT 20.895 139.325 21.065 139.495 ;
        RECT 21.855 140.045 22.025 140.215 ;
        RECT 21.855 139.685 22.025 139.855 ;
        RECT 21.855 139.325 22.025 139.495 ;
        RECT 22.815 140.045 22.985 140.215 ;
        RECT 22.815 139.685 22.985 139.855 ;
        RECT 22.815 139.325 22.985 139.495 ;
        RECT 23.775 140.045 23.945 140.215 ;
        RECT 23.775 139.685 23.945 139.855 ;
        RECT 23.775 139.325 23.945 139.495 ;
        RECT 24.735 140.045 24.905 140.215 ;
        RECT 24.735 139.685 24.905 139.855 ;
        RECT 24.735 139.325 24.905 139.495 ;
        RECT 19.935 137.205 20.105 137.375 ;
        RECT 20.895 137.205 21.065 137.375 ;
        RECT 21.855 137.205 22.025 137.375 ;
        RECT 22.815 137.205 22.985 137.375 ;
        RECT 23.775 137.205 23.945 137.375 ;
        RECT 24.735 137.205 24.905 137.375 ;
        RECT 19.935 133.610 20.105 133.780 ;
        RECT 19.935 133.250 20.105 133.420 ;
        RECT 19.935 132.890 20.105 133.060 ;
        RECT 20.895 133.610 21.065 133.780 ;
        RECT 20.895 133.250 21.065 133.420 ;
        RECT 20.895 132.890 21.065 133.060 ;
        RECT 21.855 133.610 22.025 133.780 ;
        RECT 21.855 133.250 22.025 133.420 ;
        RECT 21.855 132.890 22.025 133.060 ;
        RECT 22.815 133.610 22.985 133.780 ;
        RECT 22.815 133.250 22.985 133.420 ;
        RECT 22.815 132.890 22.985 133.060 ;
        RECT 23.775 133.610 23.945 133.780 ;
        RECT 23.775 133.250 23.945 133.420 ;
        RECT 23.775 132.890 23.945 133.060 ;
        RECT 24.735 133.610 24.905 133.780 ;
        RECT 24.735 133.250 24.905 133.420 ;
        RECT 24.735 132.890 24.905 133.060 ;
        RECT 19.935 130.770 20.105 130.940 ;
        RECT 20.895 130.770 21.065 130.940 ;
        RECT 21.855 130.770 22.025 130.940 ;
        RECT 22.815 130.770 22.985 130.940 ;
        RECT 23.775 130.770 23.945 130.940 ;
        RECT 24.735 130.770 24.905 130.940 ;
        RECT 19.935 127.175 20.105 127.345 ;
        RECT 19.935 126.815 20.105 126.985 ;
        RECT 19.935 126.455 20.105 126.625 ;
        RECT 20.895 127.175 21.065 127.345 ;
        RECT 20.895 126.815 21.065 126.985 ;
        RECT 20.895 126.455 21.065 126.625 ;
        RECT 21.855 127.175 22.025 127.345 ;
        RECT 21.855 126.815 22.025 126.985 ;
        RECT 21.855 126.455 22.025 126.625 ;
        RECT 22.815 127.175 22.985 127.345 ;
        RECT 22.815 126.815 22.985 126.985 ;
        RECT 22.815 126.455 22.985 126.625 ;
        RECT 23.775 127.175 23.945 127.345 ;
        RECT 23.775 126.815 23.945 126.985 ;
        RECT 23.775 126.455 23.945 126.625 ;
        RECT 24.735 127.175 24.905 127.345 ;
        RECT 24.735 126.815 24.905 126.985 ;
        RECT 24.735 126.455 24.905 126.625 ;
        RECT 19.935 124.335 20.105 124.505 ;
        RECT 20.895 124.335 21.065 124.505 ;
        RECT 21.855 124.335 22.025 124.505 ;
        RECT 22.815 124.335 22.985 124.505 ;
        RECT 23.775 124.335 23.945 124.505 ;
        RECT 24.735 124.335 24.905 124.505 ;
        RECT 19.935 120.740 20.105 120.910 ;
        RECT 19.935 120.380 20.105 120.550 ;
        RECT 19.935 120.020 20.105 120.190 ;
        RECT 20.895 120.740 21.065 120.910 ;
        RECT 20.895 120.380 21.065 120.550 ;
        RECT 20.895 120.020 21.065 120.190 ;
        RECT 21.855 120.740 22.025 120.910 ;
        RECT 21.855 120.380 22.025 120.550 ;
        RECT 21.855 120.020 22.025 120.190 ;
        RECT 22.815 120.740 22.985 120.910 ;
        RECT 22.815 120.380 22.985 120.550 ;
        RECT 22.815 120.020 22.985 120.190 ;
        RECT 23.775 120.740 23.945 120.910 ;
        RECT 23.775 120.380 23.945 120.550 ;
        RECT 23.775 120.020 23.945 120.190 ;
        RECT 24.735 120.740 24.905 120.910 ;
        RECT 24.735 120.380 24.905 120.550 ;
        RECT 24.735 120.020 24.905 120.190 ;
        RECT 19.935 117.900 20.105 118.070 ;
        RECT 20.895 117.900 21.065 118.070 ;
        RECT 21.855 117.900 22.025 118.070 ;
        RECT 22.815 117.900 22.985 118.070 ;
        RECT 23.775 117.900 23.945 118.070 ;
        RECT 24.735 117.900 24.905 118.070 ;
        RECT 19.935 114.305 20.105 114.475 ;
        RECT 19.935 113.945 20.105 114.115 ;
        RECT 19.935 113.585 20.105 113.755 ;
        RECT 20.895 114.305 21.065 114.475 ;
        RECT 20.895 113.945 21.065 114.115 ;
        RECT 20.895 113.585 21.065 113.755 ;
        RECT 21.855 114.305 22.025 114.475 ;
        RECT 21.855 113.945 22.025 114.115 ;
        RECT 21.855 113.585 22.025 113.755 ;
        RECT 22.815 114.305 22.985 114.475 ;
        RECT 22.815 113.945 22.985 114.115 ;
        RECT 22.815 113.585 22.985 113.755 ;
        RECT 23.775 114.305 23.945 114.475 ;
        RECT 23.775 113.945 23.945 114.115 ;
        RECT 23.775 113.585 23.945 113.755 ;
        RECT 24.735 114.305 24.905 114.475 ;
        RECT 24.735 113.945 24.905 114.115 ;
        RECT 24.735 113.585 24.905 113.755 ;
        RECT 19.935 111.465 20.105 111.635 ;
        RECT 20.895 111.465 21.065 111.635 ;
        RECT 21.855 111.465 22.025 111.635 ;
        RECT 22.815 111.465 22.985 111.635 ;
        RECT 23.775 111.465 23.945 111.635 ;
        RECT 24.735 111.465 24.905 111.635 ;
        RECT 19.935 107.870 20.105 108.040 ;
        RECT 19.935 107.510 20.105 107.680 ;
        RECT 19.935 107.150 20.105 107.320 ;
        RECT 20.895 107.870 21.065 108.040 ;
        RECT 20.895 107.510 21.065 107.680 ;
        RECT 20.895 107.150 21.065 107.320 ;
        RECT 21.855 107.870 22.025 108.040 ;
        RECT 21.855 107.510 22.025 107.680 ;
        RECT 21.855 107.150 22.025 107.320 ;
        RECT 22.815 107.870 22.985 108.040 ;
        RECT 22.815 107.510 22.985 107.680 ;
        RECT 22.815 107.150 22.985 107.320 ;
        RECT 23.775 107.870 23.945 108.040 ;
        RECT 23.775 107.510 23.945 107.680 ;
        RECT 23.775 107.150 23.945 107.320 ;
        RECT 24.735 107.870 24.905 108.040 ;
        RECT 24.735 107.510 24.905 107.680 ;
        RECT 24.735 107.150 24.905 107.320 ;
        RECT 19.935 105.030 20.105 105.200 ;
        RECT 20.895 105.030 21.065 105.200 ;
        RECT 21.855 105.030 22.025 105.200 ;
        RECT 22.815 105.030 22.985 105.200 ;
        RECT 23.775 105.030 23.945 105.200 ;
        RECT 24.735 105.030 24.905 105.200 ;
        RECT 19.935 101.435 20.105 101.605 ;
        RECT 19.935 101.075 20.105 101.245 ;
        RECT 19.935 100.715 20.105 100.885 ;
        RECT 20.895 101.435 21.065 101.605 ;
        RECT 20.895 101.075 21.065 101.245 ;
        RECT 20.895 100.715 21.065 100.885 ;
        RECT 21.855 101.435 22.025 101.605 ;
        RECT 21.855 101.075 22.025 101.245 ;
        RECT 21.855 100.715 22.025 100.885 ;
        RECT 22.815 101.435 22.985 101.605 ;
        RECT 22.815 101.075 22.985 101.245 ;
        RECT 22.815 100.715 22.985 100.885 ;
        RECT 23.775 101.435 23.945 101.605 ;
        RECT 23.775 101.075 23.945 101.245 ;
        RECT 23.775 100.715 23.945 100.885 ;
        RECT 24.735 101.435 24.905 101.605 ;
        RECT 24.735 101.075 24.905 101.245 ;
        RECT 24.735 100.715 24.905 100.885 ;
        RECT 19.935 98.595 20.105 98.765 ;
        RECT 20.895 98.595 21.065 98.765 ;
        RECT 21.855 98.595 22.025 98.765 ;
        RECT 22.815 98.595 22.985 98.765 ;
        RECT 23.775 98.595 23.945 98.765 ;
        RECT 24.735 98.595 24.905 98.765 ;
        RECT 19.935 95.000 20.105 95.170 ;
        RECT 19.935 94.640 20.105 94.810 ;
        RECT 19.935 94.280 20.105 94.450 ;
        RECT 20.895 95.000 21.065 95.170 ;
        RECT 20.895 94.640 21.065 94.810 ;
        RECT 20.895 94.280 21.065 94.450 ;
        RECT 21.855 95.000 22.025 95.170 ;
        RECT 21.855 94.640 22.025 94.810 ;
        RECT 21.855 94.280 22.025 94.450 ;
        RECT 22.815 95.000 22.985 95.170 ;
        RECT 22.815 94.640 22.985 94.810 ;
        RECT 22.815 94.280 22.985 94.450 ;
        RECT 23.775 95.000 23.945 95.170 ;
        RECT 23.775 94.640 23.945 94.810 ;
        RECT 23.775 94.280 23.945 94.450 ;
        RECT 24.735 95.000 24.905 95.170 ;
        RECT 24.735 94.640 24.905 94.810 ;
        RECT 24.735 94.280 24.905 94.450 ;
        RECT 19.935 92.160 20.105 92.330 ;
        RECT 20.895 92.160 21.065 92.330 ;
        RECT 21.855 92.160 22.025 92.330 ;
        RECT 22.815 92.160 22.985 92.330 ;
        RECT 23.775 92.160 23.945 92.330 ;
        RECT 24.735 92.160 24.905 92.330 ;
        RECT 19.935 88.565 20.105 88.735 ;
        RECT 19.935 88.205 20.105 88.375 ;
        RECT 19.935 87.845 20.105 88.015 ;
        RECT 20.895 88.565 21.065 88.735 ;
        RECT 20.895 88.205 21.065 88.375 ;
        RECT 20.895 87.845 21.065 88.015 ;
        RECT 21.855 88.565 22.025 88.735 ;
        RECT 21.855 88.205 22.025 88.375 ;
        RECT 21.855 87.845 22.025 88.015 ;
        RECT 22.815 88.565 22.985 88.735 ;
        RECT 22.815 88.205 22.985 88.375 ;
        RECT 22.815 87.845 22.985 88.015 ;
        RECT 23.775 88.565 23.945 88.735 ;
        RECT 23.775 88.205 23.945 88.375 ;
        RECT 23.775 87.845 23.945 88.015 ;
        RECT 24.735 88.565 24.905 88.735 ;
        RECT 24.735 88.205 24.905 88.375 ;
        RECT 24.735 87.845 24.905 88.015 ;
        RECT 19.935 85.725 20.105 85.895 ;
        RECT 20.895 85.725 21.065 85.895 ;
        RECT 21.855 85.725 22.025 85.895 ;
        RECT 22.815 85.725 22.985 85.895 ;
        RECT 23.775 85.725 23.945 85.895 ;
        RECT 24.735 85.725 24.905 85.895 ;
        RECT 19.935 82.130 20.105 82.300 ;
        RECT 19.935 81.770 20.105 81.940 ;
        RECT 19.935 81.410 20.105 81.580 ;
        RECT 20.895 82.130 21.065 82.300 ;
        RECT 20.895 81.770 21.065 81.940 ;
        RECT 20.895 81.410 21.065 81.580 ;
        RECT 21.855 82.130 22.025 82.300 ;
        RECT 21.855 81.770 22.025 81.940 ;
        RECT 21.855 81.410 22.025 81.580 ;
        RECT 22.815 82.130 22.985 82.300 ;
        RECT 22.815 81.770 22.985 81.940 ;
        RECT 22.815 81.410 22.985 81.580 ;
        RECT 23.775 82.130 23.945 82.300 ;
        RECT 23.775 81.770 23.945 81.940 ;
        RECT 23.775 81.410 23.945 81.580 ;
        RECT 24.735 82.130 24.905 82.300 ;
        RECT 24.735 81.770 24.905 81.940 ;
        RECT 24.735 81.410 24.905 81.580 ;
        RECT 19.935 79.290 20.105 79.460 ;
        RECT 20.895 79.290 21.065 79.460 ;
        RECT 21.855 79.290 22.025 79.460 ;
        RECT 22.815 79.290 22.985 79.460 ;
        RECT 23.775 79.290 23.945 79.460 ;
        RECT 24.735 79.290 24.905 79.460 ;
        RECT 19.935 75.695 20.105 75.865 ;
        RECT 19.935 75.335 20.105 75.505 ;
        RECT 19.935 74.975 20.105 75.145 ;
        RECT 20.895 75.695 21.065 75.865 ;
        RECT 20.895 75.335 21.065 75.505 ;
        RECT 20.895 74.975 21.065 75.145 ;
        RECT 21.855 75.695 22.025 75.865 ;
        RECT 21.855 75.335 22.025 75.505 ;
        RECT 21.855 74.975 22.025 75.145 ;
        RECT 22.815 75.695 22.985 75.865 ;
        RECT 22.815 75.335 22.985 75.505 ;
        RECT 22.815 74.975 22.985 75.145 ;
        RECT 23.775 75.695 23.945 75.865 ;
        RECT 23.775 75.335 23.945 75.505 ;
        RECT 23.775 74.975 23.945 75.145 ;
        RECT 24.735 75.695 24.905 75.865 ;
        RECT 24.735 75.335 24.905 75.505 ;
        RECT 24.735 74.975 24.905 75.145 ;
        RECT 19.935 72.855 20.105 73.025 ;
        RECT 20.895 72.855 21.065 73.025 ;
        RECT 21.855 72.855 22.025 73.025 ;
        RECT 22.815 72.855 22.985 73.025 ;
        RECT 23.775 72.855 23.945 73.025 ;
        RECT 24.735 72.855 24.905 73.025 ;
        RECT 19.935 69.260 20.105 69.430 ;
        RECT 19.935 68.900 20.105 69.070 ;
        RECT 19.935 68.540 20.105 68.710 ;
        RECT 20.895 69.260 21.065 69.430 ;
        RECT 20.895 68.900 21.065 69.070 ;
        RECT 20.895 68.540 21.065 68.710 ;
        RECT 21.855 69.260 22.025 69.430 ;
        RECT 21.855 68.900 22.025 69.070 ;
        RECT 21.855 68.540 22.025 68.710 ;
        RECT 22.815 69.260 22.985 69.430 ;
        RECT 22.815 68.900 22.985 69.070 ;
        RECT 22.815 68.540 22.985 68.710 ;
        RECT 23.775 69.260 23.945 69.430 ;
        RECT 23.775 68.900 23.945 69.070 ;
        RECT 23.775 68.540 23.945 68.710 ;
        RECT 24.735 69.260 24.905 69.430 ;
        RECT 24.735 68.900 24.905 69.070 ;
        RECT 24.735 68.540 24.905 68.710 ;
        RECT 19.935 66.420 20.105 66.590 ;
        RECT 20.895 66.420 21.065 66.590 ;
        RECT 21.855 66.420 22.025 66.590 ;
        RECT 22.815 66.420 22.985 66.590 ;
        RECT 23.775 66.420 23.945 66.590 ;
        RECT 24.735 66.420 24.905 66.590 ;
        RECT 19.935 62.825 20.105 62.995 ;
        RECT 19.935 62.465 20.105 62.635 ;
        RECT 19.935 62.105 20.105 62.275 ;
        RECT 20.895 62.825 21.065 62.995 ;
        RECT 20.895 62.465 21.065 62.635 ;
        RECT 20.895 62.105 21.065 62.275 ;
        RECT 21.855 62.825 22.025 62.995 ;
        RECT 21.855 62.465 22.025 62.635 ;
        RECT 21.855 62.105 22.025 62.275 ;
        RECT 22.815 62.825 22.985 62.995 ;
        RECT 22.815 62.465 22.985 62.635 ;
        RECT 22.815 62.105 22.985 62.275 ;
        RECT 23.775 62.825 23.945 62.995 ;
        RECT 23.775 62.465 23.945 62.635 ;
        RECT 23.775 62.105 23.945 62.275 ;
        RECT 24.735 62.825 24.905 62.995 ;
        RECT 24.735 62.465 24.905 62.635 ;
        RECT 24.735 62.105 24.905 62.275 ;
        RECT 19.935 59.985 20.105 60.155 ;
        RECT 20.895 59.985 21.065 60.155 ;
        RECT 21.855 59.985 22.025 60.155 ;
        RECT 22.815 59.985 22.985 60.155 ;
        RECT 23.775 59.985 23.945 60.155 ;
        RECT 24.735 59.985 24.905 60.155 ;
        RECT 19.935 56.390 20.105 56.560 ;
        RECT 19.935 56.030 20.105 56.200 ;
        RECT 19.935 55.670 20.105 55.840 ;
        RECT 20.895 56.390 21.065 56.560 ;
        RECT 20.895 56.030 21.065 56.200 ;
        RECT 20.895 55.670 21.065 55.840 ;
        RECT 21.855 56.390 22.025 56.560 ;
        RECT 21.855 56.030 22.025 56.200 ;
        RECT 21.855 55.670 22.025 55.840 ;
        RECT 22.815 56.390 22.985 56.560 ;
        RECT 22.815 56.030 22.985 56.200 ;
        RECT 22.815 55.670 22.985 55.840 ;
        RECT 23.775 56.390 23.945 56.560 ;
        RECT 23.775 56.030 23.945 56.200 ;
        RECT 23.775 55.670 23.945 55.840 ;
        RECT 24.735 56.390 24.905 56.560 ;
        RECT 24.735 56.030 24.905 56.200 ;
        RECT 24.735 55.670 24.905 55.840 ;
        RECT 19.935 53.550 20.105 53.720 ;
        RECT 20.895 53.550 21.065 53.720 ;
        RECT 21.855 53.550 22.025 53.720 ;
        RECT 22.815 53.550 22.985 53.720 ;
        RECT 23.775 53.550 23.945 53.720 ;
        RECT 24.735 53.550 24.905 53.720 ;
        RECT 19.935 49.955 20.105 50.125 ;
        RECT 19.935 49.595 20.105 49.765 ;
        RECT 19.935 49.235 20.105 49.405 ;
        RECT 20.895 49.955 21.065 50.125 ;
        RECT 20.895 49.595 21.065 49.765 ;
        RECT 20.895 49.235 21.065 49.405 ;
        RECT 21.855 49.955 22.025 50.125 ;
        RECT 21.855 49.595 22.025 49.765 ;
        RECT 21.855 49.235 22.025 49.405 ;
        RECT 22.815 49.955 22.985 50.125 ;
        RECT 22.815 49.595 22.985 49.765 ;
        RECT 22.815 49.235 22.985 49.405 ;
        RECT 23.775 49.955 23.945 50.125 ;
        RECT 23.775 49.595 23.945 49.765 ;
        RECT 23.775 49.235 23.945 49.405 ;
        RECT 24.735 49.955 24.905 50.125 ;
        RECT 24.735 49.595 24.905 49.765 ;
        RECT 24.735 49.235 24.905 49.405 ;
        RECT 19.935 47.115 20.105 47.285 ;
        RECT 20.895 47.115 21.065 47.285 ;
        RECT 21.855 47.115 22.025 47.285 ;
        RECT 22.815 47.115 22.985 47.285 ;
        RECT 23.775 47.115 23.945 47.285 ;
        RECT 24.735 47.115 24.905 47.285 ;
        RECT 19.935 43.520 20.105 43.690 ;
        RECT 19.935 43.160 20.105 43.330 ;
        RECT 19.935 42.800 20.105 42.970 ;
        RECT 20.895 43.520 21.065 43.690 ;
        RECT 20.895 43.160 21.065 43.330 ;
        RECT 20.895 42.800 21.065 42.970 ;
        RECT 21.855 43.520 22.025 43.690 ;
        RECT 21.855 43.160 22.025 43.330 ;
        RECT 21.855 42.800 22.025 42.970 ;
        RECT 22.815 43.520 22.985 43.690 ;
        RECT 22.815 43.160 22.985 43.330 ;
        RECT 22.815 42.800 22.985 42.970 ;
        RECT 23.775 43.520 23.945 43.690 ;
        RECT 23.775 43.160 23.945 43.330 ;
        RECT 23.775 42.800 23.945 42.970 ;
        RECT 24.735 43.520 24.905 43.690 ;
        RECT 24.735 43.160 24.905 43.330 ;
        RECT 24.735 42.800 24.905 42.970 ;
        RECT 19.935 40.680 20.105 40.850 ;
        RECT 20.895 40.680 21.065 40.850 ;
        RECT 21.855 40.680 22.025 40.850 ;
        RECT 22.815 40.680 22.985 40.850 ;
        RECT 23.775 40.680 23.945 40.850 ;
        RECT 24.735 40.680 24.905 40.850 ;
        RECT 19.935 37.085 20.105 37.255 ;
        RECT 19.935 36.725 20.105 36.895 ;
        RECT 19.935 36.365 20.105 36.535 ;
        RECT 20.895 37.085 21.065 37.255 ;
        RECT 20.895 36.725 21.065 36.895 ;
        RECT 20.895 36.365 21.065 36.535 ;
        RECT 21.855 37.085 22.025 37.255 ;
        RECT 21.855 36.725 22.025 36.895 ;
        RECT 21.855 36.365 22.025 36.535 ;
        RECT 22.815 37.085 22.985 37.255 ;
        RECT 22.815 36.725 22.985 36.895 ;
        RECT 22.815 36.365 22.985 36.535 ;
        RECT 23.775 37.085 23.945 37.255 ;
        RECT 23.775 36.725 23.945 36.895 ;
        RECT 23.775 36.365 23.945 36.535 ;
        RECT 24.735 37.085 24.905 37.255 ;
        RECT 24.735 36.725 24.905 36.895 ;
        RECT 24.735 36.365 24.905 36.535 ;
        RECT 19.935 34.245 20.105 34.415 ;
        RECT 20.895 34.245 21.065 34.415 ;
        RECT 21.855 34.245 22.025 34.415 ;
        RECT 22.815 34.245 22.985 34.415 ;
        RECT 23.775 34.245 23.945 34.415 ;
        RECT 24.735 34.245 24.905 34.415 ;
        RECT 19.935 30.650 20.105 30.820 ;
        RECT 19.935 30.290 20.105 30.460 ;
        RECT 19.935 29.930 20.105 30.100 ;
        RECT 20.895 30.650 21.065 30.820 ;
        RECT 20.895 30.290 21.065 30.460 ;
        RECT 20.895 29.930 21.065 30.100 ;
        RECT 21.855 30.650 22.025 30.820 ;
        RECT 21.855 30.290 22.025 30.460 ;
        RECT 21.855 29.930 22.025 30.100 ;
        RECT 22.815 30.650 22.985 30.820 ;
        RECT 22.815 30.290 22.985 30.460 ;
        RECT 22.815 29.930 22.985 30.100 ;
        RECT 23.775 30.650 23.945 30.820 ;
        RECT 23.775 30.290 23.945 30.460 ;
        RECT 23.775 29.930 23.945 30.100 ;
        RECT 24.735 30.650 24.905 30.820 ;
        RECT 24.735 30.290 24.905 30.460 ;
        RECT 24.735 29.930 24.905 30.100 ;
        RECT 19.935 27.810 20.105 27.980 ;
        RECT 20.895 27.810 21.065 27.980 ;
        RECT 21.855 27.810 22.025 27.980 ;
        RECT 22.815 27.810 22.985 27.980 ;
        RECT 23.775 27.810 23.945 27.980 ;
        RECT 24.735 27.810 24.905 27.980 ;
        RECT 19.935 24.215 20.105 24.385 ;
        RECT 19.935 23.855 20.105 24.025 ;
        RECT 19.935 23.495 20.105 23.665 ;
        RECT 20.895 24.215 21.065 24.385 ;
        RECT 20.895 23.855 21.065 24.025 ;
        RECT 20.895 23.495 21.065 23.665 ;
        RECT 21.855 24.215 22.025 24.385 ;
        RECT 21.855 23.855 22.025 24.025 ;
        RECT 21.855 23.495 22.025 23.665 ;
        RECT 22.815 24.215 22.985 24.385 ;
        RECT 22.815 23.855 22.985 24.025 ;
        RECT 22.815 23.495 22.985 23.665 ;
        RECT 23.775 24.215 23.945 24.385 ;
        RECT 23.775 23.855 23.945 24.025 ;
        RECT 23.775 23.495 23.945 23.665 ;
        RECT 24.735 24.215 24.905 24.385 ;
        RECT 24.735 23.855 24.905 24.025 ;
        RECT 24.735 23.495 24.905 23.665 ;
        RECT 19.935 21.375 20.105 21.545 ;
        RECT 20.895 21.375 21.065 21.545 ;
        RECT 21.855 21.375 22.025 21.545 ;
        RECT 22.815 21.375 22.985 21.545 ;
        RECT 23.775 21.375 23.945 21.545 ;
        RECT 24.735 21.375 24.905 21.545 ;
        RECT 19.935 17.780 20.105 17.950 ;
        RECT 19.935 17.420 20.105 17.590 ;
        RECT 19.935 17.060 20.105 17.230 ;
        RECT 20.895 17.780 21.065 17.950 ;
        RECT 20.895 17.420 21.065 17.590 ;
        RECT 20.895 17.060 21.065 17.230 ;
        RECT 21.855 17.780 22.025 17.950 ;
        RECT 21.855 17.420 22.025 17.590 ;
        RECT 21.855 17.060 22.025 17.230 ;
        RECT 22.815 17.780 22.985 17.950 ;
        RECT 22.815 17.420 22.985 17.590 ;
        RECT 22.815 17.060 22.985 17.230 ;
        RECT 23.775 17.780 23.945 17.950 ;
        RECT 23.775 17.420 23.945 17.590 ;
        RECT 23.775 17.060 23.945 17.230 ;
        RECT 24.735 17.780 24.905 17.950 ;
        RECT 24.735 17.420 24.905 17.590 ;
        RECT 24.735 17.060 24.905 17.230 ;
        RECT 19.935 14.940 20.105 15.110 ;
        RECT 20.895 14.940 21.065 15.110 ;
        RECT 21.855 14.940 22.025 15.110 ;
        RECT 22.815 14.940 22.985 15.110 ;
        RECT 23.775 14.940 23.945 15.110 ;
        RECT 24.735 14.940 24.905 15.110 ;
        RECT 19.935 11.345 20.105 11.515 ;
        RECT 19.935 10.985 20.105 11.155 ;
        RECT 19.935 10.625 20.105 10.795 ;
        RECT 20.895 11.345 21.065 11.515 ;
        RECT 20.895 10.985 21.065 11.155 ;
        RECT 20.895 10.625 21.065 10.795 ;
        RECT 21.855 11.345 22.025 11.515 ;
        RECT 21.855 10.985 22.025 11.155 ;
        RECT 21.855 10.625 22.025 10.795 ;
        RECT 22.815 11.345 22.985 11.515 ;
        RECT 22.815 10.985 22.985 11.155 ;
        RECT 22.815 10.625 22.985 10.795 ;
        RECT 23.775 11.345 23.945 11.515 ;
        RECT 23.775 10.985 23.945 11.155 ;
        RECT 23.775 10.625 23.945 10.795 ;
        RECT 24.735 11.345 24.905 11.515 ;
        RECT 24.735 10.985 24.905 11.155 ;
        RECT 24.735 10.625 24.905 10.795 ;
        RECT 19.935 8.505 20.105 8.675 ;
        RECT 20.895 8.505 21.065 8.675 ;
        RECT 21.855 8.505 22.025 8.675 ;
        RECT 22.815 8.505 22.985 8.675 ;
        RECT 23.775 8.505 23.945 8.675 ;
        RECT 24.735 8.505 24.905 8.675 ;
        RECT 19.935 4.910 20.105 5.080 ;
        RECT 19.935 4.550 20.105 4.720 ;
        RECT 19.935 4.190 20.105 4.360 ;
        RECT 20.895 4.910 21.065 5.080 ;
        RECT 20.895 4.550 21.065 4.720 ;
        RECT 20.895 4.190 21.065 4.360 ;
        RECT 21.855 4.910 22.025 5.080 ;
        RECT 21.855 4.550 22.025 4.720 ;
        RECT 21.855 4.190 22.025 4.360 ;
        RECT 22.815 4.910 22.985 5.080 ;
        RECT 22.815 4.550 22.985 4.720 ;
        RECT 22.815 4.190 22.985 4.360 ;
        RECT 23.775 4.910 23.945 5.080 ;
        RECT 23.775 4.550 23.945 4.720 ;
        RECT 23.775 4.190 23.945 4.360 ;
        RECT 24.735 4.910 24.905 5.080 ;
        RECT 24.735 4.550 24.905 4.720 ;
        RECT 24.735 4.190 24.905 4.360 ;
        RECT 19.935 2.070 20.105 2.240 ;
        RECT 20.895 2.070 21.065 2.240 ;
        RECT 21.855 2.070 22.025 2.240 ;
        RECT 22.815 2.070 22.985 2.240 ;
        RECT 23.775 2.070 23.945 2.240 ;
        RECT 24.735 2.070 24.905 2.240 ;
      LAYER met1 ;
        RECT 19.905 203.440 20.135 204.800 ;
        RECT 20.865 203.440 21.095 204.800 ;
        RECT 21.825 203.440 22.055 204.800 ;
        RECT 22.785 203.440 23.015 204.800 ;
        RECT 23.745 203.440 23.975 204.800 ;
        RECT 24.705 203.440 24.935 204.800 ;
        RECT 19.935 202.735 20.105 203.440 ;
        RECT 20.895 202.735 21.065 203.440 ;
        RECT 21.855 202.735 22.025 203.440 ;
        RECT 22.815 202.735 22.985 203.440 ;
        RECT 23.775 202.735 23.945 203.440 ;
        RECT 24.735 202.735 24.905 203.440 ;
        RECT 25.885 202.835 28.715 203.005 ;
        RECT 25.885 202.735 26.055 202.835 ;
        RECT 19.935 202.565 26.055 202.735 ;
        RECT 19.935 201.900 20.105 202.565 ;
        RECT 20.895 201.900 21.065 202.565 ;
        RECT 21.855 201.900 22.025 202.565 ;
        RECT 22.815 201.900 22.985 202.565 ;
        RECT 23.775 201.900 23.945 202.565 ;
        RECT 24.735 201.900 24.905 202.565 ;
        RECT 19.905 201.380 20.135 201.900 ;
        RECT 20.865 201.380 21.095 201.900 ;
        RECT 21.825 201.380 22.055 201.900 ;
        RECT 22.785 201.380 23.015 201.900 ;
        RECT 23.745 201.380 23.975 201.900 ;
        RECT 24.705 201.380 24.935 201.900 ;
        RECT 19.905 197.005 20.135 198.365 ;
        RECT 20.865 197.005 21.095 198.365 ;
        RECT 21.825 197.005 22.055 198.365 ;
        RECT 22.785 197.005 23.015 198.365 ;
        RECT 23.745 197.005 23.975 198.365 ;
        RECT 24.705 197.005 24.935 198.365 ;
        RECT 19.935 196.300 20.105 197.005 ;
        RECT 20.895 196.300 21.065 197.005 ;
        RECT 21.855 196.300 22.025 197.005 ;
        RECT 22.815 196.300 22.985 197.005 ;
        RECT 23.775 196.300 23.945 197.005 ;
        RECT 24.735 196.300 24.905 197.005 ;
        RECT 28.415 196.570 28.715 202.835 ;
        RECT 25.885 196.400 28.715 196.570 ;
        RECT 25.885 196.300 26.055 196.400 ;
        RECT 19.935 196.130 26.055 196.300 ;
        RECT 19.935 195.465 20.105 196.130 ;
        RECT 20.895 195.465 21.065 196.130 ;
        RECT 21.855 195.465 22.025 196.130 ;
        RECT 22.815 195.465 22.985 196.130 ;
        RECT 23.775 195.465 23.945 196.130 ;
        RECT 24.735 195.465 24.905 196.130 ;
        RECT 19.905 194.945 20.135 195.465 ;
        RECT 20.865 194.945 21.095 195.465 ;
        RECT 21.825 194.945 22.055 195.465 ;
        RECT 22.785 194.945 23.015 195.465 ;
        RECT 23.745 194.945 23.975 195.465 ;
        RECT 24.705 194.945 24.935 195.465 ;
        RECT 19.905 190.570 20.135 191.930 ;
        RECT 20.865 190.570 21.095 191.930 ;
        RECT 21.825 190.570 22.055 191.930 ;
        RECT 22.785 190.570 23.015 191.930 ;
        RECT 23.745 190.570 23.975 191.930 ;
        RECT 24.705 190.570 24.935 191.930 ;
        RECT 19.935 189.865 20.105 190.570 ;
        RECT 20.895 189.865 21.065 190.570 ;
        RECT 21.855 189.865 22.025 190.570 ;
        RECT 22.815 189.865 22.985 190.570 ;
        RECT 23.775 189.865 23.945 190.570 ;
        RECT 24.735 189.865 24.905 190.570 ;
        RECT 28.415 190.135 28.715 196.400 ;
        RECT 25.885 189.965 28.715 190.135 ;
        RECT 25.885 189.865 26.055 189.965 ;
        RECT 19.935 189.695 26.055 189.865 ;
        RECT 19.935 189.030 20.105 189.695 ;
        RECT 20.895 189.030 21.065 189.695 ;
        RECT 21.855 189.030 22.025 189.695 ;
        RECT 22.815 189.030 22.985 189.695 ;
        RECT 23.775 189.030 23.945 189.695 ;
        RECT 24.735 189.030 24.905 189.695 ;
        RECT 19.905 188.510 20.135 189.030 ;
        RECT 20.865 188.510 21.095 189.030 ;
        RECT 21.825 188.510 22.055 189.030 ;
        RECT 22.785 188.510 23.015 189.030 ;
        RECT 23.745 188.510 23.975 189.030 ;
        RECT 24.705 188.510 24.935 189.030 ;
        RECT 19.905 184.135 20.135 185.495 ;
        RECT 20.865 184.135 21.095 185.495 ;
        RECT 21.825 184.135 22.055 185.495 ;
        RECT 22.785 184.135 23.015 185.495 ;
        RECT 23.745 184.135 23.975 185.495 ;
        RECT 24.705 184.135 24.935 185.495 ;
        RECT 19.935 183.430 20.105 184.135 ;
        RECT 20.895 183.430 21.065 184.135 ;
        RECT 21.855 183.430 22.025 184.135 ;
        RECT 22.815 183.430 22.985 184.135 ;
        RECT 23.775 183.430 23.945 184.135 ;
        RECT 24.735 183.430 24.905 184.135 ;
        RECT 28.415 183.700 28.715 189.965 ;
        RECT 25.885 183.530 28.715 183.700 ;
        RECT 25.885 183.430 26.055 183.530 ;
        RECT 19.935 183.260 26.055 183.430 ;
        RECT 19.935 182.595 20.105 183.260 ;
        RECT 20.895 182.595 21.065 183.260 ;
        RECT 21.855 182.595 22.025 183.260 ;
        RECT 22.815 182.595 22.985 183.260 ;
        RECT 23.775 182.595 23.945 183.260 ;
        RECT 24.735 182.595 24.905 183.260 ;
        RECT 19.905 182.075 20.135 182.595 ;
        RECT 20.865 182.075 21.095 182.595 ;
        RECT 21.825 182.075 22.055 182.595 ;
        RECT 22.785 182.075 23.015 182.595 ;
        RECT 23.745 182.075 23.975 182.595 ;
        RECT 24.705 182.075 24.935 182.595 ;
        RECT 19.905 177.700 20.135 179.060 ;
        RECT 20.865 177.700 21.095 179.060 ;
        RECT 21.825 177.700 22.055 179.060 ;
        RECT 22.785 177.700 23.015 179.060 ;
        RECT 23.745 177.700 23.975 179.060 ;
        RECT 24.705 177.700 24.935 179.060 ;
        RECT 19.935 176.995 20.105 177.700 ;
        RECT 20.895 176.995 21.065 177.700 ;
        RECT 21.855 176.995 22.025 177.700 ;
        RECT 22.815 176.995 22.985 177.700 ;
        RECT 23.775 176.995 23.945 177.700 ;
        RECT 24.735 176.995 24.905 177.700 ;
        RECT 28.415 177.265 28.715 183.530 ;
        RECT 25.885 177.095 28.715 177.265 ;
        RECT 25.885 176.995 26.055 177.095 ;
        RECT 19.935 176.825 26.055 176.995 ;
        RECT 19.935 176.160 20.105 176.825 ;
        RECT 20.895 176.160 21.065 176.825 ;
        RECT 21.855 176.160 22.025 176.825 ;
        RECT 22.815 176.160 22.985 176.825 ;
        RECT 23.775 176.160 23.945 176.825 ;
        RECT 24.735 176.160 24.905 176.825 ;
        RECT 19.905 175.640 20.135 176.160 ;
        RECT 20.865 175.640 21.095 176.160 ;
        RECT 21.825 175.640 22.055 176.160 ;
        RECT 22.785 175.640 23.015 176.160 ;
        RECT 23.745 175.640 23.975 176.160 ;
        RECT 24.705 175.640 24.935 176.160 ;
        RECT 19.905 171.265 20.135 172.625 ;
        RECT 20.865 171.265 21.095 172.625 ;
        RECT 21.825 171.265 22.055 172.625 ;
        RECT 22.785 171.265 23.015 172.625 ;
        RECT 23.745 171.265 23.975 172.625 ;
        RECT 24.705 171.265 24.935 172.625 ;
        RECT 19.935 170.560 20.105 171.265 ;
        RECT 20.895 170.560 21.065 171.265 ;
        RECT 21.855 170.560 22.025 171.265 ;
        RECT 22.815 170.560 22.985 171.265 ;
        RECT 23.775 170.560 23.945 171.265 ;
        RECT 24.735 170.560 24.905 171.265 ;
        RECT 28.415 170.830 28.715 177.095 ;
        RECT 25.885 170.660 28.715 170.830 ;
        RECT 25.885 170.560 26.055 170.660 ;
        RECT 19.935 170.390 26.055 170.560 ;
        RECT 19.935 169.725 20.105 170.390 ;
        RECT 20.895 169.725 21.065 170.390 ;
        RECT 21.855 169.725 22.025 170.390 ;
        RECT 22.815 169.725 22.985 170.390 ;
        RECT 23.775 169.725 23.945 170.390 ;
        RECT 24.735 169.725 24.905 170.390 ;
        RECT 19.905 169.205 20.135 169.725 ;
        RECT 20.865 169.205 21.095 169.725 ;
        RECT 21.825 169.205 22.055 169.725 ;
        RECT 22.785 169.205 23.015 169.725 ;
        RECT 23.745 169.205 23.975 169.725 ;
        RECT 24.705 169.205 24.935 169.725 ;
        RECT 19.905 164.830 20.135 166.190 ;
        RECT 20.865 164.830 21.095 166.190 ;
        RECT 21.825 164.830 22.055 166.190 ;
        RECT 22.785 164.830 23.015 166.190 ;
        RECT 23.745 164.830 23.975 166.190 ;
        RECT 24.705 164.830 24.935 166.190 ;
        RECT 19.935 164.125 20.105 164.830 ;
        RECT 20.895 164.125 21.065 164.830 ;
        RECT 21.855 164.125 22.025 164.830 ;
        RECT 22.815 164.125 22.985 164.830 ;
        RECT 23.775 164.125 23.945 164.830 ;
        RECT 24.735 164.125 24.905 164.830 ;
        RECT 28.415 164.395 28.715 170.660 ;
        RECT 25.885 164.225 28.715 164.395 ;
        RECT 25.885 164.125 26.055 164.225 ;
        RECT 19.935 163.955 26.055 164.125 ;
        RECT 19.935 163.290 20.105 163.955 ;
        RECT 20.895 163.290 21.065 163.955 ;
        RECT 21.855 163.290 22.025 163.955 ;
        RECT 22.815 163.290 22.985 163.955 ;
        RECT 23.775 163.290 23.945 163.955 ;
        RECT 24.735 163.290 24.905 163.955 ;
        RECT 19.905 162.770 20.135 163.290 ;
        RECT 20.865 162.770 21.095 163.290 ;
        RECT 21.825 162.770 22.055 163.290 ;
        RECT 22.785 162.770 23.015 163.290 ;
        RECT 23.745 162.770 23.975 163.290 ;
        RECT 24.705 162.770 24.935 163.290 ;
        RECT 19.905 158.395 20.135 159.755 ;
        RECT 20.865 158.395 21.095 159.755 ;
        RECT 21.825 158.395 22.055 159.755 ;
        RECT 22.785 158.395 23.015 159.755 ;
        RECT 23.745 158.395 23.975 159.755 ;
        RECT 24.705 158.395 24.935 159.755 ;
        RECT 19.935 157.690 20.105 158.395 ;
        RECT 20.895 157.690 21.065 158.395 ;
        RECT 21.855 157.690 22.025 158.395 ;
        RECT 22.815 157.690 22.985 158.395 ;
        RECT 23.775 157.690 23.945 158.395 ;
        RECT 24.735 157.690 24.905 158.395 ;
        RECT 28.415 157.960 28.715 164.225 ;
        RECT 25.885 157.790 28.715 157.960 ;
        RECT 25.885 157.690 26.055 157.790 ;
        RECT 19.935 157.520 26.055 157.690 ;
        RECT 19.935 156.855 20.105 157.520 ;
        RECT 20.895 156.855 21.065 157.520 ;
        RECT 21.855 156.855 22.025 157.520 ;
        RECT 22.815 156.855 22.985 157.520 ;
        RECT 23.775 156.855 23.945 157.520 ;
        RECT 24.735 156.855 24.905 157.520 ;
        RECT 19.905 156.335 20.135 156.855 ;
        RECT 20.865 156.335 21.095 156.855 ;
        RECT 21.825 156.335 22.055 156.855 ;
        RECT 22.785 156.335 23.015 156.855 ;
        RECT 23.745 156.335 23.975 156.855 ;
        RECT 24.705 156.335 24.935 156.855 ;
        RECT 19.905 151.960 20.135 153.320 ;
        RECT 20.865 151.960 21.095 153.320 ;
        RECT 21.825 151.960 22.055 153.320 ;
        RECT 22.785 151.960 23.015 153.320 ;
        RECT 23.745 151.960 23.975 153.320 ;
        RECT 24.705 151.960 24.935 153.320 ;
        RECT 19.935 151.255 20.105 151.960 ;
        RECT 20.895 151.255 21.065 151.960 ;
        RECT 21.855 151.255 22.025 151.960 ;
        RECT 22.815 151.255 22.985 151.960 ;
        RECT 23.775 151.255 23.945 151.960 ;
        RECT 24.735 151.255 24.905 151.960 ;
        RECT 28.415 151.525 28.715 157.790 ;
        RECT 25.885 151.355 28.715 151.525 ;
        RECT 25.885 151.255 26.055 151.355 ;
        RECT 19.935 151.085 26.055 151.255 ;
        RECT 19.935 150.420 20.105 151.085 ;
        RECT 20.895 150.420 21.065 151.085 ;
        RECT 21.855 150.420 22.025 151.085 ;
        RECT 22.815 150.420 22.985 151.085 ;
        RECT 23.775 150.420 23.945 151.085 ;
        RECT 24.735 150.420 24.905 151.085 ;
        RECT 19.905 149.900 20.135 150.420 ;
        RECT 20.865 149.900 21.095 150.420 ;
        RECT 21.825 149.900 22.055 150.420 ;
        RECT 22.785 149.900 23.015 150.420 ;
        RECT 23.745 149.900 23.975 150.420 ;
        RECT 24.705 149.900 24.935 150.420 ;
        RECT 19.905 145.525 20.135 146.885 ;
        RECT 20.865 145.525 21.095 146.885 ;
        RECT 21.825 145.525 22.055 146.885 ;
        RECT 22.785 145.525 23.015 146.885 ;
        RECT 23.745 145.525 23.975 146.885 ;
        RECT 24.705 145.525 24.935 146.885 ;
        RECT 19.935 144.820 20.105 145.525 ;
        RECT 20.895 144.820 21.065 145.525 ;
        RECT 21.855 144.820 22.025 145.525 ;
        RECT 22.815 144.820 22.985 145.525 ;
        RECT 23.775 144.820 23.945 145.525 ;
        RECT 24.735 144.820 24.905 145.525 ;
        RECT 28.415 145.090 28.715 151.355 ;
        RECT 25.885 144.920 28.715 145.090 ;
        RECT 25.885 144.820 26.055 144.920 ;
        RECT 19.935 144.650 26.055 144.820 ;
        RECT 19.935 143.985 20.105 144.650 ;
        RECT 20.895 143.985 21.065 144.650 ;
        RECT 21.855 143.985 22.025 144.650 ;
        RECT 22.815 143.985 22.985 144.650 ;
        RECT 23.775 143.985 23.945 144.650 ;
        RECT 24.735 143.985 24.905 144.650 ;
        RECT 19.905 143.465 20.135 143.985 ;
        RECT 20.865 143.465 21.095 143.985 ;
        RECT 21.825 143.465 22.055 143.985 ;
        RECT 22.785 143.465 23.015 143.985 ;
        RECT 23.745 143.465 23.975 143.985 ;
        RECT 24.705 143.465 24.935 143.985 ;
        RECT 19.905 139.090 20.135 140.450 ;
        RECT 20.865 139.090 21.095 140.450 ;
        RECT 21.825 139.090 22.055 140.450 ;
        RECT 22.785 139.090 23.015 140.450 ;
        RECT 23.745 139.090 23.975 140.450 ;
        RECT 24.705 139.090 24.935 140.450 ;
        RECT 19.935 138.385 20.105 139.090 ;
        RECT 20.895 138.385 21.065 139.090 ;
        RECT 21.855 138.385 22.025 139.090 ;
        RECT 22.815 138.385 22.985 139.090 ;
        RECT 23.775 138.385 23.945 139.090 ;
        RECT 24.735 138.385 24.905 139.090 ;
        RECT 28.415 138.655 28.715 144.920 ;
        RECT 25.885 138.485 28.715 138.655 ;
        RECT 25.885 138.385 26.055 138.485 ;
        RECT 19.935 138.215 26.055 138.385 ;
        RECT 19.935 137.550 20.105 138.215 ;
        RECT 20.895 137.550 21.065 138.215 ;
        RECT 21.855 137.550 22.025 138.215 ;
        RECT 22.815 137.550 22.985 138.215 ;
        RECT 23.775 137.550 23.945 138.215 ;
        RECT 24.735 137.550 24.905 138.215 ;
        RECT 19.905 137.030 20.135 137.550 ;
        RECT 20.865 137.030 21.095 137.550 ;
        RECT 21.825 137.030 22.055 137.550 ;
        RECT 22.785 137.030 23.015 137.550 ;
        RECT 23.745 137.030 23.975 137.550 ;
        RECT 24.705 137.030 24.935 137.550 ;
        RECT 19.905 132.655 20.135 134.015 ;
        RECT 20.865 132.655 21.095 134.015 ;
        RECT 21.825 132.655 22.055 134.015 ;
        RECT 22.785 132.655 23.015 134.015 ;
        RECT 23.745 132.655 23.975 134.015 ;
        RECT 24.705 132.655 24.935 134.015 ;
        RECT 19.935 131.950 20.105 132.655 ;
        RECT 20.895 131.950 21.065 132.655 ;
        RECT 21.855 131.950 22.025 132.655 ;
        RECT 22.815 131.950 22.985 132.655 ;
        RECT 23.775 131.950 23.945 132.655 ;
        RECT 24.735 131.950 24.905 132.655 ;
        RECT 28.415 132.220 28.715 138.485 ;
        RECT 25.885 132.050 28.715 132.220 ;
        RECT 25.885 131.950 26.055 132.050 ;
        RECT 19.935 131.780 26.055 131.950 ;
        RECT 19.935 131.115 20.105 131.780 ;
        RECT 20.895 131.115 21.065 131.780 ;
        RECT 21.855 131.115 22.025 131.780 ;
        RECT 22.815 131.115 22.985 131.780 ;
        RECT 23.775 131.115 23.945 131.780 ;
        RECT 24.735 131.115 24.905 131.780 ;
        RECT 19.905 130.595 20.135 131.115 ;
        RECT 20.865 130.595 21.095 131.115 ;
        RECT 21.825 130.595 22.055 131.115 ;
        RECT 22.785 130.595 23.015 131.115 ;
        RECT 23.745 130.595 23.975 131.115 ;
        RECT 24.705 130.595 24.935 131.115 ;
        RECT 19.905 126.220 20.135 127.580 ;
        RECT 20.865 126.220 21.095 127.580 ;
        RECT 21.825 126.220 22.055 127.580 ;
        RECT 22.785 126.220 23.015 127.580 ;
        RECT 23.745 126.220 23.975 127.580 ;
        RECT 24.705 126.220 24.935 127.580 ;
        RECT 19.935 125.515 20.105 126.220 ;
        RECT 20.895 125.515 21.065 126.220 ;
        RECT 21.855 125.515 22.025 126.220 ;
        RECT 22.815 125.515 22.985 126.220 ;
        RECT 23.775 125.515 23.945 126.220 ;
        RECT 24.735 125.515 24.905 126.220 ;
        RECT 28.415 125.785 28.715 132.050 ;
        RECT 25.885 125.615 28.715 125.785 ;
        RECT 25.885 125.515 26.055 125.615 ;
        RECT 19.935 125.345 26.055 125.515 ;
        RECT 19.935 124.680 20.105 125.345 ;
        RECT 20.895 124.680 21.065 125.345 ;
        RECT 21.855 124.680 22.025 125.345 ;
        RECT 22.815 124.680 22.985 125.345 ;
        RECT 23.775 124.680 23.945 125.345 ;
        RECT 24.735 124.680 24.905 125.345 ;
        RECT 19.905 124.160 20.135 124.680 ;
        RECT 20.865 124.160 21.095 124.680 ;
        RECT 21.825 124.160 22.055 124.680 ;
        RECT 22.785 124.160 23.015 124.680 ;
        RECT 23.745 124.160 23.975 124.680 ;
        RECT 24.705 124.160 24.935 124.680 ;
        RECT 19.905 119.785 20.135 121.145 ;
        RECT 20.865 119.785 21.095 121.145 ;
        RECT 21.825 119.785 22.055 121.145 ;
        RECT 22.785 119.785 23.015 121.145 ;
        RECT 23.745 119.785 23.975 121.145 ;
        RECT 24.705 119.785 24.935 121.145 ;
        RECT 19.935 119.080 20.105 119.785 ;
        RECT 20.895 119.080 21.065 119.785 ;
        RECT 21.855 119.080 22.025 119.785 ;
        RECT 22.815 119.080 22.985 119.785 ;
        RECT 23.775 119.080 23.945 119.785 ;
        RECT 24.735 119.080 24.905 119.785 ;
        RECT 28.415 119.350 28.715 125.615 ;
        RECT 25.885 119.180 28.715 119.350 ;
        RECT 25.885 119.080 26.055 119.180 ;
        RECT 19.935 118.910 26.055 119.080 ;
        RECT 19.935 118.245 20.105 118.910 ;
        RECT 20.895 118.245 21.065 118.910 ;
        RECT 21.855 118.245 22.025 118.910 ;
        RECT 22.815 118.245 22.985 118.910 ;
        RECT 23.775 118.245 23.945 118.910 ;
        RECT 24.735 118.245 24.905 118.910 ;
        RECT 19.905 117.725 20.135 118.245 ;
        RECT 20.865 117.725 21.095 118.245 ;
        RECT 21.825 117.725 22.055 118.245 ;
        RECT 22.785 117.725 23.015 118.245 ;
        RECT 23.745 117.725 23.975 118.245 ;
        RECT 24.705 117.725 24.935 118.245 ;
        RECT 19.905 113.350 20.135 114.710 ;
        RECT 20.865 113.350 21.095 114.710 ;
        RECT 21.825 113.350 22.055 114.710 ;
        RECT 22.785 113.350 23.015 114.710 ;
        RECT 23.745 113.350 23.975 114.710 ;
        RECT 24.705 113.350 24.935 114.710 ;
        RECT 19.935 112.645 20.105 113.350 ;
        RECT 20.895 112.645 21.065 113.350 ;
        RECT 21.855 112.645 22.025 113.350 ;
        RECT 22.815 112.645 22.985 113.350 ;
        RECT 23.775 112.645 23.945 113.350 ;
        RECT 24.735 112.645 24.905 113.350 ;
        RECT 28.415 112.915 28.715 119.180 ;
        RECT 25.885 112.745 28.715 112.915 ;
        RECT 25.885 112.645 26.055 112.745 ;
        RECT 19.935 112.475 26.055 112.645 ;
        RECT 19.935 111.810 20.105 112.475 ;
        RECT 20.895 111.810 21.065 112.475 ;
        RECT 21.855 111.810 22.025 112.475 ;
        RECT 22.815 111.810 22.985 112.475 ;
        RECT 23.775 111.810 23.945 112.475 ;
        RECT 24.735 111.810 24.905 112.475 ;
        RECT 19.905 111.290 20.135 111.810 ;
        RECT 20.865 111.290 21.095 111.810 ;
        RECT 21.825 111.290 22.055 111.810 ;
        RECT 22.785 111.290 23.015 111.810 ;
        RECT 23.745 111.290 23.975 111.810 ;
        RECT 24.705 111.290 24.935 111.810 ;
        RECT 19.905 106.915 20.135 108.275 ;
        RECT 20.865 106.915 21.095 108.275 ;
        RECT 21.825 106.915 22.055 108.275 ;
        RECT 22.785 106.915 23.015 108.275 ;
        RECT 23.745 106.915 23.975 108.275 ;
        RECT 24.705 106.915 24.935 108.275 ;
        RECT 19.935 106.210 20.105 106.915 ;
        RECT 20.895 106.210 21.065 106.915 ;
        RECT 21.855 106.210 22.025 106.915 ;
        RECT 22.815 106.210 22.985 106.915 ;
        RECT 23.775 106.210 23.945 106.915 ;
        RECT 24.735 106.210 24.905 106.915 ;
        RECT 28.415 106.480 28.715 112.745 ;
        RECT 25.885 106.310 28.715 106.480 ;
        RECT 25.885 106.210 26.055 106.310 ;
        RECT 19.935 106.040 26.055 106.210 ;
        RECT 19.935 105.375 20.105 106.040 ;
        RECT 20.895 105.375 21.065 106.040 ;
        RECT 21.855 105.375 22.025 106.040 ;
        RECT 22.815 105.375 22.985 106.040 ;
        RECT 23.775 105.375 23.945 106.040 ;
        RECT 24.735 105.375 24.905 106.040 ;
        RECT 19.905 104.855 20.135 105.375 ;
        RECT 20.865 104.855 21.095 105.375 ;
        RECT 21.825 104.855 22.055 105.375 ;
        RECT 22.785 104.855 23.015 105.375 ;
        RECT 23.745 104.855 23.975 105.375 ;
        RECT 24.705 104.855 24.935 105.375 ;
        RECT 19.905 100.480 20.135 101.840 ;
        RECT 20.865 100.480 21.095 101.840 ;
        RECT 21.825 100.480 22.055 101.840 ;
        RECT 22.785 100.480 23.015 101.840 ;
        RECT 23.745 100.480 23.975 101.840 ;
        RECT 24.705 100.480 24.935 101.840 ;
        RECT 19.935 99.775 20.105 100.480 ;
        RECT 20.895 99.775 21.065 100.480 ;
        RECT 21.855 99.775 22.025 100.480 ;
        RECT 22.815 99.775 22.985 100.480 ;
        RECT 23.775 99.775 23.945 100.480 ;
        RECT 24.735 99.775 24.905 100.480 ;
        RECT 28.415 100.045 28.715 106.310 ;
        RECT 25.885 99.875 28.715 100.045 ;
        RECT 25.885 99.775 26.055 99.875 ;
        RECT 19.935 99.605 26.055 99.775 ;
        RECT 19.935 98.940 20.105 99.605 ;
        RECT 20.895 98.940 21.065 99.605 ;
        RECT 21.855 98.940 22.025 99.605 ;
        RECT 22.815 98.940 22.985 99.605 ;
        RECT 23.775 98.940 23.945 99.605 ;
        RECT 24.735 98.940 24.905 99.605 ;
        RECT 19.905 98.420 20.135 98.940 ;
        RECT 20.865 98.420 21.095 98.940 ;
        RECT 21.825 98.420 22.055 98.940 ;
        RECT 22.785 98.420 23.015 98.940 ;
        RECT 23.745 98.420 23.975 98.940 ;
        RECT 24.705 98.420 24.935 98.940 ;
        RECT 19.905 94.045 20.135 95.405 ;
        RECT 20.865 94.045 21.095 95.405 ;
        RECT 21.825 94.045 22.055 95.405 ;
        RECT 22.785 94.045 23.015 95.405 ;
        RECT 23.745 94.045 23.975 95.405 ;
        RECT 24.705 94.045 24.935 95.405 ;
        RECT 19.935 93.340 20.105 94.045 ;
        RECT 20.895 93.340 21.065 94.045 ;
        RECT 21.855 93.340 22.025 94.045 ;
        RECT 22.815 93.340 22.985 94.045 ;
        RECT 23.775 93.340 23.945 94.045 ;
        RECT 24.735 93.340 24.905 94.045 ;
        RECT 28.415 93.610 28.715 99.875 ;
        RECT 25.885 93.440 28.715 93.610 ;
        RECT 25.885 93.340 26.055 93.440 ;
        RECT 19.935 93.170 26.055 93.340 ;
        RECT 19.935 92.505 20.105 93.170 ;
        RECT 20.895 92.505 21.065 93.170 ;
        RECT 21.855 92.505 22.025 93.170 ;
        RECT 22.815 92.505 22.985 93.170 ;
        RECT 23.775 92.505 23.945 93.170 ;
        RECT 24.735 92.505 24.905 93.170 ;
        RECT 19.905 91.985 20.135 92.505 ;
        RECT 20.865 91.985 21.095 92.505 ;
        RECT 21.825 91.985 22.055 92.505 ;
        RECT 22.785 91.985 23.015 92.505 ;
        RECT 23.745 91.985 23.975 92.505 ;
        RECT 24.705 91.985 24.935 92.505 ;
        RECT 19.905 87.610 20.135 88.970 ;
        RECT 20.865 87.610 21.095 88.970 ;
        RECT 21.825 87.610 22.055 88.970 ;
        RECT 22.785 87.610 23.015 88.970 ;
        RECT 23.745 87.610 23.975 88.970 ;
        RECT 24.705 87.610 24.935 88.970 ;
        RECT 19.935 86.905 20.105 87.610 ;
        RECT 20.895 86.905 21.065 87.610 ;
        RECT 21.855 86.905 22.025 87.610 ;
        RECT 22.815 86.905 22.985 87.610 ;
        RECT 23.775 86.905 23.945 87.610 ;
        RECT 24.735 86.905 24.905 87.610 ;
        RECT 28.415 87.175 28.715 93.440 ;
        RECT 25.885 87.005 28.715 87.175 ;
        RECT 25.885 86.905 26.055 87.005 ;
        RECT 19.935 86.735 26.055 86.905 ;
        RECT 19.935 86.070 20.105 86.735 ;
        RECT 20.895 86.070 21.065 86.735 ;
        RECT 21.855 86.070 22.025 86.735 ;
        RECT 22.815 86.070 22.985 86.735 ;
        RECT 23.775 86.070 23.945 86.735 ;
        RECT 24.735 86.070 24.905 86.735 ;
        RECT 19.905 85.550 20.135 86.070 ;
        RECT 20.865 85.550 21.095 86.070 ;
        RECT 21.825 85.550 22.055 86.070 ;
        RECT 22.785 85.550 23.015 86.070 ;
        RECT 23.745 85.550 23.975 86.070 ;
        RECT 24.705 85.550 24.935 86.070 ;
        RECT 19.905 81.175 20.135 82.535 ;
        RECT 20.865 81.175 21.095 82.535 ;
        RECT 21.825 81.175 22.055 82.535 ;
        RECT 22.785 81.175 23.015 82.535 ;
        RECT 23.745 81.175 23.975 82.535 ;
        RECT 24.705 81.175 24.935 82.535 ;
        RECT 19.935 80.470 20.105 81.175 ;
        RECT 20.895 80.470 21.065 81.175 ;
        RECT 21.855 80.470 22.025 81.175 ;
        RECT 22.815 80.470 22.985 81.175 ;
        RECT 23.775 80.470 23.945 81.175 ;
        RECT 24.735 80.470 24.905 81.175 ;
        RECT 28.415 80.740 28.715 87.005 ;
        RECT 25.885 80.570 28.715 80.740 ;
        RECT 25.885 80.470 26.055 80.570 ;
        RECT 19.935 80.300 26.055 80.470 ;
        RECT 19.935 79.635 20.105 80.300 ;
        RECT 20.895 79.635 21.065 80.300 ;
        RECT 21.855 79.635 22.025 80.300 ;
        RECT 22.815 79.635 22.985 80.300 ;
        RECT 23.775 79.635 23.945 80.300 ;
        RECT 24.735 79.635 24.905 80.300 ;
        RECT 19.905 79.115 20.135 79.635 ;
        RECT 20.865 79.115 21.095 79.635 ;
        RECT 21.825 79.115 22.055 79.635 ;
        RECT 22.785 79.115 23.015 79.635 ;
        RECT 23.745 79.115 23.975 79.635 ;
        RECT 24.705 79.115 24.935 79.635 ;
        RECT 19.905 74.740 20.135 76.100 ;
        RECT 20.865 74.740 21.095 76.100 ;
        RECT 21.825 74.740 22.055 76.100 ;
        RECT 22.785 74.740 23.015 76.100 ;
        RECT 23.745 74.740 23.975 76.100 ;
        RECT 24.705 74.740 24.935 76.100 ;
        RECT 19.935 74.035 20.105 74.740 ;
        RECT 20.895 74.035 21.065 74.740 ;
        RECT 21.855 74.035 22.025 74.740 ;
        RECT 22.815 74.035 22.985 74.740 ;
        RECT 23.775 74.035 23.945 74.740 ;
        RECT 24.735 74.035 24.905 74.740 ;
        RECT 28.415 74.305 28.715 80.570 ;
        RECT 25.885 74.135 28.715 74.305 ;
        RECT 25.885 74.035 26.055 74.135 ;
        RECT 19.935 73.865 26.055 74.035 ;
        RECT 19.935 73.200 20.105 73.865 ;
        RECT 20.895 73.200 21.065 73.865 ;
        RECT 21.855 73.200 22.025 73.865 ;
        RECT 22.815 73.200 22.985 73.865 ;
        RECT 23.775 73.200 23.945 73.865 ;
        RECT 24.735 73.200 24.905 73.865 ;
        RECT 19.905 72.680 20.135 73.200 ;
        RECT 20.865 72.680 21.095 73.200 ;
        RECT 21.825 72.680 22.055 73.200 ;
        RECT 22.785 72.680 23.015 73.200 ;
        RECT 23.745 72.680 23.975 73.200 ;
        RECT 24.705 72.680 24.935 73.200 ;
        RECT 19.905 68.305 20.135 69.665 ;
        RECT 20.865 68.305 21.095 69.665 ;
        RECT 21.825 68.305 22.055 69.665 ;
        RECT 22.785 68.305 23.015 69.665 ;
        RECT 23.745 68.305 23.975 69.665 ;
        RECT 24.705 68.305 24.935 69.665 ;
        RECT 19.935 67.600 20.105 68.305 ;
        RECT 20.895 67.600 21.065 68.305 ;
        RECT 21.855 67.600 22.025 68.305 ;
        RECT 22.815 67.600 22.985 68.305 ;
        RECT 23.775 67.600 23.945 68.305 ;
        RECT 24.735 67.600 24.905 68.305 ;
        RECT 28.415 67.870 28.715 74.135 ;
        RECT 25.885 67.700 28.715 67.870 ;
        RECT 25.885 67.600 26.055 67.700 ;
        RECT 19.935 67.430 26.055 67.600 ;
        RECT 19.935 66.765 20.105 67.430 ;
        RECT 20.895 66.765 21.065 67.430 ;
        RECT 21.855 66.765 22.025 67.430 ;
        RECT 22.815 66.765 22.985 67.430 ;
        RECT 23.775 66.765 23.945 67.430 ;
        RECT 24.735 66.765 24.905 67.430 ;
        RECT 19.905 66.245 20.135 66.765 ;
        RECT 20.865 66.245 21.095 66.765 ;
        RECT 21.825 66.245 22.055 66.765 ;
        RECT 22.785 66.245 23.015 66.765 ;
        RECT 23.745 66.245 23.975 66.765 ;
        RECT 24.705 66.245 24.935 66.765 ;
        RECT 19.905 61.870 20.135 63.230 ;
        RECT 20.865 61.870 21.095 63.230 ;
        RECT 21.825 61.870 22.055 63.230 ;
        RECT 22.785 61.870 23.015 63.230 ;
        RECT 23.745 61.870 23.975 63.230 ;
        RECT 24.705 61.870 24.935 63.230 ;
        RECT 19.935 61.165 20.105 61.870 ;
        RECT 20.895 61.165 21.065 61.870 ;
        RECT 21.855 61.165 22.025 61.870 ;
        RECT 22.815 61.165 22.985 61.870 ;
        RECT 23.775 61.165 23.945 61.870 ;
        RECT 24.735 61.165 24.905 61.870 ;
        RECT 28.415 61.435 28.715 67.700 ;
        RECT 25.885 61.265 28.715 61.435 ;
        RECT 25.885 61.165 26.055 61.265 ;
        RECT 19.935 60.995 26.055 61.165 ;
        RECT 19.935 60.330 20.105 60.995 ;
        RECT 20.895 60.330 21.065 60.995 ;
        RECT 21.855 60.330 22.025 60.995 ;
        RECT 22.815 60.330 22.985 60.995 ;
        RECT 23.775 60.330 23.945 60.995 ;
        RECT 24.735 60.330 24.905 60.995 ;
        RECT 19.905 59.810 20.135 60.330 ;
        RECT 20.865 59.810 21.095 60.330 ;
        RECT 21.825 59.810 22.055 60.330 ;
        RECT 22.785 59.810 23.015 60.330 ;
        RECT 23.745 59.810 23.975 60.330 ;
        RECT 24.705 59.810 24.935 60.330 ;
        RECT 19.905 55.435 20.135 56.795 ;
        RECT 20.865 55.435 21.095 56.795 ;
        RECT 21.825 55.435 22.055 56.795 ;
        RECT 22.785 55.435 23.015 56.795 ;
        RECT 23.745 55.435 23.975 56.795 ;
        RECT 24.705 55.435 24.935 56.795 ;
        RECT 19.935 54.730 20.105 55.435 ;
        RECT 20.895 54.730 21.065 55.435 ;
        RECT 21.855 54.730 22.025 55.435 ;
        RECT 22.815 54.730 22.985 55.435 ;
        RECT 23.775 54.730 23.945 55.435 ;
        RECT 24.735 54.730 24.905 55.435 ;
        RECT 28.415 55.000 28.715 61.265 ;
        RECT 25.885 54.830 28.715 55.000 ;
        RECT 25.885 54.730 26.055 54.830 ;
        RECT 19.935 54.560 26.055 54.730 ;
        RECT 19.935 53.895 20.105 54.560 ;
        RECT 20.895 53.895 21.065 54.560 ;
        RECT 21.855 53.895 22.025 54.560 ;
        RECT 22.815 53.895 22.985 54.560 ;
        RECT 23.775 53.895 23.945 54.560 ;
        RECT 24.735 53.895 24.905 54.560 ;
        RECT 19.905 53.375 20.135 53.895 ;
        RECT 20.865 53.375 21.095 53.895 ;
        RECT 21.825 53.375 22.055 53.895 ;
        RECT 22.785 53.375 23.015 53.895 ;
        RECT 23.745 53.375 23.975 53.895 ;
        RECT 24.705 53.375 24.935 53.895 ;
        RECT 19.905 49.000 20.135 50.360 ;
        RECT 20.865 49.000 21.095 50.360 ;
        RECT 21.825 49.000 22.055 50.360 ;
        RECT 22.785 49.000 23.015 50.360 ;
        RECT 23.745 49.000 23.975 50.360 ;
        RECT 24.705 49.000 24.935 50.360 ;
        RECT 19.935 48.295 20.105 49.000 ;
        RECT 20.895 48.295 21.065 49.000 ;
        RECT 21.855 48.295 22.025 49.000 ;
        RECT 22.815 48.295 22.985 49.000 ;
        RECT 23.775 48.295 23.945 49.000 ;
        RECT 24.735 48.295 24.905 49.000 ;
        RECT 28.415 48.565 28.715 54.830 ;
        RECT 25.885 48.395 28.715 48.565 ;
        RECT 25.885 48.295 26.055 48.395 ;
        RECT 19.935 48.125 26.055 48.295 ;
        RECT 19.935 47.460 20.105 48.125 ;
        RECT 20.895 47.460 21.065 48.125 ;
        RECT 21.855 47.460 22.025 48.125 ;
        RECT 22.815 47.460 22.985 48.125 ;
        RECT 23.775 47.460 23.945 48.125 ;
        RECT 24.735 47.460 24.905 48.125 ;
        RECT 19.905 46.940 20.135 47.460 ;
        RECT 20.865 46.940 21.095 47.460 ;
        RECT 21.825 46.940 22.055 47.460 ;
        RECT 22.785 46.940 23.015 47.460 ;
        RECT 23.745 46.940 23.975 47.460 ;
        RECT 24.705 46.940 24.935 47.460 ;
        RECT 19.905 42.565 20.135 43.925 ;
        RECT 20.865 42.565 21.095 43.925 ;
        RECT 21.825 42.565 22.055 43.925 ;
        RECT 22.785 42.565 23.015 43.925 ;
        RECT 23.745 42.565 23.975 43.925 ;
        RECT 24.705 42.565 24.935 43.925 ;
        RECT 19.935 41.860 20.105 42.565 ;
        RECT 20.895 41.860 21.065 42.565 ;
        RECT 21.855 41.860 22.025 42.565 ;
        RECT 22.815 41.860 22.985 42.565 ;
        RECT 23.775 41.860 23.945 42.565 ;
        RECT 24.735 41.860 24.905 42.565 ;
        RECT 28.415 42.130 28.715 48.395 ;
        RECT 25.885 41.960 28.715 42.130 ;
        RECT 25.885 41.860 26.055 41.960 ;
        RECT 19.935 41.690 26.055 41.860 ;
        RECT 19.935 41.025 20.105 41.690 ;
        RECT 20.895 41.025 21.065 41.690 ;
        RECT 21.855 41.025 22.025 41.690 ;
        RECT 22.815 41.025 22.985 41.690 ;
        RECT 23.775 41.025 23.945 41.690 ;
        RECT 24.735 41.025 24.905 41.690 ;
        RECT 19.905 40.505 20.135 41.025 ;
        RECT 20.865 40.505 21.095 41.025 ;
        RECT 21.825 40.505 22.055 41.025 ;
        RECT 22.785 40.505 23.015 41.025 ;
        RECT 23.745 40.505 23.975 41.025 ;
        RECT 24.705 40.505 24.935 41.025 ;
        RECT 19.905 36.130 20.135 37.490 ;
        RECT 20.865 36.130 21.095 37.490 ;
        RECT 21.825 36.130 22.055 37.490 ;
        RECT 22.785 36.130 23.015 37.490 ;
        RECT 23.745 36.130 23.975 37.490 ;
        RECT 24.705 36.130 24.935 37.490 ;
        RECT 19.935 35.425 20.105 36.130 ;
        RECT 20.895 35.425 21.065 36.130 ;
        RECT 21.855 35.425 22.025 36.130 ;
        RECT 22.815 35.425 22.985 36.130 ;
        RECT 23.775 35.425 23.945 36.130 ;
        RECT 24.735 35.425 24.905 36.130 ;
        RECT 28.415 35.695 28.715 41.960 ;
        RECT 25.885 35.525 28.715 35.695 ;
        RECT 25.885 35.425 26.055 35.525 ;
        RECT 19.935 35.255 26.055 35.425 ;
        RECT 19.935 34.590 20.105 35.255 ;
        RECT 20.895 34.590 21.065 35.255 ;
        RECT 21.855 34.590 22.025 35.255 ;
        RECT 22.815 34.590 22.985 35.255 ;
        RECT 23.775 34.590 23.945 35.255 ;
        RECT 24.735 34.590 24.905 35.255 ;
        RECT 19.905 34.070 20.135 34.590 ;
        RECT 20.865 34.070 21.095 34.590 ;
        RECT 21.825 34.070 22.055 34.590 ;
        RECT 22.785 34.070 23.015 34.590 ;
        RECT 23.745 34.070 23.975 34.590 ;
        RECT 24.705 34.070 24.935 34.590 ;
        RECT 19.905 29.695 20.135 31.055 ;
        RECT 20.865 29.695 21.095 31.055 ;
        RECT 21.825 29.695 22.055 31.055 ;
        RECT 22.785 29.695 23.015 31.055 ;
        RECT 23.745 29.695 23.975 31.055 ;
        RECT 24.705 29.695 24.935 31.055 ;
        RECT 19.935 28.990 20.105 29.695 ;
        RECT 20.895 28.990 21.065 29.695 ;
        RECT 21.855 28.990 22.025 29.695 ;
        RECT 22.815 28.990 22.985 29.695 ;
        RECT 23.775 28.990 23.945 29.695 ;
        RECT 24.735 28.990 24.905 29.695 ;
        RECT 28.415 29.260 28.715 35.525 ;
        RECT 25.885 29.090 28.715 29.260 ;
        RECT 25.885 28.990 26.055 29.090 ;
        RECT 19.935 28.820 26.055 28.990 ;
        RECT 19.935 28.155 20.105 28.820 ;
        RECT 20.895 28.155 21.065 28.820 ;
        RECT 21.855 28.155 22.025 28.820 ;
        RECT 22.815 28.155 22.985 28.820 ;
        RECT 23.775 28.155 23.945 28.820 ;
        RECT 24.735 28.155 24.905 28.820 ;
        RECT 19.905 27.635 20.135 28.155 ;
        RECT 20.865 27.635 21.095 28.155 ;
        RECT 21.825 27.635 22.055 28.155 ;
        RECT 22.785 27.635 23.015 28.155 ;
        RECT 23.745 27.635 23.975 28.155 ;
        RECT 24.705 27.635 24.935 28.155 ;
        RECT 19.905 23.260 20.135 24.620 ;
        RECT 20.865 23.260 21.095 24.620 ;
        RECT 21.825 23.260 22.055 24.620 ;
        RECT 22.785 23.260 23.015 24.620 ;
        RECT 23.745 23.260 23.975 24.620 ;
        RECT 24.705 23.260 24.935 24.620 ;
        RECT 19.935 22.555 20.105 23.260 ;
        RECT 20.895 22.555 21.065 23.260 ;
        RECT 21.855 22.555 22.025 23.260 ;
        RECT 22.815 22.555 22.985 23.260 ;
        RECT 23.775 22.555 23.945 23.260 ;
        RECT 24.735 22.555 24.905 23.260 ;
        RECT 28.415 22.825 28.715 29.090 ;
        RECT 25.885 22.655 28.715 22.825 ;
        RECT 25.885 22.555 26.055 22.655 ;
        RECT 19.935 22.385 26.055 22.555 ;
        RECT 19.935 21.720 20.105 22.385 ;
        RECT 20.895 21.720 21.065 22.385 ;
        RECT 21.855 21.720 22.025 22.385 ;
        RECT 22.815 21.720 22.985 22.385 ;
        RECT 23.775 21.720 23.945 22.385 ;
        RECT 24.735 21.720 24.905 22.385 ;
        RECT 19.905 21.200 20.135 21.720 ;
        RECT 20.865 21.200 21.095 21.720 ;
        RECT 21.825 21.200 22.055 21.720 ;
        RECT 22.785 21.200 23.015 21.720 ;
        RECT 23.745 21.200 23.975 21.720 ;
        RECT 24.705 21.200 24.935 21.720 ;
        RECT 19.905 16.825 20.135 18.185 ;
        RECT 20.865 16.825 21.095 18.185 ;
        RECT 21.825 16.825 22.055 18.185 ;
        RECT 22.785 16.825 23.015 18.185 ;
        RECT 23.745 16.825 23.975 18.185 ;
        RECT 24.705 16.825 24.935 18.185 ;
        RECT 19.935 16.120 20.105 16.825 ;
        RECT 20.895 16.120 21.065 16.825 ;
        RECT 21.855 16.120 22.025 16.825 ;
        RECT 22.815 16.120 22.985 16.825 ;
        RECT 23.775 16.120 23.945 16.825 ;
        RECT 24.735 16.120 24.905 16.825 ;
        RECT 28.415 16.390 28.715 22.655 ;
        RECT 25.885 16.220 28.715 16.390 ;
        RECT 25.885 16.120 26.055 16.220 ;
        RECT 19.935 15.950 26.055 16.120 ;
        RECT 19.935 15.285 20.105 15.950 ;
        RECT 20.895 15.285 21.065 15.950 ;
        RECT 21.855 15.285 22.025 15.950 ;
        RECT 22.815 15.285 22.985 15.950 ;
        RECT 23.775 15.285 23.945 15.950 ;
        RECT 24.735 15.285 24.905 15.950 ;
        RECT 19.905 14.765 20.135 15.285 ;
        RECT 20.865 14.765 21.095 15.285 ;
        RECT 21.825 14.765 22.055 15.285 ;
        RECT 22.785 14.765 23.015 15.285 ;
        RECT 23.745 14.765 23.975 15.285 ;
        RECT 24.705 14.765 24.935 15.285 ;
        RECT 19.905 10.390 20.135 11.750 ;
        RECT 20.865 10.390 21.095 11.750 ;
        RECT 21.825 10.390 22.055 11.750 ;
        RECT 22.785 10.390 23.015 11.750 ;
        RECT 23.745 10.390 23.975 11.750 ;
        RECT 24.705 10.390 24.935 11.750 ;
        RECT 19.935 9.685 20.105 10.390 ;
        RECT 20.895 9.685 21.065 10.390 ;
        RECT 21.855 9.685 22.025 10.390 ;
        RECT 22.815 9.685 22.985 10.390 ;
        RECT 23.775 9.685 23.945 10.390 ;
        RECT 24.735 9.685 24.905 10.390 ;
        RECT 28.415 9.955 28.715 16.220 ;
        RECT 25.885 9.785 28.715 9.955 ;
        RECT 25.885 9.685 26.055 9.785 ;
        RECT 19.935 9.515 26.055 9.685 ;
        RECT 19.935 8.850 20.105 9.515 ;
        RECT 20.895 8.850 21.065 9.515 ;
        RECT 21.855 8.850 22.025 9.515 ;
        RECT 22.815 8.850 22.985 9.515 ;
        RECT 23.775 8.850 23.945 9.515 ;
        RECT 24.735 8.850 24.905 9.515 ;
        RECT 19.905 8.330 20.135 8.850 ;
        RECT 20.865 8.330 21.095 8.850 ;
        RECT 21.825 8.330 22.055 8.850 ;
        RECT 22.785 8.330 23.015 8.850 ;
        RECT 23.745 8.330 23.975 8.850 ;
        RECT 24.705 8.330 24.935 8.850 ;
        RECT 19.905 3.955 20.135 5.315 ;
        RECT 20.865 3.955 21.095 5.315 ;
        RECT 21.825 3.955 22.055 5.315 ;
        RECT 22.785 3.955 23.015 5.315 ;
        RECT 23.745 3.955 23.975 5.315 ;
        RECT 24.705 3.955 24.935 5.315 ;
        RECT 19.935 3.250 20.105 3.955 ;
        RECT 20.895 3.250 21.065 3.955 ;
        RECT 21.855 3.250 22.025 3.955 ;
        RECT 22.815 3.250 22.985 3.955 ;
        RECT 23.775 3.250 23.945 3.955 ;
        RECT 24.735 3.250 24.905 3.955 ;
        RECT 28.415 3.520 28.715 9.785 ;
        RECT 25.885 3.350 28.715 3.520 ;
        RECT 25.885 3.250 26.055 3.350 ;
        RECT 19.935 3.080 26.055 3.250 ;
        RECT 19.935 2.415 20.105 3.080 ;
        RECT 20.895 2.415 21.065 3.080 ;
        RECT 21.855 2.415 22.025 3.080 ;
        RECT 22.815 2.415 22.985 3.080 ;
        RECT 23.775 2.415 23.945 3.080 ;
        RECT 24.735 2.415 24.905 3.080 ;
        RECT 19.905 1.895 20.135 2.415 ;
        RECT 20.865 1.895 21.095 2.415 ;
        RECT 21.825 1.895 22.055 2.415 ;
        RECT 22.785 1.895 23.015 2.415 ;
        RECT 23.745 1.895 23.975 2.415 ;
        RECT 24.705 1.895 24.935 2.415 ;
        RECT 28.415 0.725 28.715 3.350 ;
    END
  END out
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 17.920 202.590 19.200 202.650 ;
        RECT 5.765 202.570 25.605 202.590 ;
        RECT 0.865 202.270 25.605 202.570 ;
        RECT 0.865 202.265 26.970 202.270 ;
        RECT 0.865 201.955 27.540 202.265 ;
        RECT 0.865 201.335 27.545 201.955 ;
        RECT 0.865 201.165 27.605 201.335 ;
        RECT 0.865 200.650 27.545 201.165 ;
        RECT 0.865 200.630 19.200 200.650 ;
        RECT 0.865 200.360 7.235 200.630 ;
        RECT 11.630 200.380 19.200 200.630 ;
        RECT 19.235 200.385 27.545 200.650 ;
        RECT 19.235 200.380 25.605 200.385 ;
        RECT 17.920 200.330 19.200 200.380 ;
        RECT 17.920 196.155 19.200 196.215 ;
        RECT 5.765 196.135 25.605 196.155 ;
        RECT 0.865 195.835 25.605 196.135 ;
        RECT 0.865 195.830 26.970 195.835 ;
        RECT 0.865 195.520 27.540 195.830 ;
        RECT 0.865 194.900 27.545 195.520 ;
        RECT 0.865 194.730 27.605 194.900 ;
        RECT 0.865 194.215 27.545 194.730 ;
        RECT 0.865 194.195 19.200 194.215 ;
        RECT 0.865 193.925 7.235 194.195 ;
        RECT 11.630 193.945 19.200 194.195 ;
        RECT 19.235 193.950 27.545 194.215 ;
        RECT 19.235 193.945 25.605 193.950 ;
        RECT 17.920 193.895 19.200 193.945 ;
        RECT 17.920 189.720 19.200 189.780 ;
        RECT 5.765 189.700 25.605 189.720 ;
        RECT 0.865 189.400 25.605 189.700 ;
        RECT 0.865 189.395 26.970 189.400 ;
        RECT 0.865 189.085 27.540 189.395 ;
        RECT 0.865 188.465 27.545 189.085 ;
        RECT 0.865 188.295 27.605 188.465 ;
        RECT 0.865 187.780 27.545 188.295 ;
        RECT 0.865 187.760 19.200 187.780 ;
        RECT 0.865 187.490 7.235 187.760 ;
        RECT 11.630 187.510 19.200 187.760 ;
        RECT 19.235 187.515 27.545 187.780 ;
        RECT 19.235 187.510 25.605 187.515 ;
        RECT 17.920 187.460 19.200 187.510 ;
        RECT 17.920 183.285 19.200 183.345 ;
        RECT 5.765 183.265 25.605 183.285 ;
        RECT 0.865 182.965 25.605 183.265 ;
        RECT 0.865 182.960 26.970 182.965 ;
        RECT 0.865 182.650 27.540 182.960 ;
        RECT 0.865 182.030 27.545 182.650 ;
        RECT 0.865 181.860 27.605 182.030 ;
        RECT 0.865 181.345 27.545 181.860 ;
        RECT 0.865 181.325 19.200 181.345 ;
        RECT 0.865 181.055 7.235 181.325 ;
        RECT 11.630 181.075 19.200 181.325 ;
        RECT 19.235 181.080 27.545 181.345 ;
        RECT 19.235 181.075 25.605 181.080 ;
        RECT 17.920 181.025 19.200 181.075 ;
        RECT 17.920 176.850 19.200 176.910 ;
        RECT 5.765 176.830 25.605 176.850 ;
        RECT 0.865 176.530 25.605 176.830 ;
        RECT 0.865 176.525 26.970 176.530 ;
        RECT 0.865 176.215 27.540 176.525 ;
        RECT 0.865 175.595 27.545 176.215 ;
        RECT 0.865 175.425 27.605 175.595 ;
        RECT 0.865 174.910 27.545 175.425 ;
        RECT 0.865 174.890 19.200 174.910 ;
        RECT 0.865 174.620 7.235 174.890 ;
        RECT 11.630 174.640 19.200 174.890 ;
        RECT 19.235 174.645 27.545 174.910 ;
        RECT 19.235 174.640 25.605 174.645 ;
        RECT 17.920 174.590 19.200 174.640 ;
        RECT 17.920 170.415 19.200 170.475 ;
        RECT 5.765 170.395 25.605 170.415 ;
        RECT 0.865 170.095 25.605 170.395 ;
        RECT 0.865 170.090 26.970 170.095 ;
        RECT 0.865 169.780 27.540 170.090 ;
        RECT 0.865 169.160 27.545 169.780 ;
        RECT 0.865 168.990 27.605 169.160 ;
        RECT 0.865 168.475 27.545 168.990 ;
        RECT 0.865 168.455 19.200 168.475 ;
        RECT 0.865 168.185 7.235 168.455 ;
        RECT 11.630 168.205 19.200 168.455 ;
        RECT 19.235 168.210 27.545 168.475 ;
        RECT 19.235 168.205 25.605 168.210 ;
        RECT 17.920 168.155 19.200 168.205 ;
        RECT 17.920 163.980 19.200 164.040 ;
        RECT 5.765 163.960 25.605 163.980 ;
        RECT 0.865 163.660 25.605 163.960 ;
        RECT 0.865 163.655 26.970 163.660 ;
        RECT 0.865 163.345 27.540 163.655 ;
        RECT 0.865 162.725 27.545 163.345 ;
        RECT 0.865 162.555 27.605 162.725 ;
        RECT 0.865 162.040 27.545 162.555 ;
        RECT 0.865 162.020 19.200 162.040 ;
        RECT 0.865 161.750 7.235 162.020 ;
        RECT 11.630 161.770 19.200 162.020 ;
        RECT 19.235 161.775 27.545 162.040 ;
        RECT 19.235 161.770 25.605 161.775 ;
        RECT 17.920 161.720 19.200 161.770 ;
        RECT 17.920 157.545 19.200 157.605 ;
        RECT 5.765 157.525 25.605 157.545 ;
        RECT 0.865 157.225 25.605 157.525 ;
        RECT 0.865 157.220 26.970 157.225 ;
        RECT 0.865 156.910 27.540 157.220 ;
        RECT 0.865 156.290 27.545 156.910 ;
        RECT 0.865 156.120 27.605 156.290 ;
        RECT 0.865 155.605 27.545 156.120 ;
        RECT 0.865 155.585 19.200 155.605 ;
        RECT 0.865 155.315 7.235 155.585 ;
        RECT 11.630 155.335 19.200 155.585 ;
        RECT 19.235 155.340 27.545 155.605 ;
        RECT 19.235 155.335 25.605 155.340 ;
        RECT 17.920 155.285 19.200 155.335 ;
        RECT 17.920 151.110 19.200 151.170 ;
        RECT 5.765 151.090 25.605 151.110 ;
        RECT 0.865 150.790 25.605 151.090 ;
        RECT 0.865 150.785 26.970 150.790 ;
        RECT 0.865 150.475 27.540 150.785 ;
        RECT 0.865 149.855 27.545 150.475 ;
        RECT 0.865 149.685 27.605 149.855 ;
        RECT 0.865 149.170 27.545 149.685 ;
        RECT 0.865 149.150 19.200 149.170 ;
        RECT 0.865 148.880 7.235 149.150 ;
        RECT 11.630 148.900 19.200 149.150 ;
        RECT 19.235 148.905 27.545 149.170 ;
        RECT 19.235 148.900 25.605 148.905 ;
        RECT 17.920 148.850 19.200 148.900 ;
        RECT 17.920 144.675 19.200 144.735 ;
        RECT 5.765 144.655 25.605 144.675 ;
        RECT 0.865 144.355 25.605 144.655 ;
        RECT 0.865 144.350 26.970 144.355 ;
        RECT 0.865 144.040 27.540 144.350 ;
        RECT 0.865 143.420 27.545 144.040 ;
        RECT 0.865 143.250 27.605 143.420 ;
        RECT 0.865 142.735 27.545 143.250 ;
        RECT 0.865 142.715 19.200 142.735 ;
        RECT 0.865 142.445 7.235 142.715 ;
        RECT 11.630 142.465 19.200 142.715 ;
        RECT 19.235 142.470 27.545 142.735 ;
        RECT 19.235 142.465 25.605 142.470 ;
        RECT 17.920 142.415 19.200 142.465 ;
        RECT 17.920 138.240 19.200 138.300 ;
        RECT 5.765 138.220 25.605 138.240 ;
        RECT 0.865 137.920 25.605 138.220 ;
        RECT 0.865 137.915 26.970 137.920 ;
        RECT 0.865 137.605 27.540 137.915 ;
        RECT 0.865 136.985 27.545 137.605 ;
        RECT 0.865 136.815 27.605 136.985 ;
        RECT 0.865 136.300 27.545 136.815 ;
        RECT 0.865 136.280 19.200 136.300 ;
        RECT 0.865 136.010 7.235 136.280 ;
        RECT 11.630 136.030 19.200 136.280 ;
        RECT 19.235 136.035 27.545 136.300 ;
        RECT 19.235 136.030 25.605 136.035 ;
        RECT 17.920 135.980 19.200 136.030 ;
        RECT 17.920 131.805 19.200 131.865 ;
        RECT 5.765 131.785 25.605 131.805 ;
        RECT 0.865 131.485 25.605 131.785 ;
        RECT 0.865 131.480 26.970 131.485 ;
        RECT 0.865 131.170 27.540 131.480 ;
        RECT 0.865 130.550 27.545 131.170 ;
        RECT 0.865 130.380 27.605 130.550 ;
        RECT 0.865 129.865 27.545 130.380 ;
        RECT 0.865 129.845 19.200 129.865 ;
        RECT 0.865 129.575 7.235 129.845 ;
        RECT 11.630 129.595 19.200 129.845 ;
        RECT 19.235 129.600 27.545 129.865 ;
        RECT 19.235 129.595 25.605 129.600 ;
        RECT 17.920 129.545 19.200 129.595 ;
        RECT 17.920 125.370 19.200 125.430 ;
        RECT 5.765 125.350 25.605 125.370 ;
        RECT 0.865 125.050 25.605 125.350 ;
        RECT 0.865 125.045 26.970 125.050 ;
        RECT 0.865 124.735 27.540 125.045 ;
        RECT 0.865 124.115 27.545 124.735 ;
        RECT 0.865 123.945 27.605 124.115 ;
        RECT 0.865 123.430 27.545 123.945 ;
        RECT 0.865 123.410 19.200 123.430 ;
        RECT 0.865 123.140 7.235 123.410 ;
        RECT 11.630 123.160 19.200 123.410 ;
        RECT 19.235 123.165 27.545 123.430 ;
        RECT 19.235 123.160 25.605 123.165 ;
        RECT 17.920 123.110 19.200 123.160 ;
        RECT 17.920 118.935 19.200 118.995 ;
        RECT 5.765 118.915 25.605 118.935 ;
        RECT 0.865 118.615 25.605 118.915 ;
        RECT 0.865 118.610 26.970 118.615 ;
        RECT 0.865 118.300 27.540 118.610 ;
        RECT 0.865 117.680 27.545 118.300 ;
        RECT 0.865 117.510 27.605 117.680 ;
        RECT 0.865 116.995 27.545 117.510 ;
        RECT 0.865 116.975 19.200 116.995 ;
        RECT 0.865 116.705 7.235 116.975 ;
        RECT 11.630 116.725 19.200 116.975 ;
        RECT 19.235 116.730 27.545 116.995 ;
        RECT 19.235 116.725 25.605 116.730 ;
        RECT 17.920 116.675 19.200 116.725 ;
        RECT 17.920 112.500 19.200 112.560 ;
        RECT 5.765 112.480 25.605 112.500 ;
        RECT 0.865 112.180 25.605 112.480 ;
        RECT 0.865 112.175 26.970 112.180 ;
        RECT 0.865 111.865 27.540 112.175 ;
        RECT 0.865 111.245 27.545 111.865 ;
        RECT 0.865 111.075 27.605 111.245 ;
        RECT 0.865 110.560 27.545 111.075 ;
        RECT 0.865 110.540 19.200 110.560 ;
        RECT 0.865 110.270 7.235 110.540 ;
        RECT 11.630 110.290 19.200 110.540 ;
        RECT 19.235 110.295 27.545 110.560 ;
        RECT 19.235 110.290 25.605 110.295 ;
        RECT 17.920 110.240 19.200 110.290 ;
        RECT 17.920 106.065 19.200 106.125 ;
        RECT 5.765 106.045 25.605 106.065 ;
        RECT 0.865 105.745 25.605 106.045 ;
        RECT 0.865 105.740 26.970 105.745 ;
        RECT 0.865 105.430 27.540 105.740 ;
        RECT 0.865 104.810 27.545 105.430 ;
        RECT 0.865 104.640 27.605 104.810 ;
        RECT 0.865 104.125 27.545 104.640 ;
        RECT 0.865 104.105 19.200 104.125 ;
        RECT 0.865 103.835 7.235 104.105 ;
        RECT 11.630 103.855 19.200 104.105 ;
        RECT 19.235 103.860 27.545 104.125 ;
        RECT 19.235 103.855 25.605 103.860 ;
        RECT 17.920 103.805 19.200 103.855 ;
        RECT 17.920 99.630 19.200 99.690 ;
        RECT 5.765 99.610 25.605 99.630 ;
        RECT 0.865 99.310 25.605 99.610 ;
        RECT 0.865 99.305 26.970 99.310 ;
        RECT 0.865 98.995 27.540 99.305 ;
        RECT 0.865 98.375 27.545 98.995 ;
        RECT 0.865 98.205 27.605 98.375 ;
        RECT 0.865 97.690 27.545 98.205 ;
        RECT 0.865 97.670 19.200 97.690 ;
        RECT 0.865 97.400 7.235 97.670 ;
        RECT 11.630 97.420 19.200 97.670 ;
        RECT 19.235 97.425 27.545 97.690 ;
        RECT 19.235 97.420 25.605 97.425 ;
        RECT 17.920 97.370 19.200 97.420 ;
        RECT 17.920 93.195 19.200 93.255 ;
        RECT 5.765 93.175 25.605 93.195 ;
        RECT 0.865 92.875 25.605 93.175 ;
        RECT 0.865 92.870 26.970 92.875 ;
        RECT 0.865 92.560 27.540 92.870 ;
        RECT 0.865 91.940 27.545 92.560 ;
        RECT 0.865 91.770 27.605 91.940 ;
        RECT 0.865 91.255 27.545 91.770 ;
        RECT 0.865 91.235 19.200 91.255 ;
        RECT 0.865 90.965 7.235 91.235 ;
        RECT 11.630 90.985 19.200 91.235 ;
        RECT 19.235 90.990 27.545 91.255 ;
        RECT 19.235 90.985 25.605 90.990 ;
        RECT 17.920 90.935 19.200 90.985 ;
        RECT 17.920 86.760 19.200 86.820 ;
        RECT 5.765 86.740 25.605 86.760 ;
        RECT 0.865 86.440 25.605 86.740 ;
        RECT 0.865 86.435 26.970 86.440 ;
        RECT 0.865 86.125 27.540 86.435 ;
        RECT 0.865 85.505 27.545 86.125 ;
        RECT 0.865 85.335 27.605 85.505 ;
        RECT 0.865 84.820 27.545 85.335 ;
        RECT 0.865 84.800 19.200 84.820 ;
        RECT 0.865 84.530 7.235 84.800 ;
        RECT 11.630 84.550 19.200 84.800 ;
        RECT 19.235 84.555 27.545 84.820 ;
        RECT 19.235 84.550 25.605 84.555 ;
        RECT 17.920 84.500 19.200 84.550 ;
        RECT 17.920 80.325 19.200 80.385 ;
        RECT 5.765 80.305 25.605 80.325 ;
        RECT 0.865 80.005 25.605 80.305 ;
        RECT 0.865 80.000 26.970 80.005 ;
        RECT 0.865 79.690 27.540 80.000 ;
        RECT 0.865 79.070 27.545 79.690 ;
        RECT 0.865 78.900 27.605 79.070 ;
        RECT 0.865 78.385 27.545 78.900 ;
        RECT 0.865 78.365 19.200 78.385 ;
        RECT 0.865 78.095 7.235 78.365 ;
        RECT 11.630 78.115 19.200 78.365 ;
        RECT 19.235 78.120 27.545 78.385 ;
        RECT 19.235 78.115 25.605 78.120 ;
        RECT 17.920 78.065 19.200 78.115 ;
        RECT 17.920 73.890 19.200 73.950 ;
        RECT 5.765 73.870 25.605 73.890 ;
        RECT 0.865 73.570 25.605 73.870 ;
        RECT 0.865 73.565 26.970 73.570 ;
        RECT 0.865 73.255 27.540 73.565 ;
        RECT 0.865 72.635 27.545 73.255 ;
        RECT 0.865 72.465 27.605 72.635 ;
        RECT 0.865 71.950 27.545 72.465 ;
        RECT 0.865 71.930 19.200 71.950 ;
        RECT 0.865 71.660 7.235 71.930 ;
        RECT 11.630 71.680 19.200 71.930 ;
        RECT 19.235 71.685 27.545 71.950 ;
        RECT 19.235 71.680 25.605 71.685 ;
        RECT 17.920 71.630 19.200 71.680 ;
        RECT 17.920 67.455 19.200 67.515 ;
        RECT 5.765 67.435 25.605 67.455 ;
        RECT 0.865 67.135 25.605 67.435 ;
        RECT 0.865 67.130 26.970 67.135 ;
        RECT 0.865 66.820 27.540 67.130 ;
        RECT 0.865 66.200 27.545 66.820 ;
        RECT 0.865 66.030 27.605 66.200 ;
        RECT 0.865 65.515 27.545 66.030 ;
        RECT 0.865 65.495 19.200 65.515 ;
        RECT 0.865 65.225 7.235 65.495 ;
        RECT 11.630 65.245 19.200 65.495 ;
        RECT 19.235 65.250 27.545 65.515 ;
        RECT 19.235 65.245 25.605 65.250 ;
        RECT 17.920 65.195 19.200 65.245 ;
        RECT 17.920 61.020 19.200 61.080 ;
        RECT 5.765 61.000 25.605 61.020 ;
        RECT 0.865 60.700 25.605 61.000 ;
        RECT 0.865 60.695 26.970 60.700 ;
        RECT 0.865 60.385 27.540 60.695 ;
        RECT 0.865 59.765 27.545 60.385 ;
        RECT 0.865 59.595 27.605 59.765 ;
        RECT 0.865 59.080 27.545 59.595 ;
        RECT 0.865 59.060 19.200 59.080 ;
        RECT 0.865 58.790 7.235 59.060 ;
        RECT 11.630 58.810 19.200 59.060 ;
        RECT 19.235 58.815 27.545 59.080 ;
        RECT 19.235 58.810 25.605 58.815 ;
        RECT 17.920 58.760 19.200 58.810 ;
        RECT 17.920 54.585 19.200 54.645 ;
        RECT 5.765 54.565 25.605 54.585 ;
        RECT 0.865 54.265 25.605 54.565 ;
        RECT 0.865 54.260 26.970 54.265 ;
        RECT 0.865 53.950 27.540 54.260 ;
        RECT 0.865 53.330 27.545 53.950 ;
        RECT 0.865 53.160 27.605 53.330 ;
        RECT 0.865 52.645 27.545 53.160 ;
        RECT 0.865 52.625 19.200 52.645 ;
        RECT 0.865 52.355 7.235 52.625 ;
        RECT 11.630 52.375 19.200 52.625 ;
        RECT 19.235 52.380 27.545 52.645 ;
        RECT 19.235 52.375 25.605 52.380 ;
        RECT 17.920 52.325 19.200 52.375 ;
        RECT 17.920 48.150 19.200 48.210 ;
        RECT 5.765 48.130 25.605 48.150 ;
        RECT 0.865 47.830 25.605 48.130 ;
        RECT 0.865 47.825 26.970 47.830 ;
        RECT 0.865 47.515 27.540 47.825 ;
        RECT 0.865 46.895 27.545 47.515 ;
        RECT 0.865 46.725 27.605 46.895 ;
        RECT 0.865 46.210 27.545 46.725 ;
        RECT 0.865 46.190 19.200 46.210 ;
        RECT 0.865 45.920 7.235 46.190 ;
        RECT 11.630 45.940 19.200 46.190 ;
        RECT 19.235 45.945 27.545 46.210 ;
        RECT 19.235 45.940 25.605 45.945 ;
        RECT 17.920 45.890 19.200 45.940 ;
        RECT 17.920 41.715 19.200 41.775 ;
        RECT 5.765 41.695 25.605 41.715 ;
        RECT 0.865 41.395 25.605 41.695 ;
        RECT 0.865 41.390 26.970 41.395 ;
        RECT 0.865 41.080 27.540 41.390 ;
        RECT 0.865 40.460 27.545 41.080 ;
        RECT 0.865 40.290 27.605 40.460 ;
        RECT 0.865 39.775 27.545 40.290 ;
        RECT 0.865 39.755 19.200 39.775 ;
        RECT 0.865 39.485 7.235 39.755 ;
        RECT 11.630 39.505 19.200 39.755 ;
        RECT 19.235 39.510 27.545 39.775 ;
        RECT 19.235 39.505 25.605 39.510 ;
        RECT 17.920 39.455 19.200 39.505 ;
        RECT 17.920 35.280 19.200 35.340 ;
        RECT 5.765 35.260 25.605 35.280 ;
        RECT 0.865 34.960 25.605 35.260 ;
        RECT 0.865 34.955 26.970 34.960 ;
        RECT 0.865 34.645 27.540 34.955 ;
        RECT 0.865 34.025 27.545 34.645 ;
        RECT 0.865 33.855 27.605 34.025 ;
        RECT 0.865 33.340 27.545 33.855 ;
        RECT 0.865 33.320 19.200 33.340 ;
        RECT 0.865 33.050 7.235 33.320 ;
        RECT 11.630 33.070 19.200 33.320 ;
        RECT 19.235 33.075 27.545 33.340 ;
        RECT 19.235 33.070 25.605 33.075 ;
        RECT 17.920 33.020 19.200 33.070 ;
        RECT 17.920 28.845 19.200 28.905 ;
        RECT 5.765 28.825 25.605 28.845 ;
        RECT 0.865 28.525 25.605 28.825 ;
        RECT 0.865 28.520 26.970 28.525 ;
        RECT 0.865 28.210 27.540 28.520 ;
        RECT 0.865 27.590 27.545 28.210 ;
        RECT 0.865 27.420 27.605 27.590 ;
        RECT 0.865 26.905 27.545 27.420 ;
        RECT 0.865 26.885 19.200 26.905 ;
        RECT 0.865 26.615 7.235 26.885 ;
        RECT 11.630 26.635 19.200 26.885 ;
        RECT 19.235 26.640 27.545 26.905 ;
        RECT 19.235 26.635 25.605 26.640 ;
        RECT 17.920 26.585 19.200 26.635 ;
        RECT 17.920 22.410 19.200 22.470 ;
        RECT 5.765 22.390 25.605 22.410 ;
        RECT 0.865 22.090 25.605 22.390 ;
        RECT 0.865 22.085 26.970 22.090 ;
        RECT 0.865 21.775 27.540 22.085 ;
        RECT 0.865 21.155 27.545 21.775 ;
        RECT 0.865 20.985 27.605 21.155 ;
        RECT 0.865 20.470 27.545 20.985 ;
        RECT 0.865 20.450 19.200 20.470 ;
        RECT 0.865 20.180 7.235 20.450 ;
        RECT 11.630 20.200 19.200 20.450 ;
        RECT 19.235 20.205 27.545 20.470 ;
        RECT 19.235 20.200 25.605 20.205 ;
        RECT 17.920 20.150 19.200 20.200 ;
        RECT 17.920 15.975 19.200 16.035 ;
        RECT 5.765 15.955 25.605 15.975 ;
        RECT 0.865 15.655 25.605 15.955 ;
        RECT 0.865 15.650 26.970 15.655 ;
        RECT 0.865 15.340 27.540 15.650 ;
        RECT 0.865 14.720 27.545 15.340 ;
        RECT 0.865 14.550 27.605 14.720 ;
        RECT 0.865 14.035 27.545 14.550 ;
        RECT 0.865 14.015 19.200 14.035 ;
        RECT 0.865 13.745 7.235 14.015 ;
        RECT 11.630 13.765 19.200 14.015 ;
        RECT 19.235 13.770 27.545 14.035 ;
        RECT 19.235 13.765 25.605 13.770 ;
        RECT 17.920 13.715 19.200 13.765 ;
        RECT 17.920 9.540 19.200 9.600 ;
        RECT 5.765 9.520 25.605 9.540 ;
        RECT 0.865 9.220 25.605 9.520 ;
        RECT 0.865 9.215 26.970 9.220 ;
        RECT 0.865 8.905 27.540 9.215 ;
        RECT 0.865 8.285 27.545 8.905 ;
        RECT 0.865 8.115 27.605 8.285 ;
        RECT 0.865 7.600 27.545 8.115 ;
        RECT 0.865 7.580 19.200 7.600 ;
        RECT 0.865 7.310 7.235 7.580 ;
        RECT 11.630 7.330 19.200 7.580 ;
        RECT 19.235 7.335 27.545 7.600 ;
        RECT 19.235 7.330 25.605 7.335 ;
        RECT 17.920 7.280 19.200 7.330 ;
        RECT 17.920 3.105 19.200 3.165 ;
        RECT 5.765 3.085 25.605 3.105 ;
        RECT 0.865 2.785 25.605 3.085 ;
        RECT 0.865 2.780 26.970 2.785 ;
        RECT 0.865 2.470 27.540 2.780 ;
        RECT 0.865 1.850 27.545 2.470 ;
        RECT 0.865 1.680 27.605 1.850 ;
        RECT 0.865 1.165 27.545 1.680 ;
        RECT 0.865 1.145 19.200 1.165 ;
        RECT 0.865 0.875 7.235 1.145 ;
        RECT 11.630 0.895 19.200 1.145 ;
        RECT 19.235 0.900 27.545 1.165 ;
        RECT 19.235 0.895 25.605 0.900 ;
        RECT 17.920 0.845 19.200 0.895 ;
      LAYER li1 ;
        RECT 0.995 202.270 7.105 202.440 ;
        RECT 0.995 200.660 1.165 202.270 ;
        RECT 6.935 200.660 7.105 202.270 ;
        RECT 0.995 200.490 7.105 200.660 ;
        RECT 11.760 202.290 17.870 202.460 ;
        RECT 11.760 200.680 11.930 202.290 ;
        RECT 17.700 200.680 17.870 202.290 ;
        RECT 19.365 202.290 25.475 202.460 ;
        RECT 18.235 201.400 18.405 201.940 ;
        RECT 11.760 200.510 17.870 200.680 ;
        RECT 19.365 200.680 19.535 202.290 ;
        RECT 25.305 200.680 25.475 202.290 ;
        RECT 27.200 201.335 27.430 202.155 ;
        RECT 26.370 201.165 27.750 201.335 ;
        RECT 19.365 200.510 25.475 200.680 ;
        RECT 0.995 195.835 7.105 196.005 ;
        RECT 0.995 194.225 1.165 195.835 ;
        RECT 6.935 194.225 7.105 195.835 ;
        RECT 0.995 194.055 7.105 194.225 ;
        RECT 11.760 195.855 17.870 196.025 ;
        RECT 11.760 194.245 11.930 195.855 ;
        RECT 17.700 194.245 17.870 195.855 ;
        RECT 19.365 195.855 25.475 196.025 ;
        RECT 18.235 194.965 18.405 195.505 ;
        RECT 11.760 194.075 17.870 194.245 ;
        RECT 19.365 194.245 19.535 195.855 ;
        RECT 25.305 194.245 25.475 195.855 ;
        RECT 27.200 194.900 27.430 195.720 ;
        RECT 26.370 194.730 27.750 194.900 ;
        RECT 19.365 194.075 25.475 194.245 ;
        RECT 0.995 189.400 7.105 189.570 ;
        RECT 0.995 187.790 1.165 189.400 ;
        RECT 6.935 187.790 7.105 189.400 ;
        RECT 0.995 187.620 7.105 187.790 ;
        RECT 11.760 189.420 17.870 189.590 ;
        RECT 11.760 187.810 11.930 189.420 ;
        RECT 17.700 187.810 17.870 189.420 ;
        RECT 19.365 189.420 25.475 189.590 ;
        RECT 18.235 188.530 18.405 189.070 ;
        RECT 11.760 187.640 17.870 187.810 ;
        RECT 19.365 187.810 19.535 189.420 ;
        RECT 25.305 187.810 25.475 189.420 ;
        RECT 27.200 188.465 27.430 189.285 ;
        RECT 26.370 188.295 27.750 188.465 ;
        RECT 19.365 187.640 25.475 187.810 ;
        RECT 0.995 182.965 7.105 183.135 ;
        RECT 0.995 181.355 1.165 182.965 ;
        RECT 6.935 181.355 7.105 182.965 ;
        RECT 0.995 181.185 7.105 181.355 ;
        RECT 11.760 182.985 17.870 183.155 ;
        RECT 11.760 181.375 11.930 182.985 ;
        RECT 17.700 181.375 17.870 182.985 ;
        RECT 19.365 182.985 25.475 183.155 ;
        RECT 18.235 182.095 18.405 182.635 ;
        RECT 11.760 181.205 17.870 181.375 ;
        RECT 19.365 181.375 19.535 182.985 ;
        RECT 25.305 181.375 25.475 182.985 ;
        RECT 27.200 182.030 27.430 182.850 ;
        RECT 26.370 181.860 27.750 182.030 ;
        RECT 19.365 181.205 25.475 181.375 ;
        RECT 0.995 176.530 7.105 176.700 ;
        RECT 0.995 174.920 1.165 176.530 ;
        RECT 6.935 174.920 7.105 176.530 ;
        RECT 0.995 174.750 7.105 174.920 ;
        RECT 11.760 176.550 17.870 176.720 ;
        RECT 11.760 174.940 11.930 176.550 ;
        RECT 17.700 174.940 17.870 176.550 ;
        RECT 19.365 176.550 25.475 176.720 ;
        RECT 18.235 175.660 18.405 176.200 ;
        RECT 11.760 174.770 17.870 174.940 ;
        RECT 19.365 174.940 19.535 176.550 ;
        RECT 25.305 174.940 25.475 176.550 ;
        RECT 27.200 175.595 27.430 176.415 ;
        RECT 26.370 175.425 27.750 175.595 ;
        RECT 19.365 174.770 25.475 174.940 ;
        RECT 0.995 170.095 7.105 170.265 ;
        RECT 0.995 168.485 1.165 170.095 ;
        RECT 6.935 168.485 7.105 170.095 ;
        RECT 0.995 168.315 7.105 168.485 ;
        RECT 11.760 170.115 17.870 170.285 ;
        RECT 11.760 168.505 11.930 170.115 ;
        RECT 17.700 168.505 17.870 170.115 ;
        RECT 19.365 170.115 25.475 170.285 ;
        RECT 18.235 169.225 18.405 169.765 ;
        RECT 11.760 168.335 17.870 168.505 ;
        RECT 19.365 168.505 19.535 170.115 ;
        RECT 25.305 168.505 25.475 170.115 ;
        RECT 27.200 169.160 27.430 169.980 ;
        RECT 26.370 168.990 27.750 169.160 ;
        RECT 19.365 168.335 25.475 168.505 ;
        RECT 0.995 163.660 7.105 163.830 ;
        RECT 0.995 162.050 1.165 163.660 ;
        RECT 6.935 162.050 7.105 163.660 ;
        RECT 0.995 161.880 7.105 162.050 ;
        RECT 11.760 163.680 17.870 163.850 ;
        RECT 11.760 162.070 11.930 163.680 ;
        RECT 17.700 162.070 17.870 163.680 ;
        RECT 19.365 163.680 25.475 163.850 ;
        RECT 18.235 162.790 18.405 163.330 ;
        RECT 11.760 161.900 17.870 162.070 ;
        RECT 19.365 162.070 19.535 163.680 ;
        RECT 25.305 162.070 25.475 163.680 ;
        RECT 27.200 162.725 27.430 163.545 ;
        RECT 26.370 162.555 27.750 162.725 ;
        RECT 19.365 161.900 25.475 162.070 ;
        RECT 0.995 157.225 7.105 157.395 ;
        RECT 0.995 155.615 1.165 157.225 ;
        RECT 6.935 155.615 7.105 157.225 ;
        RECT 0.995 155.445 7.105 155.615 ;
        RECT 11.760 157.245 17.870 157.415 ;
        RECT 11.760 155.635 11.930 157.245 ;
        RECT 17.700 155.635 17.870 157.245 ;
        RECT 19.365 157.245 25.475 157.415 ;
        RECT 18.235 156.355 18.405 156.895 ;
        RECT 11.760 155.465 17.870 155.635 ;
        RECT 19.365 155.635 19.535 157.245 ;
        RECT 25.305 155.635 25.475 157.245 ;
        RECT 27.200 156.290 27.430 157.110 ;
        RECT 26.370 156.120 27.750 156.290 ;
        RECT 19.365 155.465 25.475 155.635 ;
        RECT 0.995 150.790 7.105 150.960 ;
        RECT 0.995 149.180 1.165 150.790 ;
        RECT 6.935 149.180 7.105 150.790 ;
        RECT 0.995 149.010 7.105 149.180 ;
        RECT 11.760 150.810 17.870 150.980 ;
        RECT 11.760 149.200 11.930 150.810 ;
        RECT 17.700 149.200 17.870 150.810 ;
        RECT 19.365 150.810 25.475 150.980 ;
        RECT 18.235 149.920 18.405 150.460 ;
        RECT 11.760 149.030 17.870 149.200 ;
        RECT 19.365 149.200 19.535 150.810 ;
        RECT 25.305 149.200 25.475 150.810 ;
        RECT 27.200 149.855 27.430 150.675 ;
        RECT 26.370 149.685 27.750 149.855 ;
        RECT 19.365 149.030 25.475 149.200 ;
        RECT 0.995 144.355 7.105 144.525 ;
        RECT 0.995 142.745 1.165 144.355 ;
        RECT 6.935 142.745 7.105 144.355 ;
        RECT 0.995 142.575 7.105 142.745 ;
        RECT 11.760 144.375 17.870 144.545 ;
        RECT 11.760 142.765 11.930 144.375 ;
        RECT 17.700 142.765 17.870 144.375 ;
        RECT 19.365 144.375 25.475 144.545 ;
        RECT 18.235 143.485 18.405 144.025 ;
        RECT 11.760 142.595 17.870 142.765 ;
        RECT 19.365 142.765 19.535 144.375 ;
        RECT 25.305 142.765 25.475 144.375 ;
        RECT 27.200 143.420 27.430 144.240 ;
        RECT 26.370 143.250 27.750 143.420 ;
        RECT 19.365 142.595 25.475 142.765 ;
        RECT 0.995 137.920 7.105 138.090 ;
        RECT 0.995 136.310 1.165 137.920 ;
        RECT 6.935 136.310 7.105 137.920 ;
        RECT 0.995 136.140 7.105 136.310 ;
        RECT 11.760 137.940 17.870 138.110 ;
        RECT 11.760 136.330 11.930 137.940 ;
        RECT 17.700 136.330 17.870 137.940 ;
        RECT 19.365 137.940 25.475 138.110 ;
        RECT 18.235 137.050 18.405 137.590 ;
        RECT 11.760 136.160 17.870 136.330 ;
        RECT 19.365 136.330 19.535 137.940 ;
        RECT 25.305 136.330 25.475 137.940 ;
        RECT 27.200 136.985 27.430 137.805 ;
        RECT 26.370 136.815 27.750 136.985 ;
        RECT 19.365 136.160 25.475 136.330 ;
        RECT 0.995 131.485 7.105 131.655 ;
        RECT 0.995 129.875 1.165 131.485 ;
        RECT 6.935 129.875 7.105 131.485 ;
        RECT 0.995 129.705 7.105 129.875 ;
        RECT 11.760 131.505 17.870 131.675 ;
        RECT 11.760 129.895 11.930 131.505 ;
        RECT 17.700 129.895 17.870 131.505 ;
        RECT 19.365 131.505 25.475 131.675 ;
        RECT 18.235 130.615 18.405 131.155 ;
        RECT 11.760 129.725 17.870 129.895 ;
        RECT 19.365 129.895 19.535 131.505 ;
        RECT 25.305 129.895 25.475 131.505 ;
        RECT 27.200 130.550 27.430 131.370 ;
        RECT 26.370 130.380 27.750 130.550 ;
        RECT 19.365 129.725 25.475 129.895 ;
        RECT 0.995 125.050 7.105 125.220 ;
        RECT 0.995 123.440 1.165 125.050 ;
        RECT 6.935 123.440 7.105 125.050 ;
        RECT 0.995 123.270 7.105 123.440 ;
        RECT 11.760 125.070 17.870 125.240 ;
        RECT 11.760 123.460 11.930 125.070 ;
        RECT 17.700 123.460 17.870 125.070 ;
        RECT 19.365 125.070 25.475 125.240 ;
        RECT 18.235 124.180 18.405 124.720 ;
        RECT 11.760 123.290 17.870 123.460 ;
        RECT 19.365 123.460 19.535 125.070 ;
        RECT 25.305 123.460 25.475 125.070 ;
        RECT 27.200 124.115 27.430 124.935 ;
        RECT 26.370 123.945 27.750 124.115 ;
        RECT 19.365 123.290 25.475 123.460 ;
        RECT 0.995 118.615 7.105 118.785 ;
        RECT 0.995 117.005 1.165 118.615 ;
        RECT 6.935 117.005 7.105 118.615 ;
        RECT 0.995 116.835 7.105 117.005 ;
        RECT 11.760 118.635 17.870 118.805 ;
        RECT 11.760 117.025 11.930 118.635 ;
        RECT 17.700 117.025 17.870 118.635 ;
        RECT 19.365 118.635 25.475 118.805 ;
        RECT 18.235 117.745 18.405 118.285 ;
        RECT 11.760 116.855 17.870 117.025 ;
        RECT 19.365 117.025 19.535 118.635 ;
        RECT 25.305 117.025 25.475 118.635 ;
        RECT 27.200 117.680 27.430 118.500 ;
        RECT 26.370 117.510 27.750 117.680 ;
        RECT 19.365 116.855 25.475 117.025 ;
        RECT 0.995 112.180 7.105 112.350 ;
        RECT 0.995 110.570 1.165 112.180 ;
        RECT 6.935 110.570 7.105 112.180 ;
        RECT 0.995 110.400 7.105 110.570 ;
        RECT 11.760 112.200 17.870 112.370 ;
        RECT 11.760 110.590 11.930 112.200 ;
        RECT 17.700 110.590 17.870 112.200 ;
        RECT 19.365 112.200 25.475 112.370 ;
        RECT 18.235 111.310 18.405 111.850 ;
        RECT 11.760 110.420 17.870 110.590 ;
        RECT 19.365 110.590 19.535 112.200 ;
        RECT 25.305 110.590 25.475 112.200 ;
        RECT 27.200 111.245 27.430 112.065 ;
        RECT 26.370 111.075 27.750 111.245 ;
        RECT 19.365 110.420 25.475 110.590 ;
        RECT 0.995 105.745 7.105 105.915 ;
        RECT 0.995 104.135 1.165 105.745 ;
        RECT 6.935 104.135 7.105 105.745 ;
        RECT 0.995 103.965 7.105 104.135 ;
        RECT 11.760 105.765 17.870 105.935 ;
        RECT 11.760 104.155 11.930 105.765 ;
        RECT 17.700 104.155 17.870 105.765 ;
        RECT 19.365 105.765 25.475 105.935 ;
        RECT 18.235 104.875 18.405 105.415 ;
        RECT 11.760 103.985 17.870 104.155 ;
        RECT 19.365 104.155 19.535 105.765 ;
        RECT 25.305 104.155 25.475 105.765 ;
        RECT 27.200 104.810 27.430 105.630 ;
        RECT 26.370 104.640 27.750 104.810 ;
        RECT 19.365 103.985 25.475 104.155 ;
        RECT 0.995 99.310 7.105 99.480 ;
        RECT 0.995 97.700 1.165 99.310 ;
        RECT 6.935 97.700 7.105 99.310 ;
        RECT 0.995 97.530 7.105 97.700 ;
        RECT 11.760 99.330 17.870 99.500 ;
        RECT 11.760 97.720 11.930 99.330 ;
        RECT 17.700 97.720 17.870 99.330 ;
        RECT 19.365 99.330 25.475 99.500 ;
        RECT 18.235 98.440 18.405 98.980 ;
        RECT 11.760 97.550 17.870 97.720 ;
        RECT 19.365 97.720 19.535 99.330 ;
        RECT 25.305 97.720 25.475 99.330 ;
        RECT 27.200 98.375 27.430 99.195 ;
        RECT 26.370 98.205 27.750 98.375 ;
        RECT 19.365 97.550 25.475 97.720 ;
        RECT 0.995 92.875 7.105 93.045 ;
        RECT 0.995 91.265 1.165 92.875 ;
        RECT 6.935 91.265 7.105 92.875 ;
        RECT 0.995 91.095 7.105 91.265 ;
        RECT 11.760 92.895 17.870 93.065 ;
        RECT 11.760 91.285 11.930 92.895 ;
        RECT 17.700 91.285 17.870 92.895 ;
        RECT 19.365 92.895 25.475 93.065 ;
        RECT 18.235 92.005 18.405 92.545 ;
        RECT 11.760 91.115 17.870 91.285 ;
        RECT 19.365 91.285 19.535 92.895 ;
        RECT 25.305 91.285 25.475 92.895 ;
        RECT 27.200 91.940 27.430 92.760 ;
        RECT 26.370 91.770 27.750 91.940 ;
        RECT 19.365 91.115 25.475 91.285 ;
        RECT 0.995 86.440 7.105 86.610 ;
        RECT 0.995 84.830 1.165 86.440 ;
        RECT 6.935 84.830 7.105 86.440 ;
        RECT 0.995 84.660 7.105 84.830 ;
        RECT 11.760 86.460 17.870 86.630 ;
        RECT 11.760 84.850 11.930 86.460 ;
        RECT 17.700 84.850 17.870 86.460 ;
        RECT 19.365 86.460 25.475 86.630 ;
        RECT 18.235 85.570 18.405 86.110 ;
        RECT 11.760 84.680 17.870 84.850 ;
        RECT 19.365 84.850 19.535 86.460 ;
        RECT 25.305 84.850 25.475 86.460 ;
        RECT 27.200 85.505 27.430 86.325 ;
        RECT 26.370 85.335 27.750 85.505 ;
        RECT 19.365 84.680 25.475 84.850 ;
        RECT 0.995 80.005 7.105 80.175 ;
        RECT 0.995 78.395 1.165 80.005 ;
        RECT 6.935 78.395 7.105 80.005 ;
        RECT 0.995 78.225 7.105 78.395 ;
        RECT 11.760 80.025 17.870 80.195 ;
        RECT 11.760 78.415 11.930 80.025 ;
        RECT 17.700 78.415 17.870 80.025 ;
        RECT 19.365 80.025 25.475 80.195 ;
        RECT 18.235 79.135 18.405 79.675 ;
        RECT 11.760 78.245 17.870 78.415 ;
        RECT 19.365 78.415 19.535 80.025 ;
        RECT 25.305 78.415 25.475 80.025 ;
        RECT 27.200 79.070 27.430 79.890 ;
        RECT 26.370 78.900 27.750 79.070 ;
        RECT 19.365 78.245 25.475 78.415 ;
        RECT 0.995 73.570 7.105 73.740 ;
        RECT 0.995 71.960 1.165 73.570 ;
        RECT 6.935 71.960 7.105 73.570 ;
        RECT 0.995 71.790 7.105 71.960 ;
        RECT 11.760 73.590 17.870 73.760 ;
        RECT 11.760 71.980 11.930 73.590 ;
        RECT 17.700 71.980 17.870 73.590 ;
        RECT 19.365 73.590 25.475 73.760 ;
        RECT 18.235 72.700 18.405 73.240 ;
        RECT 11.760 71.810 17.870 71.980 ;
        RECT 19.365 71.980 19.535 73.590 ;
        RECT 25.305 71.980 25.475 73.590 ;
        RECT 27.200 72.635 27.430 73.455 ;
        RECT 26.370 72.465 27.750 72.635 ;
        RECT 19.365 71.810 25.475 71.980 ;
        RECT 0.995 67.135 7.105 67.305 ;
        RECT 0.995 65.525 1.165 67.135 ;
        RECT 6.935 65.525 7.105 67.135 ;
        RECT 0.995 65.355 7.105 65.525 ;
        RECT 11.760 67.155 17.870 67.325 ;
        RECT 11.760 65.545 11.930 67.155 ;
        RECT 17.700 65.545 17.870 67.155 ;
        RECT 19.365 67.155 25.475 67.325 ;
        RECT 18.235 66.265 18.405 66.805 ;
        RECT 11.760 65.375 17.870 65.545 ;
        RECT 19.365 65.545 19.535 67.155 ;
        RECT 25.305 65.545 25.475 67.155 ;
        RECT 27.200 66.200 27.430 67.020 ;
        RECT 26.370 66.030 27.750 66.200 ;
        RECT 19.365 65.375 25.475 65.545 ;
        RECT 0.995 60.700 7.105 60.870 ;
        RECT 0.995 59.090 1.165 60.700 ;
        RECT 6.935 59.090 7.105 60.700 ;
        RECT 0.995 58.920 7.105 59.090 ;
        RECT 11.760 60.720 17.870 60.890 ;
        RECT 11.760 59.110 11.930 60.720 ;
        RECT 17.700 59.110 17.870 60.720 ;
        RECT 19.365 60.720 25.475 60.890 ;
        RECT 18.235 59.830 18.405 60.370 ;
        RECT 11.760 58.940 17.870 59.110 ;
        RECT 19.365 59.110 19.535 60.720 ;
        RECT 25.305 59.110 25.475 60.720 ;
        RECT 27.200 59.765 27.430 60.585 ;
        RECT 26.370 59.595 27.750 59.765 ;
        RECT 19.365 58.940 25.475 59.110 ;
        RECT 0.995 54.265 7.105 54.435 ;
        RECT 0.995 52.655 1.165 54.265 ;
        RECT 6.935 52.655 7.105 54.265 ;
        RECT 0.995 52.485 7.105 52.655 ;
        RECT 11.760 54.285 17.870 54.455 ;
        RECT 11.760 52.675 11.930 54.285 ;
        RECT 17.700 52.675 17.870 54.285 ;
        RECT 19.365 54.285 25.475 54.455 ;
        RECT 18.235 53.395 18.405 53.935 ;
        RECT 11.760 52.505 17.870 52.675 ;
        RECT 19.365 52.675 19.535 54.285 ;
        RECT 25.305 52.675 25.475 54.285 ;
        RECT 27.200 53.330 27.430 54.150 ;
        RECT 26.370 53.160 27.750 53.330 ;
        RECT 19.365 52.505 25.475 52.675 ;
        RECT 0.995 47.830 7.105 48.000 ;
        RECT 0.995 46.220 1.165 47.830 ;
        RECT 6.935 46.220 7.105 47.830 ;
        RECT 0.995 46.050 7.105 46.220 ;
        RECT 11.760 47.850 17.870 48.020 ;
        RECT 11.760 46.240 11.930 47.850 ;
        RECT 17.700 46.240 17.870 47.850 ;
        RECT 19.365 47.850 25.475 48.020 ;
        RECT 18.235 46.960 18.405 47.500 ;
        RECT 11.760 46.070 17.870 46.240 ;
        RECT 19.365 46.240 19.535 47.850 ;
        RECT 25.305 46.240 25.475 47.850 ;
        RECT 27.200 46.895 27.430 47.715 ;
        RECT 26.370 46.725 27.750 46.895 ;
        RECT 19.365 46.070 25.475 46.240 ;
        RECT 0.995 41.395 7.105 41.565 ;
        RECT 0.995 39.785 1.165 41.395 ;
        RECT 6.935 39.785 7.105 41.395 ;
        RECT 0.995 39.615 7.105 39.785 ;
        RECT 11.760 41.415 17.870 41.585 ;
        RECT 11.760 39.805 11.930 41.415 ;
        RECT 17.700 39.805 17.870 41.415 ;
        RECT 19.365 41.415 25.475 41.585 ;
        RECT 18.235 40.525 18.405 41.065 ;
        RECT 11.760 39.635 17.870 39.805 ;
        RECT 19.365 39.805 19.535 41.415 ;
        RECT 25.305 39.805 25.475 41.415 ;
        RECT 27.200 40.460 27.430 41.280 ;
        RECT 26.370 40.290 27.750 40.460 ;
        RECT 19.365 39.635 25.475 39.805 ;
        RECT 0.995 34.960 7.105 35.130 ;
        RECT 0.995 33.350 1.165 34.960 ;
        RECT 6.935 33.350 7.105 34.960 ;
        RECT 0.995 33.180 7.105 33.350 ;
        RECT 11.760 34.980 17.870 35.150 ;
        RECT 11.760 33.370 11.930 34.980 ;
        RECT 17.700 33.370 17.870 34.980 ;
        RECT 19.365 34.980 25.475 35.150 ;
        RECT 18.235 34.090 18.405 34.630 ;
        RECT 11.760 33.200 17.870 33.370 ;
        RECT 19.365 33.370 19.535 34.980 ;
        RECT 25.305 33.370 25.475 34.980 ;
        RECT 27.200 34.025 27.430 34.845 ;
        RECT 26.370 33.855 27.750 34.025 ;
        RECT 19.365 33.200 25.475 33.370 ;
        RECT 0.995 28.525 7.105 28.695 ;
        RECT 0.995 26.915 1.165 28.525 ;
        RECT 6.935 26.915 7.105 28.525 ;
        RECT 0.995 26.745 7.105 26.915 ;
        RECT 11.760 28.545 17.870 28.715 ;
        RECT 11.760 26.935 11.930 28.545 ;
        RECT 17.700 26.935 17.870 28.545 ;
        RECT 19.365 28.545 25.475 28.715 ;
        RECT 18.235 27.655 18.405 28.195 ;
        RECT 11.760 26.765 17.870 26.935 ;
        RECT 19.365 26.935 19.535 28.545 ;
        RECT 25.305 26.935 25.475 28.545 ;
        RECT 27.200 27.590 27.430 28.410 ;
        RECT 26.370 27.420 27.750 27.590 ;
        RECT 19.365 26.765 25.475 26.935 ;
        RECT 0.995 22.090 7.105 22.260 ;
        RECT 0.995 20.480 1.165 22.090 ;
        RECT 6.935 20.480 7.105 22.090 ;
        RECT 0.995 20.310 7.105 20.480 ;
        RECT 11.760 22.110 17.870 22.280 ;
        RECT 11.760 20.500 11.930 22.110 ;
        RECT 17.700 20.500 17.870 22.110 ;
        RECT 19.365 22.110 25.475 22.280 ;
        RECT 18.235 21.220 18.405 21.760 ;
        RECT 11.760 20.330 17.870 20.500 ;
        RECT 19.365 20.500 19.535 22.110 ;
        RECT 25.305 20.500 25.475 22.110 ;
        RECT 27.200 21.155 27.430 21.975 ;
        RECT 26.370 20.985 27.750 21.155 ;
        RECT 19.365 20.330 25.475 20.500 ;
        RECT 0.995 15.655 7.105 15.825 ;
        RECT 0.995 14.045 1.165 15.655 ;
        RECT 6.935 14.045 7.105 15.655 ;
        RECT 0.995 13.875 7.105 14.045 ;
        RECT 11.760 15.675 17.870 15.845 ;
        RECT 11.760 14.065 11.930 15.675 ;
        RECT 17.700 14.065 17.870 15.675 ;
        RECT 19.365 15.675 25.475 15.845 ;
        RECT 18.235 14.785 18.405 15.325 ;
        RECT 11.760 13.895 17.870 14.065 ;
        RECT 19.365 14.065 19.535 15.675 ;
        RECT 25.305 14.065 25.475 15.675 ;
        RECT 27.200 14.720 27.430 15.540 ;
        RECT 26.370 14.550 27.750 14.720 ;
        RECT 19.365 13.895 25.475 14.065 ;
        RECT 0.995 9.220 7.105 9.390 ;
        RECT 0.995 7.610 1.165 9.220 ;
        RECT 6.935 7.610 7.105 9.220 ;
        RECT 0.995 7.440 7.105 7.610 ;
        RECT 11.760 9.240 17.870 9.410 ;
        RECT 11.760 7.630 11.930 9.240 ;
        RECT 17.700 7.630 17.870 9.240 ;
        RECT 19.365 9.240 25.475 9.410 ;
        RECT 18.235 8.350 18.405 8.890 ;
        RECT 11.760 7.460 17.870 7.630 ;
        RECT 19.365 7.630 19.535 9.240 ;
        RECT 25.305 7.630 25.475 9.240 ;
        RECT 27.200 8.285 27.430 9.105 ;
        RECT 26.370 8.115 27.750 8.285 ;
        RECT 19.365 7.460 25.475 7.630 ;
        RECT 0.995 2.785 7.105 2.955 ;
        RECT 0.995 1.175 1.165 2.785 ;
        RECT 6.935 1.175 7.105 2.785 ;
        RECT 0.995 1.005 7.105 1.175 ;
        RECT 11.760 2.805 17.870 2.975 ;
        RECT 11.760 1.195 11.930 2.805 ;
        RECT 17.700 1.195 17.870 2.805 ;
        RECT 19.365 2.805 25.475 2.975 ;
        RECT 18.235 1.915 18.405 2.455 ;
        RECT 11.760 1.025 17.870 1.195 ;
        RECT 19.365 1.195 19.535 2.805 ;
        RECT 25.305 1.195 25.475 2.805 ;
        RECT 27.200 1.850 27.430 2.670 ;
        RECT 26.370 1.680 27.750 1.850 ;
        RECT 19.365 1.025 25.475 1.195 ;
      LAYER mcon ;
        RECT 6.935 201.745 7.105 201.915 ;
        RECT 6.935 201.385 7.105 201.555 ;
        RECT 6.935 201.025 7.105 201.195 ;
        RECT 17.700 201.765 17.870 201.935 ;
        RECT 17.700 201.405 17.870 201.575 ;
        RECT 18.235 201.480 18.405 201.860 ;
        RECT 17.700 201.045 17.870 201.215 ;
        RECT 25.305 201.765 25.475 201.935 ;
        RECT 25.305 201.405 25.475 201.575 ;
        RECT 25.305 201.045 25.475 201.215 ;
        RECT 26.515 201.165 26.685 201.335 ;
        RECT 26.975 201.165 27.145 201.335 ;
        RECT 27.435 201.165 27.605 201.335 ;
        RECT 6.935 195.310 7.105 195.480 ;
        RECT 6.935 194.950 7.105 195.120 ;
        RECT 6.935 194.590 7.105 194.760 ;
        RECT 17.700 195.330 17.870 195.500 ;
        RECT 17.700 194.970 17.870 195.140 ;
        RECT 18.235 195.045 18.405 195.425 ;
        RECT 17.700 194.610 17.870 194.780 ;
        RECT 25.305 195.330 25.475 195.500 ;
        RECT 25.305 194.970 25.475 195.140 ;
        RECT 25.305 194.610 25.475 194.780 ;
        RECT 26.515 194.730 26.685 194.900 ;
        RECT 26.975 194.730 27.145 194.900 ;
        RECT 27.435 194.730 27.605 194.900 ;
        RECT 6.935 188.875 7.105 189.045 ;
        RECT 6.935 188.515 7.105 188.685 ;
        RECT 6.935 188.155 7.105 188.325 ;
        RECT 17.700 188.895 17.870 189.065 ;
        RECT 17.700 188.535 17.870 188.705 ;
        RECT 18.235 188.610 18.405 188.990 ;
        RECT 17.700 188.175 17.870 188.345 ;
        RECT 25.305 188.895 25.475 189.065 ;
        RECT 25.305 188.535 25.475 188.705 ;
        RECT 25.305 188.175 25.475 188.345 ;
        RECT 26.515 188.295 26.685 188.465 ;
        RECT 26.975 188.295 27.145 188.465 ;
        RECT 27.435 188.295 27.605 188.465 ;
        RECT 6.935 182.440 7.105 182.610 ;
        RECT 6.935 182.080 7.105 182.250 ;
        RECT 6.935 181.720 7.105 181.890 ;
        RECT 17.700 182.460 17.870 182.630 ;
        RECT 17.700 182.100 17.870 182.270 ;
        RECT 18.235 182.175 18.405 182.555 ;
        RECT 17.700 181.740 17.870 181.910 ;
        RECT 25.305 182.460 25.475 182.630 ;
        RECT 25.305 182.100 25.475 182.270 ;
        RECT 25.305 181.740 25.475 181.910 ;
        RECT 26.515 181.860 26.685 182.030 ;
        RECT 26.975 181.860 27.145 182.030 ;
        RECT 27.435 181.860 27.605 182.030 ;
        RECT 6.935 176.005 7.105 176.175 ;
        RECT 6.935 175.645 7.105 175.815 ;
        RECT 6.935 175.285 7.105 175.455 ;
        RECT 17.700 176.025 17.870 176.195 ;
        RECT 17.700 175.665 17.870 175.835 ;
        RECT 18.235 175.740 18.405 176.120 ;
        RECT 17.700 175.305 17.870 175.475 ;
        RECT 25.305 176.025 25.475 176.195 ;
        RECT 25.305 175.665 25.475 175.835 ;
        RECT 25.305 175.305 25.475 175.475 ;
        RECT 26.515 175.425 26.685 175.595 ;
        RECT 26.975 175.425 27.145 175.595 ;
        RECT 27.435 175.425 27.605 175.595 ;
        RECT 6.935 169.570 7.105 169.740 ;
        RECT 6.935 169.210 7.105 169.380 ;
        RECT 6.935 168.850 7.105 169.020 ;
        RECT 17.700 169.590 17.870 169.760 ;
        RECT 17.700 169.230 17.870 169.400 ;
        RECT 18.235 169.305 18.405 169.685 ;
        RECT 17.700 168.870 17.870 169.040 ;
        RECT 25.305 169.590 25.475 169.760 ;
        RECT 25.305 169.230 25.475 169.400 ;
        RECT 25.305 168.870 25.475 169.040 ;
        RECT 26.515 168.990 26.685 169.160 ;
        RECT 26.975 168.990 27.145 169.160 ;
        RECT 27.435 168.990 27.605 169.160 ;
        RECT 6.935 163.135 7.105 163.305 ;
        RECT 6.935 162.775 7.105 162.945 ;
        RECT 6.935 162.415 7.105 162.585 ;
        RECT 17.700 163.155 17.870 163.325 ;
        RECT 17.700 162.795 17.870 162.965 ;
        RECT 18.235 162.870 18.405 163.250 ;
        RECT 17.700 162.435 17.870 162.605 ;
        RECT 25.305 163.155 25.475 163.325 ;
        RECT 25.305 162.795 25.475 162.965 ;
        RECT 25.305 162.435 25.475 162.605 ;
        RECT 26.515 162.555 26.685 162.725 ;
        RECT 26.975 162.555 27.145 162.725 ;
        RECT 27.435 162.555 27.605 162.725 ;
        RECT 6.935 156.700 7.105 156.870 ;
        RECT 6.935 156.340 7.105 156.510 ;
        RECT 6.935 155.980 7.105 156.150 ;
        RECT 17.700 156.720 17.870 156.890 ;
        RECT 17.700 156.360 17.870 156.530 ;
        RECT 18.235 156.435 18.405 156.815 ;
        RECT 17.700 156.000 17.870 156.170 ;
        RECT 25.305 156.720 25.475 156.890 ;
        RECT 25.305 156.360 25.475 156.530 ;
        RECT 25.305 156.000 25.475 156.170 ;
        RECT 26.515 156.120 26.685 156.290 ;
        RECT 26.975 156.120 27.145 156.290 ;
        RECT 27.435 156.120 27.605 156.290 ;
        RECT 6.935 150.265 7.105 150.435 ;
        RECT 6.935 149.905 7.105 150.075 ;
        RECT 6.935 149.545 7.105 149.715 ;
        RECT 17.700 150.285 17.870 150.455 ;
        RECT 17.700 149.925 17.870 150.095 ;
        RECT 18.235 150.000 18.405 150.380 ;
        RECT 17.700 149.565 17.870 149.735 ;
        RECT 25.305 150.285 25.475 150.455 ;
        RECT 25.305 149.925 25.475 150.095 ;
        RECT 25.305 149.565 25.475 149.735 ;
        RECT 26.515 149.685 26.685 149.855 ;
        RECT 26.975 149.685 27.145 149.855 ;
        RECT 27.435 149.685 27.605 149.855 ;
        RECT 6.935 143.830 7.105 144.000 ;
        RECT 6.935 143.470 7.105 143.640 ;
        RECT 6.935 143.110 7.105 143.280 ;
        RECT 17.700 143.850 17.870 144.020 ;
        RECT 17.700 143.490 17.870 143.660 ;
        RECT 18.235 143.565 18.405 143.945 ;
        RECT 17.700 143.130 17.870 143.300 ;
        RECT 25.305 143.850 25.475 144.020 ;
        RECT 25.305 143.490 25.475 143.660 ;
        RECT 25.305 143.130 25.475 143.300 ;
        RECT 26.515 143.250 26.685 143.420 ;
        RECT 26.975 143.250 27.145 143.420 ;
        RECT 27.435 143.250 27.605 143.420 ;
        RECT 6.935 137.395 7.105 137.565 ;
        RECT 6.935 137.035 7.105 137.205 ;
        RECT 6.935 136.675 7.105 136.845 ;
        RECT 17.700 137.415 17.870 137.585 ;
        RECT 17.700 137.055 17.870 137.225 ;
        RECT 18.235 137.130 18.405 137.510 ;
        RECT 17.700 136.695 17.870 136.865 ;
        RECT 25.305 137.415 25.475 137.585 ;
        RECT 25.305 137.055 25.475 137.225 ;
        RECT 25.305 136.695 25.475 136.865 ;
        RECT 26.515 136.815 26.685 136.985 ;
        RECT 26.975 136.815 27.145 136.985 ;
        RECT 27.435 136.815 27.605 136.985 ;
        RECT 6.935 130.960 7.105 131.130 ;
        RECT 6.935 130.600 7.105 130.770 ;
        RECT 6.935 130.240 7.105 130.410 ;
        RECT 17.700 130.980 17.870 131.150 ;
        RECT 17.700 130.620 17.870 130.790 ;
        RECT 18.235 130.695 18.405 131.075 ;
        RECT 17.700 130.260 17.870 130.430 ;
        RECT 25.305 130.980 25.475 131.150 ;
        RECT 25.305 130.620 25.475 130.790 ;
        RECT 25.305 130.260 25.475 130.430 ;
        RECT 26.515 130.380 26.685 130.550 ;
        RECT 26.975 130.380 27.145 130.550 ;
        RECT 27.435 130.380 27.605 130.550 ;
        RECT 6.935 124.525 7.105 124.695 ;
        RECT 6.935 124.165 7.105 124.335 ;
        RECT 6.935 123.805 7.105 123.975 ;
        RECT 17.700 124.545 17.870 124.715 ;
        RECT 17.700 124.185 17.870 124.355 ;
        RECT 18.235 124.260 18.405 124.640 ;
        RECT 17.700 123.825 17.870 123.995 ;
        RECT 25.305 124.545 25.475 124.715 ;
        RECT 25.305 124.185 25.475 124.355 ;
        RECT 25.305 123.825 25.475 123.995 ;
        RECT 26.515 123.945 26.685 124.115 ;
        RECT 26.975 123.945 27.145 124.115 ;
        RECT 27.435 123.945 27.605 124.115 ;
        RECT 6.935 118.090 7.105 118.260 ;
        RECT 6.935 117.730 7.105 117.900 ;
        RECT 6.935 117.370 7.105 117.540 ;
        RECT 17.700 118.110 17.870 118.280 ;
        RECT 17.700 117.750 17.870 117.920 ;
        RECT 18.235 117.825 18.405 118.205 ;
        RECT 17.700 117.390 17.870 117.560 ;
        RECT 25.305 118.110 25.475 118.280 ;
        RECT 25.305 117.750 25.475 117.920 ;
        RECT 25.305 117.390 25.475 117.560 ;
        RECT 26.515 117.510 26.685 117.680 ;
        RECT 26.975 117.510 27.145 117.680 ;
        RECT 27.435 117.510 27.605 117.680 ;
        RECT 6.935 111.655 7.105 111.825 ;
        RECT 6.935 111.295 7.105 111.465 ;
        RECT 6.935 110.935 7.105 111.105 ;
        RECT 17.700 111.675 17.870 111.845 ;
        RECT 17.700 111.315 17.870 111.485 ;
        RECT 18.235 111.390 18.405 111.770 ;
        RECT 17.700 110.955 17.870 111.125 ;
        RECT 25.305 111.675 25.475 111.845 ;
        RECT 25.305 111.315 25.475 111.485 ;
        RECT 25.305 110.955 25.475 111.125 ;
        RECT 26.515 111.075 26.685 111.245 ;
        RECT 26.975 111.075 27.145 111.245 ;
        RECT 27.435 111.075 27.605 111.245 ;
        RECT 6.935 105.220 7.105 105.390 ;
        RECT 6.935 104.860 7.105 105.030 ;
        RECT 6.935 104.500 7.105 104.670 ;
        RECT 17.700 105.240 17.870 105.410 ;
        RECT 17.700 104.880 17.870 105.050 ;
        RECT 18.235 104.955 18.405 105.335 ;
        RECT 17.700 104.520 17.870 104.690 ;
        RECT 25.305 105.240 25.475 105.410 ;
        RECT 25.305 104.880 25.475 105.050 ;
        RECT 25.305 104.520 25.475 104.690 ;
        RECT 26.515 104.640 26.685 104.810 ;
        RECT 26.975 104.640 27.145 104.810 ;
        RECT 27.435 104.640 27.605 104.810 ;
        RECT 6.935 98.785 7.105 98.955 ;
        RECT 6.935 98.425 7.105 98.595 ;
        RECT 6.935 98.065 7.105 98.235 ;
        RECT 17.700 98.805 17.870 98.975 ;
        RECT 17.700 98.445 17.870 98.615 ;
        RECT 18.235 98.520 18.405 98.900 ;
        RECT 17.700 98.085 17.870 98.255 ;
        RECT 25.305 98.805 25.475 98.975 ;
        RECT 25.305 98.445 25.475 98.615 ;
        RECT 25.305 98.085 25.475 98.255 ;
        RECT 26.515 98.205 26.685 98.375 ;
        RECT 26.975 98.205 27.145 98.375 ;
        RECT 27.435 98.205 27.605 98.375 ;
        RECT 6.935 92.350 7.105 92.520 ;
        RECT 6.935 91.990 7.105 92.160 ;
        RECT 6.935 91.630 7.105 91.800 ;
        RECT 17.700 92.370 17.870 92.540 ;
        RECT 17.700 92.010 17.870 92.180 ;
        RECT 18.235 92.085 18.405 92.465 ;
        RECT 17.700 91.650 17.870 91.820 ;
        RECT 25.305 92.370 25.475 92.540 ;
        RECT 25.305 92.010 25.475 92.180 ;
        RECT 25.305 91.650 25.475 91.820 ;
        RECT 26.515 91.770 26.685 91.940 ;
        RECT 26.975 91.770 27.145 91.940 ;
        RECT 27.435 91.770 27.605 91.940 ;
        RECT 6.935 85.915 7.105 86.085 ;
        RECT 6.935 85.555 7.105 85.725 ;
        RECT 6.935 85.195 7.105 85.365 ;
        RECT 17.700 85.935 17.870 86.105 ;
        RECT 17.700 85.575 17.870 85.745 ;
        RECT 18.235 85.650 18.405 86.030 ;
        RECT 17.700 85.215 17.870 85.385 ;
        RECT 25.305 85.935 25.475 86.105 ;
        RECT 25.305 85.575 25.475 85.745 ;
        RECT 25.305 85.215 25.475 85.385 ;
        RECT 26.515 85.335 26.685 85.505 ;
        RECT 26.975 85.335 27.145 85.505 ;
        RECT 27.435 85.335 27.605 85.505 ;
        RECT 6.935 79.480 7.105 79.650 ;
        RECT 6.935 79.120 7.105 79.290 ;
        RECT 6.935 78.760 7.105 78.930 ;
        RECT 17.700 79.500 17.870 79.670 ;
        RECT 17.700 79.140 17.870 79.310 ;
        RECT 18.235 79.215 18.405 79.595 ;
        RECT 17.700 78.780 17.870 78.950 ;
        RECT 25.305 79.500 25.475 79.670 ;
        RECT 25.305 79.140 25.475 79.310 ;
        RECT 25.305 78.780 25.475 78.950 ;
        RECT 26.515 78.900 26.685 79.070 ;
        RECT 26.975 78.900 27.145 79.070 ;
        RECT 27.435 78.900 27.605 79.070 ;
        RECT 6.935 73.045 7.105 73.215 ;
        RECT 6.935 72.685 7.105 72.855 ;
        RECT 6.935 72.325 7.105 72.495 ;
        RECT 17.700 73.065 17.870 73.235 ;
        RECT 17.700 72.705 17.870 72.875 ;
        RECT 18.235 72.780 18.405 73.160 ;
        RECT 17.700 72.345 17.870 72.515 ;
        RECT 25.305 73.065 25.475 73.235 ;
        RECT 25.305 72.705 25.475 72.875 ;
        RECT 25.305 72.345 25.475 72.515 ;
        RECT 26.515 72.465 26.685 72.635 ;
        RECT 26.975 72.465 27.145 72.635 ;
        RECT 27.435 72.465 27.605 72.635 ;
        RECT 6.935 66.610 7.105 66.780 ;
        RECT 6.935 66.250 7.105 66.420 ;
        RECT 6.935 65.890 7.105 66.060 ;
        RECT 17.700 66.630 17.870 66.800 ;
        RECT 17.700 66.270 17.870 66.440 ;
        RECT 18.235 66.345 18.405 66.725 ;
        RECT 17.700 65.910 17.870 66.080 ;
        RECT 25.305 66.630 25.475 66.800 ;
        RECT 25.305 66.270 25.475 66.440 ;
        RECT 25.305 65.910 25.475 66.080 ;
        RECT 26.515 66.030 26.685 66.200 ;
        RECT 26.975 66.030 27.145 66.200 ;
        RECT 27.435 66.030 27.605 66.200 ;
        RECT 6.935 60.175 7.105 60.345 ;
        RECT 6.935 59.815 7.105 59.985 ;
        RECT 6.935 59.455 7.105 59.625 ;
        RECT 17.700 60.195 17.870 60.365 ;
        RECT 17.700 59.835 17.870 60.005 ;
        RECT 18.235 59.910 18.405 60.290 ;
        RECT 17.700 59.475 17.870 59.645 ;
        RECT 25.305 60.195 25.475 60.365 ;
        RECT 25.305 59.835 25.475 60.005 ;
        RECT 25.305 59.475 25.475 59.645 ;
        RECT 26.515 59.595 26.685 59.765 ;
        RECT 26.975 59.595 27.145 59.765 ;
        RECT 27.435 59.595 27.605 59.765 ;
        RECT 6.935 53.740 7.105 53.910 ;
        RECT 6.935 53.380 7.105 53.550 ;
        RECT 6.935 53.020 7.105 53.190 ;
        RECT 17.700 53.760 17.870 53.930 ;
        RECT 17.700 53.400 17.870 53.570 ;
        RECT 18.235 53.475 18.405 53.855 ;
        RECT 17.700 53.040 17.870 53.210 ;
        RECT 25.305 53.760 25.475 53.930 ;
        RECT 25.305 53.400 25.475 53.570 ;
        RECT 25.305 53.040 25.475 53.210 ;
        RECT 26.515 53.160 26.685 53.330 ;
        RECT 26.975 53.160 27.145 53.330 ;
        RECT 27.435 53.160 27.605 53.330 ;
        RECT 6.935 47.305 7.105 47.475 ;
        RECT 6.935 46.945 7.105 47.115 ;
        RECT 6.935 46.585 7.105 46.755 ;
        RECT 17.700 47.325 17.870 47.495 ;
        RECT 17.700 46.965 17.870 47.135 ;
        RECT 18.235 47.040 18.405 47.420 ;
        RECT 17.700 46.605 17.870 46.775 ;
        RECT 25.305 47.325 25.475 47.495 ;
        RECT 25.305 46.965 25.475 47.135 ;
        RECT 25.305 46.605 25.475 46.775 ;
        RECT 26.515 46.725 26.685 46.895 ;
        RECT 26.975 46.725 27.145 46.895 ;
        RECT 27.435 46.725 27.605 46.895 ;
        RECT 6.935 40.870 7.105 41.040 ;
        RECT 6.935 40.510 7.105 40.680 ;
        RECT 6.935 40.150 7.105 40.320 ;
        RECT 17.700 40.890 17.870 41.060 ;
        RECT 17.700 40.530 17.870 40.700 ;
        RECT 18.235 40.605 18.405 40.985 ;
        RECT 17.700 40.170 17.870 40.340 ;
        RECT 25.305 40.890 25.475 41.060 ;
        RECT 25.305 40.530 25.475 40.700 ;
        RECT 25.305 40.170 25.475 40.340 ;
        RECT 26.515 40.290 26.685 40.460 ;
        RECT 26.975 40.290 27.145 40.460 ;
        RECT 27.435 40.290 27.605 40.460 ;
        RECT 6.935 34.435 7.105 34.605 ;
        RECT 6.935 34.075 7.105 34.245 ;
        RECT 6.935 33.715 7.105 33.885 ;
        RECT 17.700 34.455 17.870 34.625 ;
        RECT 17.700 34.095 17.870 34.265 ;
        RECT 18.235 34.170 18.405 34.550 ;
        RECT 17.700 33.735 17.870 33.905 ;
        RECT 25.305 34.455 25.475 34.625 ;
        RECT 25.305 34.095 25.475 34.265 ;
        RECT 25.305 33.735 25.475 33.905 ;
        RECT 26.515 33.855 26.685 34.025 ;
        RECT 26.975 33.855 27.145 34.025 ;
        RECT 27.435 33.855 27.605 34.025 ;
        RECT 6.935 28.000 7.105 28.170 ;
        RECT 6.935 27.640 7.105 27.810 ;
        RECT 6.935 27.280 7.105 27.450 ;
        RECT 17.700 28.020 17.870 28.190 ;
        RECT 17.700 27.660 17.870 27.830 ;
        RECT 18.235 27.735 18.405 28.115 ;
        RECT 17.700 27.300 17.870 27.470 ;
        RECT 25.305 28.020 25.475 28.190 ;
        RECT 25.305 27.660 25.475 27.830 ;
        RECT 25.305 27.300 25.475 27.470 ;
        RECT 26.515 27.420 26.685 27.590 ;
        RECT 26.975 27.420 27.145 27.590 ;
        RECT 27.435 27.420 27.605 27.590 ;
        RECT 6.935 21.565 7.105 21.735 ;
        RECT 6.935 21.205 7.105 21.375 ;
        RECT 6.935 20.845 7.105 21.015 ;
        RECT 17.700 21.585 17.870 21.755 ;
        RECT 17.700 21.225 17.870 21.395 ;
        RECT 18.235 21.300 18.405 21.680 ;
        RECT 17.700 20.865 17.870 21.035 ;
        RECT 25.305 21.585 25.475 21.755 ;
        RECT 25.305 21.225 25.475 21.395 ;
        RECT 25.305 20.865 25.475 21.035 ;
        RECT 26.515 20.985 26.685 21.155 ;
        RECT 26.975 20.985 27.145 21.155 ;
        RECT 27.435 20.985 27.605 21.155 ;
        RECT 6.935 15.130 7.105 15.300 ;
        RECT 6.935 14.770 7.105 14.940 ;
        RECT 6.935 14.410 7.105 14.580 ;
        RECT 17.700 15.150 17.870 15.320 ;
        RECT 17.700 14.790 17.870 14.960 ;
        RECT 18.235 14.865 18.405 15.245 ;
        RECT 17.700 14.430 17.870 14.600 ;
        RECT 25.305 15.150 25.475 15.320 ;
        RECT 25.305 14.790 25.475 14.960 ;
        RECT 25.305 14.430 25.475 14.600 ;
        RECT 26.515 14.550 26.685 14.720 ;
        RECT 26.975 14.550 27.145 14.720 ;
        RECT 27.435 14.550 27.605 14.720 ;
        RECT 6.935 8.695 7.105 8.865 ;
        RECT 6.935 8.335 7.105 8.505 ;
        RECT 6.935 7.975 7.105 8.145 ;
        RECT 17.700 8.715 17.870 8.885 ;
        RECT 17.700 8.355 17.870 8.525 ;
        RECT 18.235 8.430 18.405 8.810 ;
        RECT 17.700 7.995 17.870 8.165 ;
        RECT 25.305 8.715 25.475 8.885 ;
        RECT 25.305 8.355 25.475 8.525 ;
        RECT 25.305 7.995 25.475 8.165 ;
        RECT 26.515 8.115 26.685 8.285 ;
        RECT 26.975 8.115 27.145 8.285 ;
        RECT 27.435 8.115 27.605 8.285 ;
        RECT 6.935 2.260 7.105 2.430 ;
        RECT 6.935 1.900 7.105 2.070 ;
        RECT 6.935 1.540 7.105 1.710 ;
        RECT 17.700 2.280 17.870 2.450 ;
        RECT 17.700 1.920 17.870 2.090 ;
        RECT 18.235 1.995 18.405 2.375 ;
        RECT 17.700 1.560 17.870 1.730 ;
        RECT 25.305 2.280 25.475 2.450 ;
        RECT 25.305 1.920 25.475 2.090 ;
        RECT 25.305 1.560 25.475 1.730 ;
        RECT 26.515 1.680 26.685 1.850 ;
        RECT 26.975 1.680 27.145 1.850 ;
        RECT 27.435 1.680 27.605 1.850 ;
      LAYER met1 ;
        RECT 6.905 201.430 8.650 202.030 ;
        RECT 6.905 200.090 7.135 201.430 ;
        RECT 7.800 201.420 8.650 201.430 ;
        RECT 7.990 201.410 8.650 201.420 ;
        RECT 17.670 201.925 17.900 202.050 ;
        RECT 17.670 201.920 18.400 201.925 ;
        RECT 17.670 201.425 18.435 201.920 ;
        RECT 17.670 200.350 17.900 201.425 ;
        RECT 18.205 201.420 18.435 201.425 ;
        RECT 25.275 201.490 25.505 202.050 ;
        RECT 25.275 201.010 27.750 201.490 ;
        RECT 17.640 200.140 17.910 200.350 ;
        RECT 17.670 200.110 17.900 200.140 ;
        RECT 25.275 200.110 25.505 201.010 ;
        RECT 6.905 194.995 8.650 195.595 ;
        RECT 6.905 193.655 7.135 194.995 ;
        RECT 7.800 194.985 8.650 194.995 ;
        RECT 7.990 194.975 8.650 194.985 ;
        RECT 17.670 195.490 17.900 195.615 ;
        RECT 17.670 195.485 18.400 195.490 ;
        RECT 17.670 194.990 18.435 195.485 ;
        RECT 17.670 193.915 17.900 194.990 ;
        RECT 18.205 194.985 18.435 194.990 ;
        RECT 25.275 195.055 25.505 195.615 ;
        RECT 25.275 194.575 27.750 195.055 ;
        RECT 17.640 193.705 17.910 193.915 ;
        RECT 17.670 193.675 17.900 193.705 ;
        RECT 25.275 193.675 25.505 194.575 ;
        RECT 6.905 188.560 8.650 189.160 ;
        RECT 6.905 187.220 7.135 188.560 ;
        RECT 7.800 188.550 8.650 188.560 ;
        RECT 7.990 188.540 8.650 188.550 ;
        RECT 17.670 189.055 17.900 189.180 ;
        RECT 17.670 189.050 18.400 189.055 ;
        RECT 17.670 188.555 18.435 189.050 ;
        RECT 17.670 187.480 17.900 188.555 ;
        RECT 18.205 188.550 18.435 188.555 ;
        RECT 25.275 188.620 25.505 189.180 ;
        RECT 25.275 188.140 27.750 188.620 ;
        RECT 17.640 187.270 17.910 187.480 ;
        RECT 17.670 187.240 17.900 187.270 ;
        RECT 25.275 187.240 25.505 188.140 ;
        RECT 6.905 182.125 8.650 182.725 ;
        RECT 6.905 180.785 7.135 182.125 ;
        RECT 7.800 182.115 8.650 182.125 ;
        RECT 7.990 182.105 8.650 182.115 ;
        RECT 17.670 182.620 17.900 182.745 ;
        RECT 17.670 182.615 18.400 182.620 ;
        RECT 17.670 182.120 18.435 182.615 ;
        RECT 17.670 181.045 17.900 182.120 ;
        RECT 18.205 182.115 18.435 182.120 ;
        RECT 25.275 182.185 25.505 182.745 ;
        RECT 25.275 181.705 27.750 182.185 ;
        RECT 17.640 180.835 17.910 181.045 ;
        RECT 17.670 180.805 17.900 180.835 ;
        RECT 25.275 180.805 25.505 181.705 ;
        RECT 6.905 175.690 8.650 176.290 ;
        RECT 6.905 174.350 7.135 175.690 ;
        RECT 7.800 175.680 8.650 175.690 ;
        RECT 7.990 175.670 8.650 175.680 ;
        RECT 17.670 176.185 17.900 176.310 ;
        RECT 17.670 176.180 18.400 176.185 ;
        RECT 17.670 175.685 18.435 176.180 ;
        RECT 17.670 174.610 17.900 175.685 ;
        RECT 18.205 175.680 18.435 175.685 ;
        RECT 25.275 175.750 25.505 176.310 ;
        RECT 25.275 175.270 27.750 175.750 ;
        RECT 17.640 174.400 17.910 174.610 ;
        RECT 17.670 174.370 17.900 174.400 ;
        RECT 25.275 174.370 25.505 175.270 ;
        RECT 6.905 169.255 8.650 169.855 ;
        RECT 6.905 167.915 7.135 169.255 ;
        RECT 7.800 169.245 8.650 169.255 ;
        RECT 7.990 169.235 8.650 169.245 ;
        RECT 17.670 169.750 17.900 169.875 ;
        RECT 17.670 169.745 18.400 169.750 ;
        RECT 17.670 169.250 18.435 169.745 ;
        RECT 17.670 168.175 17.900 169.250 ;
        RECT 18.205 169.245 18.435 169.250 ;
        RECT 25.275 169.315 25.505 169.875 ;
        RECT 25.275 168.835 27.750 169.315 ;
        RECT 17.640 167.965 17.910 168.175 ;
        RECT 17.670 167.935 17.900 167.965 ;
        RECT 25.275 167.935 25.505 168.835 ;
        RECT 6.905 162.820 8.650 163.420 ;
        RECT 6.905 161.480 7.135 162.820 ;
        RECT 7.800 162.810 8.650 162.820 ;
        RECT 7.990 162.800 8.650 162.810 ;
        RECT 17.670 163.315 17.900 163.440 ;
        RECT 17.670 163.310 18.400 163.315 ;
        RECT 17.670 162.815 18.435 163.310 ;
        RECT 17.670 161.740 17.900 162.815 ;
        RECT 18.205 162.810 18.435 162.815 ;
        RECT 25.275 162.880 25.505 163.440 ;
        RECT 25.275 162.400 27.750 162.880 ;
        RECT 17.640 161.530 17.910 161.740 ;
        RECT 17.670 161.500 17.900 161.530 ;
        RECT 25.275 161.500 25.505 162.400 ;
        RECT 6.905 156.385 8.650 156.985 ;
        RECT 6.905 155.045 7.135 156.385 ;
        RECT 7.800 156.375 8.650 156.385 ;
        RECT 7.990 156.365 8.650 156.375 ;
        RECT 17.670 156.880 17.900 157.005 ;
        RECT 17.670 156.875 18.400 156.880 ;
        RECT 17.670 156.380 18.435 156.875 ;
        RECT 17.670 155.305 17.900 156.380 ;
        RECT 18.205 156.375 18.435 156.380 ;
        RECT 25.275 156.445 25.505 157.005 ;
        RECT 25.275 155.965 27.750 156.445 ;
        RECT 17.640 155.095 17.910 155.305 ;
        RECT 17.670 155.065 17.900 155.095 ;
        RECT 25.275 155.065 25.505 155.965 ;
        RECT 6.905 149.950 8.650 150.550 ;
        RECT 6.905 148.610 7.135 149.950 ;
        RECT 7.800 149.940 8.650 149.950 ;
        RECT 7.990 149.930 8.650 149.940 ;
        RECT 17.670 150.445 17.900 150.570 ;
        RECT 17.670 150.440 18.400 150.445 ;
        RECT 17.670 149.945 18.435 150.440 ;
        RECT 17.670 148.870 17.900 149.945 ;
        RECT 18.205 149.940 18.435 149.945 ;
        RECT 25.275 150.010 25.505 150.570 ;
        RECT 25.275 149.530 27.750 150.010 ;
        RECT 17.640 148.660 17.910 148.870 ;
        RECT 17.670 148.630 17.900 148.660 ;
        RECT 25.275 148.630 25.505 149.530 ;
        RECT 6.905 143.515 8.650 144.115 ;
        RECT 6.905 142.175 7.135 143.515 ;
        RECT 7.800 143.505 8.650 143.515 ;
        RECT 7.990 143.495 8.650 143.505 ;
        RECT 17.670 144.010 17.900 144.135 ;
        RECT 17.670 144.005 18.400 144.010 ;
        RECT 17.670 143.510 18.435 144.005 ;
        RECT 17.670 142.435 17.900 143.510 ;
        RECT 18.205 143.505 18.435 143.510 ;
        RECT 25.275 143.575 25.505 144.135 ;
        RECT 25.275 143.095 27.750 143.575 ;
        RECT 17.640 142.225 17.910 142.435 ;
        RECT 17.670 142.195 17.900 142.225 ;
        RECT 25.275 142.195 25.505 143.095 ;
        RECT 6.905 137.080 8.650 137.680 ;
        RECT 6.905 135.740 7.135 137.080 ;
        RECT 7.800 137.070 8.650 137.080 ;
        RECT 7.990 137.060 8.650 137.070 ;
        RECT 17.670 137.575 17.900 137.700 ;
        RECT 17.670 137.570 18.400 137.575 ;
        RECT 17.670 137.075 18.435 137.570 ;
        RECT 17.670 136.000 17.900 137.075 ;
        RECT 18.205 137.070 18.435 137.075 ;
        RECT 25.275 137.140 25.505 137.700 ;
        RECT 25.275 136.660 27.750 137.140 ;
        RECT 17.640 135.790 17.910 136.000 ;
        RECT 17.670 135.760 17.900 135.790 ;
        RECT 25.275 135.760 25.505 136.660 ;
        RECT 6.905 130.645 8.650 131.245 ;
        RECT 6.905 129.305 7.135 130.645 ;
        RECT 7.800 130.635 8.650 130.645 ;
        RECT 7.990 130.625 8.650 130.635 ;
        RECT 17.670 131.140 17.900 131.265 ;
        RECT 17.670 131.135 18.400 131.140 ;
        RECT 17.670 130.640 18.435 131.135 ;
        RECT 17.670 129.565 17.900 130.640 ;
        RECT 18.205 130.635 18.435 130.640 ;
        RECT 25.275 130.705 25.505 131.265 ;
        RECT 25.275 130.225 27.750 130.705 ;
        RECT 17.640 129.355 17.910 129.565 ;
        RECT 17.670 129.325 17.900 129.355 ;
        RECT 25.275 129.325 25.505 130.225 ;
        RECT 6.905 124.210 8.650 124.810 ;
        RECT 6.905 122.870 7.135 124.210 ;
        RECT 7.800 124.200 8.650 124.210 ;
        RECT 7.990 124.190 8.650 124.200 ;
        RECT 17.670 124.705 17.900 124.830 ;
        RECT 17.670 124.700 18.400 124.705 ;
        RECT 17.670 124.205 18.435 124.700 ;
        RECT 17.670 123.130 17.900 124.205 ;
        RECT 18.205 124.200 18.435 124.205 ;
        RECT 25.275 124.270 25.505 124.830 ;
        RECT 25.275 123.790 27.750 124.270 ;
        RECT 17.640 122.920 17.910 123.130 ;
        RECT 17.670 122.890 17.900 122.920 ;
        RECT 25.275 122.890 25.505 123.790 ;
        RECT 6.905 117.775 8.650 118.375 ;
        RECT 6.905 116.435 7.135 117.775 ;
        RECT 7.800 117.765 8.650 117.775 ;
        RECT 7.990 117.755 8.650 117.765 ;
        RECT 17.670 118.270 17.900 118.395 ;
        RECT 17.670 118.265 18.400 118.270 ;
        RECT 17.670 117.770 18.435 118.265 ;
        RECT 17.670 116.695 17.900 117.770 ;
        RECT 18.205 117.765 18.435 117.770 ;
        RECT 25.275 117.835 25.505 118.395 ;
        RECT 25.275 117.355 27.750 117.835 ;
        RECT 17.640 116.485 17.910 116.695 ;
        RECT 17.670 116.455 17.900 116.485 ;
        RECT 25.275 116.455 25.505 117.355 ;
        RECT 6.905 111.340 8.650 111.940 ;
        RECT 6.905 110.000 7.135 111.340 ;
        RECT 7.800 111.330 8.650 111.340 ;
        RECT 7.990 111.320 8.650 111.330 ;
        RECT 17.670 111.835 17.900 111.960 ;
        RECT 17.670 111.830 18.400 111.835 ;
        RECT 17.670 111.335 18.435 111.830 ;
        RECT 17.670 110.260 17.900 111.335 ;
        RECT 18.205 111.330 18.435 111.335 ;
        RECT 25.275 111.400 25.505 111.960 ;
        RECT 25.275 110.920 27.750 111.400 ;
        RECT 17.640 110.050 17.910 110.260 ;
        RECT 17.670 110.020 17.900 110.050 ;
        RECT 25.275 110.020 25.505 110.920 ;
        RECT 6.905 104.905 8.650 105.505 ;
        RECT 6.905 103.565 7.135 104.905 ;
        RECT 7.800 104.895 8.650 104.905 ;
        RECT 7.990 104.885 8.650 104.895 ;
        RECT 17.670 105.400 17.900 105.525 ;
        RECT 17.670 105.395 18.400 105.400 ;
        RECT 17.670 104.900 18.435 105.395 ;
        RECT 17.670 103.825 17.900 104.900 ;
        RECT 18.205 104.895 18.435 104.900 ;
        RECT 25.275 104.965 25.505 105.525 ;
        RECT 25.275 104.485 27.750 104.965 ;
        RECT 17.640 103.615 17.910 103.825 ;
        RECT 17.670 103.585 17.900 103.615 ;
        RECT 25.275 103.585 25.505 104.485 ;
        RECT 6.905 98.470 8.650 99.070 ;
        RECT 6.905 97.130 7.135 98.470 ;
        RECT 7.800 98.460 8.650 98.470 ;
        RECT 7.990 98.450 8.650 98.460 ;
        RECT 17.670 98.965 17.900 99.090 ;
        RECT 17.670 98.960 18.400 98.965 ;
        RECT 17.670 98.465 18.435 98.960 ;
        RECT 17.670 97.390 17.900 98.465 ;
        RECT 18.205 98.460 18.435 98.465 ;
        RECT 25.275 98.530 25.505 99.090 ;
        RECT 25.275 98.050 27.750 98.530 ;
        RECT 17.640 97.180 17.910 97.390 ;
        RECT 17.670 97.150 17.900 97.180 ;
        RECT 25.275 97.150 25.505 98.050 ;
        RECT 6.905 92.035 8.650 92.635 ;
        RECT 6.905 90.695 7.135 92.035 ;
        RECT 7.800 92.025 8.650 92.035 ;
        RECT 7.990 92.015 8.650 92.025 ;
        RECT 17.670 92.530 17.900 92.655 ;
        RECT 17.670 92.525 18.400 92.530 ;
        RECT 17.670 92.030 18.435 92.525 ;
        RECT 17.670 90.955 17.900 92.030 ;
        RECT 18.205 92.025 18.435 92.030 ;
        RECT 25.275 92.095 25.505 92.655 ;
        RECT 25.275 91.615 27.750 92.095 ;
        RECT 17.640 90.745 17.910 90.955 ;
        RECT 17.670 90.715 17.900 90.745 ;
        RECT 25.275 90.715 25.505 91.615 ;
        RECT 6.905 85.600 8.650 86.200 ;
        RECT 6.905 84.260 7.135 85.600 ;
        RECT 7.800 85.590 8.650 85.600 ;
        RECT 7.990 85.580 8.650 85.590 ;
        RECT 17.670 86.095 17.900 86.220 ;
        RECT 17.670 86.090 18.400 86.095 ;
        RECT 17.670 85.595 18.435 86.090 ;
        RECT 17.670 84.520 17.900 85.595 ;
        RECT 18.205 85.590 18.435 85.595 ;
        RECT 25.275 85.660 25.505 86.220 ;
        RECT 25.275 85.180 27.750 85.660 ;
        RECT 17.640 84.310 17.910 84.520 ;
        RECT 17.670 84.280 17.900 84.310 ;
        RECT 25.275 84.280 25.505 85.180 ;
        RECT 6.905 79.165 8.650 79.765 ;
        RECT 6.905 77.825 7.135 79.165 ;
        RECT 7.800 79.155 8.650 79.165 ;
        RECT 7.990 79.145 8.650 79.155 ;
        RECT 17.670 79.660 17.900 79.785 ;
        RECT 17.670 79.655 18.400 79.660 ;
        RECT 17.670 79.160 18.435 79.655 ;
        RECT 17.670 78.085 17.900 79.160 ;
        RECT 18.205 79.155 18.435 79.160 ;
        RECT 25.275 79.225 25.505 79.785 ;
        RECT 25.275 78.745 27.750 79.225 ;
        RECT 17.640 77.875 17.910 78.085 ;
        RECT 17.670 77.845 17.900 77.875 ;
        RECT 25.275 77.845 25.505 78.745 ;
        RECT 6.905 72.730 8.650 73.330 ;
        RECT 6.905 71.390 7.135 72.730 ;
        RECT 7.800 72.720 8.650 72.730 ;
        RECT 7.990 72.710 8.650 72.720 ;
        RECT 17.670 73.225 17.900 73.350 ;
        RECT 17.670 73.220 18.400 73.225 ;
        RECT 17.670 72.725 18.435 73.220 ;
        RECT 17.670 71.650 17.900 72.725 ;
        RECT 18.205 72.720 18.435 72.725 ;
        RECT 25.275 72.790 25.505 73.350 ;
        RECT 25.275 72.310 27.750 72.790 ;
        RECT 17.640 71.440 17.910 71.650 ;
        RECT 17.670 71.410 17.900 71.440 ;
        RECT 25.275 71.410 25.505 72.310 ;
        RECT 6.905 66.295 8.650 66.895 ;
        RECT 6.905 64.955 7.135 66.295 ;
        RECT 7.800 66.285 8.650 66.295 ;
        RECT 7.990 66.275 8.650 66.285 ;
        RECT 17.670 66.790 17.900 66.915 ;
        RECT 17.670 66.785 18.400 66.790 ;
        RECT 17.670 66.290 18.435 66.785 ;
        RECT 17.670 65.215 17.900 66.290 ;
        RECT 18.205 66.285 18.435 66.290 ;
        RECT 25.275 66.355 25.505 66.915 ;
        RECT 25.275 65.875 27.750 66.355 ;
        RECT 17.640 65.005 17.910 65.215 ;
        RECT 17.670 64.975 17.900 65.005 ;
        RECT 25.275 64.975 25.505 65.875 ;
        RECT 6.905 59.860 8.650 60.460 ;
        RECT 6.905 58.520 7.135 59.860 ;
        RECT 7.800 59.850 8.650 59.860 ;
        RECT 7.990 59.840 8.650 59.850 ;
        RECT 17.670 60.355 17.900 60.480 ;
        RECT 17.670 60.350 18.400 60.355 ;
        RECT 17.670 59.855 18.435 60.350 ;
        RECT 17.670 58.780 17.900 59.855 ;
        RECT 18.205 59.850 18.435 59.855 ;
        RECT 25.275 59.920 25.505 60.480 ;
        RECT 25.275 59.440 27.750 59.920 ;
        RECT 17.640 58.570 17.910 58.780 ;
        RECT 17.670 58.540 17.900 58.570 ;
        RECT 25.275 58.540 25.505 59.440 ;
        RECT 6.905 53.425 8.650 54.025 ;
        RECT 6.905 52.085 7.135 53.425 ;
        RECT 7.800 53.415 8.650 53.425 ;
        RECT 7.990 53.405 8.650 53.415 ;
        RECT 17.670 53.920 17.900 54.045 ;
        RECT 17.670 53.915 18.400 53.920 ;
        RECT 17.670 53.420 18.435 53.915 ;
        RECT 17.670 52.345 17.900 53.420 ;
        RECT 18.205 53.415 18.435 53.420 ;
        RECT 25.275 53.485 25.505 54.045 ;
        RECT 25.275 53.005 27.750 53.485 ;
        RECT 17.640 52.135 17.910 52.345 ;
        RECT 17.670 52.105 17.900 52.135 ;
        RECT 25.275 52.105 25.505 53.005 ;
        RECT 6.905 46.990 8.650 47.590 ;
        RECT 6.905 45.650 7.135 46.990 ;
        RECT 7.800 46.980 8.650 46.990 ;
        RECT 7.990 46.970 8.650 46.980 ;
        RECT 17.670 47.485 17.900 47.610 ;
        RECT 17.670 47.480 18.400 47.485 ;
        RECT 17.670 46.985 18.435 47.480 ;
        RECT 17.670 45.910 17.900 46.985 ;
        RECT 18.205 46.980 18.435 46.985 ;
        RECT 25.275 47.050 25.505 47.610 ;
        RECT 25.275 46.570 27.750 47.050 ;
        RECT 17.640 45.700 17.910 45.910 ;
        RECT 17.670 45.670 17.900 45.700 ;
        RECT 25.275 45.670 25.505 46.570 ;
        RECT 6.905 40.555 8.650 41.155 ;
        RECT 6.905 39.215 7.135 40.555 ;
        RECT 7.800 40.545 8.650 40.555 ;
        RECT 7.990 40.535 8.650 40.545 ;
        RECT 17.670 41.050 17.900 41.175 ;
        RECT 17.670 41.045 18.400 41.050 ;
        RECT 17.670 40.550 18.435 41.045 ;
        RECT 17.670 39.475 17.900 40.550 ;
        RECT 18.205 40.545 18.435 40.550 ;
        RECT 25.275 40.615 25.505 41.175 ;
        RECT 25.275 40.135 27.750 40.615 ;
        RECT 17.640 39.265 17.910 39.475 ;
        RECT 17.670 39.235 17.900 39.265 ;
        RECT 25.275 39.235 25.505 40.135 ;
        RECT 6.905 34.120 8.650 34.720 ;
        RECT 6.905 32.780 7.135 34.120 ;
        RECT 7.800 34.110 8.650 34.120 ;
        RECT 7.990 34.100 8.650 34.110 ;
        RECT 17.670 34.615 17.900 34.740 ;
        RECT 17.670 34.610 18.400 34.615 ;
        RECT 17.670 34.115 18.435 34.610 ;
        RECT 17.670 33.040 17.900 34.115 ;
        RECT 18.205 34.110 18.435 34.115 ;
        RECT 25.275 34.180 25.505 34.740 ;
        RECT 25.275 33.700 27.750 34.180 ;
        RECT 17.640 32.830 17.910 33.040 ;
        RECT 17.670 32.800 17.900 32.830 ;
        RECT 25.275 32.800 25.505 33.700 ;
        RECT 6.905 27.685 8.650 28.285 ;
        RECT 6.905 26.345 7.135 27.685 ;
        RECT 7.800 27.675 8.650 27.685 ;
        RECT 7.990 27.665 8.650 27.675 ;
        RECT 17.670 28.180 17.900 28.305 ;
        RECT 17.670 28.175 18.400 28.180 ;
        RECT 17.670 27.680 18.435 28.175 ;
        RECT 17.670 26.605 17.900 27.680 ;
        RECT 18.205 27.675 18.435 27.680 ;
        RECT 25.275 27.745 25.505 28.305 ;
        RECT 25.275 27.265 27.750 27.745 ;
        RECT 17.640 26.395 17.910 26.605 ;
        RECT 17.670 26.365 17.900 26.395 ;
        RECT 25.275 26.365 25.505 27.265 ;
        RECT 6.905 21.250 8.650 21.850 ;
        RECT 6.905 19.910 7.135 21.250 ;
        RECT 7.800 21.240 8.650 21.250 ;
        RECT 7.990 21.230 8.650 21.240 ;
        RECT 17.670 21.745 17.900 21.870 ;
        RECT 17.670 21.740 18.400 21.745 ;
        RECT 17.670 21.245 18.435 21.740 ;
        RECT 17.670 20.170 17.900 21.245 ;
        RECT 18.205 21.240 18.435 21.245 ;
        RECT 25.275 21.310 25.505 21.870 ;
        RECT 25.275 20.830 27.750 21.310 ;
        RECT 17.640 19.960 17.910 20.170 ;
        RECT 17.670 19.930 17.900 19.960 ;
        RECT 25.275 19.930 25.505 20.830 ;
        RECT 6.905 14.815 8.650 15.415 ;
        RECT 6.905 13.475 7.135 14.815 ;
        RECT 7.800 14.805 8.650 14.815 ;
        RECT 7.990 14.795 8.650 14.805 ;
        RECT 17.670 15.310 17.900 15.435 ;
        RECT 17.670 15.305 18.400 15.310 ;
        RECT 17.670 14.810 18.435 15.305 ;
        RECT 17.670 13.735 17.900 14.810 ;
        RECT 18.205 14.805 18.435 14.810 ;
        RECT 25.275 14.875 25.505 15.435 ;
        RECT 25.275 14.395 27.750 14.875 ;
        RECT 17.640 13.525 17.910 13.735 ;
        RECT 17.670 13.495 17.900 13.525 ;
        RECT 25.275 13.495 25.505 14.395 ;
        RECT 6.905 8.380 8.650 8.980 ;
        RECT 6.905 7.040 7.135 8.380 ;
        RECT 7.800 8.370 8.650 8.380 ;
        RECT 7.990 8.360 8.650 8.370 ;
        RECT 17.670 8.875 17.900 9.000 ;
        RECT 17.670 8.870 18.400 8.875 ;
        RECT 17.670 8.375 18.435 8.870 ;
        RECT 17.670 7.300 17.900 8.375 ;
        RECT 18.205 8.370 18.435 8.375 ;
        RECT 25.275 8.440 25.505 9.000 ;
        RECT 25.275 7.960 27.750 8.440 ;
        RECT 17.640 7.090 17.910 7.300 ;
        RECT 17.670 7.060 17.900 7.090 ;
        RECT 25.275 7.060 25.505 7.960 ;
        RECT 6.905 1.945 8.650 2.545 ;
        RECT 6.905 0.230 7.135 1.945 ;
        RECT 7.800 1.935 8.650 1.945 ;
        RECT 7.990 1.925 8.650 1.935 ;
        RECT 17.670 2.440 17.900 2.565 ;
        RECT 17.670 2.435 18.400 2.440 ;
        RECT 17.670 1.940 18.435 2.435 ;
        RECT 17.670 0.880 17.900 1.940 ;
        RECT 18.205 1.935 18.435 1.940 ;
        RECT 25.275 2.005 25.505 2.565 ;
        RECT 25.275 1.525 27.750 2.005 ;
        RECT 25.275 0.980 25.505 1.525 ;
        RECT 17.670 0.865 17.925 0.880 ;
        RECT 17.640 0.655 17.925 0.865 ;
        RECT 17.670 0.625 17.925 0.655 ;
        RECT 25.275 0.625 25.525 0.980 ;
        RECT 17.695 0.230 17.925 0.625 ;
        RECT 25.295 0.230 25.525 0.625 ;
        RECT 6.905 0.000 25.525 0.230 ;
      LAYER via ;
        RECT 8.040 201.410 8.600 202.030 ;
        RECT 8.040 194.975 8.600 195.595 ;
        RECT 8.040 188.540 8.600 189.160 ;
        RECT 8.040 182.105 8.600 182.725 ;
        RECT 8.040 175.670 8.600 176.290 ;
        RECT 8.040 169.235 8.600 169.855 ;
        RECT 8.040 162.800 8.600 163.420 ;
        RECT 8.040 156.365 8.600 156.985 ;
        RECT 8.040 149.930 8.600 150.550 ;
        RECT 8.040 143.495 8.600 144.115 ;
        RECT 8.040 137.060 8.600 137.680 ;
        RECT 8.040 130.625 8.600 131.245 ;
        RECT 8.040 124.190 8.600 124.810 ;
        RECT 8.040 117.755 8.600 118.375 ;
        RECT 8.040 111.320 8.600 111.940 ;
        RECT 8.040 104.885 8.600 105.505 ;
        RECT 8.040 98.450 8.600 99.070 ;
        RECT 8.040 92.015 8.600 92.635 ;
        RECT 8.040 85.580 8.600 86.200 ;
        RECT 8.040 79.145 8.600 79.765 ;
        RECT 8.040 72.710 8.600 73.330 ;
        RECT 8.040 66.275 8.600 66.895 ;
        RECT 8.040 59.840 8.600 60.460 ;
        RECT 8.040 53.405 8.600 54.025 ;
        RECT 8.040 46.970 8.600 47.590 ;
        RECT 8.040 40.535 8.600 41.155 ;
        RECT 8.040 34.100 8.600 34.720 ;
        RECT 8.040 27.665 8.600 28.285 ;
        RECT 8.040 21.230 8.600 21.850 ;
        RECT 8.040 14.795 8.600 15.415 ;
        RECT 8.040 8.360 8.600 8.980 ;
        RECT 8.040 1.925 8.600 2.545 ;
      LAYER met2 ;
        RECT 8.050 202.080 8.610 206.475 ;
        RECT 8.040 201.360 8.610 202.080 ;
        RECT 8.050 195.645 8.610 201.360 ;
        RECT 8.040 194.925 8.610 195.645 ;
        RECT 8.050 189.210 8.610 194.925 ;
        RECT 8.040 188.490 8.610 189.210 ;
        RECT 8.050 182.775 8.610 188.490 ;
        RECT 8.040 182.055 8.610 182.775 ;
        RECT 8.050 176.340 8.610 182.055 ;
        RECT 8.040 175.620 8.610 176.340 ;
        RECT 8.050 169.905 8.610 175.620 ;
        RECT 8.040 169.185 8.610 169.905 ;
        RECT 8.050 163.470 8.610 169.185 ;
        RECT 8.040 162.750 8.610 163.470 ;
        RECT 8.050 157.035 8.610 162.750 ;
        RECT 8.040 156.315 8.610 157.035 ;
        RECT 8.050 150.600 8.610 156.315 ;
        RECT 8.040 149.880 8.610 150.600 ;
        RECT 8.050 144.165 8.610 149.880 ;
        RECT 8.040 143.445 8.610 144.165 ;
        RECT 8.050 137.730 8.610 143.445 ;
        RECT 8.040 137.010 8.610 137.730 ;
        RECT 8.050 131.295 8.610 137.010 ;
        RECT 8.040 130.575 8.610 131.295 ;
        RECT 8.050 124.860 8.610 130.575 ;
        RECT 8.040 124.140 8.610 124.860 ;
        RECT 8.050 118.425 8.610 124.140 ;
        RECT 8.040 117.705 8.610 118.425 ;
        RECT 8.050 111.990 8.610 117.705 ;
        RECT 8.040 111.270 8.610 111.990 ;
        RECT 8.050 105.555 8.610 111.270 ;
        RECT 8.040 104.835 8.610 105.555 ;
        RECT 8.050 99.120 8.610 104.835 ;
        RECT 8.040 98.400 8.610 99.120 ;
        RECT 8.050 92.685 8.610 98.400 ;
        RECT 8.040 91.965 8.610 92.685 ;
        RECT 8.050 86.250 8.610 91.965 ;
        RECT 8.040 85.530 8.610 86.250 ;
        RECT 8.050 79.815 8.610 85.530 ;
        RECT 8.040 79.095 8.610 79.815 ;
        RECT 8.050 73.380 8.610 79.095 ;
        RECT 8.040 72.660 8.610 73.380 ;
        RECT 8.050 66.945 8.610 72.660 ;
        RECT 8.040 66.225 8.610 66.945 ;
        RECT 8.050 60.510 8.610 66.225 ;
        RECT 8.040 59.790 8.610 60.510 ;
        RECT 8.050 54.075 8.610 59.790 ;
        RECT 8.040 53.355 8.610 54.075 ;
        RECT 8.050 47.640 8.610 53.355 ;
        RECT 8.040 46.920 8.610 47.640 ;
        RECT 8.050 41.205 8.610 46.920 ;
        RECT 8.040 40.485 8.610 41.205 ;
        RECT 8.050 34.770 8.610 40.485 ;
        RECT 8.040 34.050 8.610 34.770 ;
        RECT 8.050 28.335 8.610 34.050 ;
        RECT 8.040 27.615 8.610 28.335 ;
        RECT 8.050 21.900 8.610 27.615 ;
        RECT 8.040 21.180 8.610 21.900 ;
        RECT 8.050 15.465 8.610 21.180 ;
        RECT 8.040 14.745 8.610 15.465 ;
        RECT 8.050 9.030 8.610 14.745 ;
        RECT 8.040 8.310 8.610 9.030 ;
        RECT 8.050 2.595 8.610 8.310 ;
        RECT 8.040 1.875 8.610 2.595 ;
        RECT 8.050 0.725 8.610 1.875 ;
    END
  END VSS
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT 11.580 205.880 27.950 205.900 ;
        RECT 0.815 204.070 27.950 205.880 ;
        RECT 0.815 202.650 27.940 204.070 ;
        RECT 0.815 202.630 12.415 202.650 ;
        RECT 26.180 202.555 27.940 202.650 ;
        RECT 11.580 199.445 27.950 199.465 ;
        RECT 0.815 197.635 27.950 199.445 ;
        RECT 0.815 196.215 27.940 197.635 ;
        RECT 0.815 196.195 12.415 196.215 ;
        RECT 26.180 196.120 27.940 196.215 ;
        RECT 11.580 193.010 27.950 193.030 ;
        RECT 0.815 191.200 27.950 193.010 ;
        RECT 0.815 189.780 27.940 191.200 ;
        RECT 0.815 189.760 12.415 189.780 ;
        RECT 26.180 189.685 27.940 189.780 ;
        RECT 11.580 186.575 27.950 186.595 ;
        RECT 0.815 184.765 27.950 186.575 ;
        RECT 0.815 183.345 27.940 184.765 ;
        RECT 0.815 183.325 12.415 183.345 ;
        RECT 26.180 183.250 27.940 183.345 ;
        RECT 11.580 180.140 27.950 180.160 ;
        RECT 0.815 178.330 27.950 180.140 ;
        RECT 0.815 176.910 27.940 178.330 ;
        RECT 0.815 176.890 12.415 176.910 ;
        RECT 26.180 176.815 27.940 176.910 ;
        RECT 11.580 173.705 27.950 173.725 ;
        RECT 0.815 171.895 27.950 173.705 ;
        RECT 0.815 170.475 27.940 171.895 ;
        RECT 0.815 170.455 12.415 170.475 ;
        RECT 26.180 170.380 27.940 170.475 ;
        RECT 11.580 167.270 27.950 167.290 ;
        RECT 0.815 165.460 27.950 167.270 ;
        RECT 0.815 164.040 27.940 165.460 ;
        RECT 0.815 164.020 12.415 164.040 ;
        RECT 26.180 163.945 27.940 164.040 ;
        RECT 11.580 160.835 27.950 160.855 ;
        RECT 0.815 159.025 27.950 160.835 ;
        RECT 0.815 157.605 27.940 159.025 ;
        RECT 0.815 157.585 12.415 157.605 ;
        RECT 26.180 157.510 27.940 157.605 ;
        RECT 11.580 154.400 27.950 154.420 ;
        RECT 0.815 152.590 27.950 154.400 ;
        RECT 0.815 151.170 27.940 152.590 ;
        RECT 0.815 151.150 12.415 151.170 ;
        RECT 26.180 151.075 27.940 151.170 ;
        RECT 11.580 147.965 27.950 147.985 ;
        RECT 0.815 146.155 27.950 147.965 ;
        RECT 0.815 144.735 27.940 146.155 ;
        RECT 0.815 144.715 12.415 144.735 ;
        RECT 26.180 144.640 27.940 144.735 ;
        RECT 11.580 141.530 27.950 141.550 ;
        RECT 0.815 139.720 27.950 141.530 ;
        RECT 0.815 138.300 27.940 139.720 ;
        RECT 0.815 138.280 12.415 138.300 ;
        RECT 26.180 138.205 27.940 138.300 ;
        RECT 11.580 135.095 27.950 135.115 ;
        RECT 0.815 133.285 27.950 135.095 ;
        RECT 0.815 131.865 27.940 133.285 ;
        RECT 0.815 131.845 12.415 131.865 ;
        RECT 26.180 131.770 27.940 131.865 ;
        RECT 11.580 128.660 27.950 128.680 ;
        RECT 0.815 126.850 27.950 128.660 ;
        RECT 0.815 125.430 27.940 126.850 ;
        RECT 0.815 125.410 12.415 125.430 ;
        RECT 26.180 125.335 27.940 125.430 ;
        RECT 11.580 122.225 27.950 122.245 ;
        RECT 0.815 120.415 27.950 122.225 ;
        RECT 0.815 118.995 27.940 120.415 ;
        RECT 0.815 118.975 12.415 118.995 ;
        RECT 26.180 118.900 27.940 118.995 ;
        RECT 11.580 115.790 27.950 115.810 ;
        RECT 0.815 113.980 27.950 115.790 ;
        RECT 0.815 112.560 27.940 113.980 ;
        RECT 0.815 112.540 12.415 112.560 ;
        RECT 26.180 112.465 27.940 112.560 ;
        RECT 11.580 109.355 27.950 109.375 ;
        RECT 0.815 107.545 27.950 109.355 ;
        RECT 0.815 106.125 27.940 107.545 ;
        RECT 0.815 106.105 12.415 106.125 ;
        RECT 26.180 106.030 27.940 106.125 ;
        RECT 11.580 102.920 27.950 102.940 ;
        RECT 0.815 101.110 27.950 102.920 ;
        RECT 0.815 99.690 27.940 101.110 ;
        RECT 0.815 99.670 12.415 99.690 ;
        RECT 26.180 99.595 27.940 99.690 ;
        RECT 11.580 96.485 27.950 96.505 ;
        RECT 0.815 94.675 27.950 96.485 ;
        RECT 0.815 93.255 27.940 94.675 ;
        RECT 0.815 93.235 12.415 93.255 ;
        RECT 26.180 93.160 27.940 93.255 ;
        RECT 11.580 90.050 27.950 90.070 ;
        RECT 0.815 88.240 27.950 90.050 ;
        RECT 0.815 86.820 27.940 88.240 ;
        RECT 0.815 86.800 12.415 86.820 ;
        RECT 26.180 86.725 27.940 86.820 ;
        RECT 11.580 83.615 27.950 83.635 ;
        RECT 0.815 81.805 27.950 83.615 ;
        RECT 0.815 80.385 27.940 81.805 ;
        RECT 0.815 80.365 12.415 80.385 ;
        RECT 26.180 80.290 27.940 80.385 ;
        RECT 11.580 77.180 27.950 77.200 ;
        RECT 0.815 75.370 27.950 77.180 ;
        RECT 0.815 73.950 27.940 75.370 ;
        RECT 0.815 73.930 12.415 73.950 ;
        RECT 26.180 73.855 27.940 73.950 ;
        RECT 11.580 70.745 27.950 70.765 ;
        RECT 0.815 68.935 27.950 70.745 ;
        RECT 0.815 67.515 27.940 68.935 ;
        RECT 0.815 67.495 12.415 67.515 ;
        RECT 26.180 67.420 27.940 67.515 ;
        RECT 11.580 64.310 27.950 64.330 ;
        RECT 0.815 62.500 27.950 64.310 ;
        RECT 0.815 61.080 27.940 62.500 ;
        RECT 0.815 61.060 12.415 61.080 ;
        RECT 26.180 60.985 27.940 61.080 ;
        RECT 11.580 57.875 27.950 57.895 ;
        RECT 0.815 56.065 27.950 57.875 ;
        RECT 0.815 54.645 27.940 56.065 ;
        RECT 0.815 54.625 12.415 54.645 ;
        RECT 26.180 54.550 27.940 54.645 ;
        RECT 11.580 51.440 27.950 51.460 ;
        RECT 0.815 49.630 27.950 51.440 ;
        RECT 0.815 48.210 27.940 49.630 ;
        RECT 0.815 48.190 12.415 48.210 ;
        RECT 26.180 48.115 27.940 48.210 ;
        RECT 11.580 45.005 27.950 45.025 ;
        RECT 0.815 43.195 27.950 45.005 ;
        RECT 0.815 41.775 27.940 43.195 ;
        RECT 0.815 41.755 12.415 41.775 ;
        RECT 26.180 41.680 27.940 41.775 ;
        RECT 11.580 38.570 27.950 38.590 ;
        RECT 0.815 36.760 27.950 38.570 ;
        RECT 0.815 35.340 27.940 36.760 ;
        RECT 0.815 35.320 12.415 35.340 ;
        RECT 26.180 35.245 27.940 35.340 ;
        RECT 11.580 32.135 27.950 32.155 ;
        RECT 0.815 30.325 27.950 32.135 ;
        RECT 0.815 28.905 27.940 30.325 ;
        RECT 0.815 28.885 12.415 28.905 ;
        RECT 26.180 28.810 27.940 28.905 ;
        RECT 11.580 25.700 27.950 25.720 ;
        RECT 0.815 23.890 27.950 25.700 ;
        RECT 0.815 22.470 27.940 23.890 ;
        RECT 0.815 22.450 12.415 22.470 ;
        RECT 26.180 22.375 27.940 22.470 ;
        RECT 11.580 19.265 27.950 19.285 ;
        RECT 0.815 17.455 27.950 19.265 ;
        RECT 0.815 16.035 27.940 17.455 ;
        RECT 0.815 16.015 12.415 16.035 ;
        RECT 26.180 15.940 27.940 16.035 ;
        RECT 11.580 12.830 27.950 12.850 ;
        RECT 0.815 11.020 27.950 12.830 ;
        RECT 0.815 9.600 27.940 11.020 ;
        RECT 0.815 9.580 12.415 9.600 ;
        RECT 26.180 9.505 27.940 9.600 ;
        RECT 11.580 6.395 27.950 6.415 ;
        RECT 0.815 4.585 27.950 6.395 ;
        RECT 0.815 3.165 27.940 4.585 ;
        RECT 0.815 3.145 12.415 3.165 ;
        RECT 26.180 3.070 27.940 3.165 ;
      LAYER li1 ;
        RECT 0.995 205.530 7.105 205.700 ;
        RECT 0.995 202.980 1.165 205.530 ;
        RECT 6.935 202.980 7.105 205.530 ;
        RECT 0.995 202.810 7.105 202.980 ;
        RECT 11.760 205.550 17.870 205.720 ;
        RECT 11.760 203.000 11.930 205.550 ;
        RECT 17.700 203.000 17.870 205.550 ;
        RECT 11.760 202.830 17.870 203.000 ;
        RECT 19.365 205.550 25.475 205.720 ;
        RECT 19.365 203.000 19.535 205.550 ;
        RECT 25.305 203.000 25.475 205.550 ;
        RECT 26.370 203.885 27.750 204.055 ;
        RECT 19.365 202.830 25.475 203.000 ;
        RECT 27.200 202.745 27.410 203.885 ;
        RECT 0.995 199.095 7.105 199.265 ;
        RECT 0.995 196.545 1.165 199.095 ;
        RECT 6.935 196.545 7.105 199.095 ;
        RECT 0.995 196.375 7.105 196.545 ;
        RECT 11.760 199.115 17.870 199.285 ;
        RECT 11.760 196.565 11.930 199.115 ;
        RECT 17.700 196.565 17.870 199.115 ;
        RECT 11.760 196.395 17.870 196.565 ;
        RECT 19.365 199.115 25.475 199.285 ;
        RECT 19.365 196.565 19.535 199.115 ;
        RECT 25.305 196.565 25.475 199.115 ;
        RECT 26.370 197.450 27.750 197.620 ;
        RECT 19.365 196.395 25.475 196.565 ;
        RECT 27.200 196.310 27.410 197.450 ;
        RECT 0.995 192.660 7.105 192.830 ;
        RECT 0.995 190.110 1.165 192.660 ;
        RECT 6.935 190.110 7.105 192.660 ;
        RECT 0.995 189.940 7.105 190.110 ;
        RECT 11.760 192.680 17.870 192.850 ;
        RECT 11.760 190.130 11.930 192.680 ;
        RECT 17.700 190.130 17.870 192.680 ;
        RECT 11.760 189.960 17.870 190.130 ;
        RECT 19.365 192.680 25.475 192.850 ;
        RECT 19.365 190.130 19.535 192.680 ;
        RECT 25.305 190.130 25.475 192.680 ;
        RECT 26.370 191.015 27.750 191.185 ;
        RECT 19.365 189.960 25.475 190.130 ;
        RECT 27.200 189.875 27.410 191.015 ;
        RECT 0.995 186.225 7.105 186.395 ;
        RECT 0.995 183.675 1.165 186.225 ;
        RECT 6.935 183.675 7.105 186.225 ;
        RECT 0.995 183.505 7.105 183.675 ;
        RECT 11.760 186.245 17.870 186.415 ;
        RECT 11.760 183.695 11.930 186.245 ;
        RECT 17.700 183.695 17.870 186.245 ;
        RECT 11.760 183.525 17.870 183.695 ;
        RECT 19.365 186.245 25.475 186.415 ;
        RECT 19.365 183.695 19.535 186.245 ;
        RECT 25.305 183.695 25.475 186.245 ;
        RECT 26.370 184.580 27.750 184.750 ;
        RECT 19.365 183.525 25.475 183.695 ;
        RECT 27.200 183.440 27.410 184.580 ;
        RECT 0.995 179.790 7.105 179.960 ;
        RECT 0.995 177.240 1.165 179.790 ;
        RECT 6.935 177.240 7.105 179.790 ;
        RECT 0.995 177.070 7.105 177.240 ;
        RECT 11.760 179.810 17.870 179.980 ;
        RECT 11.760 177.260 11.930 179.810 ;
        RECT 17.700 177.260 17.870 179.810 ;
        RECT 11.760 177.090 17.870 177.260 ;
        RECT 19.365 179.810 25.475 179.980 ;
        RECT 19.365 177.260 19.535 179.810 ;
        RECT 25.305 177.260 25.475 179.810 ;
        RECT 26.370 178.145 27.750 178.315 ;
        RECT 19.365 177.090 25.475 177.260 ;
        RECT 27.200 177.005 27.410 178.145 ;
        RECT 0.995 173.355 7.105 173.525 ;
        RECT 0.995 170.805 1.165 173.355 ;
        RECT 6.935 170.805 7.105 173.355 ;
        RECT 0.995 170.635 7.105 170.805 ;
        RECT 11.760 173.375 17.870 173.545 ;
        RECT 11.760 170.825 11.930 173.375 ;
        RECT 17.700 170.825 17.870 173.375 ;
        RECT 11.760 170.655 17.870 170.825 ;
        RECT 19.365 173.375 25.475 173.545 ;
        RECT 19.365 170.825 19.535 173.375 ;
        RECT 25.305 170.825 25.475 173.375 ;
        RECT 26.370 171.710 27.750 171.880 ;
        RECT 19.365 170.655 25.475 170.825 ;
        RECT 27.200 170.570 27.410 171.710 ;
        RECT 0.995 166.920 7.105 167.090 ;
        RECT 0.995 164.370 1.165 166.920 ;
        RECT 6.935 164.370 7.105 166.920 ;
        RECT 0.995 164.200 7.105 164.370 ;
        RECT 11.760 166.940 17.870 167.110 ;
        RECT 11.760 164.390 11.930 166.940 ;
        RECT 17.700 164.390 17.870 166.940 ;
        RECT 11.760 164.220 17.870 164.390 ;
        RECT 19.365 166.940 25.475 167.110 ;
        RECT 19.365 164.390 19.535 166.940 ;
        RECT 25.305 164.390 25.475 166.940 ;
        RECT 26.370 165.275 27.750 165.445 ;
        RECT 19.365 164.220 25.475 164.390 ;
        RECT 27.200 164.135 27.410 165.275 ;
        RECT 0.995 160.485 7.105 160.655 ;
        RECT 0.995 157.935 1.165 160.485 ;
        RECT 6.935 157.935 7.105 160.485 ;
        RECT 0.995 157.765 7.105 157.935 ;
        RECT 11.760 160.505 17.870 160.675 ;
        RECT 11.760 157.955 11.930 160.505 ;
        RECT 17.700 157.955 17.870 160.505 ;
        RECT 11.760 157.785 17.870 157.955 ;
        RECT 19.365 160.505 25.475 160.675 ;
        RECT 19.365 157.955 19.535 160.505 ;
        RECT 25.305 157.955 25.475 160.505 ;
        RECT 26.370 158.840 27.750 159.010 ;
        RECT 19.365 157.785 25.475 157.955 ;
        RECT 27.200 157.700 27.410 158.840 ;
        RECT 0.995 154.050 7.105 154.220 ;
        RECT 0.995 151.500 1.165 154.050 ;
        RECT 6.935 151.500 7.105 154.050 ;
        RECT 0.995 151.330 7.105 151.500 ;
        RECT 11.760 154.070 17.870 154.240 ;
        RECT 11.760 151.520 11.930 154.070 ;
        RECT 17.700 151.520 17.870 154.070 ;
        RECT 11.760 151.350 17.870 151.520 ;
        RECT 19.365 154.070 25.475 154.240 ;
        RECT 19.365 151.520 19.535 154.070 ;
        RECT 25.305 151.520 25.475 154.070 ;
        RECT 26.370 152.405 27.750 152.575 ;
        RECT 19.365 151.350 25.475 151.520 ;
        RECT 27.200 151.265 27.410 152.405 ;
        RECT 0.995 147.615 7.105 147.785 ;
        RECT 0.995 145.065 1.165 147.615 ;
        RECT 6.935 145.065 7.105 147.615 ;
        RECT 0.995 144.895 7.105 145.065 ;
        RECT 11.760 147.635 17.870 147.805 ;
        RECT 11.760 145.085 11.930 147.635 ;
        RECT 17.700 145.085 17.870 147.635 ;
        RECT 11.760 144.915 17.870 145.085 ;
        RECT 19.365 147.635 25.475 147.805 ;
        RECT 19.365 145.085 19.535 147.635 ;
        RECT 25.305 145.085 25.475 147.635 ;
        RECT 26.370 145.970 27.750 146.140 ;
        RECT 19.365 144.915 25.475 145.085 ;
        RECT 27.200 144.830 27.410 145.970 ;
        RECT 0.995 141.180 7.105 141.350 ;
        RECT 0.995 138.630 1.165 141.180 ;
        RECT 6.935 138.630 7.105 141.180 ;
        RECT 0.995 138.460 7.105 138.630 ;
        RECT 11.760 141.200 17.870 141.370 ;
        RECT 11.760 138.650 11.930 141.200 ;
        RECT 17.700 138.650 17.870 141.200 ;
        RECT 11.760 138.480 17.870 138.650 ;
        RECT 19.365 141.200 25.475 141.370 ;
        RECT 19.365 138.650 19.535 141.200 ;
        RECT 25.305 138.650 25.475 141.200 ;
        RECT 26.370 139.535 27.750 139.705 ;
        RECT 19.365 138.480 25.475 138.650 ;
        RECT 27.200 138.395 27.410 139.535 ;
        RECT 0.995 134.745 7.105 134.915 ;
        RECT 0.995 132.195 1.165 134.745 ;
        RECT 6.935 132.195 7.105 134.745 ;
        RECT 0.995 132.025 7.105 132.195 ;
        RECT 11.760 134.765 17.870 134.935 ;
        RECT 11.760 132.215 11.930 134.765 ;
        RECT 17.700 132.215 17.870 134.765 ;
        RECT 11.760 132.045 17.870 132.215 ;
        RECT 19.365 134.765 25.475 134.935 ;
        RECT 19.365 132.215 19.535 134.765 ;
        RECT 25.305 132.215 25.475 134.765 ;
        RECT 26.370 133.100 27.750 133.270 ;
        RECT 19.365 132.045 25.475 132.215 ;
        RECT 27.200 131.960 27.410 133.100 ;
        RECT 0.995 128.310 7.105 128.480 ;
        RECT 0.995 125.760 1.165 128.310 ;
        RECT 6.935 125.760 7.105 128.310 ;
        RECT 0.995 125.590 7.105 125.760 ;
        RECT 11.760 128.330 17.870 128.500 ;
        RECT 11.760 125.780 11.930 128.330 ;
        RECT 17.700 125.780 17.870 128.330 ;
        RECT 11.760 125.610 17.870 125.780 ;
        RECT 19.365 128.330 25.475 128.500 ;
        RECT 19.365 125.780 19.535 128.330 ;
        RECT 25.305 125.780 25.475 128.330 ;
        RECT 26.370 126.665 27.750 126.835 ;
        RECT 19.365 125.610 25.475 125.780 ;
        RECT 27.200 125.525 27.410 126.665 ;
        RECT 0.995 121.875 7.105 122.045 ;
        RECT 0.995 119.325 1.165 121.875 ;
        RECT 6.935 119.325 7.105 121.875 ;
        RECT 0.995 119.155 7.105 119.325 ;
        RECT 11.760 121.895 17.870 122.065 ;
        RECT 11.760 119.345 11.930 121.895 ;
        RECT 17.700 119.345 17.870 121.895 ;
        RECT 11.760 119.175 17.870 119.345 ;
        RECT 19.365 121.895 25.475 122.065 ;
        RECT 19.365 119.345 19.535 121.895 ;
        RECT 25.305 119.345 25.475 121.895 ;
        RECT 26.370 120.230 27.750 120.400 ;
        RECT 19.365 119.175 25.475 119.345 ;
        RECT 27.200 119.090 27.410 120.230 ;
        RECT 0.995 115.440 7.105 115.610 ;
        RECT 0.995 112.890 1.165 115.440 ;
        RECT 6.935 112.890 7.105 115.440 ;
        RECT 0.995 112.720 7.105 112.890 ;
        RECT 11.760 115.460 17.870 115.630 ;
        RECT 11.760 112.910 11.930 115.460 ;
        RECT 17.700 112.910 17.870 115.460 ;
        RECT 11.760 112.740 17.870 112.910 ;
        RECT 19.365 115.460 25.475 115.630 ;
        RECT 19.365 112.910 19.535 115.460 ;
        RECT 25.305 112.910 25.475 115.460 ;
        RECT 26.370 113.795 27.750 113.965 ;
        RECT 19.365 112.740 25.475 112.910 ;
        RECT 27.200 112.655 27.410 113.795 ;
        RECT 0.995 109.005 7.105 109.175 ;
        RECT 0.995 106.455 1.165 109.005 ;
        RECT 6.935 106.455 7.105 109.005 ;
        RECT 0.995 106.285 7.105 106.455 ;
        RECT 11.760 109.025 17.870 109.195 ;
        RECT 11.760 106.475 11.930 109.025 ;
        RECT 17.700 106.475 17.870 109.025 ;
        RECT 11.760 106.305 17.870 106.475 ;
        RECT 19.365 109.025 25.475 109.195 ;
        RECT 19.365 106.475 19.535 109.025 ;
        RECT 25.305 106.475 25.475 109.025 ;
        RECT 26.370 107.360 27.750 107.530 ;
        RECT 19.365 106.305 25.475 106.475 ;
        RECT 27.200 106.220 27.410 107.360 ;
        RECT 0.995 102.570 7.105 102.740 ;
        RECT 0.995 100.020 1.165 102.570 ;
        RECT 6.935 100.020 7.105 102.570 ;
        RECT 0.995 99.850 7.105 100.020 ;
        RECT 11.760 102.590 17.870 102.760 ;
        RECT 11.760 100.040 11.930 102.590 ;
        RECT 17.700 100.040 17.870 102.590 ;
        RECT 11.760 99.870 17.870 100.040 ;
        RECT 19.365 102.590 25.475 102.760 ;
        RECT 19.365 100.040 19.535 102.590 ;
        RECT 25.305 100.040 25.475 102.590 ;
        RECT 26.370 100.925 27.750 101.095 ;
        RECT 19.365 99.870 25.475 100.040 ;
        RECT 27.200 99.785 27.410 100.925 ;
        RECT 0.995 96.135 7.105 96.305 ;
        RECT 0.995 93.585 1.165 96.135 ;
        RECT 6.935 93.585 7.105 96.135 ;
        RECT 0.995 93.415 7.105 93.585 ;
        RECT 11.760 96.155 17.870 96.325 ;
        RECT 11.760 93.605 11.930 96.155 ;
        RECT 17.700 93.605 17.870 96.155 ;
        RECT 11.760 93.435 17.870 93.605 ;
        RECT 19.365 96.155 25.475 96.325 ;
        RECT 19.365 93.605 19.535 96.155 ;
        RECT 25.305 93.605 25.475 96.155 ;
        RECT 26.370 94.490 27.750 94.660 ;
        RECT 19.365 93.435 25.475 93.605 ;
        RECT 27.200 93.350 27.410 94.490 ;
        RECT 0.995 89.700 7.105 89.870 ;
        RECT 0.995 87.150 1.165 89.700 ;
        RECT 6.935 87.150 7.105 89.700 ;
        RECT 0.995 86.980 7.105 87.150 ;
        RECT 11.760 89.720 17.870 89.890 ;
        RECT 11.760 87.170 11.930 89.720 ;
        RECT 17.700 87.170 17.870 89.720 ;
        RECT 11.760 87.000 17.870 87.170 ;
        RECT 19.365 89.720 25.475 89.890 ;
        RECT 19.365 87.170 19.535 89.720 ;
        RECT 25.305 87.170 25.475 89.720 ;
        RECT 26.370 88.055 27.750 88.225 ;
        RECT 19.365 87.000 25.475 87.170 ;
        RECT 27.200 86.915 27.410 88.055 ;
        RECT 0.995 83.265 7.105 83.435 ;
        RECT 0.995 80.715 1.165 83.265 ;
        RECT 6.935 80.715 7.105 83.265 ;
        RECT 0.995 80.545 7.105 80.715 ;
        RECT 11.760 83.285 17.870 83.455 ;
        RECT 11.760 80.735 11.930 83.285 ;
        RECT 17.700 80.735 17.870 83.285 ;
        RECT 11.760 80.565 17.870 80.735 ;
        RECT 19.365 83.285 25.475 83.455 ;
        RECT 19.365 80.735 19.535 83.285 ;
        RECT 25.305 80.735 25.475 83.285 ;
        RECT 26.370 81.620 27.750 81.790 ;
        RECT 19.365 80.565 25.475 80.735 ;
        RECT 27.200 80.480 27.410 81.620 ;
        RECT 0.995 76.830 7.105 77.000 ;
        RECT 0.995 74.280 1.165 76.830 ;
        RECT 6.935 74.280 7.105 76.830 ;
        RECT 0.995 74.110 7.105 74.280 ;
        RECT 11.760 76.850 17.870 77.020 ;
        RECT 11.760 74.300 11.930 76.850 ;
        RECT 17.700 74.300 17.870 76.850 ;
        RECT 11.760 74.130 17.870 74.300 ;
        RECT 19.365 76.850 25.475 77.020 ;
        RECT 19.365 74.300 19.535 76.850 ;
        RECT 25.305 74.300 25.475 76.850 ;
        RECT 26.370 75.185 27.750 75.355 ;
        RECT 19.365 74.130 25.475 74.300 ;
        RECT 27.200 74.045 27.410 75.185 ;
        RECT 0.995 70.395 7.105 70.565 ;
        RECT 0.995 67.845 1.165 70.395 ;
        RECT 6.935 67.845 7.105 70.395 ;
        RECT 0.995 67.675 7.105 67.845 ;
        RECT 11.760 70.415 17.870 70.585 ;
        RECT 11.760 67.865 11.930 70.415 ;
        RECT 17.700 67.865 17.870 70.415 ;
        RECT 11.760 67.695 17.870 67.865 ;
        RECT 19.365 70.415 25.475 70.585 ;
        RECT 19.365 67.865 19.535 70.415 ;
        RECT 25.305 67.865 25.475 70.415 ;
        RECT 26.370 68.750 27.750 68.920 ;
        RECT 19.365 67.695 25.475 67.865 ;
        RECT 27.200 67.610 27.410 68.750 ;
        RECT 0.995 63.960 7.105 64.130 ;
        RECT 0.995 61.410 1.165 63.960 ;
        RECT 6.935 61.410 7.105 63.960 ;
        RECT 0.995 61.240 7.105 61.410 ;
        RECT 11.760 63.980 17.870 64.150 ;
        RECT 11.760 61.430 11.930 63.980 ;
        RECT 17.700 61.430 17.870 63.980 ;
        RECT 11.760 61.260 17.870 61.430 ;
        RECT 19.365 63.980 25.475 64.150 ;
        RECT 19.365 61.430 19.535 63.980 ;
        RECT 25.305 61.430 25.475 63.980 ;
        RECT 26.370 62.315 27.750 62.485 ;
        RECT 19.365 61.260 25.475 61.430 ;
        RECT 27.200 61.175 27.410 62.315 ;
        RECT 0.995 57.525 7.105 57.695 ;
        RECT 0.995 54.975 1.165 57.525 ;
        RECT 6.935 54.975 7.105 57.525 ;
        RECT 0.995 54.805 7.105 54.975 ;
        RECT 11.760 57.545 17.870 57.715 ;
        RECT 11.760 54.995 11.930 57.545 ;
        RECT 17.700 54.995 17.870 57.545 ;
        RECT 11.760 54.825 17.870 54.995 ;
        RECT 19.365 57.545 25.475 57.715 ;
        RECT 19.365 54.995 19.535 57.545 ;
        RECT 25.305 54.995 25.475 57.545 ;
        RECT 26.370 55.880 27.750 56.050 ;
        RECT 19.365 54.825 25.475 54.995 ;
        RECT 27.200 54.740 27.410 55.880 ;
        RECT 0.995 51.090 7.105 51.260 ;
        RECT 0.995 48.540 1.165 51.090 ;
        RECT 6.935 48.540 7.105 51.090 ;
        RECT 0.995 48.370 7.105 48.540 ;
        RECT 11.760 51.110 17.870 51.280 ;
        RECT 11.760 48.560 11.930 51.110 ;
        RECT 17.700 48.560 17.870 51.110 ;
        RECT 11.760 48.390 17.870 48.560 ;
        RECT 19.365 51.110 25.475 51.280 ;
        RECT 19.365 48.560 19.535 51.110 ;
        RECT 25.305 48.560 25.475 51.110 ;
        RECT 26.370 49.445 27.750 49.615 ;
        RECT 19.365 48.390 25.475 48.560 ;
        RECT 27.200 48.305 27.410 49.445 ;
        RECT 0.995 44.655 7.105 44.825 ;
        RECT 0.995 42.105 1.165 44.655 ;
        RECT 6.935 42.105 7.105 44.655 ;
        RECT 0.995 41.935 7.105 42.105 ;
        RECT 11.760 44.675 17.870 44.845 ;
        RECT 11.760 42.125 11.930 44.675 ;
        RECT 17.700 42.125 17.870 44.675 ;
        RECT 11.760 41.955 17.870 42.125 ;
        RECT 19.365 44.675 25.475 44.845 ;
        RECT 19.365 42.125 19.535 44.675 ;
        RECT 25.305 42.125 25.475 44.675 ;
        RECT 26.370 43.010 27.750 43.180 ;
        RECT 19.365 41.955 25.475 42.125 ;
        RECT 27.200 41.870 27.410 43.010 ;
        RECT 0.995 38.220 7.105 38.390 ;
        RECT 0.995 35.670 1.165 38.220 ;
        RECT 6.935 35.670 7.105 38.220 ;
        RECT 0.995 35.500 7.105 35.670 ;
        RECT 11.760 38.240 17.870 38.410 ;
        RECT 11.760 35.690 11.930 38.240 ;
        RECT 17.700 35.690 17.870 38.240 ;
        RECT 11.760 35.520 17.870 35.690 ;
        RECT 19.365 38.240 25.475 38.410 ;
        RECT 19.365 35.690 19.535 38.240 ;
        RECT 25.305 35.690 25.475 38.240 ;
        RECT 26.370 36.575 27.750 36.745 ;
        RECT 19.365 35.520 25.475 35.690 ;
        RECT 27.200 35.435 27.410 36.575 ;
        RECT 0.995 31.785 7.105 31.955 ;
        RECT 0.995 29.235 1.165 31.785 ;
        RECT 6.935 29.235 7.105 31.785 ;
        RECT 0.995 29.065 7.105 29.235 ;
        RECT 11.760 31.805 17.870 31.975 ;
        RECT 11.760 29.255 11.930 31.805 ;
        RECT 17.700 29.255 17.870 31.805 ;
        RECT 11.760 29.085 17.870 29.255 ;
        RECT 19.365 31.805 25.475 31.975 ;
        RECT 19.365 29.255 19.535 31.805 ;
        RECT 25.305 29.255 25.475 31.805 ;
        RECT 26.370 30.140 27.750 30.310 ;
        RECT 19.365 29.085 25.475 29.255 ;
        RECT 27.200 29.000 27.410 30.140 ;
        RECT 0.995 25.350 7.105 25.520 ;
        RECT 0.995 22.800 1.165 25.350 ;
        RECT 6.935 22.800 7.105 25.350 ;
        RECT 0.995 22.630 7.105 22.800 ;
        RECT 11.760 25.370 17.870 25.540 ;
        RECT 11.760 22.820 11.930 25.370 ;
        RECT 17.700 22.820 17.870 25.370 ;
        RECT 11.760 22.650 17.870 22.820 ;
        RECT 19.365 25.370 25.475 25.540 ;
        RECT 19.365 22.820 19.535 25.370 ;
        RECT 25.305 22.820 25.475 25.370 ;
        RECT 26.370 23.705 27.750 23.875 ;
        RECT 19.365 22.650 25.475 22.820 ;
        RECT 27.200 22.565 27.410 23.705 ;
        RECT 0.995 18.915 7.105 19.085 ;
        RECT 0.995 16.365 1.165 18.915 ;
        RECT 6.935 16.365 7.105 18.915 ;
        RECT 0.995 16.195 7.105 16.365 ;
        RECT 11.760 18.935 17.870 19.105 ;
        RECT 11.760 16.385 11.930 18.935 ;
        RECT 17.700 16.385 17.870 18.935 ;
        RECT 11.760 16.215 17.870 16.385 ;
        RECT 19.365 18.935 25.475 19.105 ;
        RECT 19.365 16.385 19.535 18.935 ;
        RECT 25.305 16.385 25.475 18.935 ;
        RECT 26.370 17.270 27.750 17.440 ;
        RECT 19.365 16.215 25.475 16.385 ;
        RECT 27.200 16.130 27.410 17.270 ;
        RECT 0.995 12.480 7.105 12.650 ;
        RECT 0.995 9.930 1.165 12.480 ;
        RECT 6.935 9.930 7.105 12.480 ;
        RECT 0.995 9.760 7.105 9.930 ;
        RECT 11.760 12.500 17.870 12.670 ;
        RECT 11.760 9.950 11.930 12.500 ;
        RECT 17.700 9.950 17.870 12.500 ;
        RECT 11.760 9.780 17.870 9.950 ;
        RECT 19.365 12.500 25.475 12.670 ;
        RECT 19.365 9.950 19.535 12.500 ;
        RECT 25.305 9.950 25.475 12.500 ;
        RECT 26.370 10.835 27.750 11.005 ;
        RECT 19.365 9.780 25.475 9.950 ;
        RECT 27.200 9.695 27.410 10.835 ;
        RECT 0.995 6.045 7.105 6.215 ;
        RECT 0.995 3.495 1.165 6.045 ;
        RECT 6.935 3.495 7.105 6.045 ;
        RECT 0.995 3.325 7.105 3.495 ;
        RECT 11.760 6.065 17.870 6.235 ;
        RECT 11.760 3.515 11.930 6.065 ;
        RECT 17.700 3.515 17.870 6.065 ;
        RECT 11.760 3.345 17.870 3.515 ;
        RECT 19.365 6.065 25.475 6.235 ;
        RECT 19.365 3.515 19.535 6.065 ;
        RECT 25.305 3.515 25.475 6.065 ;
        RECT 26.370 4.400 27.750 4.570 ;
        RECT 19.365 3.345 25.475 3.515 ;
        RECT 27.200 3.260 27.410 4.400 ;
      LAYER mcon ;
        RECT 6.935 204.890 7.105 205.060 ;
        RECT 6.935 204.530 7.105 204.700 ;
        RECT 6.935 204.170 7.105 204.340 ;
        RECT 6.935 203.810 7.105 203.980 ;
        RECT 6.935 203.450 7.105 203.620 ;
        RECT 17.700 204.910 17.870 205.080 ;
        RECT 17.700 204.550 17.870 204.720 ;
        RECT 17.700 204.190 17.870 204.360 ;
        RECT 17.700 203.830 17.870 204.000 ;
        RECT 17.700 203.470 17.870 203.640 ;
        RECT 25.305 204.910 25.475 205.080 ;
        RECT 25.305 204.550 25.475 204.720 ;
        RECT 25.305 204.190 25.475 204.360 ;
        RECT 25.305 203.830 25.475 204.000 ;
        RECT 26.515 203.885 26.685 204.055 ;
        RECT 26.975 203.885 27.145 204.055 ;
        RECT 27.435 203.885 27.605 204.055 ;
        RECT 25.305 203.470 25.475 203.640 ;
        RECT 6.935 198.455 7.105 198.625 ;
        RECT 6.935 198.095 7.105 198.265 ;
        RECT 6.935 197.735 7.105 197.905 ;
        RECT 6.935 197.375 7.105 197.545 ;
        RECT 6.935 197.015 7.105 197.185 ;
        RECT 17.700 198.475 17.870 198.645 ;
        RECT 17.700 198.115 17.870 198.285 ;
        RECT 17.700 197.755 17.870 197.925 ;
        RECT 17.700 197.395 17.870 197.565 ;
        RECT 17.700 197.035 17.870 197.205 ;
        RECT 25.305 198.475 25.475 198.645 ;
        RECT 25.305 198.115 25.475 198.285 ;
        RECT 25.305 197.755 25.475 197.925 ;
        RECT 25.305 197.395 25.475 197.565 ;
        RECT 26.515 197.450 26.685 197.620 ;
        RECT 26.975 197.450 27.145 197.620 ;
        RECT 27.435 197.450 27.605 197.620 ;
        RECT 25.305 197.035 25.475 197.205 ;
        RECT 6.935 192.020 7.105 192.190 ;
        RECT 6.935 191.660 7.105 191.830 ;
        RECT 6.935 191.300 7.105 191.470 ;
        RECT 6.935 190.940 7.105 191.110 ;
        RECT 6.935 190.580 7.105 190.750 ;
        RECT 17.700 192.040 17.870 192.210 ;
        RECT 17.700 191.680 17.870 191.850 ;
        RECT 17.700 191.320 17.870 191.490 ;
        RECT 17.700 190.960 17.870 191.130 ;
        RECT 17.700 190.600 17.870 190.770 ;
        RECT 25.305 192.040 25.475 192.210 ;
        RECT 25.305 191.680 25.475 191.850 ;
        RECT 25.305 191.320 25.475 191.490 ;
        RECT 25.305 190.960 25.475 191.130 ;
        RECT 26.515 191.015 26.685 191.185 ;
        RECT 26.975 191.015 27.145 191.185 ;
        RECT 27.435 191.015 27.605 191.185 ;
        RECT 25.305 190.600 25.475 190.770 ;
        RECT 6.935 185.585 7.105 185.755 ;
        RECT 6.935 185.225 7.105 185.395 ;
        RECT 6.935 184.865 7.105 185.035 ;
        RECT 6.935 184.505 7.105 184.675 ;
        RECT 6.935 184.145 7.105 184.315 ;
        RECT 17.700 185.605 17.870 185.775 ;
        RECT 17.700 185.245 17.870 185.415 ;
        RECT 17.700 184.885 17.870 185.055 ;
        RECT 17.700 184.525 17.870 184.695 ;
        RECT 17.700 184.165 17.870 184.335 ;
        RECT 25.305 185.605 25.475 185.775 ;
        RECT 25.305 185.245 25.475 185.415 ;
        RECT 25.305 184.885 25.475 185.055 ;
        RECT 25.305 184.525 25.475 184.695 ;
        RECT 26.515 184.580 26.685 184.750 ;
        RECT 26.975 184.580 27.145 184.750 ;
        RECT 27.435 184.580 27.605 184.750 ;
        RECT 25.305 184.165 25.475 184.335 ;
        RECT 6.935 179.150 7.105 179.320 ;
        RECT 6.935 178.790 7.105 178.960 ;
        RECT 6.935 178.430 7.105 178.600 ;
        RECT 6.935 178.070 7.105 178.240 ;
        RECT 6.935 177.710 7.105 177.880 ;
        RECT 17.700 179.170 17.870 179.340 ;
        RECT 17.700 178.810 17.870 178.980 ;
        RECT 17.700 178.450 17.870 178.620 ;
        RECT 17.700 178.090 17.870 178.260 ;
        RECT 17.700 177.730 17.870 177.900 ;
        RECT 25.305 179.170 25.475 179.340 ;
        RECT 25.305 178.810 25.475 178.980 ;
        RECT 25.305 178.450 25.475 178.620 ;
        RECT 25.305 178.090 25.475 178.260 ;
        RECT 26.515 178.145 26.685 178.315 ;
        RECT 26.975 178.145 27.145 178.315 ;
        RECT 27.435 178.145 27.605 178.315 ;
        RECT 25.305 177.730 25.475 177.900 ;
        RECT 6.935 172.715 7.105 172.885 ;
        RECT 6.935 172.355 7.105 172.525 ;
        RECT 6.935 171.995 7.105 172.165 ;
        RECT 6.935 171.635 7.105 171.805 ;
        RECT 6.935 171.275 7.105 171.445 ;
        RECT 17.700 172.735 17.870 172.905 ;
        RECT 17.700 172.375 17.870 172.545 ;
        RECT 17.700 172.015 17.870 172.185 ;
        RECT 17.700 171.655 17.870 171.825 ;
        RECT 17.700 171.295 17.870 171.465 ;
        RECT 25.305 172.735 25.475 172.905 ;
        RECT 25.305 172.375 25.475 172.545 ;
        RECT 25.305 172.015 25.475 172.185 ;
        RECT 25.305 171.655 25.475 171.825 ;
        RECT 26.515 171.710 26.685 171.880 ;
        RECT 26.975 171.710 27.145 171.880 ;
        RECT 27.435 171.710 27.605 171.880 ;
        RECT 25.305 171.295 25.475 171.465 ;
        RECT 6.935 166.280 7.105 166.450 ;
        RECT 6.935 165.920 7.105 166.090 ;
        RECT 6.935 165.560 7.105 165.730 ;
        RECT 6.935 165.200 7.105 165.370 ;
        RECT 6.935 164.840 7.105 165.010 ;
        RECT 17.700 166.300 17.870 166.470 ;
        RECT 17.700 165.940 17.870 166.110 ;
        RECT 17.700 165.580 17.870 165.750 ;
        RECT 17.700 165.220 17.870 165.390 ;
        RECT 17.700 164.860 17.870 165.030 ;
        RECT 25.305 166.300 25.475 166.470 ;
        RECT 25.305 165.940 25.475 166.110 ;
        RECT 25.305 165.580 25.475 165.750 ;
        RECT 25.305 165.220 25.475 165.390 ;
        RECT 26.515 165.275 26.685 165.445 ;
        RECT 26.975 165.275 27.145 165.445 ;
        RECT 27.435 165.275 27.605 165.445 ;
        RECT 25.305 164.860 25.475 165.030 ;
        RECT 6.935 159.845 7.105 160.015 ;
        RECT 6.935 159.485 7.105 159.655 ;
        RECT 6.935 159.125 7.105 159.295 ;
        RECT 6.935 158.765 7.105 158.935 ;
        RECT 6.935 158.405 7.105 158.575 ;
        RECT 17.700 159.865 17.870 160.035 ;
        RECT 17.700 159.505 17.870 159.675 ;
        RECT 17.700 159.145 17.870 159.315 ;
        RECT 17.700 158.785 17.870 158.955 ;
        RECT 17.700 158.425 17.870 158.595 ;
        RECT 25.305 159.865 25.475 160.035 ;
        RECT 25.305 159.505 25.475 159.675 ;
        RECT 25.305 159.145 25.475 159.315 ;
        RECT 25.305 158.785 25.475 158.955 ;
        RECT 26.515 158.840 26.685 159.010 ;
        RECT 26.975 158.840 27.145 159.010 ;
        RECT 27.435 158.840 27.605 159.010 ;
        RECT 25.305 158.425 25.475 158.595 ;
        RECT 6.935 153.410 7.105 153.580 ;
        RECT 6.935 153.050 7.105 153.220 ;
        RECT 6.935 152.690 7.105 152.860 ;
        RECT 6.935 152.330 7.105 152.500 ;
        RECT 6.935 151.970 7.105 152.140 ;
        RECT 17.700 153.430 17.870 153.600 ;
        RECT 17.700 153.070 17.870 153.240 ;
        RECT 17.700 152.710 17.870 152.880 ;
        RECT 17.700 152.350 17.870 152.520 ;
        RECT 17.700 151.990 17.870 152.160 ;
        RECT 25.305 153.430 25.475 153.600 ;
        RECT 25.305 153.070 25.475 153.240 ;
        RECT 25.305 152.710 25.475 152.880 ;
        RECT 25.305 152.350 25.475 152.520 ;
        RECT 26.515 152.405 26.685 152.575 ;
        RECT 26.975 152.405 27.145 152.575 ;
        RECT 27.435 152.405 27.605 152.575 ;
        RECT 25.305 151.990 25.475 152.160 ;
        RECT 6.935 146.975 7.105 147.145 ;
        RECT 6.935 146.615 7.105 146.785 ;
        RECT 6.935 146.255 7.105 146.425 ;
        RECT 6.935 145.895 7.105 146.065 ;
        RECT 6.935 145.535 7.105 145.705 ;
        RECT 17.700 146.995 17.870 147.165 ;
        RECT 17.700 146.635 17.870 146.805 ;
        RECT 17.700 146.275 17.870 146.445 ;
        RECT 17.700 145.915 17.870 146.085 ;
        RECT 17.700 145.555 17.870 145.725 ;
        RECT 25.305 146.995 25.475 147.165 ;
        RECT 25.305 146.635 25.475 146.805 ;
        RECT 25.305 146.275 25.475 146.445 ;
        RECT 25.305 145.915 25.475 146.085 ;
        RECT 26.515 145.970 26.685 146.140 ;
        RECT 26.975 145.970 27.145 146.140 ;
        RECT 27.435 145.970 27.605 146.140 ;
        RECT 25.305 145.555 25.475 145.725 ;
        RECT 6.935 140.540 7.105 140.710 ;
        RECT 6.935 140.180 7.105 140.350 ;
        RECT 6.935 139.820 7.105 139.990 ;
        RECT 6.935 139.460 7.105 139.630 ;
        RECT 6.935 139.100 7.105 139.270 ;
        RECT 17.700 140.560 17.870 140.730 ;
        RECT 17.700 140.200 17.870 140.370 ;
        RECT 17.700 139.840 17.870 140.010 ;
        RECT 17.700 139.480 17.870 139.650 ;
        RECT 17.700 139.120 17.870 139.290 ;
        RECT 25.305 140.560 25.475 140.730 ;
        RECT 25.305 140.200 25.475 140.370 ;
        RECT 25.305 139.840 25.475 140.010 ;
        RECT 25.305 139.480 25.475 139.650 ;
        RECT 26.515 139.535 26.685 139.705 ;
        RECT 26.975 139.535 27.145 139.705 ;
        RECT 27.435 139.535 27.605 139.705 ;
        RECT 25.305 139.120 25.475 139.290 ;
        RECT 6.935 134.105 7.105 134.275 ;
        RECT 6.935 133.745 7.105 133.915 ;
        RECT 6.935 133.385 7.105 133.555 ;
        RECT 6.935 133.025 7.105 133.195 ;
        RECT 6.935 132.665 7.105 132.835 ;
        RECT 17.700 134.125 17.870 134.295 ;
        RECT 17.700 133.765 17.870 133.935 ;
        RECT 17.700 133.405 17.870 133.575 ;
        RECT 17.700 133.045 17.870 133.215 ;
        RECT 17.700 132.685 17.870 132.855 ;
        RECT 25.305 134.125 25.475 134.295 ;
        RECT 25.305 133.765 25.475 133.935 ;
        RECT 25.305 133.405 25.475 133.575 ;
        RECT 25.305 133.045 25.475 133.215 ;
        RECT 26.515 133.100 26.685 133.270 ;
        RECT 26.975 133.100 27.145 133.270 ;
        RECT 27.435 133.100 27.605 133.270 ;
        RECT 25.305 132.685 25.475 132.855 ;
        RECT 6.935 127.670 7.105 127.840 ;
        RECT 6.935 127.310 7.105 127.480 ;
        RECT 6.935 126.950 7.105 127.120 ;
        RECT 6.935 126.590 7.105 126.760 ;
        RECT 6.935 126.230 7.105 126.400 ;
        RECT 17.700 127.690 17.870 127.860 ;
        RECT 17.700 127.330 17.870 127.500 ;
        RECT 17.700 126.970 17.870 127.140 ;
        RECT 17.700 126.610 17.870 126.780 ;
        RECT 17.700 126.250 17.870 126.420 ;
        RECT 25.305 127.690 25.475 127.860 ;
        RECT 25.305 127.330 25.475 127.500 ;
        RECT 25.305 126.970 25.475 127.140 ;
        RECT 25.305 126.610 25.475 126.780 ;
        RECT 26.515 126.665 26.685 126.835 ;
        RECT 26.975 126.665 27.145 126.835 ;
        RECT 27.435 126.665 27.605 126.835 ;
        RECT 25.305 126.250 25.475 126.420 ;
        RECT 6.935 121.235 7.105 121.405 ;
        RECT 6.935 120.875 7.105 121.045 ;
        RECT 6.935 120.515 7.105 120.685 ;
        RECT 6.935 120.155 7.105 120.325 ;
        RECT 6.935 119.795 7.105 119.965 ;
        RECT 17.700 121.255 17.870 121.425 ;
        RECT 17.700 120.895 17.870 121.065 ;
        RECT 17.700 120.535 17.870 120.705 ;
        RECT 17.700 120.175 17.870 120.345 ;
        RECT 17.700 119.815 17.870 119.985 ;
        RECT 25.305 121.255 25.475 121.425 ;
        RECT 25.305 120.895 25.475 121.065 ;
        RECT 25.305 120.535 25.475 120.705 ;
        RECT 25.305 120.175 25.475 120.345 ;
        RECT 26.515 120.230 26.685 120.400 ;
        RECT 26.975 120.230 27.145 120.400 ;
        RECT 27.435 120.230 27.605 120.400 ;
        RECT 25.305 119.815 25.475 119.985 ;
        RECT 6.935 114.800 7.105 114.970 ;
        RECT 6.935 114.440 7.105 114.610 ;
        RECT 6.935 114.080 7.105 114.250 ;
        RECT 6.935 113.720 7.105 113.890 ;
        RECT 6.935 113.360 7.105 113.530 ;
        RECT 17.700 114.820 17.870 114.990 ;
        RECT 17.700 114.460 17.870 114.630 ;
        RECT 17.700 114.100 17.870 114.270 ;
        RECT 17.700 113.740 17.870 113.910 ;
        RECT 17.700 113.380 17.870 113.550 ;
        RECT 25.305 114.820 25.475 114.990 ;
        RECT 25.305 114.460 25.475 114.630 ;
        RECT 25.305 114.100 25.475 114.270 ;
        RECT 25.305 113.740 25.475 113.910 ;
        RECT 26.515 113.795 26.685 113.965 ;
        RECT 26.975 113.795 27.145 113.965 ;
        RECT 27.435 113.795 27.605 113.965 ;
        RECT 25.305 113.380 25.475 113.550 ;
        RECT 6.935 108.365 7.105 108.535 ;
        RECT 6.935 108.005 7.105 108.175 ;
        RECT 6.935 107.645 7.105 107.815 ;
        RECT 6.935 107.285 7.105 107.455 ;
        RECT 6.935 106.925 7.105 107.095 ;
        RECT 17.700 108.385 17.870 108.555 ;
        RECT 17.700 108.025 17.870 108.195 ;
        RECT 17.700 107.665 17.870 107.835 ;
        RECT 17.700 107.305 17.870 107.475 ;
        RECT 17.700 106.945 17.870 107.115 ;
        RECT 25.305 108.385 25.475 108.555 ;
        RECT 25.305 108.025 25.475 108.195 ;
        RECT 25.305 107.665 25.475 107.835 ;
        RECT 25.305 107.305 25.475 107.475 ;
        RECT 26.515 107.360 26.685 107.530 ;
        RECT 26.975 107.360 27.145 107.530 ;
        RECT 27.435 107.360 27.605 107.530 ;
        RECT 25.305 106.945 25.475 107.115 ;
        RECT 6.935 101.930 7.105 102.100 ;
        RECT 6.935 101.570 7.105 101.740 ;
        RECT 6.935 101.210 7.105 101.380 ;
        RECT 6.935 100.850 7.105 101.020 ;
        RECT 6.935 100.490 7.105 100.660 ;
        RECT 17.700 101.950 17.870 102.120 ;
        RECT 17.700 101.590 17.870 101.760 ;
        RECT 17.700 101.230 17.870 101.400 ;
        RECT 17.700 100.870 17.870 101.040 ;
        RECT 17.700 100.510 17.870 100.680 ;
        RECT 25.305 101.950 25.475 102.120 ;
        RECT 25.305 101.590 25.475 101.760 ;
        RECT 25.305 101.230 25.475 101.400 ;
        RECT 25.305 100.870 25.475 101.040 ;
        RECT 26.515 100.925 26.685 101.095 ;
        RECT 26.975 100.925 27.145 101.095 ;
        RECT 27.435 100.925 27.605 101.095 ;
        RECT 25.305 100.510 25.475 100.680 ;
        RECT 6.935 95.495 7.105 95.665 ;
        RECT 6.935 95.135 7.105 95.305 ;
        RECT 6.935 94.775 7.105 94.945 ;
        RECT 6.935 94.415 7.105 94.585 ;
        RECT 6.935 94.055 7.105 94.225 ;
        RECT 17.700 95.515 17.870 95.685 ;
        RECT 17.700 95.155 17.870 95.325 ;
        RECT 17.700 94.795 17.870 94.965 ;
        RECT 17.700 94.435 17.870 94.605 ;
        RECT 17.700 94.075 17.870 94.245 ;
        RECT 25.305 95.515 25.475 95.685 ;
        RECT 25.305 95.155 25.475 95.325 ;
        RECT 25.305 94.795 25.475 94.965 ;
        RECT 25.305 94.435 25.475 94.605 ;
        RECT 26.515 94.490 26.685 94.660 ;
        RECT 26.975 94.490 27.145 94.660 ;
        RECT 27.435 94.490 27.605 94.660 ;
        RECT 25.305 94.075 25.475 94.245 ;
        RECT 6.935 89.060 7.105 89.230 ;
        RECT 6.935 88.700 7.105 88.870 ;
        RECT 6.935 88.340 7.105 88.510 ;
        RECT 6.935 87.980 7.105 88.150 ;
        RECT 6.935 87.620 7.105 87.790 ;
        RECT 17.700 89.080 17.870 89.250 ;
        RECT 17.700 88.720 17.870 88.890 ;
        RECT 17.700 88.360 17.870 88.530 ;
        RECT 17.700 88.000 17.870 88.170 ;
        RECT 17.700 87.640 17.870 87.810 ;
        RECT 25.305 89.080 25.475 89.250 ;
        RECT 25.305 88.720 25.475 88.890 ;
        RECT 25.305 88.360 25.475 88.530 ;
        RECT 25.305 88.000 25.475 88.170 ;
        RECT 26.515 88.055 26.685 88.225 ;
        RECT 26.975 88.055 27.145 88.225 ;
        RECT 27.435 88.055 27.605 88.225 ;
        RECT 25.305 87.640 25.475 87.810 ;
        RECT 6.935 82.625 7.105 82.795 ;
        RECT 6.935 82.265 7.105 82.435 ;
        RECT 6.935 81.905 7.105 82.075 ;
        RECT 6.935 81.545 7.105 81.715 ;
        RECT 6.935 81.185 7.105 81.355 ;
        RECT 17.700 82.645 17.870 82.815 ;
        RECT 17.700 82.285 17.870 82.455 ;
        RECT 17.700 81.925 17.870 82.095 ;
        RECT 17.700 81.565 17.870 81.735 ;
        RECT 17.700 81.205 17.870 81.375 ;
        RECT 25.305 82.645 25.475 82.815 ;
        RECT 25.305 82.285 25.475 82.455 ;
        RECT 25.305 81.925 25.475 82.095 ;
        RECT 25.305 81.565 25.475 81.735 ;
        RECT 26.515 81.620 26.685 81.790 ;
        RECT 26.975 81.620 27.145 81.790 ;
        RECT 27.435 81.620 27.605 81.790 ;
        RECT 25.305 81.205 25.475 81.375 ;
        RECT 6.935 76.190 7.105 76.360 ;
        RECT 6.935 75.830 7.105 76.000 ;
        RECT 6.935 75.470 7.105 75.640 ;
        RECT 6.935 75.110 7.105 75.280 ;
        RECT 6.935 74.750 7.105 74.920 ;
        RECT 17.700 76.210 17.870 76.380 ;
        RECT 17.700 75.850 17.870 76.020 ;
        RECT 17.700 75.490 17.870 75.660 ;
        RECT 17.700 75.130 17.870 75.300 ;
        RECT 17.700 74.770 17.870 74.940 ;
        RECT 25.305 76.210 25.475 76.380 ;
        RECT 25.305 75.850 25.475 76.020 ;
        RECT 25.305 75.490 25.475 75.660 ;
        RECT 25.305 75.130 25.475 75.300 ;
        RECT 26.515 75.185 26.685 75.355 ;
        RECT 26.975 75.185 27.145 75.355 ;
        RECT 27.435 75.185 27.605 75.355 ;
        RECT 25.305 74.770 25.475 74.940 ;
        RECT 6.935 69.755 7.105 69.925 ;
        RECT 6.935 69.395 7.105 69.565 ;
        RECT 6.935 69.035 7.105 69.205 ;
        RECT 6.935 68.675 7.105 68.845 ;
        RECT 6.935 68.315 7.105 68.485 ;
        RECT 17.700 69.775 17.870 69.945 ;
        RECT 17.700 69.415 17.870 69.585 ;
        RECT 17.700 69.055 17.870 69.225 ;
        RECT 17.700 68.695 17.870 68.865 ;
        RECT 17.700 68.335 17.870 68.505 ;
        RECT 25.305 69.775 25.475 69.945 ;
        RECT 25.305 69.415 25.475 69.585 ;
        RECT 25.305 69.055 25.475 69.225 ;
        RECT 25.305 68.695 25.475 68.865 ;
        RECT 26.515 68.750 26.685 68.920 ;
        RECT 26.975 68.750 27.145 68.920 ;
        RECT 27.435 68.750 27.605 68.920 ;
        RECT 25.305 68.335 25.475 68.505 ;
        RECT 6.935 63.320 7.105 63.490 ;
        RECT 6.935 62.960 7.105 63.130 ;
        RECT 6.935 62.600 7.105 62.770 ;
        RECT 6.935 62.240 7.105 62.410 ;
        RECT 6.935 61.880 7.105 62.050 ;
        RECT 17.700 63.340 17.870 63.510 ;
        RECT 17.700 62.980 17.870 63.150 ;
        RECT 17.700 62.620 17.870 62.790 ;
        RECT 17.700 62.260 17.870 62.430 ;
        RECT 17.700 61.900 17.870 62.070 ;
        RECT 25.305 63.340 25.475 63.510 ;
        RECT 25.305 62.980 25.475 63.150 ;
        RECT 25.305 62.620 25.475 62.790 ;
        RECT 25.305 62.260 25.475 62.430 ;
        RECT 26.515 62.315 26.685 62.485 ;
        RECT 26.975 62.315 27.145 62.485 ;
        RECT 27.435 62.315 27.605 62.485 ;
        RECT 25.305 61.900 25.475 62.070 ;
        RECT 6.935 56.885 7.105 57.055 ;
        RECT 6.935 56.525 7.105 56.695 ;
        RECT 6.935 56.165 7.105 56.335 ;
        RECT 6.935 55.805 7.105 55.975 ;
        RECT 6.935 55.445 7.105 55.615 ;
        RECT 17.700 56.905 17.870 57.075 ;
        RECT 17.700 56.545 17.870 56.715 ;
        RECT 17.700 56.185 17.870 56.355 ;
        RECT 17.700 55.825 17.870 55.995 ;
        RECT 17.700 55.465 17.870 55.635 ;
        RECT 25.305 56.905 25.475 57.075 ;
        RECT 25.305 56.545 25.475 56.715 ;
        RECT 25.305 56.185 25.475 56.355 ;
        RECT 25.305 55.825 25.475 55.995 ;
        RECT 26.515 55.880 26.685 56.050 ;
        RECT 26.975 55.880 27.145 56.050 ;
        RECT 27.435 55.880 27.605 56.050 ;
        RECT 25.305 55.465 25.475 55.635 ;
        RECT 6.935 50.450 7.105 50.620 ;
        RECT 6.935 50.090 7.105 50.260 ;
        RECT 6.935 49.730 7.105 49.900 ;
        RECT 6.935 49.370 7.105 49.540 ;
        RECT 6.935 49.010 7.105 49.180 ;
        RECT 17.700 50.470 17.870 50.640 ;
        RECT 17.700 50.110 17.870 50.280 ;
        RECT 17.700 49.750 17.870 49.920 ;
        RECT 17.700 49.390 17.870 49.560 ;
        RECT 17.700 49.030 17.870 49.200 ;
        RECT 25.305 50.470 25.475 50.640 ;
        RECT 25.305 50.110 25.475 50.280 ;
        RECT 25.305 49.750 25.475 49.920 ;
        RECT 25.305 49.390 25.475 49.560 ;
        RECT 26.515 49.445 26.685 49.615 ;
        RECT 26.975 49.445 27.145 49.615 ;
        RECT 27.435 49.445 27.605 49.615 ;
        RECT 25.305 49.030 25.475 49.200 ;
        RECT 6.935 44.015 7.105 44.185 ;
        RECT 6.935 43.655 7.105 43.825 ;
        RECT 6.935 43.295 7.105 43.465 ;
        RECT 6.935 42.935 7.105 43.105 ;
        RECT 6.935 42.575 7.105 42.745 ;
        RECT 17.700 44.035 17.870 44.205 ;
        RECT 17.700 43.675 17.870 43.845 ;
        RECT 17.700 43.315 17.870 43.485 ;
        RECT 17.700 42.955 17.870 43.125 ;
        RECT 17.700 42.595 17.870 42.765 ;
        RECT 25.305 44.035 25.475 44.205 ;
        RECT 25.305 43.675 25.475 43.845 ;
        RECT 25.305 43.315 25.475 43.485 ;
        RECT 25.305 42.955 25.475 43.125 ;
        RECT 26.515 43.010 26.685 43.180 ;
        RECT 26.975 43.010 27.145 43.180 ;
        RECT 27.435 43.010 27.605 43.180 ;
        RECT 25.305 42.595 25.475 42.765 ;
        RECT 6.935 37.580 7.105 37.750 ;
        RECT 6.935 37.220 7.105 37.390 ;
        RECT 6.935 36.860 7.105 37.030 ;
        RECT 6.935 36.500 7.105 36.670 ;
        RECT 6.935 36.140 7.105 36.310 ;
        RECT 17.700 37.600 17.870 37.770 ;
        RECT 17.700 37.240 17.870 37.410 ;
        RECT 17.700 36.880 17.870 37.050 ;
        RECT 17.700 36.520 17.870 36.690 ;
        RECT 17.700 36.160 17.870 36.330 ;
        RECT 25.305 37.600 25.475 37.770 ;
        RECT 25.305 37.240 25.475 37.410 ;
        RECT 25.305 36.880 25.475 37.050 ;
        RECT 25.305 36.520 25.475 36.690 ;
        RECT 26.515 36.575 26.685 36.745 ;
        RECT 26.975 36.575 27.145 36.745 ;
        RECT 27.435 36.575 27.605 36.745 ;
        RECT 25.305 36.160 25.475 36.330 ;
        RECT 6.935 31.145 7.105 31.315 ;
        RECT 6.935 30.785 7.105 30.955 ;
        RECT 6.935 30.425 7.105 30.595 ;
        RECT 6.935 30.065 7.105 30.235 ;
        RECT 6.935 29.705 7.105 29.875 ;
        RECT 17.700 31.165 17.870 31.335 ;
        RECT 17.700 30.805 17.870 30.975 ;
        RECT 17.700 30.445 17.870 30.615 ;
        RECT 17.700 30.085 17.870 30.255 ;
        RECT 17.700 29.725 17.870 29.895 ;
        RECT 25.305 31.165 25.475 31.335 ;
        RECT 25.305 30.805 25.475 30.975 ;
        RECT 25.305 30.445 25.475 30.615 ;
        RECT 25.305 30.085 25.475 30.255 ;
        RECT 26.515 30.140 26.685 30.310 ;
        RECT 26.975 30.140 27.145 30.310 ;
        RECT 27.435 30.140 27.605 30.310 ;
        RECT 25.305 29.725 25.475 29.895 ;
        RECT 6.935 24.710 7.105 24.880 ;
        RECT 6.935 24.350 7.105 24.520 ;
        RECT 6.935 23.990 7.105 24.160 ;
        RECT 6.935 23.630 7.105 23.800 ;
        RECT 6.935 23.270 7.105 23.440 ;
        RECT 17.700 24.730 17.870 24.900 ;
        RECT 17.700 24.370 17.870 24.540 ;
        RECT 17.700 24.010 17.870 24.180 ;
        RECT 17.700 23.650 17.870 23.820 ;
        RECT 17.700 23.290 17.870 23.460 ;
        RECT 25.305 24.730 25.475 24.900 ;
        RECT 25.305 24.370 25.475 24.540 ;
        RECT 25.305 24.010 25.475 24.180 ;
        RECT 25.305 23.650 25.475 23.820 ;
        RECT 26.515 23.705 26.685 23.875 ;
        RECT 26.975 23.705 27.145 23.875 ;
        RECT 27.435 23.705 27.605 23.875 ;
        RECT 25.305 23.290 25.475 23.460 ;
        RECT 6.935 18.275 7.105 18.445 ;
        RECT 6.935 17.915 7.105 18.085 ;
        RECT 6.935 17.555 7.105 17.725 ;
        RECT 6.935 17.195 7.105 17.365 ;
        RECT 6.935 16.835 7.105 17.005 ;
        RECT 17.700 18.295 17.870 18.465 ;
        RECT 17.700 17.935 17.870 18.105 ;
        RECT 17.700 17.575 17.870 17.745 ;
        RECT 17.700 17.215 17.870 17.385 ;
        RECT 17.700 16.855 17.870 17.025 ;
        RECT 25.305 18.295 25.475 18.465 ;
        RECT 25.305 17.935 25.475 18.105 ;
        RECT 25.305 17.575 25.475 17.745 ;
        RECT 25.305 17.215 25.475 17.385 ;
        RECT 26.515 17.270 26.685 17.440 ;
        RECT 26.975 17.270 27.145 17.440 ;
        RECT 27.435 17.270 27.605 17.440 ;
        RECT 25.305 16.855 25.475 17.025 ;
        RECT 6.935 11.840 7.105 12.010 ;
        RECT 6.935 11.480 7.105 11.650 ;
        RECT 6.935 11.120 7.105 11.290 ;
        RECT 6.935 10.760 7.105 10.930 ;
        RECT 6.935 10.400 7.105 10.570 ;
        RECT 17.700 11.860 17.870 12.030 ;
        RECT 17.700 11.500 17.870 11.670 ;
        RECT 17.700 11.140 17.870 11.310 ;
        RECT 17.700 10.780 17.870 10.950 ;
        RECT 17.700 10.420 17.870 10.590 ;
        RECT 25.305 11.860 25.475 12.030 ;
        RECT 25.305 11.500 25.475 11.670 ;
        RECT 25.305 11.140 25.475 11.310 ;
        RECT 25.305 10.780 25.475 10.950 ;
        RECT 26.515 10.835 26.685 11.005 ;
        RECT 26.975 10.835 27.145 11.005 ;
        RECT 27.435 10.835 27.605 11.005 ;
        RECT 25.305 10.420 25.475 10.590 ;
        RECT 6.935 5.405 7.105 5.575 ;
        RECT 6.935 5.045 7.105 5.215 ;
        RECT 6.935 4.685 7.105 4.855 ;
        RECT 6.935 4.325 7.105 4.495 ;
        RECT 6.935 3.965 7.105 4.135 ;
        RECT 17.700 5.425 17.870 5.595 ;
        RECT 17.700 5.065 17.870 5.235 ;
        RECT 17.700 4.705 17.870 4.875 ;
        RECT 17.700 4.345 17.870 4.515 ;
        RECT 17.700 3.985 17.870 4.155 ;
        RECT 25.305 5.425 25.475 5.595 ;
        RECT 25.305 5.065 25.475 5.235 ;
        RECT 25.305 4.705 25.475 4.875 ;
        RECT 25.305 4.345 25.475 4.515 ;
        RECT 26.515 4.400 26.685 4.570 ;
        RECT 26.975 4.400 27.145 4.570 ;
        RECT 27.435 4.400 27.605 4.570 ;
        RECT 25.305 3.985 25.475 4.155 ;
      LAYER met1 ;
        RECT 6.905 207.150 17.915 207.160 ;
        RECT 6.905 206.930 25.545 207.150 ;
        RECT 6.905 203.760 7.135 206.930 ;
        RECT 17.685 206.920 25.545 206.930 ;
        RECT 17.685 206.190 17.915 206.920 ;
        RECT 25.315 206.190 25.545 206.920 ;
        RECT 17.670 206.050 17.915 206.190 ;
        RECT 6.905 203.750 10.800 203.760 ;
        RECT 6.905 203.495 11.000 203.750 ;
        RECT 6.900 203.210 11.000 203.495 ;
        RECT 17.670 203.250 17.900 206.050 ;
        RECT 25.275 206.030 25.545 206.190 ;
        RECT 25.275 204.205 25.505 206.030 ;
        RECT 26.370 204.205 27.750 204.210 ;
        RECT 25.275 203.730 27.750 204.205 ;
        RECT 25.275 203.250 25.505 203.730 ;
        RECT 6.900 203.200 10.800 203.210 ;
        RECT 6.905 197.325 7.135 199.735 ;
        RECT 6.905 197.315 10.800 197.325 ;
        RECT 6.905 197.060 11.000 197.315 ;
        RECT 6.900 196.775 11.000 197.060 ;
        RECT 17.670 196.815 17.900 199.755 ;
        RECT 25.275 197.770 25.505 199.755 ;
        RECT 26.370 197.770 27.750 197.775 ;
        RECT 25.275 197.295 27.750 197.770 ;
        RECT 25.275 196.815 25.505 197.295 ;
        RECT 6.900 196.765 10.800 196.775 ;
        RECT 6.905 190.890 7.135 193.300 ;
        RECT 6.905 190.880 10.800 190.890 ;
        RECT 6.905 190.625 11.000 190.880 ;
        RECT 6.900 190.340 11.000 190.625 ;
        RECT 17.670 190.380 17.900 193.320 ;
        RECT 25.275 191.335 25.505 193.320 ;
        RECT 26.370 191.335 27.750 191.340 ;
        RECT 25.275 190.860 27.750 191.335 ;
        RECT 25.275 190.380 25.505 190.860 ;
        RECT 6.900 190.330 10.800 190.340 ;
        RECT 6.905 184.455 7.135 186.865 ;
        RECT 6.905 184.445 10.800 184.455 ;
        RECT 6.905 184.190 11.000 184.445 ;
        RECT 6.900 183.905 11.000 184.190 ;
        RECT 17.670 183.945 17.900 186.885 ;
        RECT 25.275 184.900 25.505 186.885 ;
        RECT 26.370 184.900 27.750 184.905 ;
        RECT 25.275 184.425 27.750 184.900 ;
        RECT 25.275 183.945 25.505 184.425 ;
        RECT 6.900 183.895 10.800 183.905 ;
        RECT 6.905 178.020 7.135 180.430 ;
        RECT 6.905 178.010 10.800 178.020 ;
        RECT 6.905 177.755 11.000 178.010 ;
        RECT 6.900 177.470 11.000 177.755 ;
        RECT 17.670 177.510 17.900 180.450 ;
        RECT 25.275 178.465 25.505 180.450 ;
        RECT 26.370 178.465 27.750 178.470 ;
        RECT 25.275 177.990 27.750 178.465 ;
        RECT 25.275 177.510 25.505 177.990 ;
        RECT 6.900 177.460 10.800 177.470 ;
        RECT 6.905 171.585 7.135 173.995 ;
        RECT 6.905 171.575 10.800 171.585 ;
        RECT 6.905 171.320 11.000 171.575 ;
        RECT 6.900 171.035 11.000 171.320 ;
        RECT 17.670 171.075 17.900 174.015 ;
        RECT 25.275 172.030 25.505 174.015 ;
        RECT 26.370 172.030 27.750 172.035 ;
        RECT 25.275 171.555 27.750 172.030 ;
        RECT 25.275 171.075 25.505 171.555 ;
        RECT 6.900 171.025 10.800 171.035 ;
        RECT 6.905 165.150 7.135 167.560 ;
        RECT 6.905 165.140 10.800 165.150 ;
        RECT 6.905 164.885 11.000 165.140 ;
        RECT 6.900 164.600 11.000 164.885 ;
        RECT 17.670 164.640 17.900 167.580 ;
        RECT 25.275 165.595 25.505 167.580 ;
        RECT 26.370 165.595 27.750 165.600 ;
        RECT 25.275 165.120 27.750 165.595 ;
        RECT 25.275 164.640 25.505 165.120 ;
        RECT 6.900 164.590 10.800 164.600 ;
        RECT 6.905 158.715 7.135 161.125 ;
        RECT 6.905 158.705 10.800 158.715 ;
        RECT 6.905 158.450 11.000 158.705 ;
        RECT 6.900 158.165 11.000 158.450 ;
        RECT 17.670 158.205 17.900 161.145 ;
        RECT 25.275 159.160 25.505 161.145 ;
        RECT 26.370 159.160 27.750 159.165 ;
        RECT 25.275 158.685 27.750 159.160 ;
        RECT 25.275 158.205 25.505 158.685 ;
        RECT 6.900 158.155 10.800 158.165 ;
        RECT 6.905 152.280 7.135 154.690 ;
        RECT 6.905 152.270 10.800 152.280 ;
        RECT 6.905 152.015 11.000 152.270 ;
        RECT 6.900 151.730 11.000 152.015 ;
        RECT 17.670 151.770 17.900 154.710 ;
        RECT 25.275 152.725 25.505 154.710 ;
        RECT 26.370 152.725 27.750 152.730 ;
        RECT 25.275 152.250 27.750 152.725 ;
        RECT 25.275 151.770 25.505 152.250 ;
        RECT 6.900 151.720 10.800 151.730 ;
        RECT 6.905 145.845 7.135 148.255 ;
        RECT 6.905 145.835 10.800 145.845 ;
        RECT 6.905 145.580 11.000 145.835 ;
        RECT 6.900 145.295 11.000 145.580 ;
        RECT 17.670 145.335 17.900 148.275 ;
        RECT 25.275 146.290 25.505 148.275 ;
        RECT 26.370 146.290 27.750 146.295 ;
        RECT 25.275 145.815 27.750 146.290 ;
        RECT 25.275 145.335 25.505 145.815 ;
        RECT 6.900 145.285 10.800 145.295 ;
        RECT 6.905 139.410 7.135 141.820 ;
        RECT 6.905 139.400 10.800 139.410 ;
        RECT 6.905 139.145 11.000 139.400 ;
        RECT 6.900 138.860 11.000 139.145 ;
        RECT 17.670 138.900 17.900 141.840 ;
        RECT 25.275 139.855 25.505 141.840 ;
        RECT 26.370 139.855 27.750 139.860 ;
        RECT 25.275 139.380 27.750 139.855 ;
        RECT 25.275 138.900 25.505 139.380 ;
        RECT 6.900 138.850 10.800 138.860 ;
        RECT 6.905 132.975 7.135 135.385 ;
        RECT 6.905 132.965 10.800 132.975 ;
        RECT 6.905 132.710 11.000 132.965 ;
        RECT 6.900 132.425 11.000 132.710 ;
        RECT 17.670 132.465 17.900 135.405 ;
        RECT 25.275 133.420 25.505 135.405 ;
        RECT 26.370 133.420 27.750 133.425 ;
        RECT 25.275 132.945 27.750 133.420 ;
        RECT 25.275 132.465 25.505 132.945 ;
        RECT 6.900 132.415 10.800 132.425 ;
        RECT 6.905 126.540 7.135 128.950 ;
        RECT 6.905 126.530 10.800 126.540 ;
        RECT 6.905 126.275 11.000 126.530 ;
        RECT 6.900 125.990 11.000 126.275 ;
        RECT 17.670 126.030 17.900 128.970 ;
        RECT 25.275 126.985 25.505 128.970 ;
        RECT 26.370 126.985 27.750 126.990 ;
        RECT 25.275 126.510 27.750 126.985 ;
        RECT 25.275 126.030 25.505 126.510 ;
        RECT 6.900 125.980 10.800 125.990 ;
        RECT 6.905 120.105 7.135 122.515 ;
        RECT 6.905 120.095 10.800 120.105 ;
        RECT 6.905 119.840 11.000 120.095 ;
        RECT 6.900 119.555 11.000 119.840 ;
        RECT 17.670 119.595 17.900 122.535 ;
        RECT 25.275 120.550 25.505 122.535 ;
        RECT 26.370 120.550 27.750 120.555 ;
        RECT 25.275 120.075 27.750 120.550 ;
        RECT 25.275 119.595 25.505 120.075 ;
        RECT 6.900 119.545 10.800 119.555 ;
        RECT 6.905 113.670 7.135 116.080 ;
        RECT 6.905 113.660 10.800 113.670 ;
        RECT 6.905 113.405 11.000 113.660 ;
        RECT 6.900 113.120 11.000 113.405 ;
        RECT 17.670 113.160 17.900 116.100 ;
        RECT 25.275 114.115 25.505 116.100 ;
        RECT 26.370 114.115 27.750 114.120 ;
        RECT 25.275 113.640 27.750 114.115 ;
        RECT 25.275 113.160 25.505 113.640 ;
        RECT 6.900 113.110 10.800 113.120 ;
        RECT 6.905 107.235 7.135 109.645 ;
        RECT 6.905 107.225 10.800 107.235 ;
        RECT 6.905 106.970 11.000 107.225 ;
        RECT 6.900 106.685 11.000 106.970 ;
        RECT 17.670 106.725 17.900 109.665 ;
        RECT 25.275 107.680 25.505 109.665 ;
        RECT 26.370 107.680 27.750 107.685 ;
        RECT 25.275 107.205 27.750 107.680 ;
        RECT 25.275 106.725 25.505 107.205 ;
        RECT 6.900 106.675 10.800 106.685 ;
        RECT 6.905 100.800 7.135 103.210 ;
        RECT 6.905 100.790 10.800 100.800 ;
        RECT 6.905 100.535 11.000 100.790 ;
        RECT 6.900 100.250 11.000 100.535 ;
        RECT 17.670 100.290 17.900 103.230 ;
        RECT 25.275 101.245 25.505 103.230 ;
        RECT 26.370 101.245 27.750 101.250 ;
        RECT 25.275 100.770 27.750 101.245 ;
        RECT 25.275 100.290 25.505 100.770 ;
        RECT 6.900 100.240 10.800 100.250 ;
        RECT 6.905 94.365 7.135 96.775 ;
        RECT 6.905 94.355 10.800 94.365 ;
        RECT 6.905 94.100 11.000 94.355 ;
        RECT 6.900 93.815 11.000 94.100 ;
        RECT 17.670 93.855 17.900 96.795 ;
        RECT 25.275 94.810 25.505 96.795 ;
        RECT 26.370 94.810 27.750 94.815 ;
        RECT 25.275 94.335 27.750 94.810 ;
        RECT 25.275 93.855 25.505 94.335 ;
        RECT 6.900 93.805 10.800 93.815 ;
        RECT 6.905 87.930 7.135 90.340 ;
        RECT 6.905 87.920 10.800 87.930 ;
        RECT 6.905 87.665 11.000 87.920 ;
        RECT 6.900 87.380 11.000 87.665 ;
        RECT 17.670 87.420 17.900 90.360 ;
        RECT 25.275 88.375 25.505 90.360 ;
        RECT 26.370 88.375 27.750 88.380 ;
        RECT 25.275 87.900 27.750 88.375 ;
        RECT 25.275 87.420 25.505 87.900 ;
        RECT 6.900 87.370 10.800 87.380 ;
        RECT 6.905 81.495 7.135 83.905 ;
        RECT 6.905 81.485 10.800 81.495 ;
        RECT 6.905 81.230 11.000 81.485 ;
        RECT 6.900 80.945 11.000 81.230 ;
        RECT 17.670 80.985 17.900 83.925 ;
        RECT 25.275 81.940 25.505 83.925 ;
        RECT 26.370 81.940 27.750 81.945 ;
        RECT 25.275 81.465 27.750 81.940 ;
        RECT 25.275 80.985 25.505 81.465 ;
        RECT 6.900 80.935 10.800 80.945 ;
        RECT 6.905 75.060 7.135 77.470 ;
        RECT 6.905 75.050 10.800 75.060 ;
        RECT 6.905 74.795 11.000 75.050 ;
        RECT 6.900 74.510 11.000 74.795 ;
        RECT 17.670 74.550 17.900 77.490 ;
        RECT 25.275 75.505 25.505 77.490 ;
        RECT 26.370 75.505 27.750 75.510 ;
        RECT 25.275 75.030 27.750 75.505 ;
        RECT 25.275 74.550 25.505 75.030 ;
        RECT 6.900 74.500 10.800 74.510 ;
        RECT 6.905 68.625 7.135 71.035 ;
        RECT 6.905 68.615 10.800 68.625 ;
        RECT 6.905 68.360 11.000 68.615 ;
        RECT 6.900 68.075 11.000 68.360 ;
        RECT 17.670 68.115 17.900 71.055 ;
        RECT 25.275 69.070 25.505 71.055 ;
        RECT 26.370 69.070 27.750 69.075 ;
        RECT 25.275 68.595 27.750 69.070 ;
        RECT 25.275 68.115 25.505 68.595 ;
        RECT 6.900 68.065 10.800 68.075 ;
        RECT 6.905 62.190 7.135 64.600 ;
        RECT 6.905 62.180 10.800 62.190 ;
        RECT 6.905 61.925 11.000 62.180 ;
        RECT 6.900 61.640 11.000 61.925 ;
        RECT 17.670 61.680 17.900 64.620 ;
        RECT 25.275 62.635 25.505 64.620 ;
        RECT 26.370 62.635 27.750 62.640 ;
        RECT 25.275 62.160 27.750 62.635 ;
        RECT 25.275 61.680 25.505 62.160 ;
        RECT 6.900 61.630 10.800 61.640 ;
        RECT 6.905 55.755 7.135 58.165 ;
        RECT 6.905 55.745 10.800 55.755 ;
        RECT 6.905 55.490 11.000 55.745 ;
        RECT 6.900 55.205 11.000 55.490 ;
        RECT 17.670 55.245 17.900 58.185 ;
        RECT 25.275 56.200 25.505 58.185 ;
        RECT 26.370 56.200 27.750 56.205 ;
        RECT 25.275 55.725 27.750 56.200 ;
        RECT 25.275 55.245 25.505 55.725 ;
        RECT 6.900 55.195 10.800 55.205 ;
        RECT 6.905 49.320 7.135 51.730 ;
        RECT 6.905 49.310 10.800 49.320 ;
        RECT 6.905 49.055 11.000 49.310 ;
        RECT 6.900 48.770 11.000 49.055 ;
        RECT 17.670 48.810 17.900 51.750 ;
        RECT 25.275 49.765 25.505 51.750 ;
        RECT 26.370 49.765 27.750 49.770 ;
        RECT 25.275 49.290 27.750 49.765 ;
        RECT 25.275 48.810 25.505 49.290 ;
        RECT 6.900 48.760 10.800 48.770 ;
        RECT 6.905 42.885 7.135 45.295 ;
        RECT 6.905 42.875 10.800 42.885 ;
        RECT 6.905 42.620 11.000 42.875 ;
        RECT 6.900 42.335 11.000 42.620 ;
        RECT 17.670 42.375 17.900 45.315 ;
        RECT 25.275 43.330 25.505 45.315 ;
        RECT 26.370 43.330 27.750 43.335 ;
        RECT 25.275 42.855 27.750 43.330 ;
        RECT 25.275 42.375 25.505 42.855 ;
        RECT 6.900 42.325 10.800 42.335 ;
        RECT 6.905 36.450 7.135 38.860 ;
        RECT 6.905 36.440 10.800 36.450 ;
        RECT 6.905 36.185 11.000 36.440 ;
        RECT 6.900 35.900 11.000 36.185 ;
        RECT 17.670 35.940 17.900 38.880 ;
        RECT 25.275 36.895 25.505 38.880 ;
        RECT 26.370 36.895 27.750 36.900 ;
        RECT 25.275 36.420 27.750 36.895 ;
        RECT 25.275 35.940 25.505 36.420 ;
        RECT 6.900 35.890 10.800 35.900 ;
        RECT 6.905 30.015 7.135 32.425 ;
        RECT 6.905 30.005 10.800 30.015 ;
        RECT 6.905 29.750 11.000 30.005 ;
        RECT 6.900 29.465 11.000 29.750 ;
        RECT 17.670 29.505 17.900 32.445 ;
        RECT 25.275 30.460 25.505 32.445 ;
        RECT 26.370 30.460 27.750 30.465 ;
        RECT 25.275 29.985 27.750 30.460 ;
        RECT 25.275 29.505 25.505 29.985 ;
        RECT 6.900 29.455 10.800 29.465 ;
        RECT 6.905 23.580 7.135 25.990 ;
        RECT 6.905 23.570 10.800 23.580 ;
        RECT 6.905 23.315 11.000 23.570 ;
        RECT 6.900 23.030 11.000 23.315 ;
        RECT 17.670 23.070 17.900 26.010 ;
        RECT 25.275 24.025 25.505 26.010 ;
        RECT 26.370 24.025 27.750 24.030 ;
        RECT 25.275 23.550 27.750 24.025 ;
        RECT 25.275 23.070 25.505 23.550 ;
        RECT 6.900 23.020 10.800 23.030 ;
        RECT 6.905 17.145 7.135 19.555 ;
        RECT 6.905 17.135 10.800 17.145 ;
        RECT 6.905 16.880 11.000 17.135 ;
        RECT 6.900 16.595 11.000 16.880 ;
        RECT 17.670 16.635 17.900 19.575 ;
        RECT 25.275 17.590 25.505 19.575 ;
        RECT 26.370 17.590 27.750 17.595 ;
        RECT 25.275 17.115 27.750 17.590 ;
        RECT 25.275 16.635 25.505 17.115 ;
        RECT 6.900 16.585 10.800 16.595 ;
        RECT 6.905 10.710 7.135 13.120 ;
        RECT 6.905 10.700 10.800 10.710 ;
        RECT 6.905 10.445 11.000 10.700 ;
        RECT 6.900 10.160 11.000 10.445 ;
        RECT 17.670 10.200 17.900 13.140 ;
        RECT 25.275 11.155 25.505 13.140 ;
        RECT 26.370 11.155 27.750 11.160 ;
        RECT 25.275 10.680 27.750 11.155 ;
        RECT 25.275 10.200 25.505 10.680 ;
        RECT 6.900 10.150 10.800 10.160 ;
        RECT 6.905 4.275 7.135 6.685 ;
        RECT 6.905 4.265 10.800 4.275 ;
        RECT 6.905 4.010 11.000 4.265 ;
        RECT 6.900 3.725 11.000 4.010 ;
        RECT 17.670 3.765 17.900 6.705 ;
        RECT 25.275 4.720 25.505 6.705 ;
        RECT 26.370 4.720 27.750 4.725 ;
        RECT 25.275 4.245 27.750 4.720 ;
        RECT 25.275 3.765 25.505 4.245 ;
        RECT 6.900 3.715 10.800 3.725 ;
      LAYER via ;
        RECT 10.280 203.210 10.950 203.750 ;
        RECT 10.280 196.775 10.950 197.315 ;
        RECT 10.280 190.340 10.950 190.880 ;
        RECT 10.280 183.905 10.950 184.445 ;
        RECT 10.280 177.470 10.950 178.010 ;
        RECT 10.280 171.035 10.950 171.575 ;
        RECT 10.280 164.600 10.950 165.140 ;
        RECT 10.280 158.165 10.950 158.705 ;
        RECT 10.280 151.730 10.950 152.270 ;
        RECT 10.280 145.295 10.950 145.835 ;
        RECT 10.280 138.860 10.950 139.400 ;
        RECT 10.280 132.425 10.950 132.965 ;
        RECT 10.280 125.990 10.950 126.530 ;
        RECT 10.280 119.555 10.950 120.095 ;
        RECT 10.280 113.120 10.950 113.660 ;
        RECT 10.280 106.685 10.950 107.225 ;
        RECT 10.280 100.250 10.950 100.790 ;
        RECT 10.280 93.815 10.950 94.355 ;
        RECT 10.280 87.380 10.950 87.920 ;
        RECT 10.280 80.945 10.950 81.485 ;
        RECT 10.280 74.510 10.950 75.050 ;
        RECT 10.280 68.075 10.950 68.615 ;
        RECT 10.280 61.640 10.950 62.180 ;
        RECT 10.280 55.205 10.950 55.745 ;
        RECT 10.280 48.770 10.950 49.310 ;
        RECT 10.280 42.335 10.950 42.875 ;
        RECT 10.280 35.900 10.950 36.440 ;
        RECT 10.280 29.465 10.950 30.005 ;
        RECT 10.280 23.030 10.950 23.570 ;
        RECT 10.280 16.595 10.950 17.135 ;
        RECT 10.280 10.160 10.950 10.700 ;
        RECT 10.280 3.725 10.950 4.265 ;
      LAYER met2 ;
        RECT 10.280 203.800 10.930 206.470 ;
        RECT 10.280 202.560 10.950 203.800 ;
        RECT 10.280 197.365 10.930 202.560 ;
        RECT 10.280 196.125 10.950 197.365 ;
        RECT 10.280 190.930 10.930 196.125 ;
        RECT 10.280 189.690 10.950 190.930 ;
        RECT 10.280 184.495 10.930 189.690 ;
        RECT 10.280 183.255 10.950 184.495 ;
        RECT 10.280 178.060 10.930 183.255 ;
        RECT 10.280 176.820 10.950 178.060 ;
        RECT 10.280 171.625 10.930 176.820 ;
        RECT 10.280 170.385 10.950 171.625 ;
        RECT 10.280 165.190 10.930 170.385 ;
        RECT 10.280 163.950 10.950 165.190 ;
        RECT 10.280 158.755 10.930 163.950 ;
        RECT 10.280 157.515 10.950 158.755 ;
        RECT 10.280 152.320 10.930 157.515 ;
        RECT 10.280 151.080 10.950 152.320 ;
        RECT 10.280 145.885 10.930 151.080 ;
        RECT 10.280 144.645 10.950 145.885 ;
        RECT 10.280 139.450 10.930 144.645 ;
        RECT 10.280 138.210 10.950 139.450 ;
        RECT 10.280 133.015 10.930 138.210 ;
        RECT 10.280 131.775 10.950 133.015 ;
        RECT 10.280 126.580 10.930 131.775 ;
        RECT 10.280 125.340 10.950 126.580 ;
        RECT 10.280 120.145 10.930 125.340 ;
        RECT 10.280 118.905 10.950 120.145 ;
        RECT 10.280 113.710 10.930 118.905 ;
        RECT 10.280 112.470 10.950 113.710 ;
        RECT 10.280 107.275 10.930 112.470 ;
        RECT 10.280 106.035 10.950 107.275 ;
        RECT 10.280 100.840 10.930 106.035 ;
        RECT 10.280 99.600 10.950 100.840 ;
        RECT 10.280 94.405 10.930 99.600 ;
        RECT 10.280 93.165 10.950 94.405 ;
        RECT 10.280 87.970 10.930 93.165 ;
        RECT 10.280 86.730 10.950 87.970 ;
        RECT 10.280 81.535 10.930 86.730 ;
        RECT 10.280 80.295 10.950 81.535 ;
        RECT 10.280 75.100 10.930 80.295 ;
        RECT 10.280 73.860 10.950 75.100 ;
        RECT 10.280 68.665 10.930 73.860 ;
        RECT 10.280 67.425 10.950 68.665 ;
        RECT 10.280 62.230 10.930 67.425 ;
        RECT 10.280 60.990 10.950 62.230 ;
        RECT 10.280 55.795 10.930 60.990 ;
        RECT 10.280 54.555 10.950 55.795 ;
        RECT 10.280 49.360 10.930 54.555 ;
        RECT 10.280 48.120 10.950 49.360 ;
        RECT 10.280 42.925 10.930 48.120 ;
        RECT 10.280 41.685 10.950 42.925 ;
        RECT 10.280 36.490 10.930 41.685 ;
        RECT 10.280 35.250 10.950 36.490 ;
        RECT 10.280 30.055 10.930 35.250 ;
        RECT 10.280 28.815 10.950 30.055 ;
        RECT 10.280 23.620 10.930 28.815 ;
        RECT 10.280 22.380 10.950 23.620 ;
        RECT 10.280 17.185 10.930 22.380 ;
        RECT 10.280 15.945 10.950 17.185 ;
        RECT 10.280 10.750 10.930 15.945 ;
        RECT 10.280 9.510 10.950 10.750 ;
        RECT 10.280 4.315 10.930 9.510 ;
        RECT 10.280 3.075 10.950 4.315 ;
        RECT 10.280 0.725 10.930 3.075 ;
    END
  END VDD
  PIN in[0]
    DIRECTION INOUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.102000 ;
    PORT
      LAYER li1 ;
        RECT 2.045 203.400 2.215 204.800 ;
        RECT 3.005 203.400 3.175 204.800 ;
        RECT 3.965 203.400 4.135 204.800 ;
        RECT 4.925 203.400 5.095 204.800 ;
        RECT 5.885 203.400 6.055 204.800 ;
        RECT 2.045 201.340 2.215 201.900 ;
        RECT 3.005 201.340 3.175 201.900 ;
        RECT 3.965 201.340 4.135 201.900 ;
        RECT 4.925 201.340 5.095 201.900 ;
        RECT 5.885 201.340 6.055 201.900 ;
      LAYER mcon ;
        RECT 2.045 204.375 2.215 204.545 ;
        RECT 2.045 204.015 2.215 204.185 ;
        RECT 2.045 203.655 2.215 203.825 ;
        RECT 3.005 204.375 3.175 204.545 ;
        RECT 3.005 204.015 3.175 204.185 ;
        RECT 3.005 203.655 3.175 203.825 ;
        RECT 3.965 204.375 4.135 204.545 ;
        RECT 3.965 204.015 4.135 204.185 ;
        RECT 3.965 203.655 4.135 203.825 ;
        RECT 4.925 204.375 5.095 204.545 ;
        RECT 4.925 204.015 5.095 204.185 ;
        RECT 4.925 203.655 5.095 203.825 ;
        RECT 5.885 204.375 6.055 204.545 ;
        RECT 5.885 204.015 6.055 204.185 ;
        RECT 5.885 203.655 6.055 203.825 ;
        RECT 2.045 201.535 2.215 201.705 ;
        RECT 3.005 201.535 3.175 201.705 ;
        RECT 3.965 201.535 4.135 201.705 ;
        RECT 4.925 201.535 5.095 201.705 ;
        RECT 5.885 201.535 6.055 201.705 ;
      LAYER met1 ;
        RECT 0.645 205.530 6.055 205.700 ;
        RECT 0.645 202.715 0.815 205.530 ;
        RECT 2.045 204.780 2.215 205.530 ;
        RECT 3.005 204.780 3.175 205.530 ;
        RECT 3.965 204.780 4.135 205.530 ;
        RECT 4.925 204.780 5.095 205.530 ;
        RECT 5.885 204.780 6.055 205.530 ;
        RECT 2.015 203.420 2.245 204.780 ;
        RECT 2.975 203.420 3.205 204.780 ;
        RECT 3.935 203.420 4.165 204.780 ;
        RECT 4.895 203.420 5.125 204.780 ;
        RECT 5.855 203.420 6.085 204.780 ;
        RECT 0.000 202.545 0.815 202.715 ;
        RECT 0.010 202.540 0.150 202.545 ;
        RECT 0.645 200.660 0.815 202.545 ;
        RECT 2.015 201.360 2.245 201.880 ;
        RECT 2.975 201.360 3.205 201.880 ;
        RECT 3.935 201.360 4.165 201.880 ;
        RECT 4.895 201.360 5.125 201.880 ;
        RECT 5.855 201.360 6.085 201.880 ;
        RECT 2.045 200.660 2.215 201.360 ;
        RECT 3.005 200.660 3.175 201.360 ;
        RECT 3.965 200.660 4.135 201.360 ;
        RECT 4.925 200.660 5.095 201.360 ;
        RECT 5.885 200.660 6.055 201.360 ;
        RECT 0.645 200.490 6.055 200.660 ;
    END
  END in[0]
  PIN in[1]
    DIRECTION INOUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.102000 ;
    PORT
      LAYER li1 ;
        RECT 2.045 196.965 2.215 198.365 ;
        RECT 3.005 196.965 3.175 198.365 ;
        RECT 3.965 196.965 4.135 198.365 ;
        RECT 4.925 196.965 5.095 198.365 ;
        RECT 5.885 196.965 6.055 198.365 ;
        RECT 2.045 194.905 2.215 195.465 ;
        RECT 3.005 194.905 3.175 195.465 ;
        RECT 3.965 194.905 4.135 195.465 ;
        RECT 4.925 194.905 5.095 195.465 ;
        RECT 5.885 194.905 6.055 195.465 ;
      LAYER mcon ;
        RECT 2.045 197.940 2.215 198.110 ;
        RECT 2.045 197.580 2.215 197.750 ;
        RECT 2.045 197.220 2.215 197.390 ;
        RECT 3.005 197.940 3.175 198.110 ;
        RECT 3.005 197.580 3.175 197.750 ;
        RECT 3.005 197.220 3.175 197.390 ;
        RECT 3.965 197.940 4.135 198.110 ;
        RECT 3.965 197.580 4.135 197.750 ;
        RECT 3.965 197.220 4.135 197.390 ;
        RECT 4.925 197.940 5.095 198.110 ;
        RECT 4.925 197.580 5.095 197.750 ;
        RECT 4.925 197.220 5.095 197.390 ;
        RECT 5.885 197.940 6.055 198.110 ;
        RECT 5.885 197.580 6.055 197.750 ;
        RECT 5.885 197.220 6.055 197.390 ;
        RECT 2.045 195.100 2.215 195.270 ;
        RECT 3.005 195.100 3.175 195.270 ;
        RECT 3.965 195.100 4.135 195.270 ;
        RECT 4.925 195.100 5.095 195.270 ;
        RECT 5.885 195.100 6.055 195.270 ;
      LAYER met1 ;
        RECT 0.645 199.095 6.055 199.265 ;
        RECT 0.645 196.280 0.815 199.095 ;
        RECT 2.045 198.345 2.215 199.095 ;
        RECT 3.005 198.345 3.175 199.095 ;
        RECT 3.965 198.345 4.135 199.095 ;
        RECT 4.925 198.345 5.095 199.095 ;
        RECT 5.885 198.345 6.055 199.095 ;
        RECT 2.015 196.985 2.245 198.345 ;
        RECT 2.975 196.985 3.205 198.345 ;
        RECT 3.935 196.985 4.165 198.345 ;
        RECT 4.895 196.985 5.125 198.345 ;
        RECT 5.855 196.985 6.085 198.345 ;
        RECT 0.000 196.110 0.815 196.280 ;
        RECT 0.010 196.105 0.150 196.110 ;
        RECT 0.645 194.225 0.815 196.110 ;
        RECT 2.015 194.925 2.245 195.445 ;
        RECT 2.975 194.925 3.205 195.445 ;
        RECT 3.935 194.925 4.165 195.445 ;
        RECT 4.895 194.925 5.125 195.445 ;
        RECT 5.855 194.925 6.085 195.445 ;
        RECT 2.045 194.225 2.215 194.925 ;
        RECT 3.005 194.225 3.175 194.925 ;
        RECT 3.965 194.225 4.135 194.925 ;
        RECT 4.925 194.225 5.095 194.925 ;
        RECT 5.885 194.225 6.055 194.925 ;
        RECT 0.645 194.055 6.055 194.225 ;
    END
  END in[1]
  PIN in[2]
    DIRECTION INOUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.102000 ;
    PORT
      LAYER li1 ;
        RECT 2.045 190.530 2.215 191.930 ;
        RECT 3.005 190.530 3.175 191.930 ;
        RECT 3.965 190.530 4.135 191.930 ;
        RECT 4.925 190.530 5.095 191.930 ;
        RECT 5.885 190.530 6.055 191.930 ;
        RECT 2.045 188.470 2.215 189.030 ;
        RECT 3.005 188.470 3.175 189.030 ;
        RECT 3.965 188.470 4.135 189.030 ;
        RECT 4.925 188.470 5.095 189.030 ;
        RECT 5.885 188.470 6.055 189.030 ;
      LAYER mcon ;
        RECT 2.045 191.505 2.215 191.675 ;
        RECT 2.045 191.145 2.215 191.315 ;
        RECT 2.045 190.785 2.215 190.955 ;
        RECT 3.005 191.505 3.175 191.675 ;
        RECT 3.005 191.145 3.175 191.315 ;
        RECT 3.005 190.785 3.175 190.955 ;
        RECT 3.965 191.505 4.135 191.675 ;
        RECT 3.965 191.145 4.135 191.315 ;
        RECT 3.965 190.785 4.135 190.955 ;
        RECT 4.925 191.505 5.095 191.675 ;
        RECT 4.925 191.145 5.095 191.315 ;
        RECT 4.925 190.785 5.095 190.955 ;
        RECT 5.885 191.505 6.055 191.675 ;
        RECT 5.885 191.145 6.055 191.315 ;
        RECT 5.885 190.785 6.055 190.955 ;
        RECT 2.045 188.665 2.215 188.835 ;
        RECT 3.005 188.665 3.175 188.835 ;
        RECT 3.965 188.665 4.135 188.835 ;
        RECT 4.925 188.665 5.095 188.835 ;
        RECT 5.885 188.665 6.055 188.835 ;
      LAYER met1 ;
        RECT 0.645 192.660 6.055 192.830 ;
        RECT 0.645 189.845 0.815 192.660 ;
        RECT 2.045 191.910 2.215 192.660 ;
        RECT 3.005 191.910 3.175 192.660 ;
        RECT 3.965 191.910 4.135 192.660 ;
        RECT 4.925 191.910 5.095 192.660 ;
        RECT 5.885 191.910 6.055 192.660 ;
        RECT 2.015 190.550 2.245 191.910 ;
        RECT 2.975 190.550 3.205 191.910 ;
        RECT 3.935 190.550 4.165 191.910 ;
        RECT 4.895 190.550 5.125 191.910 ;
        RECT 5.855 190.550 6.085 191.910 ;
        RECT 0.000 189.675 0.815 189.845 ;
        RECT 0.010 189.670 0.150 189.675 ;
        RECT 0.645 187.790 0.815 189.675 ;
        RECT 2.015 188.490 2.245 189.010 ;
        RECT 2.975 188.490 3.205 189.010 ;
        RECT 3.935 188.490 4.165 189.010 ;
        RECT 4.895 188.490 5.125 189.010 ;
        RECT 5.855 188.490 6.085 189.010 ;
        RECT 2.045 187.790 2.215 188.490 ;
        RECT 3.005 187.790 3.175 188.490 ;
        RECT 3.965 187.790 4.135 188.490 ;
        RECT 4.925 187.790 5.095 188.490 ;
        RECT 5.885 187.790 6.055 188.490 ;
        RECT 0.645 187.620 6.055 187.790 ;
    END
  END in[2]
  PIN in[3]
    DIRECTION INOUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.102000 ;
    PORT
      LAYER li1 ;
        RECT 2.045 184.095 2.215 185.495 ;
        RECT 3.005 184.095 3.175 185.495 ;
        RECT 3.965 184.095 4.135 185.495 ;
        RECT 4.925 184.095 5.095 185.495 ;
        RECT 5.885 184.095 6.055 185.495 ;
        RECT 2.045 182.035 2.215 182.595 ;
        RECT 3.005 182.035 3.175 182.595 ;
        RECT 3.965 182.035 4.135 182.595 ;
        RECT 4.925 182.035 5.095 182.595 ;
        RECT 5.885 182.035 6.055 182.595 ;
      LAYER mcon ;
        RECT 2.045 185.070 2.215 185.240 ;
        RECT 2.045 184.710 2.215 184.880 ;
        RECT 2.045 184.350 2.215 184.520 ;
        RECT 3.005 185.070 3.175 185.240 ;
        RECT 3.005 184.710 3.175 184.880 ;
        RECT 3.005 184.350 3.175 184.520 ;
        RECT 3.965 185.070 4.135 185.240 ;
        RECT 3.965 184.710 4.135 184.880 ;
        RECT 3.965 184.350 4.135 184.520 ;
        RECT 4.925 185.070 5.095 185.240 ;
        RECT 4.925 184.710 5.095 184.880 ;
        RECT 4.925 184.350 5.095 184.520 ;
        RECT 5.885 185.070 6.055 185.240 ;
        RECT 5.885 184.710 6.055 184.880 ;
        RECT 5.885 184.350 6.055 184.520 ;
        RECT 2.045 182.230 2.215 182.400 ;
        RECT 3.005 182.230 3.175 182.400 ;
        RECT 3.965 182.230 4.135 182.400 ;
        RECT 4.925 182.230 5.095 182.400 ;
        RECT 5.885 182.230 6.055 182.400 ;
      LAYER met1 ;
        RECT 0.645 186.225 6.055 186.395 ;
        RECT 0.645 183.410 0.815 186.225 ;
        RECT 2.045 185.475 2.215 186.225 ;
        RECT 3.005 185.475 3.175 186.225 ;
        RECT 3.965 185.475 4.135 186.225 ;
        RECT 4.925 185.475 5.095 186.225 ;
        RECT 5.885 185.475 6.055 186.225 ;
        RECT 2.015 184.115 2.245 185.475 ;
        RECT 2.975 184.115 3.205 185.475 ;
        RECT 3.935 184.115 4.165 185.475 ;
        RECT 4.895 184.115 5.125 185.475 ;
        RECT 5.855 184.115 6.085 185.475 ;
        RECT 0.000 183.240 0.815 183.410 ;
        RECT 0.010 183.235 0.150 183.240 ;
        RECT 0.645 181.355 0.815 183.240 ;
        RECT 2.015 182.055 2.245 182.575 ;
        RECT 2.975 182.055 3.205 182.575 ;
        RECT 3.935 182.055 4.165 182.575 ;
        RECT 4.895 182.055 5.125 182.575 ;
        RECT 5.855 182.055 6.085 182.575 ;
        RECT 2.045 181.355 2.215 182.055 ;
        RECT 3.005 181.355 3.175 182.055 ;
        RECT 3.965 181.355 4.135 182.055 ;
        RECT 4.925 181.355 5.095 182.055 ;
        RECT 5.885 181.355 6.055 182.055 ;
        RECT 0.645 181.185 6.055 181.355 ;
    END
  END in[3]
  PIN in[4]
    DIRECTION INOUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.102000 ;
    PORT
      LAYER li1 ;
        RECT 2.045 177.660 2.215 179.060 ;
        RECT 3.005 177.660 3.175 179.060 ;
        RECT 3.965 177.660 4.135 179.060 ;
        RECT 4.925 177.660 5.095 179.060 ;
        RECT 5.885 177.660 6.055 179.060 ;
        RECT 2.045 175.600 2.215 176.160 ;
        RECT 3.005 175.600 3.175 176.160 ;
        RECT 3.965 175.600 4.135 176.160 ;
        RECT 4.925 175.600 5.095 176.160 ;
        RECT 5.885 175.600 6.055 176.160 ;
      LAYER mcon ;
        RECT 2.045 178.635 2.215 178.805 ;
        RECT 2.045 178.275 2.215 178.445 ;
        RECT 2.045 177.915 2.215 178.085 ;
        RECT 3.005 178.635 3.175 178.805 ;
        RECT 3.005 178.275 3.175 178.445 ;
        RECT 3.005 177.915 3.175 178.085 ;
        RECT 3.965 178.635 4.135 178.805 ;
        RECT 3.965 178.275 4.135 178.445 ;
        RECT 3.965 177.915 4.135 178.085 ;
        RECT 4.925 178.635 5.095 178.805 ;
        RECT 4.925 178.275 5.095 178.445 ;
        RECT 4.925 177.915 5.095 178.085 ;
        RECT 5.885 178.635 6.055 178.805 ;
        RECT 5.885 178.275 6.055 178.445 ;
        RECT 5.885 177.915 6.055 178.085 ;
        RECT 2.045 175.795 2.215 175.965 ;
        RECT 3.005 175.795 3.175 175.965 ;
        RECT 3.965 175.795 4.135 175.965 ;
        RECT 4.925 175.795 5.095 175.965 ;
        RECT 5.885 175.795 6.055 175.965 ;
      LAYER met1 ;
        RECT 0.645 179.790 6.055 179.960 ;
        RECT 0.645 176.975 0.815 179.790 ;
        RECT 2.045 179.040 2.215 179.790 ;
        RECT 3.005 179.040 3.175 179.790 ;
        RECT 3.965 179.040 4.135 179.790 ;
        RECT 4.925 179.040 5.095 179.790 ;
        RECT 5.885 179.040 6.055 179.790 ;
        RECT 2.015 177.680 2.245 179.040 ;
        RECT 2.975 177.680 3.205 179.040 ;
        RECT 3.935 177.680 4.165 179.040 ;
        RECT 4.895 177.680 5.125 179.040 ;
        RECT 5.855 177.680 6.085 179.040 ;
        RECT 0.000 176.805 0.815 176.975 ;
        RECT 0.010 176.800 0.150 176.805 ;
        RECT 0.645 174.920 0.815 176.805 ;
        RECT 2.015 175.620 2.245 176.140 ;
        RECT 2.975 175.620 3.205 176.140 ;
        RECT 3.935 175.620 4.165 176.140 ;
        RECT 4.895 175.620 5.125 176.140 ;
        RECT 5.855 175.620 6.085 176.140 ;
        RECT 2.045 174.920 2.215 175.620 ;
        RECT 3.005 174.920 3.175 175.620 ;
        RECT 3.965 174.920 4.135 175.620 ;
        RECT 4.925 174.920 5.095 175.620 ;
        RECT 5.885 174.920 6.055 175.620 ;
        RECT 0.645 174.750 6.055 174.920 ;
    END
  END in[4]
  PIN in[5]
    DIRECTION INOUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.102000 ;
    PORT
      LAYER li1 ;
        RECT 2.045 171.225 2.215 172.625 ;
        RECT 3.005 171.225 3.175 172.625 ;
        RECT 3.965 171.225 4.135 172.625 ;
        RECT 4.925 171.225 5.095 172.625 ;
        RECT 5.885 171.225 6.055 172.625 ;
        RECT 2.045 169.165 2.215 169.725 ;
        RECT 3.005 169.165 3.175 169.725 ;
        RECT 3.965 169.165 4.135 169.725 ;
        RECT 4.925 169.165 5.095 169.725 ;
        RECT 5.885 169.165 6.055 169.725 ;
      LAYER mcon ;
        RECT 2.045 172.200 2.215 172.370 ;
        RECT 2.045 171.840 2.215 172.010 ;
        RECT 2.045 171.480 2.215 171.650 ;
        RECT 3.005 172.200 3.175 172.370 ;
        RECT 3.005 171.840 3.175 172.010 ;
        RECT 3.005 171.480 3.175 171.650 ;
        RECT 3.965 172.200 4.135 172.370 ;
        RECT 3.965 171.840 4.135 172.010 ;
        RECT 3.965 171.480 4.135 171.650 ;
        RECT 4.925 172.200 5.095 172.370 ;
        RECT 4.925 171.840 5.095 172.010 ;
        RECT 4.925 171.480 5.095 171.650 ;
        RECT 5.885 172.200 6.055 172.370 ;
        RECT 5.885 171.840 6.055 172.010 ;
        RECT 5.885 171.480 6.055 171.650 ;
        RECT 2.045 169.360 2.215 169.530 ;
        RECT 3.005 169.360 3.175 169.530 ;
        RECT 3.965 169.360 4.135 169.530 ;
        RECT 4.925 169.360 5.095 169.530 ;
        RECT 5.885 169.360 6.055 169.530 ;
      LAYER met1 ;
        RECT 0.645 173.355 6.055 173.525 ;
        RECT 0.645 170.540 0.815 173.355 ;
        RECT 2.045 172.605 2.215 173.355 ;
        RECT 3.005 172.605 3.175 173.355 ;
        RECT 3.965 172.605 4.135 173.355 ;
        RECT 4.925 172.605 5.095 173.355 ;
        RECT 5.885 172.605 6.055 173.355 ;
        RECT 2.015 171.245 2.245 172.605 ;
        RECT 2.975 171.245 3.205 172.605 ;
        RECT 3.935 171.245 4.165 172.605 ;
        RECT 4.895 171.245 5.125 172.605 ;
        RECT 5.855 171.245 6.085 172.605 ;
        RECT 0.000 170.370 0.815 170.540 ;
        RECT 0.010 170.365 0.150 170.370 ;
        RECT 0.645 168.485 0.815 170.370 ;
        RECT 2.015 169.185 2.245 169.705 ;
        RECT 2.975 169.185 3.205 169.705 ;
        RECT 3.935 169.185 4.165 169.705 ;
        RECT 4.895 169.185 5.125 169.705 ;
        RECT 5.855 169.185 6.085 169.705 ;
        RECT 2.045 168.485 2.215 169.185 ;
        RECT 3.005 168.485 3.175 169.185 ;
        RECT 3.965 168.485 4.135 169.185 ;
        RECT 4.925 168.485 5.095 169.185 ;
        RECT 5.885 168.485 6.055 169.185 ;
        RECT 0.645 168.315 6.055 168.485 ;
    END
  END in[5]
  PIN in[6]
    DIRECTION INOUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.102000 ;
    PORT
      LAYER li1 ;
        RECT 2.045 164.790 2.215 166.190 ;
        RECT 3.005 164.790 3.175 166.190 ;
        RECT 3.965 164.790 4.135 166.190 ;
        RECT 4.925 164.790 5.095 166.190 ;
        RECT 5.885 164.790 6.055 166.190 ;
        RECT 2.045 162.730 2.215 163.290 ;
        RECT 3.005 162.730 3.175 163.290 ;
        RECT 3.965 162.730 4.135 163.290 ;
        RECT 4.925 162.730 5.095 163.290 ;
        RECT 5.885 162.730 6.055 163.290 ;
      LAYER mcon ;
        RECT 2.045 165.765 2.215 165.935 ;
        RECT 2.045 165.405 2.215 165.575 ;
        RECT 2.045 165.045 2.215 165.215 ;
        RECT 3.005 165.765 3.175 165.935 ;
        RECT 3.005 165.405 3.175 165.575 ;
        RECT 3.005 165.045 3.175 165.215 ;
        RECT 3.965 165.765 4.135 165.935 ;
        RECT 3.965 165.405 4.135 165.575 ;
        RECT 3.965 165.045 4.135 165.215 ;
        RECT 4.925 165.765 5.095 165.935 ;
        RECT 4.925 165.405 5.095 165.575 ;
        RECT 4.925 165.045 5.095 165.215 ;
        RECT 5.885 165.765 6.055 165.935 ;
        RECT 5.885 165.405 6.055 165.575 ;
        RECT 5.885 165.045 6.055 165.215 ;
        RECT 2.045 162.925 2.215 163.095 ;
        RECT 3.005 162.925 3.175 163.095 ;
        RECT 3.965 162.925 4.135 163.095 ;
        RECT 4.925 162.925 5.095 163.095 ;
        RECT 5.885 162.925 6.055 163.095 ;
      LAYER met1 ;
        RECT 0.645 166.920 6.055 167.090 ;
        RECT 0.645 164.105 0.815 166.920 ;
        RECT 2.045 166.170 2.215 166.920 ;
        RECT 3.005 166.170 3.175 166.920 ;
        RECT 3.965 166.170 4.135 166.920 ;
        RECT 4.925 166.170 5.095 166.920 ;
        RECT 5.885 166.170 6.055 166.920 ;
        RECT 2.015 164.810 2.245 166.170 ;
        RECT 2.975 164.810 3.205 166.170 ;
        RECT 3.935 164.810 4.165 166.170 ;
        RECT 4.895 164.810 5.125 166.170 ;
        RECT 5.855 164.810 6.085 166.170 ;
        RECT 0.000 163.935 0.815 164.105 ;
        RECT 0.010 163.930 0.150 163.935 ;
        RECT 0.645 162.050 0.815 163.935 ;
        RECT 2.015 162.750 2.245 163.270 ;
        RECT 2.975 162.750 3.205 163.270 ;
        RECT 3.935 162.750 4.165 163.270 ;
        RECT 4.895 162.750 5.125 163.270 ;
        RECT 5.855 162.750 6.085 163.270 ;
        RECT 2.045 162.050 2.215 162.750 ;
        RECT 3.005 162.050 3.175 162.750 ;
        RECT 3.965 162.050 4.135 162.750 ;
        RECT 4.925 162.050 5.095 162.750 ;
        RECT 5.885 162.050 6.055 162.750 ;
        RECT 0.645 161.880 6.055 162.050 ;
    END
  END in[6]
  PIN in[7]
    DIRECTION INOUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.102000 ;
    PORT
      LAYER li1 ;
        RECT 2.045 158.355 2.215 159.755 ;
        RECT 3.005 158.355 3.175 159.755 ;
        RECT 3.965 158.355 4.135 159.755 ;
        RECT 4.925 158.355 5.095 159.755 ;
        RECT 5.885 158.355 6.055 159.755 ;
        RECT 2.045 156.295 2.215 156.855 ;
        RECT 3.005 156.295 3.175 156.855 ;
        RECT 3.965 156.295 4.135 156.855 ;
        RECT 4.925 156.295 5.095 156.855 ;
        RECT 5.885 156.295 6.055 156.855 ;
      LAYER mcon ;
        RECT 2.045 159.330 2.215 159.500 ;
        RECT 2.045 158.970 2.215 159.140 ;
        RECT 2.045 158.610 2.215 158.780 ;
        RECT 3.005 159.330 3.175 159.500 ;
        RECT 3.005 158.970 3.175 159.140 ;
        RECT 3.005 158.610 3.175 158.780 ;
        RECT 3.965 159.330 4.135 159.500 ;
        RECT 3.965 158.970 4.135 159.140 ;
        RECT 3.965 158.610 4.135 158.780 ;
        RECT 4.925 159.330 5.095 159.500 ;
        RECT 4.925 158.970 5.095 159.140 ;
        RECT 4.925 158.610 5.095 158.780 ;
        RECT 5.885 159.330 6.055 159.500 ;
        RECT 5.885 158.970 6.055 159.140 ;
        RECT 5.885 158.610 6.055 158.780 ;
        RECT 2.045 156.490 2.215 156.660 ;
        RECT 3.005 156.490 3.175 156.660 ;
        RECT 3.965 156.490 4.135 156.660 ;
        RECT 4.925 156.490 5.095 156.660 ;
        RECT 5.885 156.490 6.055 156.660 ;
      LAYER met1 ;
        RECT 0.645 160.485 6.055 160.655 ;
        RECT 0.645 157.670 0.815 160.485 ;
        RECT 2.045 159.735 2.215 160.485 ;
        RECT 3.005 159.735 3.175 160.485 ;
        RECT 3.965 159.735 4.135 160.485 ;
        RECT 4.925 159.735 5.095 160.485 ;
        RECT 5.885 159.735 6.055 160.485 ;
        RECT 2.015 158.375 2.245 159.735 ;
        RECT 2.975 158.375 3.205 159.735 ;
        RECT 3.935 158.375 4.165 159.735 ;
        RECT 4.895 158.375 5.125 159.735 ;
        RECT 5.855 158.375 6.085 159.735 ;
        RECT 0.000 157.500 0.815 157.670 ;
        RECT 0.010 157.495 0.150 157.500 ;
        RECT 0.645 155.615 0.815 157.500 ;
        RECT 2.015 156.315 2.245 156.835 ;
        RECT 2.975 156.315 3.205 156.835 ;
        RECT 3.935 156.315 4.165 156.835 ;
        RECT 4.895 156.315 5.125 156.835 ;
        RECT 5.855 156.315 6.085 156.835 ;
        RECT 2.045 155.615 2.215 156.315 ;
        RECT 3.005 155.615 3.175 156.315 ;
        RECT 3.965 155.615 4.135 156.315 ;
        RECT 4.925 155.615 5.095 156.315 ;
        RECT 5.885 155.615 6.055 156.315 ;
        RECT 0.645 155.445 6.055 155.615 ;
    END
  END in[7]
  PIN in[8]
    DIRECTION INOUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.102000 ;
    PORT
      LAYER li1 ;
        RECT 2.045 151.920 2.215 153.320 ;
        RECT 3.005 151.920 3.175 153.320 ;
        RECT 3.965 151.920 4.135 153.320 ;
        RECT 4.925 151.920 5.095 153.320 ;
        RECT 5.885 151.920 6.055 153.320 ;
        RECT 2.045 149.860 2.215 150.420 ;
        RECT 3.005 149.860 3.175 150.420 ;
        RECT 3.965 149.860 4.135 150.420 ;
        RECT 4.925 149.860 5.095 150.420 ;
        RECT 5.885 149.860 6.055 150.420 ;
      LAYER mcon ;
        RECT 2.045 152.895 2.215 153.065 ;
        RECT 2.045 152.535 2.215 152.705 ;
        RECT 2.045 152.175 2.215 152.345 ;
        RECT 3.005 152.895 3.175 153.065 ;
        RECT 3.005 152.535 3.175 152.705 ;
        RECT 3.005 152.175 3.175 152.345 ;
        RECT 3.965 152.895 4.135 153.065 ;
        RECT 3.965 152.535 4.135 152.705 ;
        RECT 3.965 152.175 4.135 152.345 ;
        RECT 4.925 152.895 5.095 153.065 ;
        RECT 4.925 152.535 5.095 152.705 ;
        RECT 4.925 152.175 5.095 152.345 ;
        RECT 5.885 152.895 6.055 153.065 ;
        RECT 5.885 152.535 6.055 152.705 ;
        RECT 5.885 152.175 6.055 152.345 ;
        RECT 2.045 150.055 2.215 150.225 ;
        RECT 3.005 150.055 3.175 150.225 ;
        RECT 3.965 150.055 4.135 150.225 ;
        RECT 4.925 150.055 5.095 150.225 ;
        RECT 5.885 150.055 6.055 150.225 ;
      LAYER met1 ;
        RECT 0.645 154.050 6.055 154.220 ;
        RECT 0.645 151.235 0.815 154.050 ;
        RECT 2.045 153.300 2.215 154.050 ;
        RECT 3.005 153.300 3.175 154.050 ;
        RECT 3.965 153.300 4.135 154.050 ;
        RECT 4.925 153.300 5.095 154.050 ;
        RECT 5.885 153.300 6.055 154.050 ;
        RECT 2.015 151.940 2.245 153.300 ;
        RECT 2.975 151.940 3.205 153.300 ;
        RECT 3.935 151.940 4.165 153.300 ;
        RECT 4.895 151.940 5.125 153.300 ;
        RECT 5.855 151.940 6.085 153.300 ;
        RECT 0.000 151.065 0.815 151.235 ;
        RECT 0.010 151.060 0.150 151.065 ;
        RECT 0.645 149.180 0.815 151.065 ;
        RECT 2.015 149.880 2.245 150.400 ;
        RECT 2.975 149.880 3.205 150.400 ;
        RECT 3.935 149.880 4.165 150.400 ;
        RECT 4.895 149.880 5.125 150.400 ;
        RECT 5.855 149.880 6.085 150.400 ;
        RECT 2.045 149.180 2.215 149.880 ;
        RECT 3.005 149.180 3.175 149.880 ;
        RECT 3.965 149.180 4.135 149.880 ;
        RECT 4.925 149.180 5.095 149.880 ;
        RECT 5.885 149.180 6.055 149.880 ;
        RECT 0.645 149.010 6.055 149.180 ;
    END
  END in[8]
  PIN in[9]
    DIRECTION INOUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.102000 ;
    PORT
      LAYER li1 ;
        RECT 2.045 145.485 2.215 146.885 ;
        RECT 3.005 145.485 3.175 146.885 ;
        RECT 3.965 145.485 4.135 146.885 ;
        RECT 4.925 145.485 5.095 146.885 ;
        RECT 5.885 145.485 6.055 146.885 ;
        RECT 2.045 143.425 2.215 143.985 ;
        RECT 3.005 143.425 3.175 143.985 ;
        RECT 3.965 143.425 4.135 143.985 ;
        RECT 4.925 143.425 5.095 143.985 ;
        RECT 5.885 143.425 6.055 143.985 ;
      LAYER mcon ;
        RECT 2.045 146.460 2.215 146.630 ;
        RECT 2.045 146.100 2.215 146.270 ;
        RECT 2.045 145.740 2.215 145.910 ;
        RECT 3.005 146.460 3.175 146.630 ;
        RECT 3.005 146.100 3.175 146.270 ;
        RECT 3.005 145.740 3.175 145.910 ;
        RECT 3.965 146.460 4.135 146.630 ;
        RECT 3.965 146.100 4.135 146.270 ;
        RECT 3.965 145.740 4.135 145.910 ;
        RECT 4.925 146.460 5.095 146.630 ;
        RECT 4.925 146.100 5.095 146.270 ;
        RECT 4.925 145.740 5.095 145.910 ;
        RECT 5.885 146.460 6.055 146.630 ;
        RECT 5.885 146.100 6.055 146.270 ;
        RECT 5.885 145.740 6.055 145.910 ;
        RECT 2.045 143.620 2.215 143.790 ;
        RECT 3.005 143.620 3.175 143.790 ;
        RECT 3.965 143.620 4.135 143.790 ;
        RECT 4.925 143.620 5.095 143.790 ;
        RECT 5.885 143.620 6.055 143.790 ;
      LAYER met1 ;
        RECT 0.645 147.615 6.055 147.785 ;
        RECT 0.645 144.800 0.815 147.615 ;
        RECT 2.045 146.865 2.215 147.615 ;
        RECT 3.005 146.865 3.175 147.615 ;
        RECT 3.965 146.865 4.135 147.615 ;
        RECT 4.925 146.865 5.095 147.615 ;
        RECT 5.885 146.865 6.055 147.615 ;
        RECT 2.015 145.505 2.245 146.865 ;
        RECT 2.975 145.505 3.205 146.865 ;
        RECT 3.935 145.505 4.165 146.865 ;
        RECT 4.895 145.505 5.125 146.865 ;
        RECT 5.855 145.505 6.085 146.865 ;
        RECT 0.000 144.630 0.815 144.800 ;
        RECT 0.010 144.625 0.150 144.630 ;
        RECT 0.645 142.745 0.815 144.630 ;
        RECT 2.015 143.445 2.245 143.965 ;
        RECT 2.975 143.445 3.205 143.965 ;
        RECT 3.935 143.445 4.165 143.965 ;
        RECT 4.895 143.445 5.125 143.965 ;
        RECT 5.855 143.445 6.085 143.965 ;
        RECT 2.045 142.745 2.215 143.445 ;
        RECT 3.005 142.745 3.175 143.445 ;
        RECT 3.965 142.745 4.135 143.445 ;
        RECT 4.925 142.745 5.095 143.445 ;
        RECT 5.885 142.745 6.055 143.445 ;
        RECT 0.645 142.575 6.055 142.745 ;
    END
  END in[9]
  PIN in[10]
    DIRECTION INOUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.102000 ;
    PORT
      LAYER li1 ;
        RECT 2.045 139.050 2.215 140.450 ;
        RECT 3.005 139.050 3.175 140.450 ;
        RECT 3.965 139.050 4.135 140.450 ;
        RECT 4.925 139.050 5.095 140.450 ;
        RECT 5.885 139.050 6.055 140.450 ;
        RECT 2.045 136.990 2.215 137.550 ;
        RECT 3.005 136.990 3.175 137.550 ;
        RECT 3.965 136.990 4.135 137.550 ;
        RECT 4.925 136.990 5.095 137.550 ;
        RECT 5.885 136.990 6.055 137.550 ;
      LAYER mcon ;
        RECT 2.045 140.025 2.215 140.195 ;
        RECT 2.045 139.665 2.215 139.835 ;
        RECT 2.045 139.305 2.215 139.475 ;
        RECT 3.005 140.025 3.175 140.195 ;
        RECT 3.005 139.665 3.175 139.835 ;
        RECT 3.005 139.305 3.175 139.475 ;
        RECT 3.965 140.025 4.135 140.195 ;
        RECT 3.965 139.665 4.135 139.835 ;
        RECT 3.965 139.305 4.135 139.475 ;
        RECT 4.925 140.025 5.095 140.195 ;
        RECT 4.925 139.665 5.095 139.835 ;
        RECT 4.925 139.305 5.095 139.475 ;
        RECT 5.885 140.025 6.055 140.195 ;
        RECT 5.885 139.665 6.055 139.835 ;
        RECT 5.885 139.305 6.055 139.475 ;
        RECT 2.045 137.185 2.215 137.355 ;
        RECT 3.005 137.185 3.175 137.355 ;
        RECT 3.965 137.185 4.135 137.355 ;
        RECT 4.925 137.185 5.095 137.355 ;
        RECT 5.885 137.185 6.055 137.355 ;
      LAYER met1 ;
        RECT 0.645 141.180 6.055 141.350 ;
        RECT 0.645 138.365 0.815 141.180 ;
        RECT 2.045 140.430 2.215 141.180 ;
        RECT 3.005 140.430 3.175 141.180 ;
        RECT 3.965 140.430 4.135 141.180 ;
        RECT 4.925 140.430 5.095 141.180 ;
        RECT 5.885 140.430 6.055 141.180 ;
        RECT 2.015 139.070 2.245 140.430 ;
        RECT 2.975 139.070 3.205 140.430 ;
        RECT 3.935 139.070 4.165 140.430 ;
        RECT 4.895 139.070 5.125 140.430 ;
        RECT 5.855 139.070 6.085 140.430 ;
        RECT 0.000 138.195 0.815 138.365 ;
        RECT 0.010 138.190 0.150 138.195 ;
        RECT 0.645 136.310 0.815 138.195 ;
        RECT 2.015 137.010 2.245 137.530 ;
        RECT 2.975 137.010 3.205 137.530 ;
        RECT 3.935 137.010 4.165 137.530 ;
        RECT 4.895 137.010 5.125 137.530 ;
        RECT 5.855 137.010 6.085 137.530 ;
        RECT 2.045 136.310 2.215 137.010 ;
        RECT 3.005 136.310 3.175 137.010 ;
        RECT 3.965 136.310 4.135 137.010 ;
        RECT 4.925 136.310 5.095 137.010 ;
        RECT 5.885 136.310 6.055 137.010 ;
        RECT 0.645 136.140 6.055 136.310 ;
    END
  END in[10]
  PIN in[11]
    DIRECTION INOUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.102000 ;
    PORT
      LAYER li1 ;
        RECT 2.045 132.615 2.215 134.015 ;
        RECT 3.005 132.615 3.175 134.015 ;
        RECT 3.965 132.615 4.135 134.015 ;
        RECT 4.925 132.615 5.095 134.015 ;
        RECT 5.885 132.615 6.055 134.015 ;
        RECT 2.045 130.555 2.215 131.115 ;
        RECT 3.005 130.555 3.175 131.115 ;
        RECT 3.965 130.555 4.135 131.115 ;
        RECT 4.925 130.555 5.095 131.115 ;
        RECT 5.885 130.555 6.055 131.115 ;
      LAYER mcon ;
        RECT 2.045 133.590 2.215 133.760 ;
        RECT 2.045 133.230 2.215 133.400 ;
        RECT 2.045 132.870 2.215 133.040 ;
        RECT 3.005 133.590 3.175 133.760 ;
        RECT 3.005 133.230 3.175 133.400 ;
        RECT 3.005 132.870 3.175 133.040 ;
        RECT 3.965 133.590 4.135 133.760 ;
        RECT 3.965 133.230 4.135 133.400 ;
        RECT 3.965 132.870 4.135 133.040 ;
        RECT 4.925 133.590 5.095 133.760 ;
        RECT 4.925 133.230 5.095 133.400 ;
        RECT 4.925 132.870 5.095 133.040 ;
        RECT 5.885 133.590 6.055 133.760 ;
        RECT 5.885 133.230 6.055 133.400 ;
        RECT 5.885 132.870 6.055 133.040 ;
        RECT 2.045 130.750 2.215 130.920 ;
        RECT 3.005 130.750 3.175 130.920 ;
        RECT 3.965 130.750 4.135 130.920 ;
        RECT 4.925 130.750 5.095 130.920 ;
        RECT 5.885 130.750 6.055 130.920 ;
      LAYER met1 ;
        RECT 0.645 134.745 6.055 134.915 ;
        RECT 0.645 131.930 0.815 134.745 ;
        RECT 2.045 133.995 2.215 134.745 ;
        RECT 3.005 133.995 3.175 134.745 ;
        RECT 3.965 133.995 4.135 134.745 ;
        RECT 4.925 133.995 5.095 134.745 ;
        RECT 5.885 133.995 6.055 134.745 ;
        RECT 2.015 132.635 2.245 133.995 ;
        RECT 2.975 132.635 3.205 133.995 ;
        RECT 3.935 132.635 4.165 133.995 ;
        RECT 4.895 132.635 5.125 133.995 ;
        RECT 5.855 132.635 6.085 133.995 ;
        RECT 0.000 131.760 0.815 131.930 ;
        RECT 0.010 131.755 0.150 131.760 ;
        RECT 0.645 129.875 0.815 131.760 ;
        RECT 2.015 130.575 2.245 131.095 ;
        RECT 2.975 130.575 3.205 131.095 ;
        RECT 3.935 130.575 4.165 131.095 ;
        RECT 4.895 130.575 5.125 131.095 ;
        RECT 5.855 130.575 6.085 131.095 ;
        RECT 2.045 129.875 2.215 130.575 ;
        RECT 3.005 129.875 3.175 130.575 ;
        RECT 3.965 129.875 4.135 130.575 ;
        RECT 4.925 129.875 5.095 130.575 ;
        RECT 5.885 129.875 6.055 130.575 ;
        RECT 0.645 129.705 6.055 129.875 ;
    END
  END in[11]
  PIN in[12]
    DIRECTION INOUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.102000 ;
    PORT
      LAYER li1 ;
        RECT 2.045 126.180 2.215 127.580 ;
        RECT 3.005 126.180 3.175 127.580 ;
        RECT 3.965 126.180 4.135 127.580 ;
        RECT 4.925 126.180 5.095 127.580 ;
        RECT 5.885 126.180 6.055 127.580 ;
        RECT 2.045 124.120 2.215 124.680 ;
        RECT 3.005 124.120 3.175 124.680 ;
        RECT 3.965 124.120 4.135 124.680 ;
        RECT 4.925 124.120 5.095 124.680 ;
        RECT 5.885 124.120 6.055 124.680 ;
      LAYER mcon ;
        RECT 2.045 127.155 2.215 127.325 ;
        RECT 2.045 126.795 2.215 126.965 ;
        RECT 2.045 126.435 2.215 126.605 ;
        RECT 3.005 127.155 3.175 127.325 ;
        RECT 3.005 126.795 3.175 126.965 ;
        RECT 3.005 126.435 3.175 126.605 ;
        RECT 3.965 127.155 4.135 127.325 ;
        RECT 3.965 126.795 4.135 126.965 ;
        RECT 3.965 126.435 4.135 126.605 ;
        RECT 4.925 127.155 5.095 127.325 ;
        RECT 4.925 126.795 5.095 126.965 ;
        RECT 4.925 126.435 5.095 126.605 ;
        RECT 5.885 127.155 6.055 127.325 ;
        RECT 5.885 126.795 6.055 126.965 ;
        RECT 5.885 126.435 6.055 126.605 ;
        RECT 2.045 124.315 2.215 124.485 ;
        RECT 3.005 124.315 3.175 124.485 ;
        RECT 3.965 124.315 4.135 124.485 ;
        RECT 4.925 124.315 5.095 124.485 ;
        RECT 5.885 124.315 6.055 124.485 ;
      LAYER met1 ;
        RECT 0.645 128.310 6.055 128.480 ;
        RECT 0.645 125.495 0.815 128.310 ;
        RECT 2.045 127.560 2.215 128.310 ;
        RECT 3.005 127.560 3.175 128.310 ;
        RECT 3.965 127.560 4.135 128.310 ;
        RECT 4.925 127.560 5.095 128.310 ;
        RECT 5.885 127.560 6.055 128.310 ;
        RECT 2.015 126.200 2.245 127.560 ;
        RECT 2.975 126.200 3.205 127.560 ;
        RECT 3.935 126.200 4.165 127.560 ;
        RECT 4.895 126.200 5.125 127.560 ;
        RECT 5.855 126.200 6.085 127.560 ;
        RECT 0.000 125.325 0.815 125.495 ;
        RECT 0.010 125.320 0.150 125.325 ;
        RECT 0.645 123.440 0.815 125.325 ;
        RECT 2.015 124.140 2.245 124.660 ;
        RECT 2.975 124.140 3.205 124.660 ;
        RECT 3.935 124.140 4.165 124.660 ;
        RECT 4.895 124.140 5.125 124.660 ;
        RECT 5.855 124.140 6.085 124.660 ;
        RECT 2.045 123.440 2.215 124.140 ;
        RECT 3.005 123.440 3.175 124.140 ;
        RECT 3.965 123.440 4.135 124.140 ;
        RECT 4.925 123.440 5.095 124.140 ;
        RECT 5.885 123.440 6.055 124.140 ;
        RECT 0.645 123.270 6.055 123.440 ;
    END
  END in[12]
  PIN in[13]
    DIRECTION INOUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.102000 ;
    PORT
      LAYER li1 ;
        RECT 2.045 119.745 2.215 121.145 ;
        RECT 3.005 119.745 3.175 121.145 ;
        RECT 3.965 119.745 4.135 121.145 ;
        RECT 4.925 119.745 5.095 121.145 ;
        RECT 5.885 119.745 6.055 121.145 ;
        RECT 2.045 117.685 2.215 118.245 ;
        RECT 3.005 117.685 3.175 118.245 ;
        RECT 3.965 117.685 4.135 118.245 ;
        RECT 4.925 117.685 5.095 118.245 ;
        RECT 5.885 117.685 6.055 118.245 ;
      LAYER mcon ;
        RECT 2.045 120.720 2.215 120.890 ;
        RECT 2.045 120.360 2.215 120.530 ;
        RECT 2.045 120.000 2.215 120.170 ;
        RECT 3.005 120.720 3.175 120.890 ;
        RECT 3.005 120.360 3.175 120.530 ;
        RECT 3.005 120.000 3.175 120.170 ;
        RECT 3.965 120.720 4.135 120.890 ;
        RECT 3.965 120.360 4.135 120.530 ;
        RECT 3.965 120.000 4.135 120.170 ;
        RECT 4.925 120.720 5.095 120.890 ;
        RECT 4.925 120.360 5.095 120.530 ;
        RECT 4.925 120.000 5.095 120.170 ;
        RECT 5.885 120.720 6.055 120.890 ;
        RECT 5.885 120.360 6.055 120.530 ;
        RECT 5.885 120.000 6.055 120.170 ;
        RECT 2.045 117.880 2.215 118.050 ;
        RECT 3.005 117.880 3.175 118.050 ;
        RECT 3.965 117.880 4.135 118.050 ;
        RECT 4.925 117.880 5.095 118.050 ;
        RECT 5.885 117.880 6.055 118.050 ;
      LAYER met1 ;
        RECT 0.645 121.875 6.055 122.045 ;
        RECT 0.645 119.060 0.815 121.875 ;
        RECT 2.045 121.125 2.215 121.875 ;
        RECT 3.005 121.125 3.175 121.875 ;
        RECT 3.965 121.125 4.135 121.875 ;
        RECT 4.925 121.125 5.095 121.875 ;
        RECT 5.885 121.125 6.055 121.875 ;
        RECT 2.015 119.765 2.245 121.125 ;
        RECT 2.975 119.765 3.205 121.125 ;
        RECT 3.935 119.765 4.165 121.125 ;
        RECT 4.895 119.765 5.125 121.125 ;
        RECT 5.855 119.765 6.085 121.125 ;
        RECT 0.000 118.890 0.815 119.060 ;
        RECT 0.010 118.885 0.150 118.890 ;
        RECT 0.645 117.005 0.815 118.890 ;
        RECT 2.015 117.705 2.245 118.225 ;
        RECT 2.975 117.705 3.205 118.225 ;
        RECT 3.935 117.705 4.165 118.225 ;
        RECT 4.895 117.705 5.125 118.225 ;
        RECT 5.855 117.705 6.085 118.225 ;
        RECT 2.045 117.005 2.215 117.705 ;
        RECT 3.005 117.005 3.175 117.705 ;
        RECT 3.965 117.005 4.135 117.705 ;
        RECT 4.925 117.005 5.095 117.705 ;
        RECT 5.885 117.005 6.055 117.705 ;
        RECT 0.645 116.835 6.055 117.005 ;
    END
  END in[13]
  PIN in[14]
    DIRECTION INOUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.102000 ;
    PORT
      LAYER li1 ;
        RECT 2.045 113.310 2.215 114.710 ;
        RECT 3.005 113.310 3.175 114.710 ;
        RECT 3.965 113.310 4.135 114.710 ;
        RECT 4.925 113.310 5.095 114.710 ;
        RECT 5.885 113.310 6.055 114.710 ;
        RECT 2.045 111.250 2.215 111.810 ;
        RECT 3.005 111.250 3.175 111.810 ;
        RECT 3.965 111.250 4.135 111.810 ;
        RECT 4.925 111.250 5.095 111.810 ;
        RECT 5.885 111.250 6.055 111.810 ;
      LAYER mcon ;
        RECT 2.045 114.285 2.215 114.455 ;
        RECT 2.045 113.925 2.215 114.095 ;
        RECT 2.045 113.565 2.215 113.735 ;
        RECT 3.005 114.285 3.175 114.455 ;
        RECT 3.005 113.925 3.175 114.095 ;
        RECT 3.005 113.565 3.175 113.735 ;
        RECT 3.965 114.285 4.135 114.455 ;
        RECT 3.965 113.925 4.135 114.095 ;
        RECT 3.965 113.565 4.135 113.735 ;
        RECT 4.925 114.285 5.095 114.455 ;
        RECT 4.925 113.925 5.095 114.095 ;
        RECT 4.925 113.565 5.095 113.735 ;
        RECT 5.885 114.285 6.055 114.455 ;
        RECT 5.885 113.925 6.055 114.095 ;
        RECT 5.885 113.565 6.055 113.735 ;
        RECT 2.045 111.445 2.215 111.615 ;
        RECT 3.005 111.445 3.175 111.615 ;
        RECT 3.965 111.445 4.135 111.615 ;
        RECT 4.925 111.445 5.095 111.615 ;
        RECT 5.885 111.445 6.055 111.615 ;
      LAYER met1 ;
        RECT 0.645 115.440 6.055 115.610 ;
        RECT 0.645 112.625 0.815 115.440 ;
        RECT 2.045 114.690 2.215 115.440 ;
        RECT 3.005 114.690 3.175 115.440 ;
        RECT 3.965 114.690 4.135 115.440 ;
        RECT 4.925 114.690 5.095 115.440 ;
        RECT 5.885 114.690 6.055 115.440 ;
        RECT 2.015 113.330 2.245 114.690 ;
        RECT 2.975 113.330 3.205 114.690 ;
        RECT 3.935 113.330 4.165 114.690 ;
        RECT 4.895 113.330 5.125 114.690 ;
        RECT 5.855 113.330 6.085 114.690 ;
        RECT 0.000 112.455 0.815 112.625 ;
        RECT 0.010 112.450 0.150 112.455 ;
        RECT 0.645 110.570 0.815 112.455 ;
        RECT 2.015 111.270 2.245 111.790 ;
        RECT 2.975 111.270 3.205 111.790 ;
        RECT 3.935 111.270 4.165 111.790 ;
        RECT 4.895 111.270 5.125 111.790 ;
        RECT 5.855 111.270 6.085 111.790 ;
        RECT 2.045 110.570 2.215 111.270 ;
        RECT 3.005 110.570 3.175 111.270 ;
        RECT 3.965 110.570 4.135 111.270 ;
        RECT 4.925 110.570 5.095 111.270 ;
        RECT 5.885 110.570 6.055 111.270 ;
        RECT 0.645 110.400 6.055 110.570 ;
    END
  END in[14]
  PIN in[15]
    DIRECTION INOUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.102000 ;
    PORT
      LAYER li1 ;
        RECT 2.045 106.875 2.215 108.275 ;
        RECT 3.005 106.875 3.175 108.275 ;
        RECT 3.965 106.875 4.135 108.275 ;
        RECT 4.925 106.875 5.095 108.275 ;
        RECT 5.885 106.875 6.055 108.275 ;
        RECT 2.045 104.815 2.215 105.375 ;
        RECT 3.005 104.815 3.175 105.375 ;
        RECT 3.965 104.815 4.135 105.375 ;
        RECT 4.925 104.815 5.095 105.375 ;
        RECT 5.885 104.815 6.055 105.375 ;
      LAYER mcon ;
        RECT 2.045 107.850 2.215 108.020 ;
        RECT 2.045 107.490 2.215 107.660 ;
        RECT 2.045 107.130 2.215 107.300 ;
        RECT 3.005 107.850 3.175 108.020 ;
        RECT 3.005 107.490 3.175 107.660 ;
        RECT 3.005 107.130 3.175 107.300 ;
        RECT 3.965 107.850 4.135 108.020 ;
        RECT 3.965 107.490 4.135 107.660 ;
        RECT 3.965 107.130 4.135 107.300 ;
        RECT 4.925 107.850 5.095 108.020 ;
        RECT 4.925 107.490 5.095 107.660 ;
        RECT 4.925 107.130 5.095 107.300 ;
        RECT 5.885 107.850 6.055 108.020 ;
        RECT 5.885 107.490 6.055 107.660 ;
        RECT 5.885 107.130 6.055 107.300 ;
        RECT 2.045 105.010 2.215 105.180 ;
        RECT 3.005 105.010 3.175 105.180 ;
        RECT 3.965 105.010 4.135 105.180 ;
        RECT 4.925 105.010 5.095 105.180 ;
        RECT 5.885 105.010 6.055 105.180 ;
      LAYER met1 ;
        RECT 0.645 109.005 6.055 109.175 ;
        RECT 0.645 106.190 0.815 109.005 ;
        RECT 2.045 108.255 2.215 109.005 ;
        RECT 3.005 108.255 3.175 109.005 ;
        RECT 3.965 108.255 4.135 109.005 ;
        RECT 4.925 108.255 5.095 109.005 ;
        RECT 5.885 108.255 6.055 109.005 ;
        RECT 2.015 106.895 2.245 108.255 ;
        RECT 2.975 106.895 3.205 108.255 ;
        RECT 3.935 106.895 4.165 108.255 ;
        RECT 4.895 106.895 5.125 108.255 ;
        RECT 5.855 106.895 6.085 108.255 ;
        RECT 0.000 106.020 0.815 106.190 ;
        RECT 0.010 106.015 0.150 106.020 ;
        RECT 0.645 104.135 0.815 106.020 ;
        RECT 2.015 104.835 2.245 105.355 ;
        RECT 2.975 104.835 3.205 105.355 ;
        RECT 3.935 104.835 4.165 105.355 ;
        RECT 4.895 104.835 5.125 105.355 ;
        RECT 5.855 104.835 6.085 105.355 ;
        RECT 2.045 104.135 2.215 104.835 ;
        RECT 3.005 104.135 3.175 104.835 ;
        RECT 3.965 104.135 4.135 104.835 ;
        RECT 4.925 104.135 5.095 104.835 ;
        RECT 5.885 104.135 6.055 104.835 ;
        RECT 0.645 103.965 6.055 104.135 ;
    END
  END in[15]
  PIN in[16]
    DIRECTION INOUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.102000 ;
    PORT
      LAYER li1 ;
        RECT 2.045 100.440 2.215 101.840 ;
        RECT 3.005 100.440 3.175 101.840 ;
        RECT 3.965 100.440 4.135 101.840 ;
        RECT 4.925 100.440 5.095 101.840 ;
        RECT 5.885 100.440 6.055 101.840 ;
        RECT 2.045 98.380 2.215 98.940 ;
        RECT 3.005 98.380 3.175 98.940 ;
        RECT 3.965 98.380 4.135 98.940 ;
        RECT 4.925 98.380 5.095 98.940 ;
        RECT 5.885 98.380 6.055 98.940 ;
      LAYER mcon ;
        RECT 2.045 101.415 2.215 101.585 ;
        RECT 2.045 101.055 2.215 101.225 ;
        RECT 2.045 100.695 2.215 100.865 ;
        RECT 3.005 101.415 3.175 101.585 ;
        RECT 3.005 101.055 3.175 101.225 ;
        RECT 3.005 100.695 3.175 100.865 ;
        RECT 3.965 101.415 4.135 101.585 ;
        RECT 3.965 101.055 4.135 101.225 ;
        RECT 3.965 100.695 4.135 100.865 ;
        RECT 4.925 101.415 5.095 101.585 ;
        RECT 4.925 101.055 5.095 101.225 ;
        RECT 4.925 100.695 5.095 100.865 ;
        RECT 5.885 101.415 6.055 101.585 ;
        RECT 5.885 101.055 6.055 101.225 ;
        RECT 5.885 100.695 6.055 100.865 ;
        RECT 2.045 98.575 2.215 98.745 ;
        RECT 3.005 98.575 3.175 98.745 ;
        RECT 3.965 98.575 4.135 98.745 ;
        RECT 4.925 98.575 5.095 98.745 ;
        RECT 5.885 98.575 6.055 98.745 ;
      LAYER met1 ;
        RECT 0.645 102.570 6.055 102.740 ;
        RECT 0.645 99.755 0.815 102.570 ;
        RECT 2.045 101.820 2.215 102.570 ;
        RECT 3.005 101.820 3.175 102.570 ;
        RECT 3.965 101.820 4.135 102.570 ;
        RECT 4.925 101.820 5.095 102.570 ;
        RECT 5.885 101.820 6.055 102.570 ;
        RECT 2.015 100.460 2.245 101.820 ;
        RECT 2.975 100.460 3.205 101.820 ;
        RECT 3.935 100.460 4.165 101.820 ;
        RECT 4.895 100.460 5.125 101.820 ;
        RECT 5.855 100.460 6.085 101.820 ;
        RECT 0.000 99.585 0.815 99.755 ;
        RECT 0.010 99.580 0.150 99.585 ;
        RECT 0.645 97.700 0.815 99.585 ;
        RECT 2.015 98.400 2.245 98.920 ;
        RECT 2.975 98.400 3.205 98.920 ;
        RECT 3.935 98.400 4.165 98.920 ;
        RECT 4.895 98.400 5.125 98.920 ;
        RECT 5.855 98.400 6.085 98.920 ;
        RECT 2.045 97.700 2.215 98.400 ;
        RECT 3.005 97.700 3.175 98.400 ;
        RECT 3.965 97.700 4.135 98.400 ;
        RECT 4.925 97.700 5.095 98.400 ;
        RECT 5.885 97.700 6.055 98.400 ;
        RECT 0.645 97.530 6.055 97.700 ;
    END
  END in[16]
  PIN in[17]
    DIRECTION INOUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.102000 ;
    PORT
      LAYER li1 ;
        RECT 2.045 94.005 2.215 95.405 ;
        RECT 3.005 94.005 3.175 95.405 ;
        RECT 3.965 94.005 4.135 95.405 ;
        RECT 4.925 94.005 5.095 95.405 ;
        RECT 5.885 94.005 6.055 95.405 ;
        RECT 2.045 91.945 2.215 92.505 ;
        RECT 3.005 91.945 3.175 92.505 ;
        RECT 3.965 91.945 4.135 92.505 ;
        RECT 4.925 91.945 5.095 92.505 ;
        RECT 5.885 91.945 6.055 92.505 ;
      LAYER mcon ;
        RECT 2.045 94.980 2.215 95.150 ;
        RECT 2.045 94.620 2.215 94.790 ;
        RECT 2.045 94.260 2.215 94.430 ;
        RECT 3.005 94.980 3.175 95.150 ;
        RECT 3.005 94.620 3.175 94.790 ;
        RECT 3.005 94.260 3.175 94.430 ;
        RECT 3.965 94.980 4.135 95.150 ;
        RECT 3.965 94.620 4.135 94.790 ;
        RECT 3.965 94.260 4.135 94.430 ;
        RECT 4.925 94.980 5.095 95.150 ;
        RECT 4.925 94.620 5.095 94.790 ;
        RECT 4.925 94.260 5.095 94.430 ;
        RECT 5.885 94.980 6.055 95.150 ;
        RECT 5.885 94.620 6.055 94.790 ;
        RECT 5.885 94.260 6.055 94.430 ;
        RECT 2.045 92.140 2.215 92.310 ;
        RECT 3.005 92.140 3.175 92.310 ;
        RECT 3.965 92.140 4.135 92.310 ;
        RECT 4.925 92.140 5.095 92.310 ;
        RECT 5.885 92.140 6.055 92.310 ;
      LAYER met1 ;
        RECT 0.645 96.135 6.055 96.305 ;
        RECT 0.645 93.320 0.815 96.135 ;
        RECT 2.045 95.385 2.215 96.135 ;
        RECT 3.005 95.385 3.175 96.135 ;
        RECT 3.965 95.385 4.135 96.135 ;
        RECT 4.925 95.385 5.095 96.135 ;
        RECT 5.885 95.385 6.055 96.135 ;
        RECT 2.015 94.025 2.245 95.385 ;
        RECT 2.975 94.025 3.205 95.385 ;
        RECT 3.935 94.025 4.165 95.385 ;
        RECT 4.895 94.025 5.125 95.385 ;
        RECT 5.855 94.025 6.085 95.385 ;
        RECT 0.000 93.150 0.815 93.320 ;
        RECT 0.010 93.145 0.150 93.150 ;
        RECT 0.645 91.265 0.815 93.150 ;
        RECT 2.015 91.965 2.245 92.485 ;
        RECT 2.975 91.965 3.205 92.485 ;
        RECT 3.935 91.965 4.165 92.485 ;
        RECT 4.895 91.965 5.125 92.485 ;
        RECT 5.855 91.965 6.085 92.485 ;
        RECT 2.045 91.265 2.215 91.965 ;
        RECT 3.005 91.265 3.175 91.965 ;
        RECT 3.965 91.265 4.135 91.965 ;
        RECT 4.925 91.265 5.095 91.965 ;
        RECT 5.885 91.265 6.055 91.965 ;
        RECT 0.645 91.095 6.055 91.265 ;
    END
  END in[17]
  PIN in[18]
    DIRECTION INOUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.102000 ;
    PORT
      LAYER li1 ;
        RECT 2.045 87.570 2.215 88.970 ;
        RECT 3.005 87.570 3.175 88.970 ;
        RECT 3.965 87.570 4.135 88.970 ;
        RECT 4.925 87.570 5.095 88.970 ;
        RECT 5.885 87.570 6.055 88.970 ;
        RECT 2.045 85.510 2.215 86.070 ;
        RECT 3.005 85.510 3.175 86.070 ;
        RECT 3.965 85.510 4.135 86.070 ;
        RECT 4.925 85.510 5.095 86.070 ;
        RECT 5.885 85.510 6.055 86.070 ;
      LAYER mcon ;
        RECT 2.045 88.545 2.215 88.715 ;
        RECT 2.045 88.185 2.215 88.355 ;
        RECT 2.045 87.825 2.215 87.995 ;
        RECT 3.005 88.545 3.175 88.715 ;
        RECT 3.005 88.185 3.175 88.355 ;
        RECT 3.005 87.825 3.175 87.995 ;
        RECT 3.965 88.545 4.135 88.715 ;
        RECT 3.965 88.185 4.135 88.355 ;
        RECT 3.965 87.825 4.135 87.995 ;
        RECT 4.925 88.545 5.095 88.715 ;
        RECT 4.925 88.185 5.095 88.355 ;
        RECT 4.925 87.825 5.095 87.995 ;
        RECT 5.885 88.545 6.055 88.715 ;
        RECT 5.885 88.185 6.055 88.355 ;
        RECT 5.885 87.825 6.055 87.995 ;
        RECT 2.045 85.705 2.215 85.875 ;
        RECT 3.005 85.705 3.175 85.875 ;
        RECT 3.965 85.705 4.135 85.875 ;
        RECT 4.925 85.705 5.095 85.875 ;
        RECT 5.885 85.705 6.055 85.875 ;
      LAYER met1 ;
        RECT 0.645 89.700 6.055 89.870 ;
        RECT 0.645 86.885 0.815 89.700 ;
        RECT 2.045 88.950 2.215 89.700 ;
        RECT 3.005 88.950 3.175 89.700 ;
        RECT 3.965 88.950 4.135 89.700 ;
        RECT 4.925 88.950 5.095 89.700 ;
        RECT 5.885 88.950 6.055 89.700 ;
        RECT 2.015 87.590 2.245 88.950 ;
        RECT 2.975 87.590 3.205 88.950 ;
        RECT 3.935 87.590 4.165 88.950 ;
        RECT 4.895 87.590 5.125 88.950 ;
        RECT 5.855 87.590 6.085 88.950 ;
        RECT 0.000 86.715 0.815 86.885 ;
        RECT 0.010 86.710 0.150 86.715 ;
        RECT 0.645 84.830 0.815 86.715 ;
        RECT 2.015 85.530 2.245 86.050 ;
        RECT 2.975 85.530 3.205 86.050 ;
        RECT 3.935 85.530 4.165 86.050 ;
        RECT 4.895 85.530 5.125 86.050 ;
        RECT 5.855 85.530 6.085 86.050 ;
        RECT 2.045 84.830 2.215 85.530 ;
        RECT 3.005 84.830 3.175 85.530 ;
        RECT 3.965 84.830 4.135 85.530 ;
        RECT 4.925 84.830 5.095 85.530 ;
        RECT 5.885 84.830 6.055 85.530 ;
        RECT 0.645 84.660 6.055 84.830 ;
    END
  END in[18]
  PIN in[19]
    DIRECTION INOUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.102000 ;
    PORT
      LAYER li1 ;
        RECT 2.045 81.135 2.215 82.535 ;
        RECT 3.005 81.135 3.175 82.535 ;
        RECT 3.965 81.135 4.135 82.535 ;
        RECT 4.925 81.135 5.095 82.535 ;
        RECT 5.885 81.135 6.055 82.535 ;
        RECT 2.045 79.075 2.215 79.635 ;
        RECT 3.005 79.075 3.175 79.635 ;
        RECT 3.965 79.075 4.135 79.635 ;
        RECT 4.925 79.075 5.095 79.635 ;
        RECT 5.885 79.075 6.055 79.635 ;
      LAYER mcon ;
        RECT 2.045 82.110 2.215 82.280 ;
        RECT 2.045 81.750 2.215 81.920 ;
        RECT 2.045 81.390 2.215 81.560 ;
        RECT 3.005 82.110 3.175 82.280 ;
        RECT 3.005 81.750 3.175 81.920 ;
        RECT 3.005 81.390 3.175 81.560 ;
        RECT 3.965 82.110 4.135 82.280 ;
        RECT 3.965 81.750 4.135 81.920 ;
        RECT 3.965 81.390 4.135 81.560 ;
        RECT 4.925 82.110 5.095 82.280 ;
        RECT 4.925 81.750 5.095 81.920 ;
        RECT 4.925 81.390 5.095 81.560 ;
        RECT 5.885 82.110 6.055 82.280 ;
        RECT 5.885 81.750 6.055 81.920 ;
        RECT 5.885 81.390 6.055 81.560 ;
        RECT 2.045 79.270 2.215 79.440 ;
        RECT 3.005 79.270 3.175 79.440 ;
        RECT 3.965 79.270 4.135 79.440 ;
        RECT 4.925 79.270 5.095 79.440 ;
        RECT 5.885 79.270 6.055 79.440 ;
      LAYER met1 ;
        RECT 0.645 83.265 6.055 83.435 ;
        RECT 0.645 80.450 0.815 83.265 ;
        RECT 2.045 82.515 2.215 83.265 ;
        RECT 3.005 82.515 3.175 83.265 ;
        RECT 3.965 82.515 4.135 83.265 ;
        RECT 4.925 82.515 5.095 83.265 ;
        RECT 5.885 82.515 6.055 83.265 ;
        RECT 2.015 81.155 2.245 82.515 ;
        RECT 2.975 81.155 3.205 82.515 ;
        RECT 3.935 81.155 4.165 82.515 ;
        RECT 4.895 81.155 5.125 82.515 ;
        RECT 5.855 81.155 6.085 82.515 ;
        RECT 0.000 80.280 0.815 80.450 ;
        RECT 0.010 80.275 0.150 80.280 ;
        RECT 0.645 78.395 0.815 80.280 ;
        RECT 2.015 79.095 2.245 79.615 ;
        RECT 2.975 79.095 3.205 79.615 ;
        RECT 3.935 79.095 4.165 79.615 ;
        RECT 4.895 79.095 5.125 79.615 ;
        RECT 5.855 79.095 6.085 79.615 ;
        RECT 2.045 78.395 2.215 79.095 ;
        RECT 3.005 78.395 3.175 79.095 ;
        RECT 3.965 78.395 4.135 79.095 ;
        RECT 4.925 78.395 5.095 79.095 ;
        RECT 5.885 78.395 6.055 79.095 ;
        RECT 0.645 78.225 6.055 78.395 ;
    END
  END in[19]
  PIN in[20]
    DIRECTION INOUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.102000 ;
    PORT
      LAYER li1 ;
        RECT 2.045 74.700 2.215 76.100 ;
        RECT 3.005 74.700 3.175 76.100 ;
        RECT 3.965 74.700 4.135 76.100 ;
        RECT 4.925 74.700 5.095 76.100 ;
        RECT 5.885 74.700 6.055 76.100 ;
        RECT 2.045 72.640 2.215 73.200 ;
        RECT 3.005 72.640 3.175 73.200 ;
        RECT 3.965 72.640 4.135 73.200 ;
        RECT 4.925 72.640 5.095 73.200 ;
        RECT 5.885 72.640 6.055 73.200 ;
      LAYER mcon ;
        RECT 2.045 75.675 2.215 75.845 ;
        RECT 2.045 75.315 2.215 75.485 ;
        RECT 2.045 74.955 2.215 75.125 ;
        RECT 3.005 75.675 3.175 75.845 ;
        RECT 3.005 75.315 3.175 75.485 ;
        RECT 3.005 74.955 3.175 75.125 ;
        RECT 3.965 75.675 4.135 75.845 ;
        RECT 3.965 75.315 4.135 75.485 ;
        RECT 3.965 74.955 4.135 75.125 ;
        RECT 4.925 75.675 5.095 75.845 ;
        RECT 4.925 75.315 5.095 75.485 ;
        RECT 4.925 74.955 5.095 75.125 ;
        RECT 5.885 75.675 6.055 75.845 ;
        RECT 5.885 75.315 6.055 75.485 ;
        RECT 5.885 74.955 6.055 75.125 ;
        RECT 2.045 72.835 2.215 73.005 ;
        RECT 3.005 72.835 3.175 73.005 ;
        RECT 3.965 72.835 4.135 73.005 ;
        RECT 4.925 72.835 5.095 73.005 ;
        RECT 5.885 72.835 6.055 73.005 ;
      LAYER met1 ;
        RECT 0.645 76.830 6.055 77.000 ;
        RECT 0.645 74.015 0.815 76.830 ;
        RECT 2.045 76.080 2.215 76.830 ;
        RECT 3.005 76.080 3.175 76.830 ;
        RECT 3.965 76.080 4.135 76.830 ;
        RECT 4.925 76.080 5.095 76.830 ;
        RECT 5.885 76.080 6.055 76.830 ;
        RECT 2.015 74.720 2.245 76.080 ;
        RECT 2.975 74.720 3.205 76.080 ;
        RECT 3.935 74.720 4.165 76.080 ;
        RECT 4.895 74.720 5.125 76.080 ;
        RECT 5.855 74.720 6.085 76.080 ;
        RECT 0.000 73.845 0.815 74.015 ;
        RECT 0.010 73.840 0.150 73.845 ;
        RECT 0.645 71.960 0.815 73.845 ;
        RECT 2.015 72.660 2.245 73.180 ;
        RECT 2.975 72.660 3.205 73.180 ;
        RECT 3.935 72.660 4.165 73.180 ;
        RECT 4.895 72.660 5.125 73.180 ;
        RECT 5.855 72.660 6.085 73.180 ;
        RECT 2.045 71.960 2.215 72.660 ;
        RECT 3.005 71.960 3.175 72.660 ;
        RECT 3.965 71.960 4.135 72.660 ;
        RECT 4.925 71.960 5.095 72.660 ;
        RECT 5.885 71.960 6.055 72.660 ;
        RECT 0.645 71.790 6.055 71.960 ;
    END
  END in[20]
  PIN in[21]
    DIRECTION INOUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.102000 ;
    PORT
      LAYER li1 ;
        RECT 2.045 68.265 2.215 69.665 ;
        RECT 3.005 68.265 3.175 69.665 ;
        RECT 3.965 68.265 4.135 69.665 ;
        RECT 4.925 68.265 5.095 69.665 ;
        RECT 5.885 68.265 6.055 69.665 ;
        RECT 2.045 66.205 2.215 66.765 ;
        RECT 3.005 66.205 3.175 66.765 ;
        RECT 3.965 66.205 4.135 66.765 ;
        RECT 4.925 66.205 5.095 66.765 ;
        RECT 5.885 66.205 6.055 66.765 ;
      LAYER mcon ;
        RECT 2.045 69.240 2.215 69.410 ;
        RECT 2.045 68.880 2.215 69.050 ;
        RECT 2.045 68.520 2.215 68.690 ;
        RECT 3.005 69.240 3.175 69.410 ;
        RECT 3.005 68.880 3.175 69.050 ;
        RECT 3.005 68.520 3.175 68.690 ;
        RECT 3.965 69.240 4.135 69.410 ;
        RECT 3.965 68.880 4.135 69.050 ;
        RECT 3.965 68.520 4.135 68.690 ;
        RECT 4.925 69.240 5.095 69.410 ;
        RECT 4.925 68.880 5.095 69.050 ;
        RECT 4.925 68.520 5.095 68.690 ;
        RECT 5.885 69.240 6.055 69.410 ;
        RECT 5.885 68.880 6.055 69.050 ;
        RECT 5.885 68.520 6.055 68.690 ;
        RECT 2.045 66.400 2.215 66.570 ;
        RECT 3.005 66.400 3.175 66.570 ;
        RECT 3.965 66.400 4.135 66.570 ;
        RECT 4.925 66.400 5.095 66.570 ;
        RECT 5.885 66.400 6.055 66.570 ;
      LAYER met1 ;
        RECT 0.645 70.395 6.055 70.565 ;
        RECT 0.645 67.580 0.815 70.395 ;
        RECT 2.045 69.645 2.215 70.395 ;
        RECT 3.005 69.645 3.175 70.395 ;
        RECT 3.965 69.645 4.135 70.395 ;
        RECT 4.925 69.645 5.095 70.395 ;
        RECT 5.885 69.645 6.055 70.395 ;
        RECT 2.015 68.285 2.245 69.645 ;
        RECT 2.975 68.285 3.205 69.645 ;
        RECT 3.935 68.285 4.165 69.645 ;
        RECT 4.895 68.285 5.125 69.645 ;
        RECT 5.855 68.285 6.085 69.645 ;
        RECT 0.000 67.410 0.815 67.580 ;
        RECT 0.010 67.405 0.150 67.410 ;
        RECT 0.645 65.525 0.815 67.410 ;
        RECT 2.015 66.225 2.245 66.745 ;
        RECT 2.975 66.225 3.205 66.745 ;
        RECT 3.935 66.225 4.165 66.745 ;
        RECT 4.895 66.225 5.125 66.745 ;
        RECT 5.855 66.225 6.085 66.745 ;
        RECT 2.045 65.525 2.215 66.225 ;
        RECT 3.005 65.525 3.175 66.225 ;
        RECT 3.965 65.525 4.135 66.225 ;
        RECT 4.925 65.525 5.095 66.225 ;
        RECT 5.885 65.525 6.055 66.225 ;
        RECT 0.645 65.355 6.055 65.525 ;
    END
  END in[21]
  PIN in[22]
    DIRECTION INOUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.102000 ;
    PORT
      LAYER li1 ;
        RECT 2.045 61.830 2.215 63.230 ;
        RECT 3.005 61.830 3.175 63.230 ;
        RECT 3.965 61.830 4.135 63.230 ;
        RECT 4.925 61.830 5.095 63.230 ;
        RECT 5.885 61.830 6.055 63.230 ;
        RECT 2.045 59.770 2.215 60.330 ;
        RECT 3.005 59.770 3.175 60.330 ;
        RECT 3.965 59.770 4.135 60.330 ;
        RECT 4.925 59.770 5.095 60.330 ;
        RECT 5.885 59.770 6.055 60.330 ;
      LAYER mcon ;
        RECT 2.045 62.805 2.215 62.975 ;
        RECT 2.045 62.445 2.215 62.615 ;
        RECT 2.045 62.085 2.215 62.255 ;
        RECT 3.005 62.805 3.175 62.975 ;
        RECT 3.005 62.445 3.175 62.615 ;
        RECT 3.005 62.085 3.175 62.255 ;
        RECT 3.965 62.805 4.135 62.975 ;
        RECT 3.965 62.445 4.135 62.615 ;
        RECT 3.965 62.085 4.135 62.255 ;
        RECT 4.925 62.805 5.095 62.975 ;
        RECT 4.925 62.445 5.095 62.615 ;
        RECT 4.925 62.085 5.095 62.255 ;
        RECT 5.885 62.805 6.055 62.975 ;
        RECT 5.885 62.445 6.055 62.615 ;
        RECT 5.885 62.085 6.055 62.255 ;
        RECT 2.045 59.965 2.215 60.135 ;
        RECT 3.005 59.965 3.175 60.135 ;
        RECT 3.965 59.965 4.135 60.135 ;
        RECT 4.925 59.965 5.095 60.135 ;
        RECT 5.885 59.965 6.055 60.135 ;
      LAYER met1 ;
        RECT 0.645 63.960 6.055 64.130 ;
        RECT 0.645 61.145 0.815 63.960 ;
        RECT 2.045 63.210 2.215 63.960 ;
        RECT 3.005 63.210 3.175 63.960 ;
        RECT 3.965 63.210 4.135 63.960 ;
        RECT 4.925 63.210 5.095 63.960 ;
        RECT 5.885 63.210 6.055 63.960 ;
        RECT 2.015 61.850 2.245 63.210 ;
        RECT 2.975 61.850 3.205 63.210 ;
        RECT 3.935 61.850 4.165 63.210 ;
        RECT 4.895 61.850 5.125 63.210 ;
        RECT 5.855 61.850 6.085 63.210 ;
        RECT 0.000 60.975 0.815 61.145 ;
        RECT 0.010 60.970 0.150 60.975 ;
        RECT 0.645 59.090 0.815 60.975 ;
        RECT 2.015 59.790 2.245 60.310 ;
        RECT 2.975 59.790 3.205 60.310 ;
        RECT 3.935 59.790 4.165 60.310 ;
        RECT 4.895 59.790 5.125 60.310 ;
        RECT 5.855 59.790 6.085 60.310 ;
        RECT 2.045 59.090 2.215 59.790 ;
        RECT 3.005 59.090 3.175 59.790 ;
        RECT 3.965 59.090 4.135 59.790 ;
        RECT 4.925 59.090 5.095 59.790 ;
        RECT 5.885 59.090 6.055 59.790 ;
        RECT 0.645 58.920 6.055 59.090 ;
    END
  END in[22]
  PIN in[23]
    DIRECTION INOUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.102000 ;
    PORT
      LAYER li1 ;
        RECT 2.045 55.395 2.215 56.795 ;
        RECT 3.005 55.395 3.175 56.795 ;
        RECT 3.965 55.395 4.135 56.795 ;
        RECT 4.925 55.395 5.095 56.795 ;
        RECT 5.885 55.395 6.055 56.795 ;
        RECT 2.045 53.335 2.215 53.895 ;
        RECT 3.005 53.335 3.175 53.895 ;
        RECT 3.965 53.335 4.135 53.895 ;
        RECT 4.925 53.335 5.095 53.895 ;
        RECT 5.885 53.335 6.055 53.895 ;
      LAYER mcon ;
        RECT 2.045 56.370 2.215 56.540 ;
        RECT 2.045 56.010 2.215 56.180 ;
        RECT 2.045 55.650 2.215 55.820 ;
        RECT 3.005 56.370 3.175 56.540 ;
        RECT 3.005 56.010 3.175 56.180 ;
        RECT 3.005 55.650 3.175 55.820 ;
        RECT 3.965 56.370 4.135 56.540 ;
        RECT 3.965 56.010 4.135 56.180 ;
        RECT 3.965 55.650 4.135 55.820 ;
        RECT 4.925 56.370 5.095 56.540 ;
        RECT 4.925 56.010 5.095 56.180 ;
        RECT 4.925 55.650 5.095 55.820 ;
        RECT 5.885 56.370 6.055 56.540 ;
        RECT 5.885 56.010 6.055 56.180 ;
        RECT 5.885 55.650 6.055 55.820 ;
        RECT 2.045 53.530 2.215 53.700 ;
        RECT 3.005 53.530 3.175 53.700 ;
        RECT 3.965 53.530 4.135 53.700 ;
        RECT 4.925 53.530 5.095 53.700 ;
        RECT 5.885 53.530 6.055 53.700 ;
      LAYER met1 ;
        RECT 0.645 57.525 6.055 57.695 ;
        RECT 0.645 54.710 0.815 57.525 ;
        RECT 2.045 56.775 2.215 57.525 ;
        RECT 3.005 56.775 3.175 57.525 ;
        RECT 3.965 56.775 4.135 57.525 ;
        RECT 4.925 56.775 5.095 57.525 ;
        RECT 5.885 56.775 6.055 57.525 ;
        RECT 2.015 55.415 2.245 56.775 ;
        RECT 2.975 55.415 3.205 56.775 ;
        RECT 3.935 55.415 4.165 56.775 ;
        RECT 4.895 55.415 5.125 56.775 ;
        RECT 5.855 55.415 6.085 56.775 ;
        RECT 0.000 54.540 0.815 54.710 ;
        RECT 0.010 54.535 0.150 54.540 ;
        RECT 0.645 52.655 0.815 54.540 ;
        RECT 2.015 53.355 2.245 53.875 ;
        RECT 2.975 53.355 3.205 53.875 ;
        RECT 3.935 53.355 4.165 53.875 ;
        RECT 4.895 53.355 5.125 53.875 ;
        RECT 5.855 53.355 6.085 53.875 ;
        RECT 2.045 52.655 2.215 53.355 ;
        RECT 3.005 52.655 3.175 53.355 ;
        RECT 3.965 52.655 4.135 53.355 ;
        RECT 4.925 52.655 5.095 53.355 ;
        RECT 5.885 52.655 6.055 53.355 ;
        RECT 0.645 52.485 6.055 52.655 ;
    END
  END in[23]
  PIN in[24]
    DIRECTION INOUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.102000 ;
    PORT
      LAYER li1 ;
        RECT 2.045 48.960 2.215 50.360 ;
        RECT 3.005 48.960 3.175 50.360 ;
        RECT 3.965 48.960 4.135 50.360 ;
        RECT 4.925 48.960 5.095 50.360 ;
        RECT 5.885 48.960 6.055 50.360 ;
        RECT 2.045 46.900 2.215 47.460 ;
        RECT 3.005 46.900 3.175 47.460 ;
        RECT 3.965 46.900 4.135 47.460 ;
        RECT 4.925 46.900 5.095 47.460 ;
        RECT 5.885 46.900 6.055 47.460 ;
      LAYER mcon ;
        RECT 2.045 49.935 2.215 50.105 ;
        RECT 2.045 49.575 2.215 49.745 ;
        RECT 2.045 49.215 2.215 49.385 ;
        RECT 3.005 49.935 3.175 50.105 ;
        RECT 3.005 49.575 3.175 49.745 ;
        RECT 3.005 49.215 3.175 49.385 ;
        RECT 3.965 49.935 4.135 50.105 ;
        RECT 3.965 49.575 4.135 49.745 ;
        RECT 3.965 49.215 4.135 49.385 ;
        RECT 4.925 49.935 5.095 50.105 ;
        RECT 4.925 49.575 5.095 49.745 ;
        RECT 4.925 49.215 5.095 49.385 ;
        RECT 5.885 49.935 6.055 50.105 ;
        RECT 5.885 49.575 6.055 49.745 ;
        RECT 5.885 49.215 6.055 49.385 ;
        RECT 2.045 47.095 2.215 47.265 ;
        RECT 3.005 47.095 3.175 47.265 ;
        RECT 3.965 47.095 4.135 47.265 ;
        RECT 4.925 47.095 5.095 47.265 ;
        RECT 5.885 47.095 6.055 47.265 ;
      LAYER met1 ;
        RECT 0.645 51.090 6.055 51.260 ;
        RECT 0.645 48.275 0.815 51.090 ;
        RECT 2.045 50.340 2.215 51.090 ;
        RECT 3.005 50.340 3.175 51.090 ;
        RECT 3.965 50.340 4.135 51.090 ;
        RECT 4.925 50.340 5.095 51.090 ;
        RECT 5.885 50.340 6.055 51.090 ;
        RECT 2.015 48.980 2.245 50.340 ;
        RECT 2.975 48.980 3.205 50.340 ;
        RECT 3.935 48.980 4.165 50.340 ;
        RECT 4.895 48.980 5.125 50.340 ;
        RECT 5.855 48.980 6.085 50.340 ;
        RECT 0.000 48.105 0.815 48.275 ;
        RECT 0.010 48.100 0.150 48.105 ;
        RECT 0.645 46.220 0.815 48.105 ;
        RECT 2.015 46.920 2.245 47.440 ;
        RECT 2.975 46.920 3.205 47.440 ;
        RECT 3.935 46.920 4.165 47.440 ;
        RECT 4.895 46.920 5.125 47.440 ;
        RECT 5.855 46.920 6.085 47.440 ;
        RECT 2.045 46.220 2.215 46.920 ;
        RECT 3.005 46.220 3.175 46.920 ;
        RECT 3.965 46.220 4.135 46.920 ;
        RECT 4.925 46.220 5.095 46.920 ;
        RECT 5.885 46.220 6.055 46.920 ;
        RECT 0.645 46.050 6.055 46.220 ;
    END
  END in[24]
  PIN in[25]
    DIRECTION INOUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.102000 ;
    PORT
      LAYER li1 ;
        RECT 2.045 42.525 2.215 43.925 ;
        RECT 3.005 42.525 3.175 43.925 ;
        RECT 3.965 42.525 4.135 43.925 ;
        RECT 4.925 42.525 5.095 43.925 ;
        RECT 5.885 42.525 6.055 43.925 ;
        RECT 2.045 40.465 2.215 41.025 ;
        RECT 3.005 40.465 3.175 41.025 ;
        RECT 3.965 40.465 4.135 41.025 ;
        RECT 4.925 40.465 5.095 41.025 ;
        RECT 5.885 40.465 6.055 41.025 ;
      LAYER mcon ;
        RECT 2.045 43.500 2.215 43.670 ;
        RECT 2.045 43.140 2.215 43.310 ;
        RECT 2.045 42.780 2.215 42.950 ;
        RECT 3.005 43.500 3.175 43.670 ;
        RECT 3.005 43.140 3.175 43.310 ;
        RECT 3.005 42.780 3.175 42.950 ;
        RECT 3.965 43.500 4.135 43.670 ;
        RECT 3.965 43.140 4.135 43.310 ;
        RECT 3.965 42.780 4.135 42.950 ;
        RECT 4.925 43.500 5.095 43.670 ;
        RECT 4.925 43.140 5.095 43.310 ;
        RECT 4.925 42.780 5.095 42.950 ;
        RECT 5.885 43.500 6.055 43.670 ;
        RECT 5.885 43.140 6.055 43.310 ;
        RECT 5.885 42.780 6.055 42.950 ;
        RECT 2.045 40.660 2.215 40.830 ;
        RECT 3.005 40.660 3.175 40.830 ;
        RECT 3.965 40.660 4.135 40.830 ;
        RECT 4.925 40.660 5.095 40.830 ;
        RECT 5.885 40.660 6.055 40.830 ;
      LAYER met1 ;
        RECT 0.645 44.655 6.055 44.825 ;
        RECT 0.645 41.840 0.815 44.655 ;
        RECT 2.045 43.905 2.215 44.655 ;
        RECT 3.005 43.905 3.175 44.655 ;
        RECT 3.965 43.905 4.135 44.655 ;
        RECT 4.925 43.905 5.095 44.655 ;
        RECT 5.885 43.905 6.055 44.655 ;
        RECT 2.015 42.545 2.245 43.905 ;
        RECT 2.975 42.545 3.205 43.905 ;
        RECT 3.935 42.545 4.165 43.905 ;
        RECT 4.895 42.545 5.125 43.905 ;
        RECT 5.855 42.545 6.085 43.905 ;
        RECT 0.000 41.670 0.815 41.840 ;
        RECT 0.010 41.665 0.150 41.670 ;
        RECT 0.645 39.785 0.815 41.670 ;
        RECT 2.015 40.485 2.245 41.005 ;
        RECT 2.975 40.485 3.205 41.005 ;
        RECT 3.935 40.485 4.165 41.005 ;
        RECT 4.895 40.485 5.125 41.005 ;
        RECT 5.855 40.485 6.085 41.005 ;
        RECT 2.045 39.785 2.215 40.485 ;
        RECT 3.005 39.785 3.175 40.485 ;
        RECT 3.965 39.785 4.135 40.485 ;
        RECT 4.925 39.785 5.095 40.485 ;
        RECT 5.885 39.785 6.055 40.485 ;
        RECT 0.645 39.615 6.055 39.785 ;
    END
  END in[25]
  PIN in[26]
    DIRECTION INOUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.102000 ;
    PORT
      LAYER li1 ;
        RECT 2.045 36.090 2.215 37.490 ;
        RECT 3.005 36.090 3.175 37.490 ;
        RECT 3.965 36.090 4.135 37.490 ;
        RECT 4.925 36.090 5.095 37.490 ;
        RECT 5.885 36.090 6.055 37.490 ;
        RECT 2.045 34.030 2.215 34.590 ;
        RECT 3.005 34.030 3.175 34.590 ;
        RECT 3.965 34.030 4.135 34.590 ;
        RECT 4.925 34.030 5.095 34.590 ;
        RECT 5.885 34.030 6.055 34.590 ;
      LAYER mcon ;
        RECT 2.045 37.065 2.215 37.235 ;
        RECT 2.045 36.705 2.215 36.875 ;
        RECT 2.045 36.345 2.215 36.515 ;
        RECT 3.005 37.065 3.175 37.235 ;
        RECT 3.005 36.705 3.175 36.875 ;
        RECT 3.005 36.345 3.175 36.515 ;
        RECT 3.965 37.065 4.135 37.235 ;
        RECT 3.965 36.705 4.135 36.875 ;
        RECT 3.965 36.345 4.135 36.515 ;
        RECT 4.925 37.065 5.095 37.235 ;
        RECT 4.925 36.705 5.095 36.875 ;
        RECT 4.925 36.345 5.095 36.515 ;
        RECT 5.885 37.065 6.055 37.235 ;
        RECT 5.885 36.705 6.055 36.875 ;
        RECT 5.885 36.345 6.055 36.515 ;
        RECT 2.045 34.225 2.215 34.395 ;
        RECT 3.005 34.225 3.175 34.395 ;
        RECT 3.965 34.225 4.135 34.395 ;
        RECT 4.925 34.225 5.095 34.395 ;
        RECT 5.885 34.225 6.055 34.395 ;
      LAYER met1 ;
        RECT 0.645 38.220 6.055 38.390 ;
        RECT 0.645 35.405 0.815 38.220 ;
        RECT 2.045 37.470 2.215 38.220 ;
        RECT 3.005 37.470 3.175 38.220 ;
        RECT 3.965 37.470 4.135 38.220 ;
        RECT 4.925 37.470 5.095 38.220 ;
        RECT 5.885 37.470 6.055 38.220 ;
        RECT 2.015 36.110 2.245 37.470 ;
        RECT 2.975 36.110 3.205 37.470 ;
        RECT 3.935 36.110 4.165 37.470 ;
        RECT 4.895 36.110 5.125 37.470 ;
        RECT 5.855 36.110 6.085 37.470 ;
        RECT 0.000 35.235 0.815 35.405 ;
        RECT 0.010 35.230 0.150 35.235 ;
        RECT 0.645 33.350 0.815 35.235 ;
        RECT 2.015 34.050 2.245 34.570 ;
        RECT 2.975 34.050 3.205 34.570 ;
        RECT 3.935 34.050 4.165 34.570 ;
        RECT 4.895 34.050 5.125 34.570 ;
        RECT 5.855 34.050 6.085 34.570 ;
        RECT 2.045 33.350 2.215 34.050 ;
        RECT 3.005 33.350 3.175 34.050 ;
        RECT 3.965 33.350 4.135 34.050 ;
        RECT 4.925 33.350 5.095 34.050 ;
        RECT 5.885 33.350 6.055 34.050 ;
        RECT 0.645 33.180 6.055 33.350 ;
    END
  END in[26]
  PIN in[27]
    DIRECTION INOUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.102000 ;
    PORT
      LAYER li1 ;
        RECT 2.045 29.655 2.215 31.055 ;
        RECT 3.005 29.655 3.175 31.055 ;
        RECT 3.965 29.655 4.135 31.055 ;
        RECT 4.925 29.655 5.095 31.055 ;
        RECT 5.885 29.655 6.055 31.055 ;
        RECT 2.045 27.595 2.215 28.155 ;
        RECT 3.005 27.595 3.175 28.155 ;
        RECT 3.965 27.595 4.135 28.155 ;
        RECT 4.925 27.595 5.095 28.155 ;
        RECT 5.885 27.595 6.055 28.155 ;
      LAYER mcon ;
        RECT 2.045 30.630 2.215 30.800 ;
        RECT 2.045 30.270 2.215 30.440 ;
        RECT 2.045 29.910 2.215 30.080 ;
        RECT 3.005 30.630 3.175 30.800 ;
        RECT 3.005 30.270 3.175 30.440 ;
        RECT 3.005 29.910 3.175 30.080 ;
        RECT 3.965 30.630 4.135 30.800 ;
        RECT 3.965 30.270 4.135 30.440 ;
        RECT 3.965 29.910 4.135 30.080 ;
        RECT 4.925 30.630 5.095 30.800 ;
        RECT 4.925 30.270 5.095 30.440 ;
        RECT 4.925 29.910 5.095 30.080 ;
        RECT 5.885 30.630 6.055 30.800 ;
        RECT 5.885 30.270 6.055 30.440 ;
        RECT 5.885 29.910 6.055 30.080 ;
        RECT 2.045 27.790 2.215 27.960 ;
        RECT 3.005 27.790 3.175 27.960 ;
        RECT 3.965 27.790 4.135 27.960 ;
        RECT 4.925 27.790 5.095 27.960 ;
        RECT 5.885 27.790 6.055 27.960 ;
      LAYER met1 ;
        RECT 0.645 31.785 6.055 31.955 ;
        RECT 0.645 28.970 0.815 31.785 ;
        RECT 2.045 31.035 2.215 31.785 ;
        RECT 3.005 31.035 3.175 31.785 ;
        RECT 3.965 31.035 4.135 31.785 ;
        RECT 4.925 31.035 5.095 31.785 ;
        RECT 5.885 31.035 6.055 31.785 ;
        RECT 2.015 29.675 2.245 31.035 ;
        RECT 2.975 29.675 3.205 31.035 ;
        RECT 3.935 29.675 4.165 31.035 ;
        RECT 4.895 29.675 5.125 31.035 ;
        RECT 5.855 29.675 6.085 31.035 ;
        RECT 0.000 28.800 0.815 28.970 ;
        RECT 0.010 28.795 0.150 28.800 ;
        RECT 0.645 26.915 0.815 28.800 ;
        RECT 2.015 27.615 2.245 28.135 ;
        RECT 2.975 27.615 3.205 28.135 ;
        RECT 3.935 27.615 4.165 28.135 ;
        RECT 4.895 27.615 5.125 28.135 ;
        RECT 5.855 27.615 6.085 28.135 ;
        RECT 2.045 26.915 2.215 27.615 ;
        RECT 3.005 26.915 3.175 27.615 ;
        RECT 3.965 26.915 4.135 27.615 ;
        RECT 4.925 26.915 5.095 27.615 ;
        RECT 5.885 26.915 6.055 27.615 ;
        RECT 0.645 26.745 6.055 26.915 ;
    END
  END in[27]
  PIN in[28]
    DIRECTION INOUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.102000 ;
    PORT
      LAYER li1 ;
        RECT 2.045 23.220 2.215 24.620 ;
        RECT 3.005 23.220 3.175 24.620 ;
        RECT 3.965 23.220 4.135 24.620 ;
        RECT 4.925 23.220 5.095 24.620 ;
        RECT 5.885 23.220 6.055 24.620 ;
        RECT 2.045 21.160 2.215 21.720 ;
        RECT 3.005 21.160 3.175 21.720 ;
        RECT 3.965 21.160 4.135 21.720 ;
        RECT 4.925 21.160 5.095 21.720 ;
        RECT 5.885 21.160 6.055 21.720 ;
      LAYER mcon ;
        RECT 2.045 24.195 2.215 24.365 ;
        RECT 2.045 23.835 2.215 24.005 ;
        RECT 2.045 23.475 2.215 23.645 ;
        RECT 3.005 24.195 3.175 24.365 ;
        RECT 3.005 23.835 3.175 24.005 ;
        RECT 3.005 23.475 3.175 23.645 ;
        RECT 3.965 24.195 4.135 24.365 ;
        RECT 3.965 23.835 4.135 24.005 ;
        RECT 3.965 23.475 4.135 23.645 ;
        RECT 4.925 24.195 5.095 24.365 ;
        RECT 4.925 23.835 5.095 24.005 ;
        RECT 4.925 23.475 5.095 23.645 ;
        RECT 5.885 24.195 6.055 24.365 ;
        RECT 5.885 23.835 6.055 24.005 ;
        RECT 5.885 23.475 6.055 23.645 ;
        RECT 2.045 21.355 2.215 21.525 ;
        RECT 3.005 21.355 3.175 21.525 ;
        RECT 3.965 21.355 4.135 21.525 ;
        RECT 4.925 21.355 5.095 21.525 ;
        RECT 5.885 21.355 6.055 21.525 ;
      LAYER met1 ;
        RECT 0.645 25.350 6.055 25.520 ;
        RECT 0.645 22.535 0.815 25.350 ;
        RECT 2.045 24.600 2.215 25.350 ;
        RECT 3.005 24.600 3.175 25.350 ;
        RECT 3.965 24.600 4.135 25.350 ;
        RECT 4.925 24.600 5.095 25.350 ;
        RECT 5.885 24.600 6.055 25.350 ;
        RECT 2.015 23.240 2.245 24.600 ;
        RECT 2.975 23.240 3.205 24.600 ;
        RECT 3.935 23.240 4.165 24.600 ;
        RECT 4.895 23.240 5.125 24.600 ;
        RECT 5.855 23.240 6.085 24.600 ;
        RECT 0.000 22.365 0.815 22.535 ;
        RECT 0.010 22.360 0.150 22.365 ;
        RECT 0.645 20.480 0.815 22.365 ;
        RECT 2.015 21.180 2.245 21.700 ;
        RECT 2.975 21.180 3.205 21.700 ;
        RECT 3.935 21.180 4.165 21.700 ;
        RECT 4.895 21.180 5.125 21.700 ;
        RECT 5.855 21.180 6.085 21.700 ;
        RECT 2.045 20.480 2.215 21.180 ;
        RECT 3.005 20.480 3.175 21.180 ;
        RECT 3.965 20.480 4.135 21.180 ;
        RECT 4.925 20.480 5.095 21.180 ;
        RECT 5.885 20.480 6.055 21.180 ;
        RECT 0.645 20.310 6.055 20.480 ;
    END
  END in[28]
  PIN in[29]
    DIRECTION INOUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.102000 ;
    PORT
      LAYER li1 ;
        RECT 2.045 16.785 2.215 18.185 ;
        RECT 3.005 16.785 3.175 18.185 ;
        RECT 3.965 16.785 4.135 18.185 ;
        RECT 4.925 16.785 5.095 18.185 ;
        RECT 5.885 16.785 6.055 18.185 ;
        RECT 2.045 14.725 2.215 15.285 ;
        RECT 3.005 14.725 3.175 15.285 ;
        RECT 3.965 14.725 4.135 15.285 ;
        RECT 4.925 14.725 5.095 15.285 ;
        RECT 5.885 14.725 6.055 15.285 ;
      LAYER mcon ;
        RECT 2.045 17.760 2.215 17.930 ;
        RECT 2.045 17.400 2.215 17.570 ;
        RECT 2.045 17.040 2.215 17.210 ;
        RECT 3.005 17.760 3.175 17.930 ;
        RECT 3.005 17.400 3.175 17.570 ;
        RECT 3.005 17.040 3.175 17.210 ;
        RECT 3.965 17.760 4.135 17.930 ;
        RECT 3.965 17.400 4.135 17.570 ;
        RECT 3.965 17.040 4.135 17.210 ;
        RECT 4.925 17.760 5.095 17.930 ;
        RECT 4.925 17.400 5.095 17.570 ;
        RECT 4.925 17.040 5.095 17.210 ;
        RECT 5.885 17.760 6.055 17.930 ;
        RECT 5.885 17.400 6.055 17.570 ;
        RECT 5.885 17.040 6.055 17.210 ;
        RECT 2.045 14.920 2.215 15.090 ;
        RECT 3.005 14.920 3.175 15.090 ;
        RECT 3.965 14.920 4.135 15.090 ;
        RECT 4.925 14.920 5.095 15.090 ;
        RECT 5.885 14.920 6.055 15.090 ;
      LAYER met1 ;
        RECT 0.645 18.915 6.055 19.085 ;
        RECT 0.645 16.100 0.815 18.915 ;
        RECT 2.045 18.165 2.215 18.915 ;
        RECT 3.005 18.165 3.175 18.915 ;
        RECT 3.965 18.165 4.135 18.915 ;
        RECT 4.925 18.165 5.095 18.915 ;
        RECT 5.885 18.165 6.055 18.915 ;
        RECT 2.015 16.805 2.245 18.165 ;
        RECT 2.975 16.805 3.205 18.165 ;
        RECT 3.935 16.805 4.165 18.165 ;
        RECT 4.895 16.805 5.125 18.165 ;
        RECT 5.855 16.805 6.085 18.165 ;
        RECT 0.000 15.930 0.815 16.100 ;
        RECT 0.010 15.925 0.150 15.930 ;
        RECT 0.645 14.045 0.815 15.930 ;
        RECT 2.015 14.745 2.245 15.265 ;
        RECT 2.975 14.745 3.205 15.265 ;
        RECT 3.935 14.745 4.165 15.265 ;
        RECT 4.895 14.745 5.125 15.265 ;
        RECT 5.855 14.745 6.085 15.265 ;
        RECT 2.045 14.045 2.215 14.745 ;
        RECT 3.005 14.045 3.175 14.745 ;
        RECT 3.965 14.045 4.135 14.745 ;
        RECT 4.925 14.045 5.095 14.745 ;
        RECT 5.885 14.045 6.055 14.745 ;
        RECT 0.645 13.875 6.055 14.045 ;
    END
  END in[29]
  PIN in[30]
    DIRECTION INOUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.102000 ;
    PORT
      LAYER li1 ;
        RECT 2.045 10.350 2.215 11.750 ;
        RECT 3.005 10.350 3.175 11.750 ;
        RECT 3.965 10.350 4.135 11.750 ;
        RECT 4.925 10.350 5.095 11.750 ;
        RECT 5.885 10.350 6.055 11.750 ;
        RECT 2.045 8.290 2.215 8.850 ;
        RECT 3.005 8.290 3.175 8.850 ;
        RECT 3.965 8.290 4.135 8.850 ;
        RECT 4.925 8.290 5.095 8.850 ;
        RECT 5.885 8.290 6.055 8.850 ;
      LAYER mcon ;
        RECT 2.045 11.325 2.215 11.495 ;
        RECT 2.045 10.965 2.215 11.135 ;
        RECT 2.045 10.605 2.215 10.775 ;
        RECT 3.005 11.325 3.175 11.495 ;
        RECT 3.005 10.965 3.175 11.135 ;
        RECT 3.005 10.605 3.175 10.775 ;
        RECT 3.965 11.325 4.135 11.495 ;
        RECT 3.965 10.965 4.135 11.135 ;
        RECT 3.965 10.605 4.135 10.775 ;
        RECT 4.925 11.325 5.095 11.495 ;
        RECT 4.925 10.965 5.095 11.135 ;
        RECT 4.925 10.605 5.095 10.775 ;
        RECT 5.885 11.325 6.055 11.495 ;
        RECT 5.885 10.965 6.055 11.135 ;
        RECT 5.885 10.605 6.055 10.775 ;
        RECT 2.045 8.485 2.215 8.655 ;
        RECT 3.005 8.485 3.175 8.655 ;
        RECT 3.965 8.485 4.135 8.655 ;
        RECT 4.925 8.485 5.095 8.655 ;
        RECT 5.885 8.485 6.055 8.655 ;
      LAYER met1 ;
        RECT 0.645 12.480 6.055 12.650 ;
        RECT 0.645 9.665 0.815 12.480 ;
        RECT 2.045 11.730 2.215 12.480 ;
        RECT 3.005 11.730 3.175 12.480 ;
        RECT 3.965 11.730 4.135 12.480 ;
        RECT 4.925 11.730 5.095 12.480 ;
        RECT 5.885 11.730 6.055 12.480 ;
        RECT 2.015 10.370 2.245 11.730 ;
        RECT 2.975 10.370 3.205 11.730 ;
        RECT 3.935 10.370 4.165 11.730 ;
        RECT 4.895 10.370 5.125 11.730 ;
        RECT 5.855 10.370 6.085 11.730 ;
        RECT 0.000 9.495 0.815 9.665 ;
        RECT 0.010 9.490 0.150 9.495 ;
        RECT 0.645 7.610 0.815 9.495 ;
        RECT 2.015 8.310 2.245 8.830 ;
        RECT 2.975 8.310 3.205 8.830 ;
        RECT 3.935 8.310 4.165 8.830 ;
        RECT 4.895 8.310 5.125 8.830 ;
        RECT 5.855 8.310 6.085 8.830 ;
        RECT 2.045 7.610 2.215 8.310 ;
        RECT 3.005 7.610 3.175 8.310 ;
        RECT 3.965 7.610 4.135 8.310 ;
        RECT 4.925 7.610 5.095 8.310 ;
        RECT 5.885 7.610 6.055 8.310 ;
        RECT 0.645 7.440 6.055 7.610 ;
    END
  END in[30]
  PIN in[31]
    DIRECTION INOUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.102000 ;
    PORT
      LAYER li1 ;
        RECT 2.045 3.915 2.215 5.315 ;
        RECT 3.005 3.915 3.175 5.315 ;
        RECT 3.965 3.915 4.135 5.315 ;
        RECT 4.925 3.915 5.095 5.315 ;
        RECT 5.885 3.915 6.055 5.315 ;
        RECT 2.045 1.855 2.215 2.415 ;
        RECT 3.005 1.855 3.175 2.415 ;
        RECT 3.965 1.855 4.135 2.415 ;
        RECT 4.925 1.855 5.095 2.415 ;
        RECT 5.885 1.855 6.055 2.415 ;
      LAYER mcon ;
        RECT 2.045 4.890 2.215 5.060 ;
        RECT 2.045 4.530 2.215 4.700 ;
        RECT 2.045 4.170 2.215 4.340 ;
        RECT 3.005 4.890 3.175 5.060 ;
        RECT 3.005 4.530 3.175 4.700 ;
        RECT 3.005 4.170 3.175 4.340 ;
        RECT 3.965 4.890 4.135 5.060 ;
        RECT 3.965 4.530 4.135 4.700 ;
        RECT 3.965 4.170 4.135 4.340 ;
        RECT 4.925 4.890 5.095 5.060 ;
        RECT 4.925 4.530 5.095 4.700 ;
        RECT 4.925 4.170 5.095 4.340 ;
        RECT 5.885 4.890 6.055 5.060 ;
        RECT 5.885 4.530 6.055 4.700 ;
        RECT 5.885 4.170 6.055 4.340 ;
        RECT 2.045 2.050 2.215 2.220 ;
        RECT 3.005 2.050 3.175 2.220 ;
        RECT 3.965 2.050 4.135 2.220 ;
        RECT 4.925 2.050 5.095 2.220 ;
        RECT 5.885 2.050 6.055 2.220 ;
      LAYER met1 ;
        RECT 0.645 6.045 6.055 6.215 ;
        RECT 0.645 3.230 0.815 6.045 ;
        RECT 2.045 5.295 2.215 6.045 ;
        RECT 3.005 5.295 3.175 6.045 ;
        RECT 3.965 5.295 4.135 6.045 ;
        RECT 4.925 5.295 5.095 6.045 ;
        RECT 5.885 5.295 6.055 6.045 ;
        RECT 2.015 3.935 2.245 5.295 ;
        RECT 2.975 3.935 3.205 5.295 ;
        RECT 3.935 3.935 4.165 5.295 ;
        RECT 4.895 3.935 5.125 5.295 ;
        RECT 5.855 3.935 6.085 5.295 ;
        RECT 0.000 3.060 0.815 3.230 ;
        RECT 0.010 3.055 0.150 3.060 ;
        RECT 0.645 1.175 0.815 3.060 ;
        RECT 2.015 1.875 2.245 2.395 ;
        RECT 2.975 1.875 3.205 2.395 ;
        RECT 3.935 1.875 4.165 2.395 ;
        RECT 4.895 1.875 5.125 2.395 ;
        RECT 5.855 1.875 6.085 2.395 ;
        RECT 2.045 1.175 2.215 1.875 ;
        RECT 3.005 1.175 3.175 1.875 ;
        RECT 3.965 1.175 4.135 1.875 ;
        RECT 4.925 1.175 5.095 1.875 ;
        RECT 5.885 1.175 6.055 1.875 ;
        RECT 0.645 1.005 6.055 1.175 ;
    END
  END in[31]
  PIN en_b[0]
    DIRECTION INOUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 4.402500 ;
    PORT
      LAYER li1 ;
        RECT 12.250 205.040 12.580 205.210 ;
        RECT 13.210 205.040 13.540 205.210 ;
        RECT 14.170 205.040 14.500 205.210 ;
        RECT 15.130 205.040 15.460 205.210 ;
        RECT 16.090 205.040 16.420 205.210 ;
        RECT 17.050 205.040 17.380 205.210 ;
        RECT 19.855 205.040 20.185 205.210 ;
        RECT 20.815 205.040 21.145 205.210 ;
        RECT 21.775 205.040 22.105 205.210 ;
        RECT 22.735 205.040 23.065 205.210 ;
        RECT 23.695 205.040 24.025 205.210 ;
        RECT 24.655 205.040 24.985 205.210 ;
        RECT 27.100 202.325 27.430 202.565 ;
        RECT 18.375 202.110 18.705 202.280 ;
      LAYER mcon ;
        RECT 12.330 205.040 12.500 205.210 ;
        RECT 13.290 205.040 13.460 205.210 ;
        RECT 14.250 205.040 14.420 205.210 ;
        RECT 15.210 205.040 15.380 205.210 ;
        RECT 16.170 205.040 16.340 205.210 ;
        RECT 17.130 205.040 17.300 205.210 ;
        RECT 19.935 205.040 20.105 205.210 ;
        RECT 20.895 205.040 21.065 205.210 ;
        RECT 21.855 205.040 22.025 205.210 ;
        RECT 22.815 205.040 22.985 205.210 ;
        RECT 23.775 205.040 23.945 205.210 ;
        RECT 24.735 205.040 24.905 205.210 ;
        RECT 27.250 202.340 27.420 202.510 ;
        RECT 18.455 202.110 18.625 202.280 ;
      LAYER met1 ;
        RECT 12.235 205.000 12.595 205.260 ;
        RECT 13.200 205.000 13.560 205.260 ;
        RECT 14.155 205.000 14.515 205.260 ;
        RECT 15.115 205.000 15.475 205.260 ;
        RECT 16.075 205.000 16.435 205.260 ;
        RECT 17.035 205.000 17.395 205.260 ;
        RECT 19.840 205.000 20.200 205.260 ;
        RECT 20.805 205.000 21.165 205.260 ;
        RECT 21.760 205.000 22.120 205.260 ;
        RECT 22.720 205.000 23.080 205.260 ;
        RECT 23.680 205.000 24.040 205.260 ;
        RECT 24.640 205.000 25.000 205.260 ;
        RECT 18.355 202.115 18.715 202.375 ;
        RECT 27.190 202.280 27.560 202.550 ;
        RECT 18.395 202.080 18.685 202.115 ;
      LAYER via ;
        RECT 12.285 205.000 12.545 205.260 ;
        RECT 13.250 205.000 13.510 205.260 ;
        RECT 14.205 205.000 14.465 205.260 ;
        RECT 15.165 205.000 15.425 205.260 ;
        RECT 16.125 205.000 16.385 205.260 ;
        RECT 17.085 205.000 17.345 205.260 ;
        RECT 19.890 205.000 20.150 205.260 ;
        RECT 20.855 205.000 21.115 205.260 ;
        RECT 21.810 205.000 22.070 205.260 ;
        RECT 22.770 205.000 23.030 205.260 ;
        RECT 23.730 205.000 23.990 205.260 ;
        RECT 24.690 205.000 24.950 205.260 ;
        RECT 18.405 202.115 18.665 202.375 ;
        RECT 27.245 202.285 27.505 202.545 ;
      LAYER met2 ;
        RECT 12.285 205.260 12.545 205.310 ;
        RECT 13.250 205.260 13.510 205.310 ;
        RECT 14.205 205.260 14.465 205.310 ;
        RECT 15.165 205.260 15.425 205.310 ;
        RECT 16.125 205.260 16.385 205.310 ;
        RECT 17.085 205.260 17.345 205.310 ;
        RECT 19.890 205.260 20.150 205.310 ;
        RECT 20.855 205.260 21.115 205.310 ;
        RECT 21.810 205.260 22.070 205.310 ;
        RECT 22.770 205.260 23.030 205.310 ;
        RECT 23.730 205.260 23.990 205.310 ;
        RECT 24.690 205.260 24.950 205.310 ;
        RECT 11.165 205.000 29.230 205.260 ;
        RECT 12.285 204.950 12.545 205.000 ;
        RECT 13.250 204.950 13.510 205.000 ;
        RECT 14.205 204.950 14.465 205.000 ;
        RECT 15.165 204.950 15.425 205.000 ;
        RECT 16.125 204.950 16.385 205.000 ;
        RECT 17.085 204.950 17.345 205.000 ;
        RECT 18.405 202.065 18.665 205.000 ;
        RECT 19.890 204.950 20.150 205.000 ;
        RECT 20.855 204.950 21.115 205.000 ;
        RECT 21.810 204.950 22.070 205.000 ;
        RECT 22.770 204.950 23.030 205.000 ;
        RECT 23.730 204.950 23.990 205.000 ;
        RECT 24.690 204.950 24.950 205.000 ;
        RECT 27.240 202.580 27.510 202.600 ;
        RECT 28.040 202.580 28.300 205.000 ;
        RECT 27.240 202.320 28.300 202.580 ;
        RECT 27.240 202.230 27.510 202.320 ;
    END
  END en_b[0]
  PIN en_b[1]
    DIRECTION INOUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 4.402500 ;
    PORT
      LAYER li1 ;
        RECT 12.250 198.605 12.580 198.775 ;
        RECT 13.210 198.605 13.540 198.775 ;
        RECT 14.170 198.605 14.500 198.775 ;
        RECT 15.130 198.605 15.460 198.775 ;
        RECT 16.090 198.605 16.420 198.775 ;
        RECT 17.050 198.605 17.380 198.775 ;
        RECT 19.855 198.605 20.185 198.775 ;
        RECT 20.815 198.605 21.145 198.775 ;
        RECT 21.775 198.605 22.105 198.775 ;
        RECT 22.735 198.605 23.065 198.775 ;
        RECT 23.695 198.605 24.025 198.775 ;
        RECT 24.655 198.605 24.985 198.775 ;
        RECT 27.100 195.890 27.430 196.130 ;
        RECT 18.375 195.675 18.705 195.845 ;
      LAYER mcon ;
        RECT 12.330 198.605 12.500 198.775 ;
        RECT 13.290 198.605 13.460 198.775 ;
        RECT 14.250 198.605 14.420 198.775 ;
        RECT 15.210 198.605 15.380 198.775 ;
        RECT 16.170 198.605 16.340 198.775 ;
        RECT 17.130 198.605 17.300 198.775 ;
        RECT 19.935 198.605 20.105 198.775 ;
        RECT 20.895 198.605 21.065 198.775 ;
        RECT 21.855 198.605 22.025 198.775 ;
        RECT 22.815 198.605 22.985 198.775 ;
        RECT 23.775 198.605 23.945 198.775 ;
        RECT 24.735 198.605 24.905 198.775 ;
        RECT 27.250 195.905 27.420 196.075 ;
        RECT 18.455 195.675 18.625 195.845 ;
      LAYER met1 ;
        RECT 12.235 198.565 12.595 198.825 ;
        RECT 13.200 198.565 13.560 198.825 ;
        RECT 14.155 198.565 14.515 198.825 ;
        RECT 15.115 198.565 15.475 198.825 ;
        RECT 16.075 198.565 16.435 198.825 ;
        RECT 17.035 198.565 17.395 198.825 ;
        RECT 19.840 198.565 20.200 198.825 ;
        RECT 20.805 198.565 21.165 198.825 ;
        RECT 21.760 198.565 22.120 198.825 ;
        RECT 22.720 198.565 23.080 198.825 ;
        RECT 23.680 198.565 24.040 198.825 ;
        RECT 24.640 198.565 25.000 198.825 ;
        RECT 18.355 195.680 18.715 195.940 ;
        RECT 27.190 195.845 27.560 196.115 ;
        RECT 18.395 195.645 18.685 195.680 ;
      LAYER via ;
        RECT 12.285 198.565 12.545 198.825 ;
        RECT 13.250 198.565 13.510 198.825 ;
        RECT 14.205 198.565 14.465 198.825 ;
        RECT 15.165 198.565 15.425 198.825 ;
        RECT 16.125 198.565 16.385 198.825 ;
        RECT 17.085 198.565 17.345 198.825 ;
        RECT 19.890 198.565 20.150 198.825 ;
        RECT 20.855 198.565 21.115 198.825 ;
        RECT 21.810 198.565 22.070 198.825 ;
        RECT 22.770 198.565 23.030 198.825 ;
        RECT 23.730 198.565 23.990 198.825 ;
        RECT 24.690 198.565 24.950 198.825 ;
        RECT 18.405 195.680 18.665 195.940 ;
        RECT 27.245 195.850 27.505 196.110 ;
      LAYER met2 ;
        RECT 12.285 198.825 12.545 198.875 ;
        RECT 13.250 198.825 13.510 198.875 ;
        RECT 14.205 198.825 14.465 198.875 ;
        RECT 15.165 198.825 15.425 198.875 ;
        RECT 16.125 198.825 16.385 198.875 ;
        RECT 17.085 198.825 17.345 198.875 ;
        RECT 19.890 198.825 20.150 198.875 ;
        RECT 20.855 198.825 21.115 198.875 ;
        RECT 21.810 198.825 22.070 198.875 ;
        RECT 22.770 198.825 23.030 198.875 ;
        RECT 23.730 198.825 23.990 198.875 ;
        RECT 24.690 198.825 24.950 198.875 ;
        RECT 11.165 198.565 29.230 198.825 ;
        RECT 12.285 198.515 12.545 198.565 ;
        RECT 13.250 198.515 13.510 198.565 ;
        RECT 14.205 198.515 14.465 198.565 ;
        RECT 15.165 198.515 15.425 198.565 ;
        RECT 16.125 198.515 16.385 198.565 ;
        RECT 17.085 198.515 17.345 198.565 ;
        RECT 18.405 195.630 18.665 198.565 ;
        RECT 19.890 198.515 20.150 198.565 ;
        RECT 20.855 198.515 21.115 198.565 ;
        RECT 21.810 198.515 22.070 198.565 ;
        RECT 22.770 198.515 23.030 198.565 ;
        RECT 23.730 198.515 23.990 198.565 ;
        RECT 24.690 198.515 24.950 198.565 ;
        RECT 27.240 196.145 27.510 196.165 ;
        RECT 28.040 196.145 28.300 198.565 ;
        RECT 27.240 195.885 28.300 196.145 ;
        RECT 27.240 195.795 27.510 195.885 ;
    END
  END en_b[1]
  PIN en_b[2]
    DIRECTION INOUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 4.402500 ;
    PORT
      LAYER li1 ;
        RECT 12.250 192.170 12.580 192.340 ;
        RECT 13.210 192.170 13.540 192.340 ;
        RECT 14.170 192.170 14.500 192.340 ;
        RECT 15.130 192.170 15.460 192.340 ;
        RECT 16.090 192.170 16.420 192.340 ;
        RECT 17.050 192.170 17.380 192.340 ;
        RECT 19.855 192.170 20.185 192.340 ;
        RECT 20.815 192.170 21.145 192.340 ;
        RECT 21.775 192.170 22.105 192.340 ;
        RECT 22.735 192.170 23.065 192.340 ;
        RECT 23.695 192.170 24.025 192.340 ;
        RECT 24.655 192.170 24.985 192.340 ;
        RECT 27.100 189.455 27.430 189.695 ;
        RECT 18.375 189.240 18.705 189.410 ;
      LAYER mcon ;
        RECT 12.330 192.170 12.500 192.340 ;
        RECT 13.290 192.170 13.460 192.340 ;
        RECT 14.250 192.170 14.420 192.340 ;
        RECT 15.210 192.170 15.380 192.340 ;
        RECT 16.170 192.170 16.340 192.340 ;
        RECT 17.130 192.170 17.300 192.340 ;
        RECT 19.935 192.170 20.105 192.340 ;
        RECT 20.895 192.170 21.065 192.340 ;
        RECT 21.855 192.170 22.025 192.340 ;
        RECT 22.815 192.170 22.985 192.340 ;
        RECT 23.775 192.170 23.945 192.340 ;
        RECT 24.735 192.170 24.905 192.340 ;
        RECT 27.250 189.470 27.420 189.640 ;
        RECT 18.455 189.240 18.625 189.410 ;
      LAYER met1 ;
        RECT 12.235 192.130 12.595 192.390 ;
        RECT 13.200 192.130 13.560 192.390 ;
        RECT 14.155 192.130 14.515 192.390 ;
        RECT 15.115 192.130 15.475 192.390 ;
        RECT 16.075 192.130 16.435 192.390 ;
        RECT 17.035 192.130 17.395 192.390 ;
        RECT 19.840 192.130 20.200 192.390 ;
        RECT 20.805 192.130 21.165 192.390 ;
        RECT 21.760 192.130 22.120 192.390 ;
        RECT 22.720 192.130 23.080 192.390 ;
        RECT 23.680 192.130 24.040 192.390 ;
        RECT 24.640 192.130 25.000 192.390 ;
        RECT 18.355 189.245 18.715 189.505 ;
        RECT 27.190 189.410 27.560 189.680 ;
        RECT 18.395 189.210 18.685 189.245 ;
      LAYER via ;
        RECT 12.285 192.130 12.545 192.390 ;
        RECT 13.250 192.130 13.510 192.390 ;
        RECT 14.205 192.130 14.465 192.390 ;
        RECT 15.165 192.130 15.425 192.390 ;
        RECT 16.125 192.130 16.385 192.390 ;
        RECT 17.085 192.130 17.345 192.390 ;
        RECT 19.890 192.130 20.150 192.390 ;
        RECT 20.855 192.130 21.115 192.390 ;
        RECT 21.810 192.130 22.070 192.390 ;
        RECT 22.770 192.130 23.030 192.390 ;
        RECT 23.730 192.130 23.990 192.390 ;
        RECT 24.690 192.130 24.950 192.390 ;
        RECT 18.405 189.245 18.665 189.505 ;
        RECT 27.245 189.415 27.505 189.675 ;
      LAYER met2 ;
        RECT 12.285 192.390 12.545 192.440 ;
        RECT 13.250 192.390 13.510 192.440 ;
        RECT 14.205 192.390 14.465 192.440 ;
        RECT 15.165 192.390 15.425 192.440 ;
        RECT 16.125 192.390 16.385 192.440 ;
        RECT 17.085 192.390 17.345 192.440 ;
        RECT 19.890 192.390 20.150 192.440 ;
        RECT 20.855 192.390 21.115 192.440 ;
        RECT 21.810 192.390 22.070 192.440 ;
        RECT 22.770 192.390 23.030 192.440 ;
        RECT 23.730 192.390 23.990 192.440 ;
        RECT 24.690 192.390 24.950 192.440 ;
        RECT 11.165 192.130 29.230 192.390 ;
        RECT 12.285 192.080 12.545 192.130 ;
        RECT 13.250 192.080 13.510 192.130 ;
        RECT 14.205 192.080 14.465 192.130 ;
        RECT 15.165 192.080 15.425 192.130 ;
        RECT 16.125 192.080 16.385 192.130 ;
        RECT 17.085 192.080 17.345 192.130 ;
        RECT 18.405 189.195 18.665 192.130 ;
        RECT 19.890 192.080 20.150 192.130 ;
        RECT 20.855 192.080 21.115 192.130 ;
        RECT 21.810 192.080 22.070 192.130 ;
        RECT 22.770 192.080 23.030 192.130 ;
        RECT 23.730 192.080 23.990 192.130 ;
        RECT 24.690 192.080 24.950 192.130 ;
        RECT 27.240 189.710 27.510 189.730 ;
        RECT 28.040 189.710 28.300 192.130 ;
        RECT 27.240 189.450 28.300 189.710 ;
        RECT 27.240 189.360 27.510 189.450 ;
    END
  END en_b[2]
  PIN en_b[3]
    DIRECTION INOUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 4.402500 ;
    PORT
      LAYER li1 ;
        RECT 12.250 185.735 12.580 185.905 ;
        RECT 13.210 185.735 13.540 185.905 ;
        RECT 14.170 185.735 14.500 185.905 ;
        RECT 15.130 185.735 15.460 185.905 ;
        RECT 16.090 185.735 16.420 185.905 ;
        RECT 17.050 185.735 17.380 185.905 ;
        RECT 19.855 185.735 20.185 185.905 ;
        RECT 20.815 185.735 21.145 185.905 ;
        RECT 21.775 185.735 22.105 185.905 ;
        RECT 22.735 185.735 23.065 185.905 ;
        RECT 23.695 185.735 24.025 185.905 ;
        RECT 24.655 185.735 24.985 185.905 ;
        RECT 27.100 183.020 27.430 183.260 ;
        RECT 18.375 182.805 18.705 182.975 ;
      LAYER mcon ;
        RECT 12.330 185.735 12.500 185.905 ;
        RECT 13.290 185.735 13.460 185.905 ;
        RECT 14.250 185.735 14.420 185.905 ;
        RECT 15.210 185.735 15.380 185.905 ;
        RECT 16.170 185.735 16.340 185.905 ;
        RECT 17.130 185.735 17.300 185.905 ;
        RECT 19.935 185.735 20.105 185.905 ;
        RECT 20.895 185.735 21.065 185.905 ;
        RECT 21.855 185.735 22.025 185.905 ;
        RECT 22.815 185.735 22.985 185.905 ;
        RECT 23.775 185.735 23.945 185.905 ;
        RECT 24.735 185.735 24.905 185.905 ;
        RECT 27.250 183.035 27.420 183.205 ;
        RECT 18.455 182.805 18.625 182.975 ;
      LAYER met1 ;
        RECT 12.235 185.695 12.595 185.955 ;
        RECT 13.200 185.695 13.560 185.955 ;
        RECT 14.155 185.695 14.515 185.955 ;
        RECT 15.115 185.695 15.475 185.955 ;
        RECT 16.075 185.695 16.435 185.955 ;
        RECT 17.035 185.695 17.395 185.955 ;
        RECT 19.840 185.695 20.200 185.955 ;
        RECT 20.805 185.695 21.165 185.955 ;
        RECT 21.760 185.695 22.120 185.955 ;
        RECT 22.720 185.695 23.080 185.955 ;
        RECT 23.680 185.695 24.040 185.955 ;
        RECT 24.640 185.695 25.000 185.955 ;
        RECT 18.355 182.810 18.715 183.070 ;
        RECT 27.190 182.975 27.560 183.245 ;
        RECT 18.395 182.775 18.685 182.810 ;
      LAYER via ;
        RECT 12.285 185.695 12.545 185.955 ;
        RECT 13.250 185.695 13.510 185.955 ;
        RECT 14.205 185.695 14.465 185.955 ;
        RECT 15.165 185.695 15.425 185.955 ;
        RECT 16.125 185.695 16.385 185.955 ;
        RECT 17.085 185.695 17.345 185.955 ;
        RECT 19.890 185.695 20.150 185.955 ;
        RECT 20.855 185.695 21.115 185.955 ;
        RECT 21.810 185.695 22.070 185.955 ;
        RECT 22.770 185.695 23.030 185.955 ;
        RECT 23.730 185.695 23.990 185.955 ;
        RECT 24.690 185.695 24.950 185.955 ;
        RECT 18.405 182.810 18.665 183.070 ;
        RECT 27.245 182.980 27.505 183.240 ;
      LAYER met2 ;
        RECT 12.285 185.955 12.545 186.005 ;
        RECT 13.250 185.955 13.510 186.005 ;
        RECT 14.205 185.955 14.465 186.005 ;
        RECT 15.165 185.955 15.425 186.005 ;
        RECT 16.125 185.955 16.385 186.005 ;
        RECT 17.085 185.955 17.345 186.005 ;
        RECT 19.890 185.955 20.150 186.005 ;
        RECT 20.855 185.955 21.115 186.005 ;
        RECT 21.810 185.955 22.070 186.005 ;
        RECT 22.770 185.955 23.030 186.005 ;
        RECT 23.730 185.955 23.990 186.005 ;
        RECT 24.690 185.955 24.950 186.005 ;
        RECT 11.165 185.695 29.230 185.955 ;
        RECT 12.285 185.645 12.545 185.695 ;
        RECT 13.250 185.645 13.510 185.695 ;
        RECT 14.205 185.645 14.465 185.695 ;
        RECT 15.165 185.645 15.425 185.695 ;
        RECT 16.125 185.645 16.385 185.695 ;
        RECT 17.085 185.645 17.345 185.695 ;
        RECT 18.405 182.760 18.665 185.695 ;
        RECT 19.890 185.645 20.150 185.695 ;
        RECT 20.855 185.645 21.115 185.695 ;
        RECT 21.810 185.645 22.070 185.695 ;
        RECT 22.770 185.645 23.030 185.695 ;
        RECT 23.730 185.645 23.990 185.695 ;
        RECT 24.690 185.645 24.950 185.695 ;
        RECT 27.240 183.275 27.510 183.295 ;
        RECT 28.040 183.275 28.300 185.695 ;
        RECT 27.240 183.015 28.300 183.275 ;
        RECT 27.240 182.925 27.510 183.015 ;
    END
  END en_b[3]
  PIN en_b[4]
    DIRECTION INOUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 4.402500 ;
    PORT
      LAYER li1 ;
        RECT 12.250 179.300 12.580 179.470 ;
        RECT 13.210 179.300 13.540 179.470 ;
        RECT 14.170 179.300 14.500 179.470 ;
        RECT 15.130 179.300 15.460 179.470 ;
        RECT 16.090 179.300 16.420 179.470 ;
        RECT 17.050 179.300 17.380 179.470 ;
        RECT 19.855 179.300 20.185 179.470 ;
        RECT 20.815 179.300 21.145 179.470 ;
        RECT 21.775 179.300 22.105 179.470 ;
        RECT 22.735 179.300 23.065 179.470 ;
        RECT 23.695 179.300 24.025 179.470 ;
        RECT 24.655 179.300 24.985 179.470 ;
        RECT 27.100 176.585 27.430 176.825 ;
        RECT 18.375 176.370 18.705 176.540 ;
      LAYER mcon ;
        RECT 12.330 179.300 12.500 179.470 ;
        RECT 13.290 179.300 13.460 179.470 ;
        RECT 14.250 179.300 14.420 179.470 ;
        RECT 15.210 179.300 15.380 179.470 ;
        RECT 16.170 179.300 16.340 179.470 ;
        RECT 17.130 179.300 17.300 179.470 ;
        RECT 19.935 179.300 20.105 179.470 ;
        RECT 20.895 179.300 21.065 179.470 ;
        RECT 21.855 179.300 22.025 179.470 ;
        RECT 22.815 179.300 22.985 179.470 ;
        RECT 23.775 179.300 23.945 179.470 ;
        RECT 24.735 179.300 24.905 179.470 ;
        RECT 27.250 176.600 27.420 176.770 ;
        RECT 18.455 176.370 18.625 176.540 ;
      LAYER met1 ;
        RECT 12.235 179.260 12.595 179.520 ;
        RECT 13.200 179.260 13.560 179.520 ;
        RECT 14.155 179.260 14.515 179.520 ;
        RECT 15.115 179.260 15.475 179.520 ;
        RECT 16.075 179.260 16.435 179.520 ;
        RECT 17.035 179.260 17.395 179.520 ;
        RECT 19.840 179.260 20.200 179.520 ;
        RECT 20.805 179.260 21.165 179.520 ;
        RECT 21.760 179.260 22.120 179.520 ;
        RECT 22.720 179.260 23.080 179.520 ;
        RECT 23.680 179.260 24.040 179.520 ;
        RECT 24.640 179.260 25.000 179.520 ;
        RECT 18.355 176.375 18.715 176.635 ;
        RECT 27.190 176.540 27.560 176.810 ;
        RECT 18.395 176.340 18.685 176.375 ;
      LAYER via ;
        RECT 12.285 179.260 12.545 179.520 ;
        RECT 13.250 179.260 13.510 179.520 ;
        RECT 14.205 179.260 14.465 179.520 ;
        RECT 15.165 179.260 15.425 179.520 ;
        RECT 16.125 179.260 16.385 179.520 ;
        RECT 17.085 179.260 17.345 179.520 ;
        RECT 19.890 179.260 20.150 179.520 ;
        RECT 20.855 179.260 21.115 179.520 ;
        RECT 21.810 179.260 22.070 179.520 ;
        RECT 22.770 179.260 23.030 179.520 ;
        RECT 23.730 179.260 23.990 179.520 ;
        RECT 24.690 179.260 24.950 179.520 ;
        RECT 18.405 176.375 18.665 176.635 ;
        RECT 27.245 176.545 27.505 176.805 ;
      LAYER met2 ;
        RECT 12.285 179.520 12.545 179.570 ;
        RECT 13.250 179.520 13.510 179.570 ;
        RECT 14.205 179.520 14.465 179.570 ;
        RECT 15.165 179.520 15.425 179.570 ;
        RECT 16.125 179.520 16.385 179.570 ;
        RECT 17.085 179.520 17.345 179.570 ;
        RECT 19.890 179.520 20.150 179.570 ;
        RECT 20.855 179.520 21.115 179.570 ;
        RECT 21.810 179.520 22.070 179.570 ;
        RECT 22.770 179.520 23.030 179.570 ;
        RECT 23.730 179.520 23.990 179.570 ;
        RECT 24.690 179.520 24.950 179.570 ;
        RECT 11.165 179.260 29.230 179.520 ;
        RECT 12.285 179.210 12.545 179.260 ;
        RECT 13.250 179.210 13.510 179.260 ;
        RECT 14.205 179.210 14.465 179.260 ;
        RECT 15.165 179.210 15.425 179.260 ;
        RECT 16.125 179.210 16.385 179.260 ;
        RECT 17.085 179.210 17.345 179.260 ;
        RECT 18.405 176.325 18.665 179.260 ;
        RECT 19.890 179.210 20.150 179.260 ;
        RECT 20.855 179.210 21.115 179.260 ;
        RECT 21.810 179.210 22.070 179.260 ;
        RECT 22.770 179.210 23.030 179.260 ;
        RECT 23.730 179.210 23.990 179.260 ;
        RECT 24.690 179.210 24.950 179.260 ;
        RECT 27.240 176.840 27.510 176.860 ;
        RECT 28.040 176.840 28.300 179.260 ;
        RECT 27.240 176.580 28.300 176.840 ;
        RECT 27.240 176.490 27.510 176.580 ;
    END
  END en_b[4]
  PIN en_b[5]
    DIRECTION INOUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 4.402500 ;
    PORT
      LAYER li1 ;
        RECT 12.250 172.865 12.580 173.035 ;
        RECT 13.210 172.865 13.540 173.035 ;
        RECT 14.170 172.865 14.500 173.035 ;
        RECT 15.130 172.865 15.460 173.035 ;
        RECT 16.090 172.865 16.420 173.035 ;
        RECT 17.050 172.865 17.380 173.035 ;
        RECT 19.855 172.865 20.185 173.035 ;
        RECT 20.815 172.865 21.145 173.035 ;
        RECT 21.775 172.865 22.105 173.035 ;
        RECT 22.735 172.865 23.065 173.035 ;
        RECT 23.695 172.865 24.025 173.035 ;
        RECT 24.655 172.865 24.985 173.035 ;
        RECT 27.100 170.150 27.430 170.390 ;
        RECT 18.375 169.935 18.705 170.105 ;
      LAYER mcon ;
        RECT 12.330 172.865 12.500 173.035 ;
        RECT 13.290 172.865 13.460 173.035 ;
        RECT 14.250 172.865 14.420 173.035 ;
        RECT 15.210 172.865 15.380 173.035 ;
        RECT 16.170 172.865 16.340 173.035 ;
        RECT 17.130 172.865 17.300 173.035 ;
        RECT 19.935 172.865 20.105 173.035 ;
        RECT 20.895 172.865 21.065 173.035 ;
        RECT 21.855 172.865 22.025 173.035 ;
        RECT 22.815 172.865 22.985 173.035 ;
        RECT 23.775 172.865 23.945 173.035 ;
        RECT 24.735 172.865 24.905 173.035 ;
        RECT 27.250 170.165 27.420 170.335 ;
        RECT 18.455 169.935 18.625 170.105 ;
      LAYER met1 ;
        RECT 12.235 172.825 12.595 173.085 ;
        RECT 13.200 172.825 13.560 173.085 ;
        RECT 14.155 172.825 14.515 173.085 ;
        RECT 15.115 172.825 15.475 173.085 ;
        RECT 16.075 172.825 16.435 173.085 ;
        RECT 17.035 172.825 17.395 173.085 ;
        RECT 19.840 172.825 20.200 173.085 ;
        RECT 20.805 172.825 21.165 173.085 ;
        RECT 21.760 172.825 22.120 173.085 ;
        RECT 22.720 172.825 23.080 173.085 ;
        RECT 23.680 172.825 24.040 173.085 ;
        RECT 24.640 172.825 25.000 173.085 ;
        RECT 18.355 169.940 18.715 170.200 ;
        RECT 27.190 170.105 27.560 170.375 ;
        RECT 18.395 169.905 18.685 169.940 ;
      LAYER via ;
        RECT 12.285 172.825 12.545 173.085 ;
        RECT 13.250 172.825 13.510 173.085 ;
        RECT 14.205 172.825 14.465 173.085 ;
        RECT 15.165 172.825 15.425 173.085 ;
        RECT 16.125 172.825 16.385 173.085 ;
        RECT 17.085 172.825 17.345 173.085 ;
        RECT 19.890 172.825 20.150 173.085 ;
        RECT 20.855 172.825 21.115 173.085 ;
        RECT 21.810 172.825 22.070 173.085 ;
        RECT 22.770 172.825 23.030 173.085 ;
        RECT 23.730 172.825 23.990 173.085 ;
        RECT 24.690 172.825 24.950 173.085 ;
        RECT 18.405 169.940 18.665 170.200 ;
        RECT 27.245 170.110 27.505 170.370 ;
      LAYER met2 ;
        RECT 12.285 173.085 12.545 173.135 ;
        RECT 13.250 173.085 13.510 173.135 ;
        RECT 14.205 173.085 14.465 173.135 ;
        RECT 15.165 173.085 15.425 173.135 ;
        RECT 16.125 173.085 16.385 173.135 ;
        RECT 17.085 173.085 17.345 173.135 ;
        RECT 19.890 173.085 20.150 173.135 ;
        RECT 20.855 173.085 21.115 173.135 ;
        RECT 21.810 173.085 22.070 173.135 ;
        RECT 22.770 173.085 23.030 173.135 ;
        RECT 23.730 173.085 23.990 173.135 ;
        RECT 24.690 173.085 24.950 173.135 ;
        RECT 11.165 172.825 29.230 173.085 ;
        RECT 12.285 172.775 12.545 172.825 ;
        RECT 13.250 172.775 13.510 172.825 ;
        RECT 14.205 172.775 14.465 172.825 ;
        RECT 15.165 172.775 15.425 172.825 ;
        RECT 16.125 172.775 16.385 172.825 ;
        RECT 17.085 172.775 17.345 172.825 ;
        RECT 18.405 169.890 18.665 172.825 ;
        RECT 19.890 172.775 20.150 172.825 ;
        RECT 20.855 172.775 21.115 172.825 ;
        RECT 21.810 172.775 22.070 172.825 ;
        RECT 22.770 172.775 23.030 172.825 ;
        RECT 23.730 172.775 23.990 172.825 ;
        RECT 24.690 172.775 24.950 172.825 ;
        RECT 27.240 170.405 27.510 170.425 ;
        RECT 28.040 170.405 28.300 172.825 ;
        RECT 27.240 170.145 28.300 170.405 ;
        RECT 27.240 170.055 27.510 170.145 ;
    END
  END en_b[5]
  PIN en_b[6]
    DIRECTION INOUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 4.402500 ;
    PORT
      LAYER li1 ;
        RECT 12.250 166.430 12.580 166.600 ;
        RECT 13.210 166.430 13.540 166.600 ;
        RECT 14.170 166.430 14.500 166.600 ;
        RECT 15.130 166.430 15.460 166.600 ;
        RECT 16.090 166.430 16.420 166.600 ;
        RECT 17.050 166.430 17.380 166.600 ;
        RECT 19.855 166.430 20.185 166.600 ;
        RECT 20.815 166.430 21.145 166.600 ;
        RECT 21.775 166.430 22.105 166.600 ;
        RECT 22.735 166.430 23.065 166.600 ;
        RECT 23.695 166.430 24.025 166.600 ;
        RECT 24.655 166.430 24.985 166.600 ;
        RECT 27.100 163.715 27.430 163.955 ;
        RECT 18.375 163.500 18.705 163.670 ;
      LAYER mcon ;
        RECT 12.330 166.430 12.500 166.600 ;
        RECT 13.290 166.430 13.460 166.600 ;
        RECT 14.250 166.430 14.420 166.600 ;
        RECT 15.210 166.430 15.380 166.600 ;
        RECT 16.170 166.430 16.340 166.600 ;
        RECT 17.130 166.430 17.300 166.600 ;
        RECT 19.935 166.430 20.105 166.600 ;
        RECT 20.895 166.430 21.065 166.600 ;
        RECT 21.855 166.430 22.025 166.600 ;
        RECT 22.815 166.430 22.985 166.600 ;
        RECT 23.775 166.430 23.945 166.600 ;
        RECT 24.735 166.430 24.905 166.600 ;
        RECT 27.250 163.730 27.420 163.900 ;
        RECT 18.455 163.500 18.625 163.670 ;
      LAYER met1 ;
        RECT 12.235 166.390 12.595 166.650 ;
        RECT 13.200 166.390 13.560 166.650 ;
        RECT 14.155 166.390 14.515 166.650 ;
        RECT 15.115 166.390 15.475 166.650 ;
        RECT 16.075 166.390 16.435 166.650 ;
        RECT 17.035 166.390 17.395 166.650 ;
        RECT 19.840 166.390 20.200 166.650 ;
        RECT 20.805 166.390 21.165 166.650 ;
        RECT 21.760 166.390 22.120 166.650 ;
        RECT 22.720 166.390 23.080 166.650 ;
        RECT 23.680 166.390 24.040 166.650 ;
        RECT 24.640 166.390 25.000 166.650 ;
        RECT 18.355 163.505 18.715 163.765 ;
        RECT 27.190 163.670 27.560 163.940 ;
        RECT 18.395 163.470 18.685 163.505 ;
      LAYER via ;
        RECT 12.285 166.390 12.545 166.650 ;
        RECT 13.250 166.390 13.510 166.650 ;
        RECT 14.205 166.390 14.465 166.650 ;
        RECT 15.165 166.390 15.425 166.650 ;
        RECT 16.125 166.390 16.385 166.650 ;
        RECT 17.085 166.390 17.345 166.650 ;
        RECT 19.890 166.390 20.150 166.650 ;
        RECT 20.855 166.390 21.115 166.650 ;
        RECT 21.810 166.390 22.070 166.650 ;
        RECT 22.770 166.390 23.030 166.650 ;
        RECT 23.730 166.390 23.990 166.650 ;
        RECT 24.690 166.390 24.950 166.650 ;
        RECT 18.405 163.505 18.665 163.765 ;
        RECT 27.245 163.675 27.505 163.935 ;
      LAYER met2 ;
        RECT 12.285 166.650 12.545 166.700 ;
        RECT 13.250 166.650 13.510 166.700 ;
        RECT 14.205 166.650 14.465 166.700 ;
        RECT 15.165 166.650 15.425 166.700 ;
        RECT 16.125 166.650 16.385 166.700 ;
        RECT 17.085 166.650 17.345 166.700 ;
        RECT 19.890 166.650 20.150 166.700 ;
        RECT 20.855 166.650 21.115 166.700 ;
        RECT 21.810 166.650 22.070 166.700 ;
        RECT 22.770 166.650 23.030 166.700 ;
        RECT 23.730 166.650 23.990 166.700 ;
        RECT 24.690 166.650 24.950 166.700 ;
        RECT 11.165 166.390 29.230 166.650 ;
        RECT 12.285 166.340 12.545 166.390 ;
        RECT 13.250 166.340 13.510 166.390 ;
        RECT 14.205 166.340 14.465 166.390 ;
        RECT 15.165 166.340 15.425 166.390 ;
        RECT 16.125 166.340 16.385 166.390 ;
        RECT 17.085 166.340 17.345 166.390 ;
        RECT 18.405 163.455 18.665 166.390 ;
        RECT 19.890 166.340 20.150 166.390 ;
        RECT 20.855 166.340 21.115 166.390 ;
        RECT 21.810 166.340 22.070 166.390 ;
        RECT 22.770 166.340 23.030 166.390 ;
        RECT 23.730 166.340 23.990 166.390 ;
        RECT 24.690 166.340 24.950 166.390 ;
        RECT 27.240 163.970 27.510 163.990 ;
        RECT 28.040 163.970 28.300 166.390 ;
        RECT 27.240 163.710 28.300 163.970 ;
        RECT 27.240 163.620 27.510 163.710 ;
    END
  END en_b[6]
  PIN en_b[7]
    DIRECTION INOUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 4.402500 ;
    PORT
      LAYER li1 ;
        RECT 12.250 159.995 12.580 160.165 ;
        RECT 13.210 159.995 13.540 160.165 ;
        RECT 14.170 159.995 14.500 160.165 ;
        RECT 15.130 159.995 15.460 160.165 ;
        RECT 16.090 159.995 16.420 160.165 ;
        RECT 17.050 159.995 17.380 160.165 ;
        RECT 19.855 159.995 20.185 160.165 ;
        RECT 20.815 159.995 21.145 160.165 ;
        RECT 21.775 159.995 22.105 160.165 ;
        RECT 22.735 159.995 23.065 160.165 ;
        RECT 23.695 159.995 24.025 160.165 ;
        RECT 24.655 159.995 24.985 160.165 ;
        RECT 27.100 157.280 27.430 157.520 ;
        RECT 18.375 157.065 18.705 157.235 ;
      LAYER mcon ;
        RECT 12.330 159.995 12.500 160.165 ;
        RECT 13.290 159.995 13.460 160.165 ;
        RECT 14.250 159.995 14.420 160.165 ;
        RECT 15.210 159.995 15.380 160.165 ;
        RECT 16.170 159.995 16.340 160.165 ;
        RECT 17.130 159.995 17.300 160.165 ;
        RECT 19.935 159.995 20.105 160.165 ;
        RECT 20.895 159.995 21.065 160.165 ;
        RECT 21.855 159.995 22.025 160.165 ;
        RECT 22.815 159.995 22.985 160.165 ;
        RECT 23.775 159.995 23.945 160.165 ;
        RECT 24.735 159.995 24.905 160.165 ;
        RECT 27.250 157.295 27.420 157.465 ;
        RECT 18.455 157.065 18.625 157.235 ;
      LAYER met1 ;
        RECT 12.235 159.955 12.595 160.215 ;
        RECT 13.200 159.955 13.560 160.215 ;
        RECT 14.155 159.955 14.515 160.215 ;
        RECT 15.115 159.955 15.475 160.215 ;
        RECT 16.075 159.955 16.435 160.215 ;
        RECT 17.035 159.955 17.395 160.215 ;
        RECT 19.840 159.955 20.200 160.215 ;
        RECT 20.805 159.955 21.165 160.215 ;
        RECT 21.760 159.955 22.120 160.215 ;
        RECT 22.720 159.955 23.080 160.215 ;
        RECT 23.680 159.955 24.040 160.215 ;
        RECT 24.640 159.955 25.000 160.215 ;
        RECT 18.355 157.070 18.715 157.330 ;
        RECT 27.190 157.235 27.560 157.505 ;
        RECT 18.395 157.035 18.685 157.070 ;
      LAYER via ;
        RECT 12.285 159.955 12.545 160.215 ;
        RECT 13.250 159.955 13.510 160.215 ;
        RECT 14.205 159.955 14.465 160.215 ;
        RECT 15.165 159.955 15.425 160.215 ;
        RECT 16.125 159.955 16.385 160.215 ;
        RECT 17.085 159.955 17.345 160.215 ;
        RECT 19.890 159.955 20.150 160.215 ;
        RECT 20.855 159.955 21.115 160.215 ;
        RECT 21.810 159.955 22.070 160.215 ;
        RECT 22.770 159.955 23.030 160.215 ;
        RECT 23.730 159.955 23.990 160.215 ;
        RECT 24.690 159.955 24.950 160.215 ;
        RECT 18.405 157.070 18.665 157.330 ;
        RECT 27.245 157.240 27.505 157.500 ;
      LAYER met2 ;
        RECT 12.285 160.215 12.545 160.265 ;
        RECT 13.250 160.215 13.510 160.265 ;
        RECT 14.205 160.215 14.465 160.265 ;
        RECT 15.165 160.215 15.425 160.265 ;
        RECT 16.125 160.215 16.385 160.265 ;
        RECT 17.085 160.215 17.345 160.265 ;
        RECT 19.890 160.215 20.150 160.265 ;
        RECT 20.855 160.215 21.115 160.265 ;
        RECT 21.810 160.215 22.070 160.265 ;
        RECT 22.770 160.215 23.030 160.265 ;
        RECT 23.730 160.215 23.990 160.265 ;
        RECT 24.690 160.215 24.950 160.265 ;
        RECT 11.165 159.955 29.230 160.215 ;
        RECT 12.285 159.905 12.545 159.955 ;
        RECT 13.250 159.905 13.510 159.955 ;
        RECT 14.205 159.905 14.465 159.955 ;
        RECT 15.165 159.905 15.425 159.955 ;
        RECT 16.125 159.905 16.385 159.955 ;
        RECT 17.085 159.905 17.345 159.955 ;
        RECT 18.405 157.020 18.665 159.955 ;
        RECT 19.890 159.905 20.150 159.955 ;
        RECT 20.855 159.905 21.115 159.955 ;
        RECT 21.810 159.905 22.070 159.955 ;
        RECT 22.770 159.905 23.030 159.955 ;
        RECT 23.730 159.905 23.990 159.955 ;
        RECT 24.690 159.905 24.950 159.955 ;
        RECT 27.240 157.535 27.510 157.555 ;
        RECT 28.040 157.535 28.300 159.955 ;
        RECT 27.240 157.275 28.300 157.535 ;
        RECT 27.240 157.185 27.510 157.275 ;
    END
  END en_b[7]
  PIN en_b[8]
    DIRECTION INOUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 4.402500 ;
    PORT
      LAYER li1 ;
        RECT 12.250 153.560 12.580 153.730 ;
        RECT 13.210 153.560 13.540 153.730 ;
        RECT 14.170 153.560 14.500 153.730 ;
        RECT 15.130 153.560 15.460 153.730 ;
        RECT 16.090 153.560 16.420 153.730 ;
        RECT 17.050 153.560 17.380 153.730 ;
        RECT 19.855 153.560 20.185 153.730 ;
        RECT 20.815 153.560 21.145 153.730 ;
        RECT 21.775 153.560 22.105 153.730 ;
        RECT 22.735 153.560 23.065 153.730 ;
        RECT 23.695 153.560 24.025 153.730 ;
        RECT 24.655 153.560 24.985 153.730 ;
        RECT 27.100 150.845 27.430 151.085 ;
        RECT 18.375 150.630 18.705 150.800 ;
      LAYER mcon ;
        RECT 12.330 153.560 12.500 153.730 ;
        RECT 13.290 153.560 13.460 153.730 ;
        RECT 14.250 153.560 14.420 153.730 ;
        RECT 15.210 153.560 15.380 153.730 ;
        RECT 16.170 153.560 16.340 153.730 ;
        RECT 17.130 153.560 17.300 153.730 ;
        RECT 19.935 153.560 20.105 153.730 ;
        RECT 20.895 153.560 21.065 153.730 ;
        RECT 21.855 153.560 22.025 153.730 ;
        RECT 22.815 153.560 22.985 153.730 ;
        RECT 23.775 153.560 23.945 153.730 ;
        RECT 24.735 153.560 24.905 153.730 ;
        RECT 27.250 150.860 27.420 151.030 ;
        RECT 18.455 150.630 18.625 150.800 ;
      LAYER met1 ;
        RECT 12.235 153.520 12.595 153.780 ;
        RECT 13.200 153.520 13.560 153.780 ;
        RECT 14.155 153.520 14.515 153.780 ;
        RECT 15.115 153.520 15.475 153.780 ;
        RECT 16.075 153.520 16.435 153.780 ;
        RECT 17.035 153.520 17.395 153.780 ;
        RECT 19.840 153.520 20.200 153.780 ;
        RECT 20.805 153.520 21.165 153.780 ;
        RECT 21.760 153.520 22.120 153.780 ;
        RECT 22.720 153.520 23.080 153.780 ;
        RECT 23.680 153.520 24.040 153.780 ;
        RECT 24.640 153.520 25.000 153.780 ;
        RECT 18.355 150.635 18.715 150.895 ;
        RECT 27.190 150.800 27.560 151.070 ;
        RECT 18.395 150.600 18.685 150.635 ;
      LAYER via ;
        RECT 12.285 153.520 12.545 153.780 ;
        RECT 13.250 153.520 13.510 153.780 ;
        RECT 14.205 153.520 14.465 153.780 ;
        RECT 15.165 153.520 15.425 153.780 ;
        RECT 16.125 153.520 16.385 153.780 ;
        RECT 17.085 153.520 17.345 153.780 ;
        RECT 19.890 153.520 20.150 153.780 ;
        RECT 20.855 153.520 21.115 153.780 ;
        RECT 21.810 153.520 22.070 153.780 ;
        RECT 22.770 153.520 23.030 153.780 ;
        RECT 23.730 153.520 23.990 153.780 ;
        RECT 24.690 153.520 24.950 153.780 ;
        RECT 18.405 150.635 18.665 150.895 ;
        RECT 27.245 150.805 27.505 151.065 ;
      LAYER met2 ;
        RECT 12.285 153.780 12.545 153.830 ;
        RECT 13.250 153.780 13.510 153.830 ;
        RECT 14.205 153.780 14.465 153.830 ;
        RECT 15.165 153.780 15.425 153.830 ;
        RECT 16.125 153.780 16.385 153.830 ;
        RECT 17.085 153.780 17.345 153.830 ;
        RECT 19.890 153.780 20.150 153.830 ;
        RECT 20.855 153.780 21.115 153.830 ;
        RECT 21.810 153.780 22.070 153.830 ;
        RECT 22.770 153.780 23.030 153.830 ;
        RECT 23.730 153.780 23.990 153.830 ;
        RECT 24.690 153.780 24.950 153.830 ;
        RECT 11.165 153.520 29.230 153.780 ;
        RECT 12.285 153.470 12.545 153.520 ;
        RECT 13.250 153.470 13.510 153.520 ;
        RECT 14.205 153.470 14.465 153.520 ;
        RECT 15.165 153.470 15.425 153.520 ;
        RECT 16.125 153.470 16.385 153.520 ;
        RECT 17.085 153.470 17.345 153.520 ;
        RECT 18.405 150.585 18.665 153.520 ;
        RECT 19.890 153.470 20.150 153.520 ;
        RECT 20.855 153.470 21.115 153.520 ;
        RECT 21.810 153.470 22.070 153.520 ;
        RECT 22.770 153.470 23.030 153.520 ;
        RECT 23.730 153.470 23.990 153.520 ;
        RECT 24.690 153.470 24.950 153.520 ;
        RECT 27.240 151.100 27.510 151.120 ;
        RECT 28.040 151.100 28.300 153.520 ;
        RECT 27.240 150.840 28.300 151.100 ;
        RECT 27.240 150.750 27.510 150.840 ;
    END
  END en_b[8]
  PIN en_b[9]
    DIRECTION INOUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 4.402500 ;
    PORT
      LAYER li1 ;
        RECT 12.250 147.125 12.580 147.295 ;
        RECT 13.210 147.125 13.540 147.295 ;
        RECT 14.170 147.125 14.500 147.295 ;
        RECT 15.130 147.125 15.460 147.295 ;
        RECT 16.090 147.125 16.420 147.295 ;
        RECT 17.050 147.125 17.380 147.295 ;
        RECT 19.855 147.125 20.185 147.295 ;
        RECT 20.815 147.125 21.145 147.295 ;
        RECT 21.775 147.125 22.105 147.295 ;
        RECT 22.735 147.125 23.065 147.295 ;
        RECT 23.695 147.125 24.025 147.295 ;
        RECT 24.655 147.125 24.985 147.295 ;
        RECT 27.100 144.410 27.430 144.650 ;
        RECT 18.375 144.195 18.705 144.365 ;
      LAYER mcon ;
        RECT 12.330 147.125 12.500 147.295 ;
        RECT 13.290 147.125 13.460 147.295 ;
        RECT 14.250 147.125 14.420 147.295 ;
        RECT 15.210 147.125 15.380 147.295 ;
        RECT 16.170 147.125 16.340 147.295 ;
        RECT 17.130 147.125 17.300 147.295 ;
        RECT 19.935 147.125 20.105 147.295 ;
        RECT 20.895 147.125 21.065 147.295 ;
        RECT 21.855 147.125 22.025 147.295 ;
        RECT 22.815 147.125 22.985 147.295 ;
        RECT 23.775 147.125 23.945 147.295 ;
        RECT 24.735 147.125 24.905 147.295 ;
        RECT 27.250 144.425 27.420 144.595 ;
        RECT 18.455 144.195 18.625 144.365 ;
      LAYER met1 ;
        RECT 12.235 147.085 12.595 147.345 ;
        RECT 13.200 147.085 13.560 147.345 ;
        RECT 14.155 147.085 14.515 147.345 ;
        RECT 15.115 147.085 15.475 147.345 ;
        RECT 16.075 147.085 16.435 147.345 ;
        RECT 17.035 147.085 17.395 147.345 ;
        RECT 19.840 147.085 20.200 147.345 ;
        RECT 20.805 147.085 21.165 147.345 ;
        RECT 21.760 147.085 22.120 147.345 ;
        RECT 22.720 147.085 23.080 147.345 ;
        RECT 23.680 147.085 24.040 147.345 ;
        RECT 24.640 147.085 25.000 147.345 ;
        RECT 18.355 144.200 18.715 144.460 ;
        RECT 27.190 144.365 27.560 144.635 ;
        RECT 18.395 144.165 18.685 144.200 ;
      LAYER via ;
        RECT 12.285 147.085 12.545 147.345 ;
        RECT 13.250 147.085 13.510 147.345 ;
        RECT 14.205 147.085 14.465 147.345 ;
        RECT 15.165 147.085 15.425 147.345 ;
        RECT 16.125 147.085 16.385 147.345 ;
        RECT 17.085 147.085 17.345 147.345 ;
        RECT 19.890 147.085 20.150 147.345 ;
        RECT 20.855 147.085 21.115 147.345 ;
        RECT 21.810 147.085 22.070 147.345 ;
        RECT 22.770 147.085 23.030 147.345 ;
        RECT 23.730 147.085 23.990 147.345 ;
        RECT 24.690 147.085 24.950 147.345 ;
        RECT 18.405 144.200 18.665 144.460 ;
        RECT 27.245 144.370 27.505 144.630 ;
      LAYER met2 ;
        RECT 12.285 147.345 12.545 147.395 ;
        RECT 13.250 147.345 13.510 147.395 ;
        RECT 14.205 147.345 14.465 147.395 ;
        RECT 15.165 147.345 15.425 147.395 ;
        RECT 16.125 147.345 16.385 147.395 ;
        RECT 17.085 147.345 17.345 147.395 ;
        RECT 19.890 147.345 20.150 147.395 ;
        RECT 20.855 147.345 21.115 147.395 ;
        RECT 21.810 147.345 22.070 147.395 ;
        RECT 22.770 147.345 23.030 147.395 ;
        RECT 23.730 147.345 23.990 147.395 ;
        RECT 24.690 147.345 24.950 147.395 ;
        RECT 11.165 147.085 29.230 147.345 ;
        RECT 12.285 147.035 12.545 147.085 ;
        RECT 13.250 147.035 13.510 147.085 ;
        RECT 14.205 147.035 14.465 147.085 ;
        RECT 15.165 147.035 15.425 147.085 ;
        RECT 16.125 147.035 16.385 147.085 ;
        RECT 17.085 147.035 17.345 147.085 ;
        RECT 18.405 144.150 18.665 147.085 ;
        RECT 19.890 147.035 20.150 147.085 ;
        RECT 20.855 147.035 21.115 147.085 ;
        RECT 21.810 147.035 22.070 147.085 ;
        RECT 22.770 147.035 23.030 147.085 ;
        RECT 23.730 147.035 23.990 147.085 ;
        RECT 24.690 147.035 24.950 147.085 ;
        RECT 27.240 144.665 27.510 144.685 ;
        RECT 28.040 144.665 28.300 147.085 ;
        RECT 27.240 144.405 28.300 144.665 ;
        RECT 27.240 144.315 27.510 144.405 ;
    END
  END en_b[9]
  PIN en_b[10]
    DIRECTION INOUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 4.402500 ;
    PORT
      LAYER li1 ;
        RECT 12.250 140.690 12.580 140.860 ;
        RECT 13.210 140.690 13.540 140.860 ;
        RECT 14.170 140.690 14.500 140.860 ;
        RECT 15.130 140.690 15.460 140.860 ;
        RECT 16.090 140.690 16.420 140.860 ;
        RECT 17.050 140.690 17.380 140.860 ;
        RECT 19.855 140.690 20.185 140.860 ;
        RECT 20.815 140.690 21.145 140.860 ;
        RECT 21.775 140.690 22.105 140.860 ;
        RECT 22.735 140.690 23.065 140.860 ;
        RECT 23.695 140.690 24.025 140.860 ;
        RECT 24.655 140.690 24.985 140.860 ;
        RECT 27.100 137.975 27.430 138.215 ;
        RECT 18.375 137.760 18.705 137.930 ;
      LAYER mcon ;
        RECT 12.330 140.690 12.500 140.860 ;
        RECT 13.290 140.690 13.460 140.860 ;
        RECT 14.250 140.690 14.420 140.860 ;
        RECT 15.210 140.690 15.380 140.860 ;
        RECT 16.170 140.690 16.340 140.860 ;
        RECT 17.130 140.690 17.300 140.860 ;
        RECT 19.935 140.690 20.105 140.860 ;
        RECT 20.895 140.690 21.065 140.860 ;
        RECT 21.855 140.690 22.025 140.860 ;
        RECT 22.815 140.690 22.985 140.860 ;
        RECT 23.775 140.690 23.945 140.860 ;
        RECT 24.735 140.690 24.905 140.860 ;
        RECT 27.250 137.990 27.420 138.160 ;
        RECT 18.455 137.760 18.625 137.930 ;
      LAYER met1 ;
        RECT 12.235 140.650 12.595 140.910 ;
        RECT 13.200 140.650 13.560 140.910 ;
        RECT 14.155 140.650 14.515 140.910 ;
        RECT 15.115 140.650 15.475 140.910 ;
        RECT 16.075 140.650 16.435 140.910 ;
        RECT 17.035 140.650 17.395 140.910 ;
        RECT 19.840 140.650 20.200 140.910 ;
        RECT 20.805 140.650 21.165 140.910 ;
        RECT 21.760 140.650 22.120 140.910 ;
        RECT 22.720 140.650 23.080 140.910 ;
        RECT 23.680 140.650 24.040 140.910 ;
        RECT 24.640 140.650 25.000 140.910 ;
        RECT 18.355 137.765 18.715 138.025 ;
        RECT 27.190 137.930 27.560 138.200 ;
        RECT 18.395 137.730 18.685 137.765 ;
      LAYER via ;
        RECT 12.285 140.650 12.545 140.910 ;
        RECT 13.250 140.650 13.510 140.910 ;
        RECT 14.205 140.650 14.465 140.910 ;
        RECT 15.165 140.650 15.425 140.910 ;
        RECT 16.125 140.650 16.385 140.910 ;
        RECT 17.085 140.650 17.345 140.910 ;
        RECT 19.890 140.650 20.150 140.910 ;
        RECT 20.855 140.650 21.115 140.910 ;
        RECT 21.810 140.650 22.070 140.910 ;
        RECT 22.770 140.650 23.030 140.910 ;
        RECT 23.730 140.650 23.990 140.910 ;
        RECT 24.690 140.650 24.950 140.910 ;
        RECT 18.405 137.765 18.665 138.025 ;
        RECT 27.245 137.935 27.505 138.195 ;
      LAYER met2 ;
        RECT 12.285 140.910 12.545 140.960 ;
        RECT 13.250 140.910 13.510 140.960 ;
        RECT 14.205 140.910 14.465 140.960 ;
        RECT 15.165 140.910 15.425 140.960 ;
        RECT 16.125 140.910 16.385 140.960 ;
        RECT 17.085 140.910 17.345 140.960 ;
        RECT 19.890 140.910 20.150 140.960 ;
        RECT 20.855 140.910 21.115 140.960 ;
        RECT 21.810 140.910 22.070 140.960 ;
        RECT 22.770 140.910 23.030 140.960 ;
        RECT 23.730 140.910 23.990 140.960 ;
        RECT 24.690 140.910 24.950 140.960 ;
        RECT 11.165 140.650 29.230 140.910 ;
        RECT 12.285 140.600 12.545 140.650 ;
        RECT 13.250 140.600 13.510 140.650 ;
        RECT 14.205 140.600 14.465 140.650 ;
        RECT 15.165 140.600 15.425 140.650 ;
        RECT 16.125 140.600 16.385 140.650 ;
        RECT 17.085 140.600 17.345 140.650 ;
        RECT 18.405 137.715 18.665 140.650 ;
        RECT 19.890 140.600 20.150 140.650 ;
        RECT 20.855 140.600 21.115 140.650 ;
        RECT 21.810 140.600 22.070 140.650 ;
        RECT 22.770 140.600 23.030 140.650 ;
        RECT 23.730 140.600 23.990 140.650 ;
        RECT 24.690 140.600 24.950 140.650 ;
        RECT 27.240 138.230 27.510 138.250 ;
        RECT 28.040 138.230 28.300 140.650 ;
        RECT 27.240 137.970 28.300 138.230 ;
        RECT 27.240 137.880 27.510 137.970 ;
    END
  END en_b[10]
  PIN en_b[11]
    DIRECTION INOUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 4.402500 ;
    PORT
      LAYER li1 ;
        RECT 12.250 134.255 12.580 134.425 ;
        RECT 13.210 134.255 13.540 134.425 ;
        RECT 14.170 134.255 14.500 134.425 ;
        RECT 15.130 134.255 15.460 134.425 ;
        RECT 16.090 134.255 16.420 134.425 ;
        RECT 17.050 134.255 17.380 134.425 ;
        RECT 19.855 134.255 20.185 134.425 ;
        RECT 20.815 134.255 21.145 134.425 ;
        RECT 21.775 134.255 22.105 134.425 ;
        RECT 22.735 134.255 23.065 134.425 ;
        RECT 23.695 134.255 24.025 134.425 ;
        RECT 24.655 134.255 24.985 134.425 ;
        RECT 27.100 131.540 27.430 131.780 ;
        RECT 18.375 131.325 18.705 131.495 ;
      LAYER mcon ;
        RECT 12.330 134.255 12.500 134.425 ;
        RECT 13.290 134.255 13.460 134.425 ;
        RECT 14.250 134.255 14.420 134.425 ;
        RECT 15.210 134.255 15.380 134.425 ;
        RECT 16.170 134.255 16.340 134.425 ;
        RECT 17.130 134.255 17.300 134.425 ;
        RECT 19.935 134.255 20.105 134.425 ;
        RECT 20.895 134.255 21.065 134.425 ;
        RECT 21.855 134.255 22.025 134.425 ;
        RECT 22.815 134.255 22.985 134.425 ;
        RECT 23.775 134.255 23.945 134.425 ;
        RECT 24.735 134.255 24.905 134.425 ;
        RECT 27.250 131.555 27.420 131.725 ;
        RECT 18.455 131.325 18.625 131.495 ;
      LAYER met1 ;
        RECT 12.235 134.215 12.595 134.475 ;
        RECT 13.200 134.215 13.560 134.475 ;
        RECT 14.155 134.215 14.515 134.475 ;
        RECT 15.115 134.215 15.475 134.475 ;
        RECT 16.075 134.215 16.435 134.475 ;
        RECT 17.035 134.215 17.395 134.475 ;
        RECT 19.840 134.215 20.200 134.475 ;
        RECT 20.805 134.215 21.165 134.475 ;
        RECT 21.760 134.215 22.120 134.475 ;
        RECT 22.720 134.215 23.080 134.475 ;
        RECT 23.680 134.215 24.040 134.475 ;
        RECT 24.640 134.215 25.000 134.475 ;
        RECT 18.355 131.330 18.715 131.590 ;
        RECT 27.190 131.495 27.560 131.765 ;
        RECT 18.395 131.295 18.685 131.330 ;
      LAYER via ;
        RECT 12.285 134.215 12.545 134.475 ;
        RECT 13.250 134.215 13.510 134.475 ;
        RECT 14.205 134.215 14.465 134.475 ;
        RECT 15.165 134.215 15.425 134.475 ;
        RECT 16.125 134.215 16.385 134.475 ;
        RECT 17.085 134.215 17.345 134.475 ;
        RECT 19.890 134.215 20.150 134.475 ;
        RECT 20.855 134.215 21.115 134.475 ;
        RECT 21.810 134.215 22.070 134.475 ;
        RECT 22.770 134.215 23.030 134.475 ;
        RECT 23.730 134.215 23.990 134.475 ;
        RECT 24.690 134.215 24.950 134.475 ;
        RECT 18.405 131.330 18.665 131.590 ;
        RECT 27.245 131.500 27.505 131.760 ;
      LAYER met2 ;
        RECT 12.285 134.475 12.545 134.525 ;
        RECT 13.250 134.475 13.510 134.525 ;
        RECT 14.205 134.475 14.465 134.525 ;
        RECT 15.165 134.475 15.425 134.525 ;
        RECT 16.125 134.475 16.385 134.525 ;
        RECT 17.085 134.475 17.345 134.525 ;
        RECT 19.890 134.475 20.150 134.525 ;
        RECT 20.855 134.475 21.115 134.525 ;
        RECT 21.810 134.475 22.070 134.525 ;
        RECT 22.770 134.475 23.030 134.525 ;
        RECT 23.730 134.475 23.990 134.525 ;
        RECT 24.690 134.475 24.950 134.525 ;
        RECT 11.165 134.215 29.230 134.475 ;
        RECT 12.285 134.165 12.545 134.215 ;
        RECT 13.250 134.165 13.510 134.215 ;
        RECT 14.205 134.165 14.465 134.215 ;
        RECT 15.165 134.165 15.425 134.215 ;
        RECT 16.125 134.165 16.385 134.215 ;
        RECT 17.085 134.165 17.345 134.215 ;
        RECT 18.405 131.280 18.665 134.215 ;
        RECT 19.890 134.165 20.150 134.215 ;
        RECT 20.855 134.165 21.115 134.215 ;
        RECT 21.810 134.165 22.070 134.215 ;
        RECT 22.770 134.165 23.030 134.215 ;
        RECT 23.730 134.165 23.990 134.215 ;
        RECT 24.690 134.165 24.950 134.215 ;
        RECT 27.240 131.795 27.510 131.815 ;
        RECT 28.040 131.795 28.300 134.215 ;
        RECT 27.240 131.535 28.300 131.795 ;
        RECT 27.240 131.445 27.510 131.535 ;
    END
  END en_b[11]
  PIN en_b[12]
    DIRECTION INOUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 4.402500 ;
    PORT
      LAYER li1 ;
        RECT 12.250 127.820 12.580 127.990 ;
        RECT 13.210 127.820 13.540 127.990 ;
        RECT 14.170 127.820 14.500 127.990 ;
        RECT 15.130 127.820 15.460 127.990 ;
        RECT 16.090 127.820 16.420 127.990 ;
        RECT 17.050 127.820 17.380 127.990 ;
        RECT 19.855 127.820 20.185 127.990 ;
        RECT 20.815 127.820 21.145 127.990 ;
        RECT 21.775 127.820 22.105 127.990 ;
        RECT 22.735 127.820 23.065 127.990 ;
        RECT 23.695 127.820 24.025 127.990 ;
        RECT 24.655 127.820 24.985 127.990 ;
        RECT 27.100 125.105 27.430 125.345 ;
        RECT 18.375 124.890 18.705 125.060 ;
      LAYER mcon ;
        RECT 12.330 127.820 12.500 127.990 ;
        RECT 13.290 127.820 13.460 127.990 ;
        RECT 14.250 127.820 14.420 127.990 ;
        RECT 15.210 127.820 15.380 127.990 ;
        RECT 16.170 127.820 16.340 127.990 ;
        RECT 17.130 127.820 17.300 127.990 ;
        RECT 19.935 127.820 20.105 127.990 ;
        RECT 20.895 127.820 21.065 127.990 ;
        RECT 21.855 127.820 22.025 127.990 ;
        RECT 22.815 127.820 22.985 127.990 ;
        RECT 23.775 127.820 23.945 127.990 ;
        RECT 24.735 127.820 24.905 127.990 ;
        RECT 27.250 125.120 27.420 125.290 ;
        RECT 18.455 124.890 18.625 125.060 ;
      LAYER met1 ;
        RECT 12.235 127.780 12.595 128.040 ;
        RECT 13.200 127.780 13.560 128.040 ;
        RECT 14.155 127.780 14.515 128.040 ;
        RECT 15.115 127.780 15.475 128.040 ;
        RECT 16.075 127.780 16.435 128.040 ;
        RECT 17.035 127.780 17.395 128.040 ;
        RECT 19.840 127.780 20.200 128.040 ;
        RECT 20.805 127.780 21.165 128.040 ;
        RECT 21.760 127.780 22.120 128.040 ;
        RECT 22.720 127.780 23.080 128.040 ;
        RECT 23.680 127.780 24.040 128.040 ;
        RECT 24.640 127.780 25.000 128.040 ;
        RECT 18.355 124.895 18.715 125.155 ;
        RECT 27.190 125.060 27.560 125.330 ;
        RECT 18.395 124.860 18.685 124.895 ;
      LAYER via ;
        RECT 12.285 127.780 12.545 128.040 ;
        RECT 13.250 127.780 13.510 128.040 ;
        RECT 14.205 127.780 14.465 128.040 ;
        RECT 15.165 127.780 15.425 128.040 ;
        RECT 16.125 127.780 16.385 128.040 ;
        RECT 17.085 127.780 17.345 128.040 ;
        RECT 19.890 127.780 20.150 128.040 ;
        RECT 20.855 127.780 21.115 128.040 ;
        RECT 21.810 127.780 22.070 128.040 ;
        RECT 22.770 127.780 23.030 128.040 ;
        RECT 23.730 127.780 23.990 128.040 ;
        RECT 24.690 127.780 24.950 128.040 ;
        RECT 18.405 124.895 18.665 125.155 ;
        RECT 27.245 125.065 27.505 125.325 ;
      LAYER met2 ;
        RECT 12.285 128.040 12.545 128.090 ;
        RECT 13.250 128.040 13.510 128.090 ;
        RECT 14.205 128.040 14.465 128.090 ;
        RECT 15.165 128.040 15.425 128.090 ;
        RECT 16.125 128.040 16.385 128.090 ;
        RECT 17.085 128.040 17.345 128.090 ;
        RECT 19.890 128.040 20.150 128.090 ;
        RECT 20.855 128.040 21.115 128.090 ;
        RECT 21.810 128.040 22.070 128.090 ;
        RECT 22.770 128.040 23.030 128.090 ;
        RECT 23.730 128.040 23.990 128.090 ;
        RECT 24.690 128.040 24.950 128.090 ;
        RECT 11.165 127.780 29.230 128.040 ;
        RECT 12.285 127.730 12.545 127.780 ;
        RECT 13.250 127.730 13.510 127.780 ;
        RECT 14.205 127.730 14.465 127.780 ;
        RECT 15.165 127.730 15.425 127.780 ;
        RECT 16.125 127.730 16.385 127.780 ;
        RECT 17.085 127.730 17.345 127.780 ;
        RECT 18.405 124.845 18.665 127.780 ;
        RECT 19.890 127.730 20.150 127.780 ;
        RECT 20.855 127.730 21.115 127.780 ;
        RECT 21.810 127.730 22.070 127.780 ;
        RECT 22.770 127.730 23.030 127.780 ;
        RECT 23.730 127.730 23.990 127.780 ;
        RECT 24.690 127.730 24.950 127.780 ;
        RECT 27.240 125.360 27.510 125.380 ;
        RECT 28.040 125.360 28.300 127.780 ;
        RECT 27.240 125.100 28.300 125.360 ;
        RECT 27.240 125.010 27.510 125.100 ;
    END
  END en_b[12]
  PIN en_b[13]
    DIRECTION INOUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 4.402500 ;
    PORT
      LAYER li1 ;
        RECT 12.250 121.385 12.580 121.555 ;
        RECT 13.210 121.385 13.540 121.555 ;
        RECT 14.170 121.385 14.500 121.555 ;
        RECT 15.130 121.385 15.460 121.555 ;
        RECT 16.090 121.385 16.420 121.555 ;
        RECT 17.050 121.385 17.380 121.555 ;
        RECT 19.855 121.385 20.185 121.555 ;
        RECT 20.815 121.385 21.145 121.555 ;
        RECT 21.775 121.385 22.105 121.555 ;
        RECT 22.735 121.385 23.065 121.555 ;
        RECT 23.695 121.385 24.025 121.555 ;
        RECT 24.655 121.385 24.985 121.555 ;
        RECT 27.100 118.670 27.430 118.910 ;
        RECT 18.375 118.455 18.705 118.625 ;
      LAYER mcon ;
        RECT 12.330 121.385 12.500 121.555 ;
        RECT 13.290 121.385 13.460 121.555 ;
        RECT 14.250 121.385 14.420 121.555 ;
        RECT 15.210 121.385 15.380 121.555 ;
        RECT 16.170 121.385 16.340 121.555 ;
        RECT 17.130 121.385 17.300 121.555 ;
        RECT 19.935 121.385 20.105 121.555 ;
        RECT 20.895 121.385 21.065 121.555 ;
        RECT 21.855 121.385 22.025 121.555 ;
        RECT 22.815 121.385 22.985 121.555 ;
        RECT 23.775 121.385 23.945 121.555 ;
        RECT 24.735 121.385 24.905 121.555 ;
        RECT 27.250 118.685 27.420 118.855 ;
        RECT 18.455 118.455 18.625 118.625 ;
      LAYER met1 ;
        RECT 12.235 121.345 12.595 121.605 ;
        RECT 13.200 121.345 13.560 121.605 ;
        RECT 14.155 121.345 14.515 121.605 ;
        RECT 15.115 121.345 15.475 121.605 ;
        RECT 16.075 121.345 16.435 121.605 ;
        RECT 17.035 121.345 17.395 121.605 ;
        RECT 19.840 121.345 20.200 121.605 ;
        RECT 20.805 121.345 21.165 121.605 ;
        RECT 21.760 121.345 22.120 121.605 ;
        RECT 22.720 121.345 23.080 121.605 ;
        RECT 23.680 121.345 24.040 121.605 ;
        RECT 24.640 121.345 25.000 121.605 ;
        RECT 18.355 118.460 18.715 118.720 ;
        RECT 27.190 118.625 27.560 118.895 ;
        RECT 18.395 118.425 18.685 118.460 ;
      LAYER via ;
        RECT 12.285 121.345 12.545 121.605 ;
        RECT 13.250 121.345 13.510 121.605 ;
        RECT 14.205 121.345 14.465 121.605 ;
        RECT 15.165 121.345 15.425 121.605 ;
        RECT 16.125 121.345 16.385 121.605 ;
        RECT 17.085 121.345 17.345 121.605 ;
        RECT 19.890 121.345 20.150 121.605 ;
        RECT 20.855 121.345 21.115 121.605 ;
        RECT 21.810 121.345 22.070 121.605 ;
        RECT 22.770 121.345 23.030 121.605 ;
        RECT 23.730 121.345 23.990 121.605 ;
        RECT 24.690 121.345 24.950 121.605 ;
        RECT 18.405 118.460 18.665 118.720 ;
        RECT 27.245 118.630 27.505 118.890 ;
      LAYER met2 ;
        RECT 12.285 121.605 12.545 121.655 ;
        RECT 13.250 121.605 13.510 121.655 ;
        RECT 14.205 121.605 14.465 121.655 ;
        RECT 15.165 121.605 15.425 121.655 ;
        RECT 16.125 121.605 16.385 121.655 ;
        RECT 17.085 121.605 17.345 121.655 ;
        RECT 19.890 121.605 20.150 121.655 ;
        RECT 20.855 121.605 21.115 121.655 ;
        RECT 21.810 121.605 22.070 121.655 ;
        RECT 22.770 121.605 23.030 121.655 ;
        RECT 23.730 121.605 23.990 121.655 ;
        RECT 24.690 121.605 24.950 121.655 ;
        RECT 11.165 121.345 29.230 121.605 ;
        RECT 12.285 121.295 12.545 121.345 ;
        RECT 13.250 121.295 13.510 121.345 ;
        RECT 14.205 121.295 14.465 121.345 ;
        RECT 15.165 121.295 15.425 121.345 ;
        RECT 16.125 121.295 16.385 121.345 ;
        RECT 17.085 121.295 17.345 121.345 ;
        RECT 18.405 118.410 18.665 121.345 ;
        RECT 19.890 121.295 20.150 121.345 ;
        RECT 20.855 121.295 21.115 121.345 ;
        RECT 21.810 121.295 22.070 121.345 ;
        RECT 22.770 121.295 23.030 121.345 ;
        RECT 23.730 121.295 23.990 121.345 ;
        RECT 24.690 121.295 24.950 121.345 ;
        RECT 27.240 118.925 27.510 118.945 ;
        RECT 28.040 118.925 28.300 121.345 ;
        RECT 27.240 118.665 28.300 118.925 ;
        RECT 27.240 118.575 27.510 118.665 ;
    END
  END en_b[13]
  PIN en_b[14]
    DIRECTION INOUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 4.402500 ;
    PORT
      LAYER li1 ;
        RECT 12.250 114.950 12.580 115.120 ;
        RECT 13.210 114.950 13.540 115.120 ;
        RECT 14.170 114.950 14.500 115.120 ;
        RECT 15.130 114.950 15.460 115.120 ;
        RECT 16.090 114.950 16.420 115.120 ;
        RECT 17.050 114.950 17.380 115.120 ;
        RECT 19.855 114.950 20.185 115.120 ;
        RECT 20.815 114.950 21.145 115.120 ;
        RECT 21.775 114.950 22.105 115.120 ;
        RECT 22.735 114.950 23.065 115.120 ;
        RECT 23.695 114.950 24.025 115.120 ;
        RECT 24.655 114.950 24.985 115.120 ;
        RECT 27.100 112.235 27.430 112.475 ;
        RECT 18.375 112.020 18.705 112.190 ;
      LAYER mcon ;
        RECT 12.330 114.950 12.500 115.120 ;
        RECT 13.290 114.950 13.460 115.120 ;
        RECT 14.250 114.950 14.420 115.120 ;
        RECT 15.210 114.950 15.380 115.120 ;
        RECT 16.170 114.950 16.340 115.120 ;
        RECT 17.130 114.950 17.300 115.120 ;
        RECT 19.935 114.950 20.105 115.120 ;
        RECT 20.895 114.950 21.065 115.120 ;
        RECT 21.855 114.950 22.025 115.120 ;
        RECT 22.815 114.950 22.985 115.120 ;
        RECT 23.775 114.950 23.945 115.120 ;
        RECT 24.735 114.950 24.905 115.120 ;
        RECT 27.250 112.250 27.420 112.420 ;
        RECT 18.455 112.020 18.625 112.190 ;
      LAYER met1 ;
        RECT 12.235 114.910 12.595 115.170 ;
        RECT 13.200 114.910 13.560 115.170 ;
        RECT 14.155 114.910 14.515 115.170 ;
        RECT 15.115 114.910 15.475 115.170 ;
        RECT 16.075 114.910 16.435 115.170 ;
        RECT 17.035 114.910 17.395 115.170 ;
        RECT 19.840 114.910 20.200 115.170 ;
        RECT 20.805 114.910 21.165 115.170 ;
        RECT 21.760 114.910 22.120 115.170 ;
        RECT 22.720 114.910 23.080 115.170 ;
        RECT 23.680 114.910 24.040 115.170 ;
        RECT 24.640 114.910 25.000 115.170 ;
        RECT 18.355 112.025 18.715 112.285 ;
        RECT 27.190 112.190 27.560 112.460 ;
        RECT 18.395 111.990 18.685 112.025 ;
      LAYER via ;
        RECT 12.285 114.910 12.545 115.170 ;
        RECT 13.250 114.910 13.510 115.170 ;
        RECT 14.205 114.910 14.465 115.170 ;
        RECT 15.165 114.910 15.425 115.170 ;
        RECT 16.125 114.910 16.385 115.170 ;
        RECT 17.085 114.910 17.345 115.170 ;
        RECT 19.890 114.910 20.150 115.170 ;
        RECT 20.855 114.910 21.115 115.170 ;
        RECT 21.810 114.910 22.070 115.170 ;
        RECT 22.770 114.910 23.030 115.170 ;
        RECT 23.730 114.910 23.990 115.170 ;
        RECT 24.690 114.910 24.950 115.170 ;
        RECT 18.405 112.025 18.665 112.285 ;
        RECT 27.245 112.195 27.505 112.455 ;
      LAYER met2 ;
        RECT 12.285 115.170 12.545 115.220 ;
        RECT 13.250 115.170 13.510 115.220 ;
        RECT 14.205 115.170 14.465 115.220 ;
        RECT 15.165 115.170 15.425 115.220 ;
        RECT 16.125 115.170 16.385 115.220 ;
        RECT 17.085 115.170 17.345 115.220 ;
        RECT 19.890 115.170 20.150 115.220 ;
        RECT 20.855 115.170 21.115 115.220 ;
        RECT 21.810 115.170 22.070 115.220 ;
        RECT 22.770 115.170 23.030 115.220 ;
        RECT 23.730 115.170 23.990 115.220 ;
        RECT 24.690 115.170 24.950 115.220 ;
        RECT 11.165 114.910 29.230 115.170 ;
        RECT 12.285 114.860 12.545 114.910 ;
        RECT 13.250 114.860 13.510 114.910 ;
        RECT 14.205 114.860 14.465 114.910 ;
        RECT 15.165 114.860 15.425 114.910 ;
        RECT 16.125 114.860 16.385 114.910 ;
        RECT 17.085 114.860 17.345 114.910 ;
        RECT 18.405 111.975 18.665 114.910 ;
        RECT 19.890 114.860 20.150 114.910 ;
        RECT 20.855 114.860 21.115 114.910 ;
        RECT 21.810 114.860 22.070 114.910 ;
        RECT 22.770 114.860 23.030 114.910 ;
        RECT 23.730 114.860 23.990 114.910 ;
        RECT 24.690 114.860 24.950 114.910 ;
        RECT 27.240 112.490 27.510 112.510 ;
        RECT 28.040 112.490 28.300 114.910 ;
        RECT 27.240 112.230 28.300 112.490 ;
        RECT 27.240 112.140 27.510 112.230 ;
    END
  END en_b[14]
  PIN en_b[15]
    DIRECTION INOUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 4.402500 ;
    PORT
      LAYER li1 ;
        RECT 12.250 108.515 12.580 108.685 ;
        RECT 13.210 108.515 13.540 108.685 ;
        RECT 14.170 108.515 14.500 108.685 ;
        RECT 15.130 108.515 15.460 108.685 ;
        RECT 16.090 108.515 16.420 108.685 ;
        RECT 17.050 108.515 17.380 108.685 ;
        RECT 19.855 108.515 20.185 108.685 ;
        RECT 20.815 108.515 21.145 108.685 ;
        RECT 21.775 108.515 22.105 108.685 ;
        RECT 22.735 108.515 23.065 108.685 ;
        RECT 23.695 108.515 24.025 108.685 ;
        RECT 24.655 108.515 24.985 108.685 ;
        RECT 27.100 105.800 27.430 106.040 ;
        RECT 18.375 105.585 18.705 105.755 ;
      LAYER mcon ;
        RECT 12.330 108.515 12.500 108.685 ;
        RECT 13.290 108.515 13.460 108.685 ;
        RECT 14.250 108.515 14.420 108.685 ;
        RECT 15.210 108.515 15.380 108.685 ;
        RECT 16.170 108.515 16.340 108.685 ;
        RECT 17.130 108.515 17.300 108.685 ;
        RECT 19.935 108.515 20.105 108.685 ;
        RECT 20.895 108.515 21.065 108.685 ;
        RECT 21.855 108.515 22.025 108.685 ;
        RECT 22.815 108.515 22.985 108.685 ;
        RECT 23.775 108.515 23.945 108.685 ;
        RECT 24.735 108.515 24.905 108.685 ;
        RECT 27.250 105.815 27.420 105.985 ;
        RECT 18.455 105.585 18.625 105.755 ;
      LAYER met1 ;
        RECT 12.235 108.475 12.595 108.735 ;
        RECT 13.200 108.475 13.560 108.735 ;
        RECT 14.155 108.475 14.515 108.735 ;
        RECT 15.115 108.475 15.475 108.735 ;
        RECT 16.075 108.475 16.435 108.735 ;
        RECT 17.035 108.475 17.395 108.735 ;
        RECT 19.840 108.475 20.200 108.735 ;
        RECT 20.805 108.475 21.165 108.735 ;
        RECT 21.760 108.475 22.120 108.735 ;
        RECT 22.720 108.475 23.080 108.735 ;
        RECT 23.680 108.475 24.040 108.735 ;
        RECT 24.640 108.475 25.000 108.735 ;
        RECT 18.355 105.590 18.715 105.850 ;
        RECT 27.190 105.755 27.560 106.025 ;
        RECT 18.395 105.555 18.685 105.590 ;
      LAYER via ;
        RECT 12.285 108.475 12.545 108.735 ;
        RECT 13.250 108.475 13.510 108.735 ;
        RECT 14.205 108.475 14.465 108.735 ;
        RECT 15.165 108.475 15.425 108.735 ;
        RECT 16.125 108.475 16.385 108.735 ;
        RECT 17.085 108.475 17.345 108.735 ;
        RECT 19.890 108.475 20.150 108.735 ;
        RECT 20.855 108.475 21.115 108.735 ;
        RECT 21.810 108.475 22.070 108.735 ;
        RECT 22.770 108.475 23.030 108.735 ;
        RECT 23.730 108.475 23.990 108.735 ;
        RECT 24.690 108.475 24.950 108.735 ;
        RECT 18.405 105.590 18.665 105.850 ;
        RECT 27.245 105.760 27.505 106.020 ;
      LAYER met2 ;
        RECT 12.285 108.735 12.545 108.785 ;
        RECT 13.250 108.735 13.510 108.785 ;
        RECT 14.205 108.735 14.465 108.785 ;
        RECT 15.165 108.735 15.425 108.785 ;
        RECT 16.125 108.735 16.385 108.785 ;
        RECT 17.085 108.735 17.345 108.785 ;
        RECT 19.890 108.735 20.150 108.785 ;
        RECT 20.855 108.735 21.115 108.785 ;
        RECT 21.810 108.735 22.070 108.785 ;
        RECT 22.770 108.735 23.030 108.785 ;
        RECT 23.730 108.735 23.990 108.785 ;
        RECT 24.690 108.735 24.950 108.785 ;
        RECT 11.165 108.475 29.230 108.735 ;
        RECT 12.285 108.425 12.545 108.475 ;
        RECT 13.250 108.425 13.510 108.475 ;
        RECT 14.205 108.425 14.465 108.475 ;
        RECT 15.165 108.425 15.425 108.475 ;
        RECT 16.125 108.425 16.385 108.475 ;
        RECT 17.085 108.425 17.345 108.475 ;
        RECT 18.405 105.540 18.665 108.475 ;
        RECT 19.890 108.425 20.150 108.475 ;
        RECT 20.855 108.425 21.115 108.475 ;
        RECT 21.810 108.425 22.070 108.475 ;
        RECT 22.770 108.425 23.030 108.475 ;
        RECT 23.730 108.425 23.990 108.475 ;
        RECT 24.690 108.425 24.950 108.475 ;
        RECT 27.240 106.055 27.510 106.075 ;
        RECT 28.040 106.055 28.300 108.475 ;
        RECT 27.240 105.795 28.300 106.055 ;
        RECT 27.240 105.705 27.510 105.795 ;
    END
  END en_b[15]
  PIN en_b[16]
    DIRECTION INOUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 4.402500 ;
    PORT
      LAYER li1 ;
        RECT 12.250 102.080 12.580 102.250 ;
        RECT 13.210 102.080 13.540 102.250 ;
        RECT 14.170 102.080 14.500 102.250 ;
        RECT 15.130 102.080 15.460 102.250 ;
        RECT 16.090 102.080 16.420 102.250 ;
        RECT 17.050 102.080 17.380 102.250 ;
        RECT 19.855 102.080 20.185 102.250 ;
        RECT 20.815 102.080 21.145 102.250 ;
        RECT 21.775 102.080 22.105 102.250 ;
        RECT 22.735 102.080 23.065 102.250 ;
        RECT 23.695 102.080 24.025 102.250 ;
        RECT 24.655 102.080 24.985 102.250 ;
        RECT 27.100 99.365 27.430 99.605 ;
        RECT 18.375 99.150 18.705 99.320 ;
      LAYER mcon ;
        RECT 12.330 102.080 12.500 102.250 ;
        RECT 13.290 102.080 13.460 102.250 ;
        RECT 14.250 102.080 14.420 102.250 ;
        RECT 15.210 102.080 15.380 102.250 ;
        RECT 16.170 102.080 16.340 102.250 ;
        RECT 17.130 102.080 17.300 102.250 ;
        RECT 19.935 102.080 20.105 102.250 ;
        RECT 20.895 102.080 21.065 102.250 ;
        RECT 21.855 102.080 22.025 102.250 ;
        RECT 22.815 102.080 22.985 102.250 ;
        RECT 23.775 102.080 23.945 102.250 ;
        RECT 24.735 102.080 24.905 102.250 ;
        RECT 27.250 99.380 27.420 99.550 ;
        RECT 18.455 99.150 18.625 99.320 ;
      LAYER met1 ;
        RECT 12.235 102.040 12.595 102.300 ;
        RECT 13.200 102.040 13.560 102.300 ;
        RECT 14.155 102.040 14.515 102.300 ;
        RECT 15.115 102.040 15.475 102.300 ;
        RECT 16.075 102.040 16.435 102.300 ;
        RECT 17.035 102.040 17.395 102.300 ;
        RECT 19.840 102.040 20.200 102.300 ;
        RECT 20.805 102.040 21.165 102.300 ;
        RECT 21.760 102.040 22.120 102.300 ;
        RECT 22.720 102.040 23.080 102.300 ;
        RECT 23.680 102.040 24.040 102.300 ;
        RECT 24.640 102.040 25.000 102.300 ;
        RECT 18.355 99.155 18.715 99.415 ;
        RECT 27.190 99.320 27.560 99.590 ;
        RECT 18.395 99.120 18.685 99.155 ;
      LAYER via ;
        RECT 12.285 102.040 12.545 102.300 ;
        RECT 13.250 102.040 13.510 102.300 ;
        RECT 14.205 102.040 14.465 102.300 ;
        RECT 15.165 102.040 15.425 102.300 ;
        RECT 16.125 102.040 16.385 102.300 ;
        RECT 17.085 102.040 17.345 102.300 ;
        RECT 19.890 102.040 20.150 102.300 ;
        RECT 20.855 102.040 21.115 102.300 ;
        RECT 21.810 102.040 22.070 102.300 ;
        RECT 22.770 102.040 23.030 102.300 ;
        RECT 23.730 102.040 23.990 102.300 ;
        RECT 24.690 102.040 24.950 102.300 ;
        RECT 18.405 99.155 18.665 99.415 ;
        RECT 27.245 99.325 27.505 99.585 ;
      LAYER met2 ;
        RECT 12.285 102.300 12.545 102.350 ;
        RECT 13.250 102.300 13.510 102.350 ;
        RECT 14.205 102.300 14.465 102.350 ;
        RECT 15.165 102.300 15.425 102.350 ;
        RECT 16.125 102.300 16.385 102.350 ;
        RECT 17.085 102.300 17.345 102.350 ;
        RECT 19.890 102.300 20.150 102.350 ;
        RECT 20.855 102.300 21.115 102.350 ;
        RECT 21.810 102.300 22.070 102.350 ;
        RECT 22.770 102.300 23.030 102.350 ;
        RECT 23.730 102.300 23.990 102.350 ;
        RECT 24.690 102.300 24.950 102.350 ;
        RECT 11.165 102.040 29.230 102.300 ;
        RECT 12.285 101.990 12.545 102.040 ;
        RECT 13.250 101.990 13.510 102.040 ;
        RECT 14.205 101.990 14.465 102.040 ;
        RECT 15.165 101.990 15.425 102.040 ;
        RECT 16.125 101.990 16.385 102.040 ;
        RECT 17.085 101.990 17.345 102.040 ;
        RECT 18.405 99.105 18.665 102.040 ;
        RECT 19.890 101.990 20.150 102.040 ;
        RECT 20.855 101.990 21.115 102.040 ;
        RECT 21.810 101.990 22.070 102.040 ;
        RECT 22.770 101.990 23.030 102.040 ;
        RECT 23.730 101.990 23.990 102.040 ;
        RECT 24.690 101.990 24.950 102.040 ;
        RECT 27.240 99.620 27.510 99.640 ;
        RECT 28.040 99.620 28.300 102.040 ;
        RECT 27.240 99.360 28.300 99.620 ;
        RECT 27.240 99.270 27.510 99.360 ;
    END
  END en_b[16]
  PIN en_b[17]
    DIRECTION INOUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 4.402500 ;
    PORT
      LAYER li1 ;
        RECT 12.250 95.645 12.580 95.815 ;
        RECT 13.210 95.645 13.540 95.815 ;
        RECT 14.170 95.645 14.500 95.815 ;
        RECT 15.130 95.645 15.460 95.815 ;
        RECT 16.090 95.645 16.420 95.815 ;
        RECT 17.050 95.645 17.380 95.815 ;
        RECT 19.855 95.645 20.185 95.815 ;
        RECT 20.815 95.645 21.145 95.815 ;
        RECT 21.775 95.645 22.105 95.815 ;
        RECT 22.735 95.645 23.065 95.815 ;
        RECT 23.695 95.645 24.025 95.815 ;
        RECT 24.655 95.645 24.985 95.815 ;
        RECT 27.100 92.930 27.430 93.170 ;
        RECT 18.375 92.715 18.705 92.885 ;
      LAYER mcon ;
        RECT 12.330 95.645 12.500 95.815 ;
        RECT 13.290 95.645 13.460 95.815 ;
        RECT 14.250 95.645 14.420 95.815 ;
        RECT 15.210 95.645 15.380 95.815 ;
        RECT 16.170 95.645 16.340 95.815 ;
        RECT 17.130 95.645 17.300 95.815 ;
        RECT 19.935 95.645 20.105 95.815 ;
        RECT 20.895 95.645 21.065 95.815 ;
        RECT 21.855 95.645 22.025 95.815 ;
        RECT 22.815 95.645 22.985 95.815 ;
        RECT 23.775 95.645 23.945 95.815 ;
        RECT 24.735 95.645 24.905 95.815 ;
        RECT 27.250 92.945 27.420 93.115 ;
        RECT 18.455 92.715 18.625 92.885 ;
      LAYER met1 ;
        RECT 12.235 95.605 12.595 95.865 ;
        RECT 13.200 95.605 13.560 95.865 ;
        RECT 14.155 95.605 14.515 95.865 ;
        RECT 15.115 95.605 15.475 95.865 ;
        RECT 16.075 95.605 16.435 95.865 ;
        RECT 17.035 95.605 17.395 95.865 ;
        RECT 19.840 95.605 20.200 95.865 ;
        RECT 20.805 95.605 21.165 95.865 ;
        RECT 21.760 95.605 22.120 95.865 ;
        RECT 22.720 95.605 23.080 95.865 ;
        RECT 23.680 95.605 24.040 95.865 ;
        RECT 24.640 95.605 25.000 95.865 ;
        RECT 18.355 92.720 18.715 92.980 ;
        RECT 27.190 92.885 27.560 93.155 ;
        RECT 18.395 92.685 18.685 92.720 ;
      LAYER via ;
        RECT 12.285 95.605 12.545 95.865 ;
        RECT 13.250 95.605 13.510 95.865 ;
        RECT 14.205 95.605 14.465 95.865 ;
        RECT 15.165 95.605 15.425 95.865 ;
        RECT 16.125 95.605 16.385 95.865 ;
        RECT 17.085 95.605 17.345 95.865 ;
        RECT 19.890 95.605 20.150 95.865 ;
        RECT 20.855 95.605 21.115 95.865 ;
        RECT 21.810 95.605 22.070 95.865 ;
        RECT 22.770 95.605 23.030 95.865 ;
        RECT 23.730 95.605 23.990 95.865 ;
        RECT 24.690 95.605 24.950 95.865 ;
        RECT 18.405 92.720 18.665 92.980 ;
        RECT 27.245 92.890 27.505 93.150 ;
      LAYER met2 ;
        RECT 12.285 95.865 12.545 95.915 ;
        RECT 13.250 95.865 13.510 95.915 ;
        RECT 14.205 95.865 14.465 95.915 ;
        RECT 15.165 95.865 15.425 95.915 ;
        RECT 16.125 95.865 16.385 95.915 ;
        RECT 17.085 95.865 17.345 95.915 ;
        RECT 19.890 95.865 20.150 95.915 ;
        RECT 20.855 95.865 21.115 95.915 ;
        RECT 21.810 95.865 22.070 95.915 ;
        RECT 22.770 95.865 23.030 95.915 ;
        RECT 23.730 95.865 23.990 95.915 ;
        RECT 24.690 95.865 24.950 95.915 ;
        RECT 11.165 95.605 29.230 95.865 ;
        RECT 12.285 95.555 12.545 95.605 ;
        RECT 13.250 95.555 13.510 95.605 ;
        RECT 14.205 95.555 14.465 95.605 ;
        RECT 15.165 95.555 15.425 95.605 ;
        RECT 16.125 95.555 16.385 95.605 ;
        RECT 17.085 95.555 17.345 95.605 ;
        RECT 18.405 92.670 18.665 95.605 ;
        RECT 19.890 95.555 20.150 95.605 ;
        RECT 20.855 95.555 21.115 95.605 ;
        RECT 21.810 95.555 22.070 95.605 ;
        RECT 22.770 95.555 23.030 95.605 ;
        RECT 23.730 95.555 23.990 95.605 ;
        RECT 24.690 95.555 24.950 95.605 ;
        RECT 27.240 93.185 27.510 93.205 ;
        RECT 28.040 93.185 28.300 95.605 ;
        RECT 27.240 92.925 28.300 93.185 ;
        RECT 27.240 92.835 27.510 92.925 ;
    END
  END en_b[17]
  PIN en_b[18]
    DIRECTION INOUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 4.402500 ;
    PORT
      LAYER li1 ;
        RECT 12.250 89.210 12.580 89.380 ;
        RECT 13.210 89.210 13.540 89.380 ;
        RECT 14.170 89.210 14.500 89.380 ;
        RECT 15.130 89.210 15.460 89.380 ;
        RECT 16.090 89.210 16.420 89.380 ;
        RECT 17.050 89.210 17.380 89.380 ;
        RECT 19.855 89.210 20.185 89.380 ;
        RECT 20.815 89.210 21.145 89.380 ;
        RECT 21.775 89.210 22.105 89.380 ;
        RECT 22.735 89.210 23.065 89.380 ;
        RECT 23.695 89.210 24.025 89.380 ;
        RECT 24.655 89.210 24.985 89.380 ;
        RECT 27.100 86.495 27.430 86.735 ;
        RECT 18.375 86.280 18.705 86.450 ;
      LAYER mcon ;
        RECT 12.330 89.210 12.500 89.380 ;
        RECT 13.290 89.210 13.460 89.380 ;
        RECT 14.250 89.210 14.420 89.380 ;
        RECT 15.210 89.210 15.380 89.380 ;
        RECT 16.170 89.210 16.340 89.380 ;
        RECT 17.130 89.210 17.300 89.380 ;
        RECT 19.935 89.210 20.105 89.380 ;
        RECT 20.895 89.210 21.065 89.380 ;
        RECT 21.855 89.210 22.025 89.380 ;
        RECT 22.815 89.210 22.985 89.380 ;
        RECT 23.775 89.210 23.945 89.380 ;
        RECT 24.735 89.210 24.905 89.380 ;
        RECT 27.250 86.510 27.420 86.680 ;
        RECT 18.455 86.280 18.625 86.450 ;
      LAYER met1 ;
        RECT 12.235 89.170 12.595 89.430 ;
        RECT 13.200 89.170 13.560 89.430 ;
        RECT 14.155 89.170 14.515 89.430 ;
        RECT 15.115 89.170 15.475 89.430 ;
        RECT 16.075 89.170 16.435 89.430 ;
        RECT 17.035 89.170 17.395 89.430 ;
        RECT 19.840 89.170 20.200 89.430 ;
        RECT 20.805 89.170 21.165 89.430 ;
        RECT 21.760 89.170 22.120 89.430 ;
        RECT 22.720 89.170 23.080 89.430 ;
        RECT 23.680 89.170 24.040 89.430 ;
        RECT 24.640 89.170 25.000 89.430 ;
        RECT 18.355 86.285 18.715 86.545 ;
        RECT 27.190 86.450 27.560 86.720 ;
        RECT 18.395 86.250 18.685 86.285 ;
      LAYER via ;
        RECT 12.285 89.170 12.545 89.430 ;
        RECT 13.250 89.170 13.510 89.430 ;
        RECT 14.205 89.170 14.465 89.430 ;
        RECT 15.165 89.170 15.425 89.430 ;
        RECT 16.125 89.170 16.385 89.430 ;
        RECT 17.085 89.170 17.345 89.430 ;
        RECT 19.890 89.170 20.150 89.430 ;
        RECT 20.855 89.170 21.115 89.430 ;
        RECT 21.810 89.170 22.070 89.430 ;
        RECT 22.770 89.170 23.030 89.430 ;
        RECT 23.730 89.170 23.990 89.430 ;
        RECT 24.690 89.170 24.950 89.430 ;
        RECT 18.405 86.285 18.665 86.545 ;
        RECT 27.245 86.455 27.505 86.715 ;
      LAYER met2 ;
        RECT 12.285 89.430 12.545 89.480 ;
        RECT 13.250 89.430 13.510 89.480 ;
        RECT 14.205 89.430 14.465 89.480 ;
        RECT 15.165 89.430 15.425 89.480 ;
        RECT 16.125 89.430 16.385 89.480 ;
        RECT 17.085 89.430 17.345 89.480 ;
        RECT 19.890 89.430 20.150 89.480 ;
        RECT 20.855 89.430 21.115 89.480 ;
        RECT 21.810 89.430 22.070 89.480 ;
        RECT 22.770 89.430 23.030 89.480 ;
        RECT 23.730 89.430 23.990 89.480 ;
        RECT 24.690 89.430 24.950 89.480 ;
        RECT 11.165 89.170 29.230 89.430 ;
        RECT 12.285 89.120 12.545 89.170 ;
        RECT 13.250 89.120 13.510 89.170 ;
        RECT 14.205 89.120 14.465 89.170 ;
        RECT 15.165 89.120 15.425 89.170 ;
        RECT 16.125 89.120 16.385 89.170 ;
        RECT 17.085 89.120 17.345 89.170 ;
        RECT 18.405 86.235 18.665 89.170 ;
        RECT 19.890 89.120 20.150 89.170 ;
        RECT 20.855 89.120 21.115 89.170 ;
        RECT 21.810 89.120 22.070 89.170 ;
        RECT 22.770 89.120 23.030 89.170 ;
        RECT 23.730 89.120 23.990 89.170 ;
        RECT 24.690 89.120 24.950 89.170 ;
        RECT 27.240 86.750 27.510 86.770 ;
        RECT 28.040 86.750 28.300 89.170 ;
        RECT 27.240 86.490 28.300 86.750 ;
        RECT 27.240 86.400 27.510 86.490 ;
    END
  END en_b[18]
  PIN en_b[19]
    DIRECTION INOUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 4.402500 ;
    PORT
      LAYER li1 ;
        RECT 12.250 82.775 12.580 82.945 ;
        RECT 13.210 82.775 13.540 82.945 ;
        RECT 14.170 82.775 14.500 82.945 ;
        RECT 15.130 82.775 15.460 82.945 ;
        RECT 16.090 82.775 16.420 82.945 ;
        RECT 17.050 82.775 17.380 82.945 ;
        RECT 19.855 82.775 20.185 82.945 ;
        RECT 20.815 82.775 21.145 82.945 ;
        RECT 21.775 82.775 22.105 82.945 ;
        RECT 22.735 82.775 23.065 82.945 ;
        RECT 23.695 82.775 24.025 82.945 ;
        RECT 24.655 82.775 24.985 82.945 ;
        RECT 27.100 80.060 27.430 80.300 ;
        RECT 18.375 79.845 18.705 80.015 ;
      LAYER mcon ;
        RECT 12.330 82.775 12.500 82.945 ;
        RECT 13.290 82.775 13.460 82.945 ;
        RECT 14.250 82.775 14.420 82.945 ;
        RECT 15.210 82.775 15.380 82.945 ;
        RECT 16.170 82.775 16.340 82.945 ;
        RECT 17.130 82.775 17.300 82.945 ;
        RECT 19.935 82.775 20.105 82.945 ;
        RECT 20.895 82.775 21.065 82.945 ;
        RECT 21.855 82.775 22.025 82.945 ;
        RECT 22.815 82.775 22.985 82.945 ;
        RECT 23.775 82.775 23.945 82.945 ;
        RECT 24.735 82.775 24.905 82.945 ;
        RECT 27.250 80.075 27.420 80.245 ;
        RECT 18.455 79.845 18.625 80.015 ;
      LAYER met1 ;
        RECT 12.235 82.735 12.595 82.995 ;
        RECT 13.200 82.735 13.560 82.995 ;
        RECT 14.155 82.735 14.515 82.995 ;
        RECT 15.115 82.735 15.475 82.995 ;
        RECT 16.075 82.735 16.435 82.995 ;
        RECT 17.035 82.735 17.395 82.995 ;
        RECT 19.840 82.735 20.200 82.995 ;
        RECT 20.805 82.735 21.165 82.995 ;
        RECT 21.760 82.735 22.120 82.995 ;
        RECT 22.720 82.735 23.080 82.995 ;
        RECT 23.680 82.735 24.040 82.995 ;
        RECT 24.640 82.735 25.000 82.995 ;
        RECT 18.355 79.850 18.715 80.110 ;
        RECT 27.190 80.015 27.560 80.285 ;
        RECT 18.395 79.815 18.685 79.850 ;
      LAYER via ;
        RECT 12.285 82.735 12.545 82.995 ;
        RECT 13.250 82.735 13.510 82.995 ;
        RECT 14.205 82.735 14.465 82.995 ;
        RECT 15.165 82.735 15.425 82.995 ;
        RECT 16.125 82.735 16.385 82.995 ;
        RECT 17.085 82.735 17.345 82.995 ;
        RECT 19.890 82.735 20.150 82.995 ;
        RECT 20.855 82.735 21.115 82.995 ;
        RECT 21.810 82.735 22.070 82.995 ;
        RECT 22.770 82.735 23.030 82.995 ;
        RECT 23.730 82.735 23.990 82.995 ;
        RECT 24.690 82.735 24.950 82.995 ;
        RECT 18.405 79.850 18.665 80.110 ;
        RECT 27.245 80.020 27.505 80.280 ;
      LAYER met2 ;
        RECT 12.285 82.995 12.545 83.045 ;
        RECT 13.250 82.995 13.510 83.045 ;
        RECT 14.205 82.995 14.465 83.045 ;
        RECT 15.165 82.995 15.425 83.045 ;
        RECT 16.125 82.995 16.385 83.045 ;
        RECT 17.085 82.995 17.345 83.045 ;
        RECT 19.890 82.995 20.150 83.045 ;
        RECT 20.855 82.995 21.115 83.045 ;
        RECT 21.810 82.995 22.070 83.045 ;
        RECT 22.770 82.995 23.030 83.045 ;
        RECT 23.730 82.995 23.990 83.045 ;
        RECT 24.690 82.995 24.950 83.045 ;
        RECT 11.165 82.735 29.230 82.995 ;
        RECT 12.285 82.685 12.545 82.735 ;
        RECT 13.250 82.685 13.510 82.735 ;
        RECT 14.205 82.685 14.465 82.735 ;
        RECT 15.165 82.685 15.425 82.735 ;
        RECT 16.125 82.685 16.385 82.735 ;
        RECT 17.085 82.685 17.345 82.735 ;
        RECT 18.405 79.800 18.665 82.735 ;
        RECT 19.890 82.685 20.150 82.735 ;
        RECT 20.855 82.685 21.115 82.735 ;
        RECT 21.810 82.685 22.070 82.735 ;
        RECT 22.770 82.685 23.030 82.735 ;
        RECT 23.730 82.685 23.990 82.735 ;
        RECT 24.690 82.685 24.950 82.735 ;
        RECT 27.240 80.315 27.510 80.335 ;
        RECT 28.040 80.315 28.300 82.735 ;
        RECT 27.240 80.055 28.300 80.315 ;
        RECT 27.240 79.965 27.510 80.055 ;
    END
  END en_b[19]
  PIN en_b[20]
    DIRECTION INOUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 4.402500 ;
    PORT
      LAYER li1 ;
        RECT 12.250 76.340 12.580 76.510 ;
        RECT 13.210 76.340 13.540 76.510 ;
        RECT 14.170 76.340 14.500 76.510 ;
        RECT 15.130 76.340 15.460 76.510 ;
        RECT 16.090 76.340 16.420 76.510 ;
        RECT 17.050 76.340 17.380 76.510 ;
        RECT 19.855 76.340 20.185 76.510 ;
        RECT 20.815 76.340 21.145 76.510 ;
        RECT 21.775 76.340 22.105 76.510 ;
        RECT 22.735 76.340 23.065 76.510 ;
        RECT 23.695 76.340 24.025 76.510 ;
        RECT 24.655 76.340 24.985 76.510 ;
        RECT 27.100 73.625 27.430 73.865 ;
        RECT 18.375 73.410 18.705 73.580 ;
      LAYER mcon ;
        RECT 12.330 76.340 12.500 76.510 ;
        RECT 13.290 76.340 13.460 76.510 ;
        RECT 14.250 76.340 14.420 76.510 ;
        RECT 15.210 76.340 15.380 76.510 ;
        RECT 16.170 76.340 16.340 76.510 ;
        RECT 17.130 76.340 17.300 76.510 ;
        RECT 19.935 76.340 20.105 76.510 ;
        RECT 20.895 76.340 21.065 76.510 ;
        RECT 21.855 76.340 22.025 76.510 ;
        RECT 22.815 76.340 22.985 76.510 ;
        RECT 23.775 76.340 23.945 76.510 ;
        RECT 24.735 76.340 24.905 76.510 ;
        RECT 27.250 73.640 27.420 73.810 ;
        RECT 18.455 73.410 18.625 73.580 ;
      LAYER met1 ;
        RECT 12.235 76.300 12.595 76.560 ;
        RECT 13.200 76.300 13.560 76.560 ;
        RECT 14.155 76.300 14.515 76.560 ;
        RECT 15.115 76.300 15.475 76.560 ;
        RECT 16.075 76.300 16.435 76.560 ;
        RECT 17.035 76.300 17.395 76.560 ;
        RECT 19.840 76.300 20.200 76.560 ;
        RECT 20.805 76.300 21.165 76.560 ;
        RECT 21.760 76.300 22.120 76.560 ;
        RECT 22.720 76.300 23.080 76.560 ;
        RECT 23.680 76.300 24.040 76.560 ;
        RECT 24.640 76.300 25.000 76.560 ;
        RECT 18.355 73.415 18.715 73.675 ;
        RECT 27.190 73.580 27.560 73.850 ;
        RECT 18.395 73.380 18.685 73.415 ;
      LAYER via ;
        RECT 12.285 76.300 12.545 76.560 ;
        RECT 13.250 76.300 13.510 76.560 ;
        RECT 14.205 76.300 14.465 76.560 ;
        RECT 15.165 76.300 15.425 76.560 ;
        RECT 16.125 76.300 16.385 76.560 ;
        RECT 17.085 76.300 17.345 76.560 ;
        RECT 19.890 76.300 20.150 76.560 ;
        RECT 20.855 76.300 21.115 76.560 ;
        RECT 21.810 76.300 22.070 76.560 ;
        RECT 22.770 76.300 23.030 76.560 ;
        RECT 23.730 76.300 23.990 76.560 ;
        RECT 24.690 76.300 24.950 76.560 ;
        RECT 18.405 73.415 18.665 73.675 ;
        RECT 27.245 73.585 27.505 73.845 ;
      LAYER met2 ;
        RECT 12.285 76.560 12.545 76.610 ;
        RECT 13.250 76.560 13.510 76.610 ;
        RECT 14.205 76.560 14.465 76.610 ;
        RECT 15.165 76.560 15.425 76.610 ;
        RECT 16.125 76.560 16.385 76.610 ;
        RECT 17.085 76.560 17.345 76.610 ;
        RECT 19.890 76.560 20.150 76.610 ;
        RECT 20.855 76.560 21.115 76.610 ;
        RECT 21.810 76.560 22.070 76.610 ;
        RECT 22.770 76.560 23.030 76.610 ;
        RECT 23.730 76.560 23.990 76.610 ;
        RECT 24.690 76.560 24.950 76.610 ;
        RECT 11.165 76.300 29.230 76.560 ;
        RECT 12.285 76.250 12.545 76.300 ;
        RECT 13.250 76.250 13.510 76.300 ;
        RECT 14.205 76.250 14.465 76.300 ;
        RECT 15.165 76.250 15.425 76.300 ;
        RECT 16.125 76.250 16.385 76.300 ;
        RECT 17.085 76.250 17.345 76.300 ;
        RECT 18.405 73.365 18.665 76.300 ;
        RECT 19.890 76.250 20.150 76.300 ;
        RECT 20.855 76.250 21.115 76.300 ;
        RECT 21.810 76.250 22.070 76.300 ;
        RECT 22.770 76.250 23.030 76.300 ;
        RECT 23.730 76.250 23.990 76.300 ;
        RECT 24.690 76.250 24.950 76.300 ;
        RECT 27.240 73.880 27.510 73.900 ;
        RECT 28.040 73.880 28.300 76.300 ;
        RECT 27.240 73.620 28.300 73.880 ;
        RECT 27.240 73.530 27.510 73.620 ;
    END
  END en_b[20]
  PIN en_b[21]
    DIRECTION INOUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 4.402500 ;
    PORT
      LAYER li1 ;
        RECT 12.250 69.905 12.580 70.075 ;
        RECT 13.210 69.905 13.540 70.075 ;
        RECT 14.170 69.905 14.500 70.075 ;
        RECT 15.130 69.905 15.460 70.075 ;
        RECT 16.090 69.905 16.420 70.075 ;
        RECT 17.050 69.905 17.380 70.075 ;
        RECT 19.855 69.905 20.185 70.075 ;
        RECT 20.815 69.905 21.145 70.075 ;
        RECT 21.775 69.905 22.105 70.075 ;
        RECT 22.735 69.905 23.065 70.075 ;
        RECT 23.695 69.905 24.025 70.075 ;
        RECT 24.655 69.905 24.985 70.075 ;
        RECT 27.100 67.190 27.430 67.430 ;
        RECT 18.375 66.975 18.705 67.145 ;
      LAYER mcon ;
        RECT 12.330 69.905 12.500 70.075 ;
        RECT 13.290 69.905 13.460 70.075 ;
        RECT 14.250 69.905 14.420 70.075 ;
        RECT 15.210 69.905 15.380 70.075 ;
        RECT 16.170 69.905 16.340 70.075 ;
        RECT 17.130 69.905 17.300 70.075 ;
        RECT 19.935 69.905 20.105 70.075 ;
        RECT 20.895 69.905 21.065 70.075 ;
        RECT 21.855 69.905 22.025 70.075 ;
        RECT 22.815 69.905 22.985 70.075 ;
        RECT 23.775 69.905 23.945 70.075 ;
        RECT 24.735 69.905 24.905 70.075 ;
        RECT 27.250 67.205 27.420 67.375 ;
        RECT 18.455 66.975 18.625 67.145 ;
      LAYER met1 ;
        RECT 12.235 69.865 12.595 70.125 ;
        RECT 13.200 69.865 13.560 70.125 ;
        RECT 14.155 69.865 14.515 70.125 ;
        RECT 15.115 69.865 15.475 70.125 ;
        RECT 16.075 69.865 16.435 70.125 ;
        RECT 17.035 69.865 17.395 70.125 ;
        RECT 19.840 69.865 20.200 70.125 ;
        RECT 20.805 69.865 21.165 70.125 ;
        RECT 21.760 69.865 22.120 70.125 ;
        RECT 22.720 69.865 23.080 70.125 ;
        RECT 23.680 69.865 24.040 70.125 ;
        RECT 24.640 69.865 25.000 70.125 ;
        RECT 18.355 66.980 18.715 67.240 ;
        RECT 27.190 67.145 27.560 67.415 ;
        RECT 18.395 66.945 18.685 66.980 ;
      LAYER via ;
        RECT 12.285 69.865 12.545 70.125 ;
        RECT 13.250 69.865 13.510 70.125 ;
        RECT 14.205 69.865 14.465 70.125 ;
        RECT 15.165 69.865 15.425 70.125 ;
        RECT 16.125 69.865 16.385 70.125 ;
        RECT 17.085 69.865 17.345 70.125 ;
        RECT 19.890 69.865 20.150 70.125 ;
        RECT 20.855 69.865 21.115 70.125 ;
        RECT 21.810 69.865 22.070 70.125 ;
        RECT 22.770 69.865 23.030 70.125 ;
        RECT 23.730 69.865 23.990 70.125 ;
        RECT 24.690 69.865 24.950 70.125 ;
        RECT 18.405 66.980 18.665 67.240 ;
        RECT 27.245 67.150 27.505 67.410 ;
      LAYER met2 ;
        RECT 12.285 70.125 12.545 70.175 ;
        RECT 13.250 70.125 13.510 70.175 ;
        RECT 14.205 70.125 14.465 70.175 ;
        RECT 15.165 70.125 15.425 70.175 ;
        RECT 16.125 70.125 16.385 70.175 ;
        RECT 17.085 70.125 17.345 70.175 ;
        RECT 19.890 70.125 20.150 70.175 ;
        RECT 20.855 70.125 21.115 70.175 ;
        RECT 21.810 70.125 22.070 70.175 ;
        RECT 22.770 70.125 23.030 70.175 ;
        RECT 23.730 70.125 23.990 70.175 ;
        RECT 24.690 70.125 24.950 70.175 ;
        RECT 11.165 69.865 29.230 70.125 ;
        RECT 12.285 69.815 12.545 69.865 ;
        RECT 13.250 69.815 13.510 69.865 ;
        RECT 14.205 69.815 14.465 69.865 ;
        RECT 15.165 69.815 15.425 69.865 ;
        RECT 16.125 69.815 16.385 69.865 ;
        RECT 17.085 69.815 17.345 69.865 ;
        RECT 18.405 66.930 18.665 69.865 ;
        RECT 19.890 69.815 20.150 69.865 ;
        RECT 20.855 69.815 21.115 69.865 ;
        RECT 21.810 69.815 22.070 69.865 ;
        RECT 22.770 69.815 23.030 69.865 ;
        RECT 23.730 69.815 23.990 69.865 ;
        RECT 24.690 69.815 24.950 69.865 ;
        RECT 27.240 67.445 27.510 67.465 ;
        RECT 28.040 67.445 28.300 69.865 ;
        RECT 27.240 67.185 28.300 67.445 ;
        RECT 27.240 67.095 27.510 67.185 ;
    END
  END en_b[21]
  PIN en_b[22]
    DIRECTION INOUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 4.402500 ;
    PORT
      LAYER li1 ;
        RECT 12.250 63.470 12.580 63.640 ;
        RECT 13.210 63.470 13.540 63.640 ;
        RECT 14.170 63.470 14.500 63.640 ;
        RECT 15.130 63.470 15.460 63.640 ;
        RECT 16.090 63.470 16.420 63.640 ;
        RECT 17.050 63.470 17.380 63.640 ;
        RECT 19.855 63.470 20.185 63.640 ;
        RECT 20.815 63.470 21.145 63.640 ;
        RECT 21.775 63.470 22.105 63.640 ;
        RECT 22.735 63.470 23.065 63.640 ;
        RECT 23.695 63.470 24.025 63.640 ;
        RECT 24.655 63.470 24.985 63.640 ;
        RECT 27.100 60.755 27.430 60.995 ;
        RECT 18.375 60.540 18.705 60.710 ;
      LAYER mcon ;
        RECT 12.330 63.470 12.500 63.640 ;
        RECT 13.290 63.470 13.460 63.640 ;
        RECT 14.250 63.470 14.420 63.640 ;
        RECT 15.210 63.470 15.380 63.640 ;
        RECT 16.170 63.470 16.340 63.640 ;
        RECT 17.130 63.470 17.300 63.640 ;
        RECT 19.935 63.470 20.105 63.640 ;
        RECT 20.895 63.470 21.065 63.640 ;
        RECT 21.855 63.470 22.025 63.640 ;
        RECT 22.815 63.470 22.985 63.640 ;
        RECT 23.775 63.470 23.945 63.640 ;
        RECT 24.735 63.470 24.905 63.640 ;
        RECT 27.250 60.770 27.420 60.940 ;
        RECT 18.455 60.540 18.625 60.710 ;
      LAYER met1 ;
        RECT 12.235 63.430 12.595 63.690 ;
        RECT 13.200 63.430 13.560 63.690 ;
        RECT 14.155 63.430 14.515 63.690 ;
        RECT 15.115 63.430 15.475 63.690 ;
        RECT 16.075 63.430 16.435 63.690 ;
        RECT 17.035 63.430 17.395 63.690 ;
        RECT 19.840 63.430 20.200 63.690 ;
        RECT 20.805 63.430 21.165 63.690 ;
        RECT 21.760 63.430 22.120 63.690 ;
        RECT 22.720 63.430 23.080 63.690 ;
        RECT 23.680 63.430 24.040 63.690 ;
        RECT 24.640 63.430 25.000 63.690 ;
        RECT 18.355 60.545 18.715 60.805 ;
        RECT 27.190 60.710 27.560 60.980 ;
        RECT 18.395 60.510 18.685 60.545 ;
      LAYER via ;
        RECT 12.285 63.430 12.545 63.690 ;
        RECT 13.250 63.430 13.510 63.690 ;
        RECT 14.205 63.430 14.465 63.690 ;
        RECT 15.165 63.430 15.425 63.690 ;
        RECT 16.125 63.430 16.385 63.690 ;
        RECT 17.085 63.430 17.345 63.690 ;
        RECT 19.890 63.430 20.150 63.690 ;
        RECT 20.855 63.430 21.115 63.690 ;
        RECT 21.810 63.430 22.070 63.690 ;
        RECT 22.770 63.430 23.030 63.690 ;
        RECT 23.730 63.430 23.990 63.690 ;
        RECT 24.690 63.430 24.950 63.690 ;
        RECT 18.405 60.545 18.665 60.805 ;
        RECT 27.245 60.715 27.505 60.975 ;
      LAYER met2 ;
        RECT 12.285 63.690 12.545 63.740 ;
        RECT 13.250 63.690 13.510 63.740 ;
        RECT 14.205 63.690 14.465 63.740 ;
        RECT 15.165 63.690 15.425 63.740 ;
        RECT 16.125 63.690 16.385 63.740 ;
        RECT 17.085 63.690 17.345 63.740 ;
        RECT 19.890 63.690 20.150 63.740 ;
        RECT 20.855 63.690 21.115 63.740 ;
        RECT 21.810 63.690 22.070 63.740 ;
        RECT 22.770 63.690 23.030 63.740 ;
        RECT 23.730 63.690 23.990 63.740 ;
        RECT 24.690 63.690 24.950 63.740 ;
        RECT 11.165 63.430 29.230 63.690 ;
        RECT 12.285 63.380 12.545 63.430 ;
        RECT 13.250 63.380 13.510 63.430 ;
        RECT 14.205 63.380 14.465 63.430 ;
        RECT 15.165 63.380 15.425 63.430 ;
        RECT 16.125 63.380 16.385 63.430 ;
        RECT 17.085 63.380 17.345 63.430 ;
        RECT 18.405 60.495 18.665 63.430 ;
        RECT 19.890 63.380 20.150 63.430 ;
        RECT 20.855 63.380 21.115 63.430 ;
        RECT 21.810 63.380 22.070 63.430 ;
        RECT 22.770 63.380 23.030 63.430 ;
        RECT 23.730 63.380 23.990 63.430 ;
        RECT 24.690 63.380 24.950 63.430 ;
        RECT 27.240 61.010 27.510 61.030 ;
        RECT 28.040 61.010 28.300 63.430 ;
        RECT 27.240 60.750 28.300 61.010 ;
        RECT 27.240 60.660 27.510 60.750 ;
    END
  END en_b[22]
  PIN en_b[23]
    DIRECTION INOUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 4.402500 ;
    PORT
      LAYER li1 ;
        RECT 12.250 57.035 12.580 57.205 ;
        RECT 13.210 57.035 13.540 57.205 ;
        RECT 14.170 57.035 14.500 57.205 ;
        RECT 15.130 57.035 15.460 57.205 ;
        RECT 16.090 57.035 16.420 57.205 ;
        RECT 17.050 57.035 17.380 57.205 ;
        RECT 19.855 57.035 20.185 57.205 ;
        RECT 20.815 57.035 21.145 57.205 ;
        RECT 21.775 57.035 22.105 57.205 ;
        RECT 22.735 57.035 23.065 57.205 ;
        RECT 23.695 57.035 24.025 57.205 ;
        RECT 24.655 57.035 24.985 57.205 ;
        RECT 27.100 54.320 27.430 54.560 ;
        RECT 18.375 54.105 18.705 54.275 ;
      LAYER mcon ;
        RECT 12.330 57.035 12.500 57.205 ;
        RECT 13.290 57.035 13.460 57.205 ;
        RECT 14.250 57.035 14.420 57.205 ;
        RECT 15.210 57.035 15.380 57.205 ;
        RECT 16.170 57.035 16.340 57.205 ;
        RECT 17.130 57.035 17.300 57.205 ;
        RECT 19.935 57.035 20.105 57.205 ;
        RECT 20.895 57.035 21.065 57.205 ;
        RECT 21.855 57.035 22.025 57.205 ;
        RECT 22.815 57.035 22.985 57.205 ;
        RECT 23.775 57.035 23.945 57.205 ;
        RECT 24.735 57.035 24.905 57.205 ;
        RECT 27.250 54.335 27.420 54.505 ;
        RECT 18.455 54.105 18.625 54.275 ;
      LAYER met1 ;
        RECT 12.235 56.995 12.595 57.255 ;
        RECT 13.200 56.995 13.560 57.255 ;
        RECT 14.155 56.995 14.515 57.255 ;
        RECT 15.115 56.995 15.475 57.255 ;
        RECT 16.075 56.995 16.435 57.255 ;
        RECT 17.035 56.995 17.395 57.255 ;
        RECT 19.840 56.995 20.200 57.255 ;
        RECT 20.805 56.995 21.165 57.255 ;
        RECT 21.760 56.995 22.120 57.255 ;
        RECT 22.720 56.995 23.080 57.255 ;
        RECT 23.680 56.995 24.040 57.255 ;
        RECT 24.640 56.995 25.000 57.255 ;
        RECT 18.355 54.110 18.715 54.370 ;
        RECT 27.190 54.275 27.560 54.545 ;
        RECT 18.395 54.075 18.685 54.110 ;
      LAYER via ;
        RECT 12.285 56.995 12.545 57.255 ;
        RECT 13.250 56.995 13.510 57.255 ;
        RECT 14.205 56.995 14.465 57.255 ;
        RECT 15.165 56.995 15.425 57.255 ;
        RECT 16.125 56.995 16.385 57.255 ;
        RECT 17.085 56.995 17.345 57.255 ;
        RECT 19.890 56.995 20.150 57.255 ;
        RECT 20.855 56.995 21.115 57.255 ;
        RECT 21.810 56.995 22.070 57.255 ;
        RECT 22.770 56.995 23.030 57.255 ;
        RECT 23.730 56.995 23.990 57.255 ;
        RECT 24.690 56.995 24.950 57.255 ;
        RECT 18.405 54.110 18.665 54.370 ;
        RECT 27.245 54.280 27.505 54.540 ;
      LAYER met2 ;
        RECT 12.285 57.255 12.545 57.305 ;
        RECT 13.250 57.255 13.510 57.305 ;
        RECT 14.205 57.255 14.465 57.305 ;
        RECT 15.165 57.255 15.425 57.305 ;
        RECT 16.125 57.255 16.385 57.305 ;
        RECT 17.085 57.255 17.345 57.305 ;
        RECT 19.890 57.255 20.150 57.305 ;
        RECT 20.855 57.255 21.115 57.305 ;
        RECT 21.810 57.255 22.070 57.305 ;
        RECT 22.770 57.255 23.030 57.305 ;
        RECT 23.730 57.255 23.990 57.305 ;
        RECT 24.690 57.255 24.950 57.305 ;
        RECT 11.165 56.995 29.230 57.255 ;
        RECT 12.285 56.945 12.545 56.995 ;
        RECT 13.250 56.945 13.510 56.995 ;
        RECT 14.205 56.945 14.465 56.995 ;
        RECT 15.165 56.945 15.425 56.995 ;
        RECT 16.125 56.945 16.385 56.995 ;
        RECT 17.085 56.945 17.345 56.995 ;
        RECT 18.405 54.060 18.665 56.995 ;
        RECT 19.890 56.945 20.150 56.995 ;
        RECT 20.855 56.945 21.115 56.995 ;
        RECT 21.810 56.945 22.070 56.995 ;
        RECT 22.770 56.945 23.030 56.995 ;
        RECT 23.730 56.945 23.990 56.995 ;
        RECT 24.690 56.945 24.950 56.995 ;
        RECT 27.240 54.575 27.510 54.595 ;
        RECT 28.040 54.575 28.300 56.995 ;
        RECT 27.240 54.315 28.300 54.575 ;
        RECT 27.240 54.225 27.510 54.315 ;
    END
  END en_b[23]
  PIN en_b[24]
    DIRECTION INOUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 4.402500 ;
    PORT
      LAYER li1 ;
        RECT 12.250 50.600 12.580 50.770 ;
        RECT 13.210 50.600 13.540 50.770 ;
        RECT 14.170 50.600 14.500 50.770 ;
        RECT 15.130 50.600 15.460 50.770 ;
        RECT 16.090 50.600 16.420 50.770 ;
        RECT 17.050 50.600 17.380 50.770 ;
        RECT 19.855 50.600 20.185 50.770 ;
        RECT 20.815 50.600 21.145 50.770 ;
        RECT 21.775 50.600 22.105 50.770 ;
        RECT 22.735 50.600 23.065 50.770 ;
        RECT 23.695 50.600 24.025 50.770 ;
        RECT 24.655 50.600 24.985 50.770 ;
        RECT 27.100 47.885 27.430 48.125 ;
        RECT 18.375 47.670 18.705 47.840 ;
      LAYER mcon ;
        RECT 12.330 50.600 12.500 50.770 ;
        RECT 13.290 50.600 13.460 50.770 ;
        RECT 14.250 50.600 14.420 50.770 ;
        RECT 15.210 50.600 15.380 50.770 ;
        RECT 16.170 50.600 16.340 50.770 ;
        RECT 17.130 50.600 17.300 50.770 ;
        RECT 19.935 50.600 20.105 50.770 ;
        RECT 20.895 50.600 21.065 50.770 ;
        RECT 21.855 50.600 22.025 50.770 ;
        RECT 22.815 50.600 22.985 50.770 ;
        RECT 23.775 50.600 23.945 50.770 ;
        RECT 24.735 50.600 24.905 50.770 ;
        RECT 27.250 47.900 27.420 48.070 ;
        RECT 18.455 47.670 18.625 47.840 ;
      LAYER met1 ;
        RECT 12.235 50.560 12.595 50.820 ;
        RECT 13.200 50.560 13.560 50.820 ;
        RECT 14.155 50.560 14.515 50.820 ;
        RECT 15.115 50.560 15.475 50.820 ;
        RECT 16.075 50.560 16.435 50.820 ;
        RECT 17.035 50.560 17.395 50.820 ;
        RECT 19.840 50.560 20.200 50.820 ;
        RECT 20.805 50.560 21.165 50.820 ;
        RECT 21.760 50.560 22.120 50.820 ;
        RECT 22.720 50.560 23.080 50.820 ;
        RECT 23.680 50.560 24.040 50.820 ;
        RECT 24.640 50.560 25.000 50.820 ;
        RECT 18.355 47.675 18.715 47.935 ;
        RECT 27.190 47.840 27.560 48.110 ;
        RECT 18.395 47.640 18.685 47.675 ;
      LAYER via ;
        RECT 12.285 50.560 12.545 50.820 ;
        RECT 13.250 50.560 13.510 50.820 ;
        RECT 14.205 50.560 14.465 50.820 ;
        RECT 15.165 50.560 15.425 50.820 ;
        RECT 16.125 50.560 16.385 50.820 ;
        RECT 17.085 50.560 17.345 50.820 ;
        RECT 19.890 50.560 20.150 50.820 ;
        RECT 20.855 50.560 21.115 50.820 ;
        RECT 21.810 50.560 22.070 50.820 ;
        RECT 22.770 50.560 23.030 50.820 ;
        RECT 23.730 50.560 23.990 50.820 ;
        RECT 24.690 50.560 24.950 50.820 ;
        RECT 18.405 47.675 18.665 47.935 ;
        RECT 27.245 47.845 27.505 48.105 ;
      LAYER met2 ;
        RECT 12.285 50.820 12.545 50.870 ;
        RECT 13.250 50.820 13.510 50.870 ;
        RECT 14.205 50.820 14.465 50.870 ;
        RECT 15.165 50.820 15.425 50.870 ;
        RECT 16.125 50.820 16.385 50.870 ;
        RECT 17.085 50.820 17.345 50.870 ;
        RECT 19.890 50.820 20.150 50.870 ;
        RECT 20.855 50.820 21.115 50.870 ;
        RECT 21.810 50.820 22.070 50.870 ;
        RECT 22.770 50.820 23.030 50.870 ;
        RECT 23.730 50.820 23.990 50.870 ;
        RECT 24.690 50.820 24.950 50.870 ;
        RECT 11.165 50.560 29.230 50.820 ;
        RECT 12.285 50.510 12.545 50.560 ;
        RECT 13.250 50.510 13.510 50.560 ;
        RECT 14.205 50.510 14.465 50.560 ;
        RECT 15.165 50.510 15.425 50.560 ;
        RECT 16.125 50.510 16.385 50.560 ;
        RECT 17.085 50.510 17.345 50.560 ;
        RECT 18.405 47.625 18.665 50.560 ;
        RECT 19.890 50.510 20.150 50.560 ;
        RECT 20.855 50.510 21.115 50.560 ;
        RECT 21.810 50.510 22.070 50.560 ;
        RECT 22.770 50.510 23.030 50.560 ;
        RECT 23.730 50.510 23.990 50.560 ;
        RECT 24.690 50.510 24.950 50.560 ;
        RECT 27.240 48.140 27.510 48.160 ;
        RECT 28.040 48.140 28.300 50.560 ;
        RECT 27.240 47.880 28.300 48.140 ;
        RECT 27.240 47.790 27.510 47.880 ;
    END
  END en_b[24]
  PIN en_b[25]
    DIRECTION INOUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 4.402500 ;
    PORT
      LAYER li1 ;
        RECT 12.250 44.165 12.580 44.335 ;
        RECT 13.210 44.165 13.540 44.335 ;
        RECT 14.170 44.165 14.500 44.335 ;
        RECT 15.130 44.165 15.460 44.335 ;
        RECT 16.090 44.165 16.420 44.335 ;
        RECT 17.050 44.165 17.380 44.335 ;
        RECT 19.855 44.165 20.185 44.335 ;
        RECT 20.815 44.165 21.145 44.335 ;
        RECT 21.775 44.165 22.105 44.335 ;
        RECT 22.735 44.165 23.065 44.335 ;
        RECT 23.695 44.165 24.025 44.335 ;
        RECT 24.655 44.165 24.985 44.335 ;
        RECT 27.100 41.450 27.430 41.690 ;
        RECT 18.375 41.235 18.705 41.405 ;
      LAYER mcon ;
        RECT 12.330 44.165 12.500 44.335 ;
        RECT 13.290 44.165 13.460 44.335 ;
        RECT 14.250 44.165 14.420 44.335 ;
        RECT 15.210 44.165 15.380 44.335 ;
        RECT 16.170 44.165 16.340 44.335 ;
        RECT 17.130 44.165 17.300 44.335 ;
        RECT 19.935 44.165 20.105 44.335 ;
        RECT 20.895 44.165 21.065 44.335 ;
        RECT 21.855 44.165 22.025 44.335 ;
        RECT 22.815 44.165 22.985 44.335 ;
        RECT 23.775 44.165 23.945 44.335 ;
        RECT 24.735 44.165 24.905 44.335 ;
        RECT 27.250 41.465 27.420 41.635 ;
        RECT 18.455 41.235 18.625 41.405 ;
      LAYER met1 ;
        RECT 12.235 44.125 12.595 44.385 ;
        RECT 13.200 44.125 13.560 44.385 ;
        RECT 14.155 44.125 14.515 44.385 ;
        RECT 15.115 44.125 15.475 44.385 ;
        RECT 16.075 44.125 16.435 44.385 ;
        RECT 17.035 44.125 17.395 44.385 ;
        RECT 19.840 44.125 20.200 44.385 ;
        RECT 20.805 44.125 21.165 44.385 ;
        RECT 21.760 44.125 22.120 44.385 ;
        RECT 22.720 44.125 23.080 44.385 ;
        RECT 23.680 44.125 24.040 44.385 ;
        RECT 24.640 44.125 25.000 44.385 ;
        RECT 18.355 41.240 18.715 41.500 ;
        RECT 27.190 41.405 27.560 41.675 ;
        RECT 18.395 41.205 18.685 41.240 ;
      LAYER via ;
        RECT 12.285 44.125 12.545 44.385 ;
        RECT 13.250 44.125 13.510 44.385 ;
        RECT 14.205 44.125 14.465 44.385 ;
        RECT 15.165 44.125 15.425 44.385 ;
        RECT 16.125 44.125 16.385 44.385 ;
        RECT 17.085 44.125 17.345 44.385 ;
        RECT 19.890 44.125 20.150 44.385 ;
        RECT 20.855 44.125 21.115 44.385 ;
        RECT 21.810 44.125 22.070 44.385 ;
        RECT 22.770 44.125 23.030 44.385 ;
        RECT 23.730 44.125 23.990 44.385 ;
        RECT 24.690 44.125 24.950 44.385 ;
        RECT 18.405 41.240 18.665 41.500 ;
        RECT 27.245 41.410 27.505 41.670 ;
      LAYER met2 ;
        RECT 12.285 44.385 12.545 44.435 ;
        RECT 13.250 44.385 13.510 44.435 ;
        RECT 14.205 44.385 14.465 44.435 ;
        RECT 15.165 44.385 15.425 44.435 ;
        RECT 16.125 44.385 16.385 44.435 ;
        RECT 17.085 44.385 17.345 44.435 ;
        RECT 19.890 44.385 20.150 44.435 ;
        RECT 20.855 44.385 21.115 44.435 ;
        RECT 21.810 44.385 22.070 44.435 ;
        RECT 22.770 44.385 23.030 44.435 ;
        RECT 23.730 44.385 23.990 44.435 ;
        RECT 24.690 44.385 24.950 44.435 ;
        RECT 11.165 44.125 29.230 44.385 ;
        RECT 12.285 44.075 12.545 44.125 ;
        RECT 13.250 44.075 13.510 44.125 ;
        RECT 14.205 44.075 14.465 44.125 ;
        RECT 15.165 44.075 15.425 44.125 ;
        RECT 16.125 44.075 16.385 44.125 ;
        RECT 17.085 44.075 17.345 44.125 ;
        RECT 18.405 41.190 18.665 44.125 ;
        RECT 19.890 44.075 20.150 44.125 ;
        RECT 20.855 44.075 21.115 44.125 ;
        RECT 21.810 44.075 22.070 44.125 ;
        RECT 22.770 44.075 23.030 44.125 ;
        RECT 23.730 44.075 23.990 44.125 ;
        RECT 24.690 44.075 24.950 44.125 ;
        RECT 27.240 41.705 27.510 41.725 ;
        RECT 28.040 41.705 28.300 44.125 ;
        RECT 27.240 41.445 28.300 41.705 ;
        RECT 27.240 41.355 27.510 41.445 ;
    END
  END en_b[25]
  PIN en_b[26]
    DIRECTION INOUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 4.402500 ;
    PORT
      LAYER li1 ;
        RECT 12.250 37.730 12.580 37.900 ;
        RECT 13.210 37.730 13.540 37.900 ;
        RECT 14.170 37.730 14.500 37.900 ;
        RECT 15.130 37.730 15.460 37.900 ;
        RECT 16.090 37.730 16.420 37.900 ;
        RECT 17.050 37.730 17.380 37.900 ;
        RECT 19.855 37.730 20.185 37.900 ;
        RECT 20.815 37.730 21.145 37.900 ;
        RECT 21.775 37.730 22.105 37.900 ;
        RECT 22.735 37.730 23.065 37.900 ;
        RECT 23.695 37.730 24.025 37.900 ;
        RECT 24.655 37.730 24.985 37.900 ;
        RECT 27.100 35.015 27.430 35.255 ;
        RECT 18.375 34.800 18.705 34.970 ;
      LAYER mcon ;
        RECT 12.330 37.730 12.500 37.900 ;
        RECT 13.290 37.730 13.460 37.900 ;
        RECT 14.250 37.730 14.420 37.900 ;
        RECT 15.210 37.730 15.380 37.900 ;
        RECT 16.170 37.730 16.340 37.900 ;
        RECT 17.130 37.730 17.300 37.900 ;
        RECT 19.935 37.730 20.105 37.900 ;
        RECT 20.895 37.730 21.065 37.900 ;
        RECT 21.855 37.730 22.025 37.900 ;
        RECT 22.815 37.730 22.985 37.900 ;
        RECT 23.775 37.730 23.945 37.900 ;
        RECT 24.735 37.730 24.905 37.900 ;
        RECT 27.250 35.030 27.420 35.200 ;
        RECT 18.455 34.800 18.625 34.970 ;
      LAYER met1 ;
        RECT 12.235 37.690 12.595 37.950 ;
        RECT 13.200 37.690 13.560 37.950 ;
        RECT 14.155 37.690 14.515 37.950 ;
        RECT 15.115 37.690 15.475 37.950 ;
        RECT 16.075 37.690 16.435 37.950 ;
        RECT 17.035 37.690 17.395 37.950 ;
        RECT 19.840 37.690 20.200 37.950 ;
        RECT 20.805 37.690 21.165 37.950 ;
        RECT 21.760 37.690 22.120 37.950 ;
        RECT 22.720 37.690 23.080 37.950 ;
        RECT 23.680 37.690 24.040 37.950 ;
        RECT 24.640 37.690 25.000 37.950 ;
        RECT 18.355 34.805 18.715 35.065 ;
        RECT 27.190 34.970 27.560 35.240 ;
        RECT 18.395 34.770 18.685 34.805 ;
      LAYER via ;
        RECT 12.285 37.690 12.545 37.950 ;
        RECT 13.250 37.690 13.510 37.950 ;
        RECT 14.205 37.690 14.465 37.950 ;
        RECT 15.165 37.690 15.425 37.950 ;
        RECT 16.125 37.690 16.385 37.950 ;
        RECT 17.085 37.690 17.345 37.950 ;
        RECT 19.890 37.690 20.150 37.950 ;
        RECT 20.855 37.690 21.115 37.950 ;
        RECT 21.810 37.690 22.070 37.950 ;
        RECT 22.770 37.690 23.030 37.950 ;
        RECT 23.730 37.690 23.990 37.950 ;
        RECT 24.690 37.690 24.950 37.950 ;
        RECT 18.405 34.805 18.665 35.065 ;
        RECT 27.245 34.975 27.505 35.235 ;
      LAYER met2 ;
        RECT 12.285 37.950 12.545 38.000 ;
        RECT 13.250 37.950 13.510 38.000 ;
        RECT 14.205 37.950 14.465 38.000 ;
        RECT 15.165 37.950 15.425 38.000 ;
        RECT 16.125 37.950 16.385 38.000 ;
        RECT 17.085 37.950 17.345 38.000 ;
        RECT 19.890 37.950 20.150 38.000 ;
        RECT 20.855 37.950 21.115 38.000 ;
        RECT 21.810 37.950 22.070 38.000 ;
        RECT 22.770 37.950 23.030 38.000 ;
        RECT 23.730 37.950 23.990 38.000 ;
        RECT 24.690 37.950 24.950 38.000 ;
        RECT 11.165 37.690 29.230 37.950 ;
        RECT 12.285 37.640 12.545 37.690 ;
        RECT 13.250 37.640 13.510 37.690 ;
        RECT 14.205 37.640 14.465 37.690 ;
        RECT 15.165 37.640 15.425 37.690 ;
        RECT 16.125 37.640 16.385 37.690 ;
        RECT 17.085 37.640 17.345 37.690 ;
        RECT 18.405 34.755 18.665 37.690 ;
        RECT 19.890 37.640 20.150 37.690 ;
        RECT 20.855 37.640 21.115 37.690 ;
        RECT 21.810 37.640 22.070 37.690 ;
        RECT 22.770 37.640 23.030 37.690 ;
        RECT 23.730 37.640 23.990 37.690 ;
        RECT 24.690 37.640 24.950 37.690 ;
        RECT 27.240 35.270 27.510 35.290 ;
        RECT 28.040 35.270 28.300 37.690 ;
        RECT 27.240 35.010 28.300 35.270 ;
        RECT 27.240 34.920 27.510 35.010 ;
    END
  END en_b[26]
  PIN en_b[27]
    DIRECTION INOUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 4.402500 ;
    PORT
      LAYER li1 ;
        RECT 12.250 31.295 12.580 31.465 ;
        RECT 13.210 31.295 13.540 31.465 ;
        RECT 14.170 31.295 14.500 31.465 ;
        RECT 15.130 31.295 15.460 31.465 ;
        RECT 16.090 31.295 16.420 31.465 ;
        RECT 17.050 31.295 17.380 31.465 ;
        RECT 19.855 31.295 20.185 31.465 ;
        RECT 20.815 31.295 21.145 31.465 ;
        RECT 21.775 31.295 22.105 31.465 ;
        RECT 22.735 31.295 23.065 31.465 ;
        RECT 23.695 31.295 24.025 31.465 ;
        RECT 24.655 31.295 24.985 31.465 ;
        RECT 27.100 28.580 27.430 28.820 ;
        RECT 18.375 28.365 18.705 28.535 ;
      LAYER mcon ;
        RECT 12.330 31.295 12.500 31.465 ;
        RECT 13.290 31.295 13.460 31.465 ;
        RECT 14.250 31.295 14.420 31.465 ;
        RECT 15.210 31.295 15.380 31.465 ;
        RECT 16.170 31.295 16.340 31.465 ;
        RECT 17.130 31.295 17.300 31.465 ;
        RECT 19.935 31.295 20.105 31.465 ;
        RECT 20.895 31.295 21.065 31.465 ;
        RECT 21.855 31.295 22.025 31.465 ;
        RECT 22.815 31.295 22.985 31.465 ;
        RECT 23.775 31.295 23.945 31.465 ;
        RECT 24.735 31.295 24.905 31.465 ;
        RECT 27.250 28.595 27.420 28.765 ;
        RECT 18.455 28.365 18.625 28.535 ;
      LAYER met1 ;
        RECT 12.235 31.255 12.595 31.515 ;
        RECT 13.200 31.255 13.560 31.515 ;
        RECT 14.155 31.255 14.515 31.515 ;
        RECT 15.115 31.255 15.475 31.515 ;
        RECT 16.075 31.255 16.435 31.515 ;
        RECT 17.035 31.255 17.395 31.515 ;
        RECT 19.840 31.255 20.200 31.515 ;
        RECT 20.805 31.255 21.165 31.515 ;
        RECT 21.760 31.255 22.120 31.515 ;
        RECT 22.720 31.255 23.080 31.515 ;
        RECT 23.680 31.255 24.040 31.515 ;
        RECT 24.640 31.255 25.000 31.515 ;
        RECT 18.355 28.370 18.715 28.630 ;
        RECT 27.190 28.535 27.560 28.805 ;
        RECT 18.395 28.335 18.685 28.370 ;
      LAYER via ;
        RECT 12.285 31.255 12.545 31.515 ;
        RECT 13.250 31.255 13.510 31.515 ;
        RECT 14.205 31.255 14.465 31.515 ;
        RECT 15.165 31.255 15.425 31.515 ;
        RECT 16.125 31.255 16.385 31.515 ;
        RECT 17.085 31.255 17.345 31.515 ;
        RECT 19.890 31.255 20.150 31.515 ;
        RECT 20.855 31.255 21.115 31.515 ;
        RECT 21.810 31.255 22.070 31.515 ;
        RECT 22.770 31.255 23.030 31.515 ;
        RECT 23.730 31.255 23.990 31.515 ;
        RECT 24.690 31.255 24.950 31.515 ;
        RECT 18.405 28.370 18.665 28.630 ;
        RECT 27.245 28.540 27.505 28.800 ;
      LAYER met2 ;
        RECT 12.285 31.515 12.545 31.565 ;
        RECT 13.250 31.515 13.510 31.565 ;
        RECT 14.205 31.515 14.465 31.565 ;
        RECT 15.165 31.515 15.425 31.565 ;
        RECT 16.125 31.515 16.385 31.565 ;
        RECT 17.085 31.515 17.345 31.565 ;
        RECT 19.890 31.515 20.150 31.565 ;
        RECT 20.855 31.515 21.115 31.565 ;
        RECT 21.810 31.515 22.070 31.565 ;
        RECT 22.770 31.515 23.030 31.565 ;
        RECT 23.730 31.515 23.990 31.565 ;
        RECT 24.690 31.515 24.950 31.565 ;
        RECT 11.165 31.255 29.230 31.515 ;
        RECT 12.285 31.205 12.545 31.255 ;
        RECT 13.250 31.205 13.510 31.255 ;
        RECT 14.205 31.205 14.465 31.255 ;
        RECT 15.165 31.205 15.425 31.255 ;
        RECT 16.125 31.205 16.385 31.255 ;
        RECT 17.085 31.205 17.345 31.255 ;
        RECT 18.405 28.320 18.665 31.255 ;
        RECT 19.890 31.205 20.150 31.255 ;
        RECT 20.855 31.205 21.115 31.255 ;
        RECT 21.810 31.205 22.070 31.255 ;
        RECT 22.770 31.205 23.030 31.255 ;
        RECT 23.730 31.205 23.990 31.255 ;
        RECT 24.690 31.205 24.950 31.255 ;
        RECT 27.240 28.835 27.510 28.855 ;
        RECT 28.040 28.835 28.300 31.255 ;
        RECT 27.240 28.575 28.300 28.835 ;
        RECT 27.240 28.485 27.510 28.575 ;
    END
  END en_b[27]
  PIN en_b[28]
    DIRECTION INOUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 4.402500 ;
    PORT
      LAYER li1 ;
        RECT 12.250 24.860 12.580 25.030 ;
        RECT 13.210 24.860 13.540 25.030 ;
        RECT 14.170 24.860 14.500 25.030 ;
        RECT 15.130 24.860 15.460 25.030 ;
        RECT 16.090 24.860 16.420 25.030 ;
        RECT 17.050 24.860 17.380 25.030 ;
        RECT 19.855 24.860 20.185 25.030 ;
        RECT 20.815 24.860 21.145 25.030 ;
        RECT 21.775 24.860 22.105 25.030 ;
        RECT 22.735 24.860 23.065 25.030 ;
        RECT 23.695 24.860 24.025 25.030 ;
        RECT 24.655 24.860 24.985 25.030 ;
        RECT 27.100 22.145 27.430 22.385 ;
        RECT 18.375 21.930 18.705 22.100 ;
      LAYER mcon ;
        RECT 12.330 24.860 12.500 25.030 ;
        RECT 13.290 24.860 13.460 25.030 ;
        RECT 14.250 24.860 14.420 25.030 ;
        RECT 15.210 24.860 15.380 25.030 ;
        RECT 16.170 24.860 16.340 25.030 ;
        RECT 17.130 24.860 17.300 25.030 ;
        RECT 19.935 24.860 20.105 25.030 ;
        RECT 20.895 24.860 21.065 25.030 ;
        RECT 21.855 24.860 22.025 25.030 ;
        RECT 22.815 24.860 22.985 25.030 ;
        RECT 23.775 24.860 23.945 25.030 ;
        RECT 24.735 24.860 24.905 25.030 ;
        RECT 27.250 22.160 27.420 22.330 ;
        RECT 18.455 21.930 18.625 22.100 ;
      LAYER met1 ;
        RECT 12.235 24.820 12.595 25.080 ;
        RECT 13.200 24.820 13.560 25.080 ;
        RECT 14.155 24.820 14.515 25.080 ;
        RECT 15.115 24.820 15.475 25.080 ;
        RECT 16.075 24.820 16.435 25.080 ;
        RECT 17.035 24.820 17.395 25.080 ;
        RECT 19.840 24.820 20.200 25.080 ;
        RECT 20.805 24.820 21.165 25.080 ;
        RECT 21.760 24.820 22.120 25.080 ;
        RECT 22.720 24.820 23.080 25.080 ;
        RECT 23.680 24.820 24.040 25.080 ;
        RECT 24.640 24.820 25.000 25.080 ;
        RECT 18.355 21.935 18.715 22.195 ;
        RECT 27.190 22.100 27.560 22.370 ;
        RECT 18.395 21.900 18.685 21.935 ;
      LAYER via ;
        RECT 12.285 24.820 12.545 25.080 ;
        RECT 13.250 24.820 13.510 25.080 ;
        RECT 14.205 24.820 14.465 25.080 ;
        RECT 15.165 24.820 15.425 25.080 ;
        RECT 16.125 24.820 16.385 25.080 ;
        RECT 17.085 24.820 17.345 25.080 ;
        RECT 19.890 24.820 20.150 25.080 ;
        RECT 20.855 24.820 21.115 25.080 ;
        RECT 21.810 24.820 22.070 25.080 ;
        RECT 22.770 24.820 23.030 25.080 ;
        RECT 23.730 24.820 23.990 25.080 ;
        RECT 24.690 24.820 24.950 25.080 ;
        RECT 18.405 21.935 18.665 22.195 ;
        RECT 27.245 22.105 27.505 22.365 ;
      LAYER met2 ;
        RECT 12.285 25.080 12.545 25.130 ;
        RECT 13.250 25.080 13.510 25.130 ;
        RECT 14.205 25.080 14.465 25.130 ;
        RECT 15.165 25.080 15.425 25.130 ;
        RECT 16.125 25.080 16.385 25.130 ;
        RECT 17.085 25.080 17.345 25.130 ;
        RECT 19.890 25.080 20.150 25.130 ;
        RECT 20.855 25.080 21.115 25.130 ;
        RECT 21.810 25.080 22.070 25.130 ;
        RECT 22.770 25.080 23.030 25.130 ;
        RECT 23.730 25.080 23.990 25.130 ;
        RECT 24.690 25.080 24.950 25.130 ;
        RECT 11.165 24.820 29.230 25.080 ;
        RECT 12.285 24.770 12.545 24.820 ;
        RECT 13.250 24.770 13.510 24.820 ;
        RECT 14.205 24.770 14.465 24.820 ;
        RECT 15.165 24.770 15.425 24.820 ;
        RECT 16.125 24.770 16.385 24.820 ;
        RECT 17.085 24.770 17.345 24.820 ;
        RECT 18.405 21.885 18.665 24.820 ;
        RECT 19.890 24.770 20.150 24.820 ;
        RECT 20.855 24.770 21.115 24.820 ;
        RECT 21.810 24.770 22.070 24.820 ;
        RECT 22.770 24.770 23.030 24.820 ;
        RECT 23.730 24.770 23.990 24.820 ;
        RECT 24.690 24.770 24.950 24.820 ;
        RECT 27.240 22.400 27.510 22.420 ;
        RECT 28.040 22.400 28.300 24.820 ;
        RECT 27.240 22.140 28.300 22.400 ;
        RECT 27.240 22.050 27.510 22.140 ;
    END
  END en_b[28]
  PIN en_b[29]
    DIRECTION INOUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 4.402500 ;
    PORT
      LAYER li1 ;
        RECT 12.250 18.425 12.580 18.595 ;
        RECT 13.210 18.425 13.540 18.595 ;
        RECT 14.170 18.425 14.500 18.595 ;
        RECT 15.130 18.425 15.460 18.595 ;
        RECT 16.090 18.425 16.420 18.595 ;
        RECT 17.050 18.425 17.380 18.595 ;
        RECT 19.855 18.425 20.185 18.595 ;
        RECT 20.815 18.425 21.145 18.595 ;
        RECT 21.775 18.425 22.105 18.595 ;
        RECT 22.735 18.425 23.065 18.595 ;
        RECT 23.695 18.425 24.025 18.595 ;
        RECT 24.655 18.425 24.985 18.595 ;
        RECT 27.100 15.710 27.430 15.950 ;
        RECT 18.375 15.495 18.705 15.665 ;
      LAYER mcon ;
        RECT 12.330 18.425 12.500 18.595 ;
        RECT 13.290 18.425 13.460 18.595 ;
        RECT 14.250 18.425 14.420 18.595 ;
        RECT 15.210 18.425 15.380 18.595 ;
        RECT 16.170 18.425 16.340 18.595 ;
        RECT 17.130 18.425 17.300 18.595 ;
        RECT 19.935 18.425 20.105 18.595 ;
        RECT 20.895 18.425 21.065 18.595 ;
        RECT 21.855 18.425 22.025 18.595 ;
        RECT 22.815 18.425 22.985 18.595 ;
        RECT 23.775 18.425 23.945 18.595 ;
        RECT 24.735 18.425 24.905 18.595 ;
        RECT 27.250 15.725 27.420 15.895 ;
        RECT 18.455 15.495 18.625 15.665 ;
      LAYER met1 ;
        RECT 12.235 18.385 12.595 18.645 ;
        RECT 13.200 18.385 13.560 18.645 ;
        RECT 14.155 18.385 14.515 18.645 ;
        RECT 15.115 18.385 15.475 18.645 ;
        RECT 16.075 18.385 16.435 18.645 ;
        RECT 17.035 18.385 17.395 18.645 ;
        RECT 19.840 18.385 20.200 18.645 ;
        RECT 20.805 18.385 21.165 18.645 ;
        RECT 21.760 18.385 22.120 18.645 ;
        RECT 22.720 18.385 23.080 18.645 ;
        RECT 23.680 18.385 24.040 18.645 ;
        RECT 24.640 18.385 25.000 18.645 ;
        RECT 18.355 15.500 18.715 15.760 ;
        RECT 27.190 15.665 27.560 15.935 ;
        RECT 18.395 15.465 18.685 15.500 ;
      LAYER via ;
        RECT 12.285 18.385 12.545 18.645 ;
        RECT 13.250 18.385 13.510 18.645 ;
        RECT 14.205 18.385 14.465 18.645 ;
        RECT 15.165 18.385 15.425 18.645 ;
        RECT 16.125 18.385 16.385 18.645 ;
        RECT 17.085 18.385 17.345 18.645 ;
        RECT 19.890 18.385 20.150 18.645 ;
        RECT 20.855 18.385 21.115 18.645 ;
        RECT 21.810 18.385 22.070 18.645 ;
        RECT 22.770 18.385 23.030 18.645 ;
        RECT 23.730 18.385 23.990 18.645 ;
        RECT 24.690 18.385 24.950 18.645 ;
        RECT 18.405 15.500 18.665 15.760 ;
        RECT 27.245 15.670 27.505 15.930 ;
      LAYER met2 ;
        RECT 12.285 18.645 12.545 18.695 ;
        RECT 13.250 18.645 13.510 18.695 ;
        RECT 14.205 18.645 14.465 18.695 ;
        RECT 15.165 18.645 15.425 18.695 ;
        RECT 16.125 18.645 16.385 18.695 ;
        RECT 17.085 18.645 17.345 18.695 ;
        RECT 19.890 18.645 20.150 18.695 ;
        RECT 20.855 18.645 21.115 18.695 ;
        RECT 21.810 18.645 22.070 18.695 ;
        RECT 22.770 18.645 23.030 18.695 ;
        RECT 23.730 18.645 23.990 18.695 ;
        RECT 24.690 18.645 24.950 18.695 ;
        RECT 11.165 18.385 29.230 18.645 ;
        RECT 12.285 18.335 12.545 18.385 ;
        RECT 13.250 18.335 13.510 18.385 ;
        RECT 14.205 18.335 14.465 18.385 ;
        RECT 15.165 18.335 15.425 18.385 ;
        RECT 16.125 18.335 16.385 18.385 ;
        RECT 17.085 18.335 17.345 18.385 ;
        RECT 18.405 15.450 18.665 18.385 ;
        RECT 19.890 18.335 20.150 18.385 ;
        RECT 20.855 18.335 21.115 18.385 ;
        RECT 21.810 18.335 22.070 18.385 ;
        RECT 22.770 18.335 23.030 18.385 ;
        RECT 23.730 18.335 23.990 18.385 ;
        RECT 24.690 18.335 24.950 18.385 ;
        RECT 27.240 15.965 27.510 15.985 ;
        RECT 28.040 15.965 28.300 18.385 ;
        RECT 27.240 15.705 28.300 15.965 ;
        RECT 27.240 15.615 27.510 15.705 ;
    END
  END en_b[29]
  PIN en_b[30]
    DIRECTION INOUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 4.402500 ;
    PORT
      LAYER li1 ;
        RECT 12.250 11.990 12.580 12.160 ;
        RECT 13.210 11.990 13.540 12.160 ;
        RECT 14.170 11.990 14.500 12.160 ;
        RECT 15.130 11.990 15.460 12.160 ;
        RECT 16.090 11.990 16.420 12.160 ;
        RECT 17.050 11.990 17.380 12.160 ;
        RECT 19.855 11.990 20.185 12.160 ;
        RECT 20.815 11.990 21.145 12.160 ;
        RECT 21.775 11.990 22.105 12.160 ;
        RECT 22.735 11.990 23.065 12.160 ;
        RECT 23.695 11.990 24.025 12.160 ;
        RECT 24.655 11.990 24.985 12.160 ;
        RECT 27.100 9.275 27.430 9.515 ;
        RECT 18.375 9.060 18.705 9.230 ;
      LAYER mcon ;
        RECT 12.330 11.990 12.500 12.160 ;
        RECT 13.290 11.990 13.460 12.160 ;
        RECT 14.250 11.990 14.420 12.160 ;
        RECT 15.210 11.990 15.380 12.160 ;
        RECT 16.170 11.990 16.340 12.160 ;
        RECT 17.130 11.990 17.300 12.160 ;
        RECT 19.935 11.990 20.105 12.160 ;
        RECT 20.895 11.990 21.065 12.160 ;
        RECT 21.855 11.990 22.025 12.160 ;
        RECT 22.815 11.990 22.985 12.160 ;
        RECT 23.775 11.990 23.945 12.160 ;
        RECT 24.735 11.990 24.905 12.160 ;
        RECT 27.250 9.290 27.420 9.460 ;
        RECT 18.455 9.060 18.625 9.230 ;
      LAYER met1 ;
        RECT 12.235 11.950 12.595 12.210 ;
        RECT 13.200 11.950 13.560 12.210 ;
        RECT 14.155 11.950 14.515 12.210 ;
        RECT 15.115 11.950 15.475 12.210 ;
        RECT 16.075 11.950 16.435 12.210 ;
        RECT 17.035 11.950 17.395 12.210 ;
        RECT 19.840 11.950 20.200 12.210 ;
        RECT 20.805 11.950 21.165 12.210 ;
        RECT 21.760 11.950 22.120 12.210 ;
        RECT 22.720 11.950 23.080 12.210 ;
        RECT 23.680 11.950 24.040 12.210 ;
        RECT 24.640 11.950 25.000 12.210 ;
        RECT 18.355 9.065 18.715 9.325 ;
        RECT 27.190 9.230 27.560 9.500 ;
        RECT 18.395 9.030 18.685 9.065 ;
      LAYER via ;
        RECT 12.285 11.950 12.545 12.210 ;
        RECT 13.250 11.950 13.510 12.210 ;
        RECT 14.205 11.950 14.465 12.210 ;
        RECT 15.165 11.950 15.425 12.210 ;
        RECT 16.125 11.950 16.385 12.210 ;
        RECT 17.085 11.950 17.345 12.210 ;
        RECT 19.890 11.950 20.150 12.210 ;
        RECT 20.855 11.950 21.115 12.210 ;
        RECT 21.810 11.950 22.070 12.210 ;
        RECT 22.770 11.950 23.030 12.210 ;
        RECT 23.730 11.950 23.990 12.210 ;
        RECT 24.690 11.950 24.950 12.210 ;
        RECT 18.405 9.065 18.665 9.325 ;
        RECT 27.245 9.235 27.505 9.495 ;
      LAYER met2 ;
        RECT 12.285 12.210 12.545 12.260 ;
        RECT 13.250 12.210 13.510 12.260 ;
        RECT 14.205 12.210 14.465 12.260 ;
        RECT 15.165 12.210 15.425 12.260 ;
        RECT 16.125 12.210 16.385 12.260 ;
        RECT 17.085 12.210 17.345 12.260 ;
        RECT 19.890 12.210 20.150 12.260 ;
        RECT 20.855 12.210 21.115 12.260 ;
        RECT 21.810 12.210 22.070 12.260 ;
        RECT 22.770 12.210 23.030 12.260 ;
        RECT 23.730 12.210 23.990 12.260 ;
        RECT 24.690 12.210 24.950 12.260 ;
        RECT 11.165 11.950 29.230 12.210 ;
        RECT 12.285 11.900 12.545 11.950 ;
        RECT 13.250 11.900 13.510 11.950 ;
        RECT 14.205 11.900 14.465 11.950 ;
        RECT 15.165 11.900 15.425 11.950 ;
        RECT 16.125 11.900 16.385 11.950 ;
        RECT 17.085 11.900 17.345 11.950 ;
        RECT 18.405 9.015 18.665 11.950 ;
        RECT 19.890 11.900 20.150 11.950 ;
        RECT 20.855 11.900 21.115 11.950 ;
        RECT 21.810 11.900 22.070 11.950 ;
        RECT 22.770 11.900 23.030 11.950 ;
        RECT 23.730 11.900 23.990 11.950 ;
        RECT 24.690 11.900 24.950 11.950 ;
        RECT 27.240 9.530 27.510 9.550 ;
        RECT 28.040 9.530 28.300 11.950 ;
        RECT 27.240 9.270 28.300 9.530 ;
        RECT 27.240 9.180 27.510 9.270 ;
    END
  END en_b[30]
  PIN en_b[31]
    DIRECTION INOUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 4.402500 ;
    PORT
      LAYER li1 ;
        RECT 12.250 5.555 12.580 5.725 ;
        RECT 13.210 5.555 13.540 5.725 ;
        RECT 14.170 5.555 14.500 5.725 ;
        RECT 15.130 5.555 15.460 5.725 ;
        RECT 16.090 5.555 16.420 5.725 ;
        RECT 17.050 5.555 17.380 5.725 ;
        RECT 19.855 5.555 20.185 5.725 ;
        RECT 20.815 5.555 21.145 5.725 ;
        RECT 21.775 5.555 22.105 5.725 ;
        RECT 22.735 5.555 23.065 5.725 ;
        RECT 23.695 5.555 24.025 5.725 ;
        RECT 24.655 5.555 24.985 5.725 ;
        RECT 27.100 2.840 27.430 3.080 ;
        RECT 18.375 2.625 18.705 2.795 ;
      LAYER mcon ;
        RECT 12.330 5.555 12.500 5.725 ;
        RECT 13.290 5.555 13.460 5.725 ;
        RECT 14.250 5.555 14.420 5.725 ;
        RECT 15.210 5.555 15.380 5.725 ;
        RECT 16.170 5.555 16.340 5.725 ;
        RECT 17.130 5.555 17.300 5.725 ;
        RECT 19.935 5.555 20.105 5.725 ;
        RECT 20.895 5.555 21.065 5.725 ;
        RECT 21.855 5.555 22.025 5.725 ;
        RECT 22.815 5.555 22.985 5.725 ;
        RECT 23.775 5.555 23.945 5.725 ;
        RECT 24.735 5.555 24.905 5.725 ;
        RECT 27.250 2.855 27.420 3.025 ;
        RECT 18.455 2.625 18.625 2.795 ;
      LAYER met1 ;
        RECT 12.235 5.515 12.595 5.775 ;
        RECT 13.200 5.515 13.560 5.775 ;
        RECT 14.155 5.515 14.515 5.775 ;
        RECT 15.115 5.515 15.475 5.775 ;
        RECT 16.075 5.515 16.435 5.775 ;
        RECT 17.035 5.515 17.395 5.775 ;
        RECT 19.840 5.515 20.200 5.775 ;
        RECT 20.805 5.515 21.165 5.775 ;
        RECT 21.760 5.515 22.120 5.775 ;
        RECT 22.720 5.515 23.080 5.775 ;
        RECT 23.680 5.515 24.040 5.775 ;
        RECT 24.640 5.515 25.000 5.775 ;
        RECT 18.355 2.630 18.715 2.890 ;
        RECT 27.190 2.795 27.560 3.065 ;
        RECT 18.395 2.595 18.685 2.630 ;
      LAYER via ;
        RECT 12.285 5.515 12.545 5.775 ;
        RECT 13.250 5.515 13.510 5.775 ;
        RECT 14.205 5.515 14.465 5.775 ;
        RECT 15.165 5.515 15.425 5.775 ;
        RECT 16.125 5.515 16.385 5.775 ;
        RECT 17.085 5.515 17.345 5.775 ;
        RECT 19.890 5.515 20.150 5.775 ;
        RECT 20.855 5.515 21.115 5.775 ;
        RECT 21.810 5.515 22.070 5.775 ;
        RECT 22.770 5.515 23.030 5.775 ;
        RECT 23.730 5.515 23.990 5.775 ;
        RECT 24.690 5.515 24.950 5.775 ;
        RECT 18.405 2.630 18.665 2.890 ;
        RECT 27.245 2.800 27.505 3.060 ;
      LAYER met2 ;
        RECT 12.285 5.775 12.545 5.825 ;
        RECT 13.250 5.775 13.510 5.825 ;
        RECT 14.205 5.775 14.465 5.825 ;
        RECT 15.165 5.775 15.425 5.825 ;
        RECT 16.125 5.775 16.385 5.825 ;
        RECT 17.085 5.775 17.345 5.825 ;
        RECT 19.890 5.775 20.150 5.825 ;
        RECT 20.855 5.775 21.115 5.825 ;
        RECT 21.810 5.775 22.070 5.825 ;
        RECT 22.770 5.775 23.030 5.825 ;
        RECT 23.730 5.775 23.990 5.825 ;
        RECT 24.690 5.775 24.950 5.825 ;
        RECT 11.165 5.515 29.230 5.775 ;
        RECT 12.285 5.465 12.545 5.515 ;
        RECT 13.250 5.465 13.510 5.515 ;
        RECT 14.205 5.465 14.465 5.515 ;
        RECT 15.165 5.465 15.425 5.515 ;
        RECT 16.125 5.465 16.385 5.515 ;
        RECT 17.085 5.465 17.345 5.515 ;
        RECT 18.405 2.580 18.665 5.515 ;
        RECT 19.890 5.465 20.150 5.515 ;
        RECT 20.855 5.465 21.115 5.515 ;
        RECT 21.810 5.465 22.070 5.515 ;
        RECT 22.770 5.465 23.030 5.515 ;
        RECT 23.730 5.465 23.990 5.515 ;
        RECT 24.690 5.465 24.950 5.515 ;
        RECT 27.240 3.095 27.510 3.115 ;
        RECT 28.040 3.095 28.300 5.515 ;
        RECT 27.240 2.835 28.300 3.095 ;
        RECT 27.240 2.745 27.510 2.835 ;
    END
  END en_b[31]
  PIN s_en
    DIRECTION INOUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 24.959999 ;
    PORT
      LAYER li1 ;
        RECT 1.485 200.980 1.815 201.150 ;
        RECT 2.445 200.980 2.775 201.150 ;
        RECT 3.405 200.980 3.735 201.150 ;
        RECT 4.365 200.980 4.695 201.150 ;
        RECT 5.325 200.980 5.655 201.150 ;
        RECT 6.285 200.980 6.615 201.150 ;
        RECT 1.485 194.545 1.815 194.715 ;
        RECT 2.445 194.545 2.775 194.715 ;
        RECT 3.405 194.545 3.735 194.715 ;
        RECT 4.365 194.545 4.695 194.715 ;
        RECT 5.325 194.545 5.655 194.715 ;
        RECT 6.285 194.545 6.615 194.715 ;
        RECT 1.485 188.110 1.815 188.280 ;
        RECT 2.445 188.110 2.775 188.280 ;
        RECT 3.405 188.110 3.735 188.280 ;
        RECT 4.365 188.110 4.695 188.280 ;
        RECT 5.325 188.110 5.655 188.280 ;
        RECT 6.285 188.110 6.615 188.280 ;
        RECT 1.485 181.675 1.815 181.845 ;
        RECT 2.445 181.675 2.775 181.845 ;
        RECT 3.405 181.675 3.735 181.845 ;
        RECT 4.365 181.675 4.695 181.845 ;
        RECT 5.325 181.675 5.655 181.845 ;
        RECT 6.285 181.675 6.615 181.845 ;
        RECT 1.485 175.240 1.815 175.410 ;
        RECT 2.445 175.240 2.775 175.410 ;
        RECT 3.405 175.240 3.735 175.410 ;
        RECT 4.365 175.240 4.695 175.410 ;
        RECT 5.325 175.240 5.655 175.410 ;
        RECT 6.285 175.240 6.615 175.410 ;
        RECT 1.485 168.805 1.815 168.975 ;
        RECT 2.445 168.805 2.775 168.975 ;
        RECT 3.405 168.805 3.735 168.975 ;
        RECT 4.365 168.805 4.695 168.975 ;
        RECT 5.325 168.805 5.655 168.975 ;
        RECT 6.285 168.805 6.615 168.975 ;
        RECT 1.485 162.370 1.815 162.540 ;
        RECT 2.445 162.370 2.775 162.540 ;
        RECT 3.405 162.370 3.735 162.540 ;
        RECT 4.365 162.370 4.695 162.540 ;
        RECT 5.325 162.370 5.655 162.540 ;
        RECT 6.285 162.370 6.615 162.540 ;
        RECT 1.485 155.935 1.815 156.105 ;
        RECT 2.445 155.935 2.775 156.105 ;
        RECT 3.405 155.935 3.735 156.105 ;
        RECT 4.365 155.935 4.695 156.105 ;
        RECT 5.325 155.935 5.655 156.105 ;
        RECT 6.285 155.935 6.615 156.105 ;
        RECT 1.485 149.500 1.815 149.670 ;
        RECT 2.445 149.500 2.775 149.670 ;
        RECT 3.405 149.500 3.735 149.670 ;
        RECT 4.365 149.500 4.695 149.670 ;
        RECT 5.325 149.500 5.655 149.670 ;
        RECT 6.285 149.500 6.615 149.670 ;
        RECT 1.485 143.065 1.815 143.235 ;
        RECT 2.445 143.065 2.775 143.235 ;
        RECT 3.405 143.065 3.735 143.235 ;
        RECT 4.365 143.065 4.695 143.235 ;
        RECT 5.325 143.065 5.655 143.235 ;
        RECT 6.285 143.065 6.615 143.235 ;
        RECT 1.485 136.630 1.815 136.800 ;
        RECT 2.445 136.630 2.775 136.800 ;
        RECT 3.405 136.630 3.735 136.800 ;
        RECT 4.365 136.630 4.695 136.800 ;
        RECT 5.325 136.630 5.655 136.800 ;
        RECT 6.285 136.630 6.615 136.800 ;
        RECT 1.485 130.195 1.815 130.365 ;
        RECT 2.445 130.195 2.775 130.365 ;
        RECT 3.405 130.195 3.735 130.365 ;
        RECT 4.365 130.195 4.695 130.365 ;
        RECT 5.325 130.195 5.655 130.365 ;
        RECT 6.285 130.195 6.615 130.365 ;
        RECT 1.485 123.760 1.815 123.930 ;
        RECT 2.445 123.760 2.775 123.930 ;
        RECT 3.405 123.760 3.735 123.930 ;
        RECT 4.365 123.760 4.695 123.930 ;
        RECT 5.325 123.760 5.655 123.930 ;
        RECT 6.285 123.760 6.615 123.930 ;
        RECT 1.485 117.325 1.815 117.495 ;
        RECT 2.445 117.325 2.775 117.495 ;
        RECT 3.405 117.325 3.735 117.495 ;
        RECT 4.365 117.325 4.695 117.495 ;
        RECT 5.325 117.325 5.655 117.495 ;
        RECT 6.285 117.325 6.615 117.495 ;
        RECT 1.485 110.890 1.815 111.060 ;
        RECT 2.445 110.890 2.775 111.060 ;
        RECT 3.405 110.890 3.735 111.060 ;
        RECT 4.365 110.890 4.695 111.060 ;
        RECT 5.325 110.890 5.655 111.060 ;
        RECT 6.285 110.890 6.615 111.060 ;
        RECT 1.485 104.455 1.815 104.625 ;
        RECT 2.445 104.455 2.775 104.625 ;
        RECT 3.405 104.455 3.735 104.625 ;
        RECT 4.365 104.455 4.695 104.625 ;
        RECT 5.325 104.455 5.655 104.625 ;
        RECT 6.285 104.455 6.615 104.625 ;
        RECT 1.485 98.020 1.815 98.190 ;
        RECT 2.445 98.020 2.775 98.190 ;
        RECT 3.405 98.020 3.735 98.190 ;
        RECT 4.365 98.020 4.695 98.190 ;
        RECT 5.325 98.020 5.655 98.190 ;
        RECT 6.285 98.020 6.615 98.190 ;
        RECT 1.485 91.585 1.815 91.755 ;
        RECT 2.445 91.585 2.775 91.755 ;
        RECT 3.405 91.585 3.735 91.755 ;
        RECT 4.365 91.585 4.695 91.755 ;
        RECT 5.325 91.585 5.655 91.755 ;
        RECT 6.285 91.585 6.615 91.755 ;
        RECT 1.485 85.150 1.815 85.320 ;
        RECT 2.445 85.150 2.775 85.320 ;
        RECT 3.405 85.150 3.735 85.320 ;
        RECT 4.365 85.150 4.695 85.320 ;
        RECT 5.325 85.150 5.655 85.320 ;
        RECT 6.285 85.150 6.615 85.320 ;
        RECT 1.485 78.715 1.815 78.885 ;
        RECT 2.445 78.715 2.775 78.885 ;
        RECT 3.405 78.715 3.735 78.885 ;
        RECT 4.365 78.715 4.695 78.885 ;
        RECT 5.325 78.715 5.655 78.885 ;
        RECT 6.285 78.715 6.615 78.885 ;
        RECT 1.485 72.280 1.815 72.450 ;
        RECT 2.445 72.280 2.775 72.450 ;
        RECT 3.405 72.280 3.735 72.450 ;
        RECT 4.365 72.280 4.695 72.450 ;
        RECT 5.325 72.280 5.655 72.450 ;
        RECT 6.285 72.280 6.615 72.450 ;
        RECT 1.485 65.845 1.815 66.015 ;
        RECT 2.445 65.845 2.775 66.015 ;
        RECT 3.405 65.845 3.735 66.015 ;
        RECT 4.365 65.845 4.695 66.015 ;
        RECT 5.325 65.845 5.655 66.015 ;
        RECT 6.285 65.845 6.615 66.015 ;
        RECT 1.485 59.410 1.815 59.580 ;
        RECT 2.445 59.410 2.775 59.580 ;
        RECT 3.405 59.410 3.735 59.580 ;
        RECT 4.365 59.410 4.695 59.580 ;
        RECT 5.325 59.410 5.655 59.580 ;
        RECT 6.285 59.410 6.615 59.580 ;
        RECT 1.485 52.975 1.815 53.145 ;
        RECT 2.445 52.975 2.775 53.145 ;
        RECT 3.405 52.975 3.735 53.145 ;
        RECT 4.365 52.975 4.695 53.145 ;
        RECT 5.325 52.975 5.655 53.145 ;
        RECT 6.285 52.975 6.615 53.145 ;
        RECT 1.485 46.540 1.815 46.710 ;
        RECT 2.445 46.540 2.775 46.710 ;
        RECT 3.405 46.540 3.735 46.710 ;
        RECT 4.365 46.540 4.695 46.710 ;
        RECT 5.325 46.540 5.655 46.710 ;
        RECT 6.285 46.540 6.615 46.710 ;
        RECT 1.485 40.105 1.815 40.275 ;
        RECT 2.445 40.105 2.775 40.275 ;
        RECT 3.405 40.105 3.735 40.275 ;
        RECT 4.365 40.105 4.695 40.275 ;
        RECT 5.325 40.105 5.655 40.275 ;
        RECT 6.285 40.105 6.615 40.275 ;
        RECT 1.485 33.670 1.815 33.840 ;
        RECT 2.445 33.670 2.775 33.840 ;
        RECT 3.405 33.670 3.735 33.840 ;
        RECT 4.365 33.670 4.695 33.840 ;
        RECT 5.325 33.670 5.655 33.840 ;
        RECT 6.285 33.670 6.615 33.840 ;
        RECT 1.485 27.235 1.815 27.405 ;
        RECT 2.445 27.235 2.775 27.405 ;
        RECT 3.405 27.235 3.735 27.405 ;
        RECT 4.365 27.235 4.695 27.405 ;
        RECT 5.325 27.235 5.655 27.405 ;
        RECT 6.285 27.235 6.615 27.405 ;
        RECT 1.485 20.800 1.815 20.970 ;
        RECT 2.445 20.800 2.775 20.970 ;
        RECT 3.405 20.800 3.735 20.970 ;
        RECT 4.365 20.800 4.695 20.970 ;
        RECT 5.325 20.800 5.655 20.970 ;
        RECT 6.285 20.800 6.615 20.970 ;
        RECT 1.485 14.365 1.815 14.535 ;
        RECT 2.445 14.365 2.775 14.535 ;
        RECT 3.405 14.365 3.735 14.535 ;
        RECT 4.365 14.365 4.695 14.535 ;
        RECT 5.325 14.365 5.655 14.535 ;
        RECT 6.285 14.365 6.615 14.535 ;
        RECT 1.485 7.930 1.815 8.100 ;
        RECT 2.445 7.930 2.775 8.100 ;
        RECT 3.405 7.930 3.735 8.100 ;
        RECT 4.365 7.930 4.695 8.100 ;
        RECT 5.325 7.930 5.655 8.100 ;
        RECT 6.285 7.930 6.615 8.100 ;
        RECT 1.485 1.495 1.815 1.665 ;
        RECT 2.445 1.495 2.775 1.665 ;
        RECT 3.405 1.495 3.735 1.665 ;
        RECT 4.365 1.495 4.695 1.665 ;
        RECT 5.325 1.495 5.655 1.665 ;
        RECT 6.285 1.495 6.615 1.665 ;
      LAYER mcon ;
        RECT 1.565 200.980 1.735 201.150 ;
        RECT 2.525 200.980 2.695 201.150 ;
        RECT 3.485 200.980 3.655 201.150 ;
        RECT 4.445 200.980 4.615 201.150 ;
        RECT 5.405 200.980 5.575 201.150 ;
        RECT 6.365 200.980 6.535 201.150 ;
        RECT 1.565 194.545 1.735 194.715 ;
        RECT 2.525 194.545 2.695 194.715 ;
        RECT 3.485 194.545 3.655 194.715 ;
        RECT 4.445 194.545 4.615 194.715 ;
        RECT 5.405 194.545 5.575 194.715 ;
        RECT 6.365 194.545 6.535 194.715 ;
        RECT 1.565 188.110 1.735 188.280 ;
        RECT 2.525 188.110 2.695 188.280 ;
        RECT 3.485 188.110 3.655 188.280 ;
        RECT 4.445 188.110 4.615 188.280 ;
        RECT 5.405 188.110 5.575 188.280 ;
        RECT 6.365 188.110 6.535 188.280 ;
        RECT 1.565 181.675 1.735 181.845 ;
        RECT 2.525 181.675 2.695 181.845 ;
        RECT 3.485 181.675 3.655 181.845 ;
        RECT 4.445 181.675 4.615 181.845 ;
        RECT 5.405 181.675 5.575 181.845 ;
        RECT 6.365 181.675 6.535 181.845 ;
        RECT 1.565 175.240 1.735 175.410 ;
        RECT 2.525 175.240 2.695 175.410 ;
        RECT 3.485 175.240 3.655 175.410 ;
        RECT 4.445 175.240 4.615 175.410 ;
        RECT 5.405 175.240 5.575 175.410 ;
        RECT 6.365 175.240 6.535 175.410 ;
        RECT 1.565 168.805 1.735 168.975 ;
        RECT 2.525 168.805 2.695 168.975 ;
        RECT 3.485 168.805 3.655 168.975 ;
        RECT 4.445 168.805 4.615 168.975 ;
        RECT 5.405 168.805 5.575 168.975 ;
        RECT 6.365 168.805 6.535 168.975 ;
        RECT 1.565 162.370 1.735 162.540 ;
        RECT 2.525 162.370 2.695 162.540 ;
        RECT 3.485 162.370 3.655 162.540 ;
        RECT 4.445 162.370 4.615 162.540 ;
        RECT 5.405 162.370 5.575 162.540 ;
        RECT 6.365 162.370 6.535 162.540 ;
        RECT 1.565 155.935 1.735 156.105 ;
        RECT 2.525 155.935 2.695 156.105 ;
        RECT 3.485 155.935 3.655 156.105 ;
        RECT 4.445 155.935 4.615 156.105 ;
        RECT 5.405 155.935 5.575 156.105 ;
        RECT 6.365 155.935 6.535 156.105 ;
        RECT 1.565 149.500 1.735 149.670 ;
        RECT 2.525 149.500 2.695 149.670 ;
        RECT 3.485 149.500 3.655 149.670 ;
        RECT 4.445 149.500 4.615 149.670 ;
        RECT 5.405 149.500 5.575 149.670 ;
        RECT 6.365 149.500 6.535 149.670 ;
        RECT 1.565 143.065 1.735 143.235 ;
        RECT 2.525 143.065 2.695 143.235 ;
        RECT 3.485 143.065 3.655 143.235 ;
        RECT 4.445 143.065 4.615 143.235 ;
        RECT 5.405 143.065 5.575 143.235 ;
        RECT 6.365 143.065 6.535 143.235 ;
        RECT 1.565 136.630 1.735 136.800 ;
        RECT 2.525 136.630 2.695 136.800 ;
        RECT 3.485 136.630 3.655 136.800 ;
        RECT 4.445 136.630 4.615 136.800 ;
        RECT 5.405 136.630 5.575 136.800 ;
        RECT 6.365 136.630 6.535 136.800 ;
        RECT 1.565 130.195 1.735 130.365 ;
        RECT 2.525 130.195 2.695 130.365 ;
        RECT 3.485 130.195 3.655 130.365 ;
        RECT 4.445 130.195 4.615 130.365 ;
        RECT 5.405 130.195 5.575 130.365 ;
        RECT 6.365 130.195 6.535 130.365 ;
        RECT 1.565 123.760 1.735 123.930 ;
        RECT 2.525 123.760 2.695 123.930 ;
        RECT 3.485 123.760 3.655 123.930 ;
        RECT 4.445 123.760 4.615 123.930 ;
        RECT 5.405 123.760 5.575 123.930 ;
        RECT 6.365 123.760 6.535 123.930 ;
        RECT 1.565 117.325 1.735 117.495 ;
        RECT 2.525 117.325 2.695 117.495 ;
        RECT 3.485 117.325 3.655 117.495 ;
        RECT 4.445 117.325 4.615 117.495 ;
        RECT 5.405 117.325 5.575 117.495 ;
        RECT 6.365 117.325 6.535 117.495 ;
        RECT 1.565 110.890 1.735 111.060 ;
        RECT 2.525 110.890 2.695 111.060 ;
        RECT 3.485 110.890 3.655 111.060 ;
        RECT 4.445 110.890 4.615 111.060 ;
        RECT 5.405 110.890 5.575 111.060 ;
        RECT 6.365 110.890 6.535 111.060 ;
        RECT 1.565 104.455 1.735 104.625 ;
        RECT 2.525 104.455 2.695 104.625 ;
        RECT 3.485 104.455 3.655 104.625 ;
        RECT 4.445 104.455 4.615 104.625 ;
        RECT 5.405 104.455 5.575 104.625 ;
        RECT 6.365 104.455 6.535 104.625 ;
        RECT 1.565 98.020 1.735 98.190 ;
        RECT 2.525 98.020 2.695 98.190 ;
        RECT 3.485 98.020 3.655 98.190 ;
        RECT 4.445 98.020 4.615 98.190 ;
        RECT 5.405 98.020 5.575 98.190 ;
        RECT 6.365 98.020 6.535 98.190 ;
        RECT 1.565 91.585 1.735 91.755 ;
        RECT 2.525 91.585 2.695 91.755 ;
        RECT 3.485 91.585 3.655 91.755 ;
        RECT 4.445 91.585 4.615 91.755 ;
        RECT 5.405 91.585 5.575 91.755 ;
        RECT 6.365 91.585 6.535 91.755 ;
        RECT 1.565 85.150 1.735 85.320 ;
        RECT 2.525 85.150 2.695 85.320 ;
        RECT 3.485 85.150 3.655 85.320 ;
        RECT 4.445 85.150 4.615 85.320 ;
        RECT 5.405 85.150 5.575 85.320 ;
        RECT 6.365 85.150 6.535 85.320 ;
        RECT 1.565 78.715 1.735 78.885 ;
        RECT 2.525 78.715 2.695 78.885 ;
        RECT 3.485 78.715 3.655 78.885 ;
        RECT 4.445 78.715 4.615 78.885 ;
        RECT 5.405 78.715 5.575 78.885 ;
        RECT 6.365 78.715 6.535 78.885 ;
        RECT 1.565 72.280 1.735 72.450 ;
        RECT 2.525 72.280 2.695 72.450 ;
        RECT 3.485 72.280 3.655 72.450 ;
        RECT 4.445 72.280 4.615 72.450 ;
        RECT 5.405 72.280 5.575 72.450 ;
        RECT 6.365 72.280 6.535 72.450 ;
        RECT 1.565 65.845 1.735 66.015 ;
        RECT 2.525 65.845 2.695 66.015 ;
        RECT 3.485 65.845 3.655 66.015 ;
        RECT 4.445 65.845 4.615 66.015 ;
        RECT 5.405 65.845 5.575 66.015 ;
        RECT 6.365 65.845 6.535 66.015 ;
        RECT 1.565 59.410 1.735 59.580 ;
        RECT 2.525 59.410 2.695 59.580 ;
        RECT 3.485 59.410 3.655 59.580 ;
        RECT 4.445 59.410 4.615 59.580 ;
        RECT 5.405 59.410 5.575 59.580 ;
        RECT 6.365 59.410 6.535 59.580 ;
        RECT 1.565 52.975 1.735 53.145 ;
        RECT 2.525 52.975 2.695 53.145 ;
        RECT 3.485 52.975 3.655 53.145 ;
        RECT 4.445 52.975 4.615 53.145 ;
        RECT 5.405 52.975 5.575 53.145 ;
        RECT 6.365 52.975 6.535 53.145 ;
        RECT 1.565 46.540 1.735 46.710 ;
        RECT 2.525 46.540 2.695 46.710 ;
        RECT 3.485 46.540 3.655 46.710 ;
        RECT 4.445 46.540 4.615 46.710 ;
        RECT 5.405 46.540 5.575 46.710 ;
        RECT 6.365 46.540 6.535 46.710 ;
        RECT 1.565 40.105 1.735 40.275 ;
        RECT 2.525 40.105 2.695 40.275 ;
        RECT 3.485 40.105 3.655 40.275 ;
        RECT 4.445 40.105 4.615 40.275 ;
        RECT 5.405 40.105 5.575 40.275 ;
        RECT 6.365 40.105 6.535 40.275 ;
        RECT 1.565 33.670 1.735 33.840 ;
        RECT 2.525 33.670 2.695 33.840 ;
        RECT 3.485 33.670 3.655 33.840 ;
        RECT 4.445 33.670 4.615 33.840 ;
        RECT 5.405 33.670 5.575 33.840 ;
        RECT 6.365 33.670 6.535 33.840 ;
        RECT 1.565 27.235 1.735 27.405 ;
        RECT 2.525 27.235 2.695 27.405 ;
        RECT 3.485 27.235 3.655 27.405 ;
        RECT 4.445 27.235 4.615 27.405 ;
        RECT 5.405 27.235 5.575 27.405 ;
        RECT 6.365 27.235 6.535 27.405 ;
        RECT 1.565 20.800 1.735 20.970 ;
        RECT 2.525 20.800 2.695 20.970 ;
        RECT 3.485 20.800 3.655 20.970 ;
        RECT 4.445 20.800 4.615 20.970 ;
        RECT 5.405 20.800 5.575 20.970 ;
        RECT 6.365 20.800 6.535 20.970 ;
        RECT 1.565 14.365 1.735 14.535 ;
        RECT 2.525 14.365 2.695 14.535 ;
        RECT 3.485 14.365 3.655 14.535 ;
        RECT 4.445 14.365 4.615 14.535 ;
        RECT 5.405 14.365 5.575 14.535 ;
        RECT 6.365 14.365 6.535 14.535 ;
        RECT 1.565 7.930 1.735 8.100 ;
        RECT 2.525 7.930 2.695 8.100 ;
        RECT 3.485 7.930 3.655 8.100 ;
        RECT 4.445 7.930 4.615 8.100 ;
        RECT 5.405 7.930 5.575 8.100 ;
        RECT 6.365 7.930 6.535 8.100 ;
        RECT 1.565 1.495 1.735 1.665 ;
        RECT 2.525 1.495 2.695 1.665 ;
        RECT 3.485 1.495 3.655 1.665 ;
        RECT 4.445 1.495 4.615 1.665 ;
        RECT 5.405 1.495 5.575 1.665 ;
        RECT 6.365 1.495 6.535 1.665 ;
      LAYER met1 ;
        RECT 9.600 201.220 9.980 201.230 ;
        RECT 1.485 201.205 1.815 201.220 ;
        RECT 2.445 201.205 2.775 201.220 ;
        RECT 3.405 201.205 3.735 201.220 ;
        RECT 4.365 201.205 4.695 201.220 ;
        RECT 1.470 200.945 1.830 201.205 ;
        RECT 2.425 200.945 2.785 201.205 ;
        RECT 3.385 200.945 3.745 201.205 ;
        RECT 4.345 200.945 4.705 201.205 ;
        RECT 5.325 201.200 5.655 201.220 ;
        RECT 6.285 201.200 6.615 201.220 ;
        RECT 1.485 200.920 1.815 200.945 ;
        RECT 2.445 200.920 2.775 200.945 ;
        RECT 3.405 200.920 3.735 200.945 ;
        RECT 4.365 200.920 4.695 200.945 ;
        RECT 5.310 200.940 5.670 201.200 ;
        RECT 6.270 200.940 6.630 201.200 ;
        RECT 7.290 200.950 9.980 201.220 ;
        RECT 7.290 200.940 9.930 200.950 ;
        RECT 5.325 200.920 5.655 200.940 ;
        RECT 6.285 200.920 6.615 200.940 ;
        RECT 9.600 194.785 9.980 194.795 ;
        RECT 1.485 194.770 1.815 194.785 ;
        RECT 2.445 194.770 2.775 194.785 ;
        RECT 3.405 194.770 3.735 194.785 ;
        RECT 4.365 194.770 4.695 194.785 ;
        RECT 1.470 194.510 1.830 194.770 ;
        RECT 2.425 194.510 2.785 194.770 ;
        RECT 3.385 194.510 3.745 194.770 ;
        RECT 4.345 194.510 4.705 194.770 ;
        RECT 5.325 194.765 5.655 194.785 ;
        RECT 6.285 194.765 6.615 194.785 ;
        RECT 1.485 194.485 1.815 194.510 ;
        RECT 2.445 194.485 2.775 194.510 ;
        RECT 3.405 194.485 3.735 194.510 ;
        RECT 4.365 194.485 4.695 194.510 ;
        RECT 5.310 194.505 5.670 194.765 ;
        RECT 6.270 194.505 6.630 194.765 ;
        RECT 7.290 194.515 9.980 194.785 ;
        RECT 7.290 194.505 9.930 194.515 ;
        RECT 5.325 194.485 5.655 194.505 ;
        RECT 6.285 194.485 6.615 194.505 ;
        RECT 9.600 188.350 9.980 188.360 ;
        RECT 1.485 188.335 1.815 188.350 ;
        RECT 2.445 188.335 2.775 188.350 ;
        RECT 3.405 188.335 3.735 188.350 ;
        RECT 4.365 188.335 4.695 188.350 ;
        RECT 1.470 188.075 1.830 188.335 ;
        RECT 2.425 188.075 2.785 188.335 ;
        RECT 3.385 188.075 3.745 188.335 ;
        RECT 4.345 188.075 4.705 188.335 ;
        RECT 5.325 188.330 5.655 188.350 ;
        RECT 6.285 188.330 6.615 188.350 ;
        RECT 1.485 188.050 1.815 188.075 ;
        RECT 2.445 188.050 2.775 188.075 ;
        RECT 3.405 188.050 3.735 188.075 ;
        RECT 4.365 188.050 4.695 188.075 ;
        RECT 5.310 188.070 5.670 188.330 ;
        RECT 6.270 188.070 6.630 188.330 ;
        RECT 7.290 188.080 9.980 188.350 ;
        RECT 7.290 188.070 9.930 188.080 ;
        RECT 5.325 188.050 5.655 188.070 ;
        RECT 6.285 188.050 6.615 188.070 ;
        RECT 9.600 181.915 9.980 181.925 ;
        RECT 1.485 181.900 1.815 181.915 ;
        RECT 2.445 181.900 2.775 181.915 ;
        RECT 3.405 181.900 3.735 181.915 ;
        RECT 4.365 181.900 4.695 181.915 ;
        RECT 1.470 181.640 1.830 181.900 ;
        RECT 2.425 181.640 2.785 181.900 ;
        RECT 3.385 181.640 3.745 181.900 ;
        RECT 4.345 181.640 4.705 181.900 ;
        RECT 5.325 181.895 5.655 181.915 ;
        RECT 6.285 181.895 6.615 181.915 ;
        RECT 1.485 181.615 1.815 181.640 ;
        RECT 2.445 181.615 2.775 181.640 ;
        RECT 3.405 181.615 3.735 181.640 ;
        RECT 4.365 181.615 4.695 181.640 ;
        RECT 5.310 181.635 5.670 181.895 ;
        RECT 6.270 181.635 6.630 181.895 ;
        RECT 7.290 181.645 9.980 181.915 ;
        RECT 7.290 181.635 9.930 181.645 ;
        RECT 5.325 181.615 5.655 181.635 ;
        RECT 6.285 181.615 6.615 181.635 ;
        RECT 9.600 175.480 9.980 175.490 ;
        RECT 1.485 175.465 1.815 175.480 ;
        RECT 2.445 175.465 2.775 175.480 ;
        RECT 3.405 175.465 3.735 175.480 ;
        RECT 4.365 175.465 4.695 175.480 ;
        RECT 1.470 175.205 1.830 175.465 ;
        RECT 2.425 175.205 2.785 175.465 ;
        RECT 3.385 175.205 3.745 175.465 ;
        RECT 4.345 175.205 4.705 175.465 ;
        RECT 5.325 175.460 5.655 175.480 ;
        RECT 6.285 175.460 6.615 175.480 ;
        RECT 1.485 175.180 1.815 175.205 ;
        RECT 2.445 175.180 2.775 175.205 ;
        RECT 3.405 175.180 3.735 175.205 ;
        RECT 4.365 175.180 4.695 175.205 ;
        RECT 5.310 175.200 5.670 175.460 ;
        RECT 6.270 175.200 6.630 175.460 ;
        RECT 7.290 175.210 9.980 175.480 ;
        RECT 7.290 175.200 9.930 175.210 ;
        RECT 5.325 175.180 5.655 175.200 ;
        RECT 6.285 175.180 6.615 175.200 ;
        RECT 9.600 169.045 9.980 169.055 ;
        RECT 1.485 169.030 1.815 169.045 ;
        RECT 2.445 169.030 2.775 169.045 ;
        RECT 3.405 169.030 3.735 169.045 ;
        RECT 4.365 169.030 4.695 169.045 ;
        RECT 1.470 168.770 1.830 169.030 ;
        RECT 2.425 168.770 2.785 169.030 ;
        RECT 3.385 168.770 3.745 169.030 ;
        RECT 4.345 168.770 4.705 169.030 ;
        RECT 5.325 169.025 5.655 169.045 ;
        RECT 6.285 169.025 6.615 169.045 ;
        RECT 1.485 168.745 1.815 168.770 ;
        RECT 2.445 168.745 2.775 168.770 ;
        RECT 3.405 168.745 3.735 168.770 ;
        RECT 4.365 168.745 4.695 168.770 ;
        RECT 5.310 168.765 5.670 169.025 ;
        RECT 6.270 168.765 6.630 169.025 ;
        RECT 7.290 168.775 9.980 169.045 ;
        RECT 7.290 168.765 9.930 168.775 ;
        RECT 5.325 168.745 5.655 168.765 ;
        RECT 6.285 168.745 6.615 168.765 ;
        RECT 9.600 162.610 9.980 162.620 ;
        RECT 1.485 162.595 1.815 162.610 ;
        RECT 2.445 162.595 2.775 162.610 ;
        RECT 3.405 162.595 3.735 162.610 ;
        RECT 4.365 162.595 4.695 162.610 ;
        RECT 1.470 162.335 1.830 162.595 ;
        RECT 2.425 162.335 2.785 162.595 ;
        RECT 3.385 162.335 3.745 162.595 ;
        RECT 4.345 162.335 4.705 162.595 ;
        RECT 5.325 162.590 5.655 162.610 ;
        RECT 6.285 162.590 6.615 162.610 ;
        RECT 1.485 162.310 1.815 162.335 ;
        RECT 2.445 162.310 2.775 162.335 ;
        RECT 3.405 162.310 3.735 162.335 ;
        RECT 4.365 162.310 4.695 162.335 ;
        RECT 5.310 162.330 5.670 162.590 ;
        RECT 6.270 162.330 6.630 162.590 ;
        RECT 7.290 162.340 9.980 162.610 ;
        RECT 7.290 162.330 9.930 162.340 ;
        RECT 5.325 162.310 5.655 162.330 ;
        RECT 6.285 162.310 6.615 162.330 ;
        RECT 9.600 156.175 9.980 156.185 ;
        RECT 1.485 156.160 1.815 156.175 ;
        RECT 2.445 156.160 2.775 156.175 ;
        RECT 3.405 156.160 3.735 156.175 ;
        RECT 4.365 156.160 4.695 156.175 ;
        RECT 1.470 155.900 1.830 156.160 ;
        RECT 2.425 155.900 2.785 156.160 ;
        RECT 3.385 155.900 3.745 156.160 ;
        RECT 4.345 155.900 4.705 156.160 ;
        RECT 5.325 156.155 5.655 156.175 ;
        RECT 6.285 156.155 6.615 156.175 ;
        RECT 1.485 155.875 1.815 155.900 ;
        RECT 2.445 155.875 2.775 155.900 ;
        RECT 3.405 155.875 3.735 155.900 ;
        RECT 4.365 155.875 4.695 155.900 ;
        RECT 5.310 155.895 5.670 156.155 ;
        RECT 6.270 155.895 6.630 156.155 ;
        RECT 7.290 155.905 9.980 156.175 ;
        RECT 7.290 155.895 9.930 155.905 ;
        RECT 5.325 155.875 5.655 155.895 ;
        RECT 6.285 155.875 6.615 155.895 ;
        RECT 9.600 149.740 9.980 149.750 ;
        RECT 1.485 149.725 1.815 149.740 ;
        RECT 2.445 149.725 2.775 149.740 ;
        RECT 3.405 149.725 3.735 149.740 ;
        RECT 4.365 149.725 4.695 149.740 ;
        RECT 1.470 149.465 1.830 149.725 ;
        RECT 2.425 149.465 2.785 149.725 ;
        RECT 3.385 149.465 3.745 149.725 ;
        RECT 4.345 149.465 4.705 149.725 ;
        RECT 5.325 149.720 5.655 149.740 ;
        RECT 6.285 149.720 6.615 149.740 ;
        RECT 1.485 149.440 1.815 149.465 ;
        RECT 2.445 149.440 2.775 149.465 ;
        RECT 3.405 149.440 3.735 149.465 ;
        RECT 4.365 149.440 4.695 149.465 ;
        RECT 5.310 149.460 5.670 149.720 ;
        RECT 6.270 149.460 6.630 149.720 ;
        RECT 7.290 149.470 9.980 149.740 ;
        RECT 7.290 149.460 9.930 149.470 ;
        RECT 5.325 149.440 5.655 149.460 ;
        RECT 6.285 149.440 6.615 149.460 ;
        RECT 9.600 143.305 9.980 143.315 ;
        RECT 1.485 143.290 1.815 143.305 ;
        RECT 2.445 143.290 2.775 143.305 ;
        RECT 3.405 143.290 3.735 143.305 ;
        RECT 4.365 143.290 4.695 143.305 ;
        RECT 1.470 143.030 1.830 143.290 ;
        RECT 2.425 143.030 2.785 143.290 ;
        RECT 3.385 143.030 3.745 143.290 ;
        RECT 4.345 143.030 4.705 143.290 ;
        RECT 5.325 143.285 5.655 143.305 ;
        RECT 6.285 143.285 6.615 143.305 ;
        RECT 1.485 143.005 1.815 143.030 ;
        RECT 2.445 143.005 2.775 143.030 ;
        RECT 3.405 143.005 3.735 143.030 ;
        RECT 4.365 143.005 4.695 143.030 ;
        RECT 5.310 143.025 5.670 143.285 ;
        RECT 6.270 143.025 6.630 143.285 ;
        RECT 7.290 143.035 9.980 143.305 ;
        RECT 7.290 143.025 9.930 143.035 ;
        RECT 5.325 143.005 5.655 143.025 ;
        RECT 6.285 143.005 6.615 143.025 ;
        RECT 9.600 136.870 9.980 136.880 ;
        RECT 1.485 136.855 1.815 136.870 ;
        RECT 2.445 136.855 2.775 136.870 ;
        RECT 3.405 136.855 3.735 136.870 ;
        RECT 4.365 136.855 4.695 136.870 ;
        RECT 1.470 136.595 1.830 136.855 ;
        RECT 2.425 136.595 2.785 136.855 ;
        RECT 3.385 136.595 3.745 136.855 ;
        RECT 4.345 136.595 4.705 136.855 ;
        RECT 5.325 136.850 5.655 136.870 ;
        RECT 6.285 136.850 6.615 136.870 ;
        RECT 1.485 136.570 1.815 136.595 ;
        RECT 2.445 136.570 2.775 136.595 ;
        RECT 3.405 136.570 3.735 136.595 ;
        RECT 4.365 136.570 4.695 136.595 ;
        RECT 5.310 136.590 5.670 136.850 ;
        RECT 6.270 136.590 6.630 136.850 ;
        RECT 7.290 136.600 9.980 136.870 ;
        RECT 7.290 136.590 9.930 136.600 ;
        RECT 5.325 136.570 5.655 136.590 ;
        RECT 6.285 136.570 6.615 136.590 ;
        RECT 9.600 130.435 9.980 130.445 ;
        RECT 1.485 130.420 1.815 130.435 ;
        RECT 2.445 130.420 2.775 130.435 ;
        RECT 3.405 130.420 3.735 130.435 ;
        RECT 4.365 130.420 4.695 130.435 ;
        RECT 1.470 130.160 1.830 130.420 ;
        RECT 2.425 130.160 2.785 130.420 ;
        RECT 3.385 130.160 3.745 130.420 ;
        RECT 4.345 130.160 4.705 130.420 ;
        RECT 5.325 130.415 5.655 130.435 ;
        RECT 6.285 130.415 6.615 130.435 ;
        RECT 1.485 130.135 1.815 130.160 ;
        RECT 2.445 130.135 2.775 130.160 ;
        RECT 3.405 130.135 3.735 130.160 ;
        RECT 4.365 130.135 4.695 130.160 ;
        RECT 5.310 130.155 5.670 130.415 ;
        RECT 6.270 130.155 6.630 130.415 ;
        RECT 7.290 130.165 9.980 130.435 ;
        RECT 7.290 130.155 9.930 130.165 ;
        RECT 5.325 130.135 5.655 130.155 ;
        RECT 6.285 130.135 6.615 130.155 ;
        RECT 9.600 124.000 9.980 124.010 ;
        RECT 1.485 123.985 1.815 124.000 ;
        RECT 2.445 123.985 2.775 124.000 ;
        RECT 3.405 123.985 3.735 124.000 ;
        RECT 4.365 123.985 4.695 124.000 ;
        RECT 1.470 123.725 1.830 123.985 ;
        RECT 2.425 123.725 2.785 123.985 ;
        RECT 3.385 123.725 3.745 123.985 ;
        RECT 4.345 123.725 4.705 123.985 ;
        RECT 5.325 123.980 5.655 124.000 ;
        RECT 6.285 123.980 6.615 124.000 ;
        RECT 1.485 123.700 1.815 123.725 ;
        RECT 2.445 123.700 2.775 123.725 ;
        RECT 3.405 123.700 3.735 123.725 ;
        RECT 4.365 123.700 4.695 123.725 ;
        RECT 5.310 123.720 5.670 123.980 ;
        RECT 6.270 123.720 6.630 123.980 ;
        RECT 7.290 123.730 9.980 124.000 ;
        RECT 7.290 123.720 9.930 123.730 ;
        RECT 5.325 123.700 5.655 123.720 ;
        RECT 6.285 123.700 6.615 123.720 ;
        RECT 9.600 117.565 9.980 117.575 ;
        RECT 1.485 117.550 1.815 117.565 ;
        RECT 2.445 117.550 2.775 117.565 ;
        RECT 3.405 117.550 3.735 117.565 ;
        RECT 4.365 117.550 4.695 117.565 ;
        RECT 1.470 117.290 1.830 117.550 ;
        RECT 2.425 117.290 2.785 117.550 ;
        RECT 3.385 117.290 3.745 117.550 ;
        RECT 4.345 117.290 4.705 117.550 ;
        RECT 5.325 117.545 5.655 117.565 ;
        RECT 6.285 117.545 6.615 117.565 ;
        RECT 1.485 117.265 1.815 117.290 ;
        RECT 2.445 117.265 2.775 117.290 ;
        RECT 3.405 117.265 3.735 117.290 ;
        RECT 4.365 117.265 4.695 117.290 ;
        RECT 5.310 117.285 5.670 117.545 ;
        RECT 6.270 117.285 6.630 117.545 ;
        RECT 7.290 117.295 9.980 117.565 ;
        RECT 7.290 117.285 9.930 117.295 ;
        RECT 5.325 117.265 5.655 117.285 ;
        RECT 6.285 117.265 6.615 117.285 ;
        RECT 9.600 111.130 9.980 111.140 ;
        RECT 1.485 111.115 1.815 111.130 ;
        RECT 2.445 111.115 2.775 111.130 ;
        RECT 3.405 111.115 3.735 111.130 ;
        RECT 4.365 111.115 4.695 111.130 ;
        RECT 1.470 110.855 1.830 111.115 ;
        RECT 2.425 110.855 2.785 111.115 ;
        RECT 3.385 110.855 3.745 111.115 ;
        RECT 4.345 110.855 4.705 111.115 ;
        RECT 5.325 111.110 5.655 111.130 ;
        RECT 6.285 111.110 6.615 111.130 ;
        RECT 1.485 110.830 1.815 110.855 ;
        RECT 2.445 110.830 2.775 110.855 ;
        RECT 3.405 110.830 3.735 110.855 ;
        RECT 4.365 110.830 4.695 110.855 ;
        RECT 5.310 110.850 5.670 111.110 ;
        RECT 6.270 110.850 6.630 111.110 ;
        RECT 7.290 110.860 9.980 111.130 ;
        RECT 7.290 110.850 9.930 110.860 ;
        RECT 5.325 110.830 5.655 110.850 ;
        RECT 6.285 110.830 6.615 110.850 ;
        RECT 9.600 104.695 9.980 104.705 ;
        RECT 1.485 104.680 1.815 104.695 ;
        RECT 2.445 104.680 2.775 104.695 ;
        RECT 3.405 104.680 3.735 104.695 ;
        RECT 4.365 104.680 4.695 104.695 ;
        RECT 1.470 104.420 1.830 104.680 ;
        RECT 2.425 104.420 2.785 104.680 ;
        RECT 3.385 104.420 3.745 104.680 ;
        RECT 4.345 104.420 4.705 104.680 ;
        RECT 5.325 104.675 5.655 104.695 ;
        RECT 6.285 104.675 6.615 104.695 ;
        RECT 1.485 104.395 1.815 104.420 ;
        RECT 2.445 104.395 2.775 104.420 ;
        RECT 3.405 104.395 3.735 104.420 ;
        RECT 4.365 104.395 4.695 104.420 ;
        RECT 5.310 104.415 5.670 104.675 ;
        RECT 6.270 104.415 6.630 104.675 ;
        RECT 7.290 104.425 9.980 104.695 ;
        RECT 7.290 104.415 9.930 104.425 ;
        RECT 5.325 104.395 5.655 104.415 ;
        RECT 6.285 104.395 6.615 104.415 ;
        RECT 9.600 98.260 9.980 98.270 ;
        RECT 1.485 98.245 1.815 98.260 ;
        RECT 2.445 98.245 2.775 98.260 ;
        RECT 3.405 98.245 3.735 98.260 ;
        RECT 4.365 98.245 4.695 98.260 ;
        RECT 1.470 97.985 1.830 98.245 ;
        RECT 2.425 97.985 2.785 98.245 ;
        RECT 3.385 97.985 3.745 98.245 ;
        RECT 4.345 97.985 4.705 98.245 ;
        RECT 5.325 98.240 5.655 98.260 ;
        RECT 6.285 98.240 6.615 98.260 ;
        RECT 1.485 97.960 1.815 97.985 ;
        RECT 2.445 97.960 2.775 97.985 ;
        RECT 3.405 97.960 3.735 97.985 ;
        RECT 4.365 97.960 4.695 97.985 ;
        RECT 5.310 97.980 5.670 98.240 ;
        RECT 6.270 97.980 6.630 98.240 ;
        RECT 7.290 97.990 9.980 98.260 ;
        RECT 7.290 97.980 9.930 97.990 ;
        RECT 5.325 97.960 5.655 97.980 ;
        RECT 6.285 97.960 6.615 97.980 ;
        RECT 9.600 91.825 9.980 91.835 ;
        RECT 1.485 91.810 1.815 91.825 ;
        RECT 2.445 91.810 2.775 91.825 ;
        RECT 3.405 91.810 3.735 91.825 ;
        RECT 4.365 91.810 4.695 91.825 ;
        RECT 1.470 91.550 1.830 91.810 ;
        RECT 2.425 91.550 2.785 91.810 ;
        RECT 3.385 91.550 3.745 91.810 ;
        RECT 4.345 91.550 4.705 91.810 ;
        RECT 5.325 91.805 5.655 91.825 ;
        RECT 6.285 91.805 6.615 91.825 ;
        RECT 1.485 91.525 1.815 91.550 ;
        RECT 2.445 91.525 2.775 91.550 ;
        RECT 3.405 91.525 3.735 91.550 ;
        RECT 4.365 91.525 4.695 91.550 ;
        RECT 5.310 91.545 5.670 91.805 ;
        RECT 6.270 91.545 6.630 91.805 ;
        RECT 7.290 91.555 9.980 91.825 ;
        RECT 7.290 91.545 9.930 91.555 ;
        RECT 5.325 91.525 5.655 91.545 ;
        RECT 6.285 91.525 6.615 91.545 ;
        RECT 9.600 85.390 9.980 85.400 ;
        RECT 1.485 85.375 1.815 85.390 ;
        RECT 2.445 85.375 2.775 85.390 ;
        RECT 3.405 85.375 3.735 85.390 ;
        RECT 4.365 85.375 4.695 85.390 ;
        RECT 1.470 85.115 1.830 85.375 ;
        RECT 2.425 85.115 2.785 85.375 ;
        RECT 3.385 85.115 3.745 85.375 ;
        RECT 4.345 85.115 4.705 85.375 ;
        RECT 5.325 85.370 5.655 85.390 ;
        RECT 6.285 85.370 6.615 85.390 ;
        RECT 1.485 85.090 1.815 85.115 ;
        RECT 2.445 85.090 2.775 85.115 ;
        RECT 3.405 85.090 3.735 85.115 ;
        RECT 4.365 85.090 4.695 85.115 ;
        RECT 5.310 85.110 5.670 85.370 ;
        RECT 6.270 85.110 6.630 85.370 ;
        RECT 7.290 85.120 9.980 85.390 ;
        RECT 7.290 85.110 9.930 85.120 ;
        RECT 5.325 85.090 5.655 85.110 ;
        RECT 6.285 85.090 6.615 85.110 ;
        RECT 9.600 78.955 9.980 78.965 ;
        RECT 1.485 78.940 1.815 78.955 ;
        RECT 2.445 78.940 2.775 78.955 ;
        RECT 3.405 78.940 3.735 78.955 ;
        RECT 4.365 78.940 4.695 78.955 ;
        RECT 1.470 78.680 1.830 78.940 ;
        RECT 2.425 78.680 2.785 78.940 ;
        RECT 3.385 78.680 3.745 78.940 ;
        RECT 4.345 78.680 4.705 78.940 ;
        RECT 5.325 78.935 5.655 78.955 ;
        RECT 6.285 78.935 6.615 78.955 ;
        RECT 1.485 78.655 1.815 78.680 ;
        RECT 2.445 78.655 2.775 78.680 ;
        RECT 3.405 78.655 3.735 78.680 ;
        RECT 4.365 78.655 4.695 78.680 ;
        RECT 5.310 78.675 5.670 78.935 ;
        RECT 6.270 78.675 6.630 78.935 ;
        RECT 7.290 78.685 9.980 78.955 ;
        RECT 7.290 78.675 9.930 78.685 ;
        RECT 5.325 78.655 5.655 78.675 ;
        RECT 6.285 78.655 6.615 78.675 ;
        RECT 9.600 72.520 9.980 72.530 ;
        RECT 1.485 72.505 1.815 72.520 ;
        RECT 2.445 72.505 2.775 72.520 ;
        RECT 3.405 72.505 3.735 72.520 ;
        RECT 4.365 72.505 4.695 72.520 ;
        RECT 1.470 72.245 1.830 72.505 ;
        RECT 2.425 72.245 2.785 72.505 ;
        RECT 3.385 72.245 3.745 72.505 ;
        RECT 4.345 72.245 4.705 72.505 ;
        RECT 5.325 72.500 5.655 72.520 ;
        RECT 6.285 72.500 6.615 72.520 ;
        RECT 1.485 72.220 1.815 72.245 ;
        RECT 2.445 72.220 2.775 72.245 ;
        RECT 3.405 72.220 3.735 72.245 ;
        RECT 4.365 72.220 4.695 72.245 ;
        RECT 5.310 72.240 5.670 72.500 ;
        RECT 6.270 72.240 6.630 72.500 ;
        RECT 7.290 72.250 9.980 72.520 ;
        RECT 7.290 72.240 9.930 72.250 ;
        RECT 5.325 72.220 5.655 72.240 ;
        RECT 6.285 72.220 6.615 72.240 ;
        RECT 9.600 66.085 9.980 66.095 ;
        RECT 1.485 66.070 1.815 66.085 ;
        RECT 2.445 66.070 2.775 66.085 ;
        RECT 3.405 66.070 3.735 66.085 ;
        RECT 4.365 66.070 4.695 66.085 ;
        RECT 1.470 65.810 1.830 66.070 ;
        RECT 2.425 65.810 2.785 66.070 ;
        RECT 3.385 65.810 3.745 66.070 ;
        RECT 4.345 65.810 4.705 66.070 ;
        RECT 5.325 66.065 5.655 66.085 ;
        RECT 6.285 66.065 6.615 66.085 ;
        RECT 1.485 65.785 1.815 65.810 ;
        RECT 2.445 65.785 2.775 65.810 ;
        RECT 3.405 65.785 3.735 65.810 ;
        RECT 4.365 65.785 4.695 65.810 ;
        RECT 5.310 65.805 5.670 66.065 ;
        RECT 6.270 65.805 6.630 66.065 ;
        RECT 7.290 65.815 9.980 66.085 ;
        RECT 7.290 65.805 9.930 65.815 ;
        RECT 5.325 65.785 5.655 65.805 ;
        RECT 6.285 65.785 6.615 65.805 ;
        RECT 9.600 59.650 9.980 59.660 ;
        RECT 1.485 59.635 1.815 59.650 ;
        RECT 2.445 59.635 2.775 59.650 ;
        RECT 3.405 59.635 3.735 59.650 ;
        RECT 4.365 59.635 4.695 59.650 ;
        RECT 1.470 59.375 1.830 59.635 ;
        RECT 2.425 59.375 2.785 59.635 ;
        RECT 3.385 59.375 3.745 59.635 ;
        RECT 4.345 59.375 4.705 59.635 ;
        RECT 5.325 59.630 5.655 59.650 ;
        RECT 6.285 59.630 6.615 59.650 ;
        RECT 1.485 59.350 1.815 59.375 ;
        RECT 2.445 59.350 2.775 59.375 ;
        RECT 3.405 59.350 3.735 59.375 ;
        RECT 4.365 59.350 4.695 59.375 ;
        RECT 5.310 59.370 5.670 59.630 ;
        RECT 6.270 59.370 6.630 59.630 ;
        RECT 7.290 59.380 9.980 59.650 ;
        RECT 7.290 59.370 9.930 59.380 ;
        RECT 5.325 59.350 5.655 59.370 ;
        RECT 6.285 59.350 6.615 59.370 ;
        RECT 9.600 53.215 9.980 53.225 ;
        RECT 1.485 53.200 1.815 53.215 ;
        RECT 2.445 53.200 2.775 53.215 ;
        RECT 3.405 53.200 3.735 53.215 ;
        RECT 4.365 53.200 4.695 53.215 ;
        RECT 1.470 52.940 1.830 53.200 ;
        RECT 2.425 52.940 2.785 53.200 ;
        RECT 3.385 52.940 3.745 53.200 ;
        RECT 4.345 52.940 4.705 53.200 ;
        RECT 5.325 53.195 5.655 53.215 ;
        RECT 6.285 53.195 6.615 53.215 ;
        RECT 1.485 52.915 1.815 52.940 ;
        RECT 2.445 52.915 2.775 52.940 ;
        RECT 3.405 52.915 3.735 52.940 ;
        RECT 4.365 52.915 4.695 52.940 ;
        RECT 5.310 52.935 5.670 53.195 ;
        RECT 6.270 52.935 6.630 53.195 ;
        RECT 7.290 52.945 9.980 53.215 ;
        RECT 7.290 52.935 9.930 52.945 ;
        RECT 5.325 52.915 5.655 52.935 ;
        RECT 6.285 52.915 6.615 52.935 ;
        RECT 9.600 46.780 9.980 46.790 ;
        RECT 1.485 46.765 1.815 46.780 ;
        RECT 2.445 46.765 2.775 46.780 ;
        RECT 3.405 46.765 3.735 46.780 ;
        RECT 4.365 46.765 4.695 46.780 ;
        RECT 1.470 46.505 1.830 46.765 ;
        RECT 2.425 46.505 2.785 46.765 ;
        RECT 3.385 46.505 3.745 46.765 ;
        RECT 4.345 46.505 4.705 46.765 ;
        RECT 5.325 46.760 5.655 46.780 ;
        RECT 6.285 46.760 6.615 46.780 ;
        RECT 1.485 46.480 1.815 46.505 ;
        RECT 2.445 46.480 2.775 46.505 ;
        RECT 3.405 46.480 3.735 46.505 ;
        RECT 4.365 46.480 4.695 46.505 ;
        RECT 5.310 46.500 5.670 46.760 ;
        RECT 6.270 46.500 6.630 46.760 ;
        RECT 7.290 46.510 9.980 46.780 ;
        RECT 7.290 46.500 9.930 46.510 ;
        RECT 5.325 46.480 5.655 46.500 ;
        RECT 6.285 46.480 6.615 46.500 ;
        RECT 9.600 40.345 9.980 40.355 ;
        RECT 1.485 40.330 1.815 40.345 ;
        RECT 2.445 40.330 2.775 40.345 ;
        RECT 3.405 40.330 3.735 40.345 ;
        RECT 4.365 40.330 4.695 40.345 ;
        RECT 1.470 40.070 1.830 40.330 ;
        RECT 2.425 40.070 2.785 40.330 ;
        RECT 3.385 40.070 3.745 40.330 ;
        RECT 4.345 40.070 4.705 40.330 ;
        RECT 5.325 40.325 5.655 40.345 ;
        RECT 6.285 40.325 6.615 40.345 ;
        RECT 1.485 40.045 1.815 40.070 ;
        RECT 2.445 40.045 2.775 40.070 ;
        RECT 3.405 40.045 3.735 40.070 ;
        RECT 4.365 40.045 4.695 40.070 ;
        RECT 5.310 40.065 5.670 40.325 ;
        RECT 6.270 40.065 6.630 40.325 ;
        RECT 7.290 40.075 9.980 40.345 ;
        RECT 7.290 40.065 9.930 40.075 ;
        RECT 5.325 40.045 5.655 40.065 ;
        RECT 6.285 40.045 6.615 40.065 ;
        RECT 9.600 33.910 9.980 33.920 ;
        RECT 1.485 33.895 1.815 33.910 ;
        RECT 2.445 33.895 2.775 33.910 ;
        RECT 3.405 33.895 3.735 33.910 ;
        RECT 4.365 33.895 4.695 33.910 ;
        RECT 1.470 33.635 1.830 33.895 ;
        RECT 2.425 33.635 2.785 33.895 ;
        RECT 3.385 33.635 3.745 33.895 ;
        RECT 4.345 33.635 4.705 33.895 ;
        RECT 5.325 33.890 5.655 33.910 ;
        RECT 6.285 33.890 6.615 33.910 ;
        RECT 1.485 33.610 1.815 33.635 ;
        RECT 2.445 33.610 2.775 33.635 ;
        RECT 3.405 33.610 3.735 33.635 ;
        RECT 4.365 33.610 4.695 33.635 ;
        RECT 5.310 33.630 5.670 33.890 ;
        RECT 6.270 33.630 6.630 33.890 ;
        RECT 7.290 33.640 9.980 33.910 ;
        RECT 7.290 33.630 9.930 33.640 ;
        RECT 5.325 33.610 5.655 33.630 ;
        RECT 6.285 33.610 6.615 33.630 ;
        RECT 9.600 27.475 9.980 27.485 ;
        RECT 1.485 27.460 1.815 27.475 ;
        RECT 2.445 27.460 2.775 27.475 ;
        RECT 3.405 27.460 3.735 27.475 ;
        RECT 4.365 27.460 4.695 27.475 ;
        RECT 1.470 27.200 1.830 27.460 ;
        RECT 2.425 27.200 2.785 27.460 ;
        RECT 3.385 27.200 3.745 27.460 ;
        RECT 4.345 27.200 4.705 27.460 ;
        RECT 5.325 27.455 5.655 27.475 ;
        RECT 6.285 27.455 6.615 27.475 ;
        RECT 1.485 27.175 1.815 27.200 ;
        RECT 2.445 27.175 2.775 27.200 ;
        RECT 3.405 27.175 3.735 27.200 ;
        RECT 4.365 27.175 4.695 27.200 ;
        RECT 5.310 27.195 5.670 27.455 ;
        RECT 6.270 27.195 6.630 27.455 ;
        RECT 7.290 27.205 9.980 27.475 ;
        RECT 7.290 27.195 9.930 27.205 ;
        RECT 5.325 27.175 5.655 27.195 ;
        RECT 6.285 27.175 6.615 27.195 ;
        RECT 9.600 21.040 9.980 21.050 ;
        RECT 1.485 21.025 1.815 21.040 ;
        RECT 2.445 21.025 2.775 21.040 ;
        RECT 3.405 21.025 3.735 21.040 ;
        RECT 4.365 21.025 4.695 21.040 ;
        RECT 1.470 20.765 1.830 21.025 ;
        RECT 2.425 20.765 2.785 21.025 ;
        RECT 3.385 20.765 3.745 21.025 ;
        RECT 4.345 20.765 4.705 21.025 ;
        RECT 5.325 21.020 5.655 21.040 ;
        RECT 6.285 21.020 6.615 21.040 ;
        RECT 1.485 20.740 1.815 20.765 ;
        RECT 2.445 20.740 2.775 20.765 ;
        RECT 3.405 20.740 3.735 20.765 ;
        RECT 4.365 20.740 4.695 20.765 ;
        RECT 5.310 20.760 5.670 21.020 ;
        RECT 6.270 20.760 6.630 21.020 ;
        RECT 7.290 20.770 9.980 21.040 ;
        RECT 7.290 20.760 9.930 20.770 ;
        RECT 5.325 20.740 5.655 20.760 ;
        RECT 6.285 20.740 6.615 20.760 ;
        RECT 9.600 14.605 9.980 14.615 ;
        RECT 1.485 14.590 1.815 14.605 ;
        RECT 2.445 14.590 2.775 14.605 ;
        RECT 3.405 14.590 3.735 14.605 ;
        RECT 4.365 14.590 4.695 14.605 ;
        RECT 1.470 14.330 1.830 14.590 ;
        RECT 2.425 14.330 2.785 14.590 ;
        RECT 3.385 14.330 3.745 14.590 ;
        RECT 4.345 14.330 4.705 14.590 ;
        RECT 5.325 14.585 5.655 14.605 ;
        RECT 6.285 14.585 6.615 14.605 ;
        RECT 1.485 14.305 1.815 14.330 ;
        RECT 2.445 14.305 2.775 14.330 ;
        RECT 3.405 14.305 3.735 14.330 ;
        RECT 4.365 14.305 4.695 14.330 ;
        RECT 5.310 14.325 5.670 14.585 ;
        RECT 6.270 14.325 6.630 14.585 ;
        RECT 7.290 14.335 9.980 14.605 ;
        RECT 7.290 14.325 9.930 14.335 ;
        RECT 5.325 14.305 5.655 14.325 ;
        RECT 6.285 14.305 6.615 14.325 ;
        RECT 9.600 8.170 9.980 8.180 ;
        RECT 1.485 8.155 1.815 8.170 ;
        RECT 2.445 8.155 2.775 8.170 ;
        RECT 3.405 8.155 3.735 8.170 ;
        RECT 4.365 8.155 4.695 8.170 ;
        RECT 1.470 7.895 1.830 8.155 ;
        RECT 2.425 7.895 2.785 8.155 ;
        RECT 3.385 7.895 3.745 8.155 ;
        RECT 4.345 7.895 4.705 8.155 ;
        RECT 5.325 8.150 5.655 8.170 ;
        RECT 6.285 8.150 6.615 8.170 ;
        RECT 1.485 7.870 1.815 7.895 ;
        RECT 2.445 7.870 2.775 7.895 ;
        RECT 3.405 7.870 3.735 7.895 ;
        RECT 4.365 7.870 4.695 7.895 ;
        RECT 5.310 7.890 5.670 8.150 ;
        RECT 6.270 7.890 6.630 8.150 ;
        RECT 7.290 7.900 9.980 8.170 ;
        RECT 7.290 7.890 9.930 7.900 ;
        RECT 5.325 7.870 5.655 7.890 ;
        RECT 6.285 7.870 6.615 7.890 ;
        RECT 9.600 1.735 9.980 1.745 ;
        RECT 1.485 1.720 1.815 1.735 ;
        RECT 2.445 1.720 2.775 1.735 ;
        RECT 3.405 1.720 3.735 1.735 ;
        RECT 4.365 1.720 4.695 1.735 ;
        RECT 1.470 1.460 1.830 1.720 ;
        RECT 2.425 1.460 2.785 1.720 ;
        RECT 3.385 1.460 3.745 1.720 ;
        RECT 4.345 1.460 4.705 1.720 ;
        RECT 5.325 1.715 5.655 1.735 ;
        RECT 6.285 1.715 6.615 1.735 ;
        RECT 1.485 1.435 1.815 1.460 ;
        RECT 2.445 1.435 2.775 1.460 ;
        RECT 3.405 1.435 3.735 1.460 ;
        RECT 4.365 1.435 4.695 1.460 ;
        RECT 5.310 1.455 5.670 1.715 ;
        RECT 6.270 1.455 6.630 1.715 ;
        RECT 7.290 1.465 9.980 1.735 ;
        RECT 7.290 1.455 9.930 1.465 ;
        RECT 5.325 1.435 5.655 1.455 ;
        RECT 6.285 1.435 6.615 1.455 ;
      LAYER via ;
        RECT 1.520 200.945 1.780 201.205 ;
        RECT 2.475 200.945 2.735 201.205 ;
        RECT 3.435 200.945 3.695 201.205 ;
        RECT 4.395 200.945 4.655 201.205 ;
        RECT 5.360 200.940 5.620 201.200 ;
        RECT 6.320 200.940 6.580 201.200 ;
        RECT 7.340 200.940 7.620 201.220 ;
        RECT 9.650 200.950 9.930 201.230 ;
        RECT 1.520 194.510 1.780 194.770 ;
        RECT 2.475 194.510 2.735 194.770 ;
        RECT 3.435 194.510 3.695 194.770 ;
        RECT 4.395 194.510 4.655 194.770 ;
        RECT 5.360 194.505 5.620 194.765 ;
        RECT 6.320 194.505 6.580 194.765 ;
        RECT 7.340 194.505 7.620 194.785 ;
        RECT 9.650 194.515 9.930 194.795 ;
        RECT 1.520 188.075 1.780 188.335 ;
        RECT 2.475 188.075 2.735 188.335 ;
        RECT 3.435 188.075 3.695 188.335 ;
        RECT 4.395 188.075 4.655 188.335 ;
        RECT 5.360 188.070 5.620 188.330 ;
        RECT 6.320 188.070 6.580 188.330 ;
        RECT 7.340 188.070 7.620 188.350 ;
        RECT 9.650 188.080 9.930 188.360 ;
        RECT 1.520 181.640 1.780 181.900 ;
        RECT 2.475 181.640 2.735 181.900 ;
        RECT 3.435 181.640 3.695 181.900 ;
        RECT 4.395 181.640 4.655 181.900 ;
        RECT 5.360 181.635 5.620 181.895 ;
        RECT 6.320 181.635 6.580 181.895 ;
        RECT 7.340 181.635 7.620 181.915 ;
        RECT 9.650 181.645 9.930 181.925 ;
        RECT 1.520 175.205 1.780 175.465 ;
        RECT 2.475 175.205 2.735 175.465 ;
        RECT 3.435 175.205 3.695 175.465 ;
        RECT 4.395 175.205 4.655 175.465 ;
        RECT 5.360 175.200 5.620 175.460 ;
        RECT 6.320 175.200 6.580 175.460 ;
        RECT 7.340 175.200 7.620 175.480 ;
        RECT 9.650 175.210 9.930 175.490 ;
        RECT 1.520 168.770 1.780 169.030 ;
        RECT 2.475 168.770 2.735 169.030 ;
        RECT 3.435 168.770 3.695 169.030 ;
        RECT 4.395 168.770 4.655 169.030 ;
        RECT 5.360 168.765 5.620 169.025 ;
        RECT 6.320 168.765 6.580 169.025 ;
        RECT 7.340 168.765 7.620 169.045 ;
        RECT 9.650 168.775 9.930 169.055 ;
        RECT 1.520 162.335 1.780 162.595 ;
        RECT 2.475 162.335 2.735 162.595 ;
        RECT 3.435 162.335 3.695 162.595 ;
        RECT 4.395 162.335 4.655 162.595 ;
        RECT 5.360 162.330 5.620 162.590 ;
        RECT 6.320 162.330 6.580 162.590 ;
        RECT 7.340 162.330 7.620 162.610 ;
        RECT 9.650 162.340 9.930 162.620 ;
        RECT 1.520 155.900 1.780 156.160 ;
        RECT 2.475 155.900 2.735 156.160 ;
        RECT 3.435 155.900 3.695 156.160 ;
        RECT 4.395 155.900 4.655 156.160 ;
        RECT 5.360 155.895 5.620 156.155 ;
        RECT 6.320 155.895 6.580 156.155 ;
        RECT 7.340 155.895 7.620 156.175 ;
        RECT 9.650 155.905 9.930 156.185 ;
        RECT 1.520 149.465 1.780 149.725 ;
        RECT 2.475 149.465 2.735 149.725 ;
        RECT 3.435 149.465 3.695 149.725 ;
        RECT 4.395 149.465 4.655 149.725 ;
        RECT 5.360 149.460 5.620 149.720 ;
        RECT 6.320 149.460 6.580 149.720 ;
        RECT 7.340 149.460 7.620 149.740 ;
        RECT 9.650 149.470 9.930 149.750 ;
        RECT 1.520 143.030 1.780 143.290 ;
        RECT 2.475 143.030 2.735 143.290 ;
        RECT 3.435 143.030 3.695 143.290 ;
        RECT 4.395 143.030 4.655 143.290 ;
        RECT 5.360 143.025 5.620 143.285 ;
        RECT 6.320 143.025 6.580 143.285 ;
        RECT 7.340 143.025 7.620 143.305 ;
        RECT 9.650 143.035 9.930 143.315 ;
        RECT 1.520 136.595 1.780 136.855 ;
        RECT 2.475 136.595 2.735 136.855 ;
        RECT 3.435 136.595 3.695 136.855 ;
        RECT 4.395 136.595 4.655 136.855 ;
        RECT 5.360 136.590 5.620 136.850 ;
        RECT 6.320 136.590 6.580 136.850 ;
        RECT 7.340 136.590 7.620 136.870 ;
        RECT 9.650 136.600 9.930 136.880 ;
        RECT 1.520 130.160 1.780 130.420 ;
        RECT 2.475 130.160 2.735 130.420 ;
        RECT 3.435 130.160 3.695 130.420 ;
        RECT 4.395 130.160 4.655 130.420 ;
        RECT 5.360 130.155 5.620 130.415 ;
        RECT 6.320 130.155 6.580 130.415 ;
        RECT 7.340 130.155 7.620 130.435 ;
        RECT 9.650 130.165 9.930 130.445 ;
        RECT 1.520 123.725 1.780 123.985 ;
        RECT 2.475 123.725 2.735 123.985 ;
        RECT 3.435 123.725 3.695 123.985 ;
        RECT 4.395 123.725 4.655 123.985 ;
        RECT 5.360 123.720 5.620 123.980 ;
        RECT 6.320 123.720 6.580 123.980 ;
        RECT 7.340 123.720 7.620 124.000 ;
        RECT 9.650 123.730 9.930 124.010 ;
        RECT 1.520 117.290 1.780 117.550 ;
        RECT 2.475 117.290 2.735 117.550 ;
        RECT 3.435 117.290 3.695 117.550 ;
        RECT 4.395 117.290 4.655 117.550 ;
        RECT 5.360 117.285 5.620 117.545 ;
        RECT 6.320 117.285 6.580 117.545 ;
        RECT 7.340 117.285 7.620 117.565 ;
        RECT 9.650 117.295 9.930 117.575 ;
        RECT 1.520 110.855 1.780 111.115 ;
        RECT 2.475 110.855 2.735 111.115 ;
        RECT 3.435 110.855 3.695 111.115 ;
        RECT 4.395 110.855 4.655 111.115 ;
        RECT 5.360 110.850 5.620 111.110 ;
        RECT 6.320 110.850 6.580 111.110 ;
        RECT 7.340 110.850 7.620 111.130 ;
        RECT 9.650 110.860 9.930 111.140 ;
        RECT 1.520 104.420 1.780 104.680 ;
        RECT 2.475 104.420 2.735 104.680 ;
        RECT 3.435 104.420 3.695 104.680 ;
        RECT 4.395 104.420 4.655 104.680 ;
        RECT 5.360 104.415 5.620 104.675 ;
        RECT 6.320 104.415 6.580 104.675 ;
        RECT 7.340 104.415 7.620 104.695 ;
        RECT 9.650 104.425 9.930 104.705 ;
        RECT 1.520 97.985 1.780 98.245 ;
        RECT 2.475 97.985 2.735 98.245 ;
        RECT 3.435 97.985 3.695 98.245 ;
        RECT 4.395 97.985 4.655 98.245 ;
        RECT 5.360 97.980 5.620 98.240 ;
        RECT 6.320 97.980 6.580 98.240 ;
        RECT 7.340 97.980 7.620 98.260 ;
        RECT 9.650 97.990 9.930 98.270 ;
        RECT 1.520 91.550 1.780 91.810 ;
        RECT 2.475 91.550 2.735 91.810 ;
        RECT 3.435 91.550 3.695 91.810 ;
        RECT 4.395 91.550 4.655 91.810 ;
        RECT 5.360 91.545 5.620 91.805 ;
        RECT 6.320 91.545 6.580 91.805 ;
        RECT 7.340 91.545 7.620 91.825 ;
        RECT 9.650 91.555 9.930 91.835 ;
        RECT 1.520 85.115 1.780 85.375 ;
        RECT 2.475 85.115 2.735 85.375 ;
        RECT 3.435 85.115 3.695 85.375 ;
        RECT 4.395 85.115 4.655 85.375 ;
        RECT 5.360 85.110 5.620 85.370 ;
        RECT 6.320 85.110 6.580 85.370 ;
        RECT 7.340 85.110 7.620 85.390 ;
        RECT 9.650 85.120 9.930 85.400 ;
        RECT 1.520 78.680 1.780 78.940 ;
        RECT 2.475 78.680 2.735 78.940 ;
        RECT 3.435 78.680 3.695 78.940 ;
        RECT 4.395 78.680 4.655 78.940 ;
        RECT 5.360 78.675 5.620 78.935 ;
        RECT 6.320 78.675 6.580 78.935 ;
        RECT 7.340 78.675 7.620 78.955 ;
        RECT 9.650 78.685 9.930 78.965 ;
        RECT 1.520 72.245 1.780 72.505 ;
        RECT 2.475 72.245 2.735 72.505 ;
        RECT 3.435 72.245 3.695 72.505 ;
        RECT 4.395 72.245 4.655 72.505 ;
        RECT 5.360 72.240 5.620 72.500 ;
        RECT 6.320 72.240 6.580 72.500 ;
        RECT 7.340 72.240 7.620 72.520 ;
        RECT 9.650 72.250 9.930 72.530 ;
        RECT 1.520 65.810 1.780 66.070 ;
        RECT 2.475 65.810 2.735 66.070 ;
        RECT 3.435 65.810 3.695 66.070 ;
        RECT 4.395 65.810 4.655 66.070 ;
        RECT 5.360 65.805 5.620 66.065 ;
        RECT 6.320 65.805 6.580 66.065 ;
        RECT 7.340 65.805 7.620 66.085 ;
        RECT 9.650 65.815 9.930 66.095 ;
        RECT 1.520 59.375 1.780 59.635 ;
        RECT 2.475 59.375 2.735 59.635 ;
        RECT 3.435 59.375 3.695 59.635 ;
        RECT 4.395 59.375 4.655 59.635 ;
        RECT 5.360 59.370 5.620 59.630 ;
        RECT 6.320 59.370 6.580 59.630 ;
        RECT 7.340 59.370 7.620 59.650 ;
        RECT 9.650 59.380 9.930 59.660 ;
        RECT 1.520 52.940 1.780 53.200 ;
        RECT 2.475 52.940 2.735 53.200 ;
        RECT 3.435 52.940 3.695 53.200 ;
        RECT 4.395 52.940 4.655 53.200 ;
        RECT 5.360 52.935 5.620 53.195 ;
        RECT 6.320 52.935 6.580 53.195 ;
        RECT 7.340 52.935 7.620 53.215 ;
        RECT 9.650 52.945 9.930 53.225 ;
        RECT 1.520 46.505 1.780 46.765 ;
        RECT 2.475 46.505 2.735 46.765 ;
        RECT 3.435 46.505 3.695 46.765 ;
        RECT 4.395 46.505 4.655 46.765 ;
        RECT 5.360 46.500 5.620 46.760 ;
        RECT 6.320 46.500 6.580 46.760 ;
        RECT 7.340 46.500 7.620 46.780 ;
        RECT 9.650 46.510 9.930 46.790 ;
        RECT 1.520 40.070 1.780 40.330 ;
        RECT 2.475 40.070 2.735 40.330 ;
        RECT 3.435 40.070 3.695 40.330 ;
        RECT 4.395 40.070 4.655 40.330 ;
        RECT 5.360 40.065 5.620 40.325 ;
        RECT 6.320 40.065 6.580 40.325 ;
        RECT 7.340 40.065 7.620 40.345 ;
        RECT 9.650 40.075 9.930 40.355 ;
        RECT 1.520 33.635 1.780 33.895 ;
        RECT 2.475 33.635 2.735 33.895 ;
        RECT 3.435 33.635 3.695 33.895 ;
        RECT 4.395 33.635 4.655 33.895 ;
        RECT 5.360 33.630 5.620 33.890 ;
        RECT 6.320 33.630 6.580 33.890 ;
        RECT 7.340 33.630 7.620 33.910 ;
        RECT 9.650 33.640 9.930 33.920 ;
        RECT 1.520 27.200 1.780 27.460 ;
        RECT 2.475 27.200 2.735 27.460 ;
        RECT 3.435 27.200 3.695 27.460 ;
        RECT 4.395 27.200 4.655 27.460 ;
        RECT 5.360 27.195 5.620 27.455 ;
        RECT 6.320 27.195 6.580 27.455 ;
        RECT 7.340 27.195 7.620 27.475 ;
        RECT 9.650 27.205 9.930 27.485 ;
        RECT 1.520 20.765 1.780 21.025 ;
        RECT 2.475 20.765 2.735 21.025 ;
        RECT 3.435 20.765 3.695 21.025 ;
        RECT 4.395 20.765 4.655 21.025 ;
        RECT 5.360 20.760 5.620 21.020 ;
        RECT 6.320 20.760 6.580 21.020 ;
        RECT 7.340 20.760 7.620 21.040 ;
        RECT 9.650 20.770 9.930 21.050 ;
        RECT 1.520 14.330 1.780 14.590 ;
        RECT 2.475 14.330 2.735 14.590 ;
        RECT 3.435 14.330 3.695 14.590 ;
        RECT 4.395 14.330 4.655 14.590 ;
        RECT 5.360 14.325 5.620 14.585 ;
        RECT 6.320 14.325 6.580 14.585 ;
        RECT 7.340 14.325 7.620 14.605 ;
        RECT 9.650 14.335 9.930 14.615 ;
        RECT 1.520 7.895 1.780 8.155 ;
        RECT 2.475 7.895 2.735 8.155 ;
        RECT 3.435 7.895 3.695 8.155 ;
        RECT 4.395 7.895 4.655 8.155 ;
        RECT 5.360 7.890 5.620 8.150 ;
        RECT 6.320 7.890 6.580 8.150 ;
        RECT 7.340 7.890 7.620 8.170 ;
        RECT 9.650 7.900 9.930 8.180 ;
        RECT 1.520 1.460 1.780 1.720 ;
        RECT 2.475 1.460 2.735 1.720 ;
        RECT 3.435 1.460 3.695 1.720 ;
        RECT 4.395 1.460 4.655 1.720 ;
        RECT 5.360 1.455 5.620 1.715 ;
        RECT 6.320 1.455 6.580 1.715 ;
        RECT 7.340 1.455 7.620 1.735 ;
        RECT 9.650 1.465 9.930 1.745 ;
      LAYER met2 ;
        RECT 1.520 201.205 1.780 201.255 ;
        RECT 2.475 201.205 2.735 201.255 ;
        RECT 3.435 201.205 3.695 201.255 ;
        RECT 4.395 201.205 4.655 201.255 ;
        RECT 5.360 201.205 5.620 201.250 ;
        RECT 6.320 201.205 6.580 201.250 ;
        RECT 7.340 201.205 7.620 201.270 ;
        RECT 0.380 200.945 7.630 201.205 ;
        RECT 1.520 200.895 1.780 200.945 ;
        RECT 2.475 200.895 2.735 200.945 ;
        RECT 3.435 200.895 3.695 200.945 ;
        RECT 4.395 200.895 4.655 200.945 ;
        RECT 5.360 200.890 5.620 200.945 ;
        RECT 6.320 200.890 6.580 200.945 ;
        RECT 7.340 200.890 7.620 200.945 ;
        RECT 1.520 194.770 1.780 194.820 ;
        RECT 2.475 194.770 2.735 194.820 ;
        RECT 3.435 194.770 3.695 194.820 ;
        RECT 4.395 194.770 4.655 194.820 ;
        RECT 5.360 194.770 5.620 194.815 ;
        RECT 6.320 194.770 6.580 194.815 ;
        RECT 7.340 194.770 7.620 194.835 ;
        RECT 0.380 194.510 7.630 194.770 ;
        RECT 1.520 194.460 1.780 194.510 ;
        RECT 2.475 194.460 2.735 194.510 ;
        RECT 3.435 194.460 3.695 194.510 ;
        RECT 4.395 194.460 4.655 194.510 ;
        RECT 5.360 194.455 5.620 194.510 ;
        RECT 6.320 194.455 6.580 194.510 ;
        RECT 7.340 194.455 7.620 194.510 ;
        RECT 1.520 188.335 1.780 188.385 ;
        RECT 2.475 188.335 2.735 188.385 ;
        RECT 3.435 188.335 3.695 188.385 ;
        RECT 4.395 188.335 4.655 188.385 ;
        RECT 5.360 188.335 5.620 188.380 ;
        RECT 6.320 188.335 6.580 188.380 ;
        RECT 7.340 188.335 7.620 188.400 ;
        RECT 0.380 188.075 7.630 188.335 ;
        RECT 1.520 188.025 1.780 188.075 ;
        RECT 2.475 188.025 2.735 188.075 ;
        RECT 3.435 188.025 3.695 188.075 ;
        RECT 4.395 188.025 4.655 188.075 ;
        RECT 5.360 188.020 5.620 188.075 ;
        RECT 6.320 188.020 6.580 188.075 ;
        RECT 7.340 188.020 7.620 188.075 ;
        RECT 1.520 181.900 1.780 181.950 ;
        RECT 2.475 181.900 2.735 181.950 ;
        RECT 3.435 181.900 3.695 181.950 ;
        RECT 4.395 181.900 4.655 181.950 ;
        RECT 5.360 181.900 5.620 181.945 ;
        RECT 6.320 181.900 6.580 181.945 ;
        RECT 7.340 181.900 7.620 181.965 ;
        RECT 0.380 181.640 7.630 181.900 ;
        RECT 1.520 181.590 1.780 181.640 ;
        RECT 2.475 181.590 2.735 181.640 ;
        RECT 3.435 181.590 3.695 181.640 ;
        RECT 4.395 181.590 4.655 181.640 ;
        RECT 5.360 181.585 5.620 181.640 ;
        RECT 6.320 181.585 6.580 181.640 ;
        RECT 7.340 181.585 7.620 181.640 ;
        RECT 1.520 175.465 1.780 175.515 ;
        RECT 2.475 175.465 2.735 175.515 ;
        RECT 3.435 175.465 3.695 175.515 ;
        RECT 4.395 175.465 4.655 175.515 ;
        RECT 5.360 175.465 5.620 175.510 ;
        RECT 6.320 175.465 6.580 175.510 ;
        RECT 7.340 175.465 7.620 175.530 ;
        RECT 0.380 175.205 7.630 175.465 ;
        RECT 1.520 175.155 1.780 175.205 ;
        RECT 2.475 175.155 2.735 175.205 ;
        RECT 3.435 175.155 3.695 175.205 ;
        RECT 4.395 175.155 4.655 175.205 ;
        RECT 5.360 175.150 5.620 175.205 ;
        RECT 6.320 175.150 6.580 175.205 ;
        RECT 7.340 175.150 7.620 175.205 ;
        RECT 1.520 169.030 1.780 169.080 ;
        RECT 2.475 169.030 2.735 169.080 ;
        RECT 3.435 169.030 3.695 169.080 ;
        RECT 4.395 169.030 4.655 169.080 ;
        RECT 5.360 169.030 5.620 169.075 ;
        RECT 6.320 169.030 6.580 169.075 ;
        RECT 7.340 169.030 7.620 169.095 ;
        RECT 0.380 168.770 7.630 169.030 ;
        RECT 1.520 168.720 1.780 168.770 ;
        RECT 2.475 168.720 2.735 168.770 ;
        RECT 3.435 168.720 3.695 168.770 ;
        RECT 4.395 168.720 4.655 168.770 ;
        RECT 5.360 168.715 5.620 168.770 ;
        RECT 6.320 168.715 6.580 168.770 ;
        RECT 7.340 168.715 7.620 168.770 ;
        RECT 1.520 162.595 1.780 162.645 ;
        RECT 2.475 162.595 2.735 162.645 ;
        RECT 3.435 162.595 3.695 162.645 ;
        RECT 4.395 162.595 4.655 162.645 ;
        RECT 5.360 162.595 5.620 162.640 ;
        RECT 6.320 162.595 6.580 162.640 ;
        RECT 7.340 162.595 7.620 162.660 ;
        RECT 0.380 162.335 7.630 162.595 ;
        RECT 1.520 162.285 1.780 162.335 ;
        RECT 2.475 162.285 2.735 162.335 ;
        RECT 3.435 162.285 3.695 162.335 ;
        RECT 4.395 162.285 4.655 162.335 ;
        RECT 5.360 162.280 5.620 162.335 ;
        RECT 6.320 162.280 6.580 162.335 ;
        RECT 7.340 162.280 7.620 162.335 ;
        RECT 1.520 156.160 1.780 156.210 ;
        RECT 2.475 156.160 2.735 156.210 ;
        RECT 3.435 156.160 3.695 156.210 ;
        RECT 4.395 156.160 4.655 156.210 ;
        RECT 5.360 156.160 5.620 156.205 ;
        RECT 6.320 156.160 6.580 156.205 ;
        RECT 7.340 156.160 7.620 156.225 ;
        RECT 0.380 155.900 7.630 156.160 ;
        RECT 1.520 155.850 1.780 155.900 ;
        RECT 2.475 155.850 2.735 155.900 ;
        RECT 3.435 155.850 3.695 155.900 ;
        RECT 4.395 155.850 4.655 155.900 ;
        RECT 5.360 155.845 5.620 155.900 ;
        RECT 6.320 155.845 6.580 155.900 ;
        RECT 7.340 155.845 7.620 155.900 ;
        RECT 1.520 149.725 1.780 149.775 ;
        RECT 2.475 149.725 2.735 149.775 ;
        RECT 3.435 149.725 3.695 149.775 ;
        RECT 4.395 149.725 4.655 149.775 ;
        RECT 5.360 149.725 5.620 149.770 ;
        RECT 6.320 149.725 6.580 149.770 ;
        RECT 7.340 149.725 7.620 149.790 ;
        RECT 0.380 149.465 7.630 149.725 ;
        RECT 1.520 149.415 1.780 149.465 ;
        RECT 2.475 149.415 2.735 149.465 ;
        RECT 3.435 149.415 3.695 149.465 ;
        RECT 4.395 149.415 4.655 149.465 ;
        RECT 5.360 149.410 5.620 149.465 ;
        RECT 6.320 149.410 6.580 149.465 ;
        RECT 7.340 149.410 7.620 149.465 ;
        RECT 1.520 143.290 1.780 143.340 ;
        RECT 2.475 143.290 2.735 143.340 ;
        RECT 3.435 143.290 3.695 143.340 ;
        RECT 4.395 143.290 4.655 143.340 ;
        RECT 5.360 143.290 5.620 143.335 ;
        RECT 6.320 143.290 6.580 143.335 ;
        RECT 7.340 143.290 7.620 143.355 ;
        RECT 0.380 143.030 7.630 143.290 ;
        RECT 1.520 142.980 1.780 143.030 ;
        RECT 2.475 142.980 2.735 143.030 ;
        RECT 3.435 142.980 3.695 143.030 ;
        RECT 4.395 142.980 4.655 143.030 ;
        RECT 5.360 142.975 5.620 143.030 ;
        RECT 6.320 142.975 6.580 143.030 ;
        RECT 7.340 142.975 7.620 143.030 ;
        RECT 1.520 136.855 1.780 136.905 ;
        RECT 2.475 136.855 2.735 136.905 ;
        RECT 3.435 136.855 3.695 136.905 ;
        RECT 4.395 136.855 4.655 136.905 ;
        RECT 5.360 136.855 5.620 136.900 ;
        RECT 6.320 136.855 6.580 136.900 ;
        RECT 7.340 136.855 7.620 136.920 ;
        RECT 0.380 136.595 7.630 136.855 ;
        RECT 1.520 136.545 1.780 136.595 ;
        RECT 2.475 136.545 2.735 136.595 ;
        RECT 3.435 136.545 3.695 136.595 ;
        RECT 4.395 136.545 4.655 136.595 ;
        RECT 5.360 136.540 5.620 136.595 ;
        RECT 6.320 136.540 6.580 136.595 ;
        RECT 7.340 136.540 7.620 136.595 ;
        RECT 1.520 130.420 1.780 130.470 ;
        RECT 2.475 130.420 2.735 130.470 ;
        RECT 3.435 130.420 3.695 130.470 ;
        RECT 4.395 130.420 4.655 130.470 ;
        RECT 5.360 130.420 5.620 130.465 ;
        RECT 6.320 130.420 6.580 130.465 ;
        RECT 7.340 130.420 7.620 130.485 ;
        RECT 0.380 130.160 7.630 130.420 ;
        RECT 1.520 130.110 1.780 130.160 ;
        RECT 2.475 130.110 2.735 130.160 ;
        RECT 3.435 130.110 3.695 130.160 ;
        RECT 4.395 130.110 4.655 130.160 ;
        RECT 5.360 130.105 5.620 130.160 ;
        RECT 6.320 130.105 6.580 130.160 ;
        RECT 7.340 130.105 7.620 130.160 ;
        RECT 1.520 123.985 1.780 124.035 ;
        RECT 2.475 123.985 2.735 124.035 ;
        RECT 3.435 123.985 3.695 124.035 ;
        RECT 4.395 123.985 4.655 124.035 ;
        RECT 5.360 123.985 5.620 124.030 ;
        RECT 6.320 123.985 6.580 124.030 ;
        RECT 7.340 123.985 7.620 124.050 ;
        RECT 0.380 123.725 7.630 123.985 ;
        RECT 1.520 123.675 1.780 123.725 ;
        RECT 2.475 123.675 2.735 123.725 ;
        RECT 3.435 123.675 3.695 123.725 ;
        RECT 4.395 123.675 4.655 123.725 ;
        RECT 5.360 123.670 5.620 123.725 ;
        RECT 6.320 123.670 6.580 123.725 ;
        RECT 7.340 123.670 7.620 123.725 ;
        RECT 1.520 117.550 1.780 117.600 ;
        RECT 2.475 117.550 2.735 117.600 ;
        RECT 3.435 117.550 3.695 117.600 ;
        RECT 4.395 117.550 4.655 117.600 ;
        RECT 5.360 117.550 5.620 117.595 ;
        RECT 6.320 117.550 6.580 117.595 ;
        RECT 7.340 117.550 7.620 117.615 ;
        RECT 0.380 117.290 7.630 117.550 ;
        RECT 1.520 117.240 1.780 117.290 ;
        RECT 2.475 117.240 2.735 117.290 ;
        RECT 3.435 117.240 3.695 117.290 ;
        RECT 4.395 117.240 4.655 117.290 ;
        RECT 5.360 117.235 5.620 117.290 ;
        RECT 6.320 117.235 6.580 117.290 ;
        RECT 7.340 117.235 7.620 117.290 ;
        RECT 1.520 111.115 1.780 111.165 ;
        RECT 2.475 111.115 2.735 111.165 ;
        RECT 3.435 111.115 3.695 111.165 ;
        RECT 4.395 111.115 4.655 111.165 ;
        RECT 5.360 111.115 5.620 111.160 ;
        RECT 6.320 111.115 6.580 111.160 ;
        RECT 7.340 111.115 7.620 111.180 ;
        RECT 0.380 110.855 7.630 111.115 ;
        RECT 1.520 110.805 1.780 110.855 ;
        RECT 2.475 110.805 2.735 110.855 ;
        RECT 3.435 110.805 3.695 110.855 ;
        RECT 4.395 110.805 4.655 110.855 ;
        RECT 5.360 110.800 5.620 110.855 ;
        RECT 6.320 110.800 6.580 110.855 ;
        RECT 7.340 110.800 7.620 110.855 ;
        RECT 1.520 104.680 1.780 104.730 ;
        RECT 2.475 104.680 2.735 104.730 ;
        RECT 3.435 104.680 3.695 104.730 ;
        RECT 4.395 104.680 4.655 104.730 ;
        RECT 5.360 104.680 5.620 104.725 ;
        RECT 6.320 104.680 6.580 104.725 ;
        RECT 7.340 104.680 7.620 104.745 ;
        RECT 0.380 104.420 7.630 104.680 ;
        RECT 1.520 104.370 1.780 104.420 ;
        RECT 2.475 104.370 2.735 104.420 ;
        RECT 3.435 104.370 3.695 104.420 ;
        RECT 4.395 104.370 4.655 104.420 ;
        RECT 5.360 104.365 5.620 104.420 ;
        RECT 6.320 104.365 6.580 104.420 ;
        RECT 7.340 104.365 7.620 104.420 ;
        RECT 1.520 98.245 1.780 98.295 ;
        RECT 2.475 98.245 2.735 98.295 ;
        RECT 3.435 98.245 3.695 98.295 ;
        RECT 4.395 98.245 4.655 98.295 ;
        RECT 5.360 98.245 5.620 98.290 ;
        RECT 6.320 98.245 6.580 98.290 ;
        RECT 7.340 98.245 7.620 98.310 ;
        RECT 0.380 97.985 7.630 98.245 ;
        RECT 1.520 97.935 1.780 97.985 ;
        RECT 2.475 97.935 2.735 97.985 ;
        RECT 3.435 97.935 3.695 97.985 ;
        RECT 4.395 97.935 4.655 97.985 ;
        RECT 5.360 97.930 5.620 97.985 ;
        RECT 6.320 97.930 6.580 97.985 ;
        RECT 7.340 97.930 7.620 97.985 ;
        RECT 1.520 91.810 1.780 91.860 ;
        RECT 2.475 91.810 2.735 91.860 ;
        RECT 3.435 91.810 3.695 91.860 ;
        RECT 4.395 91.810 4.655 91.860 ;
        RECT 5.360 91.810 5.620 91.855 ;
        RECT 6.320 91.810 6.580 91.855 ;
        RECT 7.340 91.810 7.620 91.875 ;
        RECT 0.380 91.550 7.630 91.810 ;
        RECT 1.520 91.500 1.780 91.550 ;
        RECT 2.475 91.500 2.735 91.550 ;
        RECT 3.435 91.500 3.695 91.550 ;
        RECT 4.395 91.500 4.655 91.550 ;
        RECT 5.360 91.495 5.620 91.550 ;
        RECT 6.320 91.495 6.580 91.550 ;
        RECT 7.340 91.495 7.620 91.550 ;
        RECT 1.520 85.375 1.780 85.425 ;
        RECT 2.475 85.375 2.735 85.425 ;
        RECT 3.435 85.375 3.695 85.425 ;
        RECT 4.395 85.375 4.655 85.425 ;
        RECT 5.360 85.375 5.620 85.420 ;
        RECT 6.320 85.375 6.580 85.420 ;
        RECT 7.340 85.375 7.620 85.440 ;
        RECT 0.380 85.115 7.630 85.375 ;
        RECT 1.520 85.065 1.780 85.115 ;
        RECT 2.475 85.065 2.735 85.115 ;
        RECT 3.435 85.065 3.695 85.115 ;
        RECT 4.395 85.065 4.655 85.115 ;
        RECT 5.360 85.060 5.620 85.115 ;
        RECT 6.320 85.060 6.580 85.115 ;
        RECT 7.340 85.060 7.620 85.115 ;
        RECT 1.520 78.940 1.780 78.990 ;
        RECT 2.475 78.940 2.735 78.990 ;
        RECT 3.435 78.940 3.695 78.990 ;
        RECT 4.395 78.940 4.655 78.990 ;
        RECT 5.360 78.940 5.620 78.985 ;
        RECT 6.320 78.940 6.580 78.985 ;
        RECT 7.340 78.940 7.620 79.005 ;
        RECT 0.380 78.680 7.630 78.940 ;
        RECT 1.520 78.630 1.780 78.680 ;
        RECT 2.475 78.630 2.735 78.680 ;
        RECT 3.435 78.630 3.695 78.680 ;
        RECT 4.395 78.630 4.655 78.680 ;
        RECT 5.360 78.625 5.620 78.680 ;
        RECT 6.320 78.625 6.580 78.680 ;
        RECT 7.340 78.625 7.620 78.680 ;
        RECT 1.520 72.505 1.780 72.555 ;
        RECT 2.475 72.505 2.735 72.555 ;
        RECT 3.435 72.505 3.695 72.555 ;
        RECT 4.395 72.505 4.655 72.555 ;
        RECT 5.360 72.505 5.620 72.550 ;
        RECT 6.320 72.505 6.580 72.550 ;
        RECT 7.340 72.505 7.620 72.570 ;
        RECT 0.380 72.245 7.630 72.505 ;
        RECT 1.520 72.195 1.780 72.245 ;
        RECT 2.475 72.195 2.735 72.245 ;
        RECT 3.435 72.195 3.695 72.245 ;
        RECT 4.395 72.195 4.655 72.245 ;
        RECT 5.360 72.190 5.620 72.245 ;
        RECT 6.320 72.190 6.580 72.245 ;
        RECT 7.340 72.190 7.620 72.245 ;
        RECT 1.520 66.070 1.780 66.120 ;
        RECT 2.475 66.070 2.735 66.120 ;
        RECT 3.435 66.070 3.695 66.120 ;
        RECT 4.395 66.070 4.655 66.120 ;
        RECT 5.360 66.070 5.620 66.115 ;
        RECT 6.320 66.070 6.580 66.115 ;
        RECT 7.340 66.070 7.620 66.135 ;
        RECT 0.380 65.810 7.630 66.070 ;
        RECT 1.520 65.760 1.780 65.810 ;
        RECT 2.475 65.760 2.735 65.810 ;
        RECT 3.435 65.760 3.695 65.810 ;
        RECT 4.395 65.760 4.655 65.810 ;
        RECT 5.360 65.755 5.620 65.810 ;
        RECT 6.320 65.755 6.580 65.810 ;
        RECT 7.340 65.755 7.620 65.810 ;
        RECT 1.520 59.635 1.780 59.685 ;
        RECT 2.475 59.635 2.735 59.685 ;
        RECT 3.435 59.635 3.695 59.685 ;
        RECT 4.395 59.635 4.655 59.685 ;
        RECT 5.360 59.635 5.620 59.680 ;
        RECT 6.320 59.635 6.580 59.680 ;
        RECT 7.340 59.635 7.620 59.700 ;
        RECT 0.380 59.375 7.630 59.635 ;
        RECT 1.520 59.325 1.780 59.375 ;
        RECT 2.475 59.325 2.735 59.375 ;
        RECT 3.435 59.325 3.695 59.375 ;
        RECT 4.395 59.325 4.655 59.375 ;
        RECT 5.360 59.320 5.620 59.375 ;
        RECT 6.320 59.320 6.580 59.375 ;
        RECT 7.340 59.320 7.620 59.375 ;
        RECT 1.520 53.200 1.780 53.250 ;
        RECT 2.475 53.200 2.735 53.250 ;
        RECT 3.435 53.200 3.695 53.250 ;
        RECT 4.395 53.200 4.655 53.250 ;
        RECT 5.360 53.200 5.620 53.245 ;
        RECT 6.320 53.200 6.580 53.245 ;
        RECT 7.340 53.200 7.620 53.265 ;
        RECT 0.380 52.940 7.630 53.200 ;
        RECT 1.520 52.890 1.780 52.940 ;
        RECT 2.475 52.890 2.735 52.940 ;
        RECT 3.435 52.890 3.695 52.940 ;
        RECT 4.395 52.890 4.655 52.940 ;
        RECT 5.360 52.885 5.620 52.940 ;
        RECT 6.320 52.885 6.580 52.940 ;
        RECT 7.340 52.885 7.620 52.940 ;
        RECT 1.520 46.765 1.780 46.815 ;
        RECT 2.475 46.765 2.735 46.815 ;
        RECT 3.435 46.765 3.695 46.815 ;
        RECT 4.395 46.765 4.655 46.815 ;
        RECT 5.360 46.765 5.620 46.810 ;
        RECT 6.320 46.765 6.580 46.810 ;
        RECT 7.340 46.765 7.620 46.830 ;
        RECT 0.380 46.505 7.630 46.765 ;
        RECT 1.520 46.455 1.780 46.505 ;
        RECT 2.475 46.455 2.735 46.505 ;
        RECT 3.435 46.455 3.695 46.505 ;
        RECT 4.395 46.455 4.655 46.505 ;
        RECT 5.360 46.450 5.620 46.505 ;
        RECT 6.320 46.450 6.580 46.505 ;
        RECT 7.340 46.450 7.620 46.505 ;
        RECT 1.520 40.330 1.780 40.380 ;
        RECT 2.475 40.330 2.735 40.380 ;
        RECT 3.435 40.330 3.695 40.380 ;
        RECT 4.395 40.330 4.655 40.380 ;
        RECT 5.360 40.330 5.620 40.375 ;
        RECT 6.320 40.330 6.580 40.375 ;
        RECT 7.340 40.330 7.620 40.395 ;
        RECT 0.380 40.070 7.630 40.330 ;
        RECT 1.520 40.020 1.780 40.070 ;
        RECT 2.475 40.020 2.735 40.070 ;
        RECT 3.435 40.020 3.695 40.070 ;
        RECT 4.395 40.020 4.655 40.070 ;
        RECT 5.360 40.015 5.620 40.070 ;
        RECT 6.320 40.015 6.580 40.070 ;
        RECT 7.340 40.015 7.620 40.070 ;
        RECT 1.520 33.895 1.780 33.945 ;
        RECT 2.475 33.895 2.735 33.945 ;
        RECT 3.435 33.895 3.695 33.945 ;
        RECT 4.395 33.895 4.655 33.945 ;
        RECT 5.360 33.895 5.620 33.940 ;
        RECT 6.320 33.895 6.580 33.940 ;
        RECT 7.340 33.895 7.620 33.960 ;
        RECT 0.380 33.635 7.630 33.895 ;
        RECT 1.520 33.585 1.780 33.635 ;
        RECT 2.475 33.585 2.735 33.635 ;
        RECT 3.435 33.585 3.695 33.635 ;
        RECT 4.395 33.585 4.655 33.635 ;
        RECT 5.360 33.580 5.620 33.635 ;
        RECT 6.320 33.580 6.580 33.635 ;
        RECT 7.340 33.580 7.620 33.635 ;
        RECT 1.520 27.460 1.780 27.510 ;
        RECT 2.475 27.460 2.735 27.510 ;
        RECT 3.435 27.460 3.695 27.510 ;
        RECT 4.395 27.460 4.655 27.510 ;
        RECT 5.360 27.460 5.620 27.505 ;
        RECT 6.320 27.460 6.580 27.505 ;
        RECT 7.340 27.460 7.620 27.525 ;
        RECT 0.380 27.200 7.630 27.460 ;
        RECT 1.520 27.150 1.780 27.200 ;
        RECT 2.475 27.150 2.735 27.200 ;
        RECT 3.435 27.150 3.695 27.200 ;
        RECT 4.395 27.150 4.655 27.200 ;
        RECT 5.360 27.145 5.620 27.200 ;
        RECT 6.320 27.145 6.580 27.200 ;
        RECT 7.340 27.145 7.620 27.200 ;
        RECT 1.520 21.025 1.780 21.075 ;
        RECT 2.475 21.025 2.735 21.075 ;
        RECT 3.435 21.025 3.695 21.075 ;
        RECT 4.395 21.025 4.655 21.075 ;
        RECT 5.360 21.025 5.620 21.070 ;
        RECT 6.320 21.025 6.580 21.070 ;
        RECT 7.340 21.025 7.620 21.090 ;
        RECT 0.380 20.765 7.630 21.025 ;
        RECT 1.520 20.715 1.780 20.765 ;
        RECT 2.475 20.715 2.735 20.765 ;
        RECT 3.435 20.715 3.695 20.765 ;
        RECT 4.395 20.715 4.655 20.765 ;
        RECT 5.360 20.710 5.620 20.765 ;
        RECT 6.320 20.710 6.580 20.765 ;
        RECT 7.340 20.710 7.620 20.765 ;
        RECT 1.520 14.590 1.780 14.640 ;
        RECT 2.475 14.590 2.735 14.640 ;
        RECT 3.435 14.590 3.695 14.640 ;
        RECT 4.395 14.590 4.655 14.640 ;
        RECT 5.360 14.590 5.620 14.635 ;
        RECT 6.320 14.590 6.580 14.635 ;
        RECT 7.340 14.590 7.620 14.655 ;
        RECT 0.380 14.330 7.630 14.590 ;
        RECT 1.520 14.280 1.780 14.330 ;
        RECT 2.475 14.280 2.735 14.330 ;
        RECT 3.435 14.280 3.695 14.330 ;
        RECT 4.395 14.280 4.655 14.330 ;
        RECT 5.360 14.275 5.620 14.330 ;
        RECT 6.320 14.275 6.580 14.330 ;
        RECT 7.340 14.275 7.620 14.330 ;
        RECT 1.520 8.155 1.780 8.205 ;
        RECT 2.475 8.155 2.735 8.205 ;
        RECT 3.435 8.155 3.695 8.205 ;
        RECT 4.395 8.155 4.655 8.205 ;
        RECT 5.360 8.155 5.620 8.200 ;
        RECT 6.320 8.155 6.580 8.200 ;
        RECT 7.340 8.155 7.620 8.220 ;
        RECT 0.380 7.895 7.630 8.155 ;
        RECT 1.520 7.845 1.780 7.895 ;
        RECT 2.475 7.845 2.735 7.895 ;
        RECT 3.435 7.845 3.695 7.895 ;
        RECT 4.395 7.845 4.655 7.895 ;
        RECT 5.360 7.840 5.620 7.895 ;
        RECT 6.320 7.840 6.580 7.895 ;
        RECT 7.340 7.840 7.620 7.895 ;
        RECT 1.520 1.720 1.780 1.770 ;
        RECT 2.475 1.720 2.735 1.770 ;
        RECT 3.435 1.720 3.695 1.770 ;
        RECT 4.395 1.720 4.655 1.770 ;
        RECT 5.360 1.720 5.620 1.765 ;
        RECT 6.320 1.720 6.580 1.765 ;
        RECT 7.340 1.720 7.620 1.785 ;
        RECT 0.380 1.460 7.630 1.720 ;
        RECT 1.520 1.410 1.780 1.460 ;
        RECT 2.475 1.410 2.735 1.460 ;
        RECT 3.435 1.410 3.695 1.460 ;
        RECT 4.395 1.410 4.655 1.460 ;
        RECT 5.360 1.405 5.620 1.460 ;
        RECT 6.320 1.405 6.580 1.460 ;
        RECT 7.340 1.405 7.620 1.460 ;
        RECT 9.650 0.725 9.930 206.760 ;
    END
  END s_en
  PIN s_en_b
    DIRECTION INOUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 65.279999 ;
    PORT
      LAYER li1 ;
        RECT 1.485 205.020 1.815 205.190 ;
        RECT 2.445 205.020 2.775 205.190 ;
        RECT 3.405 205.020 3.735 205.190 ;
        RECT 4.365 205.020 4.695 205.190 ;
        RECT 5.325 205.020 5.655 205.190 ;
        RECT 6.285 205.020 6.615 205.190 ;
        RECT 1.485 198.585 1.815 198.755 ;
        RECT 2.445 198.585 2.775 198.755 ;
        RECT 3.405 198.585 3.735 198.755 ;
        RECT 4.365 198.585 4.695 198.755 ;
        RECT 5.325 198.585 5.655 198.755 ;
        RECT 6.285 198.585 6.615 198.755 ;
        RECT 1.485 192.150 1.815 192.320 ;
        RECT 2.445 192.150 2.775 192.320 ;
        RECT 3.405 192.150 3.735 192.320 ;
        RECT 4.365 192.150 4.695 192.320 ;
        RECT 5.325 192.150 5.655 192.320 ;
        RECT 6.285 192.150 6.615 192.320 ;
        RECT 1.485 185.715 1.815 185.885 ;
        RECT 2.445 185.715 2.775 185.885 ;
        RECT 3.405 185.715 3.735 185.885 ;
        RECT 4.365 185.715 4.695 185.885 ;
        RECT 5.325 185.715 5.655 185.885 ;
        RECT 6.285 185.715 6.615 185.885 ;
        RECT 1.485 179.280 1.815 179.450 ;
        RECT 2.445 179.280 2.775 179.450 ;
        RECT 3.405 179.280 3.735 179.450 ;
        RECT 4.365 179.280 4.695 179.450 ;
        RECT 5.325 179.280 5.655 179.450 ;
        RECT 6.285 179.280 6.615 179.450 ;
        RECT 1.485 172.845 1.815 173.015 ;
        RECT 2.445 172.845 2.775 173.015 ;
        RECT 3.405 172.845 3.735 173.015 ;
        RECT 4.365 172.845 4.695 173.015 ;
        RECT 5.325 172.845 5.655 173.015 ;
        RECT 6.285 172.845 6.615 173.015 ;
        RECT 1.485 166.410 1.815 166.580 ;
        RECT 2.445 166.410 2.775 166.580 ;
        RECT 3.405 166.410 3.735 166.580 ;
        RECT 4.365 166.410 4.695 166.580 ;
        RECT 5.325 166.410 5.655 166.580 ;
        RECT 6.285 166.410 6.615 166.580 ;
        RECT 1.485 159.975 1.815 160.145 ;
        RECT 2.445 159.975 2.775 160.145 ;
        RECT 3.405 159.975 3.735 160.145 ;
        RECT 4.365 159.975 4.695 160.145 ;
        RECT 5.325 159.975 5.655 160.145 ;
        RECT 6.285 159.975 6.615 160.145 ;
        RECT 1.485 153.540 1.815 153.710 ;
        RECT 2.445 153.540 2.775 153.710 ;
        RECT 3.405 153.540 3.735 153.710 ;
        RECT 4.365 153.540 4.695 153.710 ;
        RECT 5.325 153.540 5.655 153.710 ;
        RECT 6.285 153.540 6.615 153.710 ;
        RECT 1.485 147.105 1.815 147.275 ;
        RECT 2.445 147.105 2.775 147.275 ;
        RECT 3.405 147.105 3.735 147.275 ;
        RECT 4.365 147.105 4.695 147.275 ;
        RECT 5.325 147.105 5.655 147.275 ;
        RECT 6.285 147.105 6.615 147.275 ;
        RECT 1.485 140.670 1.815 140.840 ;
        RECT 2.445 140.670 2.775 140.840 ;
        RECT 3.405 140.670 3.735 140.840 ;
        RECT 4.365 140.670 4.695 140.840 ;
        RECT 5.325 140.670 5.655 140.840 ;
        RECT 6.285 140.670 6.615 140.840 ;
        RECT 1.485 134.235 1.815 134.405 ;
        RECT 2.445 134.235 2.775 134.405 ;
        RECT 3.405 134.235 3.735 134.405 ;
        RECT 4.365 134.235 4.695 134.405 ;
        RECT 5.325 134.235 5.655 134.405 ;
        RECT 6.285 134.235 6.615 134.405 ;
        RECT 1.485 127.800 1.815 127.970 ;
        RECT 2.445 127.800 2.775 127.970 ;
        RECT 3.405 127.800 3.735 127.970 ;
        RECT 4.365 127.800 4.695 127.970 ;
        RECT 5.325 127.800 5.655 127.970 ;
        RECT 6.285 127.800 6.615 127.970 ;
        RECT 1.485 121.365 1.815 121.535 ;
        RECT 2.445 121.365 2.775 121.535 ;
        RECT 3.405 121.365 3.735 121.535 ;
        RECT 4.365 121.365 4.695 121.535 ;
        RECT 5.325 121.365 5.655 121.535 ;
        RECT 6.285 121.365 6.615 121.535 ;
        RECT 1.485 114.930 1.815 115.100 ;
        RECT 2.445 114.930 2.775 115.100 ;
        RECT 3.405 114.930 3.735 115.100 ;
        RECT 4.365 114.930 4.695 115.100 ;
        RECT 5.325 114.930 5.655 115.100 ;
        RECT 6.285 114.930 6.615 115.100 ;
        RECT 1.485 108.495 1.815 108.665 ;
        RECT 2.445 108.495 2.775 108.665 ;
        RECT 3.405 108.495 3.735 108.665 ;
        RECT 4.365 108.495 4.695 108.665 ;
        RECT 5.325 108.495 5.655 108.665 ;
        RECT 6.285 108.495 6.615 108.665 ;
        RECT 1.485 102.060 1.815 102.230 ;
        RECT 2.445 102.060 2.775 102.230 ;
        RECT 3.405 102.060 3.735 102.230 ;
        RECT 4.365 102.060 4.695 102.230 ;
        RECT 5.325 102.060 5.655 102.230 ;
        RECT 6.285 102.060 6.615 102.230 ;
        RECT 1.485 95.625 1.815 95.795 ;
        RECT 2.445 95.625 2.775 95.795 ;
        RECT 3.405 95.625 3.735 95.795 ;
        RECT 4.365 95.625 4.695 95.795 ;
        RECT 5.325 95.625 5.655 95.795 ;
        RECT 6.285 95.625 6.615 95.795 ;
        RECT 1.485 89.190 1.815 89.360 ;
        RECT 2.445 89.190 2.775 89.360 ;
        RECT 3.405 89.190 3.735 89.360 ;
        RECT 4.365 89.190 4.695 89.360 ;
        RECT 5.325 89.190 5.655 89.360 ;
        RECT 6.285 89.190 6.615 89.360 ;
        RECT 1.485 82.755 1.815 82.925 ;
        RECT 2.445 82.755 2.775 82.925 ;
        RECT 3.405 82.755 3.735 82.925 ;
        RECT 4.365 82.755 4.695 82.925 ;
        RECT 5.325 82.755 5.655 82.925 ;
        RECT 6.285 82.755 6.615 82.925 ;
        RECT 1.485 76.320 1.815 76.490 ;
        RECT 2.445 76.320 2.775 76.490 ;
        RECT 3.405 76.320 3.735 76.490 ;
        RECT 4.365 76.320 4.695 76.490 ;
        RECT 5.325 76.320 5.655 76.490 ;
        RECT 6.285 76.320 6.615 76.490 ;
        RECT 1.485 69.885 1.815 70.055 ;
        RECT 2.445 69.885 2.775 70.055 ;
        RECT 3.405 69.885 3.735 70.055 ;
        RECT 4.365 69.885 4.695 70.055 ;
        RECT 5.325 69.885 5.655 70.055 ;
        RECT 6.285 69.885 6.615 70.055 ;
        RECT 1.485 63.450 1.815 63.620 ;
        RECT 2.445 63.450 2.775 63.620 ;
        RECT 3.405 63.450 3.735 63.620 ;
        RECT 4.365 63.450 4.695 63.620 ;
        RECT 5.325 63.450 5.655 63.620 ;
        RECT 6.285 63.450 6.615 63.620 ;
        RECT 1.485 57.015 1.815 57.185 ;
        RECT 2.445 57.015 2.775 57.185 ;
        RECT 3.405 57.015 3.735 57.185 ;
        RECT 4.365 57.015 4.695 57.185 ;
        RECT 5.325 57.015 5.655 57.185 ;
        RECT 6.285 57.015 6.615 57.185 ;
        RECT 1.485 50.580 1.815 50.750 ;
        RECT 2.445 50.580 2.775 50.750 ;
        RECT 3.405 50.580 3.735 50.750 ;
        RECT 4.365 50.580 4.695 50.750 ;
        RECT 5.325 50.580 5.655 50.750 ;
        RECT 6.285 50.580 6.615 50.750 ;
        RECT 1.485 44.145 1.815 44.315 ;
        RECT 2.445 44.145 2.775 44.315 ;
        RECT 3.405 44.145 3.735 44.315 ;
        RECT 4.365 44.145 4.695 44.315 ;
        RECT 5.325 44.145 5.655 44.315 ;
        RECT 6.285 44.145 6.615 44.315 ;
        RECT 1.485 37.710 1.815 37.880 ;
        RECT 2.445 37.710 2.775 37.880 ;
        RECT 3.405 37.710 3.735 37.880 ;
        RECT 4.365 37.710 4.695 37.880 ;
        RECT 5.325 37.710 5.655 37.880 ;
        RECT 6.285 37.710 6.615 37.880 ;
        RECT 1.485 31.275 1.815 31.445 ;
        RECT 2.445 31.275 2.775 31.445 ;
        RECT 3.405 31.275 3.735 31.445 ;
        RECT 4.365 31.275 4.695 31.445 ;
        RECT 5.325 31.275 5.655 31.445 ;
        RECT 6.285 31.275 6.615 31.445 ;
        RECT 1.485 24.840 1.815 25.010 ;
        RECT 2.445 24.840 2.775 25.010 ;
        RECT 3.405 24.840 3.735 25.010 ;
        RECT 4.365 24.840 4.695 25.010 ;
        RECT 5.325 24.840 5.655 25.010 ;
        RECT 6.285 24.840 6.615 25.010 ;
        RECT 1.485 18.405 1.815 18.575 ;
        RECT 2.445 18.405 2.775 18.575 ;
        RECT 3.405 18.405 3.735 18.575 ;
        RECT 4.365 18.405 4.695 18.575 ;
        RECT 5.325 18.405 5.655 18.575 ;
        RECT 6.285 18.405 6.615 18.575 ;
        RECT 1.485 11.970 1.815 12.140 ;
        RECT 2.445 11.970 2.775 12.140 ;
        RECT 3.405 11.970 3.735 12.140 ;
        RECT 4.365 11.970 4.695 12.140 ;
        RECT 5.325 11.970 5.655 12.140 ;
        RECT 6.285 11.970 6.615 12.140 ;
        RECT 1.485 5.535 1.815 5.705 ;
        RECT 2.445 5.535 2.775 5.705 ;
        RECT 3.405 5.535 3.735 5.705 ;
        RECT 4.365 5.535 4.695 5.705 ;
        RECT 5.325 5.535 5.655 5.705 ;
        RECT 6.285 5.535 6.615 5.705 ;
      LAYER mcon ;
        RECT 1.565 205.020 1.735 205.190 ;
        RECT 2.525 205.020 2.695 205.190 ;
        RECT 3.485 205.020 3.655 205.190 ;
        RECT 4.445 205.020 4.615 205.190 ;
        RECT 5.405 205.020 5.575 205.190 ;
        RECT 6.365 205.020 6.535 205.190 ;
        RECT 1.565 198.585 1.735 198.755 ;
        RECT 2.525 198.585 2.695 198.755 ;
        RECT 3.485 198.585 3.655 198.755 ;
        RECT 4.445 198.585 4.615 198.755 ;
        RECT 5.405 198.585 5.575 198.755 ;
        RECT 6.365 198.585 6.535 198.755 ;
        RECT 1.565 192.150 1.735 192.320 ;
        RECT 2.525 192.150 2.695 192.320 ;
        RECT 3.485 192.150 3.655 192.320 ;
        RECT 4.445 192.150 4.615 192.320 ;
        RECT 5.405 192.150 5.575 192.320 ;
        RECT 6.365 192.150 6.535 192.320 ;
        RECT 1.565 185.715 1.735 185.885 ;
        RECT 2.525 185.715 2.695 185.885 ;
        RECT 3.485 185.715 3.655 185.885 ;
        RECT 4.445 185.715 4.615 185.885 ;
        RECT 5.405 185.715 5.575 185.885 ;
        RECT 6.365 185.715 6.535 185.885 ;
        RECT 1.565 179.280 1.735 179.450 ;
        RECT 2.525 179.280 2.695 179.450 ;
        RECT 3.485 179.280 3.655 179.450 ;
        RECT 4.445 179.280 4.615 179.450 ;
        RECT 5.405 179.280 5.575 179.450 ;
        RECT 6.365 179.280 6.535 179.450 ;
        RECT 1.565 172.845 1.735 173.015 ;
        RECT 2.525 172.845 2.695 173.015 ;
        RECT 3.485 172.845 3.655 173.015 ;
        RECT 4.445 172.845 4.615 173.015 ;
        RECT 5.405 172.845 5.575 173.015 ;
        RECT 6.365 172.845 6.535 173.015 ;
        RECT 1.565 166.410 1.735 166.580 ;
        RECT 2.525 166.410 2.695 166.580 ;
        RECT 3.485 166.410 3.655 166.580 ;
        RECT 4.445 166.410 4.615 166.580 ;
        RECT 5.405 166.410 5.575 166.580 ;
        RECT 6.365 166.410 6.535 166.580 ;
        RECT 1.565 159.975 1.735 160.145 ;
        RECT 2.525 159.975 2.695 160.145 ;
        RECT 3.485 159.975 3.655 160.145 ;
        RECT 4.445 159.975 4.615 160.145 ;
        RECT 5.405 159.975 5.575 160.145 ;
        RECT 6.365 159.975 6.535 160.145 ;
        RECT 1.565 153.540 1.735 153.710 ;
        RECT 2.525 153.540 2.695 153.710 ;
        RECT 3.485 153.540 3.655 153.710 ;
        RECT 4.445 153.540 4.615 153.710 ;
        RECT 5.405 153.540 5.575 153.710 ;
        RECT 6.365 153.540 6.535 153.710 ;
        RECT 1.565 147.105 1.735 147.275 ;
        RECT 2.525 147.105 2.695 147.275 ;
        RECT 3.485 147.105 3.655 147.275 ;
        RECT 4.445 147.105 4.615 147.275 ;
        RECT 5.405 147.105 5.575 147.275 ;
        RECT 6.365 147.105 6.535 147.275 ;
        RECT 1.565 140.670 1.735 140.840 ;
        RECT 2.525 140.670 2.695 140.840 ;
        RECT 3.485 140.670 3.655 140.840 ;
        RECT 4.445 140.670 4.615 140.840 ;
        RECT 5.405 140.670 5.575 140.840 ;
        RECT 6.365 140.670 6.535 140.840 ;
        RECT 1.565 134.235 1.735 134.405 ;
        RECT 2.525 134.235 2.695 134.405 ;
        RECT 3.485 134.235 3.655 134.405 ;
        RECT 4.445 134.235 4.615 134.405 ;
        RECT 5.405 134.235 5.575 134.405 ;
        RECT 6.365 134.235 6.535 134.405 ;
        RECT 1.565 127.800 1.735 127.970 ;
        RECT 2.525 127.800 2.695 127.970 ;
        RECT 3.485 127.800 3.655 127.970 ;
        RECT 4.445 127.800 4.615 127.970 ;
        RECT 5.405 127.800 5.575 127.970 ;
        RECT 6.365 127.800 6.535 127.970 ;
        RECT 1.565 121.365 1.735 121.535 ;
        RECT 2.525 121.365 2.695 121.535 ;
        RECT 3.485 121.365 3.655 121.535 ;
        RECT 4.445 121.365 4.615 121.535 ;
        RECT 5.405 121.365 5.575 121.535 ;
        RECT 6.365 121.365 6.535 121.535 ;
        RECT 1.565 114.930 1.735 115.100 ;
        RECT 2.525 114.930 2.695 115.100 ;
        RECT 3.485 114.930 3.655 115.100 ;
        RECT 4.445 114.930 4.615 115.100 ;
        RECT 5.405 114.930 5.575 115.100 ;
        RECT 6.365 114.930 6.535 115.100 ;
        RECT 1.565 108.495 1.735 108.665 ;
        RECT 2.525 108.495 2.695 108.665 ;
        RECT 3.485 108.495 3.655 108.665 ;
        RECT 4.445 108.495 4.615 108.665 ;
        RECT 5.405 108.495 5.575 108.665 ;
        RECT 6.365 108.495 6.535 108.665 ;
        RECT 1.565 102.060 1.735 102.230 ;
        RECT 2.525 102.060 2.695 102.230 ;
        RECT 3.485 102.060 3.655 102.230 ;
        RECT 4.445 102.060 4.615 102.230 ;
        RECT 5.405 102.060 5.575 102.230 ;
        RECT 6.365 102.060 6.535 102.230 ;
        RECT 1.565 95.625 1.735 95.795 ;
        RECT 2.525 95.625 2.695 95.795 ;
        RECT 3.485 95.625 3.655 95.795 ;
        RECT 4.445 95.625 4.615 95.795 ;
        RECT 5.405 95.625 5.575 95.795 ;
        RECT 6.365 95.625 6.535 95.795 ;
        RECT 1.565 89.190 1.735 89.360 ;
        RECT 2.525 89.190 2.695 89.360 ;
        RECT 3.485 89.190 3.655 89.360 ;
        RECT 4.445 89.190 4.615 89.360 ;
        RECT 5.405 89.190 5.575 89.360 ;
        RECT 6.365 89.190 6.535 89.360 ;
        RECT 1.565 82.755 1.735 82.925 ;
        RECT 2.525 82.755 2.695 82.925 ;
        RECT 3.485 82.755 3.655 82.925 ;
        RECT 4.445 82.755 4.615 82.925 ;
        RECT 5.405 82.755 5.575 82.925 ;
        RECT 6.365 82.755 6.535 82.925 ;
        RECT 1.565 76.320 1.735 76.490 ;
        RECT 2.525 76.320 2.695 76.490 ;
        RECT 3.485 76.320 3.655 76.490 ;
        RECT 4.445 76.320 4.615 76.490 ;
        RECT 5.405 76.320 5.575 76.490 ;
        RECT 6.365 76.320 6.535 76.490 ;
        RECT 1.565 69.885 1.735 70.055 ;
        RECT 2.525 69.885 2.695 70.055 ;
        RECT 3.485 69.885 3.655 70.055 ;
        RECT 4.445 69.885 4.615 70.055 ;
        RECT 5.405 69.885 5.575 70.055 ;
        RECT 6.365 69.885 6.535 70.055 ;
        RECT 1.565 63.450 1.735 63.620 ;
        RECT 2.525 63.450 2.695 63.620 ;
        RECT 3.485 63.450 3.655 63.620 ;
        RECT 4.445 63.450 4.615 63.620 ;
        RECT 5.405 63.450 5.575 63.620 ;
        RECT 6.365 63.450 6.535 63.620 ;
        RECT 1.565 57.015 1.735 57.185 ;
        RECT 2.525 57.015 2.695 57.185 ;
        RECT 3.485 57.015 3.655 57.185 ;
        RECT 4.445 57.015 4.615 57.185 ;
        RECT 5.405 57.015 5.575 57.185 ;
        RECT 6.365 57.015 6.535 57.185 ;
        RECT 1.565 50.580 1.735 50.750 ;
        RECT 2.525 50.580 2.695 50.750 ;
        RECT 3.485 50.580 3.655 50.750 ;
        RECT 4.445 50.580 4.615 50.750 ;
        RECT 5.405 50.580 5.575 50.750 ;
        RECT 6.365 50.580 6.535 50.750 ;
        RECT 1.565 44.145 1.735 44.315 ;
        RECT 2.525 44.145 2.695 44.315 ;
        RECT 3.485 44.145 3.655 44.315 ;
        RECT 4.445 44.145 4.615 44.315 ;
        RECT 5.405 44.145 5.575 44.315 ;
        RECT 6.365 44.145 6.535 44.315 ;
        RECT 1.565 37.710 1.735 37.880 ;
        RECT 2.525 37.710 2.695 37.880 ;
        RECT 3.485 37.710 3.655 37.880 ;
        RECT 4.445 37.710 4.615 37.880 ;
        RECT 5.405 37.710 5.575 37.880 ;
        RECT 6.365 37.710 6.535 37.880 ;
        RECT 1.565 31.275 1.735 31.445 ;
        RECT 2.525 31.275 2.695 31.445 ;
        RECT 3.485 31.275 3.655 31.445 ;
        RECT 4.445 31.275 4.615 31.445 ;
        RECT 5.405 31.275 5.575 31.445 ;
        RECT 6.365 31.275 6.535 31.445 ;
        RECT 1.565 24.840 1.735 25.010 ;
        RECT 2.525 24.840 2.695 25.010 ;
        RECT 3.485 24.840 3.655 25.010 ;
        RECT 4.445 24.840 4.615 25.010 ;
        RECT 5.405 24.840 5.575 25.010 ;
        RECT 6.365 24.840 6.535 25.010 ;
        RECT 1.565 18.405 1.735 18.575 ;
        RECT 2.525 18.405 2.695 18.575 ;
        RECT 3.485 18.405 3.655 18.575 ;
        RECT 4.445 18.405 4.615 18.575 ;
        RECT 5.405 18.405 5.575 18.575 ;
        RECT 6.365 18.405 6.535 18.575 ;
        RECT 1.565 11.970 1.735 12.140 ;
        RECT 2.525 11.970 2.695 12.140 ;
        RECT 3.485 11.970 3.655 12.140 ;
        RECT 4.445 11.970 4.615 12.140 ;
        RECT 5.405 11.970 5.575 12.140 ;
        RECT 6.365 11.970 6.535 12.140 ;
        RECT 1.565 5.535 1.735 5.705 ;
        RECT 2.525 5.535 2.695 5.705 ;
        RECT 3.485 5.535 3.655 5.705 ;
        RECT 4.445 5.535 4.615 5.705 ;
        RECT 5.405 5.535 5.575 5.705 ;
        RECT 6.365 5.535 6.535 5.705 ;
      LAYER met1 ;
        RECT 1.470 204.980 1.830 205.240 ;
        RECT 2.435 204.980 2.795 205.240 ;
        RECT 3.390 204.980 3.750 205.240 ;
        RECT 4.350 204.980 4.710 205.240 ;
        RECT 5.310 204.980 5.670 205.240 ;
        RECT 6.270 204.980 6.630 205.240 ;
        RECT 7.380 204.980 9.300 205.250 ;
        RECT 7.380 204.970 9.260 204.980 ;
        RECT 1.470 198.545 1.830 198.805 ;
        RECT 2.435 198.545 2.795 198.805 ;
        RECT 3.390 198.545 3.750 198.805 ;
        RECT 4.350 198.545 4.710 198.805 ;
        RECT 5.310 198.545 5.670 198.805 ;
        RECT 6.270 198.545 6.630 198.805 ;
        RECT 7.380 198.545 9.300 198.815 ;
        RECT 7.380 198.535 9.260 198.545 ;
        RECT 1.470 192.110 1.830 192.370 ;
        RECT 2.435 192.110 2.795 192.370 ;
        RECT 3.390 192.110 3.750 192.370 ;
        RECT 4.350 192.110 4.710 192.370 ;
        RECT 5.310 192.110 5.670 192.370 ;
        RECT 6.270 192.110 6.630 192.370 ;
        RECT 7.380 192.110 9.300 192.380 ;
        RECT 7.380 192.100 9.260 192.110 ;
        RECT 1.470 185.675 1.830 185.935 ;
        RECT 2.435 185.675 2.795 185.935 ;
        RECT 3.390 185.675 3.750 185.935 ;
        RECT 4.350 185.675 4.710 185.935 ;
        RECT 5.310 185.675 5.670 185.935 ;
        RECT 6.270 185.675 6.630 185.935 ;
        RECT 7.380 185.675 9.300 185.945 ;
        RECT 7.380 185.665 9.260 185.675 ;
        RECT 1.470 179.240 1.830 179.500 ;
        RECT 2.435 179.240 2.795 179.500 ;
        RECT 3.390 179.240 3.750 179.500 ;
        RECT 4.350 179.240 4.710 179.500 ;
        RECT 5.310 179.240 5.670 179.500 ;
        RECT 6.270 179.240 6.630 179.500 ;
        RECT 7.380 179.240 9.300 179.510 ;
        RECT 7.380 179.230 9.260 179.240 ;
        RECT 1.470 172.805 1.830 173.065 ;
        RECT 2.435 172.805 2.795 173.065 ;
        RECT 3.390 172.805 3.750 173.065 ;
        RECT 4.350 172.805 4.710 173.065 ;
        RECT 5.310 172.805 5.670 173.065 ;
        RECT 6.270 172.805 6.630 173.065 ;
        RECT 7.380 172.805 9.300 173.075 ;
        RECT 7.380 172.795 9.260 172.805 ;
        RECT 1.470 166.370 1.830 166.630 ;
        RECT 2.435 166.370 2.795 166.630 ;
        RECT 3.390 166.370 3.750 166.630 ;
        RECT 4.350 166.370 4.710 166.630 ;
        RECT 5.310 166.370 5.670 166.630 ;
        RECT 6.270 166.370 6.630 166.630 ;
        RECT 7.380 166.370 9.300 166.640 ;
        RECT 7.380 166.360 9.260 166.370 ;
        RECT 1.470 159.935 1.830 160.195 ;
        RECT 2.435 159.935 2.795 160.195 ;
        RECT 3.390 159.935 3.750 160.195 ;
        RECT 4.350 159.935 4.710 160.195 ;
        RECT 5.310 159.935 5.670 160.195 ;
        RECT 6.270 159.935 6.630 160.195 ;
        RECT 7.380 159.935 9.300 160.205 ;
        RECT 7.380 159.925 9.260 159.935 ;
        RECT 1.470 153.500 1.830 153.760 ;
        RECT 2.435 153.500 2.795 153.760 ;
        RECT 3.390 153.500 3.750 153.760 ;
        RECT 4.350 153.500 4.710 153.760 ;
        RECT 5.310 153.500 5.670 153.760 ;
        RECT 6.270 153.500 6.630 153.760 ;
        RECT 7.380 153.500 9.300 153.770 ;
        RECT 7.380 153.490 9.260 153.500 ;
        RECT 1.470 147.065 1.830 147.325 ;
        RECT 2.435 147.065 2.795 147.325 ;
        RECT 3.390 147.065 3.750 147.325 ;
        RECT 4.350 147.065 4.710 147.325 ;
        RECT 5.310 147.065 5.670 147.325 ;
        RECT 6.270 147.065 6.630 147.325 ;
        RECT 7.380 147.065 9.300 147.335 ;
        RECT 7.380 147.055 9.260 147.065 ;
        RECT 1.470 140.630 1.830 140.890 ;
        RECT 2.435 140.630 2.795 140.890 ;
        RECT 3.390 140.630 3.750 140.890 ;
        RECT 4.350 140.630 4.710 140.890 ;
        RECT 5.310 140.630 5.670 140.890 ;
        RECT 6.270 140.630 6.630 140.890 ;
        RECT 7.380 140.630 9.300 140.900 ;
        RECT 7.380 140.620 9.260 140.630 ;
        RECT 1.470 134.195 1.830 134.455 ;
        RECT 2.435 134.195 2.795 134.455 ;
        RECT 3.390 134.195 3.750 134.455 ;
        RECT 4.350 134.195 4.710 134.455 ;
        RECT 5.310 134.195 5.670 134.455 ;
        RECT 6.270 134.195 6.630 134.455 ;
        RECT 7.380 134.195 9.300 134.465 ;
        RECT 7.380 134.185 9.260 134.195 ;
        RECT 1.470 127.760 1.830 128.020 ;
        RECT 2.435 127.760 2.795 128.020 ;
        RECT 3.390 127.760 3.750 128.020 ;
        RECT 4.350 127.760 4.710 128.020 ;
        RECT 5.310 127.760 5.670 128.020 ;
        RECT 6.270 127.760 6.630 128.020 ;
        RECT 7.380 127.760 9.300 128.030 ;
        RECT 7.380 127.750 9.260 127.760 ;
        RECT 1.470 121.325 1.830 121.585 ;
        RECT 2.435 121.325 2.795 121.585 ;
        RECT 3.390 121.325 3.750 121.585 ;
        RECT 4.350 121.325 4.710 121.585 ;
        RECT 5.310 121.325 5.670 121.585 ;
        RECT 6.270 121.325 6.630 121.585 ;
        RECT 7.380 121.325 9.300 121.595 ;
        RECT 7.380 121.315 9.260 121.325 ;
        RECT 1.470 114.890 1.830 115.150 ;
        RECT 2.435 114.890 2.795 115.150 ;
        RECT 3.390 114.890 3.750 115.150 ;
        RECT 4.350 114.890 4.710 115.150 ;
        RECT 5.310 114.890 5.670 115.150 ;
        RECT 6.270 114.890 6.630 115.150 ;
        RECT 7.380 114.890 9.300 115.160 ;
        RECT 7.380 114.880 9.260 114.890 ;
        RECT 1.470 108.455 1.830 108.715 ;
        RECT 2.435 108.455 2.795 108.715 ;
        RECT 3.390 108.455 3.750 108.715 ;
        RECT 4.350 108.455 4.710 108.715 ;
        RECT 5.310 108.455 5.670 108.715 ;
        RECT 6.270 108.455 6.630 108.715 ;
        RECT 7.380 108.455 9.300 108.725 ;
        RECT 7.380 108.445 9.260 108.455 ;
        RECT 1.470 102.020 1.830 102.280 ;
        RECT 2.435 102.020 2.795 102.280 ;
        RECT 3.390 102.020 3.750 102.280 ;
        RECT 4.350 102.020 4.710 102.280 ;
        RECT 5.310 102.020 5.670 102.280 ;
        RECT 6.270 102.020 6.630 102.280 ;
        RECT 7.380 102.020 9.300 102.290 ;
        RECT 7.380 102.010 9.260 102.020 ;
        RECT 1.470 95.585 1.830 95.845 ;
        RECT 2.435 95.585 2.795 95.845 ;
        RECT 3.390 95.585 3.750 95.845 ;
        RECT 4.350 95.585 4.710 95.845 ;
        RECT 5.310 95.585 5.670 95.845 ;
        RECT 6.270 95.585 6.630 95.845 ;
        RECT 7.380 95.585 9.300 95.855 ;
        RECT 7.380 95.575 9.260 95.585 ;
        RECT 1.470 89.150 1.830 89.410 ;
        RECT 2.435 89.150 2.795 89.410 ;
        RECT 3.390 89.150 3.750 89.410 ;
        RECT 4.350 89.150 4.710 89.410 ;
        RECT 5.310 89.150 5.670 89.410 ;
        RECT 6.270 89.150 6.630 89.410 ;
        RECT 7.380 89.150 9.300 89.420 ;
        RECT 7.380 89.140 9.260 89.150 ;
        RECT 1.470 82.715 1.830 82.975 ;
        RECT 2.435 82.715 2.795 82.975 ;
        RECT 3.390 82.715 3.750 82.975 ;
        RECT 4.350 82.715 4.710 82.975 ;
        RECT 5.310 82.715 5.670 82.975 ;
        RECT 6.270 82.715 6.630 82.975 ;
        RECT 7.380 82.715 9.300 82.985 ;
        RECT 7.380 82.705 9.260 82.715 ;
        RECT 1.470 76.280 1.830 76.540 ;
        RECT 2.435 76.280 2.795 76.540 ;
        RECT 3.390 76.280 3.750 76.540 ;
        RECT 4.350 76.280 4.710 76.540 ;
        RECT 5.310 76.280 5.670 76.540 ;
        RECT 6.270 76.280 6.630 76.540 ;
        RECT 7.380 76.280 9.300 76.550 ;
        RECT 7.380 76.270 9.260 76.280 ;
        RECT 1.470 69.845 1.830 70.105 ;
        RECT 2.435 69.845 2.795 70.105 ;
        RECT 3.390 69.845 3.750 70.105 ;
        RECT 4.350 69.845 4.710 70.105 ;
        RECT 5.310 69.845 5.670 70.105 ;
        RECT 6.270 69.845 6.630 70.105 ;
        RECT 7.380 69.845 9.300 70.115 ;
        RECT 7.380 69.835 9.260 69.845 ;
        RECT 1.470 63.410 1.830 63.670 ;
        RECT 2.435 63.410 2.795 63.670 ;
        RECT 3.390 63.410 3.750 63.670 ;
        RECT 4.350 63.410 4.710 63.670 ;
        RECT 5.310 63.410 5.670 63.670 ;
        RECT 6.270 63.410 6.630 63.670 ;
        RECT 7.380 63.410 9.300 63.680 ;
        RECT 7.380 63.400 9.260 63.410 ;
        RECT 1.470 56.975 1.830 57.235 ;
        RECT 2.435 56.975 2.795 57.235 ;
        RECT 3.390 56.975 3.750 57.235 ;
        RECT 4.350 56.975 4.710 57.235 ;
        RECT 5.310 56.975 5.670 57.235 ;
        RECT 6.270 56.975 6.630 57.235 ;
        RECT 7.380 56.975 9.300 57.245 ;
        RECT 7.380 56.965 9.260 56.975 ;
        RECT 1.470 50.540 1.830 50.800 ;
        RECT 2.435 50.540 2.795 50.800 ;
        RECT 3.390 50.540 3.750 50.800 ;
        RECT 4.350 50.540 4.710 50.800 ;
        RECT 5.310 50.540 5.670 50.800 ;
        RECT 6.270 50.540 6.630 50.800 ;
        RECT 7.380 50.540 9.300 50.810 ;
        RECT 7.380 50.530 9.260 50.540 ;
        RECT 1.470 44.105 1.830 44.365 ;
        RECT 2.435 44.105 2.795 44.365 ;
        RECT 3.390 44.105 3.750 44.365 ;
        RECT 4.350 44.105 4.710 44.365 ;
        RECT 5.310 44.105 5.670 44.365 ;
        RECT 6.270 44.105 6.630 44.365 ;
        RECT 7.380 44.105 9.300 44.375 ;
        RECT 7.380 44.095 9.260 44.105 ;
        RECT 1.470 37.670 1.830 37.930 ;
        RECT 2.435 37.670 2.795 37.930 ;
        RECT 3.390 37.670 3.750 37.930 ;
        RECT 4.350 37.670 4.710 37.930 ;
        RECT 5.310 37.670 5.670 37.930 ;
        RECT 6.270 37.670 6.630 37.930 ;
        RECT 7.380 37.670 9.300 37.940 ;
        RECT 7.380 37.660 9.260 37.670 ;
        RECT 1.470 31.235 1.830 31.495 ;
        RECT 2.435 31.235 2.795 31.495 ;
        RECT 3.390 31.235 3.750 31.495 ;
        RECT 4.350 31.235 4.710 31.495 ;
        RECT 5.310 31.235 5.670 31.495 ;
        RECT 6.270 31.235 6.630 31.495 ;
        RECT 7.380 31.235 9.300 31.505 ;
        RECT 7.380 31.225 9.260 31.235 ;
        RECT 1.470 24.800 1.830 25.060 ;
        RECT 2.435 24.800 2.795 25.060 ;
        RECT 3.390 24.800 3.750 25.060 ;
        RECT 4.350 24.800 4.710 25.060 ;
        RECT 5.310 24.800 5.670 25.060 ;
        RECT 6.270 24.800 6.630 25.060 ;
        RECT 7.380 24.800 9.300 25.070 ;
        RECT 7.380 24.790 9.260 24.800 ;
        RECT 1.470 18.365 1.830 18.625 ;
        RECT 2.435 18.365 2.795 18.625 ;
        RECT 3.390 18.365 3.750 18.625 ;
        RECT 4.350 18.365 4.710 18.625 ;
        RECT 5.310 18.365 5.670 18.625 ;
        RECT 6.270 18.365 6.630 18.625 ;
        RECT 7.380 18.365 9.300 18.635 ;
        RECT 7.380 18.355 9.260 18.365 ;
        RECT 1.470 11.930 1.830 12.190 ;
        RECT 2.435 11.930 2.795 12.190 ;
        RECT 3.390 11.930 3.750 12.190 ;
        RECT 4.350 11.930 4.710 12.190 ;
        RECT 5.310 11.930 5.670 12.190 ;
        RECT 6.270 11.930 6.630 12.190 ;
        RECT 7.380 11.930 9.300 12.200 ;
        RECT 7.380 11.920 9.260 11.930 ;
        RECT 1.470 5.495 1.830 5.755 ;
        RECT 2.435 5.495 2.795 5.755 ;
        RECT 3.390 5.495 3.750 5.755 ;
        RECT 4.350 5.495 4.710 5.755 ;
        RECT 5.310 5.495 5.670 5.755 ;
        RECT 6.270 5.495 6.630 5.755 ;
        RECT 7.380 5.495 9.300 5.765 ;
        RECT 7.380 5.485 9.260 5.495 ;
      LAYER via ;
        RECT 1.520 204.980 1.780 205.240 ;
        RECT 2.485 204.980 2.745 205.240 ;
        RECT 3.440 204.980 3.700 205.240 ;
        RECT 4.400 204.980 4.660 205.240 ;
        RECT 5.360 204.980 5.620 205.240 ;
        RECT 6.320 204.980 6.580 205.240 ;
        RECT 7.430 204.970 7.690 205.250 ;
        RECT 8.960 204.980 9.250 205.250 ;
        RECT 1.520 198.545 1.780 198.805 ;
        RECT 2.485 198.545 2.745 198.805 ;
        RECT 3.440 198.545 3.700 198.805 ;
        RECT 4.400 198.545 4.660 198.805 ;
        RECT 5.360 198.545 5.620 198.805 ;
        RECT 6.320 198.545 6.580 198.805 ;
        RECT 7.430 198.535 7.690 198.815 ;
        RECT 8.960 198.545 9.250 198.815 ;
        RECT 1.520 192.110 1.780 192.370 ;
        RECT 2.485 192.110 2.745 192.370 ;
        RECT 3.440 192.110 3.700 192.370 ;
        RECT 4.400 192.110 4.660 192.370 ;
        RECT 5.360 192.110 5.620 192.370 ;
        RECT 6.320 192.110 6.580 192.370 ;
        RECT 7.430 192.100 7.690 192.380 ;
        RECT 8.960 192.110 9.250 192.380 ;
        RECT 1.520 185.675 1.780 185.935 ;
        RECT 2.485 185.675 2.745 185.935 ;
        RECT 3.440 185.675 3.700 185.935 ;
        RECT 4.400 185.675 4.660 185.935 ;
        RECT 5.360 185.675 5.620 185.935 ;
        RECT 6.320 185.675 6.580 185.935 ;
        RECT 7.430 185.665 7.690 185.945 ;
        RECT 8.960 185.675 9.250 185.945 ;
        RECT 1.520 179.240 1.780 179.500 ;
        RECT 2.485 179.240 2.745 179.500 ;
        RECT 3.440 179.240 3.700 179.500 ;
        RECT 4.400 179.240 4.660 179.500 ;
        RECT 5.360 179.240 5.620 179.500 ;
        RECT 6.320 179.240 6.580 179.500 ;
        RECT 7.430 179.230 7.690 179.510 ;
        RECT 8.960 179.240 9.250 179.510 ;
        RECT 1.520 172.805 1.780 173.065 ;
        RECT 2.485 172.805 2.745 173.065 ;
        RECT 3.440 172.805 3.700 173.065 ;
        RECT 4.400 172.805 4.660 173.065 ;
        RECT 5.360 172.805 5.620 173.065 ;
        RECT 6.320 172.805 6.580 173.065 ;
        RECT 7.430 172.795 7.690 173.075 ;
        RECT 8.960 172.805 9.250 173.075 ;
        RECT 1.520 166.370 1.780 166.630 ;
        RECT 2.485 166.370 2.745 166.630 ;
        RECT 3.440 166.370 3.700 166.630 ;
        RECT 4.400 166.370 4.660 166.630 ;
        RECT 5.360 166.370 5.620 166.630 ;
        RECT 6.320 166.370 6.580 166.630 ;
        RECT 7.430 166.360 7.690 166.640 ;
        RECT 8.960 166.370 9.250 166.640 ;
        RECT 1.520 159.935 1.780 160.195 ;
        RECT 2.485 159.935 2.745 160.195 ;
        RECT 3.440 159.935 3.700 160.195 ;
        RECT 4.400 159.935 4.660 160.195 ;
        RECT 5.360 159.935 5.620 160.195 ;
        RECT 6.320 159.935 6.580 160.195 ;
        RECT 7.430 159.925 7.690 160.205 ;
        RECT 8.960 159.935 9.250 160.205 ;
        RECT 1.520 153.500 1.780 153.760 ;
        RECT 2.485 153.500 2.745 153.760 ;
        RECT 3.440 153.500 3.700 153.760 ;
        RECT 4.400 153.500 4.660 153.760 ;
        RECT 5.360 153.500 5.620 153.760 ;
        RECT 6.320 153.500 6.580 153.760 ;
        RECT 7.430 153.490 7.690 153.770 ;
        RECT 8.960 153.500 9.250 153.770 ;
        RECT 1.520 147.065 1.780 147.325 ;
        RECT 2.485 147.065 2.745 147.325 ;
        RECT 3.440 147.065 3.700 147.325 ;
        RECT 4.400 147.065 4.660 147.325 ;
        RECT 5.360 147.065 5.620 147.325 ;
        RECT 6.320 147.065 6.580 147.325 ;
        RECT 7.430 147.055 7.690 147.335 ;
        RECT 8.960 147.065 9.250 147.335 ;
        RECT 1.520 140.630 1.780 140.890 ;
        RECT 2.485 140.630 2.745 140.890 ;
        RECT 3.440 140.630 3.700 140.890 ;
        RECT 4.400 140.630 4.660 140.890 ;
        RECT 5.360 140.630 5.620 140.890 ;
        RECT 6.320 140.630 6.580 140.890 ;
        RECT 7.430 140.620 7.690 140.900 ;
        RECT 8.960 140.630 9.250 140.900 ;
        RECT 1.520 134.195 1.780 134.455 ;
        RECT 2.485 134.195 2.745 134.455 ;
        RECT 3.440 134.195 3.700 134.455 ;
        RECT 4.400 134.195 4.660 134.455 ;
        RECT 5.360 134.195 5.620 134.455 ;
        RECT 6.320 134.195 6.580 134.455 ;
        RECT 7.430 134.185 7.690 134.465 ;
        RECT 8.960 134.195 9.250 134.465 ;
        RECT 1.520 127.760 1.780 128.020 ;
        RECT 2.485 127.760 2.745 128.020 ;
        RECT 3.440 127.760 3.700 128.020 ;
        RECT 4.400 127.760 4.660 128.020 ;
        RECT 5.360 127.760 5.620 128.020 ;
        RECT 6.320 127.760 6.580 128.020 ;
        RECT 7.430 127.750 7.690 128.030 ;
        RECT 8.960 127.760 9.250 128.030 ;
        RECT 1.520 121.325 1.780 121.585 ;
        RECT 2.485 121.325 2.745 121.585 ;
        RECT 3.440 121.325 3.700 121.585 ;
        RECT 4.400 121.325 4.660 121.585 ;
        RECT 5.360 121.325 5.620 121.585 ;
        RECT 6.320 121.325 6.580 121.585 ;
        RECT 7.430 121.315 7.690 121.595 ;
        RECT 8.960 121.325 9.250 121.595 ;
        RECT 1.520 114.890 1.780 115.150 ;
        RECT 2.485 114.890 2.745 115.150 ;
        RECT 3.440 114.890 3.700 115.150 ;
        RECT 4.400 114.890 4.660 115.150 ;
        RECT 5.360 114.890 5.620 115.150 ;
        RECT 6.320 114.890 6.580 115.150 ;
        RECT 7.430 114.880 7.690 115.160 ;
        RECT 8.960 114.890 9.250 115.160 ;
        RECT 1.520 108.455 1.780 108.715 ;
        RECT 2.485 108.455 2.745 108.715 ;
        RECT 3.440 108.455 3.700 108.715 ;
        RECT 4.400 108.455 4.660 108.715 ;
        RECT 5.360 108.455 5.620 108.715 ;
        RECT 6.320 108.455 6.580 108.715 ;
        RECT 7.430 108.445 7.690 108.725 ;
        RECT 8.960 108.455 9.250 108.725 ;
        RECT 1.520 102.020 1.780 102.280 ;
        RECT 2.485 102.020 2.745 102.280 ;
        RECT 3.440 102.020 3.700 102.280 ;
        RECT 4.400 102.020 4.660 102.280 ;
        RECT 5.360 102.020 5.620 102.280 ;
        RECT 6.320 102.020 6.580 102.280 ;
        RECT 7.430 102.010 7.690 102.290 ;
        RECT 8.960 102.020 9.250 102.290 ;
        RECT 1.520 95.585 1.780 95.845 ;
        RECT 2.485 95.585 2.745 95.845 ;
        RECT 3.440 95.585 3.700 95.845 ;
        RECT 4.400 95.585 4.660 95.845 ;
        RECT 5.360 95.585 5.620 95.845 ;
        RECT 6.320 95.585 6.580 95.845 ;
        RECT 7.430 95.575 7.690 95.855 ;
        RECT 8.960 95.585 9.250 95.855 ;
        RECT 1.520 89.150 1.780 89.410 ;
        RECT 2.485 89.150 2.745 89.410 ;
        RECT 3.440 89.150 3.700 89.410 ;
        RECT 4.400 89.150 4.660 89.410 ;
        RECT 5.360 89.150 5.620 89.410 ;
        RECT 6.320 89.150 6.580 89.410 ;
        RECT 7.430 89.140 7.690 89.420 ;
        RECT 8.960 89.150 9.250 89.420 ;
        RECT 1.520 82.715 1.780 82.975 ;
        RECT 2.485 82.715 2.745 82.975 ;
        RECT 3.440 82.715 3.700 82.975 ;
        RECT 4.400 82.715 4.660 82.975 ;
        RECT 5.360 82.715 5.620 82.975 ;
        RECT 6.320 82.715 6.580 82.975 ;
        RECT 7.430 82.705 7.690 82.985 ;
        RECT 8.960 82.715 9.250 82.985 ;
        RECT 1.520 76.280 1.780 76.540 ;
        RECT 2.485 76.280 2.745 76.540 ;
        RECT 3.440 76.280 3.700 76.540 ;
        RECT 4.400 76.280 4.660 76.540 ;
        RECT 5.360 76.280 5.620 76.540 ;
        RECT 6.320 76.280 6.580 76.540 ;
        RECT 7.430 76.270 7.690 76.550 ;
        RECT 8.960 76.280 9.250 76.550 ;
        RECT 1.520 69.845 1.780 70.105 ;
        RECT 2.485 69.845 2.745 70.105 ;
        RECT 3.440 69.845 3.700 70.105 ;
        RECT 4.400 69.845 4.660 70.105 ;
        RECT 5.360 69.845 5.620 70.105 ;
        RECT 6.320 69.845 6.580 70.105 ;
        RECT 7.430 69.835 7.690 70.115 ;
        RECT 8.960 69.845 9.250 70.115 ;
        RECT 1.520 63.410 1.780 63.670 ;
        RECT 2.485 63.410 2.745 63.670 ;
        RECT 3.440 63.410 3.700 63.670 ;
        RECT 4.400 63.410 4.660 63.670 ;
        RECT 5.360 63.410 5.620 63.670 ;
        RECT 6.320 63.410 6.580 63.670 ;
        RECT 7.430 63.400 7.690 63.680 ;
        RECT 8.960 63.410 9.250 63.680 ;
        RECT 1.520 56.975 1.780 57.235 ;
        RECT 2.485 56.975 2.745 57.235 ;
        RECT 3.440 56.975 3.700 57.235 ;
        RECT 4.400 56.975 4.660 57.235 ;
        RECT 5.360 56.975 5.620 57.235 ;
        RECT 6.320 56.975 6.580 57.235 ;
        RECT 7.430 56.965 7.690 57.245 ;
        RECT 8.960 56.975 9.250 57.245 ;
        RECT 1.520 50.540 1.780 50.800 ;
        RECT 2.485 50.540 2.745 50.800 ;
        RECT 3.440 50.540 3.700 50.800 ;
        RECT 4.400 50.540 4.660 50.800 ;
        RECT 5.360 50.540 5.620 50.800 ;
        RECT 6.320 50.540 6.580 50.800 ;
        RECT 7.430 50.530 7.690 50.810 ;
        RECT 8.960 50.540 9.250 50.810 ;
        RECT 1.520 44.105 1.780 44.365 ;
        RECT 2.485 44.105 2.745 44.365 ;
        RECT 3.440 44.105 3.700 44.365 ;
        RECT 4.400 44.105 4.660 44.365 ;
        RECT 5.360 44.105 5.620 44.365 ;
        RECT 6.320 44.105 6.580 44.365 ;
        RECT 7.430 44.095 7.690 44.375 ;
        RECT 8.960 44.105 9.250 44.375 ;
        RECT 1.520 37.670 1.780 37.930 ;
        RECT 2.485 37.670 2.745 37.930 ;
        RECT 3.440 37.670 3.700 37.930 ;
        RECT 4.400 37.670 4.660 37.930 ;
        RECT 5.360 37.670 5.620 37.930 ;
        RECT 6.320 37.670 6.580 37.930 ;
        RECT 7.430 37.660 7.690 37.940 ;
        RECT 8.960 37.670 9.250 37.940 ;
        RECT 1.520 31.235 1.780 31.495 ;
        RECT 2.485 31.235 2.745 31.495 ;
        RECT 3.440 31.235 3.700 31.495 ;
        RECT 4.400 31.235 4.660 31.495 ;
        RECT 5.360 31.235 5.620 31.495 ;
        RECT 6.320 31.235 6.580 31.495 ;
        RECT 7.430 31.225 7.690 31.505 ;
        RECT 8.960 31.235 9.250 31.505 ;
        RECT 1.520 24.800 1.780 25.060 ;
        RECT 2.485 24.800 2.745 25.060 ;
        RECT 3.440 24.800 3.700 25.060 ;
        RECT 4.400 24.800 4.660 25.060 ;
        RECT 5.360 24.800 5.620 25.060 ;
        RECT 6.320 24.800 6.580 25.060 ;
        RECT 7.430 24.790 7.690 25.070 ;
        RECT 8.960 24.800 9.250 25.070 ;
        RECT 1.520 18.365 1.780 18.625 ;
        RECT 2.485 18.365 2.745 18.625 ;
        RECT 3.440 18.365 3.700 18.625 ;
        RECT 4.400 18.365 4.660 18.625 ;
        RECT 5.360 18.365 5.620 18.625 ;
        RECT 6.320 18.365 6.580 18.625 ;
        RECT 7.430 18.355 7.690 18.635 ;
        RECT 8.960 18.365 9.250 18.635 ;
        RECT 1.520 11.930 1.780 12.190 ;
        RECT 2.485 11.930 2.745 12.190 ;
        RECT 3.440 11.930 3.700 12.190 ;
        RECT 4.400 11.930 4.660 12.190 ;
        RECT 5.360 11.930 5.620 12.190 ;
        RECT 6.320 11.930 6.580 12.190 ;
        RECT 7.430 11.920 7.690 12.200 ;
        RECT 8.960 11.930 9.250 12.200 ;
        RECT 1.520 5.495 1.780 5.755 ;
        RECT 2.485 5.495 2.745 5.755 ;
        RECT 3.440 5.495 3.700 5.755 ;
        RECT 4.400 5.495 4.660 5.755 ;
        RECT 5.360 5.495 5.620 5.755 ;
        RECT 6.320 5.495 6.580 5.755 ;
        RECT 7.430 5.485 7.690 5.765 ;
        RECT 8.960 5.495 9.250 5.765 ;
      LAYER met2 ;
        RECT 1.520 205.240 1.780 205.290 ;
        RECT 2.485 205.240 2.745 205.290 ;
        RECT 3.440 205.240 3.700 205.290 ;
        RECT 4.400 205.240 4.660 205.290 ;
        RECT 5.360 205.240 5.620 205.290 ;
        RECT 6.320 205.240 6.580 205.290 ;
        RECT 7.430 205.240 7.690 205.300 ;
        RECT 0.400 204.980 7.870 205.240 ;
        RECT 1.520 204.930 1.780 204.980 ;
        RECT 2.485 204.930 2.745 204.980 ;
        RECT 3.440 204.930 3.700 204.980 ;
        RECT 4.400 204.930 4.660 204.980 ;
        RECT 5.360 204.930 5.620 204.980 ;
        RECT 6.320 204.930 6.580 204.980 ;
        RECT 7.430 204.920 7.690 204.980 ;
        RECT 1.520 198.805 1.780 198.855 ;
        RECT 2.485 198.805 2.745 198.855 ;
        RECT 3.440 198.805 3.700 198.855 ;
        RECT 4.400 198.805 4.660 198.855 ;
        RECT 5.360 198.805 5.620 198.855 ;
        RECT 6.320 198.805 6.580 198.855 ;
        RECT 7.430 198.805 7.690 198.865 ;
        RECT 0.400 198.545 7.870 198.805 ;
        RECT 1.520 198.495 1.780 198.545 ;
        RECT 2.485 198.495 2.745 198.545 ;
        RECT 3.440 198.495 3.700 198.545 ;
        RECT 4.400 198.495 4.660 198.545 ;
        RECT 5.360 198.495 5.620 198.545 ;
        RECT 6.320 198.495 6.580 198.545 ;
        RECT 7.430 198.485 7.690 198.545 ;
        RECT 1.520 192.370 1.780 192.420 ;
        RECT 2.485 192.370 2.745 192.420 ;
        RECT 3.440 192.370 3.700 192.420 ;
        RECT 4.400 192.370 4.660 192.420 ;
        RECT 5.360 192.370 5.620 192.420 ;
        RECT 6.320 192.370 6.580 192.420 ;
        RECT 7.430 192.370 7.690 192.430 ;
        RECT 0.400 192.110 7.870 192.370 ;
        RECT 1.520 192.060 1.780 192.110 ;
        RECT 2.485 192.060 2.745 192.110 ;
        RECT 3.440 192.060 3.700 192.110 ;
        RECT 4.400 192.060 4.660 192.110 ;
        RECT 5.360 192.060 5.620 192.110 ;
        RECT 6.320 192.060 6.580 192.110 ;
        RECT 7.430 192.050 7.690 192.110 ;
        RECT 1.520 185.935 1.780 185.985 ;
        RECT 2.485 185.935 2.745 185.985 ;
        RECT 3.440 185.935 3.700 185.985 ;
        RECT 4.400 185.935 4.660 185.985 ;
        RECT 5.360 185.935 5.620 185.985 ;
        RECT 6.320 185.935 6.580 185.985 ;
        RECT 7.430 185.935 7.690 185.995 ;
        RECT 0.400 185.675 7.870 185.935 ;
        RECT 1.520 185.625 1.780 185.675 ;
        RECT 2.485 185.625 2.745 185.675 ;
        RECT 3.440 185.625 3.700 185.675 ;
        RECT 4.400 185.625 4.660 185.675 ;
        RECT 5.360 185.625 5.620 185.675 ;
        RECT 6.320 185.625 6.580 185.675 ;
        RECT 7.430 185.615 7.690 185.675 ;
        RECT 1.520 179.500 1.780 179.550 ;
        RECT 2.485 179.500 2.745 179.550 ;
        RECT 3.440 179.500 3.700 179.550 ;
        RECT 4.400 179.500 4.660 179.550 ;
        RECT 5.360 179.500 5.620 179.550 ;
        RECT 6.320 179.500 6.580 179.550 ;
        RECT 7.430 179.500 7.690 179.560 ;
        RECT 0.400 179.240 7.870 179.500 ;
        RECT 1.520 179.190 1.780 179.240 ;
        RECT 2.485 179.190 2.745 179.240 ;
        RECT 3.440 179.190 3.700 179.240 ;
        RECT 4.400 179.190 4.660 179.240 ;
        RECT 5.360 179.190 5.620 179.240 ;
        RECT 6.320 179.190 6.580 179.240 ;
        RECT 7.430 179.180 7.690 179.240 ;
        RECT 1.520 173.065 1.780 173.115 ;
        RECT 2.485 173.065 2.745 173.115 ;
        RECT 3.440 173.065 3.700 173.115 ;
        RECT 4.400 173.065 4.660 173.115 ;
        RECT 5.360 173.065 5.620 173.115 ;
        RECT 6.320 173.065 6.580 173.115 ;
        RECT 7.430 173.065 7.690 173.125 ;
        RECT 0.400 172.805 7.870 173.065 ;
        RECT 1.520 172.755 1.780 172.805 ;
        RECT 2.485 172.755 2.745 172.805 ;
        RECT 3.440 172.755 3.700 172.805 ;
        RECT 4.400 172.755 4.660 172.805 ;
        RECT 5.360 172.755 5.620 172.805 ;
        RECT 6.320 172.755 6.580 172.805 ;
        RECT 7.430 172.745 7.690 172.805 ;
        RECT 1.520 166.630 1.780 166.680 ;
        RECT 2.485 166.630 2.745 166.680 ;
        RECT 3.440 166.630 3.700 166.680 ;
        RECT 4.400 166.630 4.660 166.680 ;
        RECT 5.360 166.630 5.620 166.680 ;
        RECT 6.320 166.630 6.580 166.680 ;
        RECT 7.430 166.630 7.690 166.690 ;
        RECT 0.400 166.370 7.870 166.630 ;
        RECT 1.520 166.320 1.780 166.370 ;
        RECT 2.485 166.320 2.745 166.370 ;
        RECT 3.440 166.320 3.700 166.370 ;
        RECT 4.400 166.320 4.660 166.370 ;
        RECT 5.360 166.320 5.620 166.370 ;
        RECT 6.320 166.320 6.580 166.370 ;
        RECT 7.430 166.310 7.690 166.370 ;
        RECT 1.520 160.195 1.780 160.245 ;
        RECT 2.485 160.195 2.745 160.245 ;
        RECT 3.440 160.195 3.700 160.245 ;
        RECT 4.400 160.195 4.660 160.245 ;
        RECT 5.360 160.195 5.620 160.245 ;
        RECT 6.320 160.195 6.580 160.245 ;
        RECT 7.430 160.195 7.690 160.255 ;
        RECT 0.400 159.935 7.870 160.195 ;
        RECT 1.520 159.885 1.780 159.935 ;
        RECT 2.485 159.885 2.745 159.935 ;
        RECT 3.440 159.885 3.700 159.935 ;
        RECT 4.400 159.885 4.660 159.935 ;
        RECT 5.360 159.885 5.620 159.935 ;
        RECT 6.320 159.885 6.580 159.935 ;
        RECT 7.430 159.875 7.690 159.935 ;
        RECT 1.520 153.760 1.780 153.810 ;
        RECT 2.485 153.760 2.745 153.810 ;
        RECT 3.440 153.760 3.700 153.810 ;
        RECT 4.400 153.760 4.660 153.810 ;
        RECT 5.360 153.760 5.620 153.810 ;
        RECT 6.320 153.760 6.580 153.810 ;
        RECT 7.430 153.760 7.690 153.820 ;
        RECT 0.400 153.500 7.870 153.760 ;
        RECT 1.520 153.450 1.780 153.500 ;
        RECT 2.485 153.450 2.745 153.500 ;
        RECT 3.440 153.450 3.700 153.500 ;
        RECT 4.400 153.450 4.660 153.500 ;
        RECT 5.360 153.450 5.620 153.500 ;
        RECT 6.320 153.450 6.580 153.500 ;
        RECT 7.430 153.440 7.690 153.500 ;
        RECT 1.520 147.325 1.780 147.375 ;
        RECT 2.485 147.325 2.745 147.375 ;
        RECT 3.440 147.325 3.700 147.375 ;
        RECT 4.400 147.325 4.660 147.375 ;
        RECT 5.360 147.325 5.620 147.375 ;
        RECT 6.320 147.325 6.580 147.375 ;
        RECT 7.430 147.325 7.690 147.385 ;
        RECT 0.400 147.065 7.870 147.325 ;
        RECT 1.520 147.015 1.780 147.065 ;
        RECT 2.485 147.015 2.745 147.065 ;
        RECT 3.440 147.015 3.700 147.065 ;
        RECT 4.400 147.015 4.660 147.065 ;
        RECT 5.360 147.015 5.620 147.065 ;
        RECT 6.320 147.015 6.580 147.065 ;
        RECT 7.430 147.005 7.690 147.065 ;
        RECT 1.520 140.890 1.780 140.940 ;
        RECT 2.485 140.890 2.745 140.940 ;
        RECT 3.440 140.890 3.700 140.940 ;
        RECT 4.400 140.890 4.660 140.940 ;
        RECT 5.360 140.890 5.620 140.940 ;
        RECT 6.320 140.890 6.580 140.940 ;
        RECT 7.430 140.890 7.690 140.950 ;
        RECT 0.400 140.630 7.870 140.890 ;
        RECT 1.520 140.580 1.780 140.630 ;
        RECT 2.485 140.580 2.745 140.630 ;
        RECT 3.440 140.580 3.700 140.630 ;
        RECT 4.400 140.580 4.660 140.630 ;
        RECT 5.360 140.580 5.620 140.630 ;
        RECT 6.320 140.580 6.580 140.630 ;
        RECT 7.430 140.570 7.690 140.630 ;
        RECT 1.520 134.455 1.780 134.505 ;
        RECT 2.485 134.455 2.745 134.505 ;
        RECT 3.440 134.455 3.700 134.505 ;
        RECT 4.400 134.455 4.660 134.505 ;
        RECT 5.360 134.455 5.620 134.505 ;
        RECT 6.320 134.455 6.580 134.505 ;
        RECT 7.430 134.455 7.690 134.515 ;
        RECT 0.400 134.195 7.870 134.455 ;
        RECT 1.520 134.145 1.780 134.195 ;
        RECT 2.485 134.145 2.745 134.195 ;
        RECT 3.440 134.145 3.700 134.195 ;
        RECT 4.400 134.145 4.660 134.195 ;
        RECT 5.360 134.145 5.620 134.195 ;
        RECT 6.320 134.145 6.580 134.195 ;
        RECT 7.430 134.135 7.690 134.195 ;
        RECT 1.520 128.020 1.780 128.070 ;
        RECT 2.485 128.020 2.745 128.070 ;
        RECT 3.440 128.020 3.700 128.070 ;
        RECT 4.400 128.020 4.660 128.070 ;
        RECT 5.360 128.020 5.620 128.070 ;
        RECT 6.320 128.020 6.580 128.070 ;
        RECT 7.430 128.020 7.690 128.080 ;
        RECT 0.400 127.760 7.870 128.020 ;
        RECT 1.520 127.710 1.780 127.760 ;
        RECT 2.485 127.710 2.745 127.760 ;
        RECT 3.440 127.710 3.700 127.760 ;
        RECT 4.400 127.710 4.660 127.760 ;
        RECT 5.360 127.710 5.620 127.760 ;
        RECT 6.320 127.710 6.580 127.760 ;
        RECT 7.430 127.700 7.690 127.760 ;
        RECT 1.520 121.585 1.780 121.635 ;
        RECT 2.485 121.585 2.745 121.635 ;
        RECT 3.440 121.585 3.700 121.635 ;
        RECT 4.400 121.585 4.660 121.635 ;
        RECT 5.360 121.585 5.620 121.635 ;
        RECT 6.320 121.585 6.580 121.635 ;
        RECT 7.430 121.585 7.690 121.645 ;
        RECT 0.400 121.325 7.870 121.585 ;
        RECT 1.520 121.275 1.780 121.325 ;
        RECT 2.485 121.275 2.745 121.325 ;
        RECT 3.440 121.275 3.700 121.325 ;
        RECT 4.400 121.275 4.660 121.325 ;
        RECT 5.360 121.275 5.620 121.325 ;
        RECT 6.320 121.275 6.580 121.325 ;
        RECT 7.430 121.265 7.690 121.325 ;
        RECT 1.520 115.150 1.780 115.200 ;
        RECT 2.485 115.150 2.745 115.200 ;
        RECT 3.440 115.150 3.700 115.200 ;
        RECT 4.400 115.150 4.660 115.200 ;
        RECT 5.360 115.150 5.620 115.200 ;
        RECT 6.320 115.150 6.580 115.200 ;
        RECT 7.430 115.150 7.690 115.210 ;
        RECT 0.400 114.890 7.870 115.150 ;
        RECT 1.520 114.840 1.780 114.890 ;
        RECT 2.485 114.840 2.745 114.890 ;
        RECT 3.440 114.840 3.700 114.890 ;
        RECT 4.400 114.840 4.660 114.890 ;
        RECT 5.360 114.840 5.620 114.890 ;
        RECT 6.320 114.840 6.580 114.890 ;
        RECT 7.430 114.830 7.690 114.890 ;
        RECT 1.520 108.715 1.780 108.765 ;
        RECT 2.485 108.715 2.745 108.765 ;
        RECT 3.440 108.715 3.700 108.765 ;
        RECT 4.400 108.715 4.660 108.765 ;
        RECT 5.360 108.715 5.620 108.765 ;
        RECT 6.320 108.715 6.580 108.765 ;
        RECT 7.430 108.715 7.690 108.775 ;
        RECT 0.400 108.455 7.870 108.715 ;
        RECT 1.520 108.405 1.780 108.455 ;
        RECT 2.485 108.405 2.745 108.455 ;
        RECT 3.440 108.405 3.700 108.455 ;
        RECT 4.400 108.405 4.660 108.455 ;
        RECT 5.360 108.405 5.620 108.455 ;
        RECT 6.320 108.405 6.580 108.455 ;
        RECT 7.430 108.395 7.690 108.455 ;
        RECT 1.520 102.280 1.780 102.330 ;
        RECT 2.485 102.280 2.745 102.330 ;
        RECT 3.440 102.280 3.700 102.330 ;
        RECT 4.400 102.280 4.660 102.330 ;
        RECT 5.360 102.280 5.620 102.330 ;
        RECT 6.320 102.280 6.580 102.330 ;
        RECT 7.430 102.280 7.690 102.340 ;
        RECT 0.400 102.020 7.870 102.280 ;
        RECT 1.520 101.970 1.780 102.020 ;
        RECT 2.485 101.970 2.745 102.020 ;
        RECT 3.440 101.970 3.700 102.020 ;
        RECT 4.400 101.970 4.660 102.020 ;
        RECT 5.360 101.970 5.620 102.020 ;
        RECT 6.320 101.970 6.580 102.020 ;
        RECT 7.430 101.960 7.690 102.020 ;
        RECT 1.520 95.845 1.780 95.895 ;
        RECT 2.485 95.845 2.745 95.895 ;
        RECT 3.440 95.845 3.700 95.895 ;
        RECT 4.400 95.845 4.660 95.895 ;
        RECT 5.360 95.845 5.620 95.895 ;
        RECT 6.320 95.845 6.580 95.895 ;
        RECT 7.430 95.845 7.690 95.905 ;
        RECT 0.400 95.585 7.870 95.845 ;
        RECT 1.520 95.535 1.780 95.585 ;
        RECT 2.485 95.535 2.745 95.585 ;
        RECT 3.440 95.535 3.700 95.585 ;
        RECT 4.400 95.535 4.660 95.585 ;
        RECT 5.360 95.535 5.620 95.585 ;
        RECT 6.320 95.535 6.580 95.585 ;
        RECT 7.430 95.525 7.690 95.585 ;
        RECT 1.520 89.410 1.780 89.460 ;
        RECT 2.485 89.410 2.745 89.460 ;
        RECT 3.440 89.410 3.700 89.460 ;
        RECT 4.400 89.410 4.660 89.460 ;
        RECT 5.360 89.410 5.620 89.460 ;
        RECT 6.320 89.410 6.580 89.460 ;
        RECT 7.430 89.410 7.690 89.470 ;
        RECT 0.400 89.150 7.870 89.410 ;
        RECT 1.520 89.100 1.780 89.150 ;
        RECT 2.485 89.100 2.745 89.150 ;
        RECT 3.440 89.100 3.700 89.150 ;
        RECT 4.400 89.100 4.660 89.150 ;
        RECT 5.360 89.100 5.620 89.150 ;
        RECT 6.320 89.100 6.580 89.150 ;
        RECT 7.430 89.090 7.690 89.150 ;
        RECT 1.520 82.975 1.780 83.025 ;
        RECT 2.485 82.975 2.745 83.025 ;
        RECT 3.440 82.975 3.700 83.025 ;
        RECT 4.400 82.975 4.660 83.025 ;
        RECT 5.360 82.975 5.620 83.025 ;
        RECT 6.320 82.975 6.580 83.025 ;
        RECT 7.430 82.975 7.690 83.035 ;
        RECT 0.400 82.715 7.870 82.975 ;
        RECT 1.520 82.665 1.780 82.715 ;
        RECT 2.485 82.665 2.745 82.715 ;
        RECT 3.440 82.665 3.700 82.715 ;
        RECT 4.400 82.665 4.660 82.715 ;
        RECT 5.360 82.665 5.620 82.715 ;
        RECT 6.320 82.665 6.580 82.715 ;
        RECT 7.430 82.655 7.690 82.715 ;
        RECT 1.520 76.540 1.780 76.590 ;
        RECT 2.485 76.540 2.745 76.590 ;
        RECT 3.440 76.540 3.700 76.590 ;
        RECT 4.400 76.540 4.660 76.590 ;
        RECT 5.360 76.540 5.620 76.590 ;
        RECT 6.320 76.540 6.580 76.590 ;
        RECT 7.430 76.540 7.690 76.600 ;
        RECT 0.400 76.280 7.870 76.540 ;
        RECT 1.520 76.230 1.780 76.280 ;
        RECT 2.485 76.230 2.745 76.280 ;
        RECT 3.440 76.230 3.700 76.280 ;
        RECT 4.400 76.230 4.660 76.280 ;
        RECT 5.360 76.230 5.620 76.280 ;
        RECT 6.320 76.230 6.580 76.280 ;
        RECT 7.430 76.220 7.690 76.280 ;
        RECT 1.520 70.105 1.780 70.155 ;
        RECT 2.485 70.105 2.745 70.155 ;
        RECT 3.440 70.105 3.700 70.155 ;
        RECT 4.400 70.105 4.660 70.155 ;
        RECT 5.360 70.105 5.620 70.155 ;
        RECT 6.320 70.105 6.580 70.155 ;
        RECT 7.430 70.105 7.690 70.165 ;
        RECT 0.400 69.845 7.870 70.105 ;
        RECT 1.520 69.795 1.780 69.845 ;
        RECT 2.485 69.795 2.745 69.845 ;
        RECT 3.440 69.795 3.700 69.845 ;
        RECT 4.400 69.795 4.660 69.845 ;
        RECT 5.360 69.795 5.620 69.845 ;
        RECT 6.320 69.795 6.580 69.845 ;
        RECT 7.430 69.785 7.690 69.845 ;
        RECT 1.520 63.670 1.780 63.720 ;
        RECT 2.485 63.670 2.745 63.720 ;
        RECT 3.440 63.670 3.700 63.720 ;
        RECT 4.400 63.670 4.660 63.720 ;
        RECT 5.360 63.670 5.620 63.720 ;
        RECT 6.320 63.670 6.580 63.720 ;
        RECT 7.430 63.670 7.690 63.730 ;
        RECT 0.400 63.410 7.870 63.670 ;
        RECT 1.520 63.360 1.780 63.410 ;
        RECT 2.485 63.360 2.745 63.410 ;
        RECT 3.440 63.360 3.700 63.410 ;
        RECT 4.400 63.360 4.660 63.410 ;
        RECT 5.360 63.360 5.620 63.410 ;
        RECT 6.320 63.360 6.580 63.410 ;
        RECT 7.430 63.350 7.690 63.410 ;
        RECT 1.520 57.235 1.780 57.285 ;
        RECT 2.485 57.235 2.745 57.285 ;
        RECT 3.440 57.235 3.700 57.285 ;
        RECT 4.400 57.235 4.660 57.285 ;
        RECT 5.360 57.235 5.620 57.285 ;
        RECT 6.320 57.235 6.580 57.285 ;
        RECT 7.430 57.235 7.690 57.295 ;
        RECT 0.400 56.975 7.870 57.235 ;
        RECT 1.520 56.925 1.780 56.975 ;
        RECT 2.485 56.925 2.745 56.975 ;
        RECT 3.440 56.925 3.700 56.975 ;
        RECT 4.400 56.925 4.660 56.975 ;
        RECT 5.360 56.925 5.620 56.975 ;
        RECT 6.320 56.925 6.580 56.975 ;
        RECT 7.430 56.915 7.690 56.975 ;
        RECT 1.520 50.800 1.780 50.850 ;
        RECT 2.485 50.800 2.745 50.850 ;
        RECT 3.440 50.800 3.700 50.850 ;
        RECT 4.400 50.800 4.660 50.850 ;
        RECT 5.360 50.800 5.620 50.850 ;
        RECT 6.320 50.800 6.580 50.850 ;
        RECT 7.430 50.800 7.690 50.860 ;
        RECT 0.400 50.540 7.870 50.800 ;
        RECT 1.520 50.490 1.780 50.540 ;
        RECT 2.485 50.490 2.745 50.540 ;
        RECT 3.440 50.490 3.700 50.540 ;
        RECT 4.400 50.490 4.660 50.540 ;
        RECT 5.360 50.490 5.620 50.540 ;
        RECT 6.320 50.490 6.580 50.540 ;
        RECT 7.430 50.480 7.690 50.540 ;
        RECT 1.520 44.365 1.780 44.415 ;
        RECT 2.485 44.365 2.745 44.415 ;
        RECT 3.440 44.365 3.700 44.415 ;
        RECT 4.400 44.365 4.660 44.415 ;
        RECT 5.360 44.365 5.620 44.415 ;
        RECT 6.320 44.365 6.580 44.415 ;
        RECT 7.430 44.365 7.690 44.425 ;
        RECT 0.400 44.105 7.870 44.365 ;
        RECT 1.520 44.055 1.780 44.105 ;
        RECT 2.485 44.055 2.745 44.105 ;
        RECT 3.440 44.055 3.700 44.105 ;
        RECT 4.400 44.055 4.660 44.105 ;
        RECT 5.360 44.055 5.620 44.105 ;
        RECT 6.320 44.055 6.580 44.105 ;
        RECT 7.430 44.045 7.690 44.105 ;
        RECT 1.520 37.930 1.780 37.980 ;
        RECT 2.485 37.930 2.745 37.980 ;
        RECT 3.440 37.930 3.700 37.980 ;
        RECT 4.400 37.930 4.660 37.980 ;
        RECT 5.360 37.930 5.620 37.980 ;
        RECT 6.320 37.930 6.580 37.980 ;
        RECT 7.430 37.930 7.690 37.990 ;
        RECT 0.400 37.670 7.870 37.930 ;
        RECT 1.520 37.620 1.780 37.670 ;
        RECT 2.485 37.620 2.745 37.670 ;
        RECT 3.440 37.620 3.700 37.670 ;
        RECT 4.400 37.620 4.660 37.670 ;
        RECT 5.360 37.620 5.620 37.670 ;
        RECT 6.320 37.620 6.580 37.670 ;
        RECT 7.430 37.610 7.690 37.670 ;
        RECT 1.520 31.495 1.780 31.545 ;
        RECT 2.485 31.495 2.745 31.545 ;
        RECT 3.440 31.495 3.700 31.545 ;
        RECT 4.400 31.495 4.660 31.545 ;
        RECT 5.360 31.495 5.620 31.545 ;
        RECT 6.320 31.495 6.580 31.545 ;
        RECT 7.430 31.495 7.690 31.555 ;
        RECT 0.400 31.235 7.870 31.495 ;
        RECT 1.520 31.185 1.780 31.235 ;
        RECT 2.485 31.185 2.745 31.235 ;
        RECT 3.440 31.185 3.700 31.235 ;
        RECT 4.400 31.185 4.660 31.235 ;
        RECT 5.360 31.185 5.620 31.235 ;
        RECT 6.320 31.185 6.580 31.235 ;
        RECT 7.430 31.175 7.690 31.235 ;
        RECT 1.520 25.060 1.780 25.110 ;
        RECT 2.485 25.060 2.745 25.110 ;
        RECT 3.440 25.060 3.700 25.110 ;
        RECT 4.400 25.060 4.660 25.110 ;
        RECT 5.360 25.060 5.620 25.110 ;
        RECT 6.320 25.060 6.580 25.110 ;
        RECT 7.430 25.060 7.690 25.120 ;
        RECT 0.400 24.800 7.870 25.060 ;
        RECT 1.520 24.750 1.780 24.800 ;
        RECT 2.485 24.750 2.745 24.800 ;
        RECT 3.440 24.750 3.700 24.800 ;
        RECT 4.400 24.750 4.660 24.800 ;
        RECT 5.360 24.750 5.620 24.800 ;
        RECT 6.320 24.750 6.580 24.800 ;
        RECT 7.430 24.740 7.690 24.800 ;
        RECT 1.520 18.625 1.780 18.675 ;
        RECT 2.485 18.625 2.745 18.675 ;
        RECT 3.440 18.625 3.700 18.675 ;
        RECT 4.400 18.625 4.660 18.675 ;
        RECT 5.360 18.625 5.620 18.675 ;
        RECT 6.320 18.625 6.580 18.675 ;
        RECT 7.430 18.625 7.690 18.685 ;
        RECT 0.400 18.365 7.870 18.625 ;
        RECT 1.520 18.315 1.780 18.365 ;
        RECT 2.485 18.315 2.745 18.365 ;
        RECT 3.440 18.315 3.700 18.365 ;
        RECT 4.400 18.315 4.660 18.365 ;
        RECT 5.360 18.315 5.620 18.365 ;
        RECT 6.320 18.315 6.580 18.365 ;
        RECT 7.430 18.305 7.690 18.365 ;
        RECT 1.520 12.190 1.780 12.240 ;
        RECT 2.485 12.190 2.745 12.240 ;
        RECT 3.440 12.190 3.700 12.240 ;
        RECT 4.400 12.190 4.660 12.240 ;
        RECT 5.360 12.190 5.620 12.240 ;
        RECT 6.320 12.190 6.580 12.240 ;
        RECT 7.430 12.190 7.690 12.250 ;
        RECT 0.400 11.930 7.870 12.190 ;
        RECT 1.520 11.880 1.780 11.930 ;
        RECT 2.485 11.880 2.745 11.930 ;
        RECT 3.440 11.880 3.700 11.930 ;
        RECT 4.400 11.880 4.660 11.930 ;
        RECT 5.360 11.880 5.620 11.930 ;
        RECT 6.320 11.880 6.580 11.930 ;
        RECT 7.430 11.870 7.690 11.930 ;
        RECT 1.520 5.755 1.780 5.805 ;
        RECT 2.485 5.755 2.745 5.805 ;
        RECT 3.440 5.755 3.700 5.805 ;
        RECT 4.400 5.755 4.660 5.805 ;
        RECT 5.360 5.755 5.620 5.805 ;
        RECT 6.320 5.755 6.580 5.805 ;
        RECT 7.430 5.755 7.690 5.815 ;
        RECT 0.400 5.495 7.870 5.755 ;
        RECT 1.520 5.445 1.780 5.495 ;
        RECT 2.485 5.445 2.745 5.495 ;
        RECT 3.440 5.445 3.700 5.495 ;
        RECT 4.400 5.445 4.660 5.495 ;
        RECT 5.360 5.445 5.620 5.495 ;
        RECT 6.320 5.445 6.580 5.495 ;
        RECT 7.430 5.435 7.690 5.495 ;
        RECT 8.960 0.725 9.260 206.760 ;
    END
  END s_en_b
  OBS
      LAYER li ;
        RECT 0.730 1.510 28.680 205.880 ;
      LAYER m1 ;
        RECT 0.730 1.510 28.680 205.880 ;
      LAYER m2 ;
        RECT 0.730 1.510 28.680 205.880 ;
      LAYER m3 ;
        RECT 0.730 1.510 28.680 205.880 ; 
      LAYER li1 ;
        RECT 1.565 203.400 1.735 204.800 ;
        RECT 2.525 203.400 2.695 204.800 ;
        RECT 3.485 203.400 3.655 204.800 ;
        RECT 4.445 203.400 4.615 204.800 ;
        RECT 5.405 203.400 5.575 204.800 ;
        RECT 6.365 203.400 6.535 204.800 ;
        RECT 12.330 203.420 12.500 204.820 ;
        RECT 12.810 203.420 12.980 204.820 ;
        RECT 13.290 203.420 13.460 204.820 ;
        RECT 13.770 203.420 13.940 204.820 ;
        RECT 14.250 203.420 14.420 204.820 ;
        RECT 14.730 203.420 14.900 204.820 ;
        RECT 15.210 203.420 15.380 204.820 ;
        RECT 15.690 203.420 15.860 204.820 ;
        RECT 16.170 203.420 16.340 204.820 ;
        RECT 16.650 203.420 16.820 204.820 ;
        RECT 17.130 203.420 17.300 204.820 ;
        RECT 20.415 203.420 20.585 204.820 ;
        RECT 21.375 203.420 21.545 204.820 ;
        RECT 22.335 203.420 22.505 204.820 ;
        RECT 23.295 203.420 23.465 204.820 ;
        RECT 24.255 203.420 24.425 204.820 ;
        RECT 26.700 202.735 27.030 203.715 ;
        RECT 26.700 202.135 26.930 202.735 ;
        RECT 1.565 201.340 1.735 201.900 ;
        RECT 2.525 201.340 2.695 201.900 ;
        RECT 3.485 201.340 3.655 201.900 ;
        RECT 4.445 201.340 4.615 201.900 ;
        RECT 5.405 201.340 5.575 201.900 ;
        RECT 6.365 201.340 6.535 201.900 ;
        RECT 12.330 201.360 12.500 201.920 ;
        RECT 12.810 201.360 12.980 201.920 ;
        RECT 13.290 201.360 13.460 201.920 ;
        RECT 13.770 201.360 13.940 201.920 ;
        RECT 14.250 201.360 14.420 201.920 ;
        RECT 14.730 201.360 14.900 201.920 ;
        RECT 15.210 201.360 15.380 201.920 ;
        RECT 15.690 201.360 15.860 201.920 ;
        RECT 16.170 201.360 16.340 201.920 ;
        RECT 16.650 201.360 16.820 201.920 ;
        RECT 17.130 201.360 17.300 201.920 ;
        RECT 18.675 201.400 18.845 201.940 ;
        RECT 20.415 201.360 20.585 201.920 ;
        RECT 21.375 201.360 21.545 201.920 ;
        RECT 22.335 201.360 22.505 201.920 ;
        RECT 23.295 201.360 23.465 201.920 ;
        RECT 24.255 201.360 24.425 201.920 ;
        RECT 26.700 201.505 27.030 202.135 ;
        RECT 12.250 201.000 12.580 201.170 ;
        RECT 13.210 201.000 13.540 201.170 ;
        RECT 14.170 201.000 14.500 201.170 ;
        RECT 15.130 201.000 15.460 201.170 ;
        RECT 16.090 201.000 16.420 201.170 ;
        RECT 17.050 201.000 17.380 201.170 ;
        RECT 19.855 201.000 20.185 201.170 ;
        RECT 20.815 201.000 21.145 201.170 ;
        RECT 21.775 201.000 22.105 201.170 ;
        RECT 22.735 201.000 23.065 201.170 ;
        RECT 23.695 201.000 24.025 201.170 ;
        RECT 24.655 201.000 24.985 201.170 ;
        RECT 1.565 196.965 1.735 198.365 ;
        RECT 2.525 196.965 2.695 198.365 ;
        RECT 3.485 196.965 3.655 198.365 ;
        RECT 4.445 196.965 4.615 198.365 ;
        RECT 5.405 196.965 5.575 198.365 ;
        RECT 6.365 196.965 6.535 198.365 ;
        RECT 12.330 196.985 12.500 198.385 ;
        RECT 12.810 196.985 12.980 198.385 ;
        RECT 13.290 196.985 13.460 198.385 ;
        RECT 13.770 196.985 13.940 198.385 ;
        RECT 14.250 196.985 14.420 198.385 ;
        RECT 14.730 196.985 14.900 198.385 ;
        RECT 15.210 196.985 15.380 198.385 ;
        RECT 15.690 196.985 15.860 198.385 ;
        RECT 16.170 196.985 16.340 198.385 ;
        RECT 16.650 196.985 16.820 198.385 ;
        RECT 17.130 196.985 17.300 198.385 ;
        RECT 20.415 196.985 20.585 198.385 ;
        RECT 21.375 196.985 21.545 198.385 ;
        RECT 22.335 196.985 22.505 198.385 ;
        RECT 23.295 196.985 23.465 198.385 ;
        RECT 24.255 196.985 24.425 198.385 ;
        RECT 26.700 196.300 27.030 197.280 ;
        RECT 26.700 195.700 26.930 196.300 ;
        RECT 1.565 194.905 1.735 195.465 ;
        RECT 2.525 194.905 2.695 195.465 ;
        RECT 3.485 194.905 3.655 195.465 ;
        RECT 4.445 194.905 4.615 195.465 ;
        RECT 5.405 194.905 5.575 195.465 ;
        RECT 6.365 194.905 6.535 195.465 ;
        RECT 12.330 194.925 12.500 195.485 ;
        RECT 12.810 194.925 12.980 195.485 ;
        RECT 13.290 194.925 13.460 195.485 ;
        RECT 13.770 194.925 13.940 195.485 ;
        RECT 14.250 194.925 14.420 195.485 ;
        RECT 14.730 194.925 14.900 195.485 ;
        RECT 15.210 194.925 15.380 195.485 ;
        RECT 15.690 194.925 15.860 195.485 ;
        RECT 16.170 194.925 16.340 195.485 ;
        RECT 16.650 194.925 16.820 195.485 ;
        RECT 17.130 194.925 17.300 195.485 ;
        RECT 18.675 194.965 18.845 195.505 ;
        RECT 20.415 194.925 20.585 195.485 ;
        RECT 21.375 194.925 21.545 195.485 ;
        RECT 22.335 194.925 22.505 195.485 ;
        RECT 23.295 194.925 23.465 195.485 ;
        RECT 24.255 194.925 24.425 195.485 ;
        RECT 26.700 195.070 27.030 195.700 ;
        RECT 12.250 194.565 12.580 194.735 ;
        RECT 13.210 194.565 13.540 194.735 ;
        RECT 14.170 194.565 14.500 194.735 ;
        RECT 15.130 194.565 15.460 194.735 ;
        RECT 16.090 194.565 16.420 194.735 ;
        RECT 17.050 194.565 17.380 194.735 ;
        RECT 19.855 194.565 20.185 194.735 ;
        RECT 20.815 194.565 21.145 194.735 ;
        RECT 21.775 194.565 22.105 194.735 ;
        RECT 22.735 194.565 23.065 194.735 ;
        RECT 23.695 194.565 24.025 194.735 ;
        RECT 24.655 194.565 24.985 194.735 ;
        RECT 1.565 190.530 1.735 191.930 ;
        RECT 2.525 190.530 2.695 191.930 ;
        RECT 3.485 190.530 3.655 191.930 ;
        RECT 4.445 190.530 4.615 191.930 ;
        RECT 5.405 190.530 5.575 191.930 ;
        RECT 6.365 190.530 6.535 191.930 ;
        RECT 12.330 190.550 12.500 191.950 ;
        RECT 12.810 190.550 12.980 191.950 ;
        RECT 13.290 190.550 13.460 191.950 ;
        RECT 13.770 190.550 13.940 191.950 ;
        RECT 14.250 190.550 14.420 191.950 ;
        RECT 14.730 190.550 14.900 191.950 ;
        RECT 15.210 190.550 15.380 191.950 ;
        RECT 15.690 190.550 15.860 191.950 ;
        RECT 16.170 190.550 16.340 191.950 ;
        RECT 16.650 190.550 16.820 191.950 ;
        RECT 17.130 190.550 17.300 191.950 ;
        RECT 20.415 190.550 20.585 191.950 ;
        RECT 21.375 190.550 21.545 191.950 ;
        RECT 22.335 190.550 22.505 191.950 ;
        RECT 23.295 190.550 23.465 191.950 ;
        RECT 24.255 190.550 24.425 191.950 ;
        RECT 26.700 189.865 27.030 190.845 ;
        RECT 26.700 189.265 26.930 189.865 ;
        RECT 1.565 188.470 1.735 189.030 ;
        RECT 2.525 188.470 2.695 189.030 ;
        RECT 3.485 188.470 3.655 189.030 ;
        RECT 4.445 188.470 4.615 189.030 ;
        RECT 5.405 188.470 5.575 189.030 ;
        RECT 6.365 188.470 6.535 189.030 ;
        RECT 12.330 188.490 12.500 189.050 ;
        RECT 12.810 188.490 12.980 189.050 ;
        RECT 13.290 188.490 13.460 189.050 ;
        RECT 13.770 188.490 13.940 189.050 ;
        RECT 14.250 188.490 14.420 189.050 ;
        RECT 14.730 188.490 14.900 189.050 ;
        RECT 15.210 188.490 15.380 189.050 ;
        RECT 15.690 188.490 15.860 189.050 ;
        RECT 16.170 188.490 16.340 189.050 ;
        RECT 16.650 188.490 16.820 189.050 ;
        RECT 17.130 188.490 17.300 189.050 ;
        RECT 18.675 188.530 18.845 189.070 ;
        RECT 20.415 188.490 20.585 189.050 ;
        RECT 21.375 188.490 21.545 189.050 ;
        RECT 22.335 188.490 22.505 189.050 ;
        RECT 23.295 188.490 23.465 189.050 ;
        RECT 24.255 188.490 24.425 189.050 ;
        RECT 26.700 188.635 27.030 189.265 ;
        RECT 12.250 188.130 12.580 188.300 ;
        RECT 13.210 188.130 13.540 188.300 ;
        RECT 14.170 188.130 14.500 188.300 ;
        RECT 15.130 188.130 15.460 188.300 ;
        RECT 16.090 188.130 16.420 188.300 ;
        RECT 17.050 188.130 17.380 188.300 ;
        RECT 19.855 188.130 20.185 188.300 ;
        RECT 20.815 188.130 21.145 188.300 ;
        RECT 21.775 188.130 22.105 188.300 ;
        RECT 22.735 188.130 23.065 188.300 ;
        RECT 23.695 188.130 24.025 188.300 ;
        RECT 24.655 188.130 24.985 188.300 ;
        RECT 1.565 184.095 1.735 185.495 ;
        RECT 2.525 184.095 2.695 185.495 ;
        RECT 3.485 184.095 3.655 185.495 ;
        RECT 4.445 184.095 4.615 185.495 ;
        RECT 5.405 184.095 5.575 185.495 ;
        RECT 6.365 184.095 6.535 185.495 ;
        RECT 12.330 184.115 12.500 185.515 ;
        RECT 12.810 184.115 12.980 185.515 ;
        RECT 13.290 184.115 13.460 185.515 ;
        RECT 13.770 184.115 13.940 185.515 ;
        RECT 14.250 184.115 14.420 185.515 ;
        RECT 14.730 184.115 14.900 185.515 ;
        RECT 15.210 184.115 15.380 185.515 ;
        RECT 15.690 184.115 15.860 185.515 ;
        RECT 16.170 184.115 16.340 185.515 ;
        RECT 16.650 184.115 16.820 185.515 ;
        RECT 17.130 184.115 17.300 185.515 ;
        RECT 20.415 184.115 20.585 185.515 ;
        RECT 21.375 184.115 21.545 185.515 ;
        RECT 22.335 184.115 22.505 185.515 ;
        RECT 23.295 184.115 23.465 185.515 ;
        RECT 24.255 184.115 24.425 185.515 ;
        RECT 26.700 183.430 27.030 184.410 ;
        RECT 26.700 182.830 26.930 183.430 ;
        RECT 1.565 182.035 1.735 182.595 ;
        RECT 2.525 182.035 2.695 182.595 ;
        RECT 3.485 182.035 3.655 182.595 ;
        RECT 4.445 182.035 4.615 182.595 ;
        RECT 5.405 182.035 5.575 182.595 ;
        RECT 6.365 182.035 6.535 182.595 ;
        RECT 12.330 182.055 12.500 182.615 ;
        RECT 12.810 182.055 12.980 182.615 ;
        RECT 13.290 182.055 13.460 182.615 ;
        RECT 13.770 182.055 13.940 182.615 ;
        RECT 14.250 182.055 14.420 182.615 ;
        RECT 14.730 182.055 14.900 182.615 ;
        RECT 15.210 182.055 15.380 182.615 ;
        RECT 15.690 182.055 15.860 182.615 ;
        RECT 16.170 182.055 16.340 182.615 ;
        RECT 16.650 182.055 16.820 182.615 ;
        RECT 17.130 182.055 17.300 182.615 ;
        RECT 18.675 182.095 18.845 182.635 ;
        RECT 20.415 182.055 20.585 182.615 ;
        RECT 21.375 182.055 21.545 182.615 ;
        RECT 22.335 182.055 22.505 182.615 ;
        RECT 23.295 182.055 23.465 182.615 ;
        RECT 24.255 182.055 24.425 182.615 ;
        RECT 26.700 182.200 27.030 182.830 ;
        RECT 12.250 181.695 12.580 181.865 ;
        RECT 13.210 181.695 13.540 181.865 ;
        RECT 14.170 181.695 14.500 181.865 ;
        RECT 15.130 181.695 15.460 181.865 ;
        RECT 16.090 181.695 16.420 181.865 ;
        RECT 17.050 181.695 17.380 181.865 ;
        RECT 19.855 181.695 20.185 181.865 ;
        RECT 20.815 181.695 21.145 181.865 ;
        RECT 21.775 181.695 22.105 181.865 ;
        RECT 22.735 181.695 23.065 181.865 ;
        RECT 23.695 181.695 24.025 181.865 ;
        RECT 24.655 181.695 24.985 181.865 ;
        RECT 1.565 177.660 1.735 179.060 ;
        RECT 2.525 177.660 2.695 179.060 ;
        RECT 3.485 177.660 3.655 179.060 ;
        RECT 4.445 177.660 4.615 179.060 ;
        RECT 5.405 177.660 5.575 179.060 ;
        RECT 6.365 177.660 6.535 179.060 ;
        RECT 12.330 177.680 12.500 179.080 ;
        RECT 12.810 177.680 12.980 179.080 ;
        RECT 13.290 177.680 13.460 179.080 ;
        RECT 13.770 177.680 13.940 179.080 ;
        RECT 14.250 177.680 14.420 179.080 ;
        RECT 14.730 177.680 14.900 179.080 ;
        RECT 15.210 177.680 15.380 179.080 ;
        RECT 15.690 177.680 15.860 179.080 ;
        RECT 16.170 177.680 16.340 179.080 ;
        RECT 16.650 177.680 16.820 179.080 ;
        RECT 17.130 177.680 17.300 179.080 ;
        RECT 20.415 177.680 20.585 179.080 ;
        RECT 21.375 177.680 21.545 179.080 ;
        RECT 22.335 177.680 22.505 179.080 ;
        RECT 23.295 177.680 23.465 179.080 ;
        RECT 24.255 177.680 24.425 179.080 ;
        RECT 26.700 176.995 27.030 177.975 ;
        RECT 26.700 176.395 26.930 176.995 ;
        RECT 1.565 175.600 1.735 176.160 ;
        RECT 2.525 175.600 2.695 176.160 ;
        RECT 3.485 175.600 3.655 176.160 ;
        RECT 4.445 175.600 4.615 176.160 ;
        RECT 5.405 175.600 5.575 176.160 ;
        RECT 6.365 175.600 6.535 176.160 ;
        RECT 12.330 175.620 12.500 176.180 ;
        RECT 12.810 175.620 12.980 176.180 ;
        RECT 13.290 175.620 13.460 176.180 ;
        RECT 13.770 175.620 13.940 176.180 ;
        RECT 14.250 175.620 14.420 176.180 ;
        RECT 14.730 175.620 14.900 176.180 ;
        RECT 15.210 175.620 15.380 176.180 ;
        RECT 15.690 175.620 15.860 176.180 ;
        RECT 16.170 175.620 16.340 176.180 ;
        RECT 16.650 175.620 16.820 176.180 ;
        RECT 17.130 175.620 17.300 176.180 ;
        RECT 18.675 175.660 18.845 176.200 ;
        RECT 20.415 175.620 20.585 176.180 ;
        RECT 21.375 175.620 21.545 176.180 ;
        RECT 22.335 175.620 22.505 176.180 ;
        RECT 23.295 175.620 23.465 176.180 ;
        RECT 24.255 175.620 24.425 176.180 ;
        RECT 26.700 175.765 27.030 176.395 ;
        RECT 12.250 175.260 12.580 175.430 ;
        RECT 13.210 175.260 13.540 175.430 ;
        RECT 14.170 175.260 14.500 175.430 ;
        RECT 15.130 175.260 15.460 175.430 ;
        RECT 16.090 175.260 16.420 175.430 ;
        RECT 17.050 175.260 17.380 175.430 ;
        RECT 19.855 175.260 20.185 175.430 ;
        RECT 20.815 175.260 21.145 175.430 ;
        RECT 21.775 175.260 22.105 175.430 ;
        RECT 22.735 175.260 23.065 175.430 ;
        RECT 23.695 175.260 24.025 175.430 ;
        RECT 24.655 175.260 24.985 175.430 ;
        RECT 1.565 171.225 1.735 172.625 ;
        RECT 2.525 171.225 2.695 172.625 ;
        RECT 3.485 171.225 3.655 172.625 ;
        RECT 4.445 171.225 4.615 172.625 ;
        RECT 5.405 171.225 5.575 172.625 ;
        RECT 6.365 171.225 6.535 172.625 ;
        RECT 12.330 171.245 12.500 172.645 ;
        RECT 12.810 171.245 12.980 172.645 ;
        RECT 13.290 171.245 13.460 172.645 ;
        RECT 13.770 171.245 13.940 172.645 ;
        RECT 14.250 171.245 14.420 172.645 ;
        RECT 14.730 171.245 14.900 172.645 ;
        RECT 15.210 171.245 15.380 172.645 ;
        RECT 15.690 171.245 15.860 172.645 ;
        RECT 16.170 171.245 16.340 172.645 ;
        RECT 16.650 171.245 16.820 172.645 ;
        RECT 17.130 171.245 17.300 172.645 ;
        RECT 20.415 171.245 20.585 172.645 ;
        RECT 21.375 171.245 21.545 172.645 ;
        RECT 22.335 171.245 22.505 172.645 ;
        RECT 23.295 171.245 23.465 172.645 ;
        RECT 24.255 171.245 24.425 172.645 ;
        RECT 26.700 170.560 27.030 171.540 ;
        RECT 26.700 169.960 26.930 170.560 ;
        RECT 1.565 169.165 1.735 169.725 ;
        RECT 2.525 169.165 2.695 169.725 ;
        RECT 3.485 169.165 3.655 169.725 ;
        RECT 4.445 169.165 4.615 169.725 ;
        RECT 5.405 169.165 5.575 169.725 ;
        RECT 6.365 169.165 6.535 169.725 ;
        RECT 12.330 169.185 12.500 169.745 ;
        RECT 12.810 169.185 12.980 169.745 ;
        RECT 13.290 169.185 13.460 169.745 ;
        RECT 13.770 169.185 13.940 169.745 ;
        RECT 14.250 169.185 14.420 169.745 ;
        RECT 14.730 169.185 14.900 169.745 ;
        RECT 15.210 169.185 15.380 169.745 ;
        RECT 15.690 169.185 15.860 169.745 ;
        RECT 16.170 169.185 16.340 169.745 ;
        RECT 16.650 169.185 16.820 169.745 ;
        RECT 17.130 169.185 17.300 169.745 ;
        RECT 18.675 169.225 18.845 169.765 ;
        RECT 20.415 169.185 20.585 169.745 ;
        RECT 21.375 169.185 21.545 169.745 ;
        RECT 22.335 169.185 22.505 169.745 ;
        RECT 23.295 169.185 23.465 169.745 ;
        RECT 24.255 169.185 24.425 169.745 ;
        RECT 26.700 169.330 27.030 169.960 ;
        RECT 12.250 168.825 12.580 168.995 ;
        RECT 13.210 168.825 13.540 168.995 ;
        RECT 14.170 168.825 14.500 168.995 ;
        RECT 15.130 168.825 15.460 168.995 ;
        RECT 16.090 168.825 16.420 168.995 ;
        RECT 17.050 168.825 17.380 168.995 ;
        RECT 19.855 168.825 20.185 168.995 ;
        RECT 20.815 168.825 21.145 168.995 ;
        RECT 21.775 168.825 22.105 168.995 ;
        RECT 22.735 168.825 23.065 168.995 ;
        RECT 23.695 168.825 24.025 168.995 ;
        RECT 24.655 168.825 24.985 168.995 ;
        RECT 1.565 164.790 1.735 166.190 ;
        RECT 2.525 164.790 2.695 166.190 ;
        RECT 3.485 164.790 3.655 166.190 ;
        RECT 4.445 164.790 4.615 166.190 ;
        RECT 5.405 164.790 5.575 166.190 ;
        RECT 6.365 164.790 6.535 166.190 ;
        RECT 12.330 164.810 12.500 166.210 ;
        RECT 12.810 164.810 12.980 166.210 ;
        RECT 13.290 164.810 13.460 166.210 ;
        RECT 13.770 164.810 13.940 166.210 ;
        RECT 14.250 164.810 14.420 166.210 ;
        RECT 14.730 164.810 14.900 166.210 ;
        RECT 15.210 164.810 15.380 166.210 ;
        RECT 15.690 164.810 15.860 166.210 ;
        RECT 16.170 164.810 16.340 166.210 ;
        RECT 16.650 164.810 16.820 166.210 ;
        RECT 17.130 164.810 17.300 166.210 ;
        RECT 20.415 164.810 20.585 166.210 ;
        RECT 21.375 164.810 21.545 166.210 ;
        RECT 22.335 164.810 22.505 166.210 ;
        RECT 23.295 164.810 23.465 166.210 ;
        RECT 24.255 164.810 24.425 166.210 ;
        RECT 26.700 164.125 27.030 165.105 ;
        RECT 26.700 163.525 26.930 164.125 ;
        RECT 1.565 162.730 1.735 163.290 ;
        RECT 2.525 162.730 2.695 163.290 ;
        RECT 3.485 162.730 3.655 163.290 ;
        RECT 4.445 162.730 4.615 163.290 ;
        RECT 5.405 162.730 5.575 163.290 ;
        RECT 6.365 162.730 6.535 163.290 ;
        RECT 12.330 162.750 12.500 163.310 ;
        RECT 12.810 162.750 12.980 163.310 ;
        RECT 13.290 162.750 13.460 163.310 ;
        RECT 13.770 162.750 13.940 163.310 ;
        RECT 14.250 162.750 14.420 163.310 ;
        RECT 14.730 162.750 14.900 163.310 ;
        RECT 15.210 162.750 15.380 163.310 ;
        RECT 15.690 162.750 15.860 163.310 ;
        RECT 16.170 162.750 16.340 163.310 ;
        RECT 16.650 162.750 16.820 163.310 ;
        RECT 17.130 162.750 17.300 163.310 ;
        RECT 18.675 162.790 18.845 163.330 ;
        RECT 20.415 162.750 20.585 163.310 ;
        RECT 21.375 162.750 21.545 163.310 ;
        RECT 22.335 162.750 22.505 163.310 ;
        RECT 23.295 162.750 23.465 163.310 ;
        RECT 24.255 162.750 24.425 163.310 ;
        RECT 26.700 162.895 27.030 163.525 ;
        RECT 12.250 162.390 12.580 162.560 ;
        RECT 13.210 162.390 13.540 162.560 ;
        RECT 14.170 162.390 14.500 162.560 ;
        RECT 15.130 162.390 15.460 162.560 ;
        RECT 16.090 162.390 16.420 162.560 ;
        RECT 17.050 162.390 17.380 162.560 ;
        RECT 19.855 162.390 20.185 162.560 ;
        RECT 20.815 162.390 21.145 162.560 ;
        RECT 21.775 162.390 22.105 162.560 ;
        RECT 22.735 162.390 23.065 162.560 ;
        RECT 23.695 162.390 24.025 162.560 ;
        RECT 24.655 162.390 24.985 162.560 ;
        RECT 1.565 158.355 1.735 159.755 ;
        RECT 2.525 158.355 2.695 159.755 ;
        RECT 3.485 158.355 3.655 159.755 ;
        RECT 4.445 158.355 4.615 159.755 ;
        RECT 5.405 158.355 5.575 159.755 ;
        RECT 6.365 158.355 6.535 159.755 ;
        RECT 12.330 158.375 12.500 159.775 ;
        RECT 12.810 158.375 12.980 159.775 ;
        RECT 13.290 158.375 13.460 159.775 ;
        RECT 13.770 158.375 13.940 159.775 ;
        RECT 14.250 158.375 14.420 159.775 ;
        RECT 14.730 158.375 14.900 159.775 ;
        RECT 15.210 158.375 15.380 159.775 ;
        RECT 15.690 158.375 15.860 159.775 ;
        RECT 16.170 158.375 16.340 159.775 ;
        RECT 16.650 158.375 16.820 159.775 ;
        RECT 17.130 158.375 17.300 159.775 ;
        RECT 20.415 158.375 20.585 159.775 ;
        RECT 21.375 158.375 21.545 159.775 ;
        RECT 22.335 158.375 22.505 159.775 ;
        RECT 23.295 158.375 23.465 159.775 ;
        RECT 24.255 158.375 24.425 159.775 ;
        RECT 26.700 157.690 27.030 158.670 ;
        RECT 26.700 157.090 26.930 157.690 ;
        RECT 1.565 156.295 1.735 156.855 ;
        RECT 2.525 156.295 2.695 156.855 ;
        RECT 3.485 156.295 3.655 156.855 ;
        RECT 4.445 156.295 4.615 156.855 ;
        RECT 5.405 156.295 5.575 156.855 ;
        RECT 6.365 156.295 6.535 156.855 ;
        RECT 12.330 156.315 12.500 156.875 ;
        RECT 12.810 156.315 12.980 156.875 ;
        RECT 13.290 156.315 13.460 156.875 ;
        RECT 13.770 156.315 13.940 156.875 ;
        RECT 14.250 156.315 14.420 156.875 ;
        RECT 14.730 156.315 14.900 156.875 ;
        RECT 15.210 156.315 15.380 156.875 ;
        RECT 15.690 156.315 15.860 156.875 ;
        RECT 16.170 156.315 16.340 156.875 ;
        RECT 16.650 156.315 16.820 156.875 ;
        RECT 17.130 156.315 17.300 156.875 ;
        RECT 18.675 156.355 18.845 156.895 ;
        RECT 20.415 156.315 20.585 156.875 ;
        RECT 21.375 156.315 21.545 156.875 ;
        RECT 22.335 156.315 22.505 156.875 ;
        RECT 23.295 156.315 23.465 156.875 ;
        RECT 24.255 156.315 24.425 156.875 ;
        RECT 26.700 156.460 27.030 157.090 ;
        RECT 12.250 155.955 12.580 156.125 ;
        RECT 13.210 155.955 13.540 156.125 ;
        RECT 14.170 155.955 14.500 156.125 ;
        RECT 15.130 155.955 15.460 156.125 ;
        RECT 16.090 155.955 16.420 156.125 ;
        RECT 17.050 155.955 17.380 156.125 ;
        RECT 19.855 155.955 20.185 156.125 ;
        RECT 20.815 155.955 21.145 156.125 ;
        RECT 21.775 155.955 22.105 156.125 ;
        RECT 22.735 155.955 23.065 156.125 ;
        RECT 23.695 155.955 24.025 156.125 ;
        RECT 24.655 155.955 24.985 156.125 ;
        RECT 1.565 151.920 1.735 153.320 ;
        RECT 2.525 151.920 2.695 153.320 ;
        RECT 3.485 151.920 3.655 153.320 ;
        RECT 4.445 151.920 4.615 153.320 ;
        RECT 5.405 151.920 5.575 153.320 ;
        RECT 6.365 151.920 6.535 153.320 ;
        RECT 12.330 151.940 12.500 153.340 ;
        RECT 12.810 151.940 12.980 153.340 ;
        RECT 13.290 151.940 13.460 153.340 ;
        RECT 13.770 151.940 13.940 153.340 ;
        RECT 14.250 151.940 14.420 153.340 ;
        RECT 14.730 151.940 14.900 153.340 ;
        RECT 15.210 151.940 15.380 153.340 ;
        RECT 15.690 151.940 15.860 153.340 ;
        RECT 16.170 151.940 16.340 153.340 ;
        RECT 16.650 151.940 16.820 153.340 ;
        RECT 17.130 151.940 17.300 153.340 ;
        RECT 20.415 151.940 20.585 153.340 ;
        RECT 21.375 151.940 21.545 153.340 ;
        RECT 22.335 151.940 22.505 153.340 ;
        RECT 23.295 151.940 23.465 153.340 ;
        RECT 24.255 151.940 24.425 153.340 ;
        RECT 26.700 151.255 27.030 152.235 ;
        RECT 26.700 150.655 26.930 151.255 ;
        RECT 1.565 149.860 1.735 150.420 ;
        RECT 2.525 149.860 2.695 150.420 ;
        RECT 3.485 149.860 3.655 150.420 ;
        RECT 4.445 149.860 4.615 150.420 ;
        RECT 5.405 149.860 5.575 150.420 ;
        RECT 6.365 149.860 6.535 150.420 ;
        RECT 12.330 149.880 12.500 150.440 ;
        RECT 12.810 149.880 12.980 150.440 ;
        RECT 13.290 149.880 13.460 150.440 ;
        RECT 13.770 149.880 13.940 150.440 ;
        RECT 14.250 149.880 14.420 150.440 ;
        RECT 14.730 149.880 14.900 150.440 ;
        RECT 15.210 149.880 15.380 150.440 ;
        RECT 15.690 149.880 15.860 150.440 ;
        RECT 16.170 149.880 16.340 150.440 ;
        RECT 16.650 149.880 16.820 150.440 ;
        RECT 17.130 149.880 17.300 150.440 ;
        RECT 18.675 149.920 18.845 150.460 ;
        RECT 20.415 149.880 20.585 150.440 ;
        RECT 21.375 149.880 21.545 150.440 ;
        RECT 22.335 149.880 22.505 150.440 ;
        RECT 23.295 149.880 23.465 150.440 ;
        RECT 24.255 149.880 24.425 150.440 ;
        RECT 26.700 150.025 27.030 150.655 ;
        RECT 12.250 149.520 12.580 149.690 ;
        RECT 13.210 149.520 13.540 149.690 ;
        RECT 14.170 149.520 14.500 149.690 ;
        RECT 15.130 149.520 15.460 149.690 ;
        RECT 16.090 149.520 16.420 149.690 ;
        RECT 17.050 149.520 17.380 149.690 ;
        RECT 19.855 149.520 20.185 149.690 ;
        RECT 20.815 149.520 21.145 149.690 ;
        RECT 21.775 149.520 22.105 149.690 ;
        RECT 22.735 149.520 23.065 149.690 ;
        RECT 23.695 149.520 24.025 149.690 ;
        RECT 24.655 149.520 24.985 149.690 ;
        RECT 1.565 145.485 1.735 146.885 ;
        RECT 2.525 145.485 2.695 146.885 ;
        RECT 3.485 145.485 3.655 146.885 ;
        RECT 4.445 145.485 4.615 146.885 ;
        RECT 5.405 145.485 5.575 146.885 ;
        RECT 6.365 145.485 6.535 146.885 ;
        RECT 12.330 145.505 12.500 146.905 ;
        RECT 12.810 145.505 12.980 146.905 ;
        RECT 13.290 145.505 13.460 146.905 ;
        RECT 13.770 145.505 13.940 146.905 ;
        RECT 14.250 145.505 14.420 146.905 ;
        RECT 14.730 145.505 14.900 146.905 ;
        RECT 15.210 145.505 15.380 146.905 ;
        RECT 15.690 145.505 15.860 146.905 ;
        RECT 16.170 145.505 16.340 146.905 ;
        RECT 16.650 145.505 16.820 146.905 ;
        RECT 17.130 145.505 17.300 146.905 ;
        RECT 20.415 145.505 20.585 146.905 ;
        RECT 21.375 145.505 21.545 146.905 ;
        RECT 22.335 145.505 22.505 146.905 ;
        RECT 23.295 145.505 23.465 146.905 ;
        RECT 24.255 145.505 24.425 146.905 ;
        RECT 26.700 144.820 27.030 145.800 ;
        RECT 26.700 144.220 26.930 144.820 ;
        RECT 1.565 143.425 1.735 143.985 ;
        RECT 2.525 143.425 2.695 143.985 ;
        RECT 3.485 143.425 3.655 143.985 ;
        RECT 4.445 143.425 4.615 143.985 ;
        RECT 5.405 143.425 5.575 143.985 ;
        RECT 6.365 143.425 6.535 143.985 ;
        RECT 12.330 143.445 12.500 144.005 ;
        RECT 12.810 143.445 12.980 144.005 ;
        RECT 13.290 143.445 13.460 144.005 ;
        RECT 13.770 143.445 13.940 144.005 ;
        RECT 14.250 143.445 14.420 144.005 ;
        RECT 14.730 143.445 14.900 144.005 ;
        RECT 15.210 143.445 15.380 144.005 ;
        RECT 15.690 143.445 15.860 144.005 ;
        RECT 16.170 143.445 16.340 144.005 ;
        RECT 16.650 143.445 16.820 144.005 ;
        RECT 17.130 143.445 17.300 144.005 ;
        RECT 18.675 143.485 18.845 144.025 ;
        RECT 20.415 143.445 20.585 144.005 ;
        RECT 21.375 143.445 21.545 144.005 ;
        RECT 22.335 143.445 22.505 144.005 ;
        RECT 23.295 143.445 23.465 144.005 ;
        RECT 24.255 143.445 24.425 144.005 ;
        RECT 26.700 143.590 27.030 144.220 ;
        RECT 12.250 143.085 12.580 143.255 ;
        RECT 13.210 143.085 13.540 143.255 ;
        RECT 14.170 143.085 14.500 143.255 ;
        RECT 15.130 143.085 15.460 143.255 ;
        RECT 16.090 143.085 16.420 143.255 ;
        RECT 17.050 143.085 17.380 143.255 ;
        RECT 19.855 143.085 20.185 143.255 ;
        RECT 20.815 143.085 21.145 143.255 ;
        RECT 21.775 143.085 22.105 143.255 ;
        RECT 22.735 143.085 23.065 143.255 ;
        RECT 23.695 143.085 24.025 143.255 ;
        RECT 24.655 143.085 24.985 143.255 ;
        RECT 1.565 139.050 1.735 140.450 ;
        RECT 2.525 139.050 2.695 140.450 ;
        RECT 3.485 139.050 3.655 140.450 ;
        RECT 4.445 139.050 4.615 140.450 ;
        RECT 5.405 139.050 5.575 140.450 ;
        RECT 6.365 139.050 6.535 140.450 ;
        RECT 12.330 139.070 12.500 140.470 ;
        RECT 12.810 139.070 12.980 140.470 ;
        RECT 13.290 139.070 13.460 140.470 ;
        RECT 13.770 139.070 13.940 140.470 ;
        RECT 14.250 139.070 14.420 140.470 ;
        RECT 14.730 139.070 14.900 140.470 ;
        RECT 15.210 139.070 15.380 140.470 ;
        RECT 15.690 139.070 15.860 140.470 ;
        RECT 16.170 139.070 16.340 140.470 ;
        RECT 16.650 139.070 16.820 140.470 ;
        RECT 17.130 139.070 17.300 140.470 ;
        RECT 20.415 139.070 20.585 140.470 ;
        RECT 21.375 139.070 21.545 140.470 ;
        RECT 22.335 139.070 22.505 140.470 ;
        RECT 23.295 139.070 23.465 140.470 ;
        RECT 24.255 139.070 24.425 140.470 ;
        RECT 26.700 138.385 27.030 139.365 ;
        RECT 26.700 137.785 26.930 138.385 ;
        RECT 1.565 136.990 1.735 137.550 ;
        RECT 2.525 136.990 2.695 137.550 ;
        RECT 3.485 136.990 3.655 137.550 ;
        RECT 4.445 136.990 4.615 137.550 ;
        RECT 5.405 136.990 5.575 137.550 ;
        RECT 6.365 136.990 6.535 137.550 ;
        RECT 12.330 137.010 12.500 137.570 ;
        RECT 12.810 137.010 12.980 137.570 ;
        RECT 13.290 137.010 13.460 137.570 ;
        RECT 13.770 137.010 13.940 137.570 ;
        RECT 14.250 137.010 14.420 137.570 ;
        RECT 14.730 137.010 14.900 137.570 ;
        RECT 15.210 137.010 15.380 137.570 ;
        RECT 15.690 137.010 15.860 137.570 ;
        RECT 16.170 137.010 16.340 137.570 ;
        RECT 16.650 137.010 16.820 137.570 ;
        RECT 17.130 137.010 17.300 137.570 ;
        RECT 18.675 137.050 18.845 137.590 ;
        RECT 20.415 137.010 20.585 137.570 ;
        RECT 21.375 137.010 21.545 137.570 ;
        RECT 22.335 137.010 22.505 137.570 ;
        RECT 23.295 137.010 23.465 137.570 ;
        RECT 24.255 137.010 24.425 137.570 ;
        RECT 26.700 137.155 27.030 137.785 ;
        RECT 12.250 136.650 12.580 136.820 ;
        RECT 13.210 136.650 13.540 136.820 ;
        RECT 14.170 136.650 14.500 136.820 ;
        RECT 15.130 136.650 15.460 136.820 ;
        RECT 16.090 136.650 16.420 136.820 ;
        RECT 17.050 136.650 17.380 136.820 ;
        RECT 19.855 136.650 20.185 136.820 ;
        RECT 20.815 136.650 21.145 136.820 ;
        RECT 21.775 136.650 22.105 136.820 ;
        RECT 22.735 136.650 23.065 136.820 ;
        RECT 23.695 136.650 24.025 136.820 ;
        RECT 24.655 136.650 24.985 136.820 ;
        RECT 1.565 132.615 1.735 134.015 ;
        RECT 2.525 132.615 2.695 134.015 ;
        RECT 3.485 132.615 3.655 134.015 ;
        RECT 4.445 132.615 4.615 134.015 ;
        RECT 5.405 132.615 5.575 134.015 ;
        RECT 6.365 132.615 6.535 134.015 ;
        RECT 12.330 132.635 12.500 134.035 ;
        RECT 12.810 132.635 12.980 134.035 ;
        RECT 13.290 132.635 13.460 134.035 ;
        RECT 13.770 132.635 13.940 134.035 ;
        RECT 14.250 132.635 14.420 134.035 ;
        RECT 14.730 132.635 14.900 134.035 ;
        RECT 15.210 132.635 15.380 134.035 ;
        RECT 15.690 132.635 15.860 134.035 ;
        RECT 16.170 132.635 16.340 134.035 ;
        RECT 16.650 132.635 16.820 134.035 ;
        RECT 17.130 132.635 17.300 134.035 ;
        RECT 20.415 132.635 20.585 134.035 ;
        RECT 21.375 132.635 21.545 134.035 ;
        RECT 22.335 132.635 22.505 134.035 ;
        RECT 23.295 132.635 23.465 134.035 ;
        RECT 24.255 132.635 24.425 134.035 ;
        RECT 26.700 131.950 27.030 132.930 ;
        RECT 26.700 131.350 26.930 131.950 ;
        RECT 1.565 130.555 1.735 131.115 ;
        RECT 2.525 130.555 2.695 131.115 ;
        RECT 3.485 130.555 3.655 131.115 ;
        RECT 4.445 130.555 4.615 131.115 ;
        RECT 5.405 130.555 5.575 131.115 ;
        RECT 6.365 130.555 6.535 131.115 ;
        RECT 12.330 130.575 12.500 131.135 ;
        RECT 12.810 130.575 12.980 131.135 ;
        RECT 13.290 130.575 13.460 131.135 ;
        RECT 13.770 130.575 13.940 131.135 ;
        RECT 14.250 130.575 14.420 131.135 ;
        RECT 14.730 130.575 14.900 131.135 ;
        RECT 15.210 130.575 15.380 131.135 ;
        RECT 15.690 130.575 15.860 131.135 ;
        RECT 16.170 130.575 16.340 131.135 ;
        RECT 16.650 130.575 16.820 131.135 ;
        RECT 17.130 130.575 17.300 131.135 ;
        RECT 18.675 130.615 18.845 131.155 ;
        RECT 20.415 130.575 20.585 131.135 ;
        RECT 21.375 130.575 21.545 131.135 ;
        RECT 22.335 130.575 22.505 131.135 ;
        RECT 23.295 130.575 23.465 131.135 ;
        RECT 24.255 130.575 24.425 131.135 ;
        RECT 26.700 130.720 27.030 131.350 ;
        RECT 12.250 130.215 12.580 130.385 ;
        RECT 13.210 130.215 13.540 130.385 ;
        RECT 14.170 130.215 14.500 130.385 ;
        RECT 15.130 130.215 15.460 130.385 ;
        RECT 16.090 130.215 16.420 130.385 ;
        RECT 17.050 130.215 17.380 130.385 ;
        RECT 19.855 130.215 20.185 130.385 ;
        RECT 20.815 130.215 21.145 130.385 ;
        RECT 21.775 130.215 22.105 130.385 ;
        RECT 22.735 130.215 23.065 130.385 ;
        RECT 23.695 130.215 24.025 130.385 ;
        RECT 24.655 130.215 24.985 130.385 ;
        RECT 1.565 126.180 1.735 127.580 ;
        RECT 2.525 126.180 2.695 127.580 ;
        RECT 3.485 126.180 3.655 127.580 ;
        RECT 4.445 126.180 4.615 127.580 ;
        RECT 5.405 126.180 5.575 127.580 ;
        RECT 6.365 126.180 6.535 127.580 ;
        RECT 12.330 126.200 12.500 127.600 ;
        RECT 12.810 126.200 12.980 127.600 ;
        RECT 13.290 126.200 13.460 127.600 ;
        RECT 13.770 126.200 13.940 127.600 ;
        RECT 14.250 126.200 14.420 127.600 ;
        RECT 14.730 126.200 14.900 127.600 ;
        RECT 15.210 126.200 15.380 127.600 ;
        RECT 15.690 126.200 15.860 127.600 ;
        RECT 16.170 126.200 16.340 127.600 ;
        RECT 16.650 126.200 16.820 127.600 ;
        RECT 17.130 126.200 17.300 127.600 ;
        RECT 20.415 126.200 20.585 127.600 ;
        RECT 21.375 126.200 21.545 127.600 ;
        RECT 22.335 126.200 22.505 127.600 ;
        RECT 23.295 126.200 23.465 127.600 ;
        RECT 24.255 126.200 24.425 127.600 ;
        RECT 26.700 125.515 27.030 126.495 ;
        RECT 26.700 124.915 26.930 125.515 ;
        RECT 1.565 124.120 1.735 124.680 ;
        RECT 2.525 124.120 2.695 124.680 ;
        RECT 3.485 124.120 3.655 124.680 ;
        RECT 4.445 124.120 4.615 124.680 ;
        RECT 5.405 124.120 5.575 124.680 ;
        RECT 6.365 124.120 6.535 124.680 ;
        RECT 12.330 124.140 12.500 124.700 ;
        RECT 12.810 124.140 12.980 124.700 ;
        RECT 13.290 124.140 13.460 124.700 ;
        RECT 13.770 124.140 13.940 124.700 ;
        RECT 14.250 124.140 14.420 124.700 ;
        RECT 14.730 124.140 14.900 124.700 ;
        RECT 15.210 124.140 15.380 124.700 ;
        RECT 15.690 124.140 15.860 124.700 ;
        RECT 16.170 124.140 16.340 124.700 ;
        RECT 16.650 124.140 16.820 124.700 ;
        RECT 17.130 124.140 17.300 124.700 ;
        RECT 18.675 124.180 18.845 124.720 ;
        RECT 20.415 124.140 20.585 124.700 ;
        RECT 21.375 124.140 21.545 124.700 ;
        RECT 22.335 124.140 22.505 124.700 ;
        RECT 23.295 124.140 23.465 124.700 ;
        RECT 24.255 124.140 24.425 124.700 ;
        RECT 26.700 124.285 27.030 124.915 ;
        RECT 12.250 123.780 12.580 123.950 ;
        RECT 13.210 123.780 13.540 123.950 ;
        RECT 14.170 123.780 14.500 123.950 ;
        RECT 15.130 123.780 15.460 123.950 ;
        RECT 16.090 123.780 16.420 123.950 ;
        RECT 17.050 123.780 17.380 123.950 ;
        RECT 19.855 123.780 20.185 123.950 ;
        RECT 20.815 123.780 21.145 123.950 ;
        RECT 21.775 123.780 22.105 123.950 ;
        RECT 22.735 123.780 23.065 123.950 ;
        RECT 23.695 123.780 24.025 123.950 ;
        RECT 24.655 123.780 24.985 123.950 ;
        RECT 1.565 119.745 1.735 121.145 ;
        RECT 2.525 119.745 2.695 121.145 ;
        RECT 3.485 119.745 3.655 121.145 ;
        RECT 4.445 119.745 4.615 121.145 ;
        RECT 5.405 119.745 5.575 121.145 ;
        RECT 6.365 119.745 6.535 121.145 ;
        RECT 12.330 119.765 12.500 121.165 ;
        RECT 12.810 119.765 12.980 121.165 ;
        RECT 13.290 119.765 13.460 121.165 ;
        RECT 13.770 119.765 13.940 121.165 ;
        RECT 14.250 119.765 14.420 121.165 ;
        RECT 14.730 119.765 14.900 121.165 ;
        RECT 15.210 119.765 15.380 121.165 ;
        RECT 15.690 119.765 15.860 121.165 ;
        RECT 16.170 119.765 16.340 121.165 ;
        RECT 16.650 119.765 16.820 121.165 ;
        RECT 17.130 119.765 17.300 121.165 ;
        RECT 20.415 119.765 20.585 121.165 ;
        RECT 21.375 119.765 21.545 121.165 ;
        RECT 22.335 119.765 22.505 121.165 ;
        RECT 23.295 119.765 23.465 121.165 ;
        RECT 24.255 119.765 24.425 121.165 ;
        RECT 26.700 119.080 27.030 120.060 ;
        RECT 26.700 118.480 26.930 119.080 ;
        RECT 1.565 117.685 1.735 118.245 ;
        RECT 2.525 117.685 2.695 118.245 ;
        RECT 3.485 117.685 3.655 118.245 ;
        RECT 4.445 117.685 4.615 118.245 ;
        RECT 5.405 117.685 5.575 118.245 ;
        RECT 6.365 117.685 6.535 118.245 ;
        RECT 12.330 117.705 12.500 118.265 ;
        RECT 12.810 117.705 12.980 118.265 ;
        RECT 13.290 117.705 13.460 118.265 ;
        RECT 13.770 117.705 13.940 118.265 ;
        RECT 14.250 117.705 14.420 118.265 ;
        RECT 14.730 117.705 14.900 118.265 ;
        RECT 15.210 117.705 15.380 118.265 ;
        RECT 15.690 117.705 15.860 118.265 ;
        RECT 16.170 117.705 16.340 118.265 ;
        RECT 16.650 117.705 16.820 118.265 ;
        RECT 17.130 117.705 17.300 118.265 ;
        RECT 18.675 117.745 18.845 118.285 ;
        RECT 20.415 117.705 20.585 118.265 ;
        RECT 21.375 117.705 21.545 118.265 ;
        RECT 22.335 117.705 22.505 118.265 ;
        RECT 23.295 117.705 23.465 118.265 ;
        RECT 24.255 117.705 24.425 118.265 ;
        RECT 26.700 117.850 27.030 118.480 ;
        RECT 12.250 117.345 12.580 117.515 ;
        RECT 13.210 117.345 13.540 117.515 ;
        RECT 14.170 117.345 14.500 117.515 ;
        RECT 15.130 117.345 15.460 117.515 ;
        RECT 16.090 117.345 16.420 117.515 ;
        RECT 17.050 117.345 17.380 117.515 ;
        RECT 19.855 117.345 20.185 117.515 ;
        RECT 20.815 117.345 21.145 117.515 ;
        RECT 21.775 117.345 22.105 117.515 ;
        RECT 22.735 117.345 23.065 117.515 ;
        RECT 23.695 117.345 24.025 117.515 ;
        RECT 24.655 117.345 24.985 117.515 ;
        RECT 1.565 113.310 1.735 114.710 ;
        RECT 2.525 113.310 2.695 114.710 ;
        RECT 3.485 113.310 3.655 114.710 ;
        RECT 4.445 113.310 4.615 114.710 ;
        RECT 5.405 113.310 5.575 114.710 ;
        RECT 6.365 113.310 6.535 114.710 ;
        RECT 12.330 113.330 12.500 114.730 ;
        RECT 12.810 113.330 12.980 114.730 ;
        RECT 13.290 113.330 13.460 114.730 ;
        RECT 13.770 113.330 13.940 114.730 ;
        RECT 14.250 113.330 14.420 114.730 ;
        RECT 14.730 113.330 14.900 114.730 ;
        RECT 15.210 113.330 15.380 114.730 ;
        RECT 15.690 113.330 15.860 114.730 ;
        RECT 16.170 113.330 16.340 114.730 ;
        RECT 16.650 113.330 16.820 114.730 ;
        RECT 17.130 113.330 17.300 114.730 ;
        RECT 20.415 113.330 20.585 114.730 ;
        RECT 21.375 113.330 21.545 114.730 ;
        RECT 22.335 113.330 22.505 114.730 ;
        RECT 23.295 113.330 23.465 114.730 ;
        RECT 24.255 113.330 24.425 114.730 ;
        RECT 26.700 112.645 27.030 113.625 ;
        RECT 26.700 112.045 26.930 112.645 ;
        RECT 1.565 111.250 1.735 111.810 ;
        RECT 2.525 111.250 2.695 111.810 ;
        RECT 3.485 111.250 3.655 111.810 ;
        RECT 4.445 111.250 4.615 111.810 ;
        RECT 5.405 111.250 5.575 111.810 ;
        RECT 6.365 111.250 6.535 111.810 ;
        RECT 12.330 111.270 12.500 111.830 ;
        RECT 12.810 111.270 12.980 111.830 ;
        RECT 13.290 111.270 13.460 111.830 ;
        RECT 13.770 111.270 13.940 111.830 ;
        RECT 14.250 111.270 14.420 111.830 ;
        RECT 14.730 111.270 14.900 111.830 ;
        RECT 15.210 111.270 15.380 111.830 ;
        RECT 15.690 111.270 15.860 111.830 ;
        RECT 16.170 111.270 16.340 111.830 ;
        RECT 16.650 111.270 16.820 111.830 ;
        RECT 17.130 111.270 17.300 111.830 ;
        RECT 18.675 111.310 18.845 111.850 ;
        RECT 20.415 111.270 20.585 111.830 ;
        RECT 21.375 111.270 21.545 111.830 ;
        RECT 22.335 111.270 22.505 111.830 ;
        RECT 23.295 111.270 23.465 111.830 ;
        RECT 24.255 111.270 24.425 111.830 ;
        RECT 26.700 111.415 27.030 112.045 ;
        RECT 12.250 110.910 12.580 111.080 ;
        RECT 13.210 110.910 13.540 111.080 ;
        RECT 14.170 110.910 14.500 111.080 ;
        RECT 15.130 110.910 15.460 111.080 ;
        RECT 16.090 110.910 16.420 111.080 ;
        RECT 17.050 110.910 17.380 111.080 ;
        RECT 19.855 110.910 20.185 111.080 ;
        RECT 20.815 110.910 21.145 111.080 ;
        RECT 21.775 110.910 22.105 111.080 ;
        RECT 22.735 110.910 23.065 111.080 ;
        RECT 23.695 110.910 24.025 111.080 ;
        RECT 24.655 110.910 24.985 111.080 ;
        RECT 1.565 106.875 1.735 108.275 ;
        RECT 2.525 106.875 2.695 108.275 ;
        RECT 3.485 106.875 3.655 108.275 ;
        RECT 4.445 106.875 4.615 108.275 ;
        RECT 5.405 106.875 5.575 108.275 ;
        RECT 6.365 106.875 6.535 108.275 ;
        RECT 12.330 106.895 12.500 108.295 ;
        RECT 12.810 106.895 12.980 108.295 ;
        RECT 13.290 106.895 13.460 108.295 ;
        RECT 13.770 106.895 13.940 108.295 ;
        RECT 14.250 106.895 14.420 108.295 ;
        RECT 14.730 106.895 14.900 108.295 ;
        RECT 15.210 106.895 15.380 108.295 ;
        RECT 15.690 106.895 15.860 108.295 ;
        RECT 16.170 106.895 16.340 108.295 ;
        RECT 16.650 106.895 16.820 108.295 ;
        RECT 17.130 106.895 17.300 108.295 ;
        RECT 20.415 106.895 20.585 108.295 ;
        RECT 21.375 106.895 21.545 108.295 ;
        RECT 22.335 106.895 22.505 108.295 ;
        RECT 23.295 106.895 23.465 108.295 ;
        RECT 24.255 106.895 24.425 108.295 ;
        RECT 26.700 106.210 27.030 107.190 ;
        RECT 26.700 105.610 26.930 106.210 ;
        RECT 1.565 104.815 1.735 105.375 ;
        RECT 2.525 104.815 2.695 105.375 ;
        RECT 3.485 104.815 3.655 105.375 ;
        RECT 4.445 104.815 4.615 105.375 ;
        RECT 5.405 104.815 5.575 105.375 ;
        RECT 6.365 104.815 6.535 105.375 ;
        RECT 12.330 104.835 12.500 105.395 ;
        RECT 12.810 104.835 12.980 105.395 ;
        RECT 13.290 104.835 13.460 105.395 ;
        RECT 13.770 104.835 13.940 105.395 ;
        RECT 14.250 104.835 14.420 105.395 ;
        RECT 14.730 104.835 14.900 105.395 ;
        RECT 15.210 104.835 15.380 105.395 ;
        RECT 15.690 104.835 15.860 105.395 ;
        RECT 16.170 104.835 16.340 105.395 ;
        RECT 16.650 104.835 16.820 105.395 ;
        RECT 17.130 104.835 17.300 105.395 ;
        RECT 18.675 104.875 18.845 105.415 ;
        RECT 20.415 104.835 20.585 105.395 ;
        RECT 21.375 104.835 21.545 105.395 ;
        RECT 22.335 104.835 22.505 105.395 ;
        RECT 23.295 104.835 23.465 105.395 ;
        RECT 24.255 104.835 24.425 105.395 ;
        RECT 26.700 104.980 27.030 105.610 ;
        RECT 12.250 104.475 12.580 104.645 ;
        RECT 13.210 104.475 13.540 104.645 ;
        RECT 14.170 104.475 14.500 104.645 ;
        RECT 15.130 104.475 15.460 104.645 ;
        RECT 16.090 104.475 16.420 104.645 ;
        RECT 17.050 104.475 17.380 104.645 ;
        RECT 19.855 104.475 20.185 104.645 ;
        RECT 20.815 104.475 21.145 104.645 ;
        RECT 21.775 104.475 22.105 104.645 ;
        RECT 22.735 104.475 23.065 104.645 ;
        RECT 23.695 104.475 24.025 104.645 ;
        RECT 24.655 104.475 24.985 104.645 ;
        RECT 1.565 100.440 1.735 101.840 ;
        RECT 2.525 100.440 2.695 101.840 ;
        RECT 3.485 100.440 3.655 101.840 ;
        RECT 4.445 100.440 4.615 101.840 ;
        RECT 5.405 100.440 5.575 101.840 ;
        RECT 6.365 100.440 6.535 101.840 ;
        RECT 12.330 100.460 12.500 101.860 ;
        RECT 12.810 100.460 12.980 101.860 ;
        RECT 13.290 100.460 13.460 101.860 ;
        RECT 13.770 100.460 13.940 101.860 ;
        RECT 14.250 100.460 14.420 101.860 ;
        RECT 14.730 100.460 14.900 101.860 ;
        RECT 15.210 100.460 15.380 101.860 ;
        RECT 15.690 100.460 15.860 101.860 ;
        RECT 16.170 100.460 16.340 101.860 ;
        RECT 16.650 100.460 16.820 101.860 ;
        RECT 17.130 100.460 17.300 101.860 ;
        RECT 20.415 100.460 20.585 101.860 ;
        RECT 21.375 100.460 21.545 101.860 ;
        RECT 22.335 100.460 22.505 101.860 ;
        RECT 23.295 100.460 23.465 101.860 ;
        RECT 24.255 100.460 24.425 101.860 ;
        RECT 26.700 99.775 27.030 100.755 ;
        RECT 26.700 99.175 26.930 99.775 ;
        RECT 1.565 98.380 1.735 98.940 ;
        RECT 2.525 98.380 2.695 98.940 ;
        RECT 3.485 98.380 3.655 98.940 ;
        RECT 4.445 98.380 4.615 98.940 ;
        RECT 5.405 98.380 5.575 98.940 ;
        RECT 6.365 98.380 6.535 98.940 ;
        RECT 12.330 98.400 12.500 98.960 ;
        RECT 12.810 98.400 12.980 98.960 ;
        RECT 13.290 98.400 13.460 98.960 ;
        RECT 13.770 98.400 13.940 98.960 ;
        RECT 14.250 98.400 14.420 98.960 ;
        RECT 14.730 98.400 14.900 98.960 ;
        RECT 15.210 98.400 15.380 98.960 ;
        RECT 15.690 98.400 15.860 98.960 ;
        RECT 16.170 98.400 16.340 98.960 ;
        RECT 16.650 98.400 16.820 98.960 ;
        RECT 17.130 98.400 17.300 98.960 ;
        RECT 18.675 98.440 18.845 98.980 ;
        RECT 20.415 98.400 20.585 98.960 ;
        RECT 21.375 98.400 21.545 98.960 ;
        RECT 22.335 98.400 22.505 98.960 ;
        RECT 23.295 98.400 23.465 98.960 ;
        RECT 24.255 98.400 24.425 98.960 ;
        RECT 26.700 98.545 27.030 99.175 ;
        RECT 12.250 98.040 12.580 98.210 ;
        RECT 13.210 98.040 13.540 98.210 ;
        RECT 14.170 98.040 14.500 98.210 ;
        RECT 15.130 98.040 15.460 98.210 ;
        RECT 16.090 98.040 16.420 98.210 ;
        RECT 17.050 98.040 17.380 98.210 ;
        RECT 19.855 98.040 20.185 98.210 ;
        RECT 20.815 98.040 21.145 98.210 ;
        RECT 21.775 98.040 22.105 98.210 ;
        RECT 22.735 98.040 23.065 98.210 ;
        RECT 23.695 98.040 24.025 98.210 ;
        RECT 24.655 98.040 24.985 98.210 ;
        RECT 1.565 94.005 1.735 95.405 ;
        RECT 2.525 94.005 2.695 95.405 ;
        RECT 3.485 94.005 3.655 95.405 ;
        RECT 4.445 94.005 4.615 95.405 ;
        RECT 5.405 94.005 5.575 95.405 ;
        RECT 6.365 94.005 6.535 95.405 ;
        RECT 12.330 94.025 12.500 95.425 ;
        RECT 12.810 94.025 12.980 95.425 ;
        RECT 13.290 94.025 13.460 95.425 ;
        RECT 13.770 94.025 13.940 95.425 ;
        RECT 14.250 94.025 14.420 95.425 ;
        RECT 14.730 94.025 14.900 95.425 ;
        RECT 15.210 94.025 15.380 95.425 ;
        RECT 15.690 94.025 15.860 95.425 ;
        RECT 16.170 94.025 16.340 95.425 ;
        RECT 16.650 94.025 16.820 95.425 ;
        RECT 17.130 94.025 17.300 95.425 ;
        RECT 20.415 94.025 20.585 95.425 ;
        RECT 21.375 94.025 21.545 95.425 ;
        RECT 22.335 94.025 22.505 95.425 ;
        RECT 23.295 94.025 23.465 95.425 ;
        RECT 24.255 94.025 24.425 95.425 ;
        RECT 26.700 93.340 27.030 94.320 ;
        RECT 26.700 92.740 26.930 93.340 ;
        RECT 1.565 91.945 1.735 92.505 ;
        RECT 2.525 91.945 2.695 92.505 ;
        RECT 3.485 91.945 3.655 92.505 ;
        RECT 4.445 91.945 4.615 92.505 ;
        RECT 5.405 91.945 5.575 92.505 ;
        RECT 6.365 91.945 6.535 92.505 ;
        RECT 12.330 91.965 12.500 92.525 ;
        RECT 12.810 91.965 12.980 92.525 ;
        RECT 13.290 91.965 13.460 92.525 ;
        RECT 13.770 91.965 13.940 92.525 ;
        RECT 14.250 91.965 14.420 92.525 ;
        RECT 14.730 91.965 14.900 92.525 ;
        RECT 15.210 91.965 15.380 92.525 ;
        RECT 15.690 91.965 15.860 92.525 ;
        RECT 16.170 91.965 16.340 92.525 ;
        RECT 16.650 91.965 16.820 92.525 ;
        RECT 17.130 91.965 17.300 92.525 ;
        RECT 18.675 92.005 18.845 92.545 ;
        RECT 20.415 91.965 20.585 92.525 ;
        RECT 21.375 91.965 21.545 92.525 ;
        RECT 22.335 91.965 22.505 92.525 ;
        RECT 23.295 91.965 23.465 92.525 ;
        RECT 24.255 91.965 24.425 92.525 ;
        RECT 26.700 92.110 27.030 92.740 ;
        RECT 12.250 91.605 12.580 91.775 ;
        RECT 13.210 91.605 13.540 91.775 ;
        RECT 14.170 91.605 14.500 91.775 ;
        RECT 15.130 91.605 15.460 91.775 ;
        RECT 16.090 91.605 16.420 91.775 ;
        RECT 17.050 91.605 17.380 91.775 ;
        RECT 19.855 91.605 20.185 91.775 ;
        RECT 20.815 91.605 21.145 91.775 ;
        RECT 21.775 91.605 22.105 91.775 ;
        RECT 22.735 91.605 23.065 91.775 ;
        RECT 23.695 91.605 24.025 91.775 ;
        RECT 24.655 91.605 24.985 91.775 ;
        RECT 1.565 87.570 1.735 88.970 ;
        RECT 2.525 87.570 2.695 88.970 ;
        RECT 3.485 87.570 3.655 88.970 ;
        RECT 4.445 87.570 4.615 88.970 ;
        RECT 5.405 87.570 5.575 88.970 ;
        RECT 6.365 87.570 6.535 88.970 ;
        RECT 12.330 87.590 12.500 88.990 ;
        RECT 12.810 87.590 12.980 88.990 ;
        RECT 13.290 87.590 13.460 88.990 ;
        RECT 13.770 87.590 13.940 88.990 ;
        RECT 14.250 87.590 14.420 88.990 ;
        RECT 14.730 87.590 14.900 88.990 ;
        RECT 15.210 87.590 15.380 88.990 ;
        RECT 15.690 87.590 15.860 88.990 ;
        RECT 16.170 87.590 16.340 88.990 ;
        RECT 16.650 87.590 16.820 88.990 ;
        RECT 17.130 87.590 17.300 88.990 ;
        RECT 20.415 87.590 20.585 88.990 ;
        RECT 21.375 87.590 21.545 88.990 ;
        RECT 22.335 87.590 22.505 88.990 ;
        RECT 23.295 87.590 23.465 88.990 ;
        RECT 24.255 87.590 24.425 88.990 ;
        RECT 26.700 86.905 27.030 87.885 ;
        RECT 26.700 86.305 26.930 86.905 ;
        RECT 1.565 85.510 1.735 86.070 ;
        RECT 2.525 85.510 2.695 86.070 ;
        RECT 3.485 85.510 3.655 86.070 ;
        RECT 4.445 85.510 4.615 86.070 ;
        RECT 5.405 85.510 5.575 86.070 ;
        RECT 6.365 85.510 6.535 86.070 ;
        RECT 12.330 85.530 12.500 86.090 ;
        RECT 12.810 85.530 12.980 86.090 ;
        RECT 13.290 85.530 13.460 86.090 ;
        RECT 13.770 85.530 13.940 86.090 ;
        RECT 14.250 85.530 14.420 86.090 ;
        RECT 14.730 85.530 14.900 86.090 ;
        RECT 15.210 85.530 15.380 86.090 ;
        RECT 15.690 85.530 15.860 86.090 ;
        RECT 16.170 85.530 16.340 86.090 ;
        RECT 16.650 85.530 16.820 86.090 ;
        RECT 17.130 85.530 17.300 86.090 ;
        RECT 18.675 85.570 18.845 86.110 ;
        RECT 20.415 85.530 20.585 86.090 ;
        RECT 21.375 85.530 21.545 86.090 ;
        RECT 22.335 85.530 22.505 86.090 ;
        RECT 23.295 85.530 23.465 86.090 ;
        RECT 24.255 85.530 24.425 86.090 ;
        RECT 26.700 85.675 27.030 86.305 ;
        RECT 12.250 85.170 12.580 85.340 ;
        RECT 13.210 85.170 13.540 85.340 ;
        RECT 14.170 85.170 14.500 85.340 ;
        RECT 15.130 85.170 15.460 85.340 ;
        RECT 16.090 85.170 16.420 85.340 ;
        RECT 17.050 85.170 17.380 85.340 ;
        RECT 19.855 85.170 20.185 85.340 ;
        RECT 20.815 85.170 21.145 85.340 ;
        RECT 21.775 85.170 22.105 85.340 ;
        RECT 22.735 85.170 23.065 85.340 ;
        RECT 23.695 85.170 24.025 85.340 ;
        RECT 24.655 85.170 24.985 85.340 ;
        RECT 1.565 81.135 1.735 82.535 ;
        RECT 2.525 81.135 2.695 82.535 ;
        RECT 3.485 81.135 3.655 82.535 ;
        RECT 4.445 81.135 4.615 82.535 ;
        RECT 5.405 81.135 5.575 82.535 ;
        RECT 6.365 81.135 6.535 82.535 ;
        RECT 12.330 81.155 12.500 82.555 ;
        RECT 12.810 81.155 12.980 82.555 ;
        RECT 13.290 81.155 13.460 82.555 ;
        RECT 13.770 81.155 13.940 82.555 ;
        RECT 14.250 81.155 14.420 82.555 ;
        RECT 14.730 81.155 14.900 82.555 ;
        RECT 15.210 81.155 15.380 82.555 ;
        RECT 15.690 81.155 15.860 82.555 ;
        RECT 16.170 81.155 16.340 82.555 ;
        RECT 16.650 81.155 16.820 82.555 ;
        RECT 17.130 81.155 17.300 82.555 ;
        RECT 20.415 81.155 20.585 82.555 ;
        RECT 21.375 81.155 21.545 82.555 ;
        RECT 22.335 81.155 22.505 82.555 ;
        RECT 23.295 81.155 23.465 82.555 ;
        RECT 24.255 81.155 24.425 82.555 ;
        RECT 26.700 80.470 27.030 81.450 ;
        RECT 26.700 79.870 26.930 80.470 ;
        RECT 1.565 79.075 1.735 79.635 ;
        RECT 2.525 79.075 2.695 79.635 ;
        RECT 3.485 79.075 3.655 79.635 ;
        RECT 4.445 79.075 4.615 79.635 ;
        RECT 5.405 79.075 5.575 79.635 ;
        RECT 6.365 79.075 6.535 79.635 ;
        RECT 12.330 79.095 12.500 79.655 ;
        RECT 12.810 79.095 12.980 79.655 ;
        RECT 13.290 79.095 13.460 79.655 ;
        RECT 13.770 79.095 13.940 79.655 ;
        RECT 14.250 79.095 14.420 79.655 ;
        RECT 14.730 79.095 14.900 79.655 ;
        RECT 15.210 79.095 15.380 79.655 ;
        RECT 15.690 79.095 15.860 79.655 ;
        RECT 16.170 79.095 16.340 79.655 ;
        RECT 16.650 79.095 16.820 79.655 ;
        RECT 17.130 79.095 17.300 79.655 ;
        RECT 18.675 79.135 18.845 79.675 ;
        RECT 20.415 79.095 20.585 79.655 ;
        RECT 21.375 79.095 21.545 79.655 ;
        RECT 22.335 79.095 22.505 79.655 ;
        RECT 23.295 79.095 23.465 79.655 ;
        RECT 24.255 79.095 24.425 79.655 ;
        RECT 26.700 79.240 27.030 79.870 ;
        RECT 12.250 78.735 12.580 78.905 ;
        RECT 13.210 78.735 13.540 78.905 ;
        RECT 14.170 78.735 14.500 78.905 ;
        RECT 15.130 78.735 15.460 78.905 ;
        RECT 16.090 78.735 16.420 78.905 ;
        RECT 17.050 78.735 17.380 78.905 ;
        RECT 19.855 78.735 20.185 78.905 ;
        RECT 20.815 78.735 21.145 78.905 ;
        RECT 21.775 78.735 22.105 78.905 ;
        RECT 22.735 78.735 23.065 78.905 ;
        RECT 23.695 78.735 24.025 78.905 ;
        RECT 24.655 78.735 24.985 78.905 ;
        RECT 1.565 74.700 1.735 76.100 ;
        RECT 2.525 74.700 2.695 76.100 ;
        RECT 3.485 74.700 3.655 76.100 ;
        RECT 4.445 74.700 4.615 76.100 ;
        RECT 5.405 74.700 5.575 76.100 ;
        RECT 6.365 74.700 6.535 76.100 ;
        RECT 12.330 74.720 12.500 76.120 ;
        RECT 12.810 74.720 12.980 76.120 ;
        RECT 13.290 74.720 13.460 76.120 ;
        RECT 13.770 74.720 13.940 76.120 ;
        RECT 14.250 74.720 14.420 76.120 ;
        RECT 14.730 74.720 14.900 76.120 ;
        RECT 15.210 74.720 15.380 76.120 ;
        RECT 15.690 74.720 15.860 76.120 ;
        RECT 16.170 74.720 16.340 76.120 ;
        RECT 16.650 74.720 16.820 76.120 ;
        RECT 17.130 74.720 17.300 76.120 ;
        RECT 20.415 74.720 20.585 76.120 ;
        RECT 21.375 74.720 21.545 76.120 ;
        RECT 22.335 74.720 22.505 76.120 ;
        RECT 23.295 74.720 23.465 76.120 ;
        RECT 24.255 74.720 24.425 76.120 ;
        RECT 26.700 74.035 27.030 75.015 ;
        RECT 26.700 73.435 26.930 74.035 ;
        RECT 1.565 72.640 1.735 73.200 ;
        RECT 2.525 72.640 2.695 73.200 ;
        RECT 3.485 72.640 3.655 73.200 ;
        RECT 4.445 72.640 4.615 73.200 ;
        RECT 5.405 72.640 5.575 73.200 ;
        RECT 6.365 72.640 6.535 73.200 ;
        RECT 12.330 72.660 12.500 73.220 ;
        RECT 12.810 72.660 12.980 73.220 ;
        RECT 13.290 72.660 13.460 73.220 ;
        RECT 13.770 72.660 13.940 73.220 ;
        RECT 14.250 72.660 14.420 73.220 ;
        RECT 14.730 72.660 14.900 73.220 ;
        RECT 15.210 72.660 15.380 73.220 ;
        RECT 15.690 72.660 15.860 73.220 ;
        RECT 16.170 72.660 16.340 73.220 ;
        RECT 16.650 72.660 16.820 73.220 ;
        RECT 17.130 72.660 17.300 73.220 ;
        RECT 18.675 72.700 18.845 73.240 ;
        RECT 20.415 72.660 20.585 73.220 ;
        RECT 21.375 72.660 21.545 73.220 ;
        RECT 22.335 72.660 22.505 73.220 ;
        RECT 23.295 72.660 23.465 73.220 ;
        RECT 24.255 72.660 24.425 73.220 ;
        RECT 26.700 72.805 27.030 73.435 ;
        RECT 12.250 72.300 12.580 72.470 ;
        RECT 13.210 72.300 13.540 72.470 ;
        RECT 14.170 72.300 14.500 72.470 ;
        RECT 15.130 72.300 15.460 72.470 ;
        RECT 16.090 72.300 16.420 72.470 ;
        RECT 17.050 72.300 17.380 72.470 ;
        RECT 19.855 72.300 20.185 72.470 ;
        RECT 20.815 72.300 21.145 72.470 ;
        RECT 21.775 72.300 22.105 72.470 ;
        RECT 22.735 72.300 23.065 72.470 ;
        RECT 23.695 72.300 24.025 72.470 ;
        RECT 24.655 72.300 24.985 72.470 ;
        RECT 1.565 68.265 1.735 69.665 ;
        RECT 2.525 68.265 2.695 69.665 ;
        RECT 3.485 68.265 3.655 69.665 ;
        RECT 4.445 68.265 4.615 69.665 ;
        RECT 5.405 68.265 5.575 69.665 ;
        RECT 6.365 68.265 6.535 69.665 ;
        RECT 12.330 68.285 12.500 69.685 ;
        RECT 12.810 68.285 12.980 69.685 ;
        RECT 13.290 68.285 13.460 69.685 ;
        RECT 13.770 68.285 13.940 69.685 ;
        RECT 14.250 68.285 14.420 69.685 ;
        RECT 14.730 68.285 14.900 69.685 ;
        RECT 15.210 68.285 15.380 69.685 ;
        RECT 15.690 68.285 15.860 69.685 ;
        RECT 16.170 68.285 16.340 69.685 ;
        RECT 16.650 68.285 16.820 69.685 ;
        RECT 17.130 68.285 17.300 69.685 ;
        RECT 20.415 68.285 20.585 69.685 ;
        RECT 21.375 68.285 21.545 69.685 ;
        RECT 22.335 68.285 22.505 69.685 ;
        RECT 23.295 68.285 23.465 69.685 ;
        RECT 24.255 68.285 24.425 69.685 ;
        RECT 26.700 67.600 27.030 68.580 ;
        RECT 26.700 67.000 26.930 67.600 ;
        RECT 1.565 66.205 1.735 66.765 ;
        RECT 2.525 66.205 2.695 66.765 ;
        RECT 3.485 66.205 3.655 66.765 ;
        RECT 4.445 66.205 4.615 66.765 ;
        RECT 5.405 66.205 5.575 66.765 ;
        RECT 6.365 66.205 6.535 66.765 ;
        RECT 12.330 66.225 12.500 66.785 ;
        RECT 12.810 66.225 12.980 66.785 ;
        RECT 13.290 66.225 13.460 66.785 ;
        RECT 13.770 66.225 13.940 66.785 ;
        RECT 14.250 66.225 14.420 66.785 ;
        RECT 14.730 66.225 14.900 66.785 ;
        RECT 15.210 66.225 15.380 66.785 ;
        RECT 15.690 66.225 15.860 66.785 ;
        RECT 16.170 66.225 16.340 66.785 ;
        RECT 16.650 66.225 16.820 66.785 ;
        RECT 17.130 66.225 17.300 66.785 ;
        RECT 18.675 66.265 18.845 66.805 ;
        RECT 20.415 66.225 20.585 66.785 ;
        RECT 21.375 66.225 21.545 66.785 ;
        RECT 22.335 66.225 22.505 66.785 ;
        RECT 23.295 66.225 23.465 66.785 ;
        RECT 24.255 66.225 24.425 66.785 ;
        RECT 26.700 66.370 27.030 67.000 ;
        RECT 12.250 65.865 12.580 66.035 ;
        RECT 13.210 65.865 13.540 66.035 ;
        RECT 14.170 65.865 14.500 66.035 ;
        RECT 15.130 65.865 15.460 66.035 ;
        RECT 16.090 65.865 16.420 66.035 ;
        RECT 17.050 65.865 17.380 66.035 ;
        RECT 19.855 65.865 20.185 66.035 ;
        RECT 20.815 65.865 21.145 66.035 ;
        RECT 21.775 65.865 22.105 66.035 ;
        RECT 22.735 65.865 23.065 66.035 ;
        RECT 23.695 65.865 24.025 66.035 ;
        RECT 24.655 65.865 24.985 66.035 ;
        RECT 1.565 61.830 1.735 63.230 ;
        RECT 2.525 61.830 2.695 63.230 ;
        RECT 3.485 61.830 3.655 63.230 ;
        RECT 4.445 61.830 4.615 63.230 ;
        RECT 5.405 61.830 5.575 63.230 ;
        RECT 6.365 61.830 6.535 63.230 ;
        RECT 12.330 61.850 12.500 63.250 ;
        RECT 12.810 61.850 12.980 63.250 ;
        RECT 13.290 61.850 13.460 63.250 ;
        RECT 13.770 61.850 13.940 63.250 ;
        RECT 14.250 61.850 14.420 63.250 ;
        RECT 14.730 61.850 14.900 63.250 ;
        RECT 15.210 61.850 15.380 63.250 ;
        RECT 15.690 61.850 15.860 63.250 ;
        RECT 16.170 61.850 16.340 63.250 ;
        RECT 16.650 61.850 16.820 63.250 ;
        RECT 17.130 61.850 17.300 63.250 ;
        RECT 20.415 61.850 20.585 63.250 ;
        RECT 21.375 61.850 21.545 63.250 ;
        RECT 22.335 61.850 22.505 63.250 ;
        RECT 23.295 61.850 23.465 63.250 ;
        RECT 24.255 61.850 24.425 63.250 ;
        RECT 26.700 61.165 27.030 62.145 ;
        RECT 26.700 60.565 26.930 61.165 ;
        RECT 1.565 59.770 1.735 60.330 ;
        RECT 2.525 59.770 2.695 60.330 ;
        RECT 3.485 59.770 3.655 60.330 ;
        RECT 4.445 59.770 4.615 60.330 ;
        RECT 5.405 59.770 5.575 60.330 ;
        RECT 6.365 59.770 6.535 60.330 ;
        RECT 12.330 59.790 12.500 60.350 ;
        RECT 12.810 59.790 12.980 60.350 ;
        RECT 13.290 59.790 13.460 60.350 ;
        RECT 13.770 59.790 13.940 60.350 ;
        RECT 14.250 59.790 14.420 60.350 ;
        RECT 14.730 59.790 14.900 60.350 ;
        RECT 15.210 59.790 15.380 60.350 ;
        RECT 15.690 59.790 15.860 60.350 ;
        RECT 16.170 59.790 16.340 60.350 ;
        RECT 16.650 59.790 16.820 60.350 ;
        RECT 17.130 59.790 17.300 60.350 ;
        RECT 18.675 59.830 18.845 60.370 ;
        RECT 20.415 59.790 20.585 60.350 ;
        RECT 21.375 59.790 21.545 60.350 ;
        RECT 22.335 59.790 22.505 60.350 ;
        RECT 23.295 59.790 23.465 60.350 ;
        RECT 24.255 59.790 24.425 60.350 ;
        RECT 26.700 59.935 27.030 60.565 ;
        RECT 12.250 59.430 12.580 59.600 ;
        RECT 13.210 59.430 13.540 59.600 ;
        RECT 14.170 59.430 14.500 59.600 ;
        RECT 15.130 59.430 15.460 59.600 ;
        RECT 16.090 59.430 16.420 59.600 ;
        RECT 17.050 59.430 17.380 59.600 ;
        RECT 19.855 59.430 20.185 59.600 ;
        RECT 20.815 59.430 21.145 59.600 ;
        RECT 21.775 59.430 22.105 59.600 ;
        RECT 22.735 59.430 23.065 59.600 ;
        RECT 23.695 59.430 24.025 59.600 ;
        RECT 24.655 59.430 24.985 59.600 ;
        RECT 1.565 55.395 1.735 56.795 ;
        RECT 2.525 55.395 2.695 56.795 ;
        RECT 3.485 55.395 3.655 56.795 ;
        RECT 4.445 55.395 4.615 56.795 ;
        RECT 5.405 55.395 5.575 56.795 ;
        RECT 6.365 55.395 6.535 56.795 ;
        RECT 12.330 55.415 12.500 56.815 ;
        RECT 12.810 55.415 12.980 56.815 ;
        RECT 13.290 55.415 13.460 56.815 ;
        RECT 13.770 55.415 13.940 56.815 ;
        RECT 14.250 55.415 14.420 56.815 ;
        RECT 14.730 55.415 14.900 56.815 ;
        RECT 15.210 55.415 15.380 56.815 ;
        RECT 15.690 55.415 15.860 56.815 ;
        RECT 16.170 55.415 16.340 56.815 ;
        RECT 16.650 55.415 16.820 56.815 ;
        RECT 17.130 55.415 17.300 56.815 ;
        RECT 20.415 55.415 20.585 56.815 ;
        RECT 21.375 55.415 21.545 56.815 ;
        RECT 22.335 55.415 22.505 56.815 ;
        RECT 23.295 55.415 23.465 56.815 ;
        RECT 24.255 55.415 24.425 56.815 ;
        RECT 26.700 54.730 27.030 55.710 ;
        RECT 26.700 54.130 26.930 54.730 ;
        RECT 1.565 53.335 1.735 53.895 ;
        RECT 2.525 53.335 2.695 53.895 ;
        RECT 3.485 53.335 3.655 53.895 ;
        RECT 4.445 53.335 4.615 53.895 ;
        RECT 5.405 53.335 5.575 53.895 ;
        RECT 6.365 53.335 6.535 53.895 ;
        RECT 12.330 53.355 12.500 53.915 ;
        RECT 12.810 53.355 12.980 53.915 ;
        RECT 13.290 53.355 13.460 53.915 ;
        RECT 13.770 53.355 13.940 53.915 ;
        RECT 14.250 53.355 14.420 53.915 ;
        RECT 14.730 53.355 14.900 53.915 ;
        RECT 15.210 53.355 15.380 53.915 ;
        RECT 15.690 53.355 15.860 53.915 ;
        RECT 16.170 53.355 16.340 53.915 ;
        RECT 16.650 53.355 16.820 53.915 ;
        RECT 17.130 53.355 17.300 53.915 ;
        RECT 18.675 53.395 18.845 53.935 ;
        RECT 20.415 53.355 20.585 53.915 ;
        RECT 21.375 53.355 21.545 53.915 ;
        RECT 22.335 53.355 22.505 53.915 ;
        RECT 23.295 53.355 23.465 53.915 ;
        RECT 24.255 53.355 24.425 53.915 ;
        RECT 26.700 53.500 27.030 54.130 ;
        RECT 12.250 52.995 12.580 53.165 ;
        RECT 13.210 52.995 13.540 53.165 ;
        RECT 14.170 52.995 14.500 53.165 ;
        RECT 15.130 52.995 15.460 53.165 ;
        RECT 16.090 52.995 16.420 53.165 ;
        RECT 17.050 52.995 17.380 53.165 ;
        RECT 19.855 52.995 20.185 53.165 ;
        RECT 20.815 52.995 21.145 53.165 ;
        RECT 21.775 52.995 22.105 53.165 ;
        RECT 22.735 52.995 23.065 53.165 ;
        RECT 23.695 52.995 24.025 53.165 ;
        RECT 24.655 52.995 24.985 53.165 ;
        RECT 1.565 48.960 1.735 50.360 ;
        RECT 2.525 48.960 2.695 50.360 ;
        RECT 3.485 48.960 3.655 50.360 ;
        RECT 4.445 48.960 4.615 50.360 ;
        RECT 5.405 48.960 5.575 50.360 ;
        RECT 6.365 48.960 6.535 50.360 ;
        RECT 12.330 48.980 12.500 50.380 ;
        RECT 12.810 48.980 12.980 50.380 ;
        RECT 13.290 48.980 13.460 50.380 ;
        RECT 13.770 48.980 13.940 50.380 ;
        RECT 14.250 48.980 14.420 50.380 ;
        RECT 14.730 48.980 14.900 50.380 ;
        RECT 15.210 48.980 15.380 50.380 ;
        RECT 15.690 48.980 15.860 50.380 ;
        RECT 16.170 48.980 16.340 50.380 ;
        RECT 16.650 48.980 16.820 50.380 ;
        RECT 17.130 48.980 17.300 50.380 ;
        RECT 20.415 48.980 20.585 50.380 ;
        RECT 21.375 48.980 21.545 50.380 ;
        RECT 22.335 48.980 22.505 50.380 ;
        RECT 23.295 48.980 23.465 50.380 ;
        RECT 24.255 48.980 24.425 50.380 ;
        RECT 26.700 48.295 27.030 49.275 ;
        RECT 26.700 47.695 26.930 48.295 ;
        RECT 1.565 46.900 1.735 47.460 ;
        RECT 2.525 46.900 2.695 47.460 ;
        RECT 3.485 46.900 3.655 47.460 ;
        RECT 4.445 46.900 4.615 47.460 ;
        RECT 5.405 46.900 5.575 47.460 ;
        RECT 6.365 46.900 6.535 47.460 ;
        RECT 12.330 46.920 12.500 47.480 ;
        RECT 12.810 46.920 12.980 47.480 ;
        RECT 13.290 46.920 13.460 47.480 ;
        RECT 13.770 46.920 13.940 47.480 ;
        RECT 14.250 46.920 14.420 47.480 ;
        RECT 14.730 46.920 14.900 47.480 ;
        RECT 15.210 46.920 15.380 47.480 ;
        RECT 15.690 46.920 15.860 47.480 ;
        RECT 16.170 46.920 16.340 47.480 ;
        RECT 16.650 46.920 16.820 47.480 ;
        RECT 17.130 46.920 17.300 47.480 ;
        RECT 18.675 46.960 18.845 47.500 ;
        RECT 20.415 46.920 20.585 47.480 ;
        RECT 21.375 46.920 21.545 47.480 ;
        RECT 22.335 46.920 22.505 47.480 ;
        RECT 23.295 46.920 23.465 47.480 ;
        RECT 24.255 46.920 24.425 47.480 ;
        RECT 26.700 47.065 27.030 47.695 ;
        RECT 12.250 46.560 12.580 46.730 ;
        RECT 13.210 46.560 13.540 46.730 ;
        RECT 14.170 46.560 14.500 46.730 ;
        RECT 15.130 46.560 15.460 46.730 ;
        RECT 16.090 46.560 16.420 46.730 ;
        RECT 17.050 46.560 17.380 46.730 ;
        RECT 19.855 46.560 20.185 46.730 ;
        RECT 20.815 46.560 21.145 46.730 ;
        RECT 21.775 46.560 22.105 46.730 ;
        RECT 22.735 46.560 23.065 46.730 ;
        RECT 23.695 46.560 24.025 46.730 ;
        RECT 24.655 46.560 24.985 46.730 ;
        RECT 1.565 42.525 1.735 43.925 ;
        RECT 2.525 42.525 2.695 43.925 ;
        RECT 3.485 42.525 3.655 43.925 ;
        RECT 4.445 42.525 4.615 43.925 ;
        RECT 5.405 42.525 5.575 43.925 ;
        RECT 6.365 42.525 6.535 43.925 ;
        RECT 12.330 42.545 12.500 43.945 ;
        RECT 12.810 42.545 12.980 43.945 ;
        RECT 13.290 42.545 13.460 43.945 ;
        RECT 13.770 42.545 13.940 43.945 ;
        RECT 14.250 42.545 14.420 43.945 ;
        RECT 14.730 42.545 14.900 43.945 ;
        RECT 15.210 42.545 15.380 43.945 ;
        RECT 15.690 42.545 15.860 43.945 ;
        RECT 16.170 42.545 16.340 43.945 ;
        RECT 16.650 42.545 16.820 43.945 ;
        RECT 17.130 42.545 17.300 43.945 ;
        RECT 20.415 42.545 20.585 43.945 ;
        RECT 21.375 42.545 21.545 43.945 ;
        RECT 22.335 42.545 22.505 43.945 ;
        RECT 23.295 42.545 23.465 43.945 ;
        RECT 24.255 42.545 24.425 43.945 ;
        RECT 26.700 41.860 27.030 42.840 ;
        RECT 26.700 41.260 26.930 41.860 ;
        RECT 1.565 40.465 1.735 41.025 ;
        RECT 2.525 40.465 2.695 41.025 ;
        RECT 3.485 40.465 3.655 41.025 ;
        RECT 4.445 40.465 4.615 41.025 ;
        RECT 5.405 40.465 5.575 41.025 ;
        RECT 6.365 40.465 6.535 41.025 ;
        RECT 12.330 40.485 12.500 41.045 ;
        RECT 12.810 40.485 12.980 41.045 ;
        RECT 13.290 40.485 13.460 41.045 ;
        RECT 13.770 40.485 13.940 41.045 ;
        RECT 14.250 40.485 14.420 41.045 ;
        RECT 14.730 40.485 14.900 41.045 ;
        RECT 15.210 40.485 15.380 41.045 ;
        RECT 15.690 40.485 15.860 41.045 ;
        RECT 16.170 40.485 16.340 41.045 ;
        RECT 16.650 40.485 16.820 41.045 ;
        RECT 17.130 40.485 17.300 41.045 ;
        RECT 18.675 40.525 18.845 41.065 ;
        RECT 20.415 40.485 20.585 41.045 ;
        RECT 21.375 40.485 21.545 41.045 ;
        RECT 22.335 40.485 22.505 41.045 ;
        RECT 23.295 40.485 23.465 41.045 ;
        RECT 24.255 40.485 24.425 41.045 ;
        RECT 26.700 40.630 27.030 41.260 ;
        RECT 12.250 40.125 12.580 40.295 ;
        RECT 13.210 40.125 13.540 40.295 ;
        RECT 14.170 40.125 14.500 40.295 ;
        RECT 15.130 40.125 15.460 40.295 ;
        RECT 16.090 40.125 16.420 40.295 ;
        RECT 17.050 40.125 17.380 40.295 ;
        RECT 19.855 40.125 20.185 40.295 ;
        RECT 20.815 40.125 21.145 40.295 ;
        RECT 21.775 40.125 22.105 40.295 ;
        RECT 22.735 40.125 23.065 40.295 ;
        RECT 23.695 40.125 24.025 40.295 ;
        RECT 24.655 40.125 24.985 40.295 ;
        RECT 1.565 36.090 1.735 37.490 ;
        RECT 2.525 36.090 2.695 37.490 ;
        RECT 3.485 36.090 3.655 37.490 ;
        RECT 4.445 36.090 4.615 37.490 ;
        RECT 5.405 36.090 5.575 37.490 ;
        RECT 6.365 36.090 6.535 37.490 ;
        RECT 12.330 36.110 12.500 37.510 ;
        RECT 12.810 36.110 12.980 37.510 ;
        RECT 13.290 36.110 13.460 37.510 ;
        RECT 13.770 36.110 13.940 37.510 ;
        RECT 14.250 36.110 14.420 37.510 ;
        RECT 14.730 36.110 14.900 37.510 ;
        RECT 15.210 36.110 15.380 37.510 ;
        RECT 15.690 36.110 15.860 37.510 ;
        RECT 16.170 36.110 16.340 37.510 ;
        RECT 16.650 36.110 16.820 37.510 ;
        RECT 17.130 36.110 17.300 37.510 ;
        RECT 20.415 36.110 20.585 37.510 ;
        RECT 21.375 36.110 21.545 37.510 ;
        RECT 22.335 36.110 22.505 37.510 ;
        RECT 23.295 36.110 23.465 37.510 ;
        RECT 24.255 36.110 24.425 37.510 ;
        RECT 26.700 35.425 27.030 36.405 ;
        RECT 26.700 34.825 26.930 35.425 ;
        RECT 1.565 34.030 1.735 34.590 ;
        RECT 2.525 34.030 2.695 34.590 ;
        RECT 3.485 34.030 3.655 34.590 ;
        RECT 4.445 34.030 4.615 34.590 ;
        RECT 5.405 34.030 5.575 34.590 ;
        RECT 6.365 34.030 6.535 34.590 ;
        RECT 12.330 34.050 12.500 34.610 ;
        RECT 12.810 34.050 12.980 34.610 ;
        RECT 13.290 34.050 13.460 34.610 ;
        RECT 13.770 34.050 13.940 34.610 ;
        RECT 14.250 34.050 14.420 34.610 ;
        RECT 14.730 34.050 14.900 34.610 ;
        RECT 15.210 34.050 15.380 34.610 ;
        RECT 15.690 34.050 15.860 34.610 ;
        RECT 16.170 34.050 16.340 34.610 ;
        RECT 16.650 34.050 16.820 34.610 ;
        RECT 17.130 34.050 17.300 34.610 ;
        RECT 18.675 34.090 18.845 34.630 ;
        RECT 20.415 34.050 20.585 34.610 ;
        RECT 21.375 34.050 21.545 34.610 ;
        RECT 22.335 34.050 22.505 34.610 ;
        RECT 23.295 34.050 23.465 34.610 ;
        RECT 24.255 34.050 24.425 34.610 ;
        RECT 26.700 34.195 27.030 34.825 ;
        RECT 12.250 33.690 12.580 33.860 ;
        RECT 13.210 33.690 13.540 33.860 ;
        RECT 14.170 33.690 14.500 33.860 ;
        RECT 15.130 33.690 15.460 33.860 ;
        RECT 16.090 33.690 16.420 33.860 ;
        RECT 17.050 33.690 17.380 33.860 ;
        RECT 19.855 33.690 20.185 33.860 ;
        RECT 20.815 33.690 21.145 33.860 ;
        RECT 21.775 33.690 22.105 33.860 ;
        RECT 22.735 33.690 23.065 33.860 ;
        RECT 23.695 33.690 24.025 33.860 ;
        RECT 24.655 33.690 24.985 33.860 ;
        RECT 1.565 29.655 1.735 31.055 ;
        RECT 2.525 29.655 2.695 31.055 ;
        RECT 3.485 29.655 3.655 31.055 ;
        RECT 4.445 29.655 4.615 31.055 ;
        RECT 5.405 29.655 5.575 31.055 ;
        RECT 6.365 29.655 6.535 31.055 ;
        RECT 12.330 29.675 12.500 31.075 ;
        RECT 12.810 29.675 12.980 31.075 ;
        RECT 13.290 29.675 13.460 31.075 ;
        RECT 13.770 29.675 13.940 31.075 ;
        RECT 14.250 29.675 14.420 31.075 ;
        RECT 14.730 29.675 14.900 31.075 ;
        RECT 15.210 29.675 15.380 31.075 ;
        RECT 15.690 29.675 15.860 31.075 ;
        RECT 16.170 29.675 16.340 31.075 ;
        RECT 16.650 29.675 16.820 31.075 ;
        RECT 17.130 29.675 17.300 31.075 ;
        RECT 20.415 29.675 20.585 31.075 ;
        RECT 21.375 29.675 21.545 31.075 ;
        RECT 22.335 29.675 22.505 31.075 ;
        RECT 23.295 29.675 23.465 31.075 ;
        RECT 24.255 29.675 24.425 31.075 ;
        RECT 26.700 28.990 27.030 29.970 ;
        RECT 26.700 28.390 26.930 28.990 ;
        RECT 1.565 27.595 1.735 28.155 ;
        RECT 2.525 27.595 2.695 28.155 ;
        RECT 3.485 27.595 3.655 28.155 ;
        RECT 4.445 27.595 4.615 28.155 ;
        RECT 5.405 27.595 5.575 28.155 ;
        RECT 6.365 27.595 6.535 28.155 ;
        RECT 12.330 27.615 12.500 28.175 ;
        RECT 12.810 27.615 12.980 28.175 ;
        RECT 13.290 27.615 13.460 28.175 ;
        RECT 13.770 27.615 13.940 28.175 ;
        RECT 14.250 27.615 14.420 28.175 ;
        RECT 14.730 27.615 14.900 28.175 ;
        RECT 15.210 27.615 15.380 28.175 ;
        RECT 15.690 27.615 15.860 28.175 ;
        RECT 16.170 27.615 16.340 28.175 ;
        RECT 16.650 27.615 16.820 28.175 ;
        RECT 17.130 27.615 17.300 28.175 ;
        RECT 18.675 27.655 18.845 28.195 ;
        RECT 20.415 27.615 20.585 28.175 ;
        RECT 21.375 27.615 21.545 28.175 ;
        RECT 22.335 27.615 22.505 28.175 ;
        RECT 23.295 27.615 23.465 28.175 ;
        RECT 24.255 27.615 24.425 28.175 ;
        RECT 26.700 27.760 27.030 28.390 ;
        RECT 12.250 27.255 12.580 27.425 ;
        RECT 13.210 27.255 13.540 27.425 ;
        RECT 14.170 27.255 14.500 27.425 ;
        RECT 15.130 27.255 15.460 27.425 ;
        RECT 16.090 27.255 16.420 27.425 ;
        RECT 17.050 27.255 17.380 27.425 ;
        RECT 19.855 27.255 20.185 27.425 ;
        RECT 20.815 27.255 21.145 27.425 ;
        RECT 21.775 27.255 22.105 27.425 ;
        RECT 22.735 27.255 23.065 27.425 ;
        RECT 23.695 27.255 24.025 27.425 ;
        RECT 24.655 27.255 24.985 27.425 ;
        RECT 1.565 23.220 1.735 24.620 ;
        RECT 2.525 23.220 2.695 24.620 ;
        RECT 3.485 23.220 3.655 24.620 ;
        RECT 4.445 23.220 4.615 24.620 ;
        RECT 5.405 23.220 5.575 24.620 ;
        RECT 6.365 23.220 6.535 24.620 ;
        RECT 12.330 23.240 12.500 24.640 ;
        RECT 12.810 23.240 12.980 24.640 ;
        RECT 13.290 23.240 13.460 24.640 ;
        RECT 13.770 23.240 13.940 24.640 ;
        RECT 14.250 23.240 14.420 24.640 ;
        RECT 14.730 23.240 14.900 24.640 ;
        RECT 15.210 23.240 15.380 24.640 ;
        RECT 15.690 23.240 15.860 24.640 ;
        RECT 16.170 23.240 16.340 24.640 ;
        RECT 16.650 23.240 16.820 24.640 ;
        RECT 17.130 23.240 17.300 24.640 ;
        RECT 20.415 23.240 20.585 24.640 ;
        RECT 21.375 23.240 21.545 24.640 ;
        RECT 22.335 23.240 22.505 24.640 ;
        RECT 23.295 23.240 23.465 24.640 ;
        RECT 24.255 23.240 24.425 24.640 ;
        RECT 26.700 22.555 27.030 23.535 ;
        RECT 26.700 21.955 26.930 22.555 ;
        RECT 1.565 21.160 1.735 21.720 ;
        RECT 2.525 21.160 2.695 21.720 ;
        RECT 3.485 21.160 3.655 21.720 ;
        RECT 4.445 21.160 4.615 21.720 ;
        RECT 5.405 21.160 5.575 21.720 ;
        RECT 6.365 21.160 6.535 21.720 ;
        RECT 12.330 21.180 12.500 21.740 ;
        RECT 12.810 21.180 12.980 21.740 ;
        RECT 13.290 21.180 13.460 21.740 ;
        RECT 13.770 21.180 13.940 21.740 ;
        RECT 14.250 21.180 14.420 21.740 ;
        RECT 14.730 21.180 14.900 21.740 ;
        RECT 15.210 21.180 15.380 21.740 ;
        RECT 15.690 21.180 15.860 21.740 ;
        RECT 16.170 21.180 16.340 21.740 ;
        RECT 16.650 21.180 16.820 21.740 ;
        RECT 17.130 21.180 17.300 21.740 ;
        RECT 18.675 21.220 18.845 21.760 ;
        RECT 20.415 21.180 20.585 21.740 ;
        RECT 21.375 21.180 21.545 21.740 ;
        RECT 22.335 21.180 22.505 21.740 ;
        RECT 23.295 21.180 23.465 21.740 ;
        RECT 24.255 21.180 24.425 21.740 ;
        RECT 26.700 21.325 27.030 21.955 ;
        RECT 12.250 20.820 12.580 20.990 ;
        RECT 13.210 20.820 13.540 20.990 ;
        RECT 14.170 20.820 14.500 20.990 ;
        RECT 15.130 20.820 15.460 20.990 ;
        RECT 16.090 20.820 16.420 20.990 ;
        RECT 17.050 20.820 17.380 20.990 ;
        RECT 19.855 20.820 20.185 20.990 ;
        RECT 20.815 20.820 21.145 20.990 ;
        RECT 21.775 20.820 22.105 20.990 ;
        RECT 22.735 20.820 23.065 20.990 ;
        RECT 23.695 20.820 24.025 20.990 ;
        RECT 24.655 20.820 24.985 20.990 ;
        RECT 1.565 16.785 1.735 18.185 ;
        RECT 2.525 16.785 2.695 18.185 ;
        RECT 3.485 16.785 3.655 18.185 ;
        RECT 4.445 16.785 4.615 18.185 ;
        RECT 5.405 16.785 5.575 18.185 ;
        RECT 6.365 16.785 6.535 18.185 ;
        RECT 12.330 16.805 12.500 18.205 ;
        RECT 12.810 16.805 12.980 18.205 ;
        RECT 13.290 16.805 13.460 18.205 ;
        RECT 13.770 16.805 13.940 18.205 ;
        RECT 14.250 16.805 14.420 18.205 ;
        RECT 14.730 16.805 14.900 18.205 ;
        RECT 15.210 16.805 15.380 18.205 ;
        RECT 15.690 16.805 15.860 18.205 ;
        RECT 16.170 16.805 16.340 18.205 ;
        RECT 16.650 16.805 16.820 18.205 ;
        RECT 17.130 16.805 17.300 18.205 ;
        RECT 20.415 16.805 20.585 18.205 ;
        RECT 21.375 16.805 21.545 18.205 ;
        RECT 22.335 16.805 22.505 18.205 ;
        RECT 23.295 16.805 23.465 18.205 ;
        RECT 24.255 16.805 24.425 18.205 ;
        RECT 26.700 16.120 27.030 17.100 ;
        RECT 26.700 15.520 26.930 16.120 ;
        RECT 1.565 14.725 1.735 15.285 ;
        RECT 2.525 14.725 2.695 15.285 ;
        RECT 3.485 14.725 3.655 15.285 ;
        RECT 4.445 14.725 4.615 15.285 ;
        RECT 5.405 14.725 5.575 15.285 ;
        RECT 6.365 14.725 6.535 15.285 ;
        RECT 12.330 14.745 12.500 15.305 ;
        RECT 12.810 14.745 12.980 15.305 ;
        RECT 13.290 14.745 13.460 15.305 ;
        RECT 13.770 14.745 13.940 15.305 ;
        RECT 14.250 14.745 14.420 15.305 ;
        RECT 14.730 14.745 14.900 15.305 ;
        RECT 15.210 14.745 15.380 15.305 ;
        RECT 15.690 14.745 15.860 15.305 ;
        RECT 16.170 14.745 16.340 15.305 ;
        RECT 16.650 14.745 16.820 15.305 ;
        RECT 17.130 14.745 17.300 15.305 ;
        RECT 18.675 14.785 18.845 15.325 ;
        RECT 20.415 14.745 20.585 15.305 ;
        RECT 21.375 14.745 21.545 15.305 ;
        RECT 22.335 14.745 22.505 15.305 ;
        RECT 23.295 14.745 23.465 15.305 ;
        RECT 24.255 14.745 24.425 15.305 ;
        RECT 26.700 14.890 27.030 15.520 ;
        RECT 12.250 14.385 12.580 14.555 ;
        RECT 13.210 14.385 13.540 14.555 ;
        RECT 14.170 14.385 14.500 14.555 ;
        RECT 15.130 14.385 15.460 14.555 ;
        RECT 16.090 14.385 16.420 14.555 ;
        RECT 17.050 14.385 17.380 14.555 ;
        RECT 19.855 14.385 20.185 14.555 ;
        RECT 20.815 14.385 21.145 14.555 ;
        RECT 21.775 14.385 22.105 14.555 ;
        RECT 22.735 14.385 23.065 14.555 ;
        RECT 23.695 14.385 24.025 14.555 ;
        RECT 24.655 14.385 24.985 14.555 ;
        RECT 1.565 10.350 1.735 11.750 ;
        RECT 2.525 10.350 2.695 11.750 ;
        RECT 3.485 10.350 3.655 11.750 ;
        RECT 4.445 10.350 4.615 11.750 ;
        RECT 5.405 10.350 5.575 11.750 ;
        RECT 6.365 10.350 6.535 11.750 ;
        RECT 12.330 10.370 12.500 11.770 ;
        RECT 12.810 10.370 12.980 11.770 ;
        RECT 13.290 10.370 13.460 11.770 ;
        RECT 13.770 10.370 13.940 11.770 ;
        RECT 14.250 10.370 14.420 11.770 ;
        RECT 14.730 10.370 14.900 11.770 ;
        RECT 15.210 10.370 15.380 11.770 ;
        RECT 15.690 10.370 15.860 11.770 ;
        RECT 16.170 10.370 16.340 11.770 ;
        RECT 16.650 10.370 16.820 11.770 ;
        RECT 17.130 10.370 17.300 11.770 ;
        RECT 20.415 10.370 20.585 11.770 ;
        RECT 21.375 10.370 21.545 11.770 ;
        RECT 22.335 10.370 22.505 11.770 ;
        RECT 23.295 10.370 23.465 11.770 ;
        RECT 24.255 10.370 24.425 11.770 ;
        RECT 26.700 9.685 27.030 10.665 ;
        RECT 26.700 9.085 26.930 9.685 ;
        RECT 1.565 8.290 1.735 8.850 ;
        RECT 2.525 8.290 2.695 8.850 ;
        RECT 3.485 8.290 3.655 8.850 ;
        RECT 4.445 8.290 4.615 8.850 ;
        RECT 5.405 8.290 5.575 8.850 ;
        RECT 6.365 8.290 6.535 8.850 ;
        RECT 12.330 8.310 12.500 8.870 ;
        RECT 12.810 8.310 12.980 8.870 ;
        RECT 13.290 8.310 13.460 8.870 ;
        RECT 13.770 8.310 13.940 8.870 ;
        RECT 14.250 8.310 14.420 8.870 ;
        RECT 14.730 8.310 14.900 8.870 ;
        RECT 15.210 8.310 15.380 8.870 ;
        RECT 15.690 8.310 15.860 8.870 ;
        RECT 16.170 8.310 16.340 8.870 ;
        RECT 16.650 8.310 16.820 8.870 ;
        RECT 17.130 8.310 17.300 8.870 ;
        RECT 18.675 8.350 18.845 8.890 ;
        RECT 20.415 8.310 20.585 8.870 ;
        RECT 21.375 8.310 21.545 8.870 ;
        RECT 22.335 8.310 22.505 8.870 ;
        RECT 23.295 8.310 23.465 8.870 ;
        RECT 24.255 8.310 24.425 8.870 ;
        RECT 26.700 8.455 27.030 9.085 ;
        RECT 12.250 7.950 12.580 8.120 ;
        RECT 13.210 7.950 13.540 8.120 ;
        RECT 14.170 7.950 14.500 8.120 ;
        RECT 15.130 7.950 15.460 8.120 ;
        RECT 16.090 7.950 16.420 8.120 ;
        RECT 17.050 7.950 17.380 8.120 ;
        RECT 19.855 7.950 20.185 8.120 ;
        RECT 20.815 7.950 21.145 8.120 ;
        RECT 21.775 7.950 22.105 8.120 ;
        RECT 22.735 7.950 23.065 8.120 ;
        RECT 23.695 7.950 24.025 8.120 ;
        RECT 24.655 7.950 24.985 8.120 ;
        RECT 1.565 3.915 1.735 5.315 ;
        RECT 2.525 3.915 2.695 5.315 ;
        RECT 3.485 3.915 3.655 5.315 ;
        RECT 4.445 3.915 4.615 5.315 ;
        RECT 5.405 3.915 5.575 5.315 ;
        RECT 6.365 3.915 6.535 5.315 ;
        RECT 12.330 3.935 12.500 5.335 ;
        RECT 12.810 3.935 12.980 5.335 ;
        RECT 13.290 3.935 13.460 5.335 ;
        RECT 13.770 3.935 13.940 5.335 ;
        RECT 14.250 3.935 14.420 5.335 ;
        RECT 14.730 3.935 14.900 5.335 ;
        RECT 15.210 3.935 15.380 5.335 ;
        RECT 15.690 3.935 15.860 5.335 ;
        RECT 16.170 3.935 16.340 5.335 ;
        RECT 16.650 3.935 16.820 5.335 ;
        RECT 17.130 3.935 17.300 5.335 ;
        RECT 20.415 3.935 20.585 5.335 ;
        RECT 21.375 3.935 21.545 5.335 ;
        RECT 22.335 3.935 22.505 5.335 ;
        RECT 23.295 3.935 23.465 5.335 ;
        RECT 24.255 3.935 24.425 5.335 ;
        RECT 26.700 3.250 27.030 4.230 ;
        RECT 26.700 2.650 26.930 3.250 ;
        RECT 1.565 1.855 1.735 2.415 ;
        RECT 2.525 1.855 2.695 2.415 ;
        RECT 3.485 1.855 3.655 2.415 ;
        RECT 4.445 1.855 4.615 2.415 ;
        RECT 5.405 1.855 5.575 2.415 ;
        RECT 6.365 1.855 6.535 2.415 ;
        RECT 12.330 1.875 12.500 2.435 ;
        RECT 12.810 1.875 12.980 2.435 ;
        RECT 13.290 1.875 13.460 2.435 ;
        RECT 13.770 1.875 13.940 2.435 ;
        RECT 14.250 1.875 14.420 2.435 ;
        RECT 14.730 1.875 14.900 2.435 ;
        RECT 15.210 1.875 15.380 2.435 ;
        RECT 15.690 1.875 15.860 2.435 ;
        RECT 16.170 1.875 16.340 2.435 ;
        RECT 16.650 1.875 16.820 2.435 ;
        RECT 17.130 1.875 17.300 2.435 ;
        RECT 18.675 1.915 18.845 2.455 ;
        RECT 20.415 1.875 20.585 2.435 ;
        RECT 21.375 1.875 21.545 2.435 ;
        RECT 22.335 1.875 22.505 2.435 ;
        RECT 23.295 1.875 23.465 2.435 ;
        RECT 24.255 1.875 24.425 2.435 ;
        RECT 26.700 2.020 27.030 2.650 ;
        RECT 12.250 1.515 12.580 1.685 ;
        RECT 13.210 1.515 13.540 1.685 ;
        RECT 14.170 1.515 14.500 1.685 ;
        RECT 15.130 1.515 15.460 1.685 ;
        RECT 16.090 1.515 16.420 1.685 ;
        RECT 17.050 1.515 17.380 1.685 ;
        RECT 19.855 1.515 20.185 1.685 ;
        RECT 20.815 1.515 21.145 1.685 ;
        RECT 21.775 1.515 22.105 1.685 ;
        RECT 22.735 1.515 23.065 1.685 ;
        RECT 23.695 1.515 24.025 1.685 ;
        RECT 24.655 1.515 24.985 1.685 ;
      LAYER mcon ;
        RECT 1.565 204.375 1.735 204.545 ;
        RECT 1.565 204.015 1.735 204.185 ;
        RECT 1.565 203.655 1.735 203.825 ;
        RECT 2.525 204.375 2.695 204.545 ;
        RECT 2.525 204.015 2.695 204.185 ;
        RECT 2.525 203.655 2.695 203.825 ;
        RECT 3.485 204.375 3.655 204.545 ;
        RECT 3.485 204.015 3.655 204.185 ;
        RECT 3.485 203.655 3.655 203.825 ;
        RECT 4.445 204.375 4.615 204.545 ;
        RECT 4.445 204.015 4.615 204.185 ;
        RECT 4.445 203.655 4.615 203.825 ;
        RECT 5.405 204.375 5.575 204.545 ;
        RECT 5.405 204.015 5.575 204.185 ;
        RECT 5.405 203.655 5.575 203.825 ;
        RECT 6.365 204.375 6.535 204.545 ;
        RECT 6.365 204.015 6.535 204.185 ;
        RECT 6.365 203.655 6.535 203.825 ;
        RECT 12.330 204.395 12.500 204.565 ;
        RECT 12.330 204.035 12.500 204.205 ;
        RECT 12.330 203.675 12.500 203.845 ;
        RECT 12.810 204.395 12.980 204.565 ;
        RECT 12.810 204.035 12.980 204.205 ;
        RECT 12.810 203.675 12.980 203.845 ;
        RECT 13.290 204.395 13.460 204.565 ;
        RECT 13.290 204.035 13.460 204.205 ;
        RECT 13.290 203.675 13.460 203.845 ;
        RECT 13.770 204.395 13.940 204.565 ;
        RECT 13.770 204.035 13.940 204.205 ;
        RECT 13.770 203.675 13.940 203.845 ;
        RECT 14.250 204.395 14.420 204.565 ;
        RECT 14.250 204.035 14.420 204.205 ;
        RECT 14.250 203.675 14.420 203.845 ;
        RECT 14.730 204.395 14.900 204.565 ;
        RECT 14.730 204.035 14.900 204.205 ;
        RECT 14.730 203.675 14.900 203.845 ;
        RECT 15.210 204.395 15.380 204.565 ;
        RECT 15.210 204.035 15.380 204.205 ;
        RECT 15.210 203.675 15.380 203.845 ;
        RECT 15.690 204.395 15.860 204.565 ;
        RECT 15.690 204.035 15.860 204.205 ;
        RECT 15.690 203.675 15.860 203.845 ;
        RECT 16.170 204.395 16.340 204.565 ;
        RECT 16.170 204.035 16.340 204.205 ;
        RECT 16.170 203.675 16.340 203.845 ;
        RECT 16.650 204.395 16.820 204.565 ;
        RECT 16.650 204.035 16.820 204.205 ;
        RECT 16.650 203.675 16.820 203.845 ;
        RECT 17.130 204.395 17.300 204.565 ;
        RECT 17.130 204.035 17.300 204.205 ;
        RECT 17.130 203.675 17.300 203.845 ;
        RECT 20.415 204.395 20.585 204.565 ;
        RECT 20.415 204.035 20.585 204.205 ;
        RECT 20.415 203.675 20.585 203.845 ;
        RECT 21.375 204.395 21.545 204.565 ;
        RECT 21.375 204.035 21.545 204.205 ;
        RECT 21.375 203.675 21.545 203.845 ;
        RECT 22.335 204.395 22.505 204.565 ;
        RECT 22.335 204.035 22.505 204.205 ;
        RECT 22.335 203.675 22.505 203.845 ;
        RECT 23.295 204.395 23.465 204.565 ;
        RECT 23.295 204.035 23.465 204.205 ;
        RECT 23.295 203.675 23.465 203.845 ;
        RECT 24.255 204.395 24.425 204.565 ;
        RECT 24.255 204.035 24.425 204.205 ;
        RECT 24.255 203.675 24.425 203.845 ;
        RECT 26.740 202.315 26.910 202.485 ;
        RECT 1.565 201.535 1.735 201.705 ;
        RECT 2.525 201.535 2.695 201.705 ;
        RECT 3.485 201.535 3.655 201.705 ;
        RECT 4.445 201.535 4.615 201.705 ;
        RECT 5.405 201.535 5.575 201.705 ;
        RECT 6.365 201.535 6.535 201.705 ;
        RECT 12.330 201.555 12.500 201.725 ;
        RECT 12.810 201.555 12.980 201.725 ;
        RECT 13.290 201.555 13.460 201.725 ;
        RECT 13.770 201.555 13.940 201.725 ;
        RECT 14.250 201.555 14.420 201.725 ;
        RECT 14.730 201.555 14.900 201.725 ;
        RECT 15.210 201.555 15.380 201.725 ;
        RECT 15.690 201.555 15.860 201.725 ;
        RECT 16.170 201.555 16.340 201.725 ;
        RECT 16.650 201.555 16.820 201.725 ;
        RECT 17.130 201.555 17.300 201.725 ;
        RECT 18.675 201.480 18.845 201.860 ;
        RECT 20.415 201.555 20.585 201.725 ;
        RECT 21.375 201.555 21.545 201.725 ;
        RECT 22.335 201.555 22.505 201.725 ;
        RECT 23.295 201.555 23.465 201.725 ;
        RECT 24.255 201.555 24.425 201.725 ;
        RECT 12.330 201.000 12.500 201.170 ;
        RECT 13.290 201.000 13.460 201.170 ;
        RECT 14.250 201.000 14.420 201.170 ;
        RECT 15.210 201.000 15.380 201.170 ;
        RECT 16.170 201.000 16.340 201.170 ;
        RECT 17.130 201.000 17.300 201.170 ;
        RECT 19.935 201.000 20.105 201.170 ;
        RECT 20.895 201.000 21.065 201.170 ;
        RECT 21.855 201.000 22.025 201.170 ;
        RECT 22.815 201.000 22.985 201.170 ;
        RECT 23.775 201.000 23.945 201.170 ;
        RECT 24.735 201.000 24.905 201.170 ;
        RECT 1.565 197.940 1.735 198.110 ;
        RECT 1.565 197.580 1.735 197.750 ;
        RECT 1.565 197.220 1.735 197.390 ;
        RECT 2.525 197.940 2.695 198.110 ;
        RECT 2.525 197.580 2.695 197.750 ;
        RECT 2.525 197.220 2.695 197.390 ;
        RECT 3.485 197.940 3.655 198.110 ;
        RECT 3.485 197.580 3.655 197.750 ;
        RECT 3.485 197.220 3.655 197.390 ;
        RECT 4.445 197.940 4.615 198.110 ;
        RECT 4.445 197.580 4.615 197.750 ;
        RECT 4.445 197.220 4.615 197.390 ;
        RECT 5.405 197.940 5.575 198.110 ;
        RECT 5.405 197.580 5.575 197.750 ;
        RECT 5.405 197.220 5.575 197.390 ;
        RECT 6.365 197.940 6.535 198.110 ;
        RECT 6.365 197.580 6.535 197.750 ;
        RECT 6.365 197.220 6.535 197.390 ;
        RECT 12.330 197.960 12.500 198.130 ;
        RECT 12.330 197.600 12.500 197.770 ;
        RECT 12.330 197.240 12.500 197.410 ;
        RECT 12.810 197.960 12.980 198.130 ;
        RECT 12.810 197.600 12.980 197.770 ;
        RECT 12.810 197.240 12.980 197.410 ;
        RECT 13.290 197.960 13.460 198.130 ;
        RECT 13.290 197.600 13.460 197.770 ;
        RECT 13.290 197.240 13.460 197.410 ;
        RECT 13.770 197.960 13.940 198.130 ;
        RECT 13.770 197.600 13.940 197.770 ;
        RECT 13.770 197.240 13.940 197.410 ;
        RECT 14.250 197.960 14.420 198.130 ;
        RECT 14.250 197.600 14.420 197.770 ;
        RECT 14.250 197.240 14.420 197.410 ;
        RECT 14.730 197.960 14.900 198.130 ;
        RECT 14.730 197.600 14.900 197.770 ;
        RECT 14.730 197.240 14.900 197.410 ;
        RECT 15.210 197.960 15.380 198.130 ;
        RECT 15.210 197.600 15.380 197.770 ;
        RECT 15.210 197.240 15.380 197.410 ;
        RECT 15.690 197.960 15.860 198.130 ;
        RECT 15.690 197.600 15.860 197.770 ;
        RECT 15.690 197.240 15.860 197.410 ;
        RECT 16.170 197.960 16.340 198.130 ;
        RECT 16.170 197.600 16.340 197.770 ;
        RECT 16.170 197.240 16.340 197.410 ;
        RECT 16.650 197.960 16.820 198.130 ;
        RECT 16.650 197.600 16.820 197.770 ;
        RECT 16.650 197.240 16.820 197.410 ;
        RECT 17.130 197.960 17.300 198.130 ;
        RECT 17.130 197.600 17.300 197.770 ;
        RECT 17.130 197.240 17.300 197.410 ;
        RECT 20.415 197.960 20.585 198.130 ;
        RECT 20.415 197.600 20.585 197.770 ;
        RECT 20.415 197.240 20.585 197.410 ;
        RECT 21.375 197.960 21.545 198.130 ;
        RECT 21.375 197.600 21.545 197.770 ;
        RECT 21.375 197.240 21.545 197.410 ;
        RECT 22.335 197.960 22.505 198.130 ;
        RECT 22.335 197.600 22.505 197.770 ;
        RECT 22.335 197.240 22.505 197.410 ;
        RECT 23.295 197.960 23.465 198.130 ;
        RECT 23.295 197.600 23.465 197.770 ;
        RECT 23.295 197.240 23.465 197.410 ;
        RECT 24.255 197.960 24.425 198.130 ;
        RECT 24.255 197.600 24.425 197.770 ;
        RECT 24.255 197.240 24.425 197.410 ;
        RECT 26.740 195.880 26.910 196.050 ;
        RECT 1.565 195.100 1.735 195.270 ;
        RECT 2.525 195.100 2.695 195.270 ;
        RECT 3.485 195.100 3.655 195.270 ;
        RECT 4.445 195.100 4.615 195.270 ;
        RECT 5.405 195.100 5.575 195.270 ;
        RECT 6.365 195.100 6.535 195.270 ;
        RECT 12.330 195.120 12.500 195.290 ;
        RECT 12.810 195.120 12.980 195.290 ;
        RECT 13.290 195.120 13.460 195.290 ;
        RECT 13.770 195.120 13.940 195.290 ;
        RECT 14.250 195.120 14.420 195.290 ;
        RECT 14.730 195.120 14.900 195.290 ;
        RECT 15.210 195.120 15.380 195.290 ;
        RECT 15.690 195.120 15.860 195.290 ;
        RECT 16.170 195.120 16.340 195.290 ;
        RECT 16.650 195.120 16.820 195.290 ;
        RECT 17.130 195.120 17.300 195.290 ;
        RECT 18.675 195.045 18.845 195.425 ;
        RECT 20.415 195.120 20.585 195.290 ;
        RECT 21.375 195.120 21.545 195.290 ;
        RECT 22.335 195.120 22.505 195.290 ;
        RECT 23.295 195.120 23.465 195.290 ;
        RECT 24.255 195.120 24.425 195.290 ;
        RECT 12.330 194.565 12.500 194.735 ;
        RECT 13.290 194.565 13.460 194.735 ;
        RECT 14.250 194.565 14.420 194.735 ;
        RECT 15.210 194.565 15.380 194.735 ;
        RECT 16.170 194.565 16.340 194.735 ;
        RECT 17.130 194.565 17.300 194.735 ;
        RECT 19.935 194.565 20.105 194.735 ;
        RECT 20.895 194.565 21.065 194.735 ;
        RECT 21.855 194.565 22.025 194.735 ;
        RECT 22.815 194.565 22.985 194.735 ;
        RECT 23.775 194.565 23.945 194.735 ;
        RECT 24.735 194.565 24.905 194.735 ;
        RECT 1.565 191.505 1.735 191.675 ;
        RECT 1.565 191.145 1.735 191.315 ;
        RECT 1.565 190.785 1.735 190.955 ;
        RECT 2.525 191.505 2.695 191.675 ;
        RECT 2.525 191.145 2.695 191.315 ;
        RECT 2.525 190.785 2.695 190.955 ;
        RECT 3.485 191.505 3.655 191.675 ;
        RECT 3.485 191.145 3.655 191.315 ;
        RECT 3.485 190.785 3.655 190.955 ;
        RECT 4.445 191.505 4.615 191.675 ;
        RECT 4.445 191.145 4.615 191.315 ;
        RECT 4.445 190.785 4.615 190.955 ;
        RECT 5.405 191.505 5.575 191.675 ;
        RECT 5.405 191.145 5.575 191.315 ;
        RECT 5.405 190.785 5.575 190.955 ;
        RECT 6.365 191.505 6.535 191.675 ;
        RECT 6.365 191.145 6.535 191.315 ;
        RECT 6.365 190.785 6.535 190.955 ;
        RECT 12.330 191.525 12.500 191.695 ;
        RECT 12.330 191.165 12.500 191.335 ;
        RECT 12.330 190.805 12.500 190.975 ;
        RECT 12.810 191.525 12.980 191.695 ;
        RECT 12.810 191.165 12.980 191.335 ;
        RECT 12.810 190.805 12.980 190.975 ;
        RECT 13.290 191.525 13.460 191.695 ;
        RECT 13.290 191.165 13.460 191.335 ;
        RECT 13.290 190.805 13.460 190.975 ;
        RECT 13.770 191.525 13.940 191.695 ;
        RECT 13.770 191.165 13.940 191.335 ;
        RECT 13.770 190.805 13.940 190.975 ;
        RECT 14.250 191.525 14.420 191.695 ;
        RECT 14.250 191.165 14.420 191.335 ;
        RECT 14.250 190.805 14.420 190.975 ;
        RECT 14.730 191.525 14.900 191.695 ;
        RECT 14.730 191.165 14.900 191.335 ;
        RECT 14.730 190.805 14.900 190.975 ;
        RECT 15.210 191.525 15.380 191.695 ;
        RECT 15.210 191.165 15.380 191.335 ;
        RECT 15.210 190.805 15.380 190.975 ;
        RECT 15.690 191.525 15.860 191.695 ;
        RECT 15.690 191.165 15.860 191.335 ;
        RECT 15.690 190.805 15.860 190.975 ;
        RECT 16.170 191.525 16.340 191.695 ;
        RECT 16.170 191.165 16.340 191.335 ;
        RECT 16.170 190.805 16.340 190.975 ;
        RECT 16.650 191.525 16.820 191.695 ;
        RECT 16.650 191.165 16.820 191.335 ;
        RECT 16.650 190.805 16.820 190.975 ;
        RECT 17.130 191.525 17.300 191.695 ;
        RECT 17.130 191.165 17.300 191.335 ;
        RECT 17.130 190.805 17.300 190.975 ;
        RECT 20.415 191.525 20.585 191.695 ;
        RECT 20.415 191.165 20.585 191.335 ;
        RECT 20.415 190.805 20.585 190.975 ;
        RECT 21.375 191.525 21.545 191.695 ;
        RECT 21.375 191.165 21.545 191.335 ;
        RECT 21.375 190.805 21.545 190.975 ;
        RECT 22.335 191.525 22.505 191.695 ;
        RECT 22.335 191.165 22.505 191.335 ;
        RECT 22.335 190.805 22.505 190.975 ;
        RECT 23.295 191.525 23.465 191.695 ;
        RECT 23.295 191.165 23.465 191.335 ;
        RECT 23.295 190.805 23.465 190.975 ;
        RECT 24.255 191.525 24.425 191.695 ;
        RECT 24.255 191.165 24.425 191.335 ;
        RECT 24.255 190.805 24.425 190.975 ;
        RECT 26.740 189.445 26.910 189.615 ;
        RECT 1.565 188.665 1.735 188.835 ;
        RECT 2.525 188.665 2.695 188.835 ;
        RECT 3.485 188.665 3.655 188.835 ;
        RECT 4.445 188.665 4.615 188.835 ;
        RECT 5.405 188.665 5.575 188.835 ;
        RECT 6.365 188.665 6.535 188.835 ;
        RECT 12.330 188.685 12.500 188.855 ;
        RECT 12.810 188.685 12.980 188.855 ;
        RECT 13.290 188.685 13.460 188.855 ;
        RECT 13.770 188.685 13.940 188.855 ;
        RECT 14.250 188.685 14.420 188.855 ;
        RECT 14.730 188.685 14.900 188.855 ;
        RECT 15.210 188.685 15.380 188.855 ;
        RECT 15.690 188.685 15.860 188.855 ;
        RECT 16.170 188.685 16.340 188.855 ;
        RECT 16.650 188.685 16.820 188.855 ;
        RECT 17.130 188.685 17.300 188.855 ;
        RECT 18.675 188.610 18.845 188.990 ;
        RECT 20.415 188.685 20.585 188.855 ;
        RECT 21.375 188.685 21.545 188.855 ;
        RECT 22.335 188.685 22.505 188.855 ;
        RECT 23.295 188.685 23.465 188.855 ;
        RECT 24.255 188.685 24.425 188.855 ;
        RECT 12.330 188.130 12.500 188.300 ;
        RECT 13.290 188.130 13.460 188.300 ;
        RECT 14.250 188.130 14.420 188.300 ;
        RECT 15.210 188.130 15.380 188.300 ;
        RECT 16.170 188.130 16.340 188.300 ;
        RECT 17.130 188.130 17.300 188.300 ;
        RECT 19.935 188.130 20.105 188.300 ;
        RECT 20.895 188.130 21.065 188.300 ;
        RECT 21.855 188.130 22.025 188.300 ;
        RECT 22.815 188.130 22.985 188.300 ;
        RECT 23.775 188.130 23.945 188.300 ;
        RECT 24.735 188.130 24.905 188.300 ;
        RECT 1.565 185.070 1.735 185.240 ;
        RECT 1.565 184.710 1.735 184.880 ;
        RECT 1.565 184.350 1.735 184.520 ;
        RECT 2.525 185.070 2.695 185.240 ;
        RECT 2.525 184.710 2.695 184.880 ;
        RECT 2.525 184.350 2.695 184.520 ;
        RECT 3.485 185.070 3.655 185.240 ;
        RECT 3.485 184.710 3.655 184.880 ;
        RECT 3.485 184.350 3.655 184.520 ;
        RECT 4.445 185.070 4.615 185.240 ;
        RECT 4.445 184.710 4.615 184.880 ;
        RECT 4.445 184.350 4.615 184.520 ;
        RECT 5.405 185.070 5.575 185.240 ;
        RECT 5.405 184.710 5.575 184.880 ;
        RECT 5.405 184.350 5.575 184.520 ;
        RECT 6.365 185.070 6.535 185.240 ;
        RECT 6.365 184.710 6.535 184.880 ;
        RECT 6.365 184.350 6.535 184.520 ;
        RECT 12.330 185.090 12.500 185.260 ;
        RECT 12.330 184.730 12.500 184.900 ;
        RECT 12.330 184.370 12.500 184.540 ;
        RECT 12.810 185.090 12.980 185.260 ;
        RECT 12.810 184.730 12.980 184.900 ;
        RECT 12.810 184.370 12.980 184.540 ;
        RECT 13.290 185.090 13.460 185.260 ;
        RECT 13.290 184.730 13.460 184.900 ;
        RECT 13.290 184.370 13.460 184.540 ;
        RECT 13.770 185.090 13.940 185.260 ;
        RECT 13.770 184.730 13.940 184.900 ;
        RECT 13.770 184.370 13.940 184.540 ;
        RECT 14.250 185.090 14.420 185.260 ;
        RECT 14.250 184.730 14.420 184.900 ;
        RECT 14.250 184.370 14.420 184.540 ;
        RECT 14.730 185.090 14.900 185.260 ;
        RECT 14.730 184.730 14.900 184.900 ;
        RECT 14.730 184.370 14.900 184.540 ;
        RECT 15.210 185.090 15.380 185.260 ;
        RECT 15.210 184.730 15.380 184.900 ;
        RECT 15.210 184.370 15.380 184.540 ;
        RECT 15.690 185.090 15.860 185.260 ;
        RECT 15.690 184.730 15.860 184.900 ;
        RECT 15.690 184.370 15.860 184.540 ;
        RECT 16.170 185.090 16.340 185.260 ;
        RECT 16.170 184.730 16.340 184.900 ;
        RECT 16.170 184.370 16.340 184.540 ;
        RECT 16.650 185.090 16.820 185.260 ;
        RECT 16.650 184.730 16.820 184.900 ;
        RECT 16.650 184.370 16.820 184.540 ;
        RECT 17.130 185.090 17.300 185.260 ;
        RECT 17.130 184.730 17.300 184.900 ;
        RECT 17.130 184.370 17.300 184.540 ;
        RECT 20.415 185.090 20.585 185.260 ;
        RECT 20.415 184.730 20.585 184.900 ;
        RECT 20.415 184.370 20.585 184.540 ;
        RECT 21.375 185.090 21.545 185.260 ;
        RECT 21.375 184.730 21.545 184.900 ;
        RECT 21.375 184.370 21.545 184.540 ;
        RECT 22.335 185.090 22.505 185.260 ;
        RECT 22.335 184.730 22.505 184.900 ;
        RECT 22.335 184.370 22.505 184.540 ;
        RECT 23.295 185.090 23.465 185.260 ;
        RECT 23.295 184.730 23.465 184.900 ;
        RECT 23.295 184.370 23.465 184.540 ;
        RECT 24.255 185.090 24.425 185.260 ;
        RECT 24.255 184.730 24.425 184.900 ;
        RECT 24.255 184.370 24.425 184.540 ;
        RECT 26.740 183.010 26.910 183.180 ;
        RECT 1.565 182.230 1.735 182.400 ;
        RECT 2.525 182.230 2.695 182.400 ;
        RECT 3.485 182.230 3.655 182.400 ;
        RECT 4.445 182.230 4.615 182.400 ;
        RECT 5.405 182.230 5.575 182.400 ;
        RECT 6.365 182.230 6.535 182.400 ;
        RECT 12.330 182.250 12.500 182.420 ;
        RECT 12.810 182.250 12.980 182.420 ;
        RECT 13.290 182.250 13.460 182.420 ;
        RECT 13.770 182.250 13.940 182.420 ;
        RECT 14.250 182.250 14.420 182.420 ;
        RECT 14.730 182.250 14.900 182.420 ;
        RECT 15.210 182.250 15.380 182.420 ;
        RECT 15.690 182.250 15.860 182.420 ;
        RECT 16.170 182.250 16.340 182.420 ;
        RECT 16.650 182.250 16.820 182.420 ;
        RECT 17.130 182.250 17.300 182.420 ;
        RECT 18.675 182.175 18.845 182.555 ;
        RECT 20.415 182.250 20.585 182.420 ;
        RECT 21.375 182.250 21.545 182.420 ;
        RECT 22.335 182.250 22.505 182.420 ;
        RECT 23.295 182.250 23.465 182.420 ;
        RECT 24.255 182.250 24.425 182.420 ;
        RECT 12.330 181.695 12.500 181.865 ;
        RECT 13.290 181.695 13.460 181.865 ;
        RECT 14.250 181.695 14.420 181.865 ;
        RECT 15.210 181.695 15.380 181.865 ;
        RECT 16.170 181.695 16.340 181.865 ;
        RECT 17.130 181.695 17.300 181.865 ;
        RECT 19.935 181.695 20.105 181.865 ;
        RECT 20.895 181.695 21.065 181.865 ;
        RECT 21.855 181.695 22.025 181.865 ;
        RECT 22.815 181.695 22.985 181.865 ;
        RECT 23.775 181.695 23.945 181.865 ;
        RECT 24.735 181.695 24.905 181.865 ;
        RECT 1.565 178.635 1.735 178.805 ;
        RECT 1.565 178.275 1.735 178.445 ;
        RECT 1.565 177.915 1.735 178.085 ;
        RECT 2.525 178.635 2.695 178.805 ;
        RECT 2.525 178.275 2.695 178.445 ;
        RECT 2.525 177.915 2.695 178.085 ;
        RECT 3.485 178.635 3.655 178.805 ;
        RECT 3.485 178.275 3.655 178.445 ;
        RECT 3.485 177.915 3.655 178.085 ;
        RECT 4.445 178.635 4.615 178.805 ;
        RECT 4.445 178.275 4.615 178.445 ;
        RECT 4.445 177.915 4.615 178.085 ;
        RECT 5.405 178.635 5.575 178.805 ;
        RECT 5.405 178.275 5.575 178.445 ;
        RECT 5.405 177.915 5.575 178.085 ;
        RECT 6.365 178.635 6.535 178.805 ;
        RECT 6.365 178.275 6.535 178.445 ;
        RECT 6.365 177.915 6.535 178.085 ;
        RECT 12.330 178.655 12.500 178.825 ;
        RECT 12.330 178.295 12.500 178.465 ;
        RECT 12.330 177.935 12.500 178.105 ;
        RECT 12.810 178.655 12.980 178.825 ;
        RECT 12.810 178.295 12.980 178.465 ;
        RECT 12.810 177.935 12.980 178.105 ;
        RECT 13.290 178.655 13.460 178.825 ;
        RECT 13.290 178.295 13.460 178.465 ;
        RECT 13.290 177.935 13.460 178.105 ;
        RECT 13.770 178.655 13.940 178.825 ;
        RECT 13.770 178.295 13.940 178.465 ;
        RECT 13.770 177.935 13.940 178.105 ;
        RECT 14.250 178.655 14.420 178.825 ;
        RECT 14.250 178.295 14.420 178.465 ;
        RECT 14.250 177.935 14.420 178.105 ;
        RECT 14.730 178.655 14.900 178.825 ;
        RECT 14.730 178.295 14.900 178.465 ;
        RECT 14.730 177.935 14.900 178.105 ;
        RECT 15.210 178.655 15.380 178.825 ;
        RECT 15.210 178.295 15.380 178.465 ;
        RECT 15.210 177.935 15.380 178.105 ;
        RECT 15.690 178.655 15.860 178.825 ;
        RECT 15.690 178.295 15.860 178.465 ;
        RECT 15.690 177.935 15.860 178.105 ;
        RECT 16.170 178.655 16.340 178.825 ;
        RECT 16.170 178.295 16.340 178.465 ;
        RECT 16.170 177.935 16.340 178.105 ;
        RECT 16.650 178.655 16.820 178.825 ;
        RECT 16.650 178.295 16.820 178.465 ;
        RECT 16.650 177.935 16.820 178.105 ;
        RECT 17.130 178.655 17.300 178.825 ;
        RECT 17.130 178.295 17.300 178.465 ;
        RECT 17.130 177.935 17.300 178.105 ;
        RECT 20.415 178.655 20.585 178.825 ;
        RECT 20.415 178.295 20.585 178.465 ;
        RECT 20.415 177.935 20.585 178.105 ;
        RECT 21.375 178.655 21.545 178.825 ;
        RECT 21.375 178.295 21.545 178.465 ;
        RECT 21.375 177.935 21.545 178.105 ;
        RECT 22.335 178.655 22.505 178.825 ;
        RECT 22.335 178.295 22.505 178.465 ;
        RECT 22.335 177.935 22.505 178.105 ;
        RECT 23.295 178.655 23.465 178.825 ;
        RECT 23.295 178.295 23.465 178.465 ;
        RECT 23.295 177.935 23.465 178.105 ;
        RECT 24.255 178.655 24.425 178.825 ;
        RECT 24.255 178.295 24.425 178.465 ;
        RECT 24.255 177.935 24.425 178.105 ;
        RECT 26.740 176.575 26.910 176.745 ;
        RECT 1.565 175.795 1.735 175.965 ;
        RECT 2.525 175.795 2.695 175.965 ;
        RECT 3.485 175.795 3.655 175.965 ;
        RECT 4.445 175.795 4.615 175.965 ;
        RECT 5.405 175.795 5.575 175.965 ;
        RECT 6.365 175.795 6.535 175.965 ;
        RECT 12.330 175.815 12.500 175.985 ;
        RECT 12.810 175.815 12.980 175.985 ;
        RECT 13.290 175.815 13.460 175.985 ;
        RECT 13.770 175.815 13.940 175.985 ;
        RECT 14.250 175.815 14.420 175.985 ;
        RECT 14.730 175.815 14.900 175.985 ;
        RECT 15.210 175.815 15.380 175.985 ;
        RECT 15.690 175.815 15.860 175.985 ;
        RECT 16.170 175.815 16.340 175.985 ;
        RECT 16.650 175.815 16.820 175.985 ;
        RECT 17.130 175.815 17.300 175.985 ;
        RECT 18.675 175.740 18.845 176.120 ;
        RECT 20.415 175.815 20.585 175.985 ;
        RECT 21.375 175.815 21.545 175.985 ;
        RECT 22.335 175.815 22.505 175.985 ;
        RECT 23.295 175.815 23.465 175.985 ;
        RECT 24.255 175.815 24.425 175.985 ;
        RECT 12.330 175.260 12.500 175.430 ;
        RECT 13.290 175.260 13.460 175.430 ;
        RECT 14.250 175.260 14.420 175.430 ;
        RECT 15.210 175.260 15.380 175.430 ;
        RECT 16.170 175.260 16.340 175.430 ;
        RECT 17.130 175.260 17.300 175.430 ;
        RECT 19.935 175.260 20.105 175.430 ;
        RECT 20.895 175.260 21.065 175.430 ;
        RECT 21.855 175.260 22.025 175.430 ;
        RECT 22.815 175.260 22.985 175.430 ;
        RECT 23.775 175.260 23.945 175.430 ;
        RECT 24.735 175.260 24.905 175.430 ;
        RECT 1.565 172.200 1.735 172.370 ;
        RECT 1.565 171.840 1.735 172.010 ;
        RECT 1.565 171.480 1.735 171.650 ;
        RECT 2.525 172.200 2.695 172.370 ;
        RECT 2.525 171.840 2.695 172.010 ;
        RECT 2.525 171.480 2.695 171.650 ;
        RECT 3.485 172.200 3.655 172.370 ;
        RECT 3.485 171.840 3.655 172.010 ;
        RECT 3.485 171.480 3.655 171.650 ;
        RECT 4.445 172.200 4.615 172.370 ;
        RECT 4.445 171.840 4.615 172.010 ;
        RECT 4.445 171.480 4.615 171.650 ;
        RECT 5.405 172.200 5.575 172.370 ;
        RECT 5.405 171.840 5.575 172.010 ;
        RECT 5.405 171.480 5.575 171.650 ;
        RECT 6.365 172.200 6.535 172.370 ;
        RECT 6.365 171.840 6.535 172.010 ;
        RECT 6.365 171.480 6.535 171.650 ;
        RECT 12.330 172.220 12.500 172.390 ;
        RECT 12.330 171.860 12.500 172.030 ;
        RECT 12.330 171.500 12.500 171.670 ;
        RECT 12.810 172.220 12.980 172.390 ;
        RECT 12.810 171.860 12.980 172.030 ;
        RECT 12.810 171.500 12.980 171.670 ;
        RECT 13.290 172.220 13.460 172.390 ;
        RECT 13.290 171.860 13.460 172.030 ;
        RECT 13.290 171.500 13.460 171.670 ;
        RECT 13.770 172.220 13.940 172.390 ;
        RECT 13.770 171.860 13.940 172.030 ;
        RECT 13.770 171.500 13.940 171.670 ;
        RECT 14.250 172.220 14.420 172.390 ;
        RECT 14.250 171.860 14.420 172.030 ;
        RECT 14.250 171.500 14.420 171.670 ;
        RECT 14.730 172.220 14.900 172.390 ;
        RECT 14.730 171.860 14.900 172.030 ;
        RECT 14.730 171.500 14.900 171.670 ;
        RECT 15.210 172.220 15.380 172.390 ;
        RECT 15.210 171.860 15.380 172.030 ;
        RECT 15.210 171.500 15.380 171.670 ;
        RECT 15.690 172.220 15.860 172.390 ;
        RECT 15.690 171.860 15.860 172.030 ;
        RECT 15.690 171.500 15.860 171.670 ;
        RECT 16.170 172.220 16.340 172.390 ;
        RECT 16.170 171.860 16.340 172.030 ;
        RECT 16.170 171.500 16.340 171.670 ;
        RECT 16.650 172.220 16.820 172.390 ;
        RECT 16.650 171.860 16.820 172.030 ;
        RECT 16.650 171.500 16.820 171.670 ;
        RECT 17.130 172.220 17.300 172.390 ;
        RECT 17.130 171.860 17.300 172.030 ;
        RECT 17.130 171.500 17.300 171.670 ;
        RECT 20.415 172.220 20.585 172.390 ;
        RECT 20.415 171.860 20.585 172.030 ;
        RECT 20.415 171.500 20.585 171.670 ;
        RECT 21.375 172.220 21.545 172.390 ;
        RECT 21.375 171.860 21.545 172.030 ;
        RECT 21.375 171.500 21.545 171.670 ;
        RECT 22.335 172.220 22.505 172.390 ;
        RECT 22.335 171.860 22.505 172.030 ;
        RECT 22.335 171.500 22.505 171.670 ;
        RECT 23.295 172.220 23.465 172.390 ;
        RECT 23.295 171.860 23.465 172.030 ;
        RECT 23.295 171.500 23.465 171.670 ;
        RECT 24.255 172.220 24.425 172.390 ;
        RECT 24.255 171.860 24.425 172.030 ;
        RECT 24.255 171.500 24.425 171.670 ;
        RECT 26.740 170.140 26.910 170.310 ;
        RECT 1.565 169.360 1.735 169.530 ;
        RECT 2.525 169.360 2.695 169.530 ;
        RECT 3.485 169.360 3.655 169.530 ;
        RECT 4.445 169.360 4.615 169.530 ;
        RECT 5.405 169.360 5.575 169.530 ;
        RECT 6.365 169.360 6.535 169.530 ;
        RECT 12.330 169.380 12.500 169.550 ;
        RECT 12.810 169.380 12.980 169.550 ;
        RECT 13.290 169.380 13.460 169.550 ;
        RECT 13.770 169.380 13.940 169.550 ;
        RECT 14.250 169.380 14.420 169.550 ;
        RECT 14.730 169.380 14.900 169.550 ;
        RECT 15.210 169.380 15.380 169.550 ;
        RECT 15.690 169.380 15.860 169.550 ;
        RECT 16.170 169.380 16.340 169.550 ;
        RECT 16.650 169.380 16.820 169.550 ;
        RECT 17.130 169.380 17.300 169.550 ;
        RECT 18.675 169.305 18.845 169.685 ;
        RECT 20.415 169.380 20.585 169.550 ;
        RECT 21.375 169.380 21.545 169.550 ;
        RECT 22.335 169.380 22.505 169.550 ;
        RECT 23.295 169.380 23.465 169.550 ;
        RECT 24.255 169.380 24.425 169.550 ;
        RECT 12.330 168.825 12.500 168.995 ;
        RECT 13.290 168.825 13.460 168.995 ;
        RECT 14.250 168.825 14.420 168.995 ;
        RECT 15.210 168.825 15.380 168.995 ;
        RECT 16.170 168.825 16.340 168.995 ;
        RECT 17.130 168.825 17.300 168.995 ;
        RECT 19.935 168.825 20.105 168.995 ;
        RECT 20.895 168.825 21.065 168.995 ;
        RECT 21.855 168.825 22.025 168.995 ;
        RECT 22.815 168.825 22.985 168.995 ;
        RECT 23.775 168.825 23.945 168.995 ;
        RECT 24.735 168.825 24.905 168.995 ;
        RECT 1.565 165.765 1.735 165.935 ;
        RECT 1.565 165.405 1.735 165.575 ;
        RECT 1.565 165.045 1.735 165.215 ;
        RECT 2.525 165.765 2.695 165.935 ;
        RECT 2.525 165.405 2.695 165.575 ;
        RECT 2.525 165.045 2.695 165.215 ;
        RECT 3.485 165.765 3.655 165.935 ;
        RECT 3.485 165.405 3.655 165.575 ;
        RECT 3.485 165.045 3.655 165.215 ;
        RECT 4.445 165.765 4.615 165.935 ;
        RECT 4.445 165.405 4.615 165.575 ;
        RECT 4.445 165.045 4.615 165.215 ;
        RECT 5.405 165.765 5.575 165.935 ;
        RECT 5.405 165.405 5.575 165.575 ;
        RECT 5.405 165.045 5.575 165.215 ;
        RECT 6.365 165.765 6.535 165.935 ;
        RECT 6.365 165.405 6.535 165.575 ;
        RECT 6.365 165.045 6.535 165.215 ;
        RECT 12.330 165.785 12.500 165.955 ;
        RECT 12.330 165.425 12.500 165.595 ;
        RECT 12.330 165.065 12.500 165.235 ;
        RECT 12.810 165.785 12.980 165.955 ;
        RECT 12.810 165.425 12.980 165.595 ;
        RECT 12.810 165.065 12.980 165.235 ;
        RECT 13.290 165.785 13.460 165.955 ;
        RECT 13.290 165.425 13.460 165.595 ;
        RECT 13.290 165.065 13.460 165.235 ;
        RECT 13.770 165.785 13.940 165.955 ;
        RECT 13.770 165.425 13.940 165.595 ;
        RECT 13.770 165.065 13.940 165.235 ;
        RECT 14.250 165.785 14.420 165.955 ;
        RECT 14.250 165.425 14.420 165.595 ;
        RECT 14.250 165.065 14.420 165.235 ;
        RECT 14.730 165.785 14.900 165.955 ;
        RECT 14.730 165.425 14.900 165.595 ;
        RECT 14.730 165.065 14.900 165.235 ;
        RECT 15.210 165.785 15.380 165.955 ;
        RECT 15.210 165.425 15.380 165.595 ;
        RECT 15.210 165.065 15.380 165.235 ;
        RECT 15.690 165.785 15.860 165.955 ;
        RECT 15.690 165.425 15.860 165.595 ;
        RECT 15.690 165.065 15.860 165.235 ;
        RECT 16.170 165.785 16.340 165.955 ;
        RECT 16.170 165.425 16.340 165.595 ;
        RECT 16.170 165.065 16.340 165.235 ;
        RECT 16.650 165.785 16.820 165.955 ;
        RECT 16.650 165.425 16.820 165.595 ;
        RECT 16.650 165.065 16.820 165.235 ;
        RECT 17.130 165.785 17.300 165.955 ;
        RECT 17.130 165.425 17.300 165.595 ;
        RECT 17.130 165.065 17.300 165.235 ;
        RECT 20.415 165.785 20.585 165.955 ;
        RECT 20.415 165.425 20.585 165.595 ;
        RECT 20.415 165.065 20.585 165.235 ;
        RECT 21.375 165.785 21.545 165.955 ;
        RECT 21.375 165.425 21.545 165.595 ;
        RECT 21.375 165.065 21.545 165.235 ;
        RECT 22.335 165.785 22.505 165.955 ;
        RECT 22.335 165.425 22.505 165.595 ;
        RECT 22.335 165.065 22.505 165.235 ;
        RECT 23.295 165.785 23.465 165.955 ;
        RECT 23.295 165.425 23.465 165.595 ;
        RECT 23.295 165.065 23.465 165.235 ;
        RECT 24.255 165.785 24.425 165.955 ;
        RECT 24.255 165.425 24.425 165.595 ;
        RECT 24.255 165.065 24.425 165.235 ;
        RECT 26.740 163.705 26.910 163.875 ;
        RECT 1.565 162.925 1.735 163.095 ;
        RECT 2.525 162.925 2.695 163.095 ;
        RECT 3.485 162.925 3.655 163.095 ;
        RECT 4.445 162.925 4.615 163.095 ;
        RECT 5.405 162.925 5.575 163.095 ;
        RECT 6.365 162.925 6.535 163.095 ;
        RECT 12.330 162.945 12.500 163.115 ;
        RECT 12.810 162.945 12.980 163.115 ;
        RECT 13.290 162.945 13.460 163.115 ;
        RECT 13.770 162.945 13.940 163.115 ;
        RECT 14.250 162.945 14.420 163.115 ;
        RECT 14.730 162.945 14.900 163.115 ;
        RECT 15.210 162.945 15.380 163.115 ;
        RECT 15.690 162.945 15.860 163.115 ;
        RECT 16.170 162.945 16.340 163.115 ;
        RECT 16.650 162.945 16.820 163.115 ;
        RECT 17.130 162.945 17.300 163.115 ;
        RECT 18.675 162.870 18.845 163.250 ;
        RECT 20.415 162.945 20.585 163.115 ;
        RECT 21.375 162.945 21.545 163.115 ;
        RECT 22.335 162.945 22.505 163.115 ;
        RECT 23.295 162.945 23.465 163.115 ;
        RECT 24.255 162.945 24.425 163.115 ;
        RECT 12.330 162.390 12.500 162.560 ;
        RECT 13.290 162.390 13.460 162.560 ;
        RECT 14.250 162.390 14.420 162.560 ;
        RECT 15.210 162.390 15.380 162.560 ;
        RECT 16.170 162.390 16.340 162.560 ;
        RECT 17.130 162.390 17.300 162.560 ;
        RECT 19.935 162.390 20.105 162.560 ;
        RECT 20.895 162.390 21.065 162.560 ;
        RECT 21.855 162.390 22.025 162.560 ;
        RECT 22.815 162.390 22.985 162.560 ;
        RECT 23.775 162.390 23.945 162.560 ;
        RECT 24.735 162.390 24.905 162.560 ;
        RECT 1.565 159.330 1.735 159.500 ;
        RECT 1.565 158.970 1.735 159.140 ;
        RECT 1.565 158.610 1.735 158.780 ;
        RECT 2.525 159.330 2.695 159.500 ;
        RECT 2.525 158.970 2.695 159.140 ;
        RECT 2.525 158.610 2.695 158.780 ;
        RECT 3.485 159.330 3.655 159.500 ;
        RECT 3.485 158.970 3.655 159.140 ;
        RECT 3.485 158.610 3.655 158.780 ;
        RECT 4.445 159.330 4.615 159.500 ;
        RECT 4.445 158.970 4.615 159.140 ;
        RECT 4.445 158.610 4.615 158.780 ;
        RECT 5.405 159.330 5.575 159.500 ;
        RECT 5.405 158.970 5.575 159.140 ;
        RECT 5.405 158.610 5.575 158.780 ;
        RECT 6.365 159.330 6.535 159.500 ;
        RECT 6.365 158.970 6.535 159.140 ;
        RECT 6.365 158.610 6.535 158.780 ;
        RECT 12.330 159.350 12.500 159.520 ;
        RECT 12.330 158.990 12.500 159.160 ;
        RECT 12.330 158.630 12.500 158.800 ;
        RECT 12.810 159.350 12.980 159.520 ;
        RECT 12.810 158.990 12.980 159.160 ;
        RECT 12.810 158.630 12.980 158.800 ;
        RECT 13.290 159.350 13.460 159.520 ;
        RECT 13.290 158.990 13.460 159.160 ;
        RECT 13.290 158.630 13.460 158.800 ;
        RECT 13.770 159.350 13.940 159.520 ;
        RECT 13.770 158.990 13.940 159.160 ;
        RECT 13.770 158.630 13.940 158.800 ;
        RECT 14.250 159.350 14.420 159.520 ;
        RECT 14.250 158.990 14.420 159.160 ;
        RECT 14.250 158.630 14.420 158.800 ;
        RECT 14.730 159.350 14.900 159.520 ;
        RECT 14.730 158.990 14.900 159.160 ;
        RECT 14.730 158.630 14.900 158.800 ;
        RECT 15.210 159.350 15.380 159.520 ;
        RECT 15.210 158.990 15.380 159.160 ;
        RECT 15.210 158.630 15.380 158.800 ;
        RECT 15.690 159.350 15.860 159.520 ;
        RECT 15.690 158.990 15.860 159.160 ;
        RECT 15.690 158.630 15.860 158.800 ;
        RECT 16.170 159.350 16.340 159.520 ;
        RECT 16.170 158.990 16.340 159.160 ;
        RECT 16.170 158.630 16.340 158.800 ;
        RECT 16.650 159.350 16.820 159.520 ;
        RECT 16.650 158.990 16.820 159.160 ;
        RECT 16.650 158.630 16.820 158.800 ;
        RECT 17.130 159.350 17.300 159.520 ;
        RECT 17.130 158.990 17.300 159.160 ;
        RECT 17.130 158.630 17.300 158.800 ;
        RECT 20.415 159.350 20.585 159.520 ;
        RECT 20.415 158.990 20.585 159.160 ;
        RECT 20.415 158.630 20.585 158.800 ;
        RECT 21.375 159.350 21.545 159.520 ;
        RECT 21.375 158.990 21.545 159.160 ;
        RECT 21.375 158.630 21.545 158.800 ;
        RECT 22.335 159.350 22.505 159.520 ;
        RECT 22.335 158.990 22.505 159.160 ;
        RECT 22.335 158.630 22.505 158.800 ;
        RECT 23.295 159.350 23.465 159.520 ;
        RECT 23.295 158.990 23.465 159.160 ;
        RECT 23.295 158.630 23.465 158.800 ;
        RECT 24.255 159.350 24.425 159.520 ;
        RECT 24.255 158.990 24.425 159.160 ;
        RECT 24.255 158.630 24.425 158.800 ;
        RECT 26.740 157.270 26.910 157.440 ;
        RECT 1.565 156.490 1.735 156.660 ;
        RECT 2.525 156.490 2.695 156.660 ;
        RECT 3.485 156.490 3.655 156.660 ;
        RECT 4.445 156.490 4.615 156.660 ;
        RECT 5.405 156.490 5.575 156.660 ;
        RECT 6.365 156.490 6.535 156.660 ;
        RECT 12.330 156.510 12.500 156.680 ;
        RECT 12.810 156.510 12.980 156.680 ;
        RECT 13.290 156.510 13.460 156.680 ;
        RECT 13.770 156.510 13.940 156.680 ;
        RECT 14.250 156.510 14.420 156.680 ;
        RECT 14.730 156.510 14.900 156.680 ;
        RECT 15.210 156.510 15.380 156.680 ;
        RECT 15.690 156.510 15.860 156.680 ;
        RECT 16.170 156.510 16.340 156.680 ;
        RECT 16.650 156.510 16.820 156.680 ;
        RECT 17.130 156.510 17.300 156.680 ;
        RECT 18.675 156.435 18.845 156.815 ;
        RECT 20.415 156.510 20.585 156.680 ;
        RECT 21.375 156.510 21.545 156.680 ;
        RECT 22.335 156.510 22.505 156.680 ;
        RECT 23.295 156.510 23.465 156.680 ;
        RECT 24.255 156.510 24.425 156.680 ;
        RECT 12.330 155.955 12.500 156.125 ;
        RECT 13.290 155.955 13.460 156.125 ;
        RECT 14.250 155.955 14.420 156.125 ;
        RECT 15.210 155.955 15.380 156.125 ;
        RECT 16.170 155.955 16.340 156.125 ;
        RECT 17.130 155.955 17.300 156.125 ;
        RECT 19.935 155.955 20.105 156.125 ;
        RECT 20.895 155.955 21.065 156.125 ;
        RECT 21.855 155.955 22.025 156.125 ;
        RECT 22.815 155.955 22.985 156.125 ;
        RECT 23.775 155.955 23.945 156.125 ;
        RECT 24.735 155.955 24.905 156.125 ;
        RECT 1.565 152.895 1.735 153.065 ;
        RECT 1.565 152.535 1.735 152.705 ;
        RECT 1.565 152.175 1.735 152.345 ;
        RECT 2.525 152.895 2.695 153.065 ;
        RECT 2.525 152.535 2.695 152.705 ;
        RECT 2.525 152.175 2.695 152.345 ;
        RECT 3.485 152.895 3.655 153.065 ;
        RECT 3.485 152.535 3.655 152.705 ;
        RECT 3.485 152.175 3.655 152.345 ;
        RECT 4.445 152.895 4.615 153.065 ;
        RECT 4.445 152.535 4.615 152.705 ;
        RECT 4.445 152.175 4.615 152.345 ;
        RECT 5.405 152.895 5.575 153.065 ;
        RECT 5.405 152.535 5.575 152.705 ;
        RECT 5.405 152.175 5.575 152.345 ;
        RECT 6.365 152.895 6.535 153.065 ;
        RECT 6.365 152.535 6.535 152.705 ;
        RECT 6.365 152.175 6.535 152.345 ;
        RECT 12.330 152.915 12.500 153.085 ;
        RECT 12.330 152.555 12.500 152.725 ;
        RECT 12.330 152.195 12.500 152.365 ;
        RECT 12.810 152.915 12.980 153.085 ;
        RECT 12.810 152.555 12.980 152.725 ;
        RECT 12.810 152.195 12.980 152.365 ;
        RECT 13.290 152.915 13.460 153.085 ;
        RECT 13.290 152.555 13.460 152.725 ;
        RECT 13.290 152.195 13.460 152.365 ;
        RECT 13.770 152.915 13.940 153.085 ;
        RECT 13.770 152.555 13.940 152.725 ;
        RECT 13.770 152.195 13.940 152.365 ;
        RECT 14.250 152.915 14.420 153.085 ;
        RECT 14.250 152.555 14.420 152.725 ;
        RECT 14.250 152.195 14.420 152.365 ;
        RECT 14.730 152.915 14.900 153.085 ;
        RECT 14.730 152.555 14.900 152.725 ;
        RECT 14.730 152.195 14.900 152.365 ;
        RECT 15.210 152.915 15.380 153.085 ;
        RECT 15.210 152.555 15.380 152.725 ;
        RECT 15.210 152.195 15.380 152.365 ;
        RECT 15.690 152.915 15.860 153.085 ;
        RECT 15.690 152.555 15.860 152.725 ;
        RECT 15.690 152.195 15.860 152.365 ;
        RECT 16.170 152.915 16.340 153.085 ;
        RECT 16.170 152.555 16.340 152.725 ;
        RECT 16.170 152.195 16.340 152.365 ;
        RECT 16.650 152.915 16.820 153.085 ;
        RECT 16.650 152.555 16.820 152.725 ;
        RECT 16.650 152.195 16.820 152.365 ;
        RECT 17.130 152.915 17.300 153.085 ;
        RECT 17.130 152.555 17.300 152.725 ;
        RECT 17.130 152.195 17.300 152.365 ;
        RECT 20.415 152.915 20.585 153.085 ;
        RECT 20.415 152.555 20.585 152.725 ;
        RECT 20.415 152.195 20.585 152.365 ;
        RECT 21.375 152.915 21.545 153.085 ;
        RECT 21.375 152.555 21.545 152.725 ;
        RECT 21.375 152.195 21.545 152.365 ;
        RECT 22.335 152.915 22.505 153.085 ;
        RECT 22.335 152.555 22.505 152.725 ;
        RECT 22.335 152.195 22.505 152.365 ;
        RECT 23.295 152.915 23.465 153.085 ;
        RECT 23.295 152.555 23.465 152.725 ;
        RECT 23.295 152.195 23.465 152.365 ;
        RECT 24.255 152.915 24.425 153.085 ;
        RECT 24.255 152.555 24.425 152.725 ;
        RECT 24.255 152.195 24.425 152.365 ;
        RECT 26.740 150.835 26.910 151.005 ;
        RECT 1.565 150.055 1.735 150.225 ;
        RECT 2.525 150.055 2.695 150.225 ;
        RECT 3.485 150.055 3.655 150.225 ;
        RECT 4.445 150.055 4.615 150.225 ;
        RECT 5.405 150.055 5.575 150.225 ;
        RECT 6.365 150.055 6.535 150.225 ;
        RECT 12.330 150.075 12.500 150.245 ;
        RECT 12.810 150.075 12.980 150.245 ;
        RECT 13.290 150.075 13.460 150.245 ;
        RECT 13.770 150.075 13.940 150.245 ;
        RECT 14.250 150.075 14.420 150.245 ;
        RECT 14.730 150.075 14.900 150.245 ;
        RECT 15.210 150.075 15.380 150.245 ;
        RECT 15.690 150.075 15.860 150.245 ;
        RECT 16.170 150.075 16.340 150.245 ;
        RECT 16.650 150.075 16.820 150.245 ;
        RECT 17.130 150.075 17.300 150.245 ;
        RECT 18.675 150.000 18.845 150.380 ;
        RECT 20.415 150.075 20.585 150.245 ;
        RECT 21.375 150.075 21.545 150.245 ;
        RECT 22.335 150.075 22.505 150.245 ;
        RECT 23.295 150.075 23.465 150.245 ;
        RECT 24.255 150.075 24.425 150.245 ;
        RECT 12.330 149.520 12.500 149.690 ;
        RECT 13.290 149.520 13.460 149.690 ;
        RECT 14.250 149.520 14.420 149.690 ;
        RECT 15.210 149.520 15.380 149.690 ;
        RECT 16.170 149.520 16.340 149.690 ;
        RECT 17.130 149.520 17.300 149.690 ;
        RECT 19.935 149.520 20.105 149.690 ;
        RECT 20.895 149.520 21.065 149.690 ;
        RECT 21.855 149.520 22.025 149.690 ;
        RECT 22.815 149.520 22.985 149.690 ;
        RECT 23.775 149.520 23.945 149.690 ;
        RECT 24.735 149.520 24.905 149.690 ;
        RECT 1.565 146.460 1.735 146.630 ;
        RECT 1.565 146.100 1.735 146.270 ;
        RECT 1.565 145.740 1.735 145.910 ;
        RECT 2.525 146.460 2.695 146.630 ;
        RECT 2.525 146.100 2.695 146.270 ;
        RECT 2.525 145.740 2.695 145.910 ;
        RECT 3.485 146.460 3.655 146.630 ;
        RECT 3.485 146.100 3.655 146.270 ;
        RECT 3.485 145.740 3.655 145.910 ;
        RECT 4.445 146.460 4.615 146.630 ;
        RECT 4.445 146.100 4.615 146.270 ;
        RECT 4.445 145.740 4.615 145.910 ;
        RECT 5.405 146.460 5.575 146.630 ;
        RECT 5.405 146.100 5.575 146.270 ;
        RECT 5.405 145.740 5.575 145.910 ;
        RECT 6.365 146.460 6.535 146.630 ;
        RECT 6.365 146.100 6.535 146.270 ;
        RECT 6.365 145.740 6.535 145.910 ;
        RECT 12.330 146.480 12.500 146.650 ;
        RECT 12.330 146.120 12.500 146.290 ;
        RECT 12.330 145.760 12.500 145.930 ;
        RECT 12.810 146.480 12.980 146.650 ;
        RECT 12.810 146.120 12.980 146.290 ;
        RECT 12.810 145.760 12.980 145.930 ;
        RECT 13.290 146.480 13.460 146.650 ;
        RECT 13.290 146.120 13.460 146.290 ;
        RECT 13.290 145.760 13.460 145.930 ;
        RECT 13.770 146.480 13.940 146.650 ;
        RECT 13.770 146.120 13.940 146.290 ;
        RECT 13.770 145.760 13.940 145.930 ;
        RECT 14.250 146.480 14.420 146.650 ;
        RECT 14.250 146.120 14.420 146.290 ;
        RECT 14.250 145.760 14.420 145.930 ;
        RECT 14.730 146.480 14.900 146.650 ;
        RECT 14.730 146.120 14.900 146.290 ;
        RECT 14.730 145.760 14.900 145.930 ;
        RECT 15.210 146.480 15.380 146.650 ;
        RECT 15.210 146.120 15.380 146.290 ;
        RECT 15.210 145.760 15.380 145.930 ;
        RECT 15.690 146.480 15.860 146.650 ;
        RECT 15.690 146.120 15.860 146.290 ;
        RECT 15.690 145.760 15.860 145.930 ;
        RECT 16.170 146.480 16.340 146.650 ;
        RECT 16.170 146.120 16.340 146.290 ;
        RECT 16.170 145.760 16.340 145.930 ;
        RECT 16.650 146.480 16.820 146.650 ;
        RECT 16.650 146.120 16.820 146.290 ;
        RECT 16.650 145.760 16.820 145.930 ;
        RECT 17.130 146.480 17.300 146.650 ;
        RECT 17.130 146.120 17.300 146.290 ;
        RECT 17.130 145.760 17.300 145.930 ;
        RECT 20.415 146.480 20.585 146.650 ;
        RECT 20.415 146.120 20.585 146.290 ;
        RECT 20.415 145.760 20.585 145.930 ;
        RECT 21.375 146.480 21.545 146.650 ;
        RECT 21.375 146.120 21.545 146.290 ;
        RECT 21.375 145.760 21.545 145.930 ;
        RECT 22.335 146.480 22.505 146.650 ;
        RECT 22.335 146.120 22.505 146.290 ;
        RECT 22.335 145.760 22.505 145.930 ;
        RECT 23.295 146.480 23.465 146.650 ;
        RECT 23.295 146.120 23.465 146.290 ;
        RECT 23.295 145.760 23.465 145.930 ;
        RECT 24.255 146.480 24.425 146.650 ;
        RECT 24.255 146.120 24.425 146.290 ;
        RECT 24.255 145.760 24.425 145.930 ;
        RECT 26.740 144.400 26.910 144.570 ;
        RECT 1.565 143.620 1.735 143.790 ;
        RECT 2.525 143.620 2.695 143.790 ;
        RECT 3.485 143.620 3.655 143.790 ;
        RECT 4.445 143.620 4.615 143.790 ;
        RECT 5.405 143.620 5.575 143.790 ;
        RECT 6.365 143.620 6.535 143.790 ;
        RECT 12.330 143.640 12.500 143.810 ;
        RECT 12.810 143.640 12.980 143.810 ;
        RECT 13.290 143.640 13.460 143.810 ;
        RECT 13.770 143.640 13.940 143.810 ;
        RECT 14.250 143.640 14.420 143.810 ;
        RECT 14.730 143.640 14.900 143.810 ;
        RECT 15.210 143.640 15.380 143.810 ;
        RECT 15.690 143.640 15.860 143.810 ;
        RECT 16.170 143.640 16.340 143.810 ;
        RECT 16.650 143.640 16.820 143.810 ;
        RECT 17.130 143.640 17.300 143.810 ;
        RECT 18.675 143.565 18.845 143.945 ;
        RECT 20.415 143.640 20.585 143.810 ;
        RECT 21.375 143.640 21.545 143.810 ;
        RECT 22.335 143.640 22.505 143.810 ;
        RECT 23.295 143.640 23.465 143.810 ;
        RECT 24.255 143.640 24.425 143.810 ;
        RECT 12.330 143.085 12.500 143.255 ;
        RECT 13.290 143.085 13.460 143.255 ;
        RECT 14.250 143.085 14.420 143.255 ;
        RECT 15.210 143.085 15.380 143.255 ;
        RECT 16.170 143.085 16.340 143.255 ;
        RECT 17.130 143.085 17.300 143.255 ;
        RECT 19.935 143.085 20.105 143.255 ;
        RECT 20.895 143.085 21.065 143.255 ;
        RECT 21.855 143.085 22.025 143.255 ;
        RECT 22.815 143.085 22.985 143.255 ;
        RECT 23.775 143.085 23.945 143.255 ;
        RECT 24.735 143.085 24.905 143.255 ;
        RECT 1.565 140.025 1.735 140.195 ;
        RECT 1.565 139.665 1.735 139.835 ;
        RECT 1.565 139.305 1.735 139.475 ;
        RECT 2.525 140.025 2.695 140.195 ;
        RECT 2.525 139.665 2.695 139.835 ;
        RECT 2.525 139.305 2.695 139.475 ;
        RECT 3.485 140.025 3.655 140.195 ;
        RECT 3.485 139.665 3.655 139.835 ;
        RECT 3.485 139.305 3.655 139.475 ;
        RECT 4.445 140.025 4.615 140.195 ;
        RECT 4.445 139.665 4.615 139.835 ;
        RECT 4.445 139.305 4.615 139.475 ;
        RECT 5.405 140.025 5.575 140.195 ;
        RECT 5.405 139.665 5.575 139.835 ;
        RECT 5.405 139.305 5.575 139.475 ;
        RECT 6.365 140.025 6.535 140.195 ;
        RECT 6.365 139.665 6.535 139.835 ;
        RECT 6.365 139.305 6.535 139.475 ;
        RECT 12.330 140.045 12.500 140.215 ;
        RECT 12.330 139.685 12.500 139.855 ;
        RECT 12.330 139.325 12.500 139.495 ;
        RECT 12.810 140.045 12.980 140.215 ;
        RECT 12.810 139.685 12.980 139.855 ;
        RECT 12.810 139.325 12.980 139.495 ;
        RECT 13.290 140.045 13.460 140.215 ;
        RECT 13.290 139.685 13.460 139.855 ;
        RECT 13.290 139.325 13.460 139.495 ;
        RECT 13.770 140.045 13.940 140.215 ;
        RECT 13.770 139.685 13.940 139.855 ;
        RECT 13.770 139.325 13.940 139.495 ;
        RECT 14.250 140.045 14.420 140.215 ;
        RECT 14.250 139.685 14.420 139.855 ;
        RECT 14.250 139.325 14.420 139.495 ;
        RECT 14.730 140.045 14.900 140.215 ;
        RECT 14.730 139.685 14.900 139.855 ;
        RECT 14.730 139.325 14.900 139.495 ;
        RECT 15.210 140.045 15.380 140.215 ;
        RECT 15.210 139.685 15.380 139.855 ;
        RECT 15.210 139.325 15.380 139.495 ;
        RECT 15.690 140.045 15.860 140.215 ;
        RECT 15.690 139.685 15.860 139.855 ;
        RECT 15.690 139.325 15.860 139.495 ;
        RECT 16.170 140.045 16.340 140.215 ;
        RECT 16.170 139.685 16.340 139.855 ;
        RECT 16.170 139.325 16.340 139.495 ;
        RECT 16.650 140.045 16.820 140.215 ;
        RECT 16.650 139.685 16.820 139.855 ;
        RECT 16.650 139.325 16.820 139.495 ;
        RECT 17.130 140.045 17.300 140.215 ;
        RECT 17.130 139.685 17.300 139.855 ;
        RECT 17.130 139.325 17.300 139.495 ;
        RECT 20.415 140.045 20.585 140.215 ;
        RECT 20.415 139.685 20.585 139.855 ;
        RECT 20.415 139.325 20.585 139.495 ;
        RECT 21.375 140.045 21.545 140.215 ;
        RECT 21.375 139.685 21.545 139.855 ;
        RECT 21.375 139.325 21.545 139.495 ;
        RECT 22.335 140.045 22.505 140.215 ;
        RECT 22.335 139.685 22.505 139.855 ;
        RECT 22.335 139.325 22.505 139.495 ;
        RECT 23.295 140.045 23.465 140.215 ;
        RECT 23.295 139.685 23.465 139.855 ;
        RECT 23.295 139.325 23.465 139.495 ;
        RECT 24.255 140.045 24.425 140.215 ;
        RECT 24.255 139.685 24.425 139.855 ;
        RECT 24.255 139.325 24.425 139.495 ;
        RECT 26.740 137.965 26.910 138.135 ;
        RECT 1.565 137.185 1.735 137.355 ;
        RECT 2.525 137.185 2.695 137.355 ;
        RECT 3.485 137.185 3.655 137.355 ;
        RECT 4.445 137.185 4.615 137.355 ;
        RECT 5.405 137.185 5.575 137.355 ;
        RECT 6.365 137.185 6.535 137.355 ;
        RECT 12.330 137.205 12.500 137.375 ;
        RECT 12.810 137.205 12.980 137.375 ;
        RECT 13.290 137.205 13.460 137.375 ;
        RECT 13.770 137.205 13.940 137.375 ;
        RECT 14.250 137.205 14.420 137.375 ;
        RECT 14.730 137.205 14.900 137.375 ;
        RECT 15.210 137.205 15.380 137.375 ;
        RECT 15.690 137.205 15.860 137.375 ;
        RECT 16.170 137.205 16.340 137.375 ;
        RECT 16.650 137.205 16.820 137.375 ;
        RECT 17.130 137.205 17.300 137.375 ;
        RECT 18.675 137.130 18.845 137.510 ;
        RECT 20.415 137.205 20.585 137.375 ;
        RECT 21.375 137.205 21.545 137.375 ;
        RECT 22.335 137.205 22.505 137.375 ;
        RECT 23.295 137.205 23.465 137.375 ;
        RECT 24.255 137.205 24.425 137.375 ;
        RECT 12.330 136.650 12.500 136.820 ;
        RECT 13.290 136.650 13.460 136.820 ;
        RECT 14.250 136.650 14.420 136.820 ;
        RECT 15.210 136.650 15.380 136.820 ;
        RECT 16.170 136.650 16.340 136.820 ;
        RECT 17.130 136.650 17.300 136.820 ;
        RECT 19.935 136.650 20.105 136.820 ;
        RECT 20.895 136.650 21.065 136.820 ;
        RECT 21.855 136.650 22.025 136.820 ;
        RECT 22.815 136.650 22.985 136.820 ;
        RECT 23.775 136.650 23.945 136.820 ;
        RECT 24.735 136.650 24.905 136.820 ;
        RECT 1.565 133.590 1.735 133.760 ;
        RECT 1.565 133.230 1.735 133.400 ;
        RECT 1.565 132.870 1.735 133.040 ;
        RECT 2.525 133.590 2.695 133.760 ;
        RECT 2.525 133.230 2.695 133.400 ;
        RECT 2.525 132.870 2.695 133.040 ;
        RECT 3.485 133.590 3.655 133.760 ;
        RECT 3.485 133.230 3.655 133.400 ;
        RECT 3.485 132.870 3.655 133.040 ;
        RECT 4.445 133.590 4.615 133.760 ;
        RECT 4.445 133.230 4.615 133.400 ;
        RECT 4.445 132.870 4.615 133.040 ;
        RECT 5.405 133.590 5.575 133.760 ;
        RECT 5.405 133.230 5.575 133.400 ;
        RECT 5.405 132.870 5.575 133.040 ;
        RECT 6.365 133.590 6.535 133.760 ;
        RECT 6.365 133.230 6.535 133.400 ;
        RECT 6.365 132.870 6.535 133.040 ;
        RECT 12.330 133.610 12.500 133.780 ;
        RECT 12.330 133.250 12.500 133.420 ;
        RECT 12.330 132.890 12.500 133.060 ;
        RECT 12.810 133.610 12.980 133.780 ;
        RECT 12.810 133.250 12.980 133.420 ;
        RECT 12.810 132.890 12.980 133.060 ;
        RECT 13.290 133.610 13.460 133.780 ;
        RECT 13.290 133.250 13.460 133.420 ;
        RECT 13.290 132.890 13.460 133.060 ;
        RECT 13.770 133.610 13.940 133.780 ;
        RECT 13.770 133.250 13.940 133.420 ;
        RECT 13.770 132.890 13.940 133.060 ;
        RECT 14.250 133.610 14.420 133.780 ;
        RECT 14.250 133.250 14.420 133.420 ;
        RECT 14.250 132.890 14.420 133.060 ;
        RECT 14.730 133.610 14.900 133.780 ;
        RECT 14.730 133.250 14.900 133.420 ;
        RECT 14.730 132.890 14.900 133.060 ;
        RECT 15.210 133.610 15.380 133.780 ;
        RECT 15.210 133.250 15.380 133.420 ;
        RECT 15.210 132.890 15.380 133.060 ;
        RECT 15.690 133.610 15.860 133.780 ;
        RECT 15.690 133.250 15.860 133.420 ;
        RECT 15.690 132.890 15.860 133.060 ;
        RECT 16.170 133.610 16.340 133.780 ;
        RECT 16.170 133.250 16.340 133.420 ;
        RECT 16.170 132.890 16.340 133.060 ;
        RECT 16.650 133.610 16.820 133.780 ;
        RECT 16.650 133.250 16.820 133.420 ;
        RECT 16.650 132.890 16.820 133.060 ;
        RECT 17.130 133.610 17.300 133.780 ;
        RECT 17.130 133.250 17.300 133.420 ;
        RECT 17.130 132.890 17.300 133.060 ;
        RECT 20.415 133.610 20.585 133.780 ;
        RECT 20.415 133.250 20.585 133.420 ;
        RECT 20.415 132.890 20.585 133.060 ;
        RECT 21.375 133.610 21.545 133.780 ;
        RECT 21.375 133.250 21.545 133.420 ;
        RECT 21.375 132.890 21.545 133.060 ;
        RECT 22.335 133.610 22.505 133.780 ;
        RECT 22.335 133.250 22.505 133.420 ;
        RECT 22.335 132.890 22.505 133.060 ;
        RECT 23.295 133.610 23.465 133.780 ;
        RECT 23.295 133.250 23.465 133.420 ;
        RECT 23.295 132.890 23.465 133.060 ;
        RECT 24.255 133.610 24.425 133.780 ;
        RECT 24.255 133.250 24.425 133.420 ;
        RECT 24.255 132.890 24.425 133.060 ;
        RECT 26.740 131.530 26.910 131.700 ;
        RECT 1.565 130.750 1.735 130.920 ;
        RECT 2.525 130.750 2.695 130.920 ;
        RECT 3.485 130.750 3.655 130.920 ;
        RECT 4.445 130.750 4.615 130.920 ;
        RECT 5.405 130.750 5.575 130.920 ;
        RECT 6.365 130.750 6.535 130.920 ;
        RECT 12.330 130.770 12.500 130.940 ;
        RECT 12.810 130.770 12.980 130.940 ;
        RECT 13.290 130.770 13.460 130.940 ;
        RECT 13.770 130.770 13.940 130.940 ;
        RECT 14.250 130.770 14.420 130.940 ;
        RECT 14.730 130.770 14.900 130.940 ;
        RECT 15.210 130.770 15.380 130.940 ;
        RECT 15.690 130.770 15.860 130.940 ;
        RECT 16.170 130.770 16.340 130.940 ;
        RECT 16.650 130.770 16.820 130.940 ;
        RECT 17.130 130.770 17.300 130.940 ;
        RECT 18.675 130.695 18.845 131.075 ;
        RECT 20.415 130.770 20.585 130.940 ;
        RECT 21.375 130.770 21.545 130.940 ;
        RECT 22.335 130.770 22.505 130.940 ;
        RECT 23.295 130.770 23.465 130.940 ;
        RECT 24.255 130.770 24.425 130.940 ;
        RECT 12.330 130.215 12.500 130.385 ;
        RECT 13.290 130.215 13.460 130.385 ;
        RECT 14.250 130.215 14.420 130.385 ;
        RECT 15.210 130.215 15.380 130.385 ;
        RECT 16.170 130.215 16.340 130.385 ;
        RECT 17.130 130.215 17.300 130.385 ;
        RECT 19.935 130.215 20.105 130.385 ;
        RECT 20.895 130.215 21.065 130.385 ;
        RECT 21.855 130.215 22.025 130.385 ;
        RECT 22.815 130.215 22.985 130.385 ;
        RECT 23.775 130.215 23.945 130.385 ;
        RECT 24.735 130.215 24.905 130.385 ;
        RECT 1.565 127.155 1.735 127.325 ;
        RECT 1.565 126.795 1.735 126.965 ;
        RECT 1.565 126.435 1.735 126.605 ;
        RECT 2.525 127.155 2.695 127.325 ;
        RECT 2.525 126.795 2.695 126.965 ;
        RECT 2.525 126.435 2.695 126.605 ;
        RECT 3.485 127.155 3.655 127.325 ;
        RECT 3.485 126.795 3.655 126.965 ;
        RECT 3.485 126.435 3.655 126.605 ;
        RECT 4.445 127.155 4.615 127.325 ;
        RECT 4.445 126.795 4.615 126.965 ;
        RECT 4.445 126.435 4.615 126.605 ;
        RECT 5.405 127.155 5.575 127.325 ;
        RECT 5.405 126.795 5.575 126.965 ;
        RECT 5.405 126.435 5.575 126.605 ;
        RECT 6.365 127.155 6.535 127.325 ;
        RECT 6.365 126.795 6.535 126.965 ;
        RECT 6.365 126.435 6.535 126.605 ;
        RECT 12.330 127.175 12.500 127.345 ;
        RECT 12.330 126.815 12.500 126.985 ;
        RECT 12.330 126.455 12.500 126.625 ;
        RECT 12.810 127.175 12.980 127.345 ;
        RECT 12.810 126.815 12.980 126.985 ;
        RECT 12.810 126.455 12.980 126.625 ;
        RECT 13.290 127.175 13.460 127.345 ;
        RECT 13.290 126.815 13.460 126.985 ;
        RECT 13.290 126.455 13.460 126.625 ;
        RECT 13.770 127.175 13.940 127.345 ;
        RECT 13.770 126.815 13.940 126.985 ;
        RECT 13.770 126.455 13.940 126.625 ;
        RECT 14.250 127.175 14.420 127.345 ;
        RECT 14.250 126.815 14.420 126.985 ;
        RECT 14.250 126.455 14.420 126.625 ;
        RECT 14.730 127.175 14.900 127.345 ;
        RECT 14.730 126.815 14.900 126.985 ;
        RECT 14.730 126.455 14.900 126.625 ;
        RECT 15.210 127.175 15.380 127.345 ;
        RECT 15.210 126.815 15.380 126.985 ;
        RECT 15.210 126.455 15.380 126.625 ;
        RECT 15.690 127.175 15.860 127.345 ;
        RECT 15.690 126.815 15.860 126.985 ;
        RECT 15.690 126.455 15.860 126.625 ;
        RECT 16.170 127.175 16.340 127.345 ;
        RECT 16.170 126.815 16.340 126.985 ;
        RECT 16.170 126.455 16.340 126.625 ;
        RECT 16.650 127.175 16.820 127.345 ;
        RECT 16.650 126.815 16.820 126.985 ;
        RECT 16.650 126.455 16.820 126.625 ;
        RECT 17.130 127.175 17.300 127.345 ;
        RECT 17.130 126.815 17.300 126.985 ;
        RECT 17.130 126.455 17.300 126.625 ;
        RECT 20.415 127.175 20.585 127.345 ;
        RECT 20.415 126.815 20.585 126.985 ;
        RECT 20.415 126.455 20.585 126.625 ;
        RECT 21.375 127.175 21.545 127.345 ;
        RECT 21.375 126.815 21.545 126.985 ;
        RECT 21.375 126.455 21.545 126.625 ;
        RECT 22.335 127.175 22.505 127.345 ;
        RECT 22.335 126.815 22.505 126.985 ;
        RECT 22.335 126.455 22.505 126.625 ;
        RECT 23.295 127.175 23.465 127.345 ;
        RECT 23.295 126.815 23.465 126.985 ;
        RECT 23.295 126.455 23.465 126.625 ;
        RECT 24.255 127.175 24.425 127.345 ;
        RECT 24.255 126.815 24.425 126.985 ;
        RECT 24.255 126.455 24.425 126.625 ;
        RECT 26.740 125.095 26.910 125.265 ;
        RECT 1.565 124.315 1.735 124.485 ;
        RECT 2.525 124.315 2.695 124.485 ;
        RECT 3.485 124.315 3.655 124.485 ;
        RECT 4.445 124.315 4.615 124.485 ;
        RECT 5.405 124.315 5.575 124.485 ;
        RECT 6.365 124.315 6.535 124.485 ;
        RECT 12.330 124.335 12.500 124.505 ;
        RECT 12.810 124.335 12.980 124.505 ;
        RECT 13.290 124.335 13.460 124.505 ;
        RECT 13.770 124.335 13.940 124.505 ;
        RECT 14.250 124.335 14.420 124.505 ;
        RECT 14.730 124.335 14.900 124.505 ;
        RECT 15.210 124.335 15.380 124.505 ;
        RECT 15.690 124.335 15.860 124.505 ;
        RECT 16.170 124.335 16.340 124.505 ;
        RECT 16.650 124.335 16.820 124.505 ;
        RECT 17.130 124.335 17.300 124.505 ;
        RECT 18.675 124.260 18.845 124.640 ;
        RECT 20.415 124.335 20.585 124.505 ;
        RECT 21.375 124.335 21.545 124.505 ;
        RECT 22.335 124.335 22.505 124.505 ;
        RECT 23.295 124.335 23.465 124.505 ;
        RECT 24.255 124.335 24.425 124.505 ;
        RECT 12.330 123.780 12.500 123.950 ;
        RECT 13.290 123.780 13.460 123.950 ;
        RECT 14.250 123.780 14.420 123.950 ;
        RECT 15.210 123.780 15.380 123.950 ;
        RECT 16.170 123.780 16.340 123.950 ;
        RECT 17.130 123.780 17.300 123.950 ;
        RECT 19.935 123.780 20.105 123.950 ;
        RECT 20.895 123.780 21.065 123.950 ;
        RECT 21.855 123.780 22.025 123.950 ;
        RECT 22.815 123.780 22.985 123.950 ;
        RECT 23.775 123.780 23.945 123.950 ;
        RECT 24.735 123.780 24.905 123.950 ;
        RECT 1.565 120.720 1.735 120.890 ;
        RECT 1.565 120.360 1.735 120.530 ;
        RECT 1.565 120.000 1.735 120.170 ;
        RECT 2.525 120.720 2.695 120.890 ;
        RECT 2.525 120.360 2.695 120.530 ;
        RECT 2.525 120.000 2.695 120.170 ;
        RECT 3.485 120.720 3.655 120.890 ;
        RECT 3.485 120.360 3.655 120.530 ;
        RECT 3.485 120.000 3.655 120.170 ;
        RECT 4.445 120.720 4.615 120.890 ;
        RECT 4.445 120.360 4.615 120.530 ;
        RECT 4.445 120.000 4.615 120.170 ;
        RECT 5.405 120.720 5.575 120.890 ;
        RECT 5.405 120.360 5.575 120.530 ;
        RECT 5.405 120.000 5.575 120.170 ;
        RECT 6.365 120.720 6.535 120.890 ;
        RECT 6.365 120.360 6.535 120.530 ;
        RECT 6.365 120.000 6.535 120.170 ;
        RECT 12.330 120.740 12.500 120.910 ;
        RECT 12.330 120.380 12.500 120.550 ;
        RECT 12.330 120.020 12.500 120.190 ;
        RECT 12.810 120.740 12.980 120.910 ;
        RECT 12.810 120.380 12.980 120.550 ;
        RECT 12.810 120.020 12.980 120.190 ;
        RECT 13.290 120.740 13.460 120.910 ;
        RECT 13.290 120.380 13.460 120.550 ;
        RECT 13.290 120.020 13.460 120.190 ;
        RECT 13.770 120.740 13.940 120.910 ;
        RECT 13.770 120.380 13.940 120.550 ;
        RECT 13.770 120.020 13.940 120.190 ;
        RECT 14.250 120.740 14.420 120.910 ;
        RECT 14.250 120.380 14.420 120.550 ;
        RECT 14.250 120.020 14.420 120.190 ;
        RECT 14.730 120.740 14.900 120.910 ;
        RECT 14.730 120.380 14.900 120.550 ;
        RECT 14.730 120.020 14.900 120.190 ;
        RECT 15.210 120.740 15.380 120.910 ;
        RECT 15.210 120.380 15.380 120.550 ;
        RECT 15.210 120.020 15.380 120.190 ;
        RECT 15.690 120.740 15.860 120.910 ;
        RECT 15.690 120.380 15.860 120.550 ;
        RECT 15.690 120.020 15.860 120.190 ;
        RECT 16.170 120.740 16.340 120.910 ;
        RECT 16.170 120.380 16.340 120.550 ;
        RECT 16.170 120.020 16.340 120.190 ;
        RECT 16.650 120.740 16.820 120.910 ;
        RECT 16.650 120.380 16.820 120.550 ;
        RECT 16.650 120.020 16.820 120.190 ;
        RECT 17.130 120.740 17.300 120.910 ;
        RECT 17.130 120.380 17.300 120.550 ;
        RECT 17.130 120.020 17.300 120.190 ;
        RECT 20.415 120.740 20.585 120.910 ;
        RECT 20.415 120.380 20.585 120.550 ;
        RECT 20.415 120.020 20.585 120.190 ;
        RECT 21.375 120.740 21.545 120.910 ;
        RECT 21.375 120.380 21.545 120.550 ;
        RECT 21.375 120.020 21.545 120.190 ;
        RECT 22.335 120.740 22.505 120.910 ;
        RECT 22.335 120.380 22.505 120.550 ;
        RECT 22.335 120.020 22.505 120.190 ;
        RECT 23.295 120.740 23.465 120.910 ;
        RECT 23.295 120.380 23.465 120.550 ;
        RECT 23.295 120.020 23.465 120.190 ;
        RECT 24.255 120.740 24.425 120.910 ;
        RECT 24.255 120.380 24.425 120.550 ;
        RECT 24.255 120.020 24.425 120.190 ;
        RECT 26.740 118.660 26.910 118.830 ;
        RECT 1.565 117.880 1.735 118.050 ;
        RECT 2.525 117.880 2.695 118.050 ;
        RECT 3.485 117.880 3.655 118.050 ;
        RECT 4.445 117.880 4.615 118.050 ;
        RECT 5.405 117.880 5.575 118.050 ;
        RECT 6.365 117.880 6.535 118.050 ;
        RECT 12.330 117.900 12.500 118.070 ;
        RECT 12.810 117.900 12.980 118.070 ;
        RECT 13.290 117.900 13.460 118.070 ;
        RECT 13.770 117.900 13.940 118.070 ;
        RECT 14.250 117.900 14.420 118.070 ;
        RECT 14.730 117.900 14.900 118.070 ;
        RECT 15.210 117.900 15.380 118.070 ;
        RECT 15.690 117.900 15.860 118.070 ;
        RECT 16.170 117.900 16.340 118.070 ;
        RECT 16.650 117.900 16.820 118.070 ;
        RECT 17.130 117.900 17.300 118.070 ;
        RECT 18.675 117.825 18.845 118.205 ;
        RECT 20.415 117.900 20.585 118.070 ;
        RECT 21.375 117.900 21.545 118.070 ;
        RECT 22.335 117.900 22.505 118.070 ;
        RECT 23.295 117.900 23.465 118.070 ;
        RECT 24.255 117.900 24.425 118.070 ;
        RECT 12.330 117.345 12.500 117.515 ;
        RECT 13.290 117.345 13.460 117.515 ;
        RECT 14.250 117.345 14.420 117.515 ;
        RECT 15.210 117.345 15.380 117.515 ;
        RECT 16.170 117.345 16.340 117.515 ;
        RECT 17.130 117.345 17.300 117.515 ;
        RECT 19.935 117.345 20.105 117.515 ;
        RECT 20.895 117.345 21.065 117.515 ;
        RECT 21.855 117.345 22.025 117.515 ;
        RECT 22.815 117.345 22.985 117.515 ;
        RECT 23.775 117.345 23.945 117.515 ;
        RECT 24.735 117.345 24.905 117.515 ;
        RECT 1.565 114.285 1.735 114.455 ;
        RECT 1.565 113.925 1.735 114.095 ;
        RECT 1.565 113.565 1.735 113.735 ;
        RECT 2.525 114.285 2.695 114.455 ;
        RECT 2.525 113.925 2.695 114.095 ;
        RECT 2.525 113.565 2.695 113.735 ;
        RECT 3.485 114.285 3.655 114.455 ;
        RECT 3.485 113.925 3.655 114.095 ;
        RECT 3.485 113.565 3.655 113.735 ;
        RECT 4.445 114.285 4.615 114.455 ;
        RECT 4.445 113.925 4.615 114.095 ;
        RECT 4.445 113.565 4.615 113.735 ;
        RECT 5.405 114.285 5.575 114.455 ;
        RECT 5.405 113.925 5.575 114.095 ;
        RECT 5.405 113.565 5.575 113.735 ;
        RECT 6.365 114.285 6.535 114.455 ;
        RECT 6.365 113.925 6.535 114.095 ;
        RECT 6.365 113.565 6.535 113.735 ;
        RECT 12.330 114.305 12.500 114.475 ;
        RECT 12.330 113.945 12.500 114.115 ;
        RECT 12.330 113.585 12.500 113.755 ;
        RECT 12.810 114.305 12.980 114.475 ;
        RECT 12.810 113.945 12.980 114.115 ;
        RECT 12.810 113.585 12.980 113.755 ;
        RECT 13.290 114.305 13.460 114.475 ;
        RECT 13.290 113.945 13.460 114.115 ;
        RECT 13.290 113.585 13.460 113.755 ;
        RECT 13.770 114.305 13.940 114.475 ;
        RECT 13.770 113.945 13.940 114.115 ;
        RECT 13.770 113.585 13.940 113.755 ;
        RECT 14.250 114.305 14.420 114.475 ;
        RECT 14.250 113.945 14.420 114.115 ;
        RECT 14.250 113.585 14.420 113.755 ;
        RECT 14.730 114.305 14.900 114.475 ;
        RECT 14.730 113.945 14.900 114.115 ;
        RECT 14.730 113.585 14.900 113.755 ;
        RECT 15.210 114.305 15.380 114.475 ;
        RECT 15.210 113.945 15.380 114.115 ;
        RECT 15.210 113.585 15.380 113.755 ;
        RECT 15.690 114.305 15.860 114.475 ;
        RECT 15.690 113.945 15.860 114.115 ;
        RECT 15.690 113.585 15.860 113.755 ;
        RECT 16.170 114.305 16.340 114.475 ;
        RECT 16.170 113.945 16.340 114.115 ;
        RECT 16.170 113.585 16.340 113.755 ;
        RECT 16.650 114.305 16.820 114.475 ;
        RECT 16.650 113.945 16.820 114.115 ;
        RECT 16.650 113.585 16.820 113.755 ;
        RECT 17.130 114.305 17.300 114.475 ;
        RECT 17.130 113.945 17.300 114.115 ;
        RECT 17.130 113.585 17.300 113.755 ;
        RECT 20.415 114.305 20.585 114.475 ;
        RECT 20.415 113.945 20.585 114.115 ;
        RECT 20.415 113.585 20.585 113.755 ;
        RECT 21.375 114.305 21.545 114.475 ;
        RECT 21.375 113.945 21.545 114.115 ;
        RECT 21.375 113.585 21.545 113.755 ;
        RECT 22.335 114.305 22.505 114.475 ;
        RECT 22.335 113.945 22.505 114.115 ;
        RECT 22.335 113.585 22.505 113.755 ;
        RECT 23.295 114.305 23.465 114.475 ;
        RECT 23.295 113.945 23.465 114.115 ;
        RECT 23.295 113.585 23.465 113.755 ;
        RECT 24.255 114.305 24.425 114.475 ;
        RECT 24.255 113.945 24.425 114.115 ;
        RECT 24.255 113.585 24.425 113.755 ;
        RECT 26.740 112.225 26.910 112.395 ;
        RECT 1.565 111.445 1.735 111.615 ;
        RECT 2.525 111.445 2.695 111.615 ;
        RECT 3.485 111.445 3.655 111.615 ;
        RECT 4.445 111.445 4.615 111.615 ;
        RECT 5.405 111.445 5.575 111.615 ;
        RECT 6.365 111.445 6.535 111.615 ;
        RECT 12.330 111.465 12.500 111.635 ;
        RECT 12.810 111.465 12.980 111.635 ;
        RECT 13.290 111.465 13.460 111.635 ;
        RECT 13.770 111.465 13.940 111.635 ;
        RECT 14.250 111.465 14.420 111.635 ;
        RECT 14.730 111.465 14.900 111.635 ;
        RECT 15.210 111.465 15.380 111.635 ;
        RECT 15.690 111.465 15.860 111.635 ;
        RECT 16.170 111.465 16.340 111.635 ;
        RECT 16.650 111.465 16.820 111.635 ;
        RECT 17.130 111.465 17.300 111.635 ;
        RECT 18.675 111.390 18.845 111.770 ;
        RECT 20.415 111.465 20.585 111.635 ;
        RECT 21.375 111.465 21.545 111.635 ;
        RECT 22.335 111.465 22.505 111.635 ;
        RECT 23.295 111.465 23.465 111.635 ;
        RECT 24.255 111.465 24.425 111.635 ;
        RECT 12.330 110.910 12.500 111.080 ;
        RECT 13.290 110.910 13.460 111.080 ;
        RECT 14.250 110.910 14.420 111.080 ;
        RECT 15.210 110.910 15.380 111.080 ;
        RECT 16.170 110.910 16.340 111.080 ;
        RECT 17.130 110.910 17.300 111.080 ;
        RECT 19.935 110.910 20.105 111.080 ;
        RECT 20.895 110.910 21.065 111.080 ;
        RECT 21.855 110.910 22.025 111.080 ;
        RECT 22.815 110.910 22.985 111.080 ;
        RECT 23.775 110.910 23.945 111.080 ;
        RECT 24.735 110.910 24.905 111.080 ;
        RECT 1.565 107.850 1.735 108.020 ;
        RECT 1.565 107.490 1.735 107.660 ;
        RECT 1.565 107.130 1.735 107.300 ;
        RECT 2.525 107.850 2.695 108.020 ;
        RECT 2.525 107.490 2.695 107.660 ;
        RECT 2.525 107.130 2.695 107.300 ;
        RECT 3.485 107.850 3.655 108.020 ;
        RECT 3.485 107.490 3.655 107.660 ;
        RECT 3.485 107.130 3.655 107.300 ;
        RECT 4.445 107.850 4.615 108.020 ;
        RECT 4.445 107.490 4.615 107.660 ;
        RECT 4.445 107.130 4.615 107.300 ;
        RECT 5.405 107.850 5.575 108.020 ;
        RECT 5.405 107.490 5.575 107.660 ;
        RECT 5.405 107.130 5.575 107.300 ;
        RECT 6.365 107.850 6.535 108.020 ;
        RECT 6.365 107.490 6.535 107.660 ;
        RECT 6.365 107.130 6.535 107.300 ;
        RECT 12.330 107.870 12.500 108.040 ;
        RECT 12.330 107.510 12.500 107.680 ;
        RECT 12.330 107.150 12.500 107.320 ;
        RECT 12.810 107.870 12.980 108.040 ;
        RECT 12.810 107.510 12.980 107.680 ;
        RECT 12.810 107.150 12.980 107.320 ;
        RECT 13.290 107.870 13.460 108.040 ;
        RECT 13.290 107.510 13.460 107.680 ;
        RECT 13.290 107.150 13.460 107.320 ;
        RECT 13.770 107.870 13.940 108.040 ;
        RECT 13.770 107.510 13.940 107.680 ;
        RECT 13.770 107.150 13.940 107.320 ;
        RECT 14.250 107.870 14.420 108.040 ;
        RECT 14.250 107.510 14.420 107.680 ;
        RECT 14.250 107.150 14.420 107.320 ;
        RECT 14.730 107.870 14.900 108.040 ;
        RECT 14.730 107.510 14.900 107.680 ;
        RECT 14.730 107.150 14.900 107.320 ;
        RECT 15.210 107.870 15.380 108.040 ;
        RECT 15.210 107.510 15.380 107.680 ;
        RECT 15.210 107.150 15.380 107.320 ;
        RECT 15.690 107.870 15.860 108.040 ;
        RECT 15.690 107.510 15.860 107.680 ;
        RECT 15.690 107.150 15.860 107.320 ;
        RECT 16.170 107.870 16.340 108.040 ;
        RECT 16.170 107.510 16.340 107.680 ;
        RECT 16.170 107.150 16.340 107.320 ;
        RECT 16.650 107.870 16.820 108.040 ;
        RECT 16.650 107.510 16.820 107.680 ;
        RECT 16.650 107.150 16.820 107.320 ;
        RECT 17.130 107.870 17.300 108.040 ;
        RECT 17.130 107.510 17.300 107.680 ;
        RECT 17.130 107.150 17.300 107.320 ;
        RECT 20.415 107.870 20.585 108.040 ;
        RECT 20.415 107.510 20.585 107.680 ;
        RECT 20.415 107.150 20.585 107.320 ;
        RECT 21.375 107.870 21.545 108.040 ;
        RECT 21.375 107.510 21.545 107.680 ;
        RECT 21.375 107.150 21.545 107.320 ;
        RECT 22.335 107.870 22.505 108.040 ;
        RECT 22.335 107.510 22.505 107.680 ;
        RECT 22.335 107.150 22.505 107.320 ;
        RECT 23.295 107.870 23.465 108.040 ;
        RECT 23.295 107.510 23.465 107.680 ;
        RECT 23.295 107.150 23.465 107.320 ;
        RECT 24.255 107.870 24.425 108.040 ;
        RECT 24.255 107.510 24.425 107.680 ;
        RECT 24.255 107.150 24.425 107.320 ;
        RECT 26.740 105.790 26.910 105.960 ;
        RECT 1.565 105.010 1.735 105.180 ;
        RECT 2.525 105.010 2.695 105.180 ;
        RECT 3.485 105.010 3.655 105.180 ;
        RECT 4.445 105.010 4.615 105.180 ;
        RECT 5.405 105.010 5.575 105.180 ;
        RECT 6.365 105.010 6.535 105.180 ;
        RECT 12.330 105.030 12.500 105.200 ;
        RECT 12.810 105.030 12.980 105.200 ;
        RECT 13.290 105.030 13.460 105.200 ;
        RECT 13.770 105.030 13.940 105.200 ;
        RECT 14.250 105.030 14.420 105.200 ;
        RECT 14.730 105.030 14.900 105.200 ;
        RECT 15.210 105.030 15.380 105.200 ;
        RECT 15.690 105.030 15.860 105.200 ;
        RECT 16.170 105.030 16.340 105.200 ;
        RECT 16.650 105.030 16.820 105.200 ;
        RECT 17.130 105.030 17.300 105.200 ;
        RECT 18.675 104.955 18.845 105.335 ;
        RECT 20.415 105.030 20.585 105.200 ;
        RECT 21.375 105.030 21.545 105.200 ;
        RECT 22.335 105.030 22.505 105.200 ;
        RECT 23.295 105.030 23.465 105.200 ;
        RECT 24.255 105.030 24.425 105.200 ;
        RECT 12.330 104.475 12.500 104.645 ;
        RECT 13.290 104.475 13.460 104.645 ;
        RECT 14.250 104.475 14.420 104.645 ;
        RECT 15.210 104.475 15.380 104.645 ;
        RECT 16.170 104.475 16.340 104.645 ;
        RECT 17.130 104.475 17.300 104.645 ;
        RECT 19.935 104.475 20.105 104.645 ;
        RECT 20.895 104.475 21.065 104.645 ;
        RECT 21.855 104.475 22.025 104.645 ;
        RECT 22.815 104.475 22.985 104.645 ;
        RECT 23.775 104.475 23.945 104.645 ;
        RECT 24.735 104.475 24.905 104.645 ;
        RECT 1.565 101.415 1.735 101.585 ;
        RECT 1.565 101.055 1.735 101.225 ;
        RECT 1.565 100.695 1.735 100.865 ;
        RECT 2.525 101.415 2.695 101.585 ;
        RECT 2.525 101.055 2.695 101.225 ;
        RECT 2.525 100.695 2.695 100.865 ;
        RECT 3.485 101.415 3.655 101.585 ;
        RECT 3.485 101.055 3.655 101.225 ;
        RECT 3.485 100.695 3.655 100.865 ;
        RECT 4.445 101.415 4.615 101.585 ;
        RECT 4.445 101.055 4.615 101.225 ;
        RECT 4.445 100.695 4.615 100.865 ;
        RECT 5.405 101.415 5.575 101.585 ;
        RECT 5.405 101.055 5.575 101.225 ;
        RECT 5.405 100.695 5.575 100.865 ;
        RECT 6.365 101.415 6.535 101.585 ;
        RECT 6.365 101.055 6.535 101.225 ;
        RECT 6.365 100.695 6.535 100.865 ;
        RECT 12.330 101.435 12.500 101.605 ;
        RECT 12.330 101.075 12.500 101.245 ;
        RECT 12.330 100.715 12.500 100.885 ;
        RECT 12.810 101.435 12.980 101.605 ;
        RECT 12.810 101.075 12.980 101.245 ;
        RECT 12.810 100.715 12.980 100.885 ;
        RECT 13.290 101.435 13.460 101.605 ;
        RECT 13.290 101.075 13.460 101.245 ;
        RECT 13.290 100.715 13.460 100.885 ;
        RECT 13.770 101.435 13.940 101.605 ;
        RECT 13.770 101.075 13.940 101.245 ;
        RECT 13.770 100.715 13.940 100.885 ;
        RECT 14.250 101.435 14.420 101.605 ;
        RECT 14.250 101.075 14.420 101.245 ;
        RECT 14.250 100.715 14.420 100.885 ;
        RECT 14.730 101.435 14.900 101.605 ;
        RECT 14.730 101.075 14.900 101.245 ;
        RECT 14.730 100.715 14.900 100.885 ;
        RECT 15.210 101.435 15.380 101.605 ;
        RECT 15.210 101.075 15.380 101.245 ;
        RECT 15.210 100.715 15.380 100.885 ;
        RECT 15.690 101.435 15.860 101.605 ;
        RECT 15.690 101.075 15.860 101.245 ;
        RECT 15.690 100.715 15.860 100.885 ;
        RECT 16.170 101.435 16.340 101.605 ;
        RECT 16.170 101.075 16.340 101.245 ;
        RECT 16.170 100.715 16.340 100.885 ;
        RECT 16.650 101.435 16.820 101.605 ;
        RECT 16.650 101.075 16.820 101.245 ;
        RECT 16.650 100.715 16.820 100.885 ;
        RECT 17.130 101.435 17.300 101.605 ;
        RECT 17.130 101.075 17.300 101.245 ;
        RECT 17.130 100.715 17.300 100.885 ;
        RECT 20.415 101.435 20.585 101.605 ;
        RECT 20.415 101.075 20.585 101.245 ;
        RECT 20.415 100.715 20.585 100.885 ;
        RECT 21.375 101.435 21.545 101.605 ;
        RECT 21.375 101.075 21.545 101.245 ;
        RECT 21.375 100.715 21.545 100.885 ;
        RECT 22.335 101.435 22.505 101.605 ;
        RECT 22.335 101.075 22.505 101.245 ;
        RECT 22.335 100.715 22.505 100.885 ;
        RECT 23.295 101.435 23.465 101.605 ;
        RECT 23.295 101.075 23.465 101.245 ;
        RECT 23.295 100.715 23.465 100.885 ;
        RECT 24.255 101.435 24.425 101.605 ;
        RECT 24.255 101.075 24.425 101.245 ;
        RECT 24.255 100.715 24.425 100.885 ;
        RECT 26.740 99.355 26.910 99.525 ;
        RECT 1.565 98.575 1.735 98.745 ;
        RECT 2.525 98.575 2.695 98.745 ;
        RECT 3.485 98.575 3.655 98.745 ;
        RECT 4.445 98.575 4.615 98.745 ;
        RECT 5.405 98.575 5.575 98.745 ;
        RECT 6.365 98.575 6.535 98.745 ;
        RECT 12.330 98.595 12.500 98.765 ;
        RECT 12.810 98.595 12.980 98.765 ;
        RECT 13.290 98.595 13.460 98.765 ;
        RECT 13.770 98.595 13.940 98.765 ;
        RECT 14.250 98.595 14.420 98.765 ;
        RECT 14.730 98.595 14.900 98.765 ;
        RECT 15.210 98.595 15.380 98.765 ;
        RECT 15.690 98.595 15.860 98.765 ;
        RECT 16.170 98.595 16.340 98.765 ;
        RECT 16.650 98.595 16.820 98.765 ;
        RECT 17.130 98.595 17.300 98.765 ;
        RECT 18.675 98.520 18.845 98.900 ;
        RECT 20.415 98.595 20.585 98.765 ;
        RECT 21.375 98.595 21.545 98.765 ;
        RECT 22.335 98.595 22.505 98.765 ;
        RECT 23.295 98.595 23.465 98.765 ;
        RECT 24.255 98.595 24.425 98.765 ;
        RECT 12.330 98.040 12.500 98.210 ;
        RECT 13.290 98.040 13.460 98.210 ;
        RECT 14.250 98.040 14.420 98.210 ;
        RECT 15.210 98.040 15.380 98.210 ;
        RECT 16.170 98.040 16.340 98.210 ;
        RECT 17.130 98.040 17.300 98.210 ;
        RECT 19.935 98.040 20.105 98.210 ;
        RECT 20.895 98.040 21.065 98.210 ;
        RECT 21.855 98.040 22.025 98.210 ;
        RECT 22.815 98.040 22.985 98.210 ;
        RECT 23.775 98.040 23.945 98.210 ;
        RECT 24.735 98.040 24.905 98.210 ;
        RECT 1.565 94.980 1.735 95.150 ;
        RECT 1.565 94.620 1.735 94.790 ;
        RECT 1.565 94.260 1.735 94.430 ;
        RECT 2.525 94.980 2.695 95.150 ;
        RECT 2.525 94.620 2.695 94.790 ;
        RECT 2.525 94.260 2.695 94.430 ;
        RECT 3.485 94.980 3.655 95.150 ;
        RECT 3.485 94.620 3.655 94.790 ;
        RECT 3.485 94.260 3.655 94.430 ;
        RECT 4.445 94.980 4.615 95.150 ;
        RECT 4.445 94.620 4.615 94.790 ;
        RECT 4.445 94.260 4.615 94.430 ;
        RECT 5.405 94.980 5.575 95.150 ;
        RECT 5.405 94.620 5.575 94.790 ;
        RECT 5.405 94.260 5.575 94.430 ;
        RECT 6.365 94.980 6.535 95.150 ;
        RECT 6.365 94.620 6.535 94.790 ;
        RECT 6.365 94.260 6.535 94.430 ;
        RECT 12.330 95.000 12.500 95.170 ;
        RECT 12.330 94.640 12.500 94.810 ;
        RECT 12.330 94.280 12.500 94.450 ;
        RECT 12.810 95.000 12.980 95.170 ;
        RECT 12.810 94.640 12.980 94.810 ;
        RECT 12.810 94.280 12.980 94.450 ;
        RECT 13.290 95.000 13.460 95.170 ;
        RECT 13.290 94.640 13.460 94.810 ;
        RECT 13.290 94.280 13.460 94.450 ;
        RECT 13.770 95.000 13.940 95.170 ;
        RECT 13.770 94.640 13.940 94.810 ;
        RECT 13.770 94.280 13.940 94.450 ;
        RECT 14.250 95.000 14.420 95.170 ;
        RECT 14.250 94.640 14.420 94.810 ;
        RECT 14.250 94.280 14.420 94.450 ;
        RECT 14.730 95.000 14.900 95.170 ;
        RECT 14.730 94.640 14.900 94.810 ;
        RECT 14.730 94.280 14.900 94.450 ;
        RECT 15.210 95.000 15.380 95.170 ;
        RECT 15.210 94.640 15.380 94.810 ;
        RECT 15.210 94.280 15.380 94.450 ;
        RECT 15.690 95.000 15.860 95.170 ;
        RECT 15.690 94.640 15.860 94.810 ;
        RECT 15.690 94.280 15.860 94.450 ;
        RECT 16.170 95.000 16.340 95.170 ;
        RECT 16.170 94.640 16.340 94.810 ;
        RECT 16.170 94.280 16.340 94.450 ;
        RECT 16.650 95.000 16.820 95.170 ;
        RECT 16.650 94.640 16.820 94.810 ;
        RECT 16.650 94.280 16.820 94.450 ;
        RECT 17.130 95.000 17.300 95.170 ;
        RECT 17.130 94.640 17.300 94.810 ;
        RECT 17.130 94.280 17.300 94.450 ;
        RECT 20.415 95.000 20.585 95.170 ;
        RECT 20.415 94.640 20.585 94.810 ;
        RECT 20.415 94.280 20.585 94.450 ;
        RECT 21.375 95.000 21.545 95.170 ;
        RECT 21.375 94.640 21.545 94.810 ;
        RECT 21.375 94.280 21.545 94.450 ;
        RECT 22.335 95.000 22.505 95.170 ;
        RECT 22.335 94.640 22.505 94.810 ;
        RECT 22.335 94.280 22.505 94.450 ;
        RECT 23.295 95.000 23.465 95.170 ;
        RECT 23.295 94.640 23.465 94.810 ;
        RECT 23.295 94.280 23.465 94.450 ;
        RECT 24.255 95.000 24.425 95.170 ;
        RECT 24.255 94.640 24.425 94.810 ;
        RECT 24.255 94.280 24.425 94.450 ;
        RECT 26.740 92.920 26.910 93.090 ;
        RECT 1.565 92.140 1.735 92.310 ;
        RECT 2.525 92.140 2.695 92.310 ;
        RECT 3.485 92.140 3.655 92.310 ;
        RECT 4.445 92.140 4.615 92.310 ;
        RECT 5.405 92.140 5.575 92.310 ;
        RECT 6.365 92.140 6.535 92.310 ;
        RECT 12.330 92.160 12.500 92.330 ;
        RECT 12.810 92.160 12.980 92.330 ;
        RECT 13.290 92.160 13.460 92.330 ;
        RECT 13.770 92.160 13.940 92.330 ;
        RECT 14.250 92.160 14.420 92.330 ;
        RECT 14.730 92.160 14.900 92.330 ;
        RECT 15.210 92.160 15.380 92.330 ;
        RECT 15.690 92.160 15.860 92.330 ;
        RECT 16.170 92.160 16.340 92.330 ;
        RECT 16.650 92.160 16.820 92.330 ;
        RECT 17.130 92.160 17.300 92.330 ;
        RECT 18.675 92.085 18.845 92.465 ;
        RECT 20.415 92.160 20.585 92.330 ;
        RECT 21.375 92.160 21.545 92.330 ;
        RECT 22.335 92.160 22.505 92.330 ;
        RECT 23.295 92.160 23.465 92.330 ;
        RECT 24.255 92.160 24.425 92.330 ;
        RECT 12.330 91.605 12.500 91.775 ;
        RECT 13.290 91.605 13.460 91.775 ;
        RECT 14.250 91.605 14.420 91.775 ;
        RECT 15.210 91.605 15.380 91.775 ;
        RECT 16.170 91.605 16.340 91.775 ;
        RECT 17.130 91.605 17.300 91.775 ;
        RECT 19.935 91.605 20.105 91.775 ;
        RECT 20.895 91.605 21.065 91.775 ;
        RECT 21.855 91.605 22.025 91.775 ;
        RECT 22.815 91.605 22.985 91.775 ;
        RECT 23.775 91.605 23.945 91.775 ;
        RECT 24.735 91.605 24.905 91.775 ;
        RECT 1.565 88.545 1.735 88.715 ;
        RECT 1.565 88.185 1.735 88.355 ;
        RECT 1.565 87.825 1.735 87.995 ;
        RECT 2.525 88.545 2.695 88.715 ;
        RECT 2.525 88.185 2.695 88.355 ;
        RECT 2.525 87.825 2.695 87.995 ;
        RECT 3.485 88.545 3.655 88.715 ;
        RECT 3.485 88.185 3.655 88.355 ;
        RECT 3.485 87.825 3.655 87.995 ;
        RECT 4.445 88.545 4.615 88.715 ;
        RECT 4.445 88.185 4.615 88.355 ;
        RECT 4.445 87.825 4.615 87.995 ;
        RECT 5.405 88.545 5.575 88.715 ;
        RECT 5.405 88.185 5.575 88.355 ;
        RECT 5.405 87.825 5.575 87.995 ;
        RECT 6.365 88.545 6.535 88.715 ;
        RECT 6.365 88.185 6.535 88.355 ;
        RECT 6.365 87.825 6.535 87.995 ;
        RECT 12.330 88.565 12.500 88.735 ;
        RECT 12.330 88.205 12.500 88.375 ;
        RECT 12.330 87.845 12.500 88.015 ;
        RECT 12.810 88.565 12.980 88.735 ;
        RECT 12.810 88.205 12.980 88.375 ;
        RECT 12.810 87.845 12.980 88.015 ;
        RECT 13.290 88.565 13.460 88.735 ;
        RECT 13.290 88.205 13.460 88.375 ;
        RECT 13.290 87.845 13.460 88.015 ;
        RECT 13.770 88.565 13.940 88.735 ;
        RECT 13.770 88.205 13.940 88.375 ;
        RECT 13.770 87.845 13.940 88.015 ;
        RECT 14.250 88.565 14.420 88.735 ;
        RECT 14.250 88.205 14.420 88.375 ;
        RECT 14.250 87.845 14.420 88.015 ;
        RECT 14.730 88.565 14.900 88.735 ;
        RECT 14.730 88.205 14.900 88.375 ;
        RECT 14.730 87.845 14.900 88.015 ;
        RECT 15.210 88.565 15.380 88.735 ;
        RECT 15.210 88.205 15.380 88.375 ;
        RECT 15.210 87.845 15.380 88.015 ;
        RECT 15.690 88.565 15.860 88.735 ;
        RECT 15.690 88.205 15.860 88.375 ;
        RECT 15.690 87.845 15.860 88.015 ;
        RECT 16.170 88.565 16.340 88.735 ;
        RECT 16.170 88.205 16.340 88.375 ;
        RECT 16.170 87.845 16.340 88.015 ;
        RECT 16.650 88.565 16.820 88.735 ;
        RECT 16.650 88.205 16.820 88.375 ;
        RECT 16.650 87.845 16.820 88.015 ;
        RECT 17.130 88.565 17.300 88.735 ;
        RECT 17.130 88.205 17.300 88.375 ;
        RECT 17.130 87.845 17.300 88.015 ;
        RECT 20.415 88.565 20.585 88.735 ;
        RECT 20.415 88.205 20.585 88.375 ;
        RECT 20.415 87.845 20.585 88.015 ;
        RECT 21.375 88.565 21.545 88.735 ;
        RECT 21.375 88.205 21.545 88.375 ;
        RECT 21.375 87.845 21.545 88.015 ;
        RECT 22.335 88.565 22.505 88.735 ;
        RECT 22.335 88.205 22.505 88.375 ;
        RECT 22.335 87.845 22.505 88.015 ;
        RECT 23.295 88.565 23.465 88.735 ;
        RECT 23.295 88.205 23.465 88.375 ;
        RECT 23.295 87.845 23.465 88.015 ;
        RECT 24.255 88.565 24.425 88.735 ;
        RECT 24.255 88.205 24.425 88.375 ;
        RECT 24.255 87.845 24.425 88.015 ;
        RECT 26.740 86.485 26.910 86.655 ;
        RECT 1.565 85.705 1.735 85.875 ;
        RECT 2.525 85.705 2.695 85.875 ;
        RECT 3.485 85.705 3.655 85.875 ;
        RECT 4.445 85.705 4.615 85.875 ;
        RECT 5.405 85.705 5.575 85.875 ;
        RECT 6.365 85.705 6.535 85.875 ;
        RECT 12.330 85.725 12.500 85.895 ;
        RECT 12.810 85.725 12.980 85.895 ;
        RECT 13.290 85.725 13.460 85.895 ;
        RECT 13.770 85.725 13.940 85.895 ;
        RECT 14.250 85.725 14.420 85.895 ;
        RECT 14.730 85.725 14.900 85.895 ;
        RECT 15.210 85.725 15.380 85.895 ;
        RECT 15.690 85.725 15.860 85.895 ;
        RECT 16.170 85.725 16.340 85.895 ;
        RECT 16.650 85.725 16.820 85.895 ;
        RECT 17.130 85.725 17.300 85.895 ;
        RECT 18.675 85.650 18.845 86.030 ;
        RECT 20.415 85.725 20.585 85.895 ;
        RECT 21.375 85.725 21.545 85.895 ;
        RECT 22.335 85.725 22.505 85.895 ;
        RECT 23.295 85.725 23.465 85.895 ;
        RECT 24.255 85.725 24.425 85.895 ;
        RECT 12.330 85.170 12.500 85.340 ;
        RECT 13.290 85.170 13.460 85.340 ;
        RECT 14.250 85.170 14.420 85.340 ;
        RECT 15.210 85.170 15.380 85.340 ;
        RECT 16.170 85.170 16.340 85.340 ;
        RECT 17.130 85.170 17.300 85.340 ;
        RECT 19.935 85.170 20.105 85.340 ;
        RECT 20.895 85.170 21.065 85.340 ;
        RECT 21.855 85.170 22.025 85.340 ;
        RECT 22.815 85.170 22.985 85.340 ;
        RECT 23.775 85.170 23.945 85.340 ;
        RECT 24.735 85.170 24.905 85.340 ;
        RECT 1.565 82.110 1.735 82.280 ;
        RECT 1.565 81.750 1.735 81.920 ;
        RECT 1.565 81.390 1.735 81.560 ;
        RECT 2.525 82.110 2.695 82.280 ;
        RECT 2.525 81.750 2.695 81.920 ;
        RECT 2.525 81.390 2.695 81.560 ;
        RECT 3.485 82.110 3.655 82.280 ;
        RECT 3.485 81.750 3.655 81.920 ;
        RECT 3.485 81.390 3.655 81.560 ;
        RECT 4.445 82.110 4.615 82.280 ;
        RECT 4.445 81.750 4.615 81.920 ;
        RECT 4.445 81.390 4.615 81.560 ;
        RECT 5.405 82.110 5.575 82.280 ;
        RECT 5.405 81.750 5.575 81.920 ;
        RECT 5.405 81.390 5.575 81.560 ;
        RECT 6.365 82.110 6.535 82.280 ;
        RECT 6.365 81.750 6.535 81.920 ;
        RECT 6.365 81.390 6.535 81.560 ;
        RECT 12.330 82.130 12.500 82.300 ;
        RECT 12.330 81.770 12.500 81.940 ;
        RECT 12.330 81.410 12.500 81.580 ;
        RECT 12.810 82.130 12.980 82.300 ;
        RECT 12.810 81.770 12.980 81.940 ;
        RECT 12.810 81.410 12.980 81.580 ;
        RECT 13.290 82.130 13.460 82.300 ;
        RECT 13.290 81.770 13.460 81.940 ;
        RECT 13.290 81.410 13.460 81.580 ;
        RECT 13.770 82.130 13.940 82.300 ;
        RECT 13.770 81.770 13.940 81.940 ;
        RECT 13.770 81.410 13.940 81.580 ;
        RECT 14.250 82.130 14.420 82.300 ;
        RECT 14.250 81.770 14.420 81.940 ;
        RECT 14.250 81.410 14.420 81.580 ;
        RECT 14.730 82.130 14.900 82.300 ;
        RECT 14.730 81.770 14.900 81.940 ;
        RECT 14.730 81.410 14.900 81.580 ;
        RECT 15.210 82.130 15.380 82.300 ;
        RECT 15.210 81.770 15.380 81.940 ;
        RECT 15.210 81.410 15.380 81.580 ;
        RECT 15.690 82.130 15.860 82.300 ;
        RECT 15.690 81.770 15.860 81.940 ;
        RECT 15.690 81.410 15.860 81.580 ;
        RECT 16.170 82.130 16.340 82.300 ;
        RECT 16.170 81.770 16.340 81.940 ;
        RECT 16.170 81.410 16.340 81.580 ;
        RECT 16.650 82.130 16.820 82.300 ;
        RECT 16.650 81.770 16.820 81.940 ;
        RECT 16.650 81.410 16.820 81.580 ;
        RECT 17.130 82.130 17.300 82.300 ;
        RECT 17.130 81.770 17.300 81.940 ;
        RECT 17.130 81.410 17.300 81.580 ;
        RECT 20.415 82.130 20.585 82.300 ;
        RECT 20.415 81.770 20.585 81.940 ;
        RECT 20.415 81.410 20.585 81.580 ;
        RECT 21.375 82.130 21.545 82.300 ;
        RECT 21.375 81.770 21.545 81.940 ;
        RECT 21.375 81.410 21.545 81.580 ;
        RECT 22.335 82.130 22.505 82.300 ;
        RECT 22.335 81.770 22.505 81.940 ;
        RECT 22.335 81.410 22.505 81.580 ;
        RECT 23.295 82.130 23.465 82.300 ;
        RECT 23.295 81.770 23.465 81.940 ;
        RECT 23.295 81.410 23.465 81.580 ;
        RECT 24.255 82.130 24.425 82.300 ;
        RECT 24.255 81.770 24.425 81.940 ;
        RECT 24.255 81.410 24.425 81.580 ;
        RECT 26.740 80.050 26.910 80.220 ;
        RECT 1.565 79.270 1.735 79.440 ;
        RECT 2.525 79.270 2.695 79.440 ;
        RECT 3.485 79.270 3.655 79.440 ;
        RECT 4.445 79.270 4.615 79.440 ;
        RECT 5.405 79.270 5.575 79.440 ;
        RECT 6.365 79.270 6.535 79.440 ;
        RECT 12.330 79.290 12.500 79.460 ;
        RECT 12.810 79.290 12.980 79.460 ;
        RECT 13.290 79.290 13.460 79.460 ;
        RECT 13.770 79.290 13.940 79.460 ;
        RECT 14.250 79.290 14.420 79.460 ;
        RECT 14.730 79.290 14.900 79.460 ;
        RECT 15.210 79.290 15.380 79.460 ;
        RECT 15.690 79.290 15.860 79.460 ;
        RECT 16.170 79.290 16.340 79.460 ;
        RECT 16.650 79.290 16.820 79.460 ;
        RECT 17.130 79.290 17.300 79.460 ;
        RECT 18.675 79.215 18.845 79.595 ;
        RECT 20.415 79.290 20.585 79.460 ;
        RECT 21.375 79.290 21.545 79.460 ;
        RECT 22.335 79.290 22.505 79.460 ;
        RECT 23.295 79.290 23.465 79.460 ;
        RECT 24.255 79.290 24.425 79.460 ;
        RECT 12.330 78.735 12.500 78.905 ;
        RECT 13.290 78.735 13.460 78.905 ;
        RECT 14.250 78.735 14.420 78.905 ;
        RECT 15.210 78.735 15.380 78.905 ;
        RECT 16.170 78.735 16.340 78.905 ;
        RECT 17.130 78.735 17.300 78.905 ;
        RECT 19.935 78.735 20.105 78.905 ;
        RECT 20.895 78.735 21.065 78.905 ;
        RECT 21.855 78.735 22.025 78.905 ;
        RECT 22.815 78.735 22.985 78.905 ;
        RECT 23.775 78.735 23.945 78.905 ;
        RECT 24.735 78.735 24.905 78.905 ;
        RECT 1.565 75.675 1.735 75.845 ;
        RECT 1.565 75.315 1.735 75.485 ;
        RECT 1.565 74.955 1.735 75.125 ;
        RECT 2.525 75.675 2.695 75.845 ;
        RECT 2.525 75.315 2.695 75.485 ;
        RECT 2.525 74.955 2.695 75.125 ;
        RECT 3.485 75.675 3.655 75.845 ;
        RECT 3.485 75.315 3.655 75.485 ;
        RECT 3.485 74.955 3.655 75.125 ;
        RECT 4.445 75.675 4.615 75.845 ;
        RECT 4.445 75.315 4.615 75.485 ;
        RECT 4.445 74.955 4.615 75.125 ;
        RECT 5.405 75.675 5.575 75.845 ;
        RECT 5.405 75.315 5.575 75.485 ;
        RECT 5.405 74.955 5.575 75.125 ;
        RECT 6.365 75.675 6.535 75.845 ;
        RECT 6.365 75.315 6.535 75.485 ;
        RECT 6.365 74.955 6.535 75.125 ;
        RECT 12.330 75.695 12.500 75.865 ;
        RECT 12.330 75.335 12.500 75.505 ;
        RECT 12.330 74.975 12.500 75.145 ;
        RECT 12.810 75.695 12.980 75.865 ;
        RECT 12.810 75.335 12.980 75.505 ;
        RECT 12.810 74.975 12.980 75.145 ;
        RECT 13.290 75.695 13.460 75.865 ;
        RECT 13.290 75.335 13.460 75.505 ;
        RECT 13.290 74.975 13.460 75.145 ;
        RECT 13.770 75.695 13.940 75.865 ;
        RECT 13.770 75.335 13.940 75.505 ;
        RECT 13.770 74.975 13.940 75.145 ;
        RECT 14.250 75.695 14.420 75.865 ;
        RECT 14.250 75.335 14.420 75.505 ;
        RECT 14.250 74.975 14.420 75.145 ;
        RECT 14.730 75.695 14.900 75.865 ;
        RECT 14.730 75.335 14.900 75.505 ;
        RECT 14.730 74.975 14.900 75.145 ;
        RECT 15.210 75.695 15.380 75.865 ;
        RECT 15.210 75.335 15.380 75.505 ;
        RECT 15.210 74.975 15.380 75.145 ;
        RECT 15.690 75.695 15.860 75.865 ;
        RECT 15.690 75.335 15.860 75.505 ;
        RECT 15.690 74.975 15.860 75.145 ;
        RECT 16.170 75.695 16.340 75.865 ;
        RECT 16.170 75.335 16.340 75.505 ;
        RECT 16.170 74.975 16.340 75.145 ;
        RECT 16.650 75.695 16.820 75.865 ;
        RECT 16.650 75.335 16.820 75.505 ;
        RECT 16.650 74.975 16.820 75.145 ;
        RECT 17.130 75.695 17.300 75.865 ;
        RECT 17.130 75.335 17.300 75.505 ;
        RECT 17.130 74.975 17.300 75.145 ;
        RECT 20.415 75.695 20.585 75.865 ;
        RECT 20.415 75.335 20.585 75.505 ;
        RECT 20.415 74.975 20.585 75.145 ;
        RECT 21.375 75.695 21.545 75.865 ;
        RECT 21.375 75.335 21.545 75.505 ;
        RECT 21.375 74.975 21.545 75.145 ;
        RECT 22.335 75.695 22.505 75.865 ;
        RECT 22.335 75.335 22.505 75.505 ;
        RECT 22.335 74.975 22.505 75.145 ;
        RECT 23.295 75.695 23.465 75.865 ;
        RECT 23.295 75.335 23.465 75.505 ;
        RECT 23.295 74.975 23.465 75.145 ;
        RECT 24.255 75.695 24.425 75.865 ;
        RECT 24.255 75.335 24.425 75.505 ;
        RECT 24.255 74.975 24.425 75.145 ;
        RECT 26.740 73.615 26.910 73.785 ;
        RECT 1.565 72.835 1.735 73.005 ;
        RECT 2.525 72.835 2.695 73.005 ;
        RECT 3.485 72.835 3.655 73.005 ;
        RECT 4.445 72.835 4.615 73.005 ;
        RECT 5.405 72.835 5.575 73.005 ;
        RECT 6.365 72.835 6.535 73.005 ;
        RECT 12.330 72.855 12.500 73.025 ;
        RECT 12.810 72.855 12.980 73.025 ;
        RECT 13.290 72.855 13.460 73.025 ;
        RECT 13.770 72.855 13.940 73.025 ;
        RECT 14.250 72.855 14.420 73.025 ;
        RECT 14.730 72.855 14.900 73.025 ;
        RECT 15.210 72.855 15.380 73.025 ;
        RECT 15.690 72.855 15.860 73.025 ;
        RECT 16.170 72.855 16.340 73.025 ;
        RECT 16.650 72.855 16.820 73.025 ;
        RECT 17.130 72.855 17.300 73.025 ;
        RECT 18.675 72.780 18.845 73.160 ;
        RECT 20.415 72.855 20.585 73.025 ;
        RECT 21.375 72.855 21.545 73.025 ;
        RECT 22.335 72.855 22.505 73.025 ;
        RECT 23.295 72.855 23.465 73.025 ;
        RECT 24.255 72.855 24.425 73.025 ;
        RECT 12.330 72.300 12.500 72.470 ;
        RECT 13.290 72.300 13.460 72.470 ;
        RECT 14.250 72.300 14.420 72.470 ;
        RECT 15.210 72.300 15.380 72.470 ;
        RECT 16.170 72.300 16.340 72.470 ;
        RECT 17.130 72.300 17.300 72.470 ;
        RECT 19.935 72.300 20.105 72.470 ;
        RECT 20.895 72.300 21.065 72.470 ;
        RECT 21.855 72.300 22.025 72.470 ;
        RECT 22.815 72.300 22.985 72.470 ;
        RECT 23.775 72.300 23.945 72.470 ;
        RECT 24.735 72.300 24.905 72.470 ;
        RECT 1.565 69.240 1.735 69.410 ;
        RECT 1.565 68.880 1.735 69.050 ;
        RECT 1.565 68.520 1.735 68.690 ;
        RECT 2.525 69.240 2.695 69.410 ;
        RECT 2.525 68.880 2.695 69.050 ;
        RECT 2.525 68.520 2.695 68.690 ;
        RECT 3.485 69.240 3.655 69.410 ;
        RECT 3.485 68.880 3.655 69.050 ;
        RECT 3.485 68.520 3.655 68.690 ;
        RECT 4.445 69.240 4.615 69.410 ;
        RECT 4.445 68.880 4.615 69.050 ;
        RECT 4.445 68.520 4.615 68.690 ;
        RECT 5.405 69.240 5.575 69.410 ;
        RECT 5.405 68.880 5.575 69.050 ;
        RECT 5.405 68.520 5.575 68.690 ;
        RECT 6.365 69.240 6.535 69.410 ;
        RECT 6.365 68.880 6.535 69.050 ;
        RECT 6.365 68.520 6.535 68.690 ;
        RECT 12.330 69.260 12.500 69.430 ;
        RECT 12.330 68.900 12.500 69.070 ;
        RECT 12.330 68.540 12.500 68.710 ;
        RECT 12.810 69.260 12.980 69.430 ;
        RECT 12.810 68.900 12.980 69.070 ;
        RECT 12.810 68.540 12.980 68.710 ;
        RECT 13.290 69.260 13.460 69.430 ;
        RECT 13.290 68.900 13.460 69.070 ;
        RECT 13.290 68.540 13.460 68.710 ;
        RECT 13.770 69.260 13.940 69.430 ;
        RECT 13.770 68.900 13.940 69.070 ;
        RECT 13.770 68.540 13.940 68.710 ;
        RECT 14.250 69.260 14.420 69.430 ;
        RECT 14.250 68.900 14.420 69.070 ;
        RECT 14.250 68.540 14.420 68.710 ;
        RECT 14.730 69.260 14.900 69.430 ;
        RECT 14.730 68.900 14.900 69.070 ;
        RECT 14.730 68.540 14.900 68.710 ;
        RECT 15.210 69.260 15.380 69.430 ;
        RECT 15.210 68.900 15.380 69.070 ;
        RECT 15.210 68.540 15.380 68.710 ;
        RECT 15.690 69.260 15.860 69.430 ;
        RECT 15.690 68.900 15.860 69.070 ;
        RECT 15.690 68.540 15.860 68.710 ;
        RECT 16.170 69.260 16.340 69.430 ;
        RECT 16.170 68.900 16.340 69.070 ;
        RECT 16.170 68.540 16.340 68.710 ;
        RECT 16.650 69.260 16.820 69.430 ;
        RECT 16.650 68.900 16.820 69.070 ;
        RECT 16.650 68.540 16.820 68.710 ;
        RECT 17.130 69.260 17.300 69.430 ;
        RECT 17.130 68.900 17.300 69.070 ;
        RECT 17.130 68.540 17.300 68.710 ;
        RECT 20.415 69.260 20.585 69.430 ;
        RECT 20.415 68.900 20.585 69.070 ;
        RECT 20.415 68.540 20.585 68.710 ;
        RECT 21.375 69.260 21.545 69.430 ;
        RECT 21.375 68.900 21.545 69.070 ;
        RECT 21.375 68.540 21.545 68.710 ;
        RECT 22.335 69.260 22.505 69.430 ;
        RECT 22.335 68.900 22.505 69.070 ;
        RECT 22.335 68.540 22.505 68.710 ;
        RECT 23.295 69.260 23.465 69.430 ;
        RECT 23.295 68.900 23.465 69.070 ;
        RECT 23.295 68.540 23.465 68.710 ;
        RECT 24.255 69.260 24.425 69.430 ;
        RECT 24.255 68.900 24.425 69.070 ;
        RECT 24.255 68.540 24.425 68.710 ;
        RECT 26.740 67.180 26.910 67.350 ;
        RECT 1.565 66.400 1.735 66.570 ;
        RECT 2.525 66.400 2.695 66.570 ;
        RECT 3.485 66.400 3.655 66.570 ;
        RECT 4.445 66.400 4.615 66.570 ;
        RECT 5.405 66.400 5.575 66.570 ;
        RECT 6.365 66.400 6.535 66.570 ;
        RECT 12.330 66.420 12.500 66.590 ;
        RECT 12.810 66.420 12.980 66.590 ;
        RECT 13.290 66.420 13.460 66.590 ;
        RECT 13.770 66.420 13.940 66.590 ;
        RECT 14.250 66.420 14.420 66.590 ;
        RECT 14.730 66.420 14.900 66.590 ;
        RECT 15.210 66.420 15.380 66.590 ;
        RECT 15.690 66.420 15.860 66.590 ;
        RECT 16.170 66.420 16.340 66.590 ;
        RECT 16.650 66.420 16.820 66.590 ;
        RECT 17.130 66.420 17.300 66.590 ;
        RECT 18.675 66.345 18.845 66.725 ;
        RECT 20.415 66.420 20.585 66.590 ;
        RECT 21.375 66.420 21.545 66.590 ;
        RECT 22.335 66.420 22.505 66.590 ;
        RECT 23.295 66.420 23.465 66.590 ;
        RECT 24.255 66.420 24.425 66.590 ;
        RECT 12.330 65.865 12.500 66.035 ;
        RECT 13.290 65.865 13.460 66.035 ;
        RECT 14.250 65.865 14.420 66.035 ;
        RECT 15.210 65.865 15.380 66.035 ;
        RECT 16.170 65.865 16.340 66.035 ;
        RECT 17.130 65.865 17.300 66.035 ;
        RECT 19.935 65.865 20.105 66.035 ;
        RECT 20.895 65.865 21.065 66.035 ;
        RECT 21.855 65.865 22.025 66.035 ;
        RECT 22.815 65.865 22.985 66.035 ;
        RECT 23.775 65.865 23.945 66.035 ;
        RECT 24.735 65.865 24.905 66.035 ;
        RECT 1.565 62.805 1.735 62.975 ;
        RECT 1.565 62.445 1.735 62.615 ;
        RECT 1.565 62.085 1.735 62.255 ;
        RECT 2.525 62.805 2.695 62.975 ;
        RECT 2.525 62.445 2.695 62.615 ;
        RECT 2.525 62.085 2.695 62.255 ;
        RECT 3.485 62.805 3.655 62.975 ;
        RECT 3.485 62.445 3.655 62.615 ;
        RECT 3.485 62.085 3.655 62.255 ;
        RECT 4.445 62.805 4.615 62.975 ;
        RECT 4.445 62.445 4.615 62.615 ;
        RECT 4.445 62.085 4.615 62.255 ;
        RECT 5.405 62.805 5.575 62.975 ;
        RECT 5.405 62.445 5.575 62.615 ;
        RECT 5.405 62.085 5.575 62.255 ;
        RECT 6.365 62.805 6.535 62.975 ;
        RECT 6.365 62.445 6.535 62.615 ;
        RECT 6.365 62.085 6.535 62.255 ;
        RECT 12.330 62.825 12.500 62.995 ;
        RECT 12.330 62.465 12.500 62.635 ;
        RECT 12.330 62.105 12.500 62.275 ;
        RECT 12.810 62.825 12.980 62.995 ;
        RECT 12.810 62.465 12.980 62.635 ;
        RECT 12.810 62.105 12.980 62.275 ;
        RECT 13.290 62.825 13.460 62.995 ;
        RECT 13.290 62.465 13.460 62.635 ;
        RECT 13.290 62.105 13.460 62.275 ;
        RECT 13.770 62.825 13.940 62.995 ;
        RECT 13.770 62.465 13.940 62.635 ;
        RECT 13.770 62.105 13.940 62.275 ;
        RECT 14.250 62.825 14.420 62.995 ;
        RECT 14.250 62.465 14.420 62.635 ;
        RECT 14.250 62.105 14.420 62.275 ;
        RECT 14.730 62.825 14.900 62.995 ;
        RECT 14.730 62.465 14.900 62.635 ;
        RECT 14.730 62.105 14.900 62.275 ;
        RECT 15.210 62.825 15.380 62.995 ;
        RECT 15.210 62.465 15.380 62.635 ;
        RECT 15.210 62.105 15.380 62.275 ;
        RECT 15.690 62.825 15.860 62.995 ;
        RECT 15.690 62.465 15.860 62.635 ;
        RECT 15.690 62.105 15.860 62.275 ;
        RECT 16.170 62.825 16.340 62.995 ;
        RECT 16.170 62.465 16.340 62.635 ;
        RECT 16.170 62.105 16.340 62.275 ;
        RECT 16.650 62.825 16.820 62.995 ;
        RECT 16.650 62.465 16.820 62.635 ;
        RECT 16.650 62.105 16.820 62.275 ;
        RECT 17.130 62.825 17.300 62.995 ;
        RECT 17.130 62.465 17.300 62.635 ;
        RECT 17.130 62.105 17.300 62.275 ;
        RECT 20.415 62.825 20.585 62.995 ;
        RECT 20.415 62.465 20.585 62.635 ;
        RECT 20.415 62.105 20.585 62.275 ;
        RECT 21.375 62.825 21.545 62.995 ;
        RECT 21.375 62.465 21.545 62.635 ;
        RECT 21.375 62.105 21.545 62.275 ;
        RECT 22.335 62.825 22.505 62.995 ;
        RECT 22.335 62.465 22.505 62.635 ;
        RECT 22.335 62.105 22.505 62.275 ;
        RECT 23.295 62.825 23.465 62.995 ;
        RECT 23.295 62.465 23.465 62.635 ;
        RECT 23.295 62.105 23.465 62.275 ;
        RECT 24.255 62.825 24.425 62.995 ;
        RECT 24.255 62.465 24.425 62.635 ;
        RECT 24.255 62.105 24.425 62.275 ;
        RECT 26.740 60.745 26.910 60.915 ;
        RECT 1.565 59.965 1.735 60.135 ;
        RECT 2.525 59.965 2.695 60.135 ;
        RECT 3.485 59.965 3.655 60.135 ;
        RECT 4.445 59.965 4.615 60.135 ;
        RECT 5.405 59.965 5.575 60.135 ;
        RECT 6.365 59.965 6.535 60.135 ;
        RECT 12.330 59.985 12.500 60.155 ;
        RECT 12.810 59.985 12.980 60.155 ;
        RECT 13.290 59.985 13.460 60.155 ;
        RECT 13.770 59.985 13.940 60.155 ;
        RECT 14.250 59.985 14.420 60.155 ;
        RECT 14.730 59.985 14.900 60.155 ;
        RECT 15.210 59.985 15.380 60.155 ;
        RECT 15.690 59.985 15.860 60.155 ;
        RECT 16.170 59.985 16.340 60.155 ;
        RECT 16.650 59.985 16.820 60.155 ;
        RECT 17.130 59.985 17.300 60.155 ;
        RECT 18.675 59.910 18.845 60.290 ;
        RECT 20.415 59.985 20.585 60.155 ;
        RECT 21.375 59.985 21.545 60.155 ;
        RECT 22.335 59.985 22.505 60.155 ;
        RECT 23.295 59.985 23.465 60.155 ;
        RECT 24.255 59.985 24.425 60.155 ;
        RECT 12.330 59.430 12.500 59.600 ;
        RECT 13.290 59.430 13.460 59.600 ;
        RECT 14.250 59.430 14.420 59.600 ;
        RECT 15.210 59.430 15.380 59.600 ;
        RECT 16.170 59.430 16.340 59.600 ;
        RECT 17.130 59.430 17.300 59.600 ;
        RECT 19.935 59.430 20.105 59.600 ;
        RECT 20.895 59.430 21.065 59.600 ;
        RECT 21.855 59.430 22.025 59.600 ;
        RECT 22.815 59.430 22.985 59.600 ;
        RECT 23.775 59.430 23.945 59.600 ;
        RECT 24.735 59.430 24.905 59.600 ;
        RECT 1.565 56.370 1.735 56.540 ;
        RECT 1.565 56.010 1.735 56.180 ;
        RECT 1.565 55.650 1.735 55.820 ;
        RECT 2.525 56.370 2.695 56.540 ;
        RECT 2.525 56.010 2.695 56.180 ;
        RECT 2.525 55.650 2.695 55.820 ;
        RECT 3.485 56.370 3.655 56.540 ;
        RECT 3.485 56.010 3.655 56.180 ;
        RECT 3.485 55.650 3.655 55.820 ;
        RECT 4.445 56.370 4.615 56.540 ;
        RECT 4.445 56.010 4.615 56.180 ;
        RECT 4.445 55.650 4.615 55.820 ;
        RECT 5.405 56.370 5.575 56.540 ;
        RECT 5.405 56.010 5.575 56.180 ;
        RECT 5.405 55.650 5.575 55.820 ;
        RECT 6.365 56.370 6.535 56.540 ;
        RECT 6.365 56.010 6.535 56.180 ;
        RECT 6.365 55.650 6.535 55.820 ;
        RECT 12.330 56.390 12.500 56.560 ;
        RECT 12.330 56.030 12.500 56.200 ;
        RECT 12.330 55.670 12.500 55.840 ;
        RECT 12.810 56.390 12.980 56.560 ;
        RECT 12.810 56.030 12.980 56.200 ;
        RECT 12.810 55.670 12.980 55.840 ;
        RECT 13.290 56.390 13.460 56.560 ;
        RECT 13.290 56.030 13.460 56.200 ;
        RECT 13.290 55.670 13.460 55.840 ;
        RECT 13.770 56.390 13.940 56.560 ;
        RECT 13.770 56.030 13.940 56.200 ;
        RECT 13.770 55.670 13.940 55.840 ;
        RECT 14.250 56.390 14.420 56.560 ;
        RECT 14.250 56.030 14.420 56.200 ;
        RECT 14.250 55.670 14.420 55.840 ;
        RECT 14.730 56.390 14.900 56.560 ;
        RECT 14.730 56.030 14.900 56.200 ;
        RECT 14.730 55.670 14.900 55.840 ;
        RECT 15.210 56.390 15.380 56.560 ;
        RECT 15.210 56.030 15.380 56.200 ;
        RECT 15.210 55.670 15.380 55.840 ;
        RECT 15.690 56.390 15.860 56.560 ;
        RECT 15.690 56.030 15.860 56.200 ;
        RECT 15.690 55.670 15.860 55.840 ;
        RECT 16.170 56.390 16.340 56.560 ;
        RECT 16.170 56.030 16.340 56.200 ;
        RECT 16.170 55.670 16.340 55.840 ;
        RECT 16.650 56.390 16.820 56.560 ;
        RECT 16.650 56.030 16.820 56.200 ;
        RECT 16.650 55.670 16.820 55.840 ;
        RECT 17.130 56.390 17.300 56.560 ;
        RECT 17.130 56.030 17.300 56.200 ;
        RECT 17.130 55.670 17.300 55.840 ;
        RECT 20.415 56.390 20.585 56.560 ;
        RECT 20.415 56.030 20.585 56.200 ;
        RECT 20.415 55.670 20.585 55.840 ;
        RECT 21.375 56.390 21.545 56.560 ;
        RECT 21.375 56.030 21.545 56.200 ;
        RECT 21.375 55.670 21.545 55.840 ;
        RECT 22.335 56.390 22.505 56.560 ;
        RECT 22.335 56.030 22.505 56.200 ;
        RECT 22.335 55.670 22.505 55.840 ;
        RECT 23.295 56.390 23.465 56.560 ;
        RECT 23.295 56.030 23.465 56.200 ;
        RECT 23.295 55.670 23.465 55.840 ;
        RECT 24.255 56.390 24.425 56.560 ;
        RECT 24.255 56.030 24.425 56.200 ;
        RECT 24.255 55.670 24.425 55.840 ;
        RECT 26.740 54.310 26.910 54.480 ;
        RECT 1.565 53.530 1.735 53.700 ;
        RECT 2.525 53.530 2.695 53.700 ;
        RECT 3.485 53.530 3.655 53.700 ;
        RECT 4.445 53.530 4.615 53.700 ;
        RECT 5.405 53.530 5.575 53.700 ;
        RECT 6.365 53.530 6.535 53.700 ;
        RECT 12.330 53.550 12.500 53.720 ;
        RECT 12.810 53.550 12.980 53.720 ;
        RECT 13.290 53.550 13.460 53.720 ;
        RECT 13.770 53.550 13.940 53.720 ;
        RECT 14.250 53.550 14.420 53.720 ;
        RECT 14.730 53.550 14.900 53.720 ;
        RECT 15.210 53.550 15.380 53.720 ;
        RECT 15.690 53.550 15.860 53.720 ;
        RECT 16.170 53.550 16.340 53.720 ;
        RECT 16.650 53.550 16.820 53.720 ;
        RECT 17.130 53.550 17.300 53.720 ;
        RECT 18.675 53.475 18.845 53.855 ;
        RECT 20.415 53.550 20.585 53.720 ;
        RECT 21.375 53.550 21.545 53.720 ;
        RECT 22.335 53.550 22.505 53.720 ;
        RECT 23.295 53.550 23.465 53.720 ;
        RECT 24.255 53.550 24.425 53.720 ;
        RECT 12.330 52.995 12.500 53.165 ;
        RECT 13.290 52.995 13.460 53.165 ;
        RECT 14.250 52.995 14.420 53.165 ;
        RECT 15.210 52.995 15.380 53.165 ;
        RECT 16.170 52.995 16.340 53.165 ;
        RECT 17.130 52.995 17.300 53.165 ;
        RECT 19.935 52.995 20.105 53.165 ;
        RECT 20.895 52.995 21.065 53.165 ;
        RECT 21.855 52.995 22.025 53.165 ;
        RECT 22.815 52.995 22.985 53.165 ;
        RECT 23.775 52.995 23.945 53.165 ;
        RECT 24.735 52.995 24.905 53.165 ;
        RECT 1.565 49.935 1.735 50.105 ;
        RECT 1.565 49.575 1.735 49.745 ;
        RECT 1.565 49.215 1.735 49.385 ;
        RECT 2.525 49.935 2.695 50.105 ;
        RECT 2.525 49.575 2.695 49.745 ;
        RECT 2.525 49.215 2.695 49.385 ;
        RECT 3.485 49.935 3.655 50.105 ;
        RECT 3.485 49.575 3.655 49.745 ;
        RECT 3.485 49.215 3.655 49.385 ;
        RECT 4.445 49.935 4.615 50.105 ;
        RECT 4.445 49.575 4.615 49.745 ;
        RECT 4.445 49.215 4.615 49.385 ;
        RECT 5.405 49.935 5.575 50.105 ;
        RECT 5.405 49.575 5.575 49.745 ;
        RECT 5.405 49.215 5.575 49.385 ;
        RECT 6.365 49.935 6.535 50.105 ;
        RECT 6.365 49.575 6.535 49.745 ;
        RECT 6.365 49.215 6.535 49.385 ;
        RECT 12.330 49.955 12.500 50.125 ;
        RECT 12.330 49.595 12.500 49.765 ;
        RECT 12.330 49.235 12.500 49.405 ;
        RECT 12.810 49.955 12.980 50.125 ;
        RECT 12.810 49.595 12.980 49.765 ;
        RECT 12.810 49.235 12.980 49.405 ;
        RECT 13.290 49.955 13.460 50.125 ;
        RECT 13.290 49.595 13.460 49.765 ;
        RECT 13.290 49.235 13.460 49.405 ;
        RECT 13.770 49.955 13.940 50.125 ;
        RECT 13.770 49.595 13.940 49.765 ;
        RECT 13.770 49.235 13.940 49.405 ;
        RECT 14.250 49.955 14.420 50.125 ;
        RECT 14.250 49.595 14.420 49.765 ;
        RECT 14.250 49.235 14.420 49.405 ;
        RECT 14.730 49.955 14.900 50.125 ;
        RECT 14.730 49.595 14.900 49.765 ;
        RECT 14.730 49.235 14.900 49.405 ;
        RECT 15.210 49.955 15.380 50.125 ;
        RECT 15.210 49.595 15.380 49.765 ;
        RECT 15.210 49.235 15.380 49.405 ;
        RECT 15.690 49.955 15.860 50.125 ;
        RECT 15.690 49.595 15.860 49.765 ;
        RECT 15.690 49.235 15.860 49.405 ;
        RECT 16.170 49.955 16.340 50.125 ;
        RECT 16.170 49.595 16.340 49.765 ;
        RECT 16.170 49.235 16.340 49.405 ;
        RECT 16.650 49.955 16.820 50.125 ;
        RECT 16.650 49.595 16.820 49.765 ;
        RECT 16.650 49.235 16.820 49.405 ;
        RECT 17.130 49.955 17.300 50.125 ;
        RECT 17.130 49.595 17.300 49.765 ;
        RECT 17.130 49.235 17.300 49.405 ;
        RECT 20.415 49.955 20.585 50.125 ;
        RECT 20.415 49.595 20.585 49.765 ;
        RECT 20.415 49.235 20.585 49.405 ;
        RECT 21.375 49.955 21.545 50.125 ;
        RECT 21.375 49.595 21.545 49.765 ;
        RECT 21.375 49.235 21.545 49.405 ;
        RECT 22.335 49.955 22.505 50.125 ;
        RECT 22.335 49.595 22.505 49.765 ;
        RECT 22.335 49.235 22.505 49.405 ;
        RECT 23.295 49.955 23.465 50.125 ;
        RECT 23.295 49.595 23.465 49.765 ;
        RECT 23.295 49.235 23.465 49.405 ;
        RECT 24.255 49.955 24.425 50.125 ;
        RECT 24.255 49.595 24.425 49.765 ;
        RECT 24.255 49.235 24.425 49.405 ;
        RECT 26.740 47.875 26.910 48.045 ;
        RECT 1.565 47.095 1.735 47.265 ;
        RECT 2.525 47.095 2.695 47.265 ;
        RECT 3.485 47.095 3.655 47.265 ;
        RECT 4.445 47.095 4.615 47.265 ;
        RECT 5.405 47.095 5.575 47.265 ;
        RECT 6.365 47.095 6.535 47.265 ;
        RECT 12.330 47.115 12.500 47.285 ;
        RECT 12.810 47.115 12.980 47.285 ;
        RECT 13.290 47.115 13.460 47.285 ;
        RECT 13.770 47.115 13.940 47.285 ;
        RECT 14.250 47.115 14.420 47.285 ;
        RECT 14.730 47.115 14.900 47.285 ;
        RECT 15.210 47.115 15.380 47.285 ;
        RECT 15.690 47.115 15.860 47.285 ;
        RECT 16.170 47.115 16.340 47.285 ;
        RECT 16.650 47.115 16.820 47.285 ;
        RECT 17.130 47.115 17.300 47.285 ;
        RECT 18.675 47.040 18.845 47.420 ;
        RECT 20.415 47.115 20.585 47.285 ;
        RECT 21.375 47.115 21.545 47.285 ;
        RECT 22.335 47.115 22.505 47.285 ;
        RECT 23.295 47.115 23.465 47.285 ;
        RECT 24.255 47.115 24.425 47.285 ;
        RECT 12.330 46.560 12.500 46.730 ;
        RECT 13.290 46.560 13.460 46.730 ;
        RECT 14.250 46.560 14.420 46.730 ;
        RECT 15.210 46.560 15.380 46.730 ;
        RECT 16.170 46.560 16.340 46.730 ;
        RECT 17.130 46.560 17.300 46.730 ;
        RECT 19.935 46.560 20.105 46.730 ;
        RECT 20.895 46.560 21.065 46.730 ;
        RECT 21.855 46.560 22.025 46.730 ;
        RECT 22.815 46.560 22.985 46.730 ;
        RECT 23.775 46.560 23.945 46.730 ;
        RECT 24.735 46.560 24.905 46.730 ;
        RECT 1.565 43.500 1.735 43.670 ;
        RECT 1.565 43.140 1.735 43.310 ;
        RECT 1.565 42.780 1.735 42.950 ;
        RECT 2.525 43.500 2.695 43.670 ;
        RECT 2.525 43.140 2.695 43.310 ;
        RECT 2.525 42.780 2.695 42.950 ;
        RECT 3.485 43.500 3.655 43.670 ;
        RECT 3.485 43.140 3.655 43.310 ;
        RECT 3.485 42.780 3.655 42.950 ;
        RECT 4.445 43.500 4.615 43.670 ;
        RECT 4.445 43.140 4.615 43.310 ;
        RECT 4.445 42.780 4.615 42.950 ;
        RECT 5.405 43.500 5.575 43.670 ;
        RECT 5.405 43.140 5.575 43.310 ;
        RECT 5.405 42.780 5.575 42.950 ;
        RECT 6.365 43.500 6.535 43.670 ;
        RECT 6.365 43.140 6.535 43.310 ;
        RECT 6.365 42.780 6.535 42.950 ;
        RECT 12.330 43.520 12.500 43.690 ;
        RECT 12.330 43.160 12.500 43.330 ;
        RECT 12.330 42.800 12.500 42.970 ;
        RECT 12.810 43.520 12.980 43.690 ;
        RECT 12.810 43.160 12.980 43.330 ;
        RECT 12.810 42.800 12.980 42.970 ;
        RECT 13.290 43.520 13.460 43.690 ;
        RECT 13.290 43.160 13.460 43.330 ;
        RECT 13.290 42.800 13.460 42.970 ;
        RECT 13.770 43.520 13.940 43.690 ;
        RECT 13.770 43.160 13.940 43.330 ;
        RECT 13.770 42.800 13.940 42.970 ;
        RECT 14.250 43.520 14.420 43.690 ;
        RECT 14.250 43.160 14.420 43.330 ;
        RECT 14.250 42.800 14.420 42.970 ;
        RECT 14.730 43.520 14.900 43.690 ;
        RECT 14.730 43.160 14.900 43.330 ;
        RECT 14.730 42.800 14.900 42.970 ;
        RECT 15.210 43.520 15.380 43.690 ;
        RECT 15.210 43.160 15.380 43.330 ;
        RECT 15.210 42.800 15.380 42.970 ;
        RECT 15.690 43.520 15.860 43.690 ;
        RECT 15.690 43.160 15.860 43.330 ;
        RECT 15.690 42.800 15.860 42.970 ;
        RECT 16.170 43.520 16.340 43.690 ;
        RECT 16.170 43.160 16.340 43.330 ;
        RECT 16.170 42.800 16.340 42.970 ;
        RECT 16.650 43.520 16.820 43.690 ;
        RECT 16.650 43.160 16.820 43.330 ;
        RECT 16.650 42.800 16.820 42.970 ;
        RECT 17.130 43.520 17.300 43.690 ;
        RECT 17.130 43.160 17.300 43.330 ;
        RECT 17.130 42.800 17.300 42.970 ;
        RECT 20.415 43.520 20.585 43.690 ;
        RECT 20.415 43.160 20.585 43.330 ;
        RECT 20.415 42.800 20.585 42.970 ;
        RECT 21.375 43.520 21.545 43.690 ;
        RECT 21.375 43.160 21.545 43.330 ;
        RECT 21.375 42.800 21.545 42.970 ;
        RECT 22.335 43.520 22.505 43.690 ;
        RECT 22.335 43.160 22.505 43.330 ;
        RECT 22.335 42.800 22.505 42.970 ;
        RECT 23.295 43.520 23.465 43.690 ;
        RECT 23.295 43.160 23.465 43.330 ;
        RECT 23.295 42.800 23.465 42.970 ;
        RECT 24.255 43.520 24.425 43.690 ;
        RECT 24.255 43.160 24.425 43.330 ;
        RECT 24.255 42.800 24.425 42.970 ;
        RECT 26.740 41.440 26.910 41.610 ;
        RECT 1.565 40.660 1.735 40.830 ;
        RECT 2.525 40.660 2.695 40.830 ;
        RECT 3.485 40.660 3.655 40.830 ;
        RECT 4.445 40.660 4.615 40.830 ;
        RECT 5.405 40.660 5.575 40.830 ;
        RECT 6.365 40.660 6.535 40.830 ;
        RECT 12.330 40.680 12.500 40.850 ;
        RECT 12.810 40.680 12.980 40.850 ;
        RECT 13.290 40.680 13.460 40.850 ;
        RECT 13.770 40.680 13.940 40.850 ;
        RECT 14.250 40.680 14.420 40.850 ;
        RECT 14.730 40.680 14.900 40.850 ;
        RECT 15.210 40.680 15.380 40.850 ;
        RECT 15.690 40.680 15.860 40.850 ;
        RECT 16.170 40.680 16.340 40.850 ;
        RECT 16.650 40.680 16.820 40.850 ;
        RECT 17.130 40.680 17.300 40.850 ;
        RECT 18.675 40.605 18.845 40.985 ;
        RECT 20.415 40.680 20.585 40.850 ;
        RECT 21.375 40.680 21.545 40.850 ;
        RECT 22.335 40.680 22.505 40.850 ;
        RECT 23.295 40.680 23.465 40.850 ;
        RECT 24.255 40.680 24.425 40.850 ;
        RECT 12.330 40.125 12.500 40.295 ;
        RECT 13.290 40.125 13.460 40.295 ;
        RECT 14.250 40.125 14.420 40.295 ;
        RECT 15.210 40.125 15.380 40.295 ;
        RECT 16.170 40.125 16.340 40.295 ;
        RECT 17.130 40.125 17.300 40.295 ;
        RECT 19.935 40.125 20.105 40.295 ;
        RECT 20.895 40.125 21.065 40.295 ;
        RECT 21.855 40.125 22.025 40.295 ;
        RECT 22.815 40.125 22.985 40.295 ;
        RECT 23.775 40.125 23.945 40.295 ;
        RECT 24.735 40.125 24.905 40.295 ;
        RECT 1.565 37.065 1.735 37.235 ;
        RECT 1.565 36.705 1.735 36.875 ;
        RECT 1.565 36.345 1.735 36.515 ;
        RECT 2.525 37.065 2.695 37.235 ;
        RECT 2.525 36.705 2.695 36.875 ;
        RECT 2.525 36.345 2.695 36.515 ;
        RECT 3.485 37.065 3.655 37.235 ;
        RECT 3.485 36.705 3.655 36.875 ;
        RECT 3.485 36.345 3.655 36.515 ;
        RECT 4.445 37.065 4.615 37.235 ;
        RECT 4.445 36.705 4.615 36.875 ;
        RECT 4.445 36.345 4.615 36.515 ;
        RECT 5.405 37.065 5.575 37.235 ;
        RECT 5.405 36.705 5.575 36.875 ;
        RECT 5.405 36.345 5.575 36.515 ;
        RECT 6.365 37.065 6.535 37.235 ;
        RECT 6.365 36.705 6.535 36.875 ;
        RECT 6.365 36.345 6.535 36.515 ;
        RECT 12.330 37.085 12.500 37.255 ;
        RECT 12.330 36.725 12.500 36.895 ;
        RECT 12.330 36.365 12.500 36.535 ;
        RECT 12.810 37.085 12.980 37.255 ;
        RECT 12.810 36.725 12.980 36.895 ;
        RECT 12.810 36.365 12.980 36.535 ;
        RECT 13.290 37.085 13.460 37.255 ;
        RECT 13.290 36.725 13.460 36.895 ;
        RECT 13.290 36.365 13.460 36.535 ;
        RECT 13.770 37.085 13.940 37.255 ;
        RECT 13.770 36.725 13.940 36.895 ;
        RECT 13.770 36.365 13.940 36.535 ;
        RECT 14.250 37.085 14.420 37.255 ;
        RECT 14.250 36.725 14.420 36.895 ;
        RECT 14.250 36.365 14.420 36.535 ;
        RECT 14.730 37.085 14.900 37.255 ;
        RECT 14.730 36.725 14.900 36.895 ;
        RECT 14.730 36.365 14.900 36.535 ;
        RECT 15.210 37.085 15.380 37.255 ;
        RECT 15.210 36.725 15.380 36.895 ;
        RECT 15.210 36.365 15.380 36.535 ;
        RECT 15.690 37.085 15.860 37.255 ;
        RECT 15.690 36.725 15.860 36.895 ;
        RECT 15.690 36.365 15.860 36.535 ;
        RECT 16.170 37.085 16.340 37.255 ;
        RECT 16.170 36.725 16.340 36.895 ;
        RECT 16.170 36.365 16.340 36.535 ;
        RECT 16.650 37.085 16.820 37.255 ;
        RECT 16.650 36.725 16.820 36.895 ;
        RECT 16.650 36.365 16.820 36.535 ;
        RECT 17.130 37.085 17.300 37.255 ;
        RECT 17.130 36.725 17.300 36.895 ;
        RECT 17.130 36.365 17.300 36.535 ;
        RECT 20.415 37.085 20.585 37.255 ;
        RECT 20.415 36.725 20.585 36.895 ;
        RECT 20.415 36.365 20.585 36.535 ;
        RECT 21.375 37.085 21.545 37.255 ;
        RECT 21.375 36.725 21.545 36.895 ;
        RECT 21.375 36.365 21.545 36.535 ;
        RECT 22.335 37.085 22.505 37.255 ;
        RECT 22.335 36.725 22.505 36.895 ;
        RECT 22.335 36.365 22.505 36.535 ;
        RECT 23.295 37.085 23.465 37.255 ;
        RECT 23.295 36.725 23.465 36.895 ;
        RECT 23.295 36.365 23.465 36.535 ;
        RECT 24.255 37.085 24.425 37.255 ;
        RECT 24.255 36.725 24.425 36.895 ;
        RECT 24.255 36.365 24.425 36.535 ;
        RECT 26.740 35.005 26.910 35.175 ;
        RECT 1.565 34.225 1.735 34.395 ;
        RECT 2.525 34.225 2.695 34.395 ;
        RECT 3.485 34.225 3.655 34.395 ;
        RECT 4.445 34.225 4.615 34.395 ;
        RECT 5.405 34.225 5.575 34.395 ;
        RECT 6.365 34.225 6.535 34.395 ;
        RECT 12.330 34.245 12.500 34.415 ;
        RECT 12.810 34.245 12.980 34.415 ;
        RECT 13.290 34.245 13.460 34.415 ;
        RECT 13.770 34.245 13.940 34.415 ;
        RECT 14.250 34.245 14.420 34.415 ;
        RECT 14.730 34.245 14.900 34.415 ;
        RECT 15.210 34.245 15.380 34.415 ;
        RECT 15.690 34.245 15.860 34.415 ;
        RECT 16.170 34.245 16.340 34.415 ;
        RECT 16.650 34.245 16.820 34.415 ;
        RECT 17.130 34.245 17.300 34.415 ;
        RECT 18.675 34.170 18.845 34.550 ;
        RECT 20.415 34.245 20.585 34.415 ;
        RECT 21.375 34.245 21.545 34.415 ;
        RECT 22.335 34.245 22.505 34.415 ;
        RECT 23.295 34.245 23.465 34.415 ;
        RECT 24.255 34.245 24.425 34.415 ;
        RECT 12.330 33.690 12.500 33.860 ;
        RECT 13.290 33.690 13.460 33.860 ;
        RECT 14.250 33.690 14.420 33.860 ;
        RECT 15.210 33.690 15.380 33.860 ;
        RECT 16.170 33.690 16.340 33.860 ;
        RECT 17.130 33.690 17.300 33.860 ;
        RECT 19.935 33.690 20.105 33.860 ;
        RECT 20.895 33.690 21.065 33.860 ;
        RECT 21.855 33.690 22.025 33.860 ;
        RECT 22.815 33.690 22.985 33.860 ;
        RECT 23.775 33.690 23.945 33.860 ;
        RECT 24.735 33.690 24.905 33.860 ;
        RECT 1.565 30.630 1.735 30.800 ;
        RECT 1.565 30.270 1.735 30.440 ;
        RECT 1.565 29.910 1.735 30.080 ;
        RECT 2.525 30.630 2.695 30.800 ;
        RECT 2.525 30.270 2.695 30.440 ;
        RECT 2.525 29.910 2.695 30.080 ;
        RECT 3.485 30.630 3.655 30.800 ;
        RECT 3.485 30.270 3.655 30.440 ;
        RECT 3.485 29.910 3.655 30.080 ;
        RECT 4.445 30.630 4.615 30.800 ;
        RECT 4.445 30.270 4.615 30.440 ;
        RECT 4.445 29.910 4.615 30.080 ;
        RECT 5.405 30.630 5.575 30.800 ;
        RECT 5.405 30.270 5.575 30.440 ;
        RECT 5.405 29.910 5.575 30.080 ;
        RECT 6.365 30.630 6.535 30.800 ;
        RECT 6.365 30.270 6.535 30.440 ;
        RECT 6.365 29.910 6.535 30.080 ;
        RECT 12.330 30.650 12.500 30.820 ;
        RECT 12.330 30.290 12.500 30.460 ;
        RECT 12.330 29.930 12.500 30.100 ;
        RECT 12.810 30.650 12.980 30.820 ;
        RECT 12.810 30.290 12.980 30.460 ;
        RECT 12.810 29.930 12.980 30.100 ;
        RECT 13.290 30.650 13.460 30.820 ;
        RECT 13.290 30.290 13.460 30.460 ;
        RECT 13.290 29.930 13.460 30.100 ;
        RECT 13.770 30.650 13.940 30.820 ;
        RECT 13.770 30.290 13.940 30.460 ;
        RECT 13.770 29.930 13.940 30.100 ;
        RECT 14.250 30.650 14.420 30.820 ;
        RECT 14.250 30.290 14.420 30.460 ;
        RECT 14.250 29.930 14.420 30.100 ;
        RECT 14.730 30.650 14.900 30.820 ;
        RECT 14.730 30.290 14.900 30.460 ;
        RECT 14.730 29.930 14.900 30.100 ;
        RECT 15.210 30.650 15.380 30.820 ;
        RECT 15.210 30.290 15.380 30.460 ;
        RECT 15.210 29.930 15.380 30.100 ;
        RECT 15.690 30.650 15.860 30.820 ;
        RECT 15.690 30.290 15.860 30.460 ;
        RECT 15.690 29.930 15.860 30.100 ;
        RECT 16.170 30.650 16.340 30.820 ;
        RECT 16.170 30.290 16.340 30.460 ;
        RECT 16.170 29.930 16.340 30.100 ;
        RECT 16.650 30.650 16.820 30.820 ;
        RECT 16.650 30.290 16.820 30.460 ;
        RECT 16.650 29.930 16.820 30.100 ;
        RECT 17.130 30.650 17.300 30.820 ;
        RECT 17.130 30.290 17.300 30.460 ;
        RECT 17.130 29.930 17.300 30.100 ;
        RECT 20.415 30.650 20.585 30.820 ;
        RECT 20.415 30.290 20.585 30.460 ;
        RECT 20.415 29.930 20.585 30.100 ;
        RECT 21.375 30.650 21.545 30.820 ;
        RECT 21.375 30.290 21.545 30.460 ;
        RECT 21.375 29.930 21.545 30.100 ;
        RECT 22.335 30.650 22.505 30.820 ;
        RECT 22.335 30.290 22.505 30.460 ;
        RECT 22.335 29.930 22.505 30.100 ;
        RECT 23.295 30.650 23.465 30.820 ;
        RECT 23.295 30.290 23.465 30.460 ;
        RECT 23.295 29.930 23.465 30.100 ;
        RECT 24.255 30.650 24.425 30.820 ;
        RECT 24.255 30.290 24.425 30.460 ;
        RECT 24.255 29.930 24.425 30.100 ;
        RECT 26.740 28.570 26.910 28.740 ;
        RECT 1.565 27.790 1.735 27.960 ;
        RECT 2.525 27.790 2.695 27.960 ;
        RECT 3.485 27.790 3.655 27.960 ;
        RECT 4.445 27.790 4.615 27.960 ;
        RECT 5.405 27.790 5.575 27.960 ;
        RECT 6.365 27.790 6.535 27.960 ;
        RECT 12.330 27.810 12.500 27.980 ;
        RECT 12.810 27.810 12.980 27.980 ;
        RECT 13.290 27.810 13.460 27.980 ;
        RECT 13.770 27.810 13.940 27.980 ;
        RECT 14.250 27.810 14.420 27.980 ;
        RECT 14.730 27.810 14.900 27.980 ;
        RECT 15.210 27.810 15.380 27.980 ;
        RECT 15.690 27.810 15.860 27.980 ;
        RECT 16.170 27.810 16.340 27.980 ;
        RECT 16.650 27.810 16.820 27.980 ;
        RECT 17.130 27.810 17.300 27.980 ;
        RECT 18.675 27.735 18.845 28.115 ;
        RECT 20.415 27.810 20.585 27.980 ;
        RECT 21.375 27.810 21.545 27.980 ;
        RECT 22.335 27.810 22.505 27.980 ;
        RECT 23.295 27.810 23.465 27.980 ;
        RECT 24.255 27.810 24.425 27.980 ;
        RECT 12.330 27.255 12.500 27.425 ;
        RECT 13.290 27.255 13.460 27.425 ;
        RECT 14.250 27.255 14.420 27.425 ;
        RECT 15.210 27.255 15.380 27.425 ;
        RECT 16.170 27.255 16.340 27.425 ;
        RECT 17.130 27.255 17.300 27.425 ;
        RECT 19.935 27.255 20.105 27.425 ;
        RECT 20.895 27.255 21.065 27.425 ;
        RECT 21.855 27.255 22.025 27.425 ;
        RECT 22.815 27.255 22.985 27.425 ;
        RECT 23.775 27.255 23.945 27.425 ;
        RECT 24.735 27.255 24.905 27.425 ;
        RECT 1.565 24.195 1.735 24.365 ;
        RECT 1.565 23.835 1.735 24.005 ;
        RECT 1.565 23.475 1.735 23.645 ;
        RECT 2.525 24.195 2.695 24.365 ;
        RECT 2.525 23.835 2.695 24.005 ;
        RECT 2.525 23.475 2.695 23.645 ;
        RECT 3.485 24.195 3.655 24.365 ;
        RECT 3.485 23.835 3.655 24.005 ;
        RECT 3.485 23.475 3.655 23.645 ;
        RECT 4.445 24.195 4.615 24.365 ;
        RECT 4.445 23.835 4.615 24.005 ;
        RECT 4.445 23.475 4.615 23.645 ;
        RECT 5.405 24.195 5.575 24.365 ;
        RECT 5.405 23.835 5.575 24.005 ;
        RECT 5.405 23.475 5.575 23.645 ;
        RECT 6.365 24.195 6.535 24.365 ;
        RECT 6.365 23.835 6.535 24.005 ;
        RECT 6.365 23.475 6.535 23.645 ;
        RECT 12.330 24.215 12.500 24.385 ;
        RECT 12.330 23.855 12.500 24.025 ;
        RECT 12.330 23.495 12.500 23.665 ;
        RECT 12.810 24.215 12.980 24.385 ;
        RECT 12.810 23.855 12.980 24.025 ;
        RECT 12.810 23.495 12.980 23.665 ;
        RECT 13.290 24.215 13.460 24.385 ;
        RECT 13.290 23.855 13.460 24.025 ;
        RECT 13.290 23.495 13.460 23.665 ;
        RECT 13.770 24.215 13.940 24.385 ;
        RECT 13.770 23.855 13.940 24.025 ;
        RECT 13.770 23.495 13.940 23.665 ;
        RECT 14.250 24.215 14.420 24.385 ;
        RECT 14.250 23.855 14.420 24.025 ;
        RECT 14.250 23.495 14.420 23.665 ;
        RECT 14.730 24.215 14.900 24.385 ;
        RECT 14.730 23.855 14.900 24.025 ;
        RECT 14.730 23.495 14.900 23.665 ;
        RECT 15.210 24.215 15.380 24.385 ;
        RECT 15.210 23.855 15.380 24.025 ;
        RECT 15.210 23.495 15.380 23.665 ;
        RECT 15.690 24.215 15.860 24.385 ;
        RECT 15.690 23.855 15.860 24.025 ;
        RECT 15.690 23.495 15.860 23.665 ;
        RECT 16.170 24.215 16.340 24.385 ;
        RECT 16.170 23.855 16.340 24.025 ;
        RECT 16.170 23.495 16.340 23.665 ;
        RECT 16.650 24.215 16.820 24.385 ;
        RECT 16.650 23.855 16.820 24.025 ;
        RECT 16.650 23.495 16.820 23.665 ;
        RECT 17.130 24.215 17.300 24.385 ;
        RECT 17.130 23.855 17.300 24.025 ;
        RECT 17.130 23.495 17.300 23.665 ;
        RECT 20.415 24.215 20.585 24.385 ;
        RECT 20.415 23.855 20.585 24.025 ;
        RECT 20.415 23.495 20.585 23.665 ;
        RECT 21.375 24.215 21.545 24.385 ;
        RECT 21.375 23.855 21.545 24.025 ;
        RECT 21.375 23.495 21.545 23.665 ;
        RECT 22.335 24.215 22.505 24.385 ;
        RECT 22.335 23.855 22.505 24.025 ;
        RECT 22.335 23.495 22.505 23.665 ;
        RECT 23.295 24.215 23.465 24.385 ;
        RECT 23.295 23.855 23.465 24.025 ;
        RECT 23.295 23.495 23.465 23.665 ;
        RECT 24.255 24.215 24.425 24.385 ;
        RECT 24.255 23.855 24.425 24.025 ;
        RECT 24.255 23.495 24.425 23.665 ;
        RECT 26.740 22.135 26.910 22.305 ;
        RECT 1.565 21.355 1.735 21.525 ;
        RECT 2.525 21.355 2.695 21.525 ;
        RECT 3.485 21.355 3.655 21.525 ;
        RECT 4.445 21.355 4.615 21.525 ;
        RECT 5.405 21.355 5.575 21.525 ;
        RECT 6.365 21.355 6.535 21.525 ;
        RECT 12.330 21.375 12.500 21.545 ;
        RECT 12.810 21.375 12.980 21.545 ;
        RECT 13.290 21.375 13.460 21.545 ;
        RECT 13.770 21.375 13.940 21.545 ;
        RECT 14.250 21.375 14.420 21.545 ;
        RECT 14.730 21.375 14.900 21.545 ;
        RECT 15.210 21.375 15.380 21.545 ;
        RECT 15.690 21.375 15.860 21.545 ;
        RECT 16.170 21.375 16.340 21.545 ;
        RECT 16.650 21.375 16.820 21.545 ;
        RECT 17.130 21.375 17.300 21.545 ;
        RECT 18.675 21.300 18.845 21.680 ;
        RECT 20.415 21.375 20.585 21.545 ;
        RECT 21.375 21.375 21.545 21.545 ;
        RECT 22.335 21.375 22.505 21.545 ;
        RECT 23.295 21.375 23.465 21.545 ;
        RECT 24.255 21.375 24.425 21.545 ;
        RECT 12.330 20.820 12.500 20.990 ;
        RECT 13.290 20.820 13.460 20.990 ;
        RECT 14.250 20.820 14.420 20.990 ;
        RECT 15.210 20.820 15.380 20.990 ;
        RECT 16.170 20.820 16.340 20.990 ;
        RECT 17.130 20.820 17.300 20.990 ;
        RECT 19.935 20.820 20.105 20.990 ;
        RECT 20.895 20.820 21.065 20.990 ;
        RECT 21.855 20.820 22.025 20.990 ;
        RECT 22.815 20.820 22.985 20.990 ;
        RECT 23.775 20.820 23.945 20.990 ;
        RECT 24.735 20.820 24.905 20.990 ;
        RECT 1.565 17.760 1.735 17.930 ;
        RECT 1.565 17.400 1.735 17.570 ;
        RECT 1.565 17.040 1.735 17.210 ;
        RECT 2.525 17.760 2.695 17.930 ;
        RECT 2.525 17.400 2.695 17.570 ;
        RECT 2.525 17.040 2.695 17.210 ;
        RECT 3.485 17.760 3.655 17.930 ;
        RECT 3.485 17.400 3.655 17.570 ;
        RECT 3.485 17.040 3.655 17.210 ;
        RECT 4.445 17.760 4.615 17.930 ;
        RECT 4.445 17.400 4.615 17.570 ;
        RECT 4.445 17.040 4.615 17.210 ;
        RECT 5.405 17.760 5.575 17.930 ;
        RECT 5.405 17.400 5.575 17.570 ;
        RECT 5.405 17.040 5.575 17.210 ;
        RECT 6.365 17.760 6.535 17.930 ;
        RECT 6.365 17.400 6.535 17.570 ;
        RECT 6.365 17.040 6.535 17.210 ;
        RECT 12.330 17.780 12.500 17.950 ;
        RECT 12.330 17.420 12.500 17.590 ;
        RECT 12.330 17.060 12.500 17.230 ;
        RECT 12.810 17.780 12.980 17.950 ;
        RECT 12.810 17.420 12.980 17.590 ;
        RECT 12.810 17.060 12.980 17.230 ;
        RECT 13.290 17.780 13.460 17.950 ;
        RECT 13.290 17.420 13.460 17.590 ;
        RECT 13.290 17.060 13.460 17.230 ;
        RECT 13.770 17.780 13.940 17.950 ;
        RECT 13.770 17.420 13.940 17.590 ;
        RECT 13.770 17.060 13.940 17.230 ;
        RECT 14.250 17.780 14.420 17.950 ;
        RECT 14.250 17.420 14.420 17.590 ;
        RECT 14.250 17.060 14.420 17.230 ;
        RECT 14.730 17.780 14.900 17.950 ;
        RECT 14.730 17.420 14.900 17.590 ;
        RECT 14.730 17.060 14.900 17.230 ;
        RECT 15.210 17.780 15.380 17.950 ;
        RECT 15.210 17.420 15.380 17.590 ;
        RECT 15.210 17.060 15.380 17.230 ;
        RECT 15.690 17.780 15.860 17.950 ;
        RECT 15.690 17.420 15.860 17.590 ;
        RECT 15.690 17.060 15.860 17.230 ;
        RECT 16.170 17.780 16.340 17.950 ;
        RECT 16.170 17.420 16.340 17.590 ;
        RECT 16.170 17.060 16.340 17.230 ;
        RECT 16.650 17.780 16.820 17.950 ;
        RECT 16.650 17.420 16.820 17.590 ;
        RECT 16.650 17.060 16.820 17.230 ;
        RECT 17.130 17.780 17.300 17.950 ;
        RECT 17.130 17.420 17.300 17.590 ;
        RECT 17.130 17.060 17.300 17.230 ;
        RECT 20.415 17.780 20.585 17.950 ;
        RECT 20.415 17.420 20.585 17.590 ;
        RECT 20.415 17.060 20.585 17.230 ;
        RECT 21.375 17.780 21.545 17.950 ;
        RECT 21.375 17.420 21.545 17.590 ;
        RECT 21.375 17.060 21.545 17.230 ;
        RECT 22.335 17.780 22.505 17.950 ;
        RECT 22.335 17.420 22.505 17.590 ;
        RECT 22.335 17.060 22.505 17.230 ;
        RECT 23.295 17.780 23.465 17.950 ;
        RECT 23.295 17.420 23.465 17.590 ;
        RECT 23.295 17.060 23.465 17.230 ;
        RECT 24.255 17.780 24.425 17.950 ;
        RECT 24.255 17.420 24.425 17.590 ;
        RECT 24.255 17.060 24.425 17.230 ;
        RECT 26.740 15.700 26.910 15.870 ;
        RECT 1.565 14.920 1.735 15.090 ;
        RECT 2.525 14.920 2.695 15.090 ;
        RECT 3.485 14.920 3.655 15.090 ;
        RECT 4.445 14.920 4.615 15.090 ;
        RECT 5.405 14.920 5.575 15.090 ;
        RECT 6.365 14.920 6.535 15.090 ;
        RECT 12.330 14.940 12.500 15.110 ;
        RECT 12.810 14.940 12.980 15.110 ;
        RECT 13.290 14.940 13.460 15.110 ;
        RECT 13.770 14.940 13.940 15.110 ;
        RECT 14.250 14.940 14.420 15.110 ;
        RECT 14.730 14.940 14.900 15.110 ;
        RECT 15.210 14.940 15.380 15.110 ;
        RECT 15.690 14.940 15.860 15.110 ;
        RECT 16.170 14.940 16.340 15.110 ;
        RECT 16.650 14.940 16.820 15.110 ;
        RECT 17.130 14.940 17.300 15.110 ;
        RECT 18.675 14.865 18.845 15.245 ;
        RECT 20.415 14.940 20.585 15.110 ;
        RECT 21.375 14.940 21.545 15.110 ;
        RECT 22.335 14.940 22.505 15.110 ;
        RECT 23.295 14.940 23.465 15.110 ;
        RECT 24.255 14.940 24.425 15.110 ;
        RECT 12.330 14.385 12.500 14.555 ;
        RECT 13.290 14.385 13.460 14.555 ;
        RECT 14.250 14.385 14.420 14.555 ;
        RECT 15.210 14.385 15.380 14.555 ;
        RECT 16.170 14.385 16.340 14.555 ;
        RECT 17.130 14.385 17.300 14.555 ;
        RECT 19.935 14.385 20.105 14.555 ;
        RECT 20.895 14.385 21.065 14.555 ;
        RECT 21.855 14.385 22.025 14.555 ;
        RECT 22.815 14.385 22.985 14.555 ;
        RECT 23.775 14.385 23.945 14.555 ;
        RECT 24.735 14.385 24.905 14.555 ;
        RECT 1.565 11.325 1.735 11.495 ;
        RECT 1.565 10.965 1.735 11.135 ;
        RECT 1.565 10.605 1.735 10.775 ;
        RECT 2.525 11.325 2.695 11.495 ;
        RECT 2.525 10.965 2.695 11.135 ;
        RECT 2.525 10.605 2.695 10.775 ;
        RECT 3.485 11.325 3.655 11.495 ;
        RECT 3.485 10.965 3.655 11.135 ;
        RECT 3.485 10.605 3.655 10.775 ;
        RECT 4.445 11.325 4.615 11.495 ;
        RECT 4.445 10.965 4.615 11.135 ;
        RECT 4.445 10.605 4.615 10.775 ;
        RECT 5.405 11.325 5.575 11.495 ;
        RECT 5.405 10.965 5.575 11.135 ;
        RECT 5.405 10.605 5.575 10.775 ;
        RECT 6.365 11.325 6.535 11.495 ;
        RECT 6.365 10.965 6.535 11.135 ;
        RECT 6.365 10.605 6.535 10.775 ;
        RECT 12.330 11.345 12.500 11.515 ;
        RECT 12.330 10.985 12.500 11.155 ;
        RECT 12.330 10.625 12.500 10.795 ;
        RECT 12.810 11.345 12.980 11.515 ;
        RECT 12.810 10.985 12.980 11.155 ;
        RECT 12.810 10.625 12.980 10.795 ;
        RECT 13.290 11.345 13.460 11.515 ;
        RECT 13.290 10.985 13.460 11.155 ;
        RECT 13.290 10.625 13.460 10.795 ;
        RECT 13.770 11.345 13.940 11.515 ;
        RECT 13.770 10.985 13.940 11.155 ;
        RECT 13.770 10.625 13.940 10.795 ;
        RECT 14.250 11.345 14.420 11.515 ;
        RECT 14.250 10.985 14.420 11.155 ;
        RECT 14.250 10.625 14.420 10.795 ;
        RECT 14.730 11.345 14.900 11.515 ;
        RECT 14.730 10.985 14.900 11.155 ;
        RECT 14.730 10.625 14.900 10.795 ;
        RECT 15.210 11.345 15.380 11.515 ;
        RECT 15.210 10.985 15.380 11.155 ;
        RECT 15.210 10.625 15.380 10.795 ;
        RECT 15.690 11.345 15.860 11.515 ;
        RECT 15.690 10.985 15.860 11.155 ;
        RECT 15.690 10.625 15.860 10.795 ;
        RECT 16.170 11.345 16.340 11.515 ;
        RECT 16.170 10.985 16.340 11.155 ;
        RECT 16.170 10.625 16.340 10.795 ;
        RECT 16.650 11.345 16.820 11.515 ;
        RECT 16.650 10.985 16.820 11.155 ;
        RECT 16.650 10.625 16.820 10.795 ;
        RECT 17.130 11.345 17.300 11.515 ;
        RECT 17.130 10.985 17.300 11.155 ;
        RECT 17.130 10.625 17.300 10.795 ;
        RECT 20.415 11.345 20.585 11.515 ;
        RECT 20.415 10.985 20.585 11.155 ;
        RECT 20.415 10.625 20.585 10.795 ;
        RECT 21.375 11.345 21.545 11.515 ;
        RECT 21.375 10.985 21.545 11.155 ;
        RECT 21.375 10.625 21.545 10.795 ;
        RECT 22.335 11.345 22.505 11.515 ;
        RECT 22.335 10.985 22.505 11.155 ;
        RECT 22.335 10.625 22.505 10.795 ;
        RECT 23.295 11.345 23.465 11.515 ;
        RECT 23.295 10.985 23.465 11.155 ;
        RECT 23.295 10.625 23.465 10.795 ;
        RECT 24.255 11.345 24.425 11.515 ;
        RECT 24.255 10.985 24.425 11.155 ;
        RECT 24.255 10.625 24.425 10.795 ;
        RECT 26.740 9.265 26.910 9.435 ;
        RECT 1.565 8.485 1.735 8.655 ;
        RECT 2.525 8.485 2.695 8.655 ;
        RECT 3.485 8.485 3.655 8.655 ;
        RECT 4.445 8.485 4.615 8.655 ;
        RECT 5.405 8.485 5.575 8.655 ;
        RECT 6.365 8.485 6.535 8.655 ;
        RECT 12.330 8.505 12.500 8.675 ;
        RECT 12.810 8.505 12.980 8.675 ;
        RECT 13.290 8.505 13.460 8.675 ;
        RECT 13.770 8.505 13.940 8.675 ;
        RECT 14.250 8.505 14.420 8.675 ;
        RECT 14.730 8.505 14.900 8.675 ;
        RECT 15.210 8.505 15.380 8.675 ;
        RECT 15.690 8.505 15.860 8.675 ;
        RECT 16.170 8.505 16.340 8.675 ;
        RECT 16.650 8.505 16.820 8.675 ;
        RECT 17.130 8.505 17.300 8.675 ;
        RECT 18.675 8.430 18.845 8.810 ;
        RECT 20.415 8.505 20.585 8.675 ;
        RECT 21.375 8.505 21.545 8.675 ;
        RECT 22.335 8.505 22.505 8.675 ;
        RECT 23.295 8.505 23.465 8.675 ;
        RECT 24.255 8.505 24.425 8.675 ;
        RECT 12.330 7.950 12.500 8.120 ;
        RECT 13.290 7.950 13.460 8.120 ;
        RECT 14.250 7.950 14.420 8.120 ;
        RECT 15.210 7.950 15.380 8.120 ;
        RECT 16.170 7.950 16.340 8.120 ;
        RECT 17.130 7.950 17.300 8.120 ;
        RECT 19.935 7.950 20.105 8.120 ;
        RECT 20.895 7.950 21.065 8.120 ;
        RECT 21.855 7.950 22.025 8.120 ;
        RECT 22.815 7.950 22.985 8.120 ;
        RECT 23.775 7.950 23.945 8.120 ;
        RECT 24.735 7.950 24.905 8.120 ;
        RECT 1.565 4.890 1.735 5.060 ;
        RECT 1.565 4.530 1.735 4.700 ;
        RECT 1.565 4.170 1.735 4.340 ;
        RECT 2.525 4.890 2.695 5.060 ;
        RECT 2.525 4.530 2.695 4.700 ;
        RECT 2.525 4.170 2.695 4.340 ;
        RECT 3.485 4.890 3.655 5.060 ;
        RECT 3.485 4.530 3.655 4.700 ;
        RECT 3.485 4.170 3.655 4.340 ;
        RECT 4.445 4.890 4.615 5.060 ;
        RECT 4.445 4.530 4.615 4.700 ;
        RECT 4.445 4.170 4.615 4.340 ;
        RECT 5.405 4.890 5.575 5.060 ;
        RECT 5.405 4.530 5.575 4.700 ;
        RECT 5.405 4.170 5.575 4.340 ;
        RECT 6.365 4.890 6.535 5.060 ;
        RECT 6.365 4.530 6.535 4.700 ;
        RECT 6.365 4.170 6.535 4.340 ;
        RECT 12.330 4.910 12.500 5.080 ;
        RECT 12.330 4.550 12.500 4.720 ;
        RECT 12.330 4.190 12.500 4.360 ;
        RECT 12.810 4.910 12.980 5.080 ;
        RECT 12.810 4.550 12.980 4.720 ;
        RECT 12.810 4.190 12.980 4.360 ;
        RECT 13.290 4.910 13.460 5.080 ;
        RECT 13.290 4.550 13.460 4.720 ;
        RECT 13.290 4.190 13.460 4.360 ;
        RECT 13.770 4.910 13.940 5.080 ;
        RECT 13.770 4.550 13.940 4.720 ;
        RECT 13.770 4.190 13.940 4.360 ;
        RECT 14.250 4.910 14.420 5.080 ;
        RECT 14.250 4.550 14.420 4.720 ;
        RECT 14.250 4.190 14.420 4.360 ;
        RECT 14.730 4.910 14.900 5.080 ;
        RECT 14.730 4.550 14.900 4.720 ;
        RECT 14.730 4.190 14.900 4.360 ;
        RECT 15.210 4.910 15.380 5.080 ;
        RECT 15.210 4.550 15.380 4.720 ;
        RECT 15.210 4.190 15.380 4.360 ;
        RECT 15.690 4.910 15.860 5.080 ;
        RECT 15.690 4.550 15.860 4.720 ;
        RECT 15.690 4.190 15.860 4.360 ;
        RECT 16.170 4.910 16.340 5.080 ;
        RECT 16.170 4.550 16.340 4.720 ;
        RECT 16.170 4.190 16.340 4.360 ;
        RECT 16.650 4.910 16.820 5.080 ;
        RECT 16.650 4.550 16.820 4.720 ;
        RECT 16.650 4.190 16.820 4.360 ;
        RECT 17.130 4.910 17.300 5.080 ;
        RECT 17.130 4.550 17.300 4.720 ;
        RECT 17.130 4.190 17.300 4.360 ;
        RECT 20.415 4.910 20.585 5.080 ;
        RECT 20.415 4.550 20.585 4.720 ;
        RECT 20.415 4.190 20.585 4.360 ;
        RECT 21.375 4.910 21.545 5.080 ;
        RECT 21.375 4.550 21.545 4.720 ;
        RECT 21.375 4.190 21.545 4.360 ;
        RECT 22.335 4.910 22.505 5.080 ;
        RECT 22.335 4.550 22.505 4.720 ;
        RECT 22.335 4.190 22.505 4.360 ;
        RECT 23.295 4.910 23.465 5.080 ;
        RECT 23.295 4.550 23.465 4.720 ;
        RECT 23.295 4.190 23.465 4.360 ;
        RECT 24.255 4.910 24.425 5.080 ;
        RECT 24.255 4.550 24.425 4.720 ;
        RECT 24.255 4.190 24.425 4.360 ;
        RECT 26.740 2.830 26.910 3.000 ;
        RECT 1.565 2.050 1.735 2.220 ;
        RECT 2.525 2.050 2.695 2.220 ;
        RECT 3.485 2.050 3.655 2.220 ;
        RECT 4.445 2.050 4.615 2.220 ;
        RECT 5.405 2.050 5.575 2.220 ;
        RECT 6.365 2.050 6.535 2.220 ;
        RECT 12.330 2.070 12.500 2.240 ;
        RECT 12.810 2.070 12.980 2.240 ;
        RECT 13.290 2.070 13.460 2.240 ;
        RECT 13.770 2.070 13.940 2.240 ;
        RECT 14.250 2.070 14.420 2.240 ;
        RECT 14.730 2.070 14.900 2.240 ;
        RECT 15.210 2.070 15.380 2.240 ;
        RECT 15.690 2.070 15.860 2.240 ;
        RECT 16.170 2.070 16.340 2.240 ;
        RECT 16.650 2.070 16.820 2.240 ;
        RECT 17.130 2.070 17.300 2.240 ;
        RECT 18.675 1.995 18.845 2.375 ;
        RECT 20.415 2.070 20.585 2.240 ;
        RECT 21.375 2.070 21.545 2.240 ;
        RECT 22.335 2.070 22.505 2.240 ;
        RECT 23.295 2.070 23.465 2.240 ;
        RECT 24.255 2.070 24.425 2.240 ;
        RECT 12.330 1.515 12.500 1.685 ;
        RECT 13.290 1.515 13.460 1.685 ;
        RECT 14.250 1.515 14.420 1.685 ;
        RECT 15.210 1.515 15.380 1.685 ;
        RECT 16.170 1.515 16.340 1.685 ;
        RECT 17.130 1.515 17.300 1.685 ;
        RECT 19.935 1.515 20.105 1.685 ;
        RECT 20.895 1.515 21.065 1.685 ;
        RECT 21.855 1.515 22.025 1.685 ;
        RECT 22.815 1.515 22.985 1.685 ;
        RECT 23.775 1.515 23.945 1.685 ;
        RECT 24.735 1.515 24.905 1.685 ;
      LAYER met1 ;
        RECT 11.410 205.550 16.820 205.720 ;
        RECT 1.535 203.420 1.765 204.780 ;
        RECT 2.495 203.420 2.725 204.780 ;
        RECT 3.455 203.420 3.685 204.780 ;
        RECT 4.415 203.420 4.645 204.780 ;
        RECT 5.375 203.420 5.605 204.780 ;
        RECT 6.335 203.420 6.565 204.780 ;
        RECT 1.565 202.715 1.735 203.420 ;
        RECT 2.525 202.715 2.695 203.420 ;
        RECT 3.485 202.715 3.655 203.420 ;
        RECT 4.445 202.715 4.615 203.420 ;
        RECT 5.405 202.715 5.575 203.420 ;
        RECT 6.365 202.715 6.535 203.420 ;
        RECT 11.410 202.735 11.580 205.550 ;
        RECT 12.810 204.800 12.980 205.550 ;
        RECT 13.770 204.800 13.940 205.550 ;
        RECT 14.730 204.800 14.900 205.550 ;
        RECT 15.690 204.800 15.860 205.550 ;
        RECT 16.650 204.800 16.820 205.550 ;
        RECT 19.015 205.550 24.425 205.720 ;
        RECT 12.300 203.440 12.530 204.800 ;
        RECT 12.780 203.440 13.010 204.800 ;
        RECT 13.260 203.440 13.490 204.800 ;
        RECT 13.740 203.440 13.970 204.800 ;
        RECT 14.220 203.440 14.450 204.800 ;
        RECT 14.700 203.440 14.930 204.800 ;
        RECT 15.180 203.440 15.410 204.800 ;
        RECT 15.660 203.440 15.890 204.800 ;
        RECT 16.140 203.440 16.370 204.800 ;
        RECT 16.620 203.440 16.850 204.800 ;
        RECT 17.100 203.440 17.330 204.800 ;
        RECT 10.505 202.715 11.580 202.735 ;
        RECT 1.565 202.565 11.580 202.715 ;
        RECT 1.565 202.545 10.705 202.565 ;
        RECT 1.565 201.880 1.735 202.545 ;
        RECT 2.525 201.880 2.695 202.545 ;
        RECT 3.485 201.880 3.655 202.545 ;
        RECT 4.445 201.880 4.615 202.545 ;
        RECT 5.405 201.880 5.575 202.545 ;
        RECT 6.365 201.880 6.535 202.545 ;
        RECT 1.535 201.360 1.765 201.880 ;
        RECT 2.495 201.360 2.725 201.880 ;
        RECT 3.455 201.360 3.685 201.880 ;
        RECT 4.415 201.360 4.645 201.880 ;
        RECT 5.375 201.360 5.605 201.880 ;
        RECT 6.335 201.360 6.565 201.880 ;
        RECT 11.410 200.680 11.580 202.565 ;
        RECT 12.330 202.735 12.500 203.440 ;
        RECT 13.290 202.735 13.460 203.440 ;
        RECT 14.250 202.735 14.420 203.440 ;
        RECT 15.210 202.735 15.380 203.440 ;
        RECT 16.170 202.735 16.340 203.440 ;
        RECT 17.130 202.735 17.300 203.440 ;
        RECT 19.015 202.735 19.185 205.550 ;
        RECT 20.415 204.800 20.585 205.550 ;
        RECT 21.375 204.800 21.545 205.550 ;
        RECT 22.335 204.800 22.505 205.550 ;
        RECT 23.295 204.800 23.465 205.550 ;
        RECT 24.255 204.800 24.425 205.550 ;
        RECT 20.385 203.440 20.615 204.800 ;
        RECT 21.345 203.440 21.575 204.800 ;
        RECT 22.305 203.440 22.535 204.800 ;
        RECT 23.265 203.440 23.495 204.800 ;
        RECT 24.225 203.440 24.455 204.800 ;
        RECT 12.330 202.565 19.185 202.735 ;
        RECT 12.330 201.900 12.500 202.565 ;
        RECT 13.290 201.900 13.460 202.565 ;
        RECT 14.250 201.900 14.420 202.565 ;
        RECT 15.210 201.900 15.380 202.565 ;
        RECT 16.170 201.900 16.340 202.565 ;
        RECT 17.130 201.900 17.300 202.565 ;
        RECT 19.015 201.925 19.185 202.565 ;
        RECT 26.630 202.270 27.000 202.540 ;
        RECT 18.670 201.920 19.185 201.925 ;
        RECT 12.300 201.380 12.530 201.900 ;
        RECT 12.780 201.380 13.010 201.900 ;
        RECT 13.260 201.380 13.490 201.900 ;
        RECT 13.740 201.380 13.970 201.900 ;
        RECT 14.220 201.380 14.450 201.900 ;
        RECT 14.700 201.380 14.930 201.900 ;
        RECT 15.180 201.380 15.410 201.900 ;
        RECT 15.660 201.380 15.890 201.900 ;
        RECT 16.140 201.380 16.370 201.900 ;
        RECT 16.620 201.380 16.850 201.900 ;
        RECT 17.100 201.380 17.330 201.900 ;
        RECT 18.645 201.425 19.185 201.920 ;
        RECT 18.645 201.420 18.875 201.425 ;
        RECT 12.250 201.225 12.580 201.240 ;
        RECT 12.235 200.965 12.595 201.225 ;
        RECT 12.250 200.940 12.580 200.965 ;
        RECT 12.810 200.680 12.980 201.380 ;
        RECT 13.210 201.225 13.540 201.240 ;
        RECT 13.190 200.965 13.550 201.225 ;
        RECT 13.210 200.940 13.540 200.965 ;
        RECT 13.770 200.680 13.940 201.380 ;
        RECT 14.170 201.225 14.500 201.240 ;
        RECT 14.150 200.965 14.510 201.225 ;
        RECT 14.170 200.940 14.500 200.965 ;
        RECT 14.730 200.680 14.900 201.380 ;
        RECT 15.130 201.225 15.460 201.240 ;
        RECT 15.110 200.965 15.470 201.225 ;
        RECT 15.130 200.940 15.460 200.965 ;
        RECT 15.690 200.680 15.860 201.380 ;
        RECT 16.090 201.220 16.420 201.240 ;
        RECT 16.075 200.960 16.435 201.220 ;
        RECT 16.090 200.940 16.420 200.960 ;
        RECT 16.650 200.680 16.820 201.380 ;
        RECT 17.050 201.220 17.380 201.240 ;
        RECT 17.035 200.960 17.395 201.220 ;
        RECT 17.050 200.940 17.380 200.960 ;
        RECT 11.410 200.510 16.820 200.680 ;
        RECT 19.015 200.680 19.185 201.425 ;
        RECT 20.385 201.380 20.615 201.900 ;
        RECT 21.345 201.380 21.575 201.900 ;
        RECT 22.305 201.380 22.535 201.900 ;
        RECT 23.265 201.380 23.495 201.900 ;
        RECT 24.225 201.380 24.455 201.900 ;
        RECT 19.855 201.225 20.185 201.240 ;
        RECT 19.840 200.965 20.200 201.225 ;
        RECT 19.855 200.940 20.185 200.965 ;
        RECT 20.415 200.680 20.585 201.380 ;
        RECT 20.815 201.225 21.145 201.240 ;
        RECT 20.795 200.965 21.155 201.225 ;
        RECT 20.815 200.940 21.145 200.965 ;
        RECT 21.375 200.680 21.545 201.380 ;
        RECT 21.775 201.225 22.105 201.240 ;
        RECT 21.755 200.965 22.115 201.225 ;
        RECT 21.775 200.940 22.105 200.965 ;
        RECT 22.335 200.680 22.505 201.380 ;
        RECT 22.735 201.225 23.065 201.240 ;
        RECT 22.715 200.965 23.075 201.225 ;
        RECT 22.735 200.940 23.065 200.965 ;
        RECT 23.295 200.680 23.465 201.380 ;
        RECT 23.695 201.220 24.025 201.240 ;
        RECT 23.680 200.960 24.040 201.220 ;
        RECT 23.695 200.940 24.025 200.960 ;
        RECT 24.255 200.680 24.425 201.380 ;
        RECT 24.655 201.220 24.985 201.240 ;
        RECT 24.640 200.960 25.000 201.220 ;
        RECT 24.655 200.940 24.985 200.960 ;
        RECT 19.015 200.510 24.425 200.680 ;
        RECT 11.410 199.115 16.820 199.285 ;
        RECT 1.535 196.985 1.765 198.345 ;
        RECT 2.495 196.985 2.725 198.345 ;
        RECT 3.455 196.985 3.685 198.345 ;
        RECT 4.415 196.985 4.645 198.345 ;
        RECT 5.375 196.985 5.605 198.345 ;
        RECT 6.335 196.985 6.565 198.345 ;
        RECT 1.565 196.280 1.735 196.985 ;
        RECT 2.525 196.280 2.695 196.985 ;
        RECT 3.485 196.280 3.655 196.985 ;
        RECT 4.445 196.280 4.615 196.985 ;
        RECT 5.405 196.280 5.575 196.985 ;
        RECT 6.365 196.280 6.535 196.985 ;
        RECT 11.410 196.300 11.580 199.115 ;
        RECT 12.810 198.365 12.980 199.115 ;
        RECT 13.770 198.365 13.940 199.115 ;
        RECT 14.730 198.365 14.900 199.115 ;
        RECT 15.690 198.365 15.860 199.115 ;
        RECT 16.650 198.365 16.820 199.115 ;
        RECT 19.015 199.115 24.425 199.285 ;
        RECT 12.300 197.005 12.530 198.365 ;
        RECT 12.780 197.005 13.010 198.365 ;
        RECT 13.260 197.005 13.490 198.365 ;
        RECT 13.740 197.005 13.970 198.365 ;
        RECT 14.220 197.005 14.450 198.365 ;
        RECT 14.700 197.005 14.930 198.365 ;
        RECT 15.180 197.005 15.410 198.365 ;
        RECT 15.660 197.005 15.890 198.365 ;
        RECT 16.140 197.005 16.370 198.365 ;
        RECT 16.620 197.005 16.850 198.365 ;
        RECT 17.100 197.005 17.330 198.365 ;
        RECT 10.505 196.280 11.580 196.300 ;
        RECT 1.565 196.130 11.580 196.280 ;
        RECT 1.565 196.110 10.705 196.130 ;
        RECT 1.565 195.445 1.735 196.110 ;
        RECT 2.525 195.445 2.695 196.110 ;
        RECT 3.485 195.445 3.655 196.110 ;
        RECT 4.445 195.445 4.615 196.110 ;
        RECT 5.405 195.445 5.575 196.110 ;
        RECT 6.365 195.445 6.535 196.110 ;
        RECT 1.535 194.925 1.765 195.445 ;
        RECT 2.495 194.925 2.725 195.445 ;
        RECT 3.455 194.925 3.685 195.445 ;
        RECT 4.415 194.925 4.645 195.445 ;
        RECT 5.375 194.925 5.605 195.445 ;
        RECT 6.335 194.925 6.565 195.445 ;
        RECT 11.410 194.245 11.580 196.130 ;
        RECT 12.330 196.300 12.500 197.005 ;
        RECT 13.290 196.300 13.460 197.005 ;
        RECT 14.250 196.300 14.420 197.005 ;
        RECT 15.210 196.300 15.380 197.005 ;
        RECT 16.170 196.300 16.340 197.005 ;
        RECT 17.130 196.300 17.300 197.005 ;
        RECT 19.015 196.300 19.185 199.115 ;
        RECT 20.415 198.365 20.585 199.115 ;
        RECT 21.375 198.365 21.545 199.115 ;
        RECT 22.335 198.365 22.505 199.115 ;
        RECT 23.295 198.365 23.465 199.115 ;
        RECT 24.255 198.365 24.425 199.115 ;
        RECT 20.385 197.005 20.615 198.365 ;
        RECT 21.345 197.005 21.575 198.365 ;
        RECT 22.305 197.005 22.535 198.365 ;
        RECT 23.265 197.005 23.495 198.365 ;
        RECT 24.225 197.005 24.455 198.365 ;
        RECT 12.330 196.130 19.185 196.300 ;
        RECT 12.330 195.465 12.500 196.130 ;
        RECT 13.290 195.465 13.460 196.130 ;
        RECT 14.250 195.465 14.420 196.130 ;
        RECT 15.210 195.465 15.380 196.130 ;
        RECT 16.170 195.465 16.340 196.130 ;
        RECT 17.130 195.465 17.300 196.130 ;
        RECT 19.015 195.490 19.185 196.130 ;
        RECT 26.630 195.835 27.000 196.105 ;
        RECT 18.670 195.485 19.185 195.490 ;
        RECT 12.300 194.945 12.530 195.465 ;
        RECT 12.780 194.945 13.010 195.465 ;
        RECT 13.260 194.945 13.490 195.465 ;
        RECT 13.740 194.945 13.970 195.465 ;
        RECT 14.220 194.945 14.450 195.465 ;
        RECT 14.700 194.945 14.930 195.465 ;
        RECT 15.180 194.945 15.410 195.465 ;
        RECT 15.660 194.945 15.890 195.465 ;
        RECT 16.140 194.945 16.370 195.465 ;
        RECT 16.620 194.945 16.850 195.465 ;
        RECT 17.100 194.945 17.330 195.465 ;
        RECT 18.645 194.990 19.185 195.485 ;
        RECT 18.645 194.985 18.875 194.990 ;
        RECT 12.250 194.790 12.580 194.805 ;
        RECT 12.235 194.530 12.595 194.790 ;
        RECT 12.250 194.505 12.580 194.530 ;
        RECT 12.810 194.245 12.980 194.945 ;
        RECT 13.210 194.790 13.540 194.805 ;
        RECT 13.190 194.530 13.550 194.790 ;
        RECT 13.210 194.505 13.540 194.530 ;
        RECT 13.770 194.245 13.940 194.945 ;
        RECT 14.170 194.790 14.500 194.805 ;
        RECT 14.150 194.530 14.510 194.790 ;
        RECT 14.170 194.505 14.500 194.530 ;
        RECT 14.730 194.245 14.900 194.945 ;
        RECT 15.130 194.790 15.460 194.805 ;
        RECT 15.110 194.530 15.470 194.790 ;
        RECT 15.130 194.505 15.460 194.530 ;
        RECT 15.690 194.245 15.860 194.945 ;
        RECT 16.090 194.785 16.420 194.805 ;
        RECT 16.075 194.525 16.435 194.785 ;
        RECT 16.090 194.505 16.420 194.525 ;
        RECT 16.650 194.245 16.820 194.945 ;
        RECT 17.050 194.785 17.380 194.805 ;
        RECT 17.035 194.525 17.395 194.785 ;
        RECT 17.050 194.505 17.380 194.525 ;
        RECT 11.410 194.075 16.820 194.245 ;
        RECT 19.015 194.245 19.185 194.990 ;
        RECT 20.385 194.945 20.615 195.465 ;
        RECT 21.345 194.945 21.575 195.465 ;
        RECT 22.305 194.945 22.535 195.465 ;
        RECT 23.265 194.945 23.495 195.465 ;
        RECT 24.225 194.945 24.455 195.465 ;
        RECT 19.855 194.790 20.185 194.805 ;
        RECT 19.840 194.530 20.200 194.790 ;
        RECT 19.855 194.505 20.185 194.530 ;
        RECT 20.415 194.245 20.585 194.945 ;
        RECT 20.815 194.790 21.145 194.805 ;
        RECT 20.795 194.530 21.155 194.790 ;
        RECT 20.815 194.505 21.145 194.530 ;
        RECT 21.375 194.245 21.545 194.945 ;
        RECT 21.775 194.790 22.105 194.805 ;
        RECT 21.755 194.530 22.115 194.790 ;
        RECT 21.775 194.505 22.105 194.530 ;
        RECT 22.335 194.245 22.505 194.945 ;
        RECT 22.735 194.790 23.065 194.805 ;
        RECT 22.715 194.530 23.075 194.790 ;
        RECT 22.735 194.505 23.065 194.530 ;
        RECT 23.295 194.245 23.465 194.945 ;
        RECT 23.695 194.785 24.025 194.805 ;
        RECT 23.680 194.525 24.040 194.785 ;
        RECT 23.695 194.505 24.025 194.525 ;
        RECT 24.255 194.245 24.425 194.945 ;
        RECT 24.655 194.785 24.985 194.805 ;
        RECT 24.640 194.525 25.000 194.785 ;
        RECT 24.655 194.505 24.985 194.525 ;
        RECT 19.015 194.075 24.425 194.245 ;
        RECT 11.410 192.680 16.820 192.850 ;
        RECT 1.535 190.550 1.765 191.910 ;
        RECT 2.495 190.550 2.725 191.910 ;
        RECT 3.455 190.550 3.685 191.910 ;
        RECT 4.415 190.550 4.645 191.910 ;
        RECT 5.375 190.550 5.605 191.910 ;
        RECT 6.335 190.550 6.565 191.910 ;
        RECT 1.565 189.845 1.735 190.550 ;
        RECT 2.525 189.845 2.695 190.550 ;
        RECT 3.485 189.845 3.655 190.550 ;
        RECT 4.445 189.845 4.615 190.550 ;
        RECT 5.405 189.845 5.575 190.550 ;
        RECT 6.365 189.845 6.535 190.550 ;
        RECT 11.410 189.865 11.580 192.680 ;
        RECT 12.810 191.930 12.980 192.680 ;
        RECT 13.770 191.930 13.940 192.680 ;
        RECT 14.730 191.930 14.900 192.680 ;
        RECT 15.690 191.930 15.860 192.680 ;
        RECT 16.650 191.930 16.820 192.680 ;
        RECT 19.015 192.680 24.425 192.850 ;
        RECT 12.300 190.570 12.530 191.930 ;
        RECT 12.780 190.570 13.010 191.930 ;
        RECT 13.260 190.570 13.490 191.930 ;
        RECT 13.740 190.570 13.970 191.930 ;
        RECT 14.220 190.570 14.450 191.930 ;
        RECT 14.700 190.570 14.930 191.930 ;
        RECT 15.180 190.570 15.410 191.930 ;
        RECT 15.660 190.570 15.890 191.930 ;
        RECT 16.140 190.570 16.370 191.930 ;
        RECT 16.620 190.570 16.850 191.930 ;
        RECT 17.100 190.570 17.330 191.930 ;
        RECT 10.505 189.845 11.580 189.865 ;
        RECT 1.565 189.695 11.580 189.845 ;
        RECT 1.565 189.675 10.705 189.695 ;
        RECT 1.565 189.010 1.735 189.675 ;
        RECT 2.525 189.010 2.695 189.675 ;
        RECT 3.485 189.010 3.655 189.675 ;
        RECT 4.445 189.010 4.615 189.675 ;
        RECT 5.405 189.010 5.575 189.675 ;
        RECT 6.365 189.010 6.535 189.675 ;
        RECT 1.535 188.490 1.765 189.010 ;
        RECT 2.495 188.490 2.725 189.010 ;
        RECT 3.455 188.490 3.685 189.010 ;
        RECT 4.415 188.490 4.645 189.010 ;
        RECT 5.375 188.490 5.605 189.010 ;
        RECT 6.335 188.490 6.565 189.010 ;
        RECT 11.410 187.810 11.580 189.695 ;
        RECT 12.330 189.865 12.500 190.570 ;
        RECT 13.290 189.865 13.460 190.570 ;
        RECT 14.250 189.865 14.420 190.570 ;
        RECT 15.210 189.865 15.380 190.570 ;
        RECT 16.170 189.865 16.340 190.570 ;
        RECT 17.130 189.865 17.300 190.570 ;
        RECT 19.015 189.865 19.185 192.680 ;
        RECT 20.415 191.930 20.585 192.680 ;
        RECT 21.375 191.930 21.545 192.680 ;
        RECT 22.335 191.930 22.505 192.680 ;
        RECT 23.295 191.930 23.465 192.680 ;
        RECT 24.255 191.930 24.425 192.680 ;
        RECT 20.385 190.570 20.615 191.930 ;
        RECT 21.345 190.570 21.575 191.930 ;
        RECT 22.305 190.570 22.535 191.930 ;
        RECT 23.265 190.570 23.495 191.930 ;
        RECT 24.225 190.570 24.455 191.930 ;
        RECT 12.330 189.695 19.185 189.865 ;
        RECT 12.330 189.030 12.500 189.695 ;
        RECT 13.290 189.030 13.460 189.695 ;
        RECT 14.250 189.030 14.420 189.695 ;
        RECT 15.210 189.030 15.380 189.695 ;
        RECT 16.170 189.030 16.340 189.695 ;
        RECT 17.130 189.030 17.300 189.695 ;
        RECT 19.015 189.055 19.185 189.695 ;
        RECT 26.630 189.400 27.000 189.670 ;
        RECT 18.670 189.050 19.185 189.055 ;
        RECT 12.300 188.510 12.530 189.030 ;
        RECT 12.780 188.510 13.010 189.030 ;
        RECT 13.260 188.510 13.490 189.030 ;
        RECT 13.740 188.510 13.970 189.030 ;
        RECT 14.220 188.510 14.450 189.030 ;
        RECT 14.700 188.510 14.930 189.030 ;
        RECT 15.180 188.510 15.410 189.030 ;
        RECT 15.660 188.510 15.890 189.030 ;
        RECT 16.140 188.510 16.370 189.030 ;
        RECT 16.620 188.510 16.850 189.030 ;
        RECT 17.100 188.510 17.330 189.030 ;
        RECT 18.645 188.555 19.185 189.050 ;
        RECT 18.645 188.550 18.875 188.555 ;
        RECT 12.250 188.355 12.580 188.370 ;
        RECT 12.235 188.095 12.595 188.355 ;
        RECT 12.250 188.070 12.580 188.095 ;
        RECT 12.810 187.810 12.980 188.510 ;
        RECT 13.210 188.355 13.540 188.370 ;
        RECT 13.190 188.095 13.550 188.355 ;
        RECT 13.210 188.070 13.540 188.095 ;
        RECT 13.770 187.810 13.940 188.510 ;
        RECT 14.170 188.355 14.500 188.370 ;
        RECT 14.150 188.095 14.510 188.355 ;
        RECT 14.170 188.070 14.500 188.095 ;
        RECT 14.730 187.810 14.900 188.510 ;
        RECT 15.130 188.355 15.460 188.370 ;
        RECT 15.110 188.095 15.470 188.355 ;
        RECT 15.130 188.070 15.460 188.095 ;
        RECT 15.690 187.810 15.860 188.510 ;
        RECT 16.090 188.350 16.420 188.370 ;
        RECT 16.075 188.090 16.435 188.350 ;
        RECT 16.090 188.070 16.420 188.090 ;
        RECT 16.650 187.810 16.820 188.510 ;
        RECT 17.050 188.350 17.380 188.370 ;
        RECT 17.035 188.090 17.395 188.350 ;
        RECT 17.050 188.070 17.380 188.090 ;
        RECT 11.410 187.640 16.820 187.810 ;
        RECT 19.015 187.810 19.185 188.555 ;
        RECT 20.385 188.510 20.615 189.030 ;
        RECT 21.345 188.510 21.575 189.030 ;
        RECT 22.305 188.510 22.535 189.030 ;
        RECT 23.265 188.510 23.495 189.030 ;
        RECT 24.225 188.510 24.455 189.030 ;
        RECT 19.855 188.355 20.185 188.370 ;
        RECT 19.840 188.095 20.200 188.355 ;
        RECT 19.855 188.070 20.185 188.095 ;
        RECT 20.415 187.810 20.585 188.510 ;
        RECT 20.815 188.355 21.145 188.370 ;
        RECT 20.795 188.095 21.155 188.355 ;
        RECT 20.815 188.070 21.145 188.095 ;
        RECT 21.375 187.810 21.545 188.510 ;
        RECT 21.775 188.355 22.105 188.370 ;
        RECT 21.755 188.095 22.115 188.355 ;
        RECT 21.775 188.070 22.105 188.095 ;
        RECT 22.335 187.810 22.505 188.510 ;
        RECT 22.735 188.355 23.065 188.370 ;
        RECT 22.715 188.095 23.075 188.355 ;
        RECT 22.735 188.070 23.065 188.095 ;
        RECT 23.295 187.810 23.465 188.510 ;
        RECT 23.695 188.350 24.025 188.370 ;
        RECT 23.680 188.090 24.040 188.350 ;
        RECT 23.695 188.070 24.025 188.090 ;
        RECT 24.255 187.810 24.425 188.510 ;
        RECT 24.655 188.350 24.985 188.370 ;
        RECT 24.640 188.090 25.000 188.350 ;
        RECT 24.655 188.070 24.985 188.090 ;
        RECT 19.015 187.640 24.425 187.810 ;
        RECT 11.410 186.245 16.820 186.415 ;
        RECT 1.535 184.115 1.765 185.475 ;
        RECT 2.495 184.115 2.725 185.475 ;
        RECT 3.455 184.115 3.685 185.475 ;
        RECT 4.415 184.115 4.645 185.475 ;
        RECT 5.375 184.115 5.605 185.475 ;
        RECT 6.335 184.115 6.565 185.475 ;
        RECT 1.565 183.410 1.735 184.115 ;
        RECT 2.525 183.410 2.695 184.115 ;
        RECT 3.485 183.410 3.655 184.115 ;
        RECT 4.445 183.410 4.615 184.115 ;
        RECT 5.405 183.410 5.575 184.115 ;
        RECT 6.365 183.410 6.535 184.115 ;
        RECT 11.410 183.430 11.580 186.245 ;
        RECT 12.810 185.495 12.980 186.245 ;
        RECT 13.770 185.495 13.940 186.245 ;
        RECT 14.730 185.495 14.900 186.245 ;
        RECT 15.690 185.495 15.860 186.245 ;
        RECT 16.650 185.495 16.820 186.245 ;
        RECT 19.015 186.245 24.425 186.415 ;
        RECT 12.300 184.135 12.530 185.495 ;
        RECT 12.780 184.135 13.010 185.495 ;
        RECT 13.260 184.135 13.490 185.495 ;
        RECT 13.740 184.135 13.970 185.495 ;
        RECT 14.220 184.135 14.450 185.495 ;
        RECT 14.700 184.135 14.930 185.495 ;
        RECT 15.180 184.135 15.410 185.495 ;
        RECT 15.660 184.135 15.890 185.495 ;
        RECT 16.140 184.135 16.370 185.495 ;
        RECT 16.620 184.135 16.850 185.495 ;
        RECT 17.100 184.135 17.330 185.495 ;
        RECT 10.505 183.410 11.580 183.430 ;
        RECT 1.565 183.260 11.580 183.410 ;
        RECT 1.565 183.240 10.705 183.260 ;
        RECT 1.565 182.575 1.735 183.240 ;
        RECT 2.525 182.575 2.695 183.240 ;
        RECT 3.485 182.575 3.655 183.240 ;
        RECT 4.445 182.575 4.615 183.240 ;
        RECT 5.405 182.575 5.575 183.240 ;
        RECT 6.365 182.575 6.535 183.240 ;
        RECT 1.535 182.055 1.765 182.575 ;
        RECT 2.495 182.055 2.725 182.575 ;
        RECT 3.455 182.055 3.685 182.575 ;
        RECT 4.415 182.055 4.645 182.575 ;
        RECT 5.375 182.055 5.605 182.575 ;
        RECT 6.335 182.055 6.565 182.575 ;
        RECT 11.410 181.375 11.580 183.260 ;
        RECT 12.330 183.430 12.500 184.135 ;
        RECT 13.290 183.430 13.460 184.135 ;
        RECT 14.250 183.430 14.420 184.135 ;
        RECT 15.210 183.430 15.380 184.135 ;
        RECT 16.170 183.430 16.340 184.135 ;
        RECT 17.130 183.430 17.300 184.135 ;
        RECT 19.015 183.430 19.185 186.245 ;
        RECT 20.415 185.495 20.585 186.245 ;
        RECT 21.375 185.495 21.545 186.245 ;
        RECT 22.335 185.495 22.505 186.245 ;
        RECT 23.295 185.495 23.465 186.245 ;
        RECT 24.255 185.495 24.425 186.245 ;
        RECT 20.385 184.135 20.615 185.495 ;
        RECT 21.345 184.135 21.575 185.495 ;
        RECT 22.305 184.135 22.535 185.495 ;
        RECT 23.265 184.135 23.495 185.495 ;
        RECT 24.225 184.135 24.455 185.495 ;
        RECT 12.330 183.260 19.185 183.430 ;
        RECT 12.330 182.595 12.500 183.260 ;
        RECT 13.290 182.595 13.460 183.260 ;
        RECT 14.250 182.595 14.420 183.260 ;
        RECT 15.210 182.595 15.380 183.260 ;
        RECT 16.170 182.595 16.340 183.260 ;
        RECT 17.130 182.595 17.300 183.260 ;
        RECT 19.015 182.620 19.185 183.260 ;
        RECT 26.630 182.965 27.000 183.235 ;
        RECT 18.670 182.615 19.185 182.620 ;
        RECT 12.300 182.075 12.530 182.595 ;
        RECT 12.780 182.075 13.010 182.595 ;
        RECT 13.260 182.075 13.490 182.595 ;
        RECT 13.740 182.075 13.970 182.595 ;
        RECT 14.220 182.075 14.450 182.595 ;
        RECT 14.700 182.075 14.930 182.595 ;
        RECT 15.180 182.075 15.410 182.595 ;
        RECT 15.660 182.075 15.890 182.595 ;
        RECT 16.140 182.075 16.370 182.595 ;
        RECT 16.620 182.075 16.850 182.595 ;
        RECT 17.100 182.075 17.330 182.595 ;
        RECT 18.645 182.120 19.185 182.615 ;
        RECT 18.645 182.115 18.875 182.120 ;
        RECT 12.250 181.920 12.580 181.935 ;
        RECT 12.235 181.660 12.595 181.920 ;
        RECT 12.250 181.635 12.580 181.660 ;
        RECT 12.810 181.375 12.980 182.075 ;
        RECT 13.210 181.920 13.540 181.935 ;
        RECT 13.190 181.660 13.550 181.920 ;
        RECT 13.210 181.635 13.540 181.660 ;
        RECT 13.770 181.375 13.940 182.075 ;
        RECT 14.170 181.920 14.500 181.935 ;
        RECT 14.150 181.660 14.510 181.920 ;
        RECT 14.170 181.635 14.500 181.660 ;
        RECT 14.730 181.375 14.900 182.075 ;
        RECT 15.130 181.920 15.460 181.935 ;
        RECT 15.110 181.660 15.470 181.920 ;
        RECT 15.130 181.635 15.460 181.660 ;
        RECT 15.690 181.375 15.860 182.075 ;
        RECT 16.090 181.915 16.420 181.935 ;
        RECT 16.075 181.655 16.435 181.915 ;
        RECT 16.090 181.635 16.420 181.655 ;
        RECT 16.650 181.375 16.820 182.075 ;
        RECT 17.050 181.915 17.380 181.935 ;
        RECT 17.035 181.655 17.395 181.915 ;
        RECT 17.050 181.635 17.380 181.655 ;
        RECT 11.410 181.205 16.820 181.375 ;
        RECT 19.015 181.375 19.185 182.120 ;
        RECT 20.385 182.075 20.615 182.595 ;
        RECT 21.345 182.075 21.575 182.595 ;
        RECT 22.305 182.075 22.535 182.595 ;
        RECT 23.265 182.075 23.495 182.595 ;
        RECT 24.225 182.075 24.455 182.595 ;
        RECT 19.855 181.920 20.185 181.935 ;
        RECT 19.840 181.660 20.200 181.920 ;
        RECT 19.855 181.635 20.185 181.660 ;
        RECT 20.415 181.375 20.585 182.075 ;
        RECT 20.815 181.920 21.145 181.935 ;
        RECT 20.795 181.660 21.155 181.920 ;
        RECT 20.815 181.635 21.145 181.660 ;
        RECT 21.375 181.375 21.545 182.075 ;
        RECT 21.775 181.920 22.105 181.935 ;
        RECT 21.755 181.660 22.115 181.920 ;
        RECT 21.775 181.635 22.105 181.660 ;
        RECT 22.335 181.375 22.505 182.075 ;
        RECT 22.735 181.920 23.065 181.935 ;
        RECT 22.715 181.660 23.075 181.920 ;
        RECT 22.735 181.635 23.065 181.660 ;
        RECT 23.295 181.375 23.465 182.075 ;
        RECT 23.695 181.915 24.025 181.935 ;
        RECT 23.680 181.655 24.040 181.915 ;
        RECT 23.695 181.635 24.025 181.655 ;
        RECT 24.255 181.375 24.425 182.075 ;
        RECT 24.655 181.915 24.985 181.935 ;
        RECT 24.640 181.655 25.000 181.915 ;
        RECT 24.655 181.635 24.985 181.655 ;
        RECT 19.015 181.205 24.425 181.375 ;
        RECT 11.410 179.810 16.820 179.980 ;
        RECT 1.535 177.680 1.765 179.040 ;
        RECT 2.495 177.680 2.725 179.040 ;
        RECT 3.455 177.680 3.685 179.040 ;
        RECT 4.415 177.680 4.645 179.040 ;
        RECT 5.375 177.680 5.605 179.040 ;
        RECT 6.335 177.680 6.565 179.040 ;
        RECT 1.565 176.975 1.735 177.680 ;
        RECT 2.525 176.975 2.695 177.680 ;
        RECT 3.485 176.975 3.655 177.680 ;
        RECT 4.445 176.975 4.615 177.680 ;
        RECT 5.405 176.975 5.575 177.680 ;
        RECT 6.365 176.975 6.535 177.680 ;
        RECT 11.410 176.995 11.580 179.810 ;
        RECT 12.810 179.060 12.980 179.810 ;
        RECT 13.770 179.060 13.940 179.810 ;
        RECT 14.730 179.060 14.900 179.810 ;
        RECT 15.690 179.060 15.860 179.810 ;
        RECT 16.650 179.060 16.820 179.810 ;
        RECT 19.015 179.810 24.425 179.980 ;
        RECT 12.300 177.700 12.530 179.060 ;
        RECT 12.780 177.700 13.010 179.060 ;
        RECT 13.260 177.700 13.490 179.060 ;
        RECT 13.740 177.700 13.970 179.060 ;
        RECT 14.220 177.700 14.450 179.060 ;
        RECT 14.700 177.700 14.930 179.060 ;
        RECT 15.180 177.700 15.410 179.060 ;
        RECT 15.660 177.700 15.890 179.060 ;
        RECT 16.140 177.700 16.370 179.060 ;
        RECT 16.620 177.700 16.850 179.060 ;
        RECT 17.100 177.700 17.330 179.060 ;
        RECT 10.505 176.975 11.580 176.995 ;
        RECT 1.565 176.825 11.580 176.975 ;
        RECT 1.565 176.805 10.705 176.825 ;
        RECT 1.565 176.140 1.735 176.805 ;
        RECT 2.525 176.140 2.695 176.805 ;
        RECT 3.485 176.140 3.655 176.805 ;
        RECT 4.445 176.140 4.615 176.805 ;
        RECT 5.405 176.140 5.575 176.805 ;
        RECT 6.365 176.140 6.535 176.805 ;
        RECT 1.535 175.620 1.765 176.140 ;
        RECT 2.495 175.620 2.725 176.140 ;
        RECT 3.455 175.620 3.685 176.140 ;
        RECT 4.415 175.620 4.645 176.140 ;
        RECT 5.375 175.620 5.605 176.140 ;
        RECT 6.335 175.620 6.565 176.140 ;
        RECT 11.410 174.940 11.580 176.825 ;
        RECT 12.330 176.995 12.500 177.700 ;
        RECT 13.290 176.995 13.460 177.700 ;
        RECT 14.250 176.995 14.420 177.700 ;
        RECT 15.210 176.995 15.380 177.700 ;
        RECT 16.170 176.995 16.340 177.700 ;
        RECT 17.130 176.995 17.300 177.700 ;
        RECT 19.015 176.995 19.185 179.810 ;
        RECT 20.415 179.060 20.585 179.810 ;
        RECT 21.375 179.060 21.545 179.810 ;
        RECT 22.335 179.060 22.505 179.810 ;
        RECT 23.295 179.060 23.465 179.810 ;
        RECT 24.255 179.060 24.425 179.810 ;
        RECT 20.385 177.700 20.615 179.060 ;
        RECT 21.345 177.700 21.575 179.060 ;
        RECT 22.305 177.700 22.535 179.060 ;
        RECT 23.265 177.700 23.495 179.060 ;
        RECT 24.225 177.700 24.455 179.060 ;
        RECT 12.330 176.825 19.185 176.995 ;
        RECT 12.330 176.160 12.500 176.825 ;
        RECT 13.290 176.160 13.460 176.825 ;
        RECT 14.250 176.160 14.420 176.825 ;
        RECT 15.210 176.160 15.380 176.825 ;
        RECT 16.170 176.160 16.340 176.825 ;
        RECT 17.130 176.160 17.300 176.825 ;
        RECT 19.015 176.185 19.185 176.825 ;
        RECT 26.630 176.530 27.000 176.800 ;
        RECT 18.670 176.180 19.185 176.185 ;
        RECT 12.300 175.640 12.530 176.160 ;
        RECT 12.780 175.640 13.010 176.160 ;
        RECT 13.260 175.640 13.490 176.160 ;
        RECT 13.740 175.640 13.970 176.160 ;
        RECT 14.220 175.640 14.450 176.160 ;
        RECT 14.700 175.640 14.930 176.160 ;
        RECT 15.180 175.640 15.410 176.160 ;
        RECT 15.660 175.640 15.890 176.160 ;
        RECT 16.140 175.640 16.370 176.160 ;
        RECT 16.620 175.640 16.850 176.160 ;
        RECT 17.100 175.640 17.330 176.160 ;
        RECT 18.645 175.685 19.185 176.180 ;
        RECT 18.645 175.680 18.875 175.685 ;
        RECT 12.250 175.485 12.580 175.500 ;
        RECT 12.235 175.225 12.595 175.485 ;
        RECT 12.250 175.200 12.580 175.225 ;
        RECT 12.810 174.940 12.980 175.640 ;
        RECT 13.210 175.485 13.540 175.500 ;
        RECT 13.190 175.225 13.550 175.485 ;
        RECT 13.210 175.200 13.540 175.225 ;
        RECT 13.770 174.940 13.940 175.640 ;
        RECT 14.170 175.485 14.500 175.500 ;
        RECT 14.150 175.225 14.510 175.485 ;
        RECT 14.170 175.200 14.500 175.225 ;
        RECT 14.730 174.940 14.900 175.640 ;
        RECT 15.130 175.485 15.460 175.500 ;
        RECT 15.110 175.225 15.470 175.485 ;
        RECT 15.130 175.200 15.460 175.225 ;
        RECT 15.690 174.940 15.860 175.640 ;
        RECT 16.090 175.480 16.420 175.500 ;
        RECT 16.075 175.220 16.435 175.480 ;
        RECT 16.090 175.200 16.420 175.220 ;
        RECT 16.650 174.940 16.820 175.640 ;
        RECT 17.050 175.480 17.380 175.500 ;
        RECT 17.035 175.220 17.395 175.480 ;
        RECT 17.050 175.200 17.380 175.220 ;
        RECT 11.410 174.770 16.820 174.940 ;
        RECT 19.015 174.940 19.185 175.685 ;
        RECT 20.385 175.640 20.615 176.160 ;
        RECT 21.345 175.640 21.575 176.160 ;
        RECT 22.305 175.640 22.535 176.160 ;
        RECT 23.265 175.640 23.495 176.160 ;
        RECT 24.225 175.640 24.455 176.160 ;
        RECT 19.855 175.485 20.185 175.500 ;
        RECT 19.840 175.225 20.200 175.485 ;
        RECT 19.855 175.200 20.185 175.225 ;
        RECT 20.415 174.940 20.585 175.640 ;
        RECT 20.815 175.485 21.145 175.500 ;
        RECT 20.795 175.225 21.155 175.485 ;
        RECT 20.815 175.200 21.145 175.225 ;
        RECT 21.375 174.940 21.545 175.640 ;
        RECT 21.775 175.485 22.105 175.500 ;
        RECT 21.755 175.225 22.115 175.485 ;
        RECT 21.775 175.200 22.105 175.225 ;
        RECT 22.335 174.940 22.505 175.640 ;
        RECT 22.735 175.485 23.065 175.500 ;
        RECT 22.715 175.225 23.075 175.485 ;
        RECT 22.735 175.200 23.065 175.225 ;
        RECT 23.295 174.940 23.465 175.640 ;
        RECT 23.695 175.480 24.025 175.500 ;
        RECT 23.680 175.220 24.040 175.480 ;
        RECT 23.695 175.200 24.025 175.220 ;
        RECT 24.255 174.940 24.425 175.640 ;
        RECT 24.655 175.480 24.985 175.500 ;
        RECT 24.640 175.220 25.000 175.480 ;
        RECT 24.655 175.200 24.985 175.220 ;
        RECT 19.015 174.770 24.425 174.940 ;
        RECT 11.410 173.375 16.820 173.545 ;
        RECT 1.535 171.245 1.765 172.605 ;
        RECT 2.495 171.245 2.725 172.605 ;
        RECT 3.455 171.245 3.685 172.605 ;
        RECT 4.415 171.245 4.645 172.605 ;
        RECT 5.375 171.245 5.605 172.605 ;
        RECT 6.335 171.245 6.565 172.605 ;
        RECT 1.565 170.540 1.735 171.245 ;
        RECT 2.525 170.540 2.695 171.245 ;
        RECT 3.485 170.540 3.655 171.245 ;
        RECT 4.445 170.540 4.615 171.245 ;
        RECT 5.405 170.540 5.575 171.245 ;
        RECT 6.365 170.540 6.535 171.245 ;
        RECT 11.410 170.560 11.580 173.375 ;
        RECT 12.810 172.625 12.980 173.375 ;
        RECT 13.770 172.625 13.940 173.375 ;
        RECT 14.730 172.625 14.900 173.375 ;
        RECT 15.690 172.625 15.860 173.375 ;
        RECT 16.650 172.625 16.820 173.375 ;
        RECT 19.015 173.375 24.425 173.545 ;
        RECT 12.300 171.265 12.530 172.625 ;
        RECT 12.780 171.265 13.010 172.625 ;
        RECT 13.260 171.265 13.490 172.625 ;
        RECT 13.740 171.265 13.970 172.625 ;
        RECT 14.220 171.265 14.450 172.625 ;
        RECT 14.700 171.265 14.930 172.625 ;
        RECT 15.180 171.265 15.410 172.625 ;
        RECT 15.660 171.265 15.890 172.625 ;
        RECT 16.140 171.265 16.370 172.625 ;
        RECT 16.620 171.265 16.850 172.625 ;
        RECT 17.100 171.265 17.330 172.625 ;
        RECT 10.505 170.540 11.580 170.560 ;
        RECT 1.565 170.390 11.580 170.540 ;
        RECT 1.565 170.370 10.705 170.390 ;
        RECT 1.565 169.705 1.735 170.370 ;
        RECT 2.525 169.705 2.695 170.370 ;
        RECT 3.485 169.705 3.655 170.370 ;
        RECT 4.445 169.705 4.615 170.370 ;
        RECT 5.405 169.705 5.575 170.370 ;
        RECT 6.365 169.705 6.535 170.370 ;
        RECT 1.535 169.185 1.765 169.705 ;
        RECT 2.495 169.185 2.725 169.705 ;
        RECT 3.455 169.185 3.685 169.705 ;
        RECT 4.415 169.185 4.645 169.705 ;
        RECT 5.375 169.185 5.605 169.705 ;
        RECT 6.335 169.185 6.565 169.705 ;
        RECT 11.410 168.505 11.580 170.390 ;
        RECT 12.330 170.560 12.500 171.265 ;
        RECT 13.290 170.560 13.460 171.265 ;
        RECT 14.250 170.560 14.420 171.265 ;
        RECT 15.210 170.560 15.380 171.265 ;
        RECT 16.170 170.560 16.340 171.265 ;
        RECT 17.130 170.560 17.300 171.265 ;
        RECT 19.015 170.560 19.185 173.375 ;
        RECT 20.415 172.625 20.585 173.375 ;
        RECT 21.375 172.625 21.545 173.375 ;
        RECT 22.335 172.625 22.505 173.375 ;
        RECT 23.295 172.625 23.465 173.375 ;
        RECT 24.255 172.625 24.425 173.375 ;
        RECT 20.385 171.265 20.615 172.625 ;
        RECT 21.345 171.265 21.575 172.625 ;
        RECT 22.305 171.265 22.535 172.625 ;
        RECT 23.265 171.265 23.495 172.625 ;
        RECT 24.225 171.265 24.455 172.625 ;
        RECT 12.330 170.390 19.185 170.560 ;
        RECT 12.330 169.725 12.500 170.390 ;
        RECT 13.290 169.725 13.460 170.390 ;
        RECT 14.250 169.725 14.420 170.390 ;
        RECT 15.210 169.725 15.380 170.390 ;
        RECT 16.170 169.725 16.340 170.390 ;
        RECT 17.130 169.725 17.300 170.390 ;
        RECT 19.015 169.750 19.185 170.390 ;
        RECT 26.630 170.095 27.000 170.365 ;
        RECT 18.670 169.745 19.185 169.750 ;
        RECT 12.300 169.205 12.530 169.725 ;
        RECT 12.780 169.205 13.010 169.725 ;
        RECT 13.260 169.205 13.490 169.725 ;
        RECT 13.740 169.205 13.970 169.725 ;
        RECT 14.220 169.205 14.450 169.725 ;
        RECT 14.700 169.205 14.930 169.725 ;
        RECT 15.180 169.205 15.410 169.725 ;
        RECT 15.660 169.205 15.890 169.725 ;
        RECT 16.140 169.205 16.370 169.725 ;
        RECT 16.620 169.205 16.850 169.725 ;
        RECT 17.100 169.205 17.330 169.725 ;
        RECT 18.645 169.250 19.185 169.745 ;
        RECT 18.645 169.245 18.875 169.250 ;
        RECT 12.250 169.050 12.580 169.065 ;
        RECT 12.235 168.790 12.595 169.050 ;
        RECT 12.250 168.765 12.580 168.790 ;
        RECT 12.810 168.505 12.980 169.205 ;
        RECT 13.210 169.050 13.540 169.065 ;
        RECT 13.190 168.790 13.550 169.050 ;
        RECT 13.210 168.765 13.540 168.790 ;
        RECT 13.770 168.505 13.940 169.205 ;
        RECT 14.170 169.050 14.500 169.065 ;
        RECT 14.150 168.790 14.510 169.050 ;
        RECT 14.170 168.765 14.500 168.790 ;
        RECT 14.730 168.505 14.900 169.205 ;
        RECT 15.130 169.050 15.460 169.065 ;
        RECT 15.110 168.790 15.470 169.050 ;
        RECT 15.130 168.765 15.460 168.790 ;
        RECT 15.690 168.505 15.860 169.205 ;
        RECT 16.090 169.045 16.420 169.065 ;
        RECT 16.075 168.785 16.435 169.045 ;
        RECT 16.090 168.765 16.420 168.785 ;
        RECT 16.650 168.505 16.820 169.205 ;
        RECT 17.050 169.045 17.380 169.065 ;
        RECT 17.035 168.785 17.395 169.045 ;
        RECT 17.050 168.765 17.380 168.785 ;
        RECT 11.410 168.335 16.820 168.505 ;
        RECT 19.015 168.505 19.185 169.250 ;
        RECT 20.385 169.205 20.615 169.725 ;
        RECT 21.345 169.205 21.575 169.725 ;
        RECT 22.305 169.205 22.535 169.725 ;
        RECT 23.265 169.205 23.495 169.725 ;
        RECT 24.225 169.205 24.455 169.725 ;
        RECT 19.855 169.050 20.185 169.065 ;
        RECT 19.840 168.790 20.200 169.050 ;
        RECT 19.855 168.765 20.185 168.790 ;
        RECT 20.415 168.505 20.585 169.205 ;
        RECT 20.815 169.050 21.145 169.065 ;
        RECT 20.795 168.790 21.155 169.050 ;
        RECT 20.815 168.765 21.145 168.790 ;
        RECT 21.375 168.505 21.545 169.205 ;
        RECT 21.775 169.050 22.105 169.065 ;
        RECT 21.755 168.790 22.115 169.050 ;
        RECT 21.775 168.765 22.105 168.790 ;
        RECT 22.335 168.505 22.505 169.205 ;
        RECT 22.735 169.050 23.065 169.065 ;
        RECT 22.715 168.790 23.075 169.050 ;
        RECT 22.735 168.765 23.065 168.790 ;
        RECT 23.295 168.505 23.465 169.205 ;
        RECT 23.695 169.045 24.025 169.065 ;
        RECT 23.680 168.785 24.040 169.045 ;
        RECT 23.695 168.765 24.025 168.785 ;
        RECT 24.255 168.505 24.425 169.205 ;
        RECT 24.655 169.045 24.985 169.065 ;
        RECT 24.640 168.785 25.000 169.045 ;
        RECT 24.655 168.765 24.985 168.785 ;
        RECT 19.015 168.335 24.425 168.505 ;
        RECT 11.410 166.940 16.820 167.110 ;
        RECT 1.535 164.810 1.765 166.170 ;
        RECT 2.495 164.810 2.725 166.170 ;
        RECT 3.455 164.810 3.685 166.170 ;
        RECT 4.415 164.810 4.645 166.170 ;
        RECT 5.375 164.810 5.605 166.170 ;
        RECT 6.335 164.810 6.565 166.170 ;
        RECT 1.565 164.105 1.735 164.810 ;
        RECT 2.525 164.105 2.695 164.810 ;
        RECT 3.485 164.105 3.655 164.810 ;
        RECT 4.445 164.105 4.615 164.810 ;
        RECT 5.405 164.105 5.575 164.810 ;
        RECT 6.365 164.105 6.535 164.810 ;
        RECT 11.410 164.125 11.580 166.940 ;
        RECT 12.810 166.190 12.980 166.940 ;
        RECT 13.770 166.190 13.940 166.940 ;
        RECT 14.730 166.190 14.900 166.940 ;
        RECT 15.690 166.190 15.860 166.940 ;
        RECT 16.650 166.190 16.820 166.940 ;
        RECT 19.015 166.940 24.425 167.110 ;
        RECT 12.300 164.830 12.530 166.190 ;
        RECT 12.780 164.830 13.010 166.190 ;
        RECT 13.260 164.830 13.490 166.190 ;
        RECT 13.740 164.830 13.970 166.190 ;
        RECT 14.220 164.830 14.450 166.190 ;
        RECT 14.700 164.830 14.930 166.190 ;
        RECT 15.180 164.830 15.410 166.190 ;
        RECT 15.660 164.830 15.890 166.190 ;
        RECT 16.140 164.830 16.370 166.190 ;
        RECT 16.620 164.830 16.850 166.190 ;
        RECT 17.100 164.830 17.330 166.190 ;
        RECT 10.505 164.105 11.580 164.125 ;
        RECT 1.565 163.955 11.580 164.105 ;
        RECT 1.565 163.935 10.705 163.955 ;
        RECT 1.565 163.270 1.735 163.935 ;
        RECT 2.525 163.270 2.695 163.935 ;
        RECT 3.485 163.270 3.655 163.935 ;
        RECT 4.445 163.270 4.615 163.935 ;
        RECT 5.405 163.270 5.575 163.935 ;
        RECT 6.365 163.270 6.535 163.935 ;
        RECT 1.535 162.750 1.765 163.270 ;
        RECT 2.495 162.750 2.725 163.270 ;
        RECT 3.455 162.750 3.685 163.270 ;
        RECT 4.415 162.750 4.645 163.270 ;
        RECT 5.375 162.750 5.605 163.270 ;
        RECT 6.335 162.750 6.565 163.270 ;
        RECT 11.410 162.070 11.580 163.955 ;
        RECT 12.330 164.125 12.500 164.830 ;
        RECT 13.290 164.125 13.460 164.830 ;
        RECT 14.250 164.125 14.420 164.830 ;
        RECT 15.210 164.125 15.380 164.830 ;
        RECT 16.170 164.125 16.340 164.830 ;
        RECT 17.130 164.125 17.300 164.830 ;
        RECT 19.015 164.125 19.185 166.940 ;
        RECT 20.415 166.190 20.585 166.940 ;
        RECT 21.375 166.190 21.545 166.940 ;
        RECT 22.335 166.190 22.505 166.940 ;
        RECT 23.295 166.190 23.465 166.940 ;
        RECT 24.255 166.190 24.425 166.940 ;
        RECT 20.385 164.830 20.615 166.190 ;
        RECT 21.345 164.830 21.575 166.190 ;
        RECT 22.305 164.830 22.535 166.190 ;
        RECT 23.265 164.830 23.495 166.190 ;
        RECT 24.225 164.830 24.455 166.190 ;
        RECT 12.330 163.955 19.185 164.125 ;
        RECT 12.330 163.290 12.500 163.955 ;
        RECT 13.290 163.290 13.460 163.955 ;
        RECT 14.250 163.290 14.420 163.955 ;
        RECT 15.210 163.290 15.380 163.955 ;
        RECT 16.170 163.290 16.340 163.955 ;
        RECT 17.130 163.290 17.300 163.955 ;
        RECT 19.015 163.315 19.185 163.955 ;
        RECT 26.630 163.660 27.000 163.930 ;
        RECT 18.670 163.310 19.185 163.315 ;
        RECT 12.300 162.770 12.530 163.290 ;
        RECT 12.780 162.770 13.010 163.290 ;
        RECT 13.260 162.770 13.490 163.290 ;
        RECT 13.740 162.770 13.970 163.290 ;
        RECT 14.220 162.770 14.450 163.290 ;
        RECT 14.700 162.770 14.930 163.290 ;
        RECT 15.180 162.770 15.410 163.290 ;
        RECT 15.660 162.770 15.890 163.290 ;
        RECT 16.140 162.770 16.370 163.290 ;
        RECT 16.620 162.770 16.850 163.290 ;
        RECT 17.100 162.770 17.330 163.290 ;
        RECT 18.645 162.815 19.185 163.310 ;
        RECT 18.645 162.810 18.875 162.815 ;
        RECT 12.250 162.615 12.580 162.630 ;
        RECT 12.235 162.355 12.595 162.615 ;
        RECT 12.250 162.330 12.580 162.355 ;
        RECT 12.810 162.070 12.980 162.770 ;
        RECT 13.210 162.615 13.540 162.630 ;
        RECT 13.190 162.355 13.550 162.615 ;
        RECT 13.210 162.330 13.540 162.355 ;
        RECT 13.770 162.070 13.940 162.770 ;
        RECT 14.170 162.615 14.500 162.630 ;
        RECT 14.150 162.355 14.510 162.615 ;
        RECT 14.170 162.330 14.500 162.355 ;
        RECT 14.730 162.070 14.900 162.770 ;
        RECT 15.130 162.615 15.460 162.630 ;
        RECT 15.110 162.355 15.470 162.615 ;
        RECT 15.130 162.330 15.460 162.355 ;
        RECT 15.690 162.070 15.860 162.770 ;
        RECT 16.090 162.610 16.420 162.630 ;
        RECT 16.075 162.350 16.435 162.610 ;
        RECT 16.090 162.330 16.420 162.350 ;
        RECT 16.650 162.070 16.820 162.770 ;
        RECT 17.050 162.610 17.380 162.630 ;
        RECT 17.035 162.350 17.395 162.610 ;
        RECT 17.050 162.330 17.380 162.350 ;
        RECT 11.410 161.900 16.820 162.070 ;
        RECT 19.015 162.070 19.185 162.815 ;
        RECT 20.385 162.770 20.615 163.290 ;
        RECT 21.345 162.770 21.575 163.290 ;
        RECT 22.305 162.770 22.535 163.290 ;
        RECT 23.265 162.770 23.495 163.290 ;
        RECT 24.225 162.770 24.455 163.290 ;
        RECT 19.855 162.615 20.185 162.630 ;
        RECT 19.840 162.355 20.200 162.615 ;
        RECT 19.855 162.330 20.185 162.355 ;
        RECT 20.415 162.070 20.585 162.770 ;
        RECT 20.815 162.615 21.145 162.630 ;
        RECT 20.795 162.355 21.155 162.615 ;
        RECT 20.815 162.330 21.145 162.355 ;
        RECT 21.375 162.070 21.545 162.770 ;
        RECT 21.775 162.615 22.105 162.630 ;
        RECT 21.755 162.355 22.115 162.615 ;
        RECT 21.775 162.330 22.105 162.355 ;
        RECT 22.335 162.070 22.505 162.770 ;
        RECT 22.735 162.615 23.065 162.630 ;
        RECT 22.715 162.355 23.075 162.615 ;
        RECT 22.735 162.330 23.065 162.355 ;
        RECT 23.295 162.070 23.465 162.770 ;
        RECT 23.695 162.610 24.025 162.630 ;
        RECT 23.680 162.350 24.040 162.610 ;
        RECT 23.695 162.330 24.025 162.350 ;
        RECT 24.255 162.070 24.425 162.770 ;
        RECT 24.655 162.610 24.985 162.630 ;
        RECT 24.640 162.350 25.000 162.610 ;
        RECT 24.655 162.330 24.985 162.350 ;
        RECT 19.015 161.900 24.425 162.070 ;
        RECT 11.410 160.505 16.820 160.675 ;
        RECT 1.535 158.375 1.765 159.735 ;
        RECT 2.495 158.375 2.725 159.735 ;
        RECT 3.455 158.375 3.685 159.735 ;
        RECT 4.415 158.375 4.645 159.735 ;
        RECT 5.375 158.375 5.605 159.735 ;
        RECT 6.335 158.375 6.565 159.735 ;
        RECT 1.565 157.670 1.735 158.375 ;
        RECT 2.525 157.670 2.695 158.375 ;
        RECT 3.485 157.670 3.655 158.375 ;
        RECT 4.445 157.670 4.615 158.375 ;
        RECT 5.405 157.670 5.575 158.375 ;
        RECT 6.365 157.670 6.535 158.375 ;
        RECT 11.410 157.690 11.580 160.505 ;
        RECT 12.810 159.755 12.980 160.505 ;
        RECT 13.770 159.755 13.940 160.505 ;
        RECT 14.730 159.755 14.900 160.505 ;
        RECT 15.690 159.755 15.860 160.505 ;
        RECT 16.650 159.755 16.820 160.505 ;
        RECT 19.015 160.505 24.425 160.675 ;
        RECT 12.300 158.395 12.530 159.755 ;
        RECT 12.780 158.395 13.010 159.755 ;
        RECT 13.260 158.395 13.490 159.755 ;
        RECT 13.740 158.395 13.970 159.755 ;
        RECT 14.220 158.395 14.450 159.755 ;
        RECT 14.700 158.395 14.930 159.755 ;
        RECT 15.180 158.395 15.410 159.755 ;
        RECT 15.660 158.395 15.890 159.755 ;
        RECT 16.140 158.395 16.370 159.755 ;
        RECT 16.620 158.395 16.850 159.755 ;
        RECT 17.100 158.395 17.330 159.755 ;
        RECT 10.505 157.670 11.580 157.690 ;
        RECT 1.565 157.520 11.580 157.670 ;
        RECT 1.565 157.500 10.705 157.520 ;
        RECT 1.565 156.835 1.735 157.500 ;
        RECT 2.525 156.835 2.695 157.500 ;
        RECT 3.485 156.835 3.655 157.500 ;
        RECT 4.445 156.835 4.615 157.500 ;
        RECT 5.405 156.835 5.575 157.500 ;
        RECT 6.365 156.835 6.535 157.500 ;
        RECT 1.535 156.315 1.765 156.835 ;
        RECT 2.495 156.315 2.725 156.835 ;
        RECT 3.455 156.315 3.685 156.835 ;
        RECT 4.415 156.315 4.645 156.835 ;
        RECT 5.375 156.315 5.605 156.835 ;
        RECT 6.335 156.315 6.565 156.835 ;
        RECT 11.410 155.635 11.580 157.520 ;
        RECT 12.330 157.690 12.500 158.395 ;
        RECT 13.290 157.690 13.460 158.395 ;
        RECT 14.250 157.690 14.420 158.395 ;
        RECT 15.210 157.690 15.380 158.395 ;
        RECT 16.170 157.690 16.340 158.395 ;
        RECT 17.130 157.690 17.300 158.395 ;
        RECT 19.015 157.690 19.185 160.505 ;
        RECT 20.415 159.755 20.585 160.505 ;
        RECT 21.375 159.755 21.545 160.505 ;
        RECT 22.335 159.755 22.505 160.505 ;
        RECT 23.295 159.755 23.465 160.505 ;
        RECT 24.255 159.755 24.425 160.505 ;
        RECT 20.385 158.395 20.615 159.755 ;
        RECT 21.345 158.395 21.575 159.755 ;
        RECT 22.305 158.395 22.535 159.755 ;
        RECT 23.265 158.395 23.495 159.755 ;
        RECT 24.225 158.395 24.455 159.755 ;
        RECT 12.330 157.520 19.185 157.690 ;
        RECT 12.330 156.855 12.500 157.520 ;
        RECT 13.290 156.855 13.460 157.520 ;
        RECT 14.250 156.855 14.420 157.520 ;
        RECT 15.210 156.855 15.380 157.520 ;
        RECT 16.170 156.855 16.340 157.520 ;
        RECT 17.130 156.855 17.300 157.520 ;
        RECT 19.015 156.880 19.185 157.520 ;
        RECT 26.630 157.225 27.000 157.495 ;
        RECT 18.670 156.875 19.185 156.880 ;
        RECT 12.300 156.335 12.530 156.855 ;
        RECT 12.780 156.335 13.010 156.855 ;
        RECT 13.260 156.335 13.490 156.855 ;
        RECT 13.740 156.335 13.970 156.855 ;
        RECT 14.220 156.335 14.450 156.855 ;
        RECT 14.700 156.335 14.930 156.855 ;
        RECT 15.180 156.335 15.410 156.855 ;
        RECT 15.660 156.335 15.890 156.855 ;
        RECT 16.140 156.335 16.370 156.855 ;
        RECT 16.620 156.335 16.850 156.855 ;
        RECT 17.100 156.335 17.330 156.855 ;
        RECT 18.645 156.380 19.185 156.875 ;
        RECT 18.645 156.375 18.875 156.380 ;
        RECT 12.250 156.180 12.580 156.195 ;
        RECT 12.235 155.920 12.595 156.180 ;
        RECT 12.250 155.895 12.580 155.920 ;
        RECT 12.810 155.635 12.980 156.335 ;
        RECT 13.210 156.180 13.540 156.195 ;
        RECT 13.190 155.920 13.550 156.180 ;
        RECT 13.210 155.895 13.540 155.920 ;
        RECT 13.770 155.635 13.940 156.335 ;
        RECT 14.170 156.180 14.500 156.195 ;
        RECT 14.150 155.920 14.510 156.180 ;
        RECT 14.170 155.895 14.500 155.920 ;
        RECT 14.730 155.635 14.900 156.335 ;
        RECT 15.130 156.180 15.460 156.195 ;
        RECT 15.110 155.920 15.470 156.180 ;
        RECT 15.130 155.895 15.460 155.920 ;
        RECT 15.690 155.635 15.860 156.335 ;
        RECT 16.090 156.175 16.420 156.195 ;
        RECT 16.075 155.915 16.435 156.175 ;
        RECT 16.090 155.895 16.420 155.915 ;
        RECT 16.650 155.635 16.820 156.335 ;
        RECT 17.050 156.175 17.380 156.195 ;
        RECT 17.035 155.915 17.395 156.175 ;
        RECT 17.050 155.895 17.380 155.915 ;
        RECT 11.410 155.465 16.820 155.635 ;
        RECT 19.015 155.635 19.185 156.380 ;
        RECT 20.385 156.335 20.615 156.855 ;
        RECT 21.345 156.335 21.575 156.855 ;
        RECT 22.305 156.335 22.535 156.855 ;
        RECT 23.265 156.335 23.495 156.855 ;
        RECT 24.225 156.335 24.455 156.855 ;
        RECT 19.855 156.180 20.185 156.195 ;
        RECT 19.840 155.920 20.200 156.180 ;
        RECT 19.855 155.895 20.185 155.920 ;
        RECT 20.415 155.635 20.585 156.335 ;
        RECT 20.815 156.180 21.145 156.195 ;
        RECT 20.795 155.920 21.155 156.180 ;
        RECT 20.815 155.895 21.145 155.920 ;
        RECT 21.375 155.635 21.545 156.335 ;
        RECT 21.775 156.180 22.105 156.195 ;
        RECT 21.755 155.920 22.115 156.180 ;
        RECT 21.775 155.895 22.105 155.920 ;
        RECT 22.335 155.635 22.505 156.335 ;
        RECT 22.735 156.180 23.065 156.195 ;
        RECT 22.715 155.920 23.075 156.180 ;
        RECT 22.735 155.895 23.065 155.920 ;
        RECT 23.295 155.635 23.465 156.335 ;
        RECT 23.695 156.175 24.025 156.195 ;
        RECT 23.680 155.915 24.040 156.175 ;
        RECT 23.695 155.895 24.025 155.915 ;
        RECT 24.255 155.635 24.425 156.335 ;
        RECT 24.655 156.175 24.985 156.195 ;
        RECT 24.640 155.915 25.000 156.175 ;
        RECT 24.655 155.895 24.985 155.915 ;
        RECT 19.015 155.465 24.425 155.635 ;
        RECT 11.410 154.070 16.820 154.240 ;
        RECT 1.535 151.940 1.765 153.300 ;
        RECT 2.495 151.940 2.725 153.300 ;
        RECT 3.455 151.940 3.685 153.300 ;
        RECT 4.415 151.940 4.645 153.300 ;
        RECT 5.375 151.940 5.605 153.300 ;
        RECT 6.335 151.940 6.565 153.300 ;
        RECT 1.565 151.235 1.735 151.940 ;
        RECT 2.525 151.235 2.695 151.940 ;
        RECT 3.485 151.235 3.655 151.940 ;
        RECT 4.445 151.235 4.615 151.940 ;
        RECT 5.405 151.235 5.575 151.940 ;
        RECT 6.365 151.235 6.535 151.940 ;
        RECT 11.410 151.255 11.580 154.070 ;
        RECT 12.810 153.320 12.980 154.070 ;
        RECT 13.770 153.320 13.940 154.070 ;
        RECT 14.730 153.320 14.900 154.070 ;
        RECT 15.690 153.320 15.860 154.070 ;
        RECT 16.650 153.320 16.820 154.070 ;
        RECT 19.015 154.070 24.425 154.240 ;
        RECT 12.300 151.960 12.530 153.320 ;
        RECT 12.780 151.960 13.010 153.320 ;
        RECT 13.260 151.960 13.490 153.320 ;
        RECT 13.740 151.960 13.970 153.320 ;
        RECT 14.220 151.960 14.450 153.320 ;
        RECT 14.700 151.960 14.930 153.320 ;
        RECT 15.180 151.960 15.410 153.320 ;
        RECT 15.660 151.960 15.890 153.320 ;
        RECT 16.140 151.960 16.370 153.320 ;
        RECT 16.620 151.960 16.850 153.320 ;
        RECT 17.100 151.960 17.330 153.320 ;
        RECT 10.505 151.235 11.580 151.255 ;
        RECT 1.565 151.085 11.580 151.235 ;
        RECT 1.565 151.065 10.705 151.085 ;
        RECT 1.565 150.400 1.735 151.065 ;
        RECT 2.525 150.400 2.695 151.065 ;
        RECT 3.485 150.400 3.655 151.065 ;
        RECT 4.445 150.400 4.615 151.065 ;
        RECT 5.405 150.400 5.575 151.065 ;
        RECT 6.365 150.400 6.535 151.065 ;
        RECT 1.535 149.880 1.765 150.400 ;
        RECT 2.495 149.880 2.725 150.400 ;
        RECT 3.455 149.880 3.685 150.400 ;
        RECT 4.415 149.880 4.645 150.400 ;
        RECT 5.375 149.880 5.605 150.400 ;
        RECT 6.335 149.880 6.565 150.400 ;
        RECT 11.410 149.200 11.580 151.085 ;
        RECT 12.330 151.255 12.500 151.960 ;
        RECT 13.290 151.255 13.460 151.960 ;
        RECT 14.250 151.255 14.420 151.960 ;
        RECT 15.210 151.255 15.380 151.960 ;
        RECT 16.170 151.255 16.340 151.960 ;
        RECT 17.130 151.255 17.300 151.960 ;
        RECT 19.015 151.255 19.185 154.070 ;
        RECT 20.415 153.320 20.585 154.070 ;
        RECT 21.375 153.320 21.545 154.070 ;
        RECT 22.335 153.320 22.505 154.070 ;
        RECT 23.295 153.320 23.465 154.070 ;
        RECT 24.255 153.320 24.425 154.070 ;
        RECT 20.385 151.960 20.615 153.320 ;
        RECT 21.345 151.960 21.575 153.320 ;
        RECT 22.305 151.960 22.535 153.320 ;
        RECT 23.265 151.960 23.495 153.320 ;
        RECT 24.225 151.960 24.455 153.320 ;
        RECT 12.330 151.085 19.185 151.255 ;
        RECT 12.330 150.420 12.500 151.085 ;
        RECT 13.290 150.420 13.460 151.085 ;
        RECT 14.250 150.420 14.420 151.085 ;
        RECT 15.210 150.420 15.380 151.085 ;
        RECT 16.170 150.420 16.340 151.085 ;
        RECT 17.130 150.420 17.300 151.085 ;
        RECT 19.015 150.445 19.185 151.085 ;
        RECT 26.630 150.790 27.000 151.060 ;
        RECT 18.670 150.440 19.185 150.445 ;
        RECT 12.300 149.900 12.530 150.420 ;
        RECT 12.780 149.900 13.010 150.420 ;
        RECT 13.260 149.900 13.490 150.420 ;
        RECT 13.740 149.900 13.970 150.420 ;
        RECT 14.220 149.900 14.450 150.420 ;
        RECT 14.700 149.900 14.930 150.420 ;
        RECT 15.180 149.900 15.410 150.420 ;
        RECT 15.660 149.900 15.890 150.420 ;
        RECT 16.140 149.900 16.370 150.420 ;
        RECT 16.620 149.900 16.850 150.420 ;
        RECT 17.100 149.900 17.330 150.420 ;
        RECT 18.645 149.945 19.185 150.440 ;
        RECT 18.645 149.940 18.875 149.945 ;
        RECT 12.250 149.745 12.580 149.760 ;
        RECT 12.235 149.485 12.595 149.745 ;
        RECT 12.250 149.460 12.580 149.485 ;
        RECT 12.810 149.200 12.980 149.900 ;
        RECT 13.210 149.745 13.540 149.760 ;
        RECT 13.190 149.485 13.550 149.745 ;
        RECT 13.210 149.460 13.540 149.485 ;
        RECT 13.770 149.200 13.940 149.900 ;
        RECT 14.170 149.745 14.500 149.760 ;
        RECT 14.150 149.485 14.510 149.745 ;
        RECT 14.170 149.460 14.500 149.485 ;
        RECT 14.730 149.200 14.900 149.900 ;
        RECT 15.130 149.745 15.460 149.760 ;
        RECT 15.110 149.485 15.470 149.745 ;
        RECT 15.130 149.460 15.460 149.485 ;
        RECT 15.690 149.200 15.860 149.900 ;
        RECT 16.090 149.740 16.420 149.760 ;
        RECT 16.075 149.480 16.435 149.740 ;
        RECT 16.090 149.460 16.420 149.480 ;
        RECT 16.650 149.200 16.820 149.900 ;
        RECT 17.050 149.740 17.380 149.760 ;
        RECT 17.035 149.480 17.395 149.740 ;
        RECT 17.050 149.460 17.380 149.480 ;
        RECT 11.410 149.030 16.820 149.200 ;
        RECT 19.015 149.200 19.185 149.945 ;
        RECT 20.385 149.900 20.615 150.420 ;
        RECT 21.345 149.900 21.575 150.420 ;
        RECT 22.305 149.900 22.535 150.420 ;
        RECT 23.265 149.900 23.495 150.420 ;
        RECT 24.225 149.900 24.455 150.420 ;
        RECT 19.855 149.745 20.185 149.760 ;
        RECT 19.840 149.485 20.200 149.745 ;
        RECT 19.855 149.460 20.185 149.485 ;
        RECT 20.415 149.200 20.585 149.900 ;
        RECT 20.815 149.745 21.145 149.760 ;
        RECT 20.795 149.485 21.155 149.745 ;
        RECT 20.815 149.460 21.145 149.485 ;
        RECT 21.375 149.200 21.545 149.900 ;
        RECT 21.775 149.745 22.105 149.760 ;
        RECT 21.755 149.485 22.115 149.745 ;
        RECT 21.775 149.460 22.105 149.485 ;
        RECT 22.335 149.200 22.505 149.900 ;
        RECT 22.735 149.745 23.065 149.760 ;
        RECT 22.715 149.485 23.075 149.745 ;
        RECT 22.735 149.460 23.065 149.485 ;
        RECT 23.295 149.200 23.465 149.900 ;
        RECT 23.695 149.740 24.025 149.760 ;
        RECT 23.680 149.480 24.040 149.740 ;
        RECT 23.695 149.460 24.025 149.480 ;
        RECT 24.255 149.200 24.425 149.900 ;
        RECT 24.655 149.740 24.985 149.760 ;
        RECT 24.640 149.480 25.000 149.740 ;
        RECT 24.655 149.460 24.985 149.480 ;
        RECT 19.015 149.030 24.425 149.200 ;
        RECT 11.410 147.635 16.820 147.805 ;
        RECT 1.535 145.505 1.765 146.865 ;
        RECT 2.495 145.505 2.725 146.865 ;
        RECT 3.455 145.505 3.685 146.865 ;
        RECT 4.415 145.505 4.645 146.865 ;
        RECT 5.375 145.505 5.605 146.865 ;
        RECT 6.335 145.505 6.565 146.865 ;
        RECT 1.565 144.800 1.735 145.505 ;
        RECT 2.525 144.800 2.695 145.505 ;
        RECT 3.485 144.800 3.655 145.505 ;
        RECT 4.445 144.800 4.615 145.505 ;
        RECT 5.405 144.800 5.575 145.505 ;
        RECT 6.365 144.800 6.535 145.505 ;
        RECT 11.410 144.820 11.580 147.635 ;
        RECT 12.810 146.885 12.980 147.635 ;
        RECT 13.770 146.885 13.940 147.635 ;
        RECT 14.730 146.885 14.900 147.635 ;
        RECT 15.690 146.885 15.860 147.635 ;
        RECT 16.650 146.885 16.820 147.635 ;
        RECT 19.015 147.635 24.425 147.805 ;
        RECT 12.300 145.525 12.530 146.885 ;
        RECT 12.780 145.525 13.010 146.885 ;
        RECT 13.260 145.525 13.490 146.885 ;
        RECT 13.740 145.525 13.970 146.885 ;
        RECT 14.220 145.525 14.450 146.885 ;
        RECT 14.700 145.525 14.930 146.885 ;
        RECT 15.180 145.525 15.410 146.885 ;
        RECT 15.660 145.525 15.890 146.885 ;
        RECT 16.140 145.525 16.370 146.885 ;
        RECT 16.620 145.525 16.850 146.885 ;
        RECT 17.100 145.525 17.330 146.885 ;
        RECT 10.505 144.800 11.580 144.820 ;
        RECT 1.565 144.650 11.580 144.800 ;
        RECT 1.565 144.630 10.705 144.650 ;
        RECT 1.565 143.965 1.735 144.630 ;
        RECT 2.525 143.965 2.695 144.630 ;
        RECT 3.485 143.965 3.655 144.630 ;
        RECT 4.445 143.965 4.615 144.630 ;
        RECT 5.405 143.965 5.575 144.630 ;
        RECT 6.365 143.965 6.535 144.630 ;
        RECT 1.535 143.445 1.765 143.965 ;
        RECT 2.495 143.445 2.725 143.965 ;
        RECT 3.455 143.445 3.685 143.965 ;
        RECT 4.415 143.445 4.645 143.965 ;
        RECT 5.375 143.445 5.605 143.965 ;
        RECT 6.335 143.445 6.565 143.965 ;
        RECT 11.410 142.765 11.580 144.650 ;
        RECT 12.330 144.820 12.500 145.525 ;
        RECT 13.290 144.820 13.460 145.525 ;
        RECT 14.250 144.820 14.420 145.525 ;
        RECT 15.210 144.820 15.380 145.525 ;
        RECT 16.170 144.820 16.340 145.525 ;
        RECT 17.130 144.820 17.300 145.525 ;
        RECT 19.015 144.820 19.185 147.635 ;
        RECT 20.415 146.885 20.585 147.635 ;
        RECT 21.375 146.885 21.545 147.635 ;
        RECT 22.335 146.885 22.505 147.635 ;
        RECT 23.295 146.885 23.465 147.635 ;
        RECT 24.255 146.885 24.425 147.635 ;
        RECT 20.385 145.525 20.615 146.885 ;
        RECT 21.345 145.525 21.575 146.885 ;
        RECT 22.305 145.525 22.535 146.885 ;
        RECT 23.265 145.525 23.495 146.885 ;
        RECT 24.225 145.525 24.455 146.885 ;
        RECT 12.330 144.650 19.185 144.820 ;
        RECT 12.330 143.985 12.500 144.650 ;
        RECT 13.290 143.985 13.460 144.650 ;
        RECT 14.250 143.985 14.420 144.650 ;
        RECT 15.210 143.985 15.380 144.650 ;
        RECT 16.170 143.985 16.340 144.650 ;
        RECT 17.130 143.985 17.300 144.650 ;
        RECT 19.015 144.010 19.185 144.650 ;
        RECT 26.630 144.355 27.000 144.625 ;
        RECT 18.670 144.005 19.185 144.010 ;
        RECT 12.300 143.465 12.530 143.985 ;
        RECT 12.780 143.465 13.010 143.985 ;
        RECT 13.260 143.465 13.490 143.985 ;
        RECT 13.740 143.465 13.970 143.985 ;
        RECT 14.220 143.465 14.450 143.985 ;
        RECT 14.700 143.465 14.930 143.985 ;
        RECT 15.180 143.465 15.410 143.985 ;
        RECT 15.660 143.465 15.890 143.985 ;
        RECT 16.140 143.465 16.370 143.985 ;
        RECT 16.620 143.465 16.850 143.985 ;
        RECT 17.100 143.465 17.330 143.985 ;
        RECT 18.645 143.510 19.185 144.005 ;
        RECT 18.645 143.505 18.875 143.510 ;
        RECT 12.250 143.310 12.580 143.325 ;
        RECT 12.235 143.050 12.595 143.310 ;
        RECT 12.250 143.025 12.580 143.050 ;
        RECT 12.810 142.765 12.980 143.465 ;
        RECT 13.210 143.310 13.540 143.325 ;
        RECT 13.190 143.050 13.550 143.310 ;
        RECT 13.210 143.025 13.540 143.050 ;
        RECT 13.770 142.765 13.940 143.465 ;
        RECT 14.170 143.310 14.500 143.325 ;
        RECT 14.150 143.050 14.510 143.310 ;
        RECT 14.170 143.025 14.500 143.050 ;
        RECT 14.730 142.765 14.900 143.465 ;
        RECT 15.130 143.310 15.460 143.325 ;
        RECT 15.110 143.050 15.470 143.310 ;
        RECT 15.130 143.025 15.460 143.050 ;
        RECT 15.690 142.765 15.860 143.465 ;
        RECT 16.090 143.305 16.420 143.325 ;
        RECT 16.075 143.045 16.435 143.305 ;
        RECT 16.090 143.025 16.420 143.045 ;
        RECT 16.650 142.765 16.820 143.465 ;
        RECT 17.050 143.305 17.380 143.325 ;
        RECT 17.035 143.045 17.395 143.305 ;
        RECT 17.050 143.025 17.380 143.045 ;
        RECT 11.410 142.595 16.820 142.765 ;
        RECT 19.015 142.765 19.185 143.510 ;
        RECT 20.385 143.465 20.615 143.985 ;
        RECT 21.345 143.465 21.575 143.985 ;
        RECT 22.305 143.465 22.535 143.985 ;
        RECT 23.265 143.465 23.495 143.985 ;
        RECT 24.225 143.465 24.455 143.985 ;
        RECT 19.855 143.310 20.185 143.325 ;
        RECT 19.840 143.050 20.200 143.310 ;
        RECT 19.855 143.025 20.185 143.050 ;
        RECT 20.415 142.765 20.585 143.465 ;
        RECT 20.815 143.310 21.145 143.325 ;
        RECT 20.795 143.050 21.155 143.310 ;
        RECT 20.815 143.025 21.145 143.050 ;
        RECT 21.375 142.765 21.545 143.465 ;
        RECT 21.775 143.310 22.105 143.325 ;
        RECT 21.755 143.050 22.115 143.310 ;
        RECT 21.775 143.025 22.105 143.050 ;
        RECT 22.335 142.765 22.505 143.465 ;
        RECT 22.735 143.310 23.065 143.325 ;
        RECT 22.715 143.050 23.075 143.310 ;
        RECT 22.735 143.025 23.065 143.050 ;
        RECT 23.295 142.765 23.465 143.465 ;
        RECT 23.695 143.305 24.025 143.325 ;
        RECT 23.680 143.045 24.040 143.305 ;
        RECT 23.695 143.025 24.025 143.045 ;
        RECT 24.255 142.765 24.425 143.465 ;
        RECT 24.655 143.305 24.985 143.325 ;
        RECT 24.640 143.045 25.000 143.305 ;
        RECT 24.655 143.025 24.985 143.045 ;
        RECT 19.015 142.595 24.425 142.765 ;
        RECT 11.410 141.200 16.820 141.370 ;
        RECT 1.535 139.070 1.765 140.430 ;
        RECT 2.495 139.070 2.725 140.430 ;
        RECT 3.455 139.070 3.685 140.430 ;
        RECT 4.415 139.070 4.645 140.430 ;
        RECT 5.375 139.070 5.605 140.430 ;
        RECT 6.335 139.070 6.565 140.430 ;
        RECT 1.565 138.365 1.735 139.070 ;
        RECT 2.525 138.365 2.695 139.070 ;
        RECT 3.485 138.365 3.655 139.070 ;
        RECT 4.445 138.365 4.615 139.070 ;
        RECT 5.405 138.365 5.575 139.070 ;
        RECT 6.365 138.365 6.535 139.070 ;
        RECT 11.410 138.385 11.580 141.200 ;
        RECT 12.810 140.450 12.980 141.200 ;
        RECT 13.770 140.450 13.940 141.200 ;
        RECT 14.730 140.450 14.900 141.200 ;
        RECT 15.690 140.450 15.860 141.200 ;
        RECT 16.650 140.450 16.820 141.200 ;
        RECT 19.015 141.200 24.425 141.370 ;
        RECT 12.300 139.090 12.530 140.450 ;
        RECT 12.780 139.090 13.010 140.450 ;
        RECT 13.260 139.090 13.490 140.450 ;
        RECT 13.740 139.090 13.970 140.450 ;
        RECT 14.220 139.090 14.450 140.450 ;
        RECT 14.700 139.090 14.930 140.450 ;
        RECT 15.180 139.090 15.410 140.450 ;
        RECT 15.660 139.090 15.890 140.450 ;
        RECT 16.140 139.090 16.370 140.450 ;
        RECT 16.620 139.090 16.850 140.450 ;
        RECT 17.100 139.090 17.330 140.450 ;
        RECT 10.505 138.365 11.580 138.385 ;
        RECT 1.565 138.215 11.580 138.365 ;
        RECT 1.565 138.195 10.705 138.215 ;
        RECT 1.565 137.530 1.735 138.195 ;
        RECT 2.525 137.530 2.695 138.195 ;
        RECT 3.485 137.530 3.655 138.195 ;
        RECT 4.445 137.530 4.615 138.195 ;
        RECT 5.405 137.530 5.575 138.195 ;
        RECT 6.365 137.530 6.535 138.195 ;
        RECT 1.535 137.010 1.765 137.530 ;
        RECT 2.495 137.010 2.725 137.530 ;
        RECT 3.455 137.010 3.685 137.530 ;
        RECT 4.415 137.010 4.645 137.530 ;
        RECT 5.375 137.010 5.605 137.530 ;
        RECT 6.335 137.010 6.565 137.530 ;
        RECT 11.410 136.330 11.580 138.215 ;
        RECT 12.330 138.385 12.500 139.090 ;
        RECT 13.290 138.385 13.460 139.090 ;
        RECT 14.250 138.385 14.420 139.090 ;
        RECT 15.210 138.385 15.380 139.090 ;
        RECT 16.170 138.385 16.340 139.090 ;
        RECT 17.130 138.385 17.300 139.090 ;
        RECT 19.015 138.385 19.185 141.200 ;
        RECT 20.415 140.450 20.585 141.200 ;
        RECT 21.375 140.450 21.545 141.200 ;
        RECT 22.335 140.450 22.505 141.200 ;
        RECT 23.295 140.450 23.465 141.200 ;
        RECT 24.255 140.450 24.425 141.200 ;
        RECT 20.385 139.090 20.615 140.450 ;
        RECT 21.345 139.090 21.575 140.450 ;
        RECT 22.305 139.090 22.535 140.450 ;
        RECT 23.265 139.090 23.495 140.450 ;
        RECT 24.225 139.090 24.455 140.450 ;
        RECT 12.330 138.215 19.185 138.385 ;
        RECT 12.330 137.550 12.500 138.215 ;
        RECT 13.290 137.550 13.460 138.215 ;
        RECT 14.250 137.550 14.420 138.215 ;
        RECT 15.210 137.550 15.380 138.215 ;
        RECT 16.170 137.550 16.340 138.215 ;
        RECT 17.130 137.550 17.300 138.215 ;
        RECT 19.015 137.575 19.185 138.215 ;
        RECT 26.630 137.920 27.000 138.190 ;
        RECT 18.670 137.570 19.185 137.575 ;
        RECT 12.300 137.030 12.530 137.550 ;
        RECT 12.780 137.030 13.010 137.550 ;
        RECT 13.260 137.030 13.490 137.550 ;
        RECT 13.740 137.030 13.970 137.550 ;
        RECT 14.220 137.030 14.450 137.550 ;
        RECT 14.700 137.030 14.930 137.550 ;
        RECT 15.180 137.030 15.410 137.550 ;
        RECT 15.660 137.030 15.890 137.550 ;
        RECT 16.140 137.030 16.370 137.550 ;
        RECT 16.620 137.030 16.850 137.550 ;
        RECT 17.100 137.030 17.330 137.550 ;
        RECT 18.645 137.075 19.185 137.570 ;
        RECT 18.645 137.070 18.875 137.075 ;
        RECT 12.250 136.875 12.580 136.890 ;
        RECT 12.235 136.615 12.595 136.875 ;
        RECT 12.250 136.590 12.580 136.615 ;
        RECT 12.810 136.330 12.980 137.030 ;
        RECT 13.210 136.875 13.540 136.890 ;
        RECT 13.190 136.615 13.550 136.875 ;
        RECT 13.210 136.590 13.540 136.615 ;
        RECT 13.770 136.330 13.940 137.030 ;
        RECT 14.170 136.875 14.500 136.890 ;
        RECT 14.150 136.615 14.510 136.875 ;
        RECT 14.170 136.590 14.500 136.615 ;
        RECT 14.730 136.330 14.900 137.030 ;
        RECT 15.130 136.875 15.460 136.890 ;
        RECT 15.110 136.615 15.470 136.875 ;
        RECT 15.130 136.590 15.460 136.615 ;
        RECT 15.690 136.330 15.860 137.030 ;
        RECT 16.090 136.870 16.420 136.890 ;
        RECT 16.075 136.610 16.435 136.870 ;
        RECT 16.090 136.590 16.420 136.610 ;
        RECT 16.650 136.330 16.820 137.030 ;
        RECT 17.050 136.870 17.380 136.890 ;
        RECT 17.035 136.610 17.395 136.870 ;
        RECT 17.050 136.590 17.380 136.610 ;
        RECT 11.410 136.160 16.820 136.330 ;
        RECT 19.015 136.330 19.185 137.075 ;
        RECT 20.385 137.030 20.615 137.550 ;
        RECT 21.345 137.030 21.575 137.550 ;
        RECT 22.305 137.030 22.535 137.550 ;
        RECT 23.265 137.030 23.495 137.550 ;
        RECT 24.225 137.030 24.455 137.550 ;
        RECT 19.855 136.875 20.185 136.890 ;
        RECT 19.840 136.615 20.200 136.875 ;
        RECT 19.855 136.590 20.185 136.615 ;
        RECT 20.415 136.330 20.585 137.030 ;
        RECT 20.815 136.875 21.145 136.890 ;
        RECT 20.795 136.615 21.155 136.875 ;
        RECT 20.815 136.590 21.145 136.615 ;
        RECT 21.375 136.330 21.545 137.030 ;
        RECT 21.775 136.875 22.105 136.890 ;
        RECT 21.755 136.615 22.115 136.875 ;
        RECT 21.775 136.590 22.105 136.615 ;
        RECT 22.335 136.330 22.505 137.030 ;
        RECT 22.735 136.875 23.065 136.890 ;
        RECT 22.715 136.615 23.075 136.875 ;
        RECT 22.735 136.590 23.065 136.615 ;
        RECT 23.295 136.330 23.465 137.030 ;
        RECT 23.695 136.870 24.025 136.890 ;
        RECT 23.680 136.610 24.040 136.870 ;
        RECT 23.695 136.590 24.025 136.610 ;
        RECT 24.255 136.330 24.425 137.030 ;
        RECT 24.655 136.870 24.985 136.890 ;
        RECT 24.640 136.610 25.000 136.870 ;
        RECT 24.655 136.590 24.985 136.610 ;
        RECT 19.015 136.160 24.425 136.330 ;
        RECT 11.410 134.765 16.820 134.935 ;
        RECT 1.535 132.635 1.765 133.995 ;
        RECT 2.495 132.635 2.725 133.995 ;
        RECT 3.455 132.635 3.685 133.995 ;
        RECT 4.415 132.635 4.645 133.995 ;
        RECT 5.375 132.635 5.605 133.995 ;
        RECT 6.335 132.635 6.565 133.995 ;
        RECT 1.565 131.930 1.735 132.635 ;
        RECT 2.525 131.930 2.695 132.635 ;
        RECT 3.485 131.930 3.655 132.635 ;
        RECT 4.445 131.930 4.615 132.635 ;
        RECT 5.405 131.930 5.575 132.635 ;
        RECT 6.365 131.930 6.535 132.635 ;
        RECT 11.410 131.950 11.580 134.765 ;
        RECT 12.810 134.015 12.980 134.765 ;
        RECT 13.770 134.015 13.940 134.765 ;
        RECT 14.730 134.015 14.900 134.765 ;
        RECT 15.690 134.015 15.860 134.765 ;
        RECT 16.650 134.015 16.820 134.765 ;
        RECT 19.015 134.765 24.425 134.935 ;
        RECT 12.300 132.655 12.530 134.015 ;
        RECT 12.780 132.655 13.010 134.015 ;
        RECT 13.260 132.655 13.490 134.015 ;
        RECT 13.740 132.655 13.970 134.015 ;
        RECT 14.220 132.655 14.450 134.015 ;
        RECT 14.700 132.655 14.930 134.015 ;
        RECT 15.180 132.655 15.410 134.015 ;
        RECT 15.660 132.655 15.890 134.015 ;
        RECT 16.140 132.655 16.370 134.015 ;
        RECT 16.620 132.655 16.850 134.015 ;
        RECT 17.100 132.655 17.330 134.015 ;
        RECT 10.505 131.930 11.580 131.950 ;
        RECT 1.565 131.780 11.580 131.930 ;
        RECT 1.565 131.760 10.705 131.780 ;
        RECT 1.565 131.095 1.735 131.760 ;
        RECT 2.525 131.095 2.695 131.760 ;
        RECT 3.485 131.095 3.655 131.760 ;
        RECT 4.445 131.095 4.615 131.760 ;
        RECT 5.405 131.095 5.575 131.760 ;
        RECT 6.365 131.095 6.535 131.760 ;
        RECT 1.535 130.575 1.765 131.095 ;
        RECT 2.495 130.575 2.725 131.095 ;
        RECT 3.455 130.575 3.685 131.095 ;
        RECT 4.415 130.575 4.645 131.095 ;
        RECT 5.375 130.575 5.605 131.095 ;
        RECT 6.335 130.575 6.565 131.095 ;
        RECT 11.410 129.895 11.580 131.780 ;
        RECT 12.330 131.950 12.500 132.655 ;
        RECT 13.290 131.950 13.460 132.655 ;
        RECT 14.250 131.950 14.420 132.655 ;
        RECT 15.210 131.950 15.380 132.655 ;
        RECT 16.170 131.950 16.340 132.655 ;
        RECT 17.130 131.950 17.300 132.655 ;
        RECT 19.015 131.950 19.185 134.765 ;
        RECT 20.415 134.015 20.585 134.765 ;
        RECT 21.375 134.015 21.545 134.765 ;
        RECT 22.335 134.015 22.505 134.765 ;
        RECT 23.295 134.015 23.465 134.765 ;
        RECT 24.255 134.015 24.425 134.765 ;
        RECT 20.385 132.655 20.615 134.015 ;
        RECT 21.345 132.655 21.575 134.015 ;
        RECT 22.305 132.655 22.535 134.015 ;
        RECT 23.265 132.655 23.495 134.015 ;
        RECT 24.225 132.655 24.455 134.015 ;
        RECT 12.330 131.780 19.185 131.950 ;
        RECT 12.330 131.115 12.500 131.780 ;
        RECT 13.290 131.115 13.460 131.780 ;
        RECT 14.250 131.115 14.420 131.780 ;
        RECT 15.210 131.115 15.380 131.780 ;
        RECT 16.170 131.115 16.340 131.780 ;
        RECT 17.130 131.115 17.300 131.780 ;
        RECT 19.015 131.140 19.185 131.780 ;
        RECT 26.630 131.485 27.000 131.755 ;
        RECT 18.670 131.135 19.185 131.140 ;
        RECT 12.300 130.595 12.530 131.115 ;
        RECT 12.780 130.595 13.010 131.115 ;
        RECT 13.260 130.595 13.490 131.115 ;
        RECT 13.740 130.595 13.970 131.115 ;
        RECT 14.220 130.595 14.450 131.115 ;
        RECT 14.700 130.595 14.930 131.115 ;
        RECT 15.180 130.595 15.410 131.115 ;
        RECT 15.660 130.595 15.890 131.115 ;
        RECT 16.140 130.595 16.370 131.115 ;
        RECT 16.620 130.595 16.850 131.115 ;
        RECT 17.100 130.595 17.330 131.115 ;
        RECT 18.645 130.640 19.185 131.135 ;
        RECT 18.645 130.635 18.875 130.640 ;
        RECT 12.250 130.440 12.580 130.455 ;
        RECT 12.235 130.180 12.595 130.440 ;
        RECT 12.250 130.155 12.580 130.180 ;
        RECT 12.810 129.895 12.980 130.595 ;
        RECT 13.210 130.440 13.540 130.455 ;
        RECT 13.190 130.180 13.550 130.440 ;
        RECT 13.210 130.155 13.540 130.180 ;
        RECT 13.770 129.895 13.940 130.595 ;
        RECT 14.170 130.440 14.500 130.455 ;
        RECT 14.150 130.180 14.510 130.440 ;
        RECT 14.170 130.155 14.500 130.180 ;
        RECT 14.730 129.895 14.900 130.595 ;
        RECT 15.130 130.440 15.460 130.455 ;
        RECT 15.110 130.180 15.470 130.440 ;
        RECT 15.130 130.155 15.460 130.180 ;
        RECT 15.690 129.895 15.860 130.595 ;
        RECT 16.090 130.435 16.420 130.455 ;
        RECT 16.075 130.175 16.435 130.435 ;
        RECT 16.090 130.155 16.420 130.175 ;
        RECT 16.650 129.895 16.820 130.595 ;
        RECT 17.050 130.435 17.380 130.455 ;
        RECT 17.035 130.175 17.395 130.435 ;
        RECT 17.050 130.155 17.380 130.175 ;
        RECT 11.410 129.725 16.820 129.895 ;
        RECT 19.015 129.895 19.185 130.640 ;
        RECT 20.385 130.595 20.615 131.115 ;
        RECT 21.345 130.595 21.575 131.115 ;
        RECT 22.305 130.595 22.535 131.115 ;
        RECT 23.265 130.595 23.495 131.115 ;
        RECT 24.225 130.595 24.455 131.115 ;
        RECT 19.855 130.440 20.185 130.455 ;
        RECT 19.840 130.180 20.200 130.440 ;
        RECT 19.855 130.155 20.185 130.180 ;
        RECT 20.415 129.895 20.585 130.595 ;
        RECT 20.815 130.440 21.145 130.455 ;
        RECT 20.795 130.180 21.155 130.440 ;
        RECT 20.815 130.155 21.145 130.180 ;
        RECT 21.375 129.895 21.545 130.595 ;
        RECT 21.775 130.440 22.105 130.455 ;
        RECT 21.755 130.180 22.115 130.440 ;
        RECT 21.775 130.155 22.105 130.180 ;
        RECT 22.335 129.895 22.505 130.595 ;
        RECT 22.735 130.440 23.065 130.455 ;
        RECT 22.715 130.180 23.075 130.440 ;
        RECT 22.735 130.155 23.065 130.180 ;
        RECT 23.295 129.895 23.465 130.595 ;
        RECT 23.695 130.435 24.025 130.455 ;
        RECT 23.680 130.175 24.040 130.435 ;
        RECT 23.695 130.155 24.025 130.175 ;
        RECT 24.255 129.895 24.425 130.595 ;
        RECT 24.655 130.435 24.985 130.455 ;
        RECT 24.640 130.175 25.000 130.435 ;
        RECT 24.655 130.155 24.985 130.175 ;
        RECT 19.015 129.725 24.425 129.895 ;
        RECT 11.410 128.330 16.820 128.500 ;
        RECT 1.535 126.200 1.765 127.560 ;
        RECT 2.495 126.200 2.725 127.560 ;
        RECT 3.455 126.200 3.685 127.560 ;
        RECT 4.415 126.200 4.645 127.560 ;
        RECT 5.375 126.200 5.605 127.560 ;
        RECT 6.335 126.200 6.565 127.560 ;
        RECT 1.565 125.495 1.735 126.200 ;
        RECT 2.525 125.495 2.695 126.200 ;
        RECT 3.485 125.495 3.655 126.200 ;
        RECT 4.445 125.495 4.615 126.200 ;
        RECT 5.405 125.495 5.575 126.200 ;
        RECT 6.365 125.495 6.535 126.200 ;
        RECT 11.410 125.515 11.580 128.330 ;
        RECT 12.810 127.580 12.980 128.330 ;
        RECT 13.770 127.580 13.940 128.330 ;
        RECT 14.730 127.580 14.900 128.330 ;
        RECT 15.690 127.580 15.860 128.330 ;
        RECT 16.650 127.580 16.820 128.330 ;
        RECT 19.015 128.330 24.425 128.500 ;
        RECT 12.300 126.220 12.530 127.580 ;
        RECT 12.780 126.220 13.010 127.580 ;
        RECT 13.260 126.220 13.490 127.580 ;
        RECT 13.740 126.220 13.970 127.580 ;
        RECT 14.220 126.220 14.450 127.580 ;
        RECT 14.700 126.220 14.930 127.580 ;
        RECT 15.180 126.220 15.410 127.580 ;
        RECT 15.660 126.220 15.890 127.580 ;
        RECT 16.140 126.220 16.370 127.580 ;
        RECT 16.620 126.220 16.850 127.580 ;
        RECT 17.100 126.220 17.330 127.580 ;
        RECT 10.505 125.495 11.580 125.515 ;
        RECT 1.565 125.345 11.580 125.495 ;
        RECT 1.565 125.325 10.705 125.345 ;
        RECT 1.565 124.660 1.735 125.325 ;
        RECT 2.525 124.660 2.695 125.325 ;
        RECT 3.485 124.660 3.655 125.325 ;
        RECT 4.445 124.660 4.615 125.325 ;
        RECT 5.405 124.660 5.575 125.325 ;
        RECT 6.365 124.660 6.535 125.325 ;
        RECT 1.535 124.140 1.765 124.660 ;
        RECT 2.495 124.140 2.725 124.660 ;
        RECT 3.455 124.140 3.685 124.660 ;
        RECT 4.415 124.140 4.645 124.660 ;
        RECT 5.375 124.140 5.605 124.660 ;
        RECT 6.335 124.140 6.565 124.660 ;
        RECT 11.410 123.460 11.580 125.345 ;
        RECT 12.330 125.515 12.500 126.220 ;
        RECT 13.290 125.515 13.460 126.220 ;
        RECT 14.250 125.515 14.420 126.220 ;
        RECT 15.210 125.515 15.380 126.220 ;
        RECT 16.170 125.515 16.340 126.220 ;
        RECT 17.130 125.515 17.300 126.220 ;
        RECT 19.015 125.515 19.185 128.330 ;
        RECT 20.415 127.580 20.585 128.330 ;
        RECT 21.375 127.580 21.545 128.330 ;
        RECT 22.335 127.580 22.505 128.330 ;
        RECT 23.295 127.580 23.465 128.330 ;
        RECT 24.255 127.580 24.425 128.330 ;
        RECT 20.385 126.220 20.615 127.580 ;
        RECT 21.345 126.220 21.575 127.580 ;
        RECT 22.305 126.220 22.535 127.580 ;
        RECT 23.265 126.220 23.495 127.580 ;
        RECT 24.225 126.220 24.455 127.580 ;
        RECT 12.330 125.345 19.185 125.515 ;
        RECT 12.330 124.680 12.500 125.345 ;
        RECT 13.290 124.680 13.460 125.345 ;
        RECT 14.250 124.680 14.420 125.345 ;
        RECT 15.210 124.680 15.380 125.345 ;
        RECT 16.170 124.680 16.340 125.345 ;
        RECT 17.130 124.680 17.300 125.345 ;
        RECT 19.015 124.705 19.185 125.345 ;
        RECT 26.630 125.050 27.000 125.320 ;
        RECT 18.670 124.700 19.185 124.705 ;
        RECT 12.300 124.160 12.530 124.680 ;
        RECT 12.780 124.160 13.010 124.680 ;
        RECT 13.260 124.160 13.490 124.680 ;
        RECT 13.740 124.160 13.970 124.680 ;
        RECT 14.220 124.160 14.450 124.680 ;
        RECT 14.700 124.160 14.930 124.680 ;
        RECT 15.180 124.160 15.410 124.680 ;
        RECT 15.660 124.160 15.890 124.680 ;
        RECT 16.140 124.160 16.370 124.680 ;
        RECT 16.620 124.160 16.850 124.680 ;
        RECT 17.100 124.160 17.330 124.680 ;
        RECT 18.645 124.205 19.185 124.700 ;
        RECT 18.645 124.200 18.875 124.205 ;
        RECT 12.250 124.005 12.580 124.020 ;
        RECT 12.235 123.745 12.595 124.005 ;
        RECT 12.250 123.720 12.580 123.745 ;
        RECT 12.810 123.460 12.980 124.160 ;
        RECT 13.210 124.005 13.540 124.020 ;
        RECT 13.190 123.745 13.550 124.005 ;
        RECT 13.210 123.720 13.540 123.745 ;
        RECT 13.770 123.460 13.940 124.160 ;
        RECT 14.170 124.005 14.500 124.020 ;
        RECT 14.150 123.745 14.510 124.005 ;
        RECT 14.170 123.720 14.500 123.745 ;
        RECT 14.730 123.460 14.900 124.160 ;
        RECT 15.130 124.005 15.460 124.020 ;
        RECT 15.110 123.745 15.470 124.005 ;
        RECT 15.130 123.720 15.460 123.745 ;
        RECT 15.690 123.460 15.860 124.160 ;
        RECT 16.090 124.000 16.420 124.020 ;
        RECT 16.075 123.740 16.435 124.000 ;
        RECT 16.090 123.720 16.420 123.740 ;
        RECT 16.650 123.460 16.820 124.160 ;
        RECT 17.050 124.000 17.380 124.020 ;
        RECT 17.035 123.740 17.395 124.000 ;
        RECT 17.050 123.720 17.380 123.740 ;
        RECT 11.410 123.290 16.820 123.460 ;
        RECT 19.015 123.460 19.185 124.205 ;
        RECT 20.385 124.160 20.615 124.680 ;
        RECT 21.345 124.160 21.575 124.680 ;
        RECT 22.305 124.160 22.535 124.680 ;
        RECT 23.265 124.160 23.495 124.680 ;
        RECT 24.225 124.160 24.455 124.680 ;
        RECT 19.855 124.005 20.185 124.020 ;
        RECT 19.840 123.745 20.200 124.005 ;
        RECT 19.855 123.720 20.185 123.745 ;
        RECT 20.415 123.460 20.585 124.160 ;
        RECT 20.815 124.005 21.145 124.020 ;
        RECT 20.795 123.745 21.155 124.005 ;
        RECT 20.815 123.720 21.145 123.745 ;
        RECT 21.375 123.460 21.545 124.160 ;
        RECT 21.775 124.005 22.105 124.020 ;
        RECT 21.755 123.745 22.115 124.005 ;
        RECT 21.775 123.720 22.105 123.745 ;
        RECT 22.335 123.460 22.505 124.160 ;
        RECT 22.735 124.005 23.065 124.020 ;
        RECT 22.715 123.745 23.075 124.005 ;
        RECT 22.735 123.720 23.065 123.745 ;
        RECT 23.295 123.460 23.465 124.160 ;
        RECT 23.695 124.000 24.025 124.020 ;
        RECT 23.680 123.740 24.040 124.000 ;
        RECT 23.695 123.720 24.025 123.740 ;
        RECT 24.255 123.460 24.425 124.160 ;
        RECT 24.655 124.000 24.985 124.020 ;
        RECT 24.640 123.740 25.000 124.000 ;
        RECT 24.655 123.720 24.985 123.740 ;
        RECT 19.015 123.290 24.425 123.460 ;
        RECT 11.410 121.895 16.820 122.065 ;
        RECT 1.535 119.765 1.765 121.125 ;
        RECT 2.495 119.765 2.725 121.125 ;
        RECT 3.455 119.765 3.685 121.125 ;
        RECT 4.415 119.765 4.645 121.125 ;
        RECT 5.375 119.765 5.605 121.125 ;
        RECT 6.335 119.765 6.565 121.125 ;
        RECT 1.565 119.060 1.735 119.765 ;
        RECT 2.525 119.060 2.695 119.765 ;
        RECT 3.485 119.060 3.655 119.765 ;
        RECT 4.445 119.060 4.615 119.765 ;
        RECT 5.405 119.060 5.575 119.765 ;
        RECT 6.365 119.060 6.535 119.765 ;
        RECT 11.410 119.080 11.580 121.895 ;
        RECT 12.810 121.145 12.980 121.895 ;
        RECT 13.770 121.145 13.940 121.895 ;
        RECT 14.730 121.145 14.900 121.895 ;
        RECT 15.690 121.145 15.860 121.895 ;
        RECT 16.650 121.145 16.820 121.895 ;
        RECT 19.015 121.895 24.425 122.065 ;
        RECT 12.300 119.785 12.530 121.145 ;
        RECT 12.780 119.785 13.010 121.145 ;
        RECT 13.260 119.785 13.490 121.145 ;
        RECT 13.740 119.785 13.970 121.145 ;
        RECT 14.220 119.785 14.450 121.145 ;
        RECT 14.700 119.785 14.930 121.145 ;
        RECT 15.180 119.785 15.410 121.145 ;
        RECT 15.660 119.785 15.890 121.145 ;
        RECT 16.140 119.785 16.370 121.145 ;
        RECT 16.620 119.785 16.850 121.145 ;
        RECT 17.100 119.785 17.330 121.145 ;
        RECT 10.505 119.060 11.580 119.080 ;
        RECT 1.565 118.910 11.580 119.060 ;
        RECT 1.565 118.890 10.705 118.910 ;
        RECT 1.565 118.225 1.735 118.890 ;
        RECT 2.525 118.225 2.695 118.890 ;
        RECT 3.485 118.225 3.655 118.890 ;
        RECT 4.445 118.225 4.615 118.890 ;
        RECT 5.405 118.225 5.575 118.890 ;
        RECT 6.365 118.225 6.535 118.890 ;
        RECT 1.535 117.705 1.765 118.225 ;
        RECT 2.495 117.705 2.725 118.225 ;
        RECT 3.455 117.705 3.685 118.225 ;
        RECT 4.415 117.705 4.645 118.225 ;
        RECT 5.375 117.705 5.605 118.225 ;
        RECT 6.335 117.705 6.565 118.225 ;
        RECT 11.410 117.025 11.580 118.910 ;
        RECT 12.330 119.080 12.500 119.785 ;
        RECT 13.290 119.080 13.460 119.785 ;
        RECT 14.250 119.080 14.420 119.785 ;
        RECT 15.210 119.080 15.380 119.785 ;
        RECT 16.170 119.080 16.340 119.785 ;
        RECT 17.130 119.080 17.300 119.785 ;
        RECT 19.015 119.080 19.185 121.895 ;
        RECT 20.415 121.145 20.585 121.895 ;
        RECT 21.375 121.145 21.545 121.895 ;
        RECT 22.335 121.145 22.505 121.895 ;
        RECT 23.295 121.145 23.465 121.895 ;
        RECT 24.255 121.145 24.425 121.895 ;
        RECT 20.385 119.785 20.615 121.145 ;
        RECT 21.345 119.785 21.575 121.145 ;
        RECT 22.305 119.785 22.535 121.145 ;
        RECT 23.265 119.785 23.495 121.145 ;
        RECT 24.225 119.785 24.455 121.145 ;
        RECT 12.330 118.910 19.185 119.080 ;
        RECT 12.330 118.245 12.500 118.910 ;
        RECT 13.290 118.245 13.460 118.910 ;
        RECT 14.250 118.245 14.420 118.910 ;
        RECT 15.210 118.245 15.380 118.910 ;
        RECT 16.170 118.245 16.340 118.910 ;
        RECT 17.130 118.245 17.300 118.910 ;
        RECT 19.015 118.270 19.185 118.910 ;
        RECT 26.630 118.615 27.000 118.885 ;
        RECT 18.670 118.265 19.185 118.270 ;
        RECT 12.300 117.725 12.530 118.245 ;
        RECT 12.780 117.725 13.010 118.245 ;
        RECT 13.260 117.725 13.490 118.245 ;
        RECT 13.740 117.725 13.970 118.245 ;
        RECT 14.220 117.725 14.450 118.245 ;
        RECT 14.700 117.725 14.930 118.245 ;
        RECT 15.180 117.725 15.410 118.245 ;
        RECT 15.660 117.725 15.890 118.245 ;
        RECT 16.140 117.725 16.370 118.245 ;
        RECT 16.620 117.725 16.850 118.245 ;
        RECT 17.100 117.725 17.330 118.245 ;
        RECT 18.645 117.770 19.185 118.265 ;
        RECT 18.645 117.765 18.875 117.770 ;
        RECT 12.250 117.570 12.580 117.585 ;
        RECT 12.235 117.310 12.595 117.570 ;
        RECT 12.250 117.285 12.580 117.310 ;
        RECT 12.810 117.025 12.980 117.725 ;
        RECT 13.210 117.570 13.540 117.585 ;
        RECT 13.190 117.310 13.550 117.570 ;
        RECT 13.210 117.285 13.540 117.310 ;
        RECT 13.770 117.025 13.940 117.725 ;
        RECT 14.170 117.570 14.500 117.585 ;
        RECT 14.150 117.310 14.510 117.570 ;
        RECT 14.170 117.285 14.500 117.310 ;
        RECT 14.730 117.025 14.900 117.725 ;
        RECT 15.130 117.570 15.460 117.585 ;
        RECT 15.110 117.310 15.470 117.570 ;
        RECT 15.130 117.285 15.460 117.310 ;
        RECT 15.690 117.025 15.860 117.725 ;
        RECT 16.090 117.565 16.420 117.585 ;
        RECT 16.075 117.305 16.435 117.565 ;
        RECT 16.090 117.285 16.420 117.305 ;
        RECT 16.650 117.025 16.820 117.725 ;
        RECT 17.050 117.565 17.380 117.585 ;
        RECT 17.035 117.305 17.395 117.565 ;
        RECT 17.050 117.285 17.380 117.305 ;
        RECT 11.410 116.855 16.820 117.025 ;
        RECT 19.015 117.025 19.185 117.770 ;
        RECT 20.385 117.725 20.615 118.245 ;
        RECT 21.345 117.725 21.575 118.245 ;
        RECT 22.305 117.725 22.535 118.245 ;
        RECT 23.265 117.725 23.495 118.245 ;
        RECT 24.225 117.725 24.455 118.245 ;
        RECT 19.855 117.570 20.185 117.585 ;
        RECT 19.840 117.310 20.200 117.570 ;
        RECT 19.855 117.285 20.185 117.310 ;
        RECT 20.415 117.025 20.585 117.725 ;
        RECT 20.815 117.570 21.145 117.585 ;
        RECT 20.795 117.310 21.155 117.570 ;
        RECT 20.815 117.285 21.145 117.310 ;
        RECT 21.375 117.025 21.545 117.725 ;
        RECT 21.775 117.570 22.105 117.585 ;
        RECT 21.755 117.310 22.115 117.570 ;
        RECT 21.775 117.285 22.105 117.310 ;
        RECT 22.335 117.025 22.505 117.725 ;
        RECT 22.735 117.570 23.065 117.585 ;
        RECT 22.715 117.310 23.075 117.570 ;
        RECT 22.735 117.285 23.065 117.310 ;
        RECT 23.295 117.025 23.465 117.725 ;
        RECT 23.695 117.565 24.025 117.585 ;
        RECT 23.680 117.305 24.040 117.565 ;
        RECT 23.695 117.285 24.025 117.305 ;
        RECT 24.255 117.025 24.425 117.725 ;
        RECT 24.655 117.565 24.985 117.585 ;
        RECT 24.640 117.305 25.000 117.565 ;
        RECT 24.655 117.285 24.985 117.305 ;
        RECT 19.015 116.855 24.425 117.025 ;
        RECT 11.410 115.460 16.820 115.630 ;
        RECT 1.535 113.330 1.765 114.690 ;
        RECT 2.495 113.330 2.725 114.690 ;
        RECT 3.455 113.330 3.685 114.690 ;
        RECT 4.415 113.330 4.645 114.690 ;
        RECT 5.375 113.330 5.605 114.690 ;
        RECT 6.335 113.330 6.565 114.690 ;
        RECT 1.565 112.625 1.735 113.330 ;
        RECT 2.525 112.625 2.695 113.330 ;
        RECT 3.485 112.625 3.655 113.330 ;
        RECT 4.445 112.625 4.615 113.330 ;
        RECT 5.405 112.625 5.575 113.330 ;
        RECT 6.365 112.625 6.535 113.330 ;
        RECT 11.410 112.645 11.580 115.460 ;
        RECT 12.810 114.710 12.980 115.460 ;
        RECT 13.770 114.710 13.940 115.460 ;
        RECT 14.730 114.710 14.900 115.460 ;
        RECT 15.690 114.710 15.860 115.460 ;
        RECT 16.650 114.710 16.820 115.460 ;
        RECT 19.015 115.460 24.425 115.630 ;
        RECT 12.300 113.350 12.530 114.710 ;
        RECT 12.780 113.350 13.010 114.710 ;
        RECT 13.260 113.350 13.490 114.710 ;
        RECT 13.740 113.350 13.970 114.710 ;
        RECT 14.220 113.350 14.450 114.710 ;
        RECT 14.700 113.350 14.930 114.710 ;
        RECT 15.180 113.350 15.410 114.710 ;
        RECT 15.660 113.350 15.890 114.710 ;
        RECT 16.140 113.350 16.370 114.710 ;
        RECT 16.620 113.350 16.850 114.710 ;
        RECT 17.100 113.350 17.330 114.710 ;
        RECT 10.505 112.625 11.580 112.645 ;
        RECT 1.565 112.475 11.580 112.625 ;
        RECT 1.565 112.455 10.705 112.475 ;
        RECT 1.565 111.790 1.735 112.455 ;
        RECT 2.525 111.790 2.695 112.455 ;
        RECT 3.485 111.790 3.655 112.455 ;
        RECT 4.445 111.790 4.615 112.455 ;
        RECT 5.405 111.790 5.575 112.455 ;
        RECT 6.365 111.790 6.535 112.455 ;
        RECT 1.535 111.270 1.765 111.790 ;
        RECT 2.495 111.270 2.725 111.790 ;
        RECT 3.455 111.270 3.685 111.790 ;
        RECT 4.415 111.270 4.645 111.790 ;
        RECT 5.375 111.270 5.605 111.790 ;
        RECT 6.335 111.270 6.565 111.790 ;
        RECT 11.410 110.590 11.580 112.475 ;
        RECT 12.330 112.645 12.500 113.350 ;
        RECT 13.290 112.645 13.460 113.350 ;
        RECT 14.250 112.645 14.420 113.350 ;
        RECT 15.210 112.645 15.380 113.350 ;
        RECT 16.170 112.645 16.340 113.350 ;
        RECT 17.130 112.645 17.300 113.350 ;
        RECT 19.015 112.645 19.185 115.460 ;
        RECT 20.415 114.710 20.585 115.460 ;
        RECT 21.375 114.710 21.545 115.460 ;
        RECT 22.335 114.710 22.505 115.460 ;
        RECT 23.295 114.710 23.465 115.460 ;
        RECT 24.255 114.710 24.425 115.460 ;
        RECT 20.385 113.350 20.615 114.710 ;
        RECT 21.345 113.350 21.575 114.710 ;
        RECT 22.305 113.350 22.535 114.710 ;
        RECT 23.265 113.350 23.495 114.710 ;
        RECT 24.225 113.350 24.455 114.710 ;
        RECT 12.330 112.475 19.185 112.645 ;
        RECT 12.330 111.810 12.500 112.475 ;
        RECT 13.290 111.810 13.460 112.475 ;
        RECT 14.250 111.810 14.420 112.475 ;
        RECT 15.210 111.810 15.380 112.475 ;
        RECT 16.170 111.810 16.340 112.475 ;
        RECT 17.130 111.810 17.300 112.475 ;
        RECT 19.015 111.835 19.185 112.475 ;
        RECT 26.630 112.180 27.000 112.450 ;
        RECT 18.670 111.830 19.185 111.835 ;
        RECT 12.300 111.290 12.530 111.810 ;
        RECT 12.780 111.290 13.010 111.810 ;
        RECT 13.260 111.290 13.490 111.810 ;
        RECT 13.740 111.290 13.970 111.810 ;
        RECT 14.220 111.290 14.450 111.810 ;
        RECT 14.700 111.290 14.930 111.810 ;
        RECT 15.180 111.290 15.410 111.810 ;
        RECT 15.660 111.290 15.890 111.810 ;
        RECT 16.140 111.290 16.370 111.810 ;
        RECT 16.620 111.290 16.850 111.810 ;
        RECT 17.100 111.290 17.330 111.810 ;
        RECT 18.645 111.335 19.185 111.830 ;
        RECT 18.645 111.330 18.875 111.335 ;
        RECT 12.250 111.135 12.580 111.150 ;
        RECT 12.235 110.875 12.595 111.135 ;
        RECT 12.250 110.850 12.580 110.875 ;
        RECT 12.810 110.590 12.980 111.290 ;
        RECT 13.210 111.135 13.540 111.150 ;
        RECT 13.190 110.875 13.550 111.135 ;
        RECT 13.210 110.850 13.540 110.875 ;
        RECT 13.770 110.590 13.940 111.290 ;
        RECT 14.170 111.135 14.500 111.150 ;
        RECT 14.150 110.875 14.510 111.135 ;
        RECT 14.170 110.850 14.500 110.875 ;
        RECT 14.730 110.590 14.900 111.290 ;
        RECT 15.130 111.135 15.460 111.150 ;
        RECT 15.110 110.875 15.470 111.135 ;
        RECT 15.130 110.850 15.460 110.875 ;
        RECT 15.690 110.590 15.860 111.290 ;
        RECT 16.090 111.130 16.420 111.150 ;
        RECT 16.075 110.870 16.435 111.130 ;
        RECT 16.090 110.850 16.420 110.870 ;
        RECT 16.650 110.590 16.820 111.290 ;
        RECT 17.050 111.130 17.380 111.150 ;
        RECT 17.035 110.870 17.395 111.130 ;
        RECT 17.050 110.850 17.380 110.870 ;
        RECT 11.410 110.420 16.820 110.590 ;
        RECT 19.015 110.590 19.185 111.335 ;
        RECT 20.385 111.290 20.615 111.810 ;
        RECT 21.345 111.290 21.575 111.810 ;
        RECT 22.305 111.290 22.535 111.810 ;
        RECT 23.265 111.290 23.495 111.810 ;
        RECT 24.225 111.290 24.455 111.810 ;
        RECT 19.855 111.135 20.185 111.150 ;
        RECT 19.840 110.875 20.200 111.135 ;
        RECT 19.855 110.850 20.185 110.875 ;
        RECT 20.415 110.590 20.585 111.290 ;
        RECT 20.815 111.135 21.145 111.150 ;
        RECT 20.795 110.875 21.155 111.135 ;
        RECT 20.815 110.850 21.145 110.875 ;
        RECT 21.375 110.590 21.545 111.290 ;
        RECT 21.775 111.135 22.105 111.150 ;
        RECT 21.755 110.875 22.115 111.135 ;
        RECT 21.775 110.850 22.105 110.875 ;
        RECT 22.335 110.590 22.505 111.290 ;
        RECT 22.735 111.135 23.065 111.150 ;
        RECT 22.715 110.875 23.075 111.135 ;
        RECT 22.735 110.850 23.065 110.875 ;
        RECT 23.295 110.590 23.465 111.290 ;
        RECT 23.695 111.130 24.025 111.150 ;
        RECT 23.680 110.870 24.040 111.130 ;
        RECT 23.695 110.850 24.025 110.870 ;
        RECT 24.255 110.590 24.425 111.290 ;
        RECT 24.655 111.130 24.985 111.150 ;
        RECT 24.640 110.870 25.000 111.130 ;
        RECT 24.655 110.850 24.985 110.870 ;
        RECT 19.015 110.420 24.425 110.590 ;
        RECT 11.410 109.025 16.820 109.195 ;
        RECT 1.535 106.895 1.765 108.255 ;
        RECT 2.495 106.895 2.725 108.255 ;
        RECT 3.455 106.895 3.685 108.255 ;
        RECT 4.415 106.895 4.645 108.255 ;
        RECT 5.375 106.895 5.605 108.255 ;
        RECT 6.335 106.895 6.565 108.255 ;
        RECT 1.565 106.190 1.735 106.895 ;
        RECT 2.525 106.190 2.695 106.895 ;
        RECT 3.485 106.190 3.655 106.895 ;
        RECT 4.445 106.190 4.615 106.895 ;
        RECT 5.405 106.190 5.575 106.895 ;
        RECT 6.365 106.190 6.535 106.895 ;
        RECT 11.410 106.210 11.580 109.025 ;
        RECT 12.810 108.275 12.980 109.025 ;
        RECT 13.770 108.275 13.940 109.025 ;
        RECT 14.730 108.275 14.900 109.025 ;
        RECT 15.690 108.275 15.860 109.025 ;
        RECT 16.650 108.275 16.820 109.025 ;
        RECT 19.015 109.025 24.425 109.195 ;
        RECT 12.300 106.915 12.530 108.275 ;
        RECT 12.780 106.915 13.010 108.275 ;
        RECT 13.260 106.915 13.490 108.275 ;
        RECT 13.740 106.915 13.970 108.275 ;
        RECT 14.220 106.915 14.450 108.275 ;
        RECT 14.700 106.915 14.930 108.275 ;
        RECT 15.180 106.915 15.410 108.275 ;
        RECT 15.660 106.915 15.890 108.275 ;
        RECT 16.140 106.915 16.370 108.275 ;
        RECT 16.620 106.915 16.850 108.275 ;
        RECT 17.100 106.915 17.330 108.275 ;
        RECT 10.505 106.190 11.580 106.210 ;
        RECT 1.565 106.040 11.580 106.190 ;
        RECT 1.565 106.020 10.705 106.040 ;
        RECT 1.565 105.355 1.735 106.020 ;
        RECT 2.525 105.355 2.695 106.020 ;
        RECT 3.485 105.355 3.655 106.020 ;
        RECT 4.445 105.355 4.615 106.020 ;
        RECT 5.405 105.355 5.575 106.020 ;
        RECT 6.365 105.355 6.535 106.020 ;
        RECT 1.535 104.835 1.765 105.355 ;
        RECT 2.495 104.835 2.725 105.355 ;
        RECT 3.455 104.835 3.685 105.355 ;
        RECT 4.415 104.835 4.645 105.355 ;
        RECT 5.375 104.835 5.605 105.355 ;
        RECT 6.335 104.835 6.565 105.355 ;
        RECT 11.410 104.155 11.580 106.040 ;
        RECT 12.330 106.210 12.500 106.915 ;
        RECT 13.290 106.210 13.460 106.915 ;
        RECT 14.250 106.210 14.420 106.915 ;
        RECT 15.210 106.210 15.380 106.915 ;
        RECT 16.170 106.210 16.340 106.915 ;
        RECT 17.130 106.210 17.300 106.915 ;
        RECT 19.015 106.210 19.185 109.025 ;
        RECT 20.415 108.275 20.585 109.025 ;
        RECT 21.375 108.275 21.545 109.025 ;
        RECT 22.335 108.275 22.505 109.025 ;
        RECT 23.295 108.275 23.465 109.025 ;
        RECT 24.255 108.275 24.425 109.025 ;
        RECT 20.385 106.915 20.615 108.275 ;
        RECT 21.345 106.915 21.575 108.275 ;
        RECT 22.305 106.915 22.535 108.275 ;
        RECT 23.265 106.915 23.495 108.275 ;
        RECT 24.225 106.915 24.455 108.275 ;
        RECT 12.330 106.040 19.185 106.210 ;
        RECT 12.330 105.375 12.500 106.040 ;
        RECT 13.290 105.375 13.460 106.040 ;
        RECT 14.250 105.375 14.420 106.040 ;
        RECT 15.210 105.375 15.380 106.040 ;
        RECT 16.170 105.375 16.340 106.040 ;
        RECT 17.130 105.375 17.300 106.040 ;
        RECT 19.015 105.400 19.185 106.040 ;
        RECT 26.630 105.745 27.000 106.015 ;
        RECT 18.670 105.395 19.185 105.400 ;
        RECT 12.300 104.855 12.530 105.375 ;
        RECT 12.780 104.855 13.010 105.375 ;
        RECT 13.260 104.855 13.490 105.375 ;
        RECT 13.740 104.855 13.970 105.375 ;
        RECT 14.220 104.855 14.450 105.375 ;
        RECT 14.700 104.855 14.930 105.375 ;
        RECT 15.180 104.855 15.410 105.375 ;
        RECT 15.660 104.855 15.890 105.375 ;
        RECT 16.140 104.855 16.370 105.375 ;
        RECT 16.620 104.855 16.850 105.375 ;
        RECT 17.100 104.855 17.330 105.375 ;
        RECT 18.645 104.900 19.185 105.395 ;
        RECT 18.645 104.895 18.875 104.900 ;
        RECT 12.250 104.700 12.580 104.715 ;
        RECT 12.235 104.440 12.595 104.700 ;
        RECT 12.250 104.415 12.580 104.440 ;
        RECT 12.810 104.155 12.980 104.855 ;
        RECT 13.210 104.700 13.540 104.715 ;
        RECT 13.190 104.440 13.550 104.700 ;
        RECT 13.210 104.415 13.540 104.440 ;
        RECT 13.770 104.155 13.940 104.855 ;
        RECT 14.170 104.700 14.500 104.715 ;
        RECT 14.150 104.440 14.510 104.700 ;
        RECT 14.170 104.415 14.500 104.440 ;
        RECT 14.730 104.155 14.900 104.855 ;
        RECT 15.130 104.700 15.460 104.715 ;
        RECT 15.110 104.440 15.470 104.700 ;
        RECT 15.130 104.415 15.460 104.440 ;
        RECT 15.690 104.155 15.860 104.855 ;
        RECT 16.090 104.695 16.420 104.715 ;
        RECT 16.075 104.435 16.435 104.695 ;
        RECT 16.090 104.415 16.420 104.435 ;
        RECT 16.650 104.155 16.820 104.855 ;
        RECT 17.050 104.695 17.380 104.715 ;
        RECT 17.035 104.435 17.395 104.695 ;
        RECT 17.050 104.415 17.380 104.435 ;
        RECT 11.410 103.985 16.820 104.155 ;
        RECT 19.015 104.155 19.185 104.900 ;
        RECT 20.385 104.855 20.615 105.375 ;
        RECT 21.345 104.855 21.575 105.375 ;
        RECT 22.305 104.855 22.535 105.375 ;
        RECT 23.265 104.855 23.495 105.375 ;
        RECT 24.225 104.855 24.455 105.375 ;
        RECT 19.855 104.700 20.185 104.715 ;
        RECT 19.840 104.440 20.200 104.700 ;
        RECT 19.855 104.415 20.185 104.440 ;
        RECT 20.415 104.155 20.585 104.855 ;
        RECT 20.815 104.700 21.145 104.715 ;
        RECT 20.795 104.440 21.155 104.700 ;
        RECT 20.815 104.415 21.145 104.440 ;
        RECT 21.375 104.155 21.545 104.855 ;
        RECT 21.775 104.700 22.105 104.715 ;
        RECT 21.755 104.440 22.115 104.700 ;
        RECT 21.775 104.415 22.105 104.440 ;
        RECT 22.335 104.155 22.505 104.855 ;
        RECT 22.735 104.700 23.065 104.715 ;
        RECT 22.715 104.440 23.075 104.700 ;
        RECT 22.735 104.415 23.065 104.440 ;
        RECT 23.295 104.155 23.465 104.855 ;
        RECT 23.695 104.695 24.025 104.715 ;
        RECT 23.680 104.435 24.040 104.695 ;
        RECT 23.695 104.415 24.025 104.435 ;
        RECT 24.255 104.155 24.425 104.855 ;
        RECT 24.655 104.695 24.985 104.715 ;
        RECT 24.640 104.435 25.000 104.695 ;
        RECT 24.655 104.415 24.985 104.435 ;
        RECT 19.015 103.985 24.425 104.155 ;
        RECT 11.410 102.590 16.820 102.760 ;
        RECT 1.535 100.460 1.765 101.820 ;
        RECT 2.495 100.460 2.725 101.820 ;
        RECT 3.455 100.460 3.685 101.820 ;
        RECT 4.415 100.460 4.645 101.820 ;
        RECT 5.375 100.460 5.605 101.820 ;
        RECT 6.335 100.460 6.565 101.820 ;
        RECT 1.565 99.755 1.735 100.460 ;
        RECT 2.525 99.755 2.695 100.460 ;
        RECT 3.485 99.755 3.655 100.460 ;
        RECT 4.445 99.755 4.615 100.460 ;
        RECT 5.405 99.755 5.575 100.460 ;
        RECT 6.365 99.755 6.535 100.460 ;
        RECT 11.410 99.775 11.580 102.590 ;
        RECT 12.810 101.840 12.980 102.590 ;
        RECT 13.770 101.840 13.940 102.590 ;
        RECT 14.730 101.840 14.900 102.590 ;
        RECT 15.690 101.840 15.860 102.590 ;
        RECT 16.650 101.840 16.820 102.590 ;
        RECT 19.015 102.590 24.425 102.760 ;
        RECT 12.300 100.480 12.530 101.840 ;
        RECT 12.780 100.480 13.010 101.840 ;
        RECT 13.260 100.480 13.490 101.840 ;
        RECT 13.740 100.480 13.970 101.840 ;
        RECT 14.220 100.480 14.450 101.840 ;
        RECT 14.700 100.480 14.930 101.840 ;
        RECT 15.180 100.480 15.410 101.840 ;
        RECT 15.660 100.480 15.890 101.840 ;
        RECT 16.140 100.480 16.370 101.840 ;
        RECT 16.620 100.480 16.850 101.840 ;
        RECT 17.100 100.480 17.330 101.840 ;
        RECT 10.505 99.755 11.580 99.775 ;
        RECT 1.565 99.605 11.580 99.755 ;
        RECT 1.565 99.585 10.705 99.605 ;
        RECT 1.565 98.920 1.735 99.585 ;
        RECT 2.525 98.920 2.695 99.585 ;
        RECT 3.485 98.920 3.655 99.585 ;
        RECT 4.445 98.920 4.615 99.585 ;
        RECT 5.405 98.920 5.575 99.585 ;
        RECT 6.365 98.920 6.535 99.585 ;
        RECT 1.535 98.400 1.765 98.920 ;
        RECT 2.495 98.400 2.725 98.920 ;
        RECT 3.455 98.400 3.685 98.920 ;
        RECT 4.415 98.400 4.645 98.920 ;
        RECT 5.375 98.400 5.605 98.920 ;
        RECT 6.335 98.400 6.565 98.920 ;
        RECT 11.410 97.720 11.580 99.605 ;
        RECT 12.330 99.775 12.500 100.480 ;
        RECT 13.290 99.775 13.460 100.480 ;
        RECT 14.250 99.775 14.420 100.480 ;
        RECT 15.210 99.775 15.380 100.480 ;
        RECT 16.170 99.775 16.340 100.480 ;
        RECT 17.130 99.775 17.300 100.480 ;
        RECT 19.015 99.775 19.185 102.590 ;
        RECT 20.415 101.840 20.585 102.590 ;
        RECT 21.375 101.840 21.545 102.590 ;
        RECT 22.335 101.840 22.505 102.590 ;
        RECT 23.295 101.840 23.465 102.590 ;
        RECT 24.255 101.840 24.425 102.590 ;
        RECT 20.385 100.480 20.615 101.840 ;
        RECT 21.345 100.480 21.575 101.840 ;
        RECT 22.305 100.480 22.535 101.840 ;
        RECT 23.265 100.480 23.495 101.840 ;
        RECT 24.225 100.480 24.455 101.840 ;
        RECT 12.330 99.605 19.185 99.775 ;
        RECT 12.330 98.940 12.500 99.605 ;
        RECT 13.290 98.940 13.460 99.605 ;
        RECT 14.250 98.940 14.420 99.605 ;
        RECT 15.210 98.940 15.380 99.605 ;
        RECT 16.170 98.940 16.340 99.605 ;
        RECT 17.130 98.940 17.300 99.605 ;
        RECT 19.015 98.965 19.185 99.605 ;
        RECT 26.630 99.310 27.000 99.580 ;
        RECT 18.670 98.960 19.185 98.965 ;
        RECT 12.300 98.420 12.530 98.940 ;
        RECT 12.780 98.420 13.010 98.940 ;
        RECT 13.260 98.420 13.490 98.940 ;
        RECT 13.740 98.420 13.970 98.940 ;
        RECT 14.220 98.420 14.450 98.940 ;
        RECT 14.700 98.420 14.930 98.940 ;
        RECT 15.180 98.420 15.410 98.940 ;
        RECT 15.660 98.420 15.890 98.940 ;
        RECT 16.140 98.420 16.370 98.940 ;
        RECT 16.620 98.420 16.850 98.940 ;
        RECT 17.100 98.420 17.330 98.940 ;
        RECT 18.645 98.465 19.185 98.960 ;
        RECT 18.645 98.460 18.875 98.465 ;
        RECT 12.250 98.265 12.580 98.280 ;
        RECT 12.235 98.005 12.595 98.265 ;
        RECT 12.250 97.980 12.580 98.005 ;
        RECT 12.810 97.720 12.980 98.420 ;
        RECT 13.210 98.265 13.540 98.280 ;
        RECT 13.190 98.005 13.550 98.265 ;
        RECT 13.210 97.980 13.540 98.005 ;
        RECT 13.770 97.720 13.940 98.420 ;
        RECT 14.170 98.265 14.500 98.280 ;
        RECT 14.150 98.005 14.510 98.265 ;
        RECT 14.170 97.980 14.500 98.005 ;
        RECT 14.730 97.720 14.900 98.420 ;
        RECT 15.130 98.265 15.460 98.280 ;
        RECT 15.110 98.005 15.470 98.265 ;
        RECT 15.130 97.980 15.460 98.005 ;
        RECT 15.690 97.720 15.860 98.420 ;
        RECT 16.090 98.260 16.420 98.280 ;
        RECT 16.075 98.000 16.435 98.260 ;
        RECT 16.090 97.980 16.420 98.000 ;
        RECT 16.650 97.720 16.820 98.420 ;
        RECT 17.050 98.260 17.380 98.280 ;
        RECT 17.035 98.000 17.395 98.260 ;
        RECT 17.050 97.980 17.380 98.000 ;
        RECT 11.410 97.550 16.820 97.720 ;
        RECT 19.015 97.720 19.185 98.465 ;
        RECT 20.385 98.420 20.615 98.940 ;
        RECT 21.345 98.420 21.575 98.940 ;
        RECT 22.305 98.420 22.535 98.940 ;
        RECT 23.265 98.420 23.495 98.940 ;
        RECT 24.225 98.420 24.455 98.940 ;
        RECT 19.855 98.265 20.185 98.280 ;
        RECT 19.840 98.005 20.200 98.265 ;
        RECT 19.855 97.980 20.185 98.005 ;
        RECT 20.415 97.720 20.585 98.420 ;
        RECT 20.815 98.265 21.145 98.280 ;
        RECT 20.795 98.005 21.155 98.265 ;
        RECT 20.815 97.980 21.145 98.005 ;
        RECT 21.375 97.720 21.545 98.420 ;
        RECT 21.775 98.265 22.105 98.280 ;
        RECT 21.755 98.005 22.115 98.265 ;
        RECT 21.775 97.980 22.105 98.005 ;
        RECT 22.335 97.720 22.505 98.420 ;
        RECT 22.735 98.265 23.065 98.280 ;
        RECT 22.715 98.005 23.075 98.265 ;
        RECT 22.735 97.980 23.065 98.005 ;
        RECT 23.295 97.720 23.465 98.420 ;
        RECT 23.695 98.260 24.025 98.280 ;
        RECT 23.680 98.000 24.040 98.260 ;
        RECT 23.695 97.980 24.025 98.000 ;
        RECT 24.255 97.720 24.425 98.420 ;
        RECT 24.655 98.260 24.985 98.280 ;
        RECT 24.640 98.000 25.000 98.260 ;
        RECT 24.655 97.980 24.985 98.000 ;
        RECT 19.015 97.550 24.425 97.720 ;
        RECT 11.410 96.155 16.820 96.325 ;
        RECT 1.535 94.025 1.765 95.385 ;
        RECT 2.495 94.025 2.725 95.385 ;
        RECT 3.455 94.025 3.685 95.385 ;
        RECT 4.415 94.025 4.645 95.385 ;
        RECT 5.375 94.025 5.605 95.385 ;
        RECT 6.335 94.025 6.565 95.385 ;
        RECT 1.565 93.320 1.735 94.025 ;
        RECT 2.525 93.320 2.695 94.025 ;
        RECT 3.485 93.320 3.655 94.025 ;
        RECT 4.445 93.320 4.615 94.025 ;
        RECT 5.405 93.320 5.575 94.025 ;
        RECT 6.365 93.320 6.535 94.025 ;
        RECT 11.410 93.340 11.580 96.155 ;
        RECT 12.810 95.405 12.980 96.155 ;
        RECT 13.770 95.405 13.940 96.155 ;
        RECT 14.730 95.405 14.900 96.155 ;
        RECT 15.690 95.405 15.860 96.155 ;
        RECT 16.650 95.405 16.820 96.155 ;
        RECT 19.015 96.155 24.425 96.325 ;
        RECT 12.300 94.045 12.530 95.405 ;
        RECT 12.780 94.045 13.010 95.405 ;
        RECT 13.260 94.045 13.490 95.405 ;
        RECT 13.740 94.045 13.970 95.405 ;
        RECT 14.220 94.045 14.450 95.405 ;
        RECT 14.700 94.045 14.930 95.405 ;
        RECT 15.180 94.045 15.410 95.405 ;
        RECT 15.660 94.045 15.890 95.405 ;
        RECT 16.140 94.045 16.370 95.405 ;
        RECT 16.620 94.045 16.850 95.405 ;
        RECT 17.100 94.045 17.330 95.405 ;
        RECT 10.505 93.320 11.580 93.340 ;
        RECT 1.565 93.170 11.580 93.320 ;
        RECT 1.565 93.150 10.705 93.170 ;
        RECT 1.565 92.485 1.735 93.150 ;
        RECT 2.525 92.485 2.695 93.150 ;
        RECT 3.485 92.485 3.655 93.150 ;
        RECT 4.445 92.485 4.615 93.150 ;
        RECT 5.405 92.485 5.575 93.150 ;
        RECT 6.365 92.485 6.535 93.150 ;
        RECT 1.535 91.965 1.765 92.485 ;
        RECT 2.495 91.965 2.725 92.485 ;
        RECT 3.455 91.965 3.685 92.485 ;
        RECT 4.415 91.965 4.645 92.485 ;
        RECT 5.375 91.965 5.605 92.485 ;
        RECT 6.335 91.965 6.565 92.485 ;
        RECT 11.410 91.285 11.580 93.170 ;
        RECT 12.330 93.340 12.500 94.045 ;
        RECT 13.290 93.340 13.460 94.045 ;
        RECT 14.250 93.340 14.420 94.045 ;
        RECT 15.210 93.340 15.380 94.045 ;
        RECT 16.170 93.340 16.340 94.045 ;
        RECT 17.130 93.340 17.300 94.045 ;
        RECT 19.015 93.340 19.185 96.155 ;
        RECT 20.415 95.405 20.585 96.155 ;
        RECT 21.375 95.405 21.545 96.155 ;
        RECT 22.335 95.405 22.505 96.155 ;
        RECT 23.295 95.405 23.465 96.155 ;
        RECT 24.255 95.405 24.425 96.155 ;
        RECT 20.385 94.045 20.615 95.405 ;
        RECT 21.345 94.045 21.575 95.405 ;
        RECT 22.305 94.045 22.535 95.405 ;
        RECT 23.265 94.045 23.495 95.405 ;
        RECT 24.225 94.045 24.455 95.405 ;
        RECT 12.330 93.170 19.185 93.340 ;
        RECT 12.330 92.505 12.500 93.170 ;
        RECT 13.290 92.505 13.460 93.170 ;
        RECT 14.250 92.505 14.420 93.170 ;
        RECT 15.210 92.505 15.380 93.170 ;
        RECT 16.170 92.505 16.340 93.170 ;
        RECT 17.130 92.505 17.300 93.170 ;
        RECT 19.015 92.530 19.185 93.170 ;
        RECT 26.630 92.875 27.000 93.145 ;
        RECT 18.670 92.525 19.185 92.530 ;
        RECT 12.300 91.985 12.530 92.505 ;
        RECT 12.780 91.985 13.010 92.505 ;
        RECT 13.260 91.985 13.490 92.505 ;
        RECT 13.740 91.985 13.970 92.505 ;
        RECT 14.220 91.985 14.450 92.505 ;
        RECT 14.700 91.985 14.930 92.505 ;
        RECT 15.180 91.985 15.410 92.505 ;
        RECT 15.660 91.985 15.890 92.505 ;
        RECT 16.140 91.985 16.370 92.505 ;
        RECT 16.620 91.985 16.850 92.505 ;
        RECT 17.100 91.985 17.330 92.505 ;
        RECT 18.645 92.030 19.185 92.525 ;
        RECT 18.645 92.025 18.875 92.030 ;
        RECT 12.250 91.830 12.580 91.845 ;
        RECT 12.235 91.570 12.595 91.830 ;
        RECT 12.250 91.545 12.580 91.570 ;
        RECT 12.810 91.285 12.980 91.985 ;
        RECT 13.210 91.830 13.540 91.845 ;
        RECT 13.190 91.570 13.550 91.830 ;
        RECT 13.210 91.545 13.540 91.570 ;
        RECT 13.770 91.285 13.940 91.985 ;
        RECT 14.170 91.830 14.500 91.845 ;
        RECT 14.150 91.570 14.510 91.830 ;
        RECT 14.170 91.545 14.500 91.570 ;
        RECT 14.730 91.285 14.900 91.985 ;
        RECT 15.130 91.830 15.460 91.845 ;
        RECT 15.110 91.570 15.470 91.830 ;
        RECT 15.130 91.545 15.460 91.570 ;
        RECT 15.690 91.285 15.860 91.985 ;
        RECT 16.090 91.825 16.420 91.845 ;
        RECT 16.075 91.565 16.435 91.825 ;
        RECT 16.090 91.545 16.420 91.565 ;
        RECT 16.650 91.285 16.820 91.985 ;
        RECT 17.050 91.825 17.380 91.845 ;
        RECT 17.035 91.565 17.395 91.825 ;
        RECT 17.050 91.545 17.380 91.565 ;
        RECT 11.410 91.115 16.820 91.285 ;
        RECT 19.015 91.285 19.185 92.030 ;
        RECT 20.385 91.985 20.615 92.505 ;
        RECT 21.345 91.985 21.575 92.505 ;
        RECT 22.305 91.985 22.535 92.505 ;
        RECT 23.265 91.985 23.495 92.505 ;
        RECT 24.225 91.985 24.455 92.505 ;
        RECT 19.855 91.830 20.185 91.845 ;
        RECT 19.840 91.570 20.200 91.830 ;
        RECT 19.855 91.545 20.185 91.570 ;
        RECT 20.415 91.285 20.585 91.985 ;
        RECT 20.815 91.830 21.145 91.845 ;
        RECT 20.795 91.570 21.155 91.830 ;
        RECT 20.815 91.545 21.145 91.570 ;
        RECT 21.375 91.285 21.545 91.985 ;
        RECT 21.775 91.830 22.105 91.845 ;
        RECT 21.755 91.570 22.115 91.830 ;
        RECT 21.775 91.545 22.105 91.570 ;
        RECT 22.335 91.285 22.505 91.985 ;
        RECT 22.735 91.830 23.065 91.845 ;
        RECT 22.715 91.570 23.075 91.830 ;
        RECT 22.735 91.545 23.065 91.570 ;
        RECT 23.295 91.285 23.465 91.985 ;
        RECT 23.695 91.825 24.025 91.845 ;
        RECT 23.680 91.565 24.040 91.825 ;
        RECT 23.695 91.545 24.025 91.565 ;
        RECT 24.255 91.285 24.425 91.985 ;
        RECT 24.655 91.825 24.985 91.845 ;
        RECT 24.640 91.565 25.000 91.825 ;
        RECT 24.655 91.545 24.985 91.565 ;
        RECT 19.015 91.115 24.425 91.285 ;
        RECT 11.410 89.720 16.820 89.890 ;
        RECT 1.535 87.590 1.765 88.950 ;
        RECT 2.495 87.590 2.725 88.950 ;
        RECT 3.455 87.590 3.685 88.950 ;
        RECT 4.415 87.590 4.645 88.950 ;
        RECT 5.375 87.590 5.605 88.950 ;
        RECT 6.335 87.590 6.565 88.950 ;
        RECT 1.565 86.885 1.735 87.590 ;
        RECT 2.525 86.885 2.695 87.590 ;
        RECT 3.485 86.885 3.655 87.590 ;
        RECT 4.445 86.885 4.615 87.590 ;
        RECT 5.405 86.885 5.575 87.590 ;
        RECT 6.365 86.885 6.535 87.590 ;
        RECT 11.410 86.905 11.580 89.720 ;
        RECT 12.810 88.970 12.980 89.720 ;
        RECT 13.770 88.970 13.940 89.720 ;
        RECT 14.730 88.970 14.900 89.720 ;
        RECT 15.690 88.970 15.860 89.720 ;
        RECT 16.650 88.970 16.820 89.720 ;
        RECT 19.015 89.720 24.425 89.890 ;
        RECT 12.300 87.610 12.530 88.970 ;
        RECT 12.780 87.610 13.010 88.970 ;
        RECT 13.260 87.610 13.490 88.970 ;
        RECT 13.740 87.610 13.970 88.970 ;
        RECT 14.220 87.610 14.450 88.970 ;
        RECT 14.700 87.610 14.930 88.970 ;
        RECT 15.180 87.610 15.410 88.970 ;
        RECT 15.660 87.610 15.890 88.970 ;
        RECT 16.140 87.610 16.370 88.970 ;
        RECT 16.620 87.610 16.850 88.970 ;
        RECT 17.100 87.610 17.330 88.970 ;
        RECT 10.505 86.885 11.580 86.905 ;
        RECT 1.565 86.735 11.580 86.885 ;
        RECT 1.565 86.715 10.705 86.735 ;
        RECT 1.565 86.050 1.735 86.715 ;
        RECT 2.525 86.050 2.695 86.715 ;
        RECT 3.485 86.050 3.655 86.715 ;
        RECT 4.445 86.050 4.615 86.715 ;
        RECT 5.405 86.050 5.575 86.715 ;
        RECT 6.365 86.050 6.535 86.715 ;
        RECT 1.535 85.530 1.765 86.050 ;
        RECT 2.495 85.530 2.725 86.050 ;
        RECT 3.455 85.530 3.685 86.050 ;
        RECT 4.415 85.530 4.645 86.050 ;
        RECT 5.375 85.530 5.605 86.050 ;
        RECT 6.335 85.530 6.565 86.050 ;
        RECT 11.410 84.850 11.580 86.735 ;
        RECT 12.330 86.905 12.500 87.610 ;
        RECT 13.290 86.905 13.460 87.610 ;
        RECT 14.250 86.905 14.420 87.610 ;
        RECT 15.210 86.905 15.380 87.610 ;
        RECT 16.170 86.905 16.340 87.610 ;
        RECT 17.130 86.905 17.300 87.610 ;
        RECT 19.015 86.905 19.185 89.720 ;
        RECT 20.415 88.970 20.585 89.720 ;
        RECT 21.375 88.970 21.545 89.720 ;
        RECT 22.335 88.970 22.505 89.720 ;
        RECT 23.295 88.970 23.465 89.720 ;
        RECT 24.255 88.970 24.425 89.720 ;
        RECT 20.385 87.610 20.615 88.970 ;
        RECT 21.345 87.610 21.575 88.970 ;
        RECT 22.305 87.610 22.535 88.970 ;
        RECT 23.265 87.610 23.495 88.970 ;
        RECT 24.225 87.610 24.455 88.970 ;
        RECT 12.330 86.735 19.185 86.905 ;
        RECT 12.330 86.070 12.500 86.735 ;
        RECT 13.290 86.070 13.460 86.735 ;
        RECT 14.250 86.070 14.420 86.735 ;
        RECT 15.210 86.070 15.380 86.735 ;
        RECT 16.170 86.070 16.340 86.735 ;
        RECT 17.130 86.070 17.300 86.735 ;
        RECT 19.015 86.095 19.185 86.735 ;
        RECT 26.630 86.440 27.000 86.710 ;
        RECT 18.670 86.090 19.185 86.095 ;
        RECT 12.300 85.550 12.530 86.070 ;
        RECT 12.780 85.550 13.010 86.070 ;
        RECT 13.260 85.550 13.490 86.070 ;
        RECT 13.740 85.550 13.970 86.070 ;
        RECT 14.220 85.550 14.450 86.070 ;
        RECT 14.700 85.550 14.930 86.070 ;
        RECT 15.180 85.550 15.410 86.070 ;
        RECT 15.660 85.550 15.890 86.070 ;
        RECT 16.140 85.550 16.370 86.070 ;
        RECT 16.620 85.550 16.850 86.070 ;
        RECT 17.100 85.550 17.330 86.070 ;
        RECT 18.645 85.595 19.185 86.090 ;
        RECT 18.645 85.590 18.875 85.595 ;
        RECT 12.250 85.395 12.580 85.410 ;
        RECT 12.235 85.135 12.595 85.395 ;
        RECT 12.250 85.110 12.580 85.135 ;
        RECT 12.810 84.850 12.980 85.550 ;
        RECT 13.210 85.395 13.540 85.410 ;
        RECT 13.190 85.135 13.550 85.395 ;
        RECT 13.210 85.110 13.540 85.135 ;
        RECT 13.770 84.850 13.940 85.550 ;
        RECT 14.170 85.395 14.500 85.410 ;
        RECT 14.150 85.135 14.510 85.395 ;
        RECT 14.170 85.110 14.500 85.135 ;
        RECT 14.730 84.850 14.900 85.550 ;
        RECT 15.130 85.395 15.460 85.410 ;
        RECT 15.110 85.135 15.470 85.395 ;
        RECT 15.130 85.110 15.460 85.135 ;
        RECT 15.690 84.850 15.860 85.550 ;
        RECT 16.090 85.390 16.420 85.410 ;
        RECT 16.075 85.130 16.435 85.390 ;
        RECT 16.090 85.110 16.420 85.130 ;
        RECT 16.650 84.850 16.820 85.550 ;
        RECT 17.050 85.390 17.380 85.410 ;
        RECT 17.035 85.130 17.395 85.390 ;
        RECT 17.050 85.110 17.380 85.130 ;
        RECT 11.410 84.680 16.820 84.850 ;
        RECT 19.015 84.850 19.185 85.595 ;
        RECT 20.385 85.550 20.615 86.070 ;
        RECT 21.345 85.550 21.575 86.070 ;
        RECT 22.305 85.550 22.535 86.070 ;
        RECT 23.265 85.550 23.495 86.070 ;
        RECT 24.225 85.550 24.455 86.070 ;
        RECT 19.855 85.395 20.185 85.410 ;
        RECT 19.840 85.135 20.200 85.395 ;
        RECT 19.855 85.110 20.185 85.135 ;
        RECT 20.415 84.850 20.585 85.550 ;
        RECT 20.815 85.395 21.145 85.410 ;
        RECT 20.795 85.135 21.155 85.395 ;
        RECT 20.815 85.110 21.145 85.135 ;
        RECT 21.375 84.850 21.545 85.550 ;
        RECT 21.775 85.395 22.105 85.410 ;
        RECT 21.755 85.135 22.115 85.395 ;
        RECT 21.775 85.110 22.105 85.135 ;
        RECT 22.335 84.850 22.505 85.550 ;
        RECT 22.735 85.395 23.065 85.410 ;
        RECT 22.715 85.135 23.075 85.395 ;
        RECT 22.735 85.110 23.065 85.135 ;
        RECT 23.295 84.850 23.465 85.550 ;
        RECT 23.695 85.390 24.025 85.410 ;
        RECT 23.680 85.130 24.040 85.390 ;
        RECT 23.695 85.110 24.025 85.130 ;
        RECT 24.255 84.850 24.425 85.550 ;
        RECT 24.655 85.390 24.985 85.410 ;
        RECT 24.640 85.130 25.000 85.390 ;
        RECT 24.655 85.110 24.985 85.130 ;
        RECT 19.015 84.680 24.425 84.850 ;
        RECT 11.410 83.285 16.820 83.455 ;
        RECT 1.535 81.155 1.765 82.515 ;
        RECT 2.495 81.155 2.725 82.515 ;
        RECT 3.455 81.155 3.685 82.515 ;
        RECT 4.415 81.155 4.645 82.515 ;
        RECT 5.375 81.155 5.605 82.515 ;
        RECT 6.335 81.155 6.565 82.515 ;
        RECT 1.565 80.450 1.735 81.155 ;
        RECT 2.525 80.450 2.695 81.155 ;
        RECT 3.485 80.450 3.655 81.155 ;
        RECT 4.445 80.450 4.615 81.155 ;
        RECT 5.405 80.450 5.575 81.155 ;
        RECT 6.365 80.450 6.535 81.155 ;
        RECT 11.410 80.470 11.580 83.285 ;
        RECT 12.810 82.535 12.980 83.285 ;
        RECT 13.770 82.535 13.940 83.285 ;
        RECT 14.730 82.535 14.900 83.285 ;
        RECT 15.690 82.535 15.860 83.285 ;
        RECT 16.650 82.535 16.820 83.285 ;
        RECT 19.015 83.285 24.425 83.455 ;
        RECT 12.300 81.175 12.530 82.535 ;
        RECT 12.780 81.175 13.010 82.535 ;
        RECT 13.260 81.175 13.490 82.535 ;
        RECT 13.740 81.175 13.970 82.535 ;
        RECT 14.220 81.175 14.450 82.535 ;
        RECT 14.700 81.175 14.930 82.535 ;
        RECT 15.180 81.175 15.410 82.535 ;
        RECT 15.660 81.175 15.890 82.535 ;
        RECT 16.140 81.175 16.370 82.535 ;
        RECT 16.620 81.175 16.850 82.535 ;
        RECT 17.100 81.175 17.330 82.535 ;
        RECT 10.505 80.450 11.580 80.470 ;
        RECT 1.565 80.300 11.580 80.450 ;
        RECT 1.565 80.280 10.705 80.300 ;
        RECT 1.565 79.615 1.735 80.280 ;
        RECT 2.525 79.615 2.695 80.280 ;
        RECT 3.485 79.615 3.655 80.280 ;
        RECT 4.445 79.615 4.615 80.280 ;
        RECT 5.405 79.615 5.575 80.280 ;
        RECT 6.365 79.615 6.535 80.280 ;
        RECT 1.535 79.095 1.765 79.615 ;
        RECT 2.495 79.095 2.725 79.615 ;
        RECT 3.455 79.095 3.685 79.615 ;
        RECT 4.415 79.095 4.645 79.615 ;
        RECT 5.375 79.095 5.605 79.615 ;
        RECT 6.335 79.095 6.565 79.615 ;
        RECT 11.410 78.415 11.580 80.300 ;
        RECT 12.330 80.470 12.500 81.175 ;
        RECT 13.290 80.470 13.460 81.175 ;
        RECT 14.250 80.470 14.420 81.175 ;
        RECT 15.210 80.470 15.380 81.175 ;
        RECT 16.170 80.470 16.340 81.175 ;
        RECT 17.130 80.470 17.300 81.175 ;
        RECT 19.015 80.470 19.185 83.285 ;
        RECT 20.415 82.535 20.585 83.285 ;
        RECT 21.375 82.535 21.545 83.285 ;
        RECT 22.335 82.535 22.505 83.285 ;
        RECT 23.295 82.535 23.465 83.285 ;
        RECT 24.255 82.535 24.425 83.285 ;
        RECT 20.385 81.175 20.615 82.535 ;
        RECT 21.345 81.175 21.575 82.535 ;
        RECT 22.305 81.175 22.535 82.535 ;
        RECT 23.265 81.175 23.495 82.535 ;
        RECT 24.225 81.175 24.455 82.535 ;
        RECT 12.330 80.300 19.185 80.470 ;
        RECT 12.330 79.635 12.500 80.300 ;
        RECT 13.290 79.635 13.460 80.300 ;
        RECT 14.250 79.635 14.420 80.300 ;
        RECT 15.210 79.635 15.380 80.300 ;
        RECT 16.170 79.635 16.340 80.300 ;
        RECT 17.130 79.635 17.300 80.300 ;
        RECT 19.015 79.660 19.185 80.300 ;
        RECT 26.630 80.005 27.000 80.275 ;
        RECT 18.670 79.655 19.185 79.660 ;
        RECT 12.300 79.115 12.530 79.635 ;
        RECT 12.780 79.115 13.010 79.635 ;
        RECT 13.260 79.115 13.490 79.635 ;
        RECT 13.740 79.115 13.970 79.635 ;
        RECT 14.220 79.115 14.450 79.635 ;
        RECT 14.700 79.115 14.930 79.635 ;
        RECT 15.180 79.115 15.410 79.635 ;
        RECT 15.660 79.115 15.890 79.635 ;
        RECT 16.140 79.115 16.370 79.635 ;
        RECT 16.620 79.115 16.850 79.635 ;
        RECT 17.100 79.115 17.330 79.635 ;
        RECT 18.645 79.160 19.185 79.655 ;
        RECT 18.645 79.155 18.875 79.160 ;
        RECT 12.250 78.960 12.580 78.975 ;
        RECT 12.235 78.700 12.595 78.960 ;
        RECT 12.250 78.675 12.580 78.700 ;
        RECT 12.810 78.415 12.980 79.115 ;
        RECT 13.210 78.960 13.540 78.975 ;
        RECT 13.190 78.700 13.550 78.960 ;
        RECT 13.210 78.675 13.540 78.700 ;
        RECT 13.770 78.415 13.940 79.115 ;
        RECT 14.170 78.960 14.500 78.975 ;
        RECT 14.150 78.700 14.510 78.960 ;
        RECT 14.170 78.675 14.500 78.700 ;
        RECT 14.730 78.415 14.900 79.115 ;
        RECT 15.130 78.960 15.460 78.975 ;
        RECT 15.110 78.700 15.470 78.960 ;
        RECT 15.130 78.675 15.460 78.700 ;
        RECT 15.690 78.415 15.860 79.115 ;
        RECT 16.090 78.955 16.420 78.975 ;
        RECT 16.075 78.695 16.435 78.955 ;
        RECT 16.090 78.675 16.420 78.695 ;
        RECT 16.650 78.415 16.820 79.115 ;
        RECT 17.050 78.955 17.380 78.975 ;
        RECT 17.035 78.695 17.395 78.955 ;
        RECT 17.050 78.675 17.380 78.695 ;
        RECT 11.410 78.245 16.820 78.415 ;
        RECT 19.015 78.415 19.185 79.160 ;
        RECT 20.385 79.115 20.615 79.635 ;
        RECT 21.345 79.115 21.575 79.635 ;
        RECT 22.305 79.115 22.535 79.635 ;
        RECT 23.265 79.115 23.495 79.635 ;
        RECT 24.225 79.115 24.455 79.635 ;
        RECT 19.855 78.960 20.185 78.975 ;
        RECT 19.840 78.700 20.200 78.960 ;
        RECT 19.855 78.675 20.185 78.700 ;
        RECT 20.415 78.415 20.585 79.115 ;
        RECT 20.815 78.960 21.145 78.975 ;
        RECT 20.795 78.700 21.155 78.960 ;
        RECT 20.815 78.675 21.145 78.700 ;
        RECT 21.375 78.415 21.545 79.115 ;
        RECT 21.775 78.960 22.105 78.975 ;
        RECT 21.755 78.700 22.115 78.960 ;
        RECT 21.775 78.675 22.105 78.700 ;
        RECT 22.335 78.415 22.505 79.115 ;
        RECT 22.735 78.960 23.065 78.975 ;
        RECT 22.715 78.700 23.075 78.960 ;
        RECT 22.735 78.675 23.065 78.700 ;
        RECT 23.295 78.415 23.465 79.115 ;
        RECT 23.695 78.955 24.025 78.975 ;
        RECT 23.680 78.695 24.040 78.955 ;
        RECT 23.695 78.675 24.025 78.695 ;
        RECT 24.255 78.415 24.425 79.115 ;
        RECT 24.655 78.955 24.985 78.975 ;
        RECT 24.640 78.695 25.000 78.955 ;
        RECT 24.655 78.675 24.985 78.695 ;
        RECT 19.015 78.245 24.425 78.415 ;
        RECT 11.410 76.850 16.820 77.020 ;
        RECT 1.535 74.720 1.765 76.080 ;
        RECT 2.495 74.720 2.725 76.080 ;
        RECT 3.455 74.720 3.685 76.080 ;
        RECT 4.415 74.720 4.645 76.080 ;
        RECT 5.375 74.720 5.605 76.080 ;
        RECT 6.335 74.720 6.565 76.080 ;
        RECT 1.565 74.015 1.735 74.720 ;
        RECT 2.525 74.015 2.695 74.720 ;
        RECT 3.485 74.015 3.655 74.720 ;
        RECT 4.445 74.015 4.615 74.720 ;
        RECT 5.405 74.015 5.575 74.720 ;
        RECT 6.365 74.015 6.535 74.720 ;
        RECT 11.410 74.035 11.580 76.850 ;
        RECT 12.810 76.100 12.980 76.850 ;
        RECT 13.770 76.100 13.940 76.850 ;
        RECT 14.730 76.100 14.900 76.850 ;
        RECT 15.690 76.100 15.860 76.850 ;
        RECT 16.650 76.100 16.820 76.850 ;
        RECT 19.015 76.850 24.425 77.020 ;
        RECT 12.300 74.740 12.530 76.100 ;
        RECT 12.780 74.740 13.010 76.100 ;
        RECT 13.260 74.740 13.490 76.100 ;
        RECT 13.740 74.740 13.970 76.100 ;
        RECT 14.220 74.740 14.450 76.100 ;
        RECT 14.700 74.740 14.930 76.100 ;
        RECT 15.180 74.740 15.410 76.100 ;
        RECT 15.660 74.740 15.890 76.100 ;
        RECT 16.140 74.740 16.370 76.100 ;
        RECT 16.620 74.740 16.850 76.100 ;
        RECT 17.100 74.740 17.330 76.100 ;
        RECT 10.505 74.015 11.580 74.035 ;
        RECT 1.565 73.865 11.580 74.015 ;
        RECT 1.565 73.845 10.705 73.865 ;
        RECT 1.565 73.180 1.735 73.845 ;
        RECT 2.525 73.180 2.695 73.845 ;
        RECT 3.485 73.180 3.655 73.845 ;
        RECT 4.445 73.180 4.615 73.845 ;
        RECT 5.405 73.180 5.575 73.845 ;
        RECT 6.365 73.180 6.535 73.845 ;
        RECT 1.535 72.660 1.765 73.180 ;
        RECT 2.495 72.660 2.725 73.180 ;
        RECT 3.455 72.660 3.685 73.180 ;
        RECT 4.415 72.660 4.645 73.180 ;
        RECT 5.375 72.660 5.605 73.180 ;
        RECT 6.335 72.660 6.565 73.180 ;
        RECT 11.410 71.980 11.580 73.865 ;
        RECT 12.330 74.035 12.500 74.740 ;
        RECT 13.290 74.035 13.460 74.740 ;
        RECT 14.250 74.035 14.420 74.740 ;
        RECT 15.210 74.035 15.380 74.740 ;
        RECT 16.170 74.035 16.340 74.740 ;
        RECT 17.130 74.035 17.300 74.740 ;
        RECT 19.015 74.035 19.185 76.850 ;
        RECT 20.415 76.100 20.585 76.850 ;
        RECT 21.375 76.100 21.545 76.850 ;
        RECT 22.335 76.100 22.505 76.850 ;
        RECT 23.295 76.100 23.465 76.850 ;
        RECT 24.255 76.100 24.425 76.850 ;
        RECT 20.385 74.740 20.615 76.100 ;
        RECT 21.345 74.740 21.575 76.100 ;
        RECT 22.305 74.740 22.535 76.100 ;
        RECT 23.265 74.740 23.495 76.100 ;
        RECT 24.225 74.740 24.455 76.100 ;
        RECT 12.330 73.865 19.185 74.035 ;
        RECT 12.330 73.200 12.500 73.865 ;
        RECT 13.290 73.200 13.460 73.865 ;
        RECT 14.250 73.200 14.420 73.865 ;
        RECT 15.210 73.200 15.380 73.865 ;
        RECT 16.170 73.200 16.340 73.865 ;
        RECT 17.130 73.200 17.300 73.865 ;
        RECT 19.015 73.225 19.185 73.865 ;
        RECT 26.630 73.570 27.000 73.840 ;
        RECT 18.670 73.220 19.185 73.225 ;
        RECT 12.300 72.680 12.530 73.200 ;
        RECT 12.780 72.680 13.010 73.200 ;
        RECT 13.260 72.680 13.490 73.200 ;
        RECT 13.740 72.680 13.970 73.200 ;
        RECT 14.220 72.680 14.450 73.200 ;
        RECT 14.700 72.680 14.930 73.200 ;
        RECT 15.180 72.680 15.410 73.200 ;
        RECT 15.660 72.680 15.890 73.200 ;
        RECT 16.140 72.680 16.370 73.200 ;
        RECT 16.620 72.680 16.850 73.200 ;
        RECT 17.100 72.680 17.330 73.200 ;
        RECT 18.645 72.725 19.185 73.220 ;
        RECT 18.645 72.720 18.875 72.725 ;
        RECT 12.250 72.525 12.580 72.540 ;
        RECT 12.235 72.265 12.595 72.525 ;
        RECT 12.250 72.240 12.580 72.265 ;
        RECT 12.810 71.980 12.980 72.680 ;
        RECT 13.210 72.525 13.540 72.540 ;
        RECT 13.190 72.265 13.550 72.525 ;
        RECT 13.210 72.240 13.540 72.265 ;
        RECT 13.770 71.980 13.940 72.680 ;
        RECT 14.170 72.525 14.500 72.540 ;
        RECT 14.150 72.265 14.510 72.525 ;
        RECT 14.170 72.240 14.500 72.265 ;
        RECT 14.730 71.980 14.900 72.680 ;
        RECT 15.130 72.525 15.460 72.540 ;
        RECT 15.110 72.265 15.470 72.525 ;
        RECT 15.130 72.240 15.460 72.265 ;
        RECT 15.690 71.980 15.860 72.680 ;
        RECT 16.090 72.520 16.420 72.540 ;
        RECT 16.075 72.260 16.435 72.520 ;
        RECT 16.090 72.240 16.420 72.260 ;
        RECT 16.650 71.980 16.820 72.680 ;
        RECT 17.050 72.520 17.380 72.540 ;
        RECT 17.035 72.260 17.395 72.520 ;
        RECT 17.050 72.240 17.380 72.260 ;
        RECT 11.410 71.810 16.820 71.980 ;
        RECT 19.015 71.980 19.185 72.725 ;
        RECT 20.385 72.680 20.615 73.200 ;
        RECT 21.345 72.680 21.575 73.200 ;
        RECT 22.305 72.680 22.535 73.200 ;
        RECT 23.265 72.680 23.495 73.200 ;
        RECT 24.225 72.680 24.455 73.200 ;
        RECT 19.855 72.525 20.185 72.540 ;
        RECT 19.840 72.265 20.200 72.525 ;
        RECT 19.855 72.240 20.185 72.265 ;
        RECT 20.415 71.980 20.585 72.680 ;
        RECT 20.815 72.525 21.145 72.540 ;
        RECT 20.795 72.265 21.155 72.525 ;
        RECT 20.815 72.240 21.145 72.265 ;
        RECT 21.375 71.980 21.545 72.680 ;
        RECT 21.775 72.525 22.105 72.540 ;
        RECT 21.755 72.265 22.115 72.525 ;
        RECT 21.775 72.240 22.105 72.265 ;
        RECT 22.335 71.980 22.505 72.680 ;
        RECT 22.735 72.525 23.065 72.540 ;
        RECT 22.715 72.265 23.075 72.525 ;
        RECT 22.735 72.240 23.065 72.265 ;
        RECT 23.295 71.980 23.465 72.680 ;
        RECT 23.695 72.520 24.025 72.540 ;
        RECT 23.680 72.260 24.040 72.520 ;
        RECT 23.695 72.240 24.025 72.260 ;
        RECT 24.255 71.980 24.425 72.680 ;
        RECT 24.655 72.520 24.985 72.540 ;
        RECT 24.640 72.260 25.000 72.520 ;
        RECT 24.655 72.240 24.985 72.260 ;
        RECT 19.015 71.810 24.425 71.980 ;
        RECT 11.410 70.415 16.820 70.585 ;
        RECT 1.535 68.285 1.765 69.645 ;
        RECT 2.495 68.285 2.725 69.645 ;
        RECT 3.455 68.285 3.685 69.645 ;
        RECT 4.415 68.285 4.645 69.645 ;
        RECT 5.375 68.285 5.605 69.645 ;
        RECT 6.335 68.285 6.565 69.645 ;
        RECT 1.565 67.580 1.735 68.285 ;
        RECT 2.525 67.580 2.695 68.285 ;
        RECT 3.485 67.580 3.655 68.285 ;
        RECT 4.445 67.580 4.615 68.285 ;
        RECT 5.405 67.580 5.575 68.285 ;
        RECT 6.365 67.580 6.535 68.285 ;
        RECT 11.410 67.600 11.580 70.415 ;
        RECT 12.810 69.665 12.980 70.415 ;
        RECT 13.770 69.665 13.940 70.415 ;
        RECT 14.730 69.665 14.900 70.415 ;
        RECT 15.690 69.665 15.860 70.415 ;
        RECT 16.650 69.665 16.820 70.415 ;
        RECT 19.015 70.415 24.425 70.585 ;
        RECT 12.300 68.305 12.530 69.665 ;
        RECT 12.780 68.305 13.010 69.665 ;
        RECT 13.260 68.305 13.490 69.665 ;
        RECT 13.740 68.305 13.970 69.665 ;
        RECT 14.220 68.305 14.450 69.665 ;
        RECT 14.700 68.305 14.930 69.665 ;
        RECT 15.180 68.305 15.410 69.665 ;
        RECT 15.660 68.305 15.890 69.665 ;
        RECT 16.140 68.305 16.370 69.665 ;
        RECT 16.620 68.305 16.850 69.665 ;
        RECT 17.100 68.305 17.330 69.665 ;
        RECT 10.505 67.580 11.580 67.600 ;
        RECT 1.565 67.430 11.580 67.580 ;
        RECT 1.565 67.410 10.705 67.430 ;
        RECT 1.565 66.745 1.735 67.410 ;
        RECT 2.525 66.745 2.695 67.410 ;
        RECT 3.485 66.745 3.655 67.410 ;
        RECT 4.445 66.745 4.615 67.410 ;
        RECT 5.405 66.745 5.575 67.410 ;
        RECT 6.365 66.745 6.535 67.410 ;
        RECT 1.535 66.225 1.765 66.745 ;
        RECT 2.495 66.225 2.725 66.745 ;
        RECT 3.455 66.225 3.685 66.745 ;
        RECT 4.415 66.225 4.645 66.745 ;
        RECT 5.375 66.225 5.605 66.745 ;
        RECT 6.335 66.225 6.565 66.745 ;
        RECT 11.410 65.545 11.580 67.430 ;
        RECT 12.330 67.600 12.500 68.305 ;
        RECT 13.290 67.600 13.460 68.305 ;
        RECT 14.250 67.600 14.420 68.305 ;
        RECT 15.210 67.600 15.380 68.305 ;
        RECT 16.170 67.600 16.340 68.305 ;
        RECT 17.130 67.600 17.300 68.305 ;
        RECT 19.015 67.600 19.185 70.415 ;
        RECT 20.415 69.665 20.585 70.415 ;
        RECT 21.375 69.665 21.545 70.415 ;
        RECT 22.335 69.665 22.505 70.415 ;
        RECT 23.295 69.665 23.465 70.415 ;
        RECT 24.255 69.665 24.425 70.415 ;
        RECT 20.385 68.305 20.615 69.665 ;
        RECT 21.345 68.305 21.575 69.665 ;
        RECT 22.305 68.305 22.535 69.665 ;
        RECT 23.265 68.305 23.495 69.665 ;
        RECT 24.225 68.305 24.455 69.665 ;
        RECT 12.330 67.430 19.185 67.600 ;
        RECT 12.330 66.765 12.500 67.430 ;
        RECT 13.290 66.765 13.460 67.430 ;
        RECT 14.250 66.765 14.420 67.430 ;
        RECT 15.210 66.765 15.380 67.430 ;
        RECT 16.170 66.765 16.340 67.430 ;
        RECT 17.130 66.765 17.300 67.430 ;
        RECT 19.015 66.790 19.185 67.430 ;
        RECT 26.630 67.135 27.000 67.405 ;
        RECT 18.670 66.785 19.185 66.790 ;
        RECT 12.300 66.245 12.530 66.765 ;
        RECT 12.780 66.245 13.010 66.765 ;
        RECT 13.260 66.245 13.490 66.765 ;
        RECT 13.740 66.245 13.970 66.765 ;
        RECT 14.220 66.245 14.450 66.765 ;
        RECT 14.700 66.245 14.930 66.765 ;
        RECT 15.180 66.245 15.410 66.765 ;
        RECT 15.660 66.245 15.890 66.765 ;
        RECT 16.140 66.245 16.370 66.765 ;
        RECT 16.620 66.245 16.850 66.765 ;
        RECT 17.100 66.245 17.330 66.765 ;
        RECT 18.645 66.290 19.185 66.785 ;
        RECT 18.645 66.285 18.875 66.290 ;
        RECT 12.250 66.090 12.580 66.105 ;
        RECT 12.235 65.830 12.595 66.090 ;
        RECT 12.250 65.805 12.580 65.830 ;
        RECT 12.810 65.545 12.980 66.245 ;
        RECT 13.210 66.090 13.540 66.105 ;
        RECT 13.190 65.830 13.550 66.090 ;
        RECT 13.210 65.805 13.540 65.830 ;
        RECT 13.770 65.545 13.940 66.245 ;
        RECT 14.170 66.090 14.500 66.105 ;
        RECT 14.150 65.830 14.510 66.090 ;
        RECT 14.170 65.805 14.500 65.830 ;
        RECT 14.730 65.545 14.900 66.245 ;
        RECT 15.130 66.090 15.460 66.105 ;
        RECT 15.110 65.830 15.470 66.090 ;
        RECT 15.130 65.805 15.460 65.830 ;
        RECT 15.690 65.545 15.860 66.245 ;
        RECT 16.090 66.085 16.420 66.105 ;
        RECT 16.075 65.825 16.435 66.085 ;
        RECT 16.090 65.805 16.420 65.825 ;
        RECT 16.650 65.545 16.820 66.245 ;
        RECT 17.050 66.085 17.380 66.105 ;
        RECT 17.035 65.825 17.395 66.085 ;
        RECT 17.050 65.805 17.380 65.825 ;
        RECT 11.410 65.375 16.820 65.545 ;
        RECT 19.015 65.545 19.185 66.290 ;
        RECT 20.385 66.245 20.615 66.765 ;
        RECT 21.345 66.245 21.575 66.765 ;
        RECT 22.305 66.245 22.535 66.765 ;
        RECT 23.265 66.245 23.495 66.765 ;
        RECT 24.225 66.245 24.455 66.765 ;
        RECT 19.855 66.090 20.185 66.105 ;
        RECT 19.840 65.830 20.200 66.090 ;
        RECT 19.855 65.805 20.185 65.830 ;
        RECT 20.415 65.545 20.585 66.245 ;
        RECT 20.815 66.090 21.145 66.105 ;
        RECT 20.795 65.830 21.155 66.090 ;
        RECT 20.815 65.805 21.145 65.830 ;
        RECT 21.375 65.545 21.545 66.245 ;
        RECT 21.775 66.090 22.105 66.105 ;
        RECT 21.755 65.830 22.115 66.090 ;
        RECT 21.775 65.805 22.105 65.830 ;
        RECT 22.335 65.545 22.505 66.245 ;
        RECT 22.735 66.090 23.065 66.105 ;
        RECT 22.715 65.830 23.075 66.090 ;
        RECT 22.735 65.805 23.065 65.830 ;
        RECT 23.295 65.545 23.465 66.245 ;
        RECT 23.695 66.085 24.025 66.105 ;
        RECT 23.680 65.825 24.040 66.085 ;
        RECT 23.695 65.805 24.025 65.825 ;
        RECT 24.255 65.545 24.425 66.245 ;
        RECT 24.655 66.085 24.985 66.105 ;
        RECT 24.640 65.825 25.000 66.085 ;
        RECT 24.655 65.805 24.985 65.825 ;
        RECT 19.015 65.375 24.425 65.545 ;
        RECT 11.410 63.980 16.820 64.150 ;
        RECT 1.535 61.850 1.765 63.210 ;
        RECT 2.495 61.850 2.725 63.210 ;
        RECT 3.455 61.850 3.685 63.210 ;
        RECT 4.415 61.850 4.645 63.210 ;
        RECT 5.375 61.850 5.605 63.210 ;
        RECT 6.335 61.850 6.565 63.210 ;
        RECT 1.565 61.145 1.735 61.850 ;
        RECT 2.525 61.145 2.695 61.850 ;
        RECT 3.485 61.145 3.655 61.850 ;
        RECT 4.445 61.145 4.615 61.850 ;
        RECT 5.405 61.145 5.575 61.850 ;
        RECT 6.365 61.145 6.535 61.850 ;
        RECT 11.410 61.165 11.580 63.980 ;
        RECT 12.810 63.230 12.980 63.980 ;
        RECT 13.770 63.230 13.940 63.980 ;
        RECT 14.730 63.230 14.900 63.980 ;
        RECT 15.690 63.230 15.860 63.980 ;
        RECT 16.650 63.230 16.820 63.980 ;
        RECT 19.015 63.980 24.425 64.150 ;
        RECT 12.300 61.870 12.530 63.230 ;
        RECT 12.780 61.870 13.010 63.230 ;
        RECT 13.260 61.870 13.490 63.230 ;
        RECT 13.740 61.870 13.970 63.230 ;
        RECT 14.220 61.870 14.450 63.230 ;
        RECT 14.700 61.870 14.930 63.230 ;
        RECT 15.180 61.870 15.410 63.230 ;
        RECT 15.660 61.870 15.890 63.230 ;
        RECT 16.140 61.870 16.370 63.230 ;
        RECT 16.620 61.870 16.850 63.230 ;
        RECT 17.100 61.870 17.330 63.230 ;
        RECT 10.505 61.145 11.580 61.165 ;
        RECT 1.565 60.995 11.580 61.145 ;
        RECT 1.565 60.975 10.705 60.995 ;
        RECT 1.565 60.310 1.735 60.975 ;
        RECT 2.525 60.310 2.695 60.975 ;
        RECT 3.485 60.310 3.655 60.975 ;
        RECT 4.445 60.310 4.615 60.975 ;
        RECT 5.405 60.310 5.575 60.975 ;
        RECT 6.365 60.310 6.535 60.975 ;
        RECT 1.535 59.790 1.765 60.310 ;
        RECT 2.495 59.790 2.725 60.310 ;
        RECT 3.455 59.790 3.685 60.310 ;
        RECT 4.415 59.790 4.645 60.310 ;
        RECT 5.375 59.790 5.605 60.310 ;
        RECT 6.335 59.790 6.565 60.310 ;
        RECT 11.410 59.110 11.580 60.995 ;
        RECT 12.330 61.165 12.500 61.870 ;
        RECT 13.290 61.165 13.460 61.870 ;
        RECT 14.250 61.165 14.420 61.870 ;
        RECT 15.210 61.165 15.380 61.870 ;
        RECT 16.170 61.165 16.340 61.870 ;
        RECT 17.130 61.165 17.300 61.870 ;
        RECT 19.015 61.165 19.185 63.980 ;
        RECT 20.415 63.230 20.585 63.980 ;
        RECT 21.375 63.230 21.545 63.980 ;
        RECT 22.335 63.230 22.505 63.980 ;
        RECT 23.295 63.230 23.465 63.980 ;
        RECT 24.255 63.230 24.425 63.980 ;
        RECT 20.385 61.870 20.615 63.230 ;
        RECT 21.345 61.870 21.575 63.230 ;
        RECT 22.305 61.870 22.535 63.230 ;
        RECT 23.265 61.870 23.495 63.230 ;
        RECT 24.225 61.870 24.455 63.230 ;
        RECT 12.330 60.995 19.185 61.165 ;
        RECT 12.330 60.330 12.500 60.995 ;
        RECT 13.290 60.330 13.460 60.995 ;
        RECT 14.250 60.330 14.420 60.995 ;
        RECT 15.210 60.330 15.380 60.995 ;
        RECT 16.170 60.330 16.340 60.995 ;
        RECT 17.130 60.330 17.300 60.995 ;
        RECT 19.015 60.355 19.185 60.995 ;
        RECT 26.630 60.700 27.000 60.970 ;
        RECT 18.670 60.350 19.185 60.355 ;
        RECT 12.300 59.810 12.530 60.330 ;
        RECT 12.780 59.810 13.010 60.330 ;
        RECT 13.260 59.810 13.490 60.330 ;
        RECT 13.740 59.810 13.970 60.330 ;
        RECT 14.220 59.810 14.450 60.330 ;
        RECT 14.700 59.810 14.930 60.330 ;
        RECT 15.180 59.810 15.410 60.330 ;
        RECT 15.660 59.810 15.890 60.330 ;
        RECT 16.140 59.810 16.370 60.330 ;
        RECT 16.620 59.810 16.850 60.330 ;
        RECT 17.100 59.810 17.330 60.330 ;
        RECT 18.645 59.855 19.185 60.350 ;
        RECT 18.645 59.850 18.875 59.855 ;
        RECT 12.250 59.655 12.580 59.670 ;
        RECT 12.235 59.395 12.595 59.655 ;
        RECT 12.250 59.370 12.580 59.395 ;
        RECT 12.810 59.110 12.980 59.810 ;
        RECT 13.210 59.655 13.540 59.670 ;
        RECT 13.190 59.395 13.550 59.655 ;
        RECT 13.210 59.370 13.540 59.395 ;
        RECT 13.770 59.110 13.940 59.810 ;
        RECT 14.170 59.655 14.500 59.670 ;
        RECT 14.150 59.395 14.510 59.655 ;
        RECT 14.170 59.370 14.500 59.395 ;
        RECT 14.730 59.110 14.900 59.810 ;
        RECT 15.130 59.655 15.460 59.670 ;
        RECT 15.110 59.395 15.470 59.655 ;
        RECT 15.130 59.370 15.460 59.395 ;
        RECT 15.690 59.110 15.860 59.810 ;
        RECT 16.090 59.650 16.420 59.670 ;
        RECT 16.075 59.390 16.435 59.650 ;
        RECT 16.090 59.370 16.420 59.390 ;
        RECT 16.650 59.110 16.820 59.810 ;
        RECT 17.050 59.650 17.380 59.670 ;
        RECT 17.035 59.390 17.395 59.650 ;
        RECT 17.050 59.370 17.380 59.390 ;
        RECT 11.410 58.940 16.820 59.110 ;
        RECT 19.015 59.110 19.185 59.855 ;
        RECT 20.385 59.810 20.615 60.330 ;
        RECT 21.345 59.810 21.575 60.330 ;
        RECT 22.305 59.810 22.535 60.330 ;
        RECT 23.265 59.810 23.495 60.330 ;
        RECT 24.225 59.810 24.455 60.330 ;
        RECT 19.855 59.655 20.185 59.670 ;
        RECT 19.840 59.395 20.200 59.655 ;
        RECT 19.855 59.370 20.185 59.395 ;
        RECT 20.415 59.110 20.585 59.810 ;
        RECT 20.815 59.655 21.145 59.670 ;
        RECT 20.795 59.395 21.155 59.655 ;
        RECT 20.815 59.370 21.145 59.395 ;
        RECT 21.375 59.110 21.545 59.810 ;
        RECT 21.775 59.655 22.105 59.670 ;
        RECT 21.755 59.395 22.115 59.655 ;
        RECT 21.775 59.370 22.105 59.395 ;
        RECT 22.335 59.110 22.505 59.810 ;
        RECT 22.735 59.655 23.065 59.670 ;
        RECT 22.715 59.395 23.075 59.655 ;
        RECT 22.735 59.370 23.065 59.395 ;
        RECT 23.295 59.110 23.465 59.810 ;
        RECT 23.695 59.650 24.025 59.670 ;
        RECT 23.680 59.390 24.040 59.650 ;
        RECT 23.695 59.370 24.025 59.390 ;
        RECT 24.255 59.110 24.425 59.810 ;
        RECT 24.655 59.650 24.985 59.670 ;
        RECT 24.640 59.390 25.000 59.650 ;
        RECT 24.655 59.370 24.985 59.390 ;
        RECT 19.015 58.940 24.425 59.110 ;
        RECT 11.410 57.545 16.820 57.715 ;
        RECT 1.535 55.415 1.765 56.775 ;
        RECT 2.495 55.415 2.725 56.775 ;
        RECT 3.455 55.415 3.685 56.775 ;
        RECT 4.415 55.415 4.645 56.775 ;
        RECT 5.375 55.415 5.605 56.775 ;
        RECT 6.335 55.415 6.565 56.775 ;
        RECT 1.565 54.710 1.735 55.415 ;
        RECT 2.525 54.710 2.695 55.415 ;
        RECT 3.485 54.710 3.655 55.415 ;
        RECT 4.445 54.710 4.615 55.415 ;
        RECT 5.405 54.710 5.575 55.415 ;
        RECT 6.365 54.710 6.535 55.415 ;
        RECT 11.410 54.730 11.580 57.545 ;
        RECT 12.810 56.795 12.980 57.545 ;
        RECT 13.770 56.795 13.940 57.545 ;
        RECT 14.730 56.795 14.900 57.545 ;
        RECT 15.690 56.795 15.860 57.545 ;
        RECT 16.650 56.795 16.820 57.545 ;
        RECT 19.015 57.545 24.425 57.715 ;
        RECT 12.300 55.435 12.530 56.795 ;
        RECT 12.780 55.435 13.010 56.795 ;
        RECT 13.260 55.435 13.490 56.795 ;
        RECT 13.740 55.435 13.970 56.795 ;
        RECT 14.220 55.435 14.450 56.795 ;
        RECT 14.700 55.435 14.930 56.795 ;
        RECT 15.180 55.435 15.410 56.795 ;
        RECT 15.660 55.435 15.890 56.795 ;
        RECT 16.140 55.435 16.370 56.795 ;
        RECT 16.620 55.435 16.850 56.795 ;
        RECT 17.100 55.435 17.330 56.795 ;
        RECT 10.505 54.710 11.580 54.730 ;
        RECT 1.565 54.560 11.580 54.710 ;
        RECT 1.565 54.540 10.705 54.560 ;
        RECT 1.565 53.875 1.735 54.540 ;
        RECT 2.525 53.875 2.695 54.540 ;
        RECT 3.485 53.875 3.655 54.540 ;
        RECT 4.445 53.875 4.615 54.540 ;
        RECT 5.405 53.875 5.575 54.540 ;
        RECT 6.365 53.875 6.535 54.540 ;
        RECT 1.535 53.355 1.765 53.875 ;
        RECT 2.495 53.355 2.725 53.875 ;
        RECT 3.455 53.355 3.685 53.875 ;
        RECT 4.415 53.355 4.645 53.875 ;
        RECT 5.375 53.355 5.605 53.875 ;
        RECT 6.335 53.355 6.565 53.875 ;
        RECT 11.410 52.675 11.580 54.560 ;
        RECT 12.330 54.730 12.500 55.435 ;
        RECT 13.290 54.730 13.460 55.435 ;
        RECT 14.250 54.730 14.420 55.435 ;
        RECT 15.210 54.730 15.380 55.435 ;
        RECT 16.170 54.730 16.340 55.435 ;
        RECT 17.130 54.730 17.300 55.435 ;
        RECT 19.015 54.730 19.185 57.545 ;
        RECT 20.415 56.795 20.585 57.545 ;
        RECT 21.375 56.795 21.545 57.545 ;
        RECT 22.335 56.795 22.505 57.545 ;
        RECT 23.295 56.795 23.465 57.545 ;
        RECT 24.255 56.795 24.425 57.545 ;
        RECT 20.385 55.435 20.615 56.795 ;
        RECT 21.345 55.435 21.575 56.795 ;
        RECT 22.305 55.435 22.535 56.795 ;
        RECT 23.265 55.435 23.495 56.795 ;
        RECT 24.225 55.435 24.455 56.795 ;
        RECT 12.330 54.560 19.185 54.730 ;
        RECT 12.330 53.895 12.500 54.560 ;
        RECT 13.290 53.895 13.460 54.560 ;
        RECT 14.250 53.895 14.420 54.560 ;
        RECT 15.210 53.895 15.380 54.560 ;
        RECT 16.170 53.895 16.340 54.560 ;
        RECT 17.130 53.895 17.300 54.560 ;
        RECT 19.015 53.920 19.185 54.560 ;
        RECT 26.630 54.265 27.000 54.535 ;
        RECT 18.670 53.915 19.185 53.920 ;
        RECT 12.300 53.375 12.530 53.895 ;
        RECT 12.780 53.375 13.010 53.895 ;
        RECT 13.260 53.375 13.490 53.895 ;
        RECT 13.740 53.375 13.970 53.895 ;
        RECT 14.220 53.375 14.450 53.895 ;
        RECT 14.700 53.375 14.930 53.895 ;
        RECT 15.180 53.375 15.410 53.895 ;
        RECT 15.660 53.375 15.890 53.895 ;
        RECT 16.140 53.375 16.370 53.895 ;
        RECT 16.620 53.375 16.850 53.895 ;
        RECT 17.100 53.375 17.330 53.895 ;
        RECT 18.645 53.420 19.185 53.915 ;
        RECT 18.645 53.415 18.875 53.420 ;
        RECT 12.250 53.220 12.580 53.235 ;
        RECT 12.235 52.960 12.595 53.220 ;
        RECT 12.250 52.935 12.580 52.960 ;
        RECT 12.810 52.675 12.980 53.375 ;
        RECT 13.210 53.220 13.540 53.235 ;
        RECT 13.190 52.960 13.550 53.220 ;
        RECT 13.210 52.935 13.540 52.960 ;
        RECT 13.770 52.675 13.940 53.375 ;
        RECT 14.170 53.220 14.500 53.235 ;
        RECT 14.150 52.960 14.510 53.220 ;
        RECT 14.170 52.935 14.500 52.960 ;
        RECT 14.730 52.675 14.900 53.375 ;
        RECT 15.130 53.220 15.460 53.235 ;
        RECT 15.110 52.960 15.470 53.220 ;
        RECT 15.130 52.935 15.460 52.960 ;
        RECT 15.690 52.675 15.860 53.375 ;
        RECT 16.090 53.215 16.420 53.235 ;
        RECT 16.075 52.955 16.435 53.215 ;
        RECT 16.090 52.935 16.420 52.955 ;
        RECT 16.650 52.675 16.820 53.375 ;
        RECT 17.050 53.215 17.380 53.235 ;
        RECT 17.035 52.955 17.395 53.215 ;
        RECT 17.050 52.935 17.380 52.955 ;
        RECT 11.410 52.505 16.820 52.675 ;
        RECT 19.015 52.675 19.185 53.420 ;
        RECT 20.385 53.375 20.615 53.895 ;
        RECT 21.345 53.375 21.575 53.895 ;
        RECT 22.305 53.375 22.535 53.895 ;
        RECT 23.265 53.375 23.495 53.895 ;
        RECT 24.225 53.375 24.455 53.895 ;
        RECT 19.855 53.220 20.185 53.235 ;
        RECT 19.840 52.960 20.200 53.220 ;
        RECT 19.855 52.935 20.185 52.960 ;
        RECT 20.415 52.675 20.585 53.375 ;
        RECT 20.815 53.220 21.145 53.235 ;
        RECT 20.795 52.960 21.155 53.220 ;
        RECT 20.815 52.935 21.145 52.960 ;
        RECT 21.375 52.675 21.545 53.375 ;
        RECT 21.775 53.220 22.105 53.235 ;
        RECT 21.755 52.960 22.115 53.220 ;
        RECT 21.775 52.935 22.105 52.960 ;
        RECT 22.335 52.675 22.505 53.375 ;
        RECT 22.735 53.220 23.065 53.235 ;
        RECT 22.715 52.960 23.075 53.220 ;
        RECT 22.735 52.935 23.065 52.960 ;
        RECT 23.295 52.675 23.465 53.375 ;
        RECT 23.695 53.215 24.025 53.235 ;
        RECT 23.680 52.955 24.040 53.215 ;
        RECT 23.695 52.935 24.025 52.955 ;
        RECT 24.255 52.675 24.425 53.375 ;
        RECT 24.655 53.215 24.985 53.235 ;
        RECT 24.640 52.955 25.000 53.215 ;
        RECT 24.655 52.935 24.985 52.955 ;
        RECT 19.015 52.505 24.425 52.675 ;
        RECT 11.410 51.110 16.820 51.280 ;
        RECT 1.535 48.980 1.765 50.340 ;
        RECT 2.495 48.980 2.725 50.340 ;
        RECT 3.455 48.980 3.685 50.340 ;
        RECT 4.415 48.980 4.645 50.340 ;
        RECT 5.375 48.980 5.605 50.340 ;
        RECT 6.335 48.980 6.565 50.340 ;
        RECT 1.565 48.275 1.735 48.980 ;
        RECT 2.525 48.275 2.695 48.980 ;
        RECT 3.485 48.275 3.655 48.980 ;
        RECT 4.445 48.275 4.615 48.980 ;
        RECT 5.405 48.275 5.575 48.980 ;
        RECT 6.365 48.275 6.535 48.980 ;
        RECT 11.410 48.295 11.580 51.110 ;
        RECT 12.810 50.360 12.980 51.110 ;
        RECT 13.770 50.360 13.940 51.110 ;
        RECT 14.730 50.360 14.900 51.110 ;
        RECT 15.690 50.360 15.860 51.110 ;
        RECT 16.650 50.360 16.820 51.110 ;
        RECT 19.015 51.110 24.425 51.280 ;
        RECT 12.300 49.000 12.530 50.360 ;
        RECT 12.780 49.000 13.010 50.360 ;
        RECT 13.260 49.000 13.490 50.360 ;
        RECT 13.740 49.000 13.970 50.360 ;
        RECT 14.220 49.000 14.450 50.360 ;
        RECT 14.700 49.000 14.930 50.360 ;
        RECT 15.180 49.000 15.410 50.360 ;
        RECT 15.660 49.000 15.890 50.360 ;
        RECT 16.140 49.000 16.370 50.360 ;
        RECT 16.620 49.000 16.850 50.360 ;
        RECT 17.100 49.000 17.330 50.360 ;
        RECT 10.505 48.275 11.580 48.295 ;
        RECT 1.565 48.125 11.580 48.275 ;
        RECT 1.565 48.105 10.705 48.125 ;
        RECT 1.565 47.440 1.735 48.105 ;
        RECT 2.525 47.440 2.695 48.105 ;
        RECT 3.485 47.440 3.655 48.105 ;
        RECT 4.445 47.440 4.615 48.105 ;
        RECT 5.405 47.440 5.575 48.105 ;
        RECT 6.365 47.440 6.535 48.105 ;
        RECT 1.535 46.920 1.765 47.440 ;
        RECT 2.495 46.920 2.725 47.440 ;
        RECT 3.455 46.920 3.685 47.440 ;
        RECT 4.415 46.920 4.645 47.440 ;
        RECT 5.375 46.920 5.605 47.440 ;
        RECT 6.335 46.920 6.565 47.440 ;
        RECT 11.410 46.240 11.580 48.125 ;
        RECT 12.330 48.295 12.500 49.000 ;
        RECT 13.290 48.295 13.460 49.000 ;
        RECT 14.250 48.295 14.420 49.000 ;
        RECT 15.210 48.295 15.380 49.000 ;
        RECT 16.170 48.295 16.340 49.000 ;
        RECT 17.130 48.295 17.300 49.000 ;
        RECT 19.015 48.295 19.185 51.110 ;
        RECT 20.415 50.360 20.585 51.110 ;
        RECT 21.375 50.360 21.545 51.110 ;
        RECT 22.335 50.360 22.505 51.110 ;
        RECT 23.295 50.360 23.465 51.110 ;
        RECT 24.255 50.360 24.425 51.110 ;
        RECT 20.385 49.000 20.615 50.360 ;
        RECT 21.345 49.000 21.575 50.360 ;
        RECT 22.305 49.000 22.535 50.360 ;
        RECT 23.265 49.000 23.495 50.360 ;
        RECT 24.225 49.000 24.455 50.360 ;
        RECT 12.330 48.125 19.185 48.295 ;
        RECT 12.330 47.460 12.500 48.125 ;
        RECT 13.290 47.460 13.460 48.125 ;
        RECT 14.250 47.460 14.420 48.125 ;
        RECT 15.210 47.460 15.380 48.125 ;
        RECT 16.170 47.460 16.340 48.125 ;
        RECT 17.130 47.460 17.300 48.125 ;
        RECT 19.015 47.485 19.185 48.125 ;
        RECT 26.630 47.830 27.000 48.100 ;
        RECT 18.670 47.480 19.185 47.485 ;
        RECT 12.300 46.940 12.530 47.460 ;
        RECT 12.780 46.940 13.010 47.460 ;
        RECT 13.260 46.940 13.490 47.460 ;
        RECT 13.740 46.940 13.970 47.460 ;
        RECT 14.220 46.940 14.450 47.460 ;
        RECT 14.700 46.940 14.930 47.460 ;
        RECT 15.180 46.940 15.410 47.460 ;
        RECT 15.660 46.940 15.890 47.460 ;
        RECT 16.140 46.940 16.370 47.460 ;
        RECT 16.620 46.940 16.850 47.460 ;
        RECT 17.100 46.940 17.330 47.460 ;
        RECT 18.645 46.985 19.185 47.480 ;
        RECT 18.645 46.980 18.875 46.985 ;
        RECT 12.250 46.785 12.580 46.800 ;
        RECT 12.235 46.525 12.595 46.785 ;
        RECT 12.250 46.500 12.580 46.525 ;
        RECT 12.810 46.240 12.980 46.940 ;
        RECT 13.210 46.785 13.540 46.800 ;
        RECT 13.190 46.525 13.550 46.785 ;
        RECT 13.210 46.500 13.540 46.525 ;
        RECT 13.770 46.240 13.940 46.940 ;
        RECT 14.170 46.785 14.500 46.800 ;
        RECT 14.150 46.525 14.510 46.785 ;
        RECT 14.170 46.500 14.500 46.525 ;
        RECT 14.730 46.240 14.900 46.940 ;
        RECT 15.130 46.785 15.460 46.800 ;
        RECT 15.110 46.525 15.470 46.785 ;
        RECT 15.130 46.500 15.460 46.525 ;
        RECT 15.690 46.240 15.860 46.940 ;
        RECT 16.090 46.780 16.420 46.800 ;
        RECT 16.075 46.520 16.435 46.780 ;
        RECT 16.090 46.500 16.420 46.520 ;
        RECT 16.650 46.240 16.820 46.940 ;
        RECT 17.050 46.780 17.380 46.800 ;
        RECT 17.035 46.520 17.395 46.780 ;
        RECT 17.050 46.500 17.380 46.520 ;
        RECT 11.410 46.070 16.820 46.240 ;
        RECT 19.015 46.240 19.185 46.985 ;
        RECT 20.385 46.940 20.615 47.460 ;
        RECT 21.345 46.940 21.575 47.460 ;
        RECT 22.305 46.940 22.535 47.460 ;
        RECT 23.265 46.940 23.495 47.460 ;
        RECT 24.225 46.940 24.455 47.460 ;
        RECT 19.855 46.785 20.185 46.800 ;
        RECT 19.840 46.525 20.200 46.785 ;
        RECT 19.855 46.500 20.185 46.525 ;
        RECT 20.415 46.240 20.585 46.940 ;
        RECT 20.815 46.785 21.145 46.800 ;
        RECT 20.795 46.525 21.155 46.785 ;
        RECT 20.815 46.500 21.145 46.525 ;
        RECT 21.375 46.240 21.545 46.940 ;
        RECT 21.775 46.785 22.105 46.800 ;
        RECT 21.755 46.525 22.115 46.785 ;
        RECT 21.775 46.500 22.105 46.525 ;
        RECT 22.335 46.240 22.505 46.940 ;
        RECT 22.735 46.785 23.065 46.800 ;
        RECT 22.715 46.525 23.075 46.785 ;
        RECT 22.735 46.500 23.065 46.525 ;
        RECT 23.295 46.240 23.465 46.940 ;
        RECT 23.695 46.780 24.025 46.800 ;
        RECT 23.680 46.520 24.040 46.780 ;
        RECT 23.695 46.500 24.025 46.520 ;
        RECT 24.255 46.240 24.425 46.940 ;
        RECT 24.655 46.780 24.985 46.800 ;
        RECT 24.640 46.520 25.000 46.780 ;
        RECT 24.655 46.500 24.985 46.520 ;
        RECT 19.015 46.070 24.425 46.240 ;
        RECT 11.410 44.675 16.820 44.845 ;
        RECT 1.535 42.545 1.765 43.905 ;
        RECT 2.495 42.545 2.725 43.905 ;
        RECT 3.455 42.545 3.685 43.905 ;
        RECT 4.415 42.545 4.645 43.905 ;
        RECT 5.375 42.545 5.605 43.905 ;
        RECT 6.335 42.545 6.565 43.905 ;
        RECT 1.565 41.840 1.735 42.545 ;
        RECT 2.525 41.840 2.695 42.545 ;
        RECT 3.485 41.840 3.655 42.545 ;
        RECT 4.445 41.840 4.615 42.545 ;
        RECT 5.405 41.840 5.575 42.545 ;
        RECT 6.365 41.840 6.535 42.545 ;
        RECT 11.410 41.860 11.580 44.675 ;
        RECT 12.810 43.925 12.980 44.675 ;
        RECT 13.770 43.925 13.940 44.675 ;
        RECT 14.730 43.925 14.900 44.675 ;
        RECT 15.690 43.925 15.860 44.675 ;
        RECT 16.650 43.925 16.820 44.675 ;
        RECT 19.015 44.675 24.425 44.845 ;
        RECT 12.300 42.565 12.530 43.925 ;
        RECT 12.780 42.565 13.010 43.925 ;
        RECT 13.260 42.565 13.490 43.925 ;
        RECT 13.740 42.565 13.970 43.925 ;
        RECT 14.220 42.565 14.450 43.925 ;
        RECT 14.700 42.565 14.930 43.925 ;
        RECT 15.180 42.565 15.410 43.925 ;
        RECT 15.660 42.565 15.890 43.925 ;
        RECT 16.140 42.565 16.370 43.925 ;
        RECT 16.620 42.565 16.850 43.925 ;
        RECT 17.100 42.565 17.330 43.925 ;
        RECT 10.505 41.840 11.580 41.860 ;
        RECT 1.565 41.690 11.580 41.840 ;
        RECT 1.565 41.670 10.705 41.690 ;
        RECT 1.565 41.005 1.735 41.670 ;
        RECT 2.525 41.005 2.695 41.670 ;
        RECT 3.485 41.005 3.655 41.670 ;
        RECT 4.445 41.005 4.615 41.670 ;
        RECT 5.405 41.005 5.575 41.670 ;
        RECT 6.365 41.005 6.535 41.670 ;
        RECT 1.535 40.485 1.765 41.005 ;
        RECT 2.495 40.485 2.725 41.005 ;
        RECT 3.455 40.485 3.685 41.005 ;
        RECT 4.415 40.485 4.645 41.005 ;
        RECT 5.375 40.485 5.605 41.005 ;
        RECT 6.335 40.485 6.565 41.005 ;
        RECT 11.410 39.805 11.580 41.690 ;
        RECT 12.330 41.860 12.500 42.565 ;
        RECT 13.290 41.860 13.460 42.565 ;
        RECT 14.250 41.860 14.420 42.565 ;
        RECT 15.210 41.860 15.380 42.565 ;
        RECT 16.170 41.860 16.340 42.565 ;
        RECT 17.130 41.860 17.300 42.565 ;
        RECT 19.015 41.860 19.185 44.675 ;
        RECT 20.415 43.925 20.585 44.675 ;
        RECT 21.375 43.925 21.545 44.675 ;
        RECT 22.335 43.925 22.505 44.675 ;
        RECT 23.295 43.925 23.465 44.675 ;
        RECT 24.255 43.925 24.425 44.675 ;
        RECT 20.385 42.565 20.615 43.925 ;
        RECT 21.345 42.565 21.575 43.925 ;
        RECT 22.305 42.565 22.535 43.925 ;
        RECT 23.265 42.565 23.495 43.925 ;
        RECT 24.225 42.565 24.455 43.925 ;
        RECT 12.330 41.690 19.185 41.860 ;
        RECT 12.330 41.025 12.500 41.690 ;
        RECT 13.290 41.025 13.460 41.690 ;
        RECT 14.250 41.025 14.420 41.690 ;
        RECT 15.210 41.025 15.380 41.690 ;
        RECT 16.170 41.025 16.340 41.690 ;
        RECT 17.130 41.025 17.300 41.690 ;
        RECT 19.015 41.050 19.185 41.690 ;
        RECT 26.630 41.395 27.000 41.665 ;
        RECT 18.670 41.045 19.185 41.050 ;
        RECT 12.300 40.505 12.530 41.025 ;
        RECT 12.780 40.505 13.010 41.025 ;
        RECT 13.260 40.505 13.490 41.025 ;
        RECT 13.740 40.505 13.970 41.025 ;
        RECT 14.220 40.505 14.450 41.025 ;
        RECT 14.700 40.505 14.930 41.025 ;
        RECT 15.180 40.505 15.410 41.025 ;
        RECT 15.660 40.505 15.890 41.025 ;
        RECT 16.140 40.505 16.370 41.025 ;
        RECT 16.620 40.505 16.850 41.025 ;
        RECT 17.100 40.505 17.330 41.025 ;
        RECT 18.645 40.550 19.185 41.045 ;
        RECT 18.645 40.545 18.875 40.550 ;
        RECT 12.250 40.350 12.580 40.365 ;
        RECT 12.235 40.090 12.595 40.350 ;
        RECT 12.250 40.065 12.580 40.090 ;
        RECT 12.810 39.805 12.980 40.505 ;
        RECT 13.210 40.350 13.540 40.365 ;
        RECT 13.190 40.090 13.550 40.350 ;
        RECT 13.210 40.065 13.540 40.090 ;
        RECT 13.770 39.805 13.940 40.505 ;
        RECT 14.170 40.350 14.500 40.365 ;
        RECT 14.150 40.090 14.510 40.350 ;
        RECT 14.170 40.065 14.500 40.090 ;
        RECT 14.730 39.805 14.900 40.505 ;
        RECT 15.130 40.350 15.460 40.365 ;
        RECT 15.110 40.090 15.470 40.350 ;
        RECT 15.130 40.065 15.460 40.090 ;
        RECT 15.690 39.805 15.860 40.505 ;
        RECT 16.090 40.345 16.420 40.365 ;
        RECT 16.075 40.085 16.435 40.345 ;
        RECT 16.090 40.065 16.420 40.085 ;
        RECT 16.650 39.805 16.820 40.505 ;
        RECT 17.050 40.345 17.380 40.365 ;
        RECT 17.035 40.085 17.395 40.345 ;
        RECT 17.050 40.065 17.380 40.085 ;
        RECT 11.410 39.635 16.820 39.805 ;
        RECT 19.015 39.805 19.185 40.550 ;
        RECT 20.385 40.505 20.615 41.025 ;
        RECT 21.345 40.505 21.575 41.025 ;
        RECT 22.305 40.505 22.535 41.025 ;
        RECT 23.265 40.505 23.495 41.025 ;
        RECT 24.225 40.505 24.455 41.025 ;
        RECT 19.855 40.350 20.185 40.365 ;
        RECT 19.840 40.090 20.200 40.350 ;
        RECT 19.855 40.065 20.185 40.090 ;
        RECT 20.415 39.805 20.585 40.505 ;
        RECT 20.815 40.350 21.145 40.365 ;
        RECT 20.795 40.090 21.155 40.350 ;
        RECT 20.815 40.065 21.145 40.090 ;
        RECT 21.375 39.805 21.545 40.505 ;
        RECT 21.775 40.350 22.105 40.365 ;
        RECT 21.755 40.090 22.115 40.350 ;
        RECT 21.775 40.065 22.105 40.090 ;
        RECT 22.335 39.805 22.505 40.505 ;
        RECT 22.735 40.350 23.065 40.365 ;
        RECT 22.715 40.090 23.075 40.350 ;
        RECT 22.735 40.065 23.065 40.090 ;
        RECT 23.295 39.805 23.465 40.505 ;
        RECT 23.695 40.345 24.025 40.365 ;
        RECT 23.680 40.085 24.040 40.345 ;
        RECT 23.695 40.065 24.025 40.085 ;
        RECT 24.255 39.805 24.425 40.505 ;
        RECT 24.655 40.345 24.985 40.365 ;
        RECT 24.640 40.085 25.000 40.345 ;
        RECT 24.655 40.065 24.985 40.085 ;
        RECT 19.015 39.635 24.425 39.805 ;
        RECT 11.410 38.240 16.820 38.410 ;
        RECT 1.535 36.110 1.765 37.470 ;
        RECT 2.495 36.110 2.725 37.470 ;
        RECT 3.455 36.110 3.685 37.470 ;
        RECT 4.415 36.110 4.645 37.470 ;
        RECT 5.375 36.110 5.605 37.470 ;
        RECT 6.335 36.110 6.565 37.470 ;
        RECT 1.565 35.405 1.735 36.110 ;
        RECT 2.525 35.405 2.695 36.110 ;
        RECT 3.485 35.405 3.655 36.110 ;
        RECT 4.445 35.405 4.615 36.110 ;
        RECT 5.405 35.405 5.575 36.110 ;
        RECT 6.365 35.405 6.535 36.110 ;
        RECT 11.410 35.425 11.580 38.240 ;
        RECT 12.810 37.490 12.980 38.240 ;
        RECT 13.770 37.490 13.940 38.240 ;
        RECT 14.730 37.490 14.900 38.240 ;
        RECT 15.690 37.490 15.860 38.240 ;
        RECT 16.650 37.490 16.820 38.240 ;
        RECT 19.015 38.240 24.425 38.410 ;
        RECT 12.300 36.130 12.530 37.490 ;
        RECT 12.780 36.130 13.010 37.490 ;
        RECT 13.260 36.130 13.490 37.490 ;
        RECT 13.740 36.130 13.970 37.490 ;
        RECT 14.220 36.130 14.450 37.490 ;
        RECT 14.700 36.130 14.930 37.490 ;
        RECT 15.180 36.130 15.410 37.490 ;
        RECT 15.660 36.130 15.890 37.490 ;
        RECT 16.140 36.130 16.370 37.490 ;
        RECT 16.620 36.130 16.850 37.490 ;
        RECT 17.100 36.130 17.330 37.490 ;
        RECT 10.505 35.405 11.580 35.425 ;
        RECT 1.565 35.255 11.580 35.405 ;
        RECT 1.565 35.235 10.705 35.255 ;
        RECT 1.565 34.570 1.735 35.235 ;
        RECT 2.525 34.570 2.695 35.235 ;
        RECT 3.485 34.570 3.655 35.235 ;
        RECT 4.445 34.570 4.615 35.235 ;
        RECT 5.405 34.570 5.575 35.235 ;
        RECT 6.365 34.570 6.535 35.235 ;
        RECT 1.535 34.050 1.765 34.570 ;
        RECT 2.495 34.050 2.725 34.570 ;
        RECT 3.455 34.050 3.685 34.570 ;
        RECT 4.415 34.050 4.645 34.570 ;
        RECT 5.375 34.050 5.605 34.570 ;
        RECT 6.335 34.050 6.565 34.570 ;
        RECT 11.410 33.370 11.580 35.255 ;
        RECT 12.330 35.425 12.500 36.130 ;
        RECT 13.290 35.425 13.460 36.130 ;
        RECT 14.250 35.425 14.420 36.130 ;
        RECT 15.210 35.425 15.380 36.130 ;
        RECT 16.170 35.425 16.340 36.130 ;
        RECT 17.130 35.425 17.300 36.130 ;
        RECT 19.015 35.425 19.185 38.240 ;
        RECT 20.415 37.490 20.585 38.240 ;
        RECT 21.375 37.490 21.545 38.240 ;
        RECT 22.335 37.490 22.505 38.240 ;
        RECT 23.295 37.490 23.465 38.240 ;
        RECT 24.255 37.490 24.425 38.240 ;
        RECT 20.385 36.130 20.615 37.490 ;
        RECT 21.345 36.130 21.575 37.490 ;
        RECT 22.305 36.130 22.535 37.490 ;
        RECT 23.265 36.130 23.495 37.490 ;
        RECT 24.225 36.130 24.455 37.490 ;
        RECT 12.330 35.255 19.185 35.425 ;
        RECT 12.330 34.590 12.500 35.255 ;
        RECT 13.290 34.590 13.460 35.255 ;
        RECT 14.250 34.590 14.420 35.255 ;
        RECT 15.210 34.590 15.380 35.255 ;
        RECT 16.170 34.590 16.340 35.255 ;
        RECT 17.130 34.590 17.300 35.255 ;
        RECT 19.015 34.615 19.185 35.255 ;
        RECT 26.630 34.960 27.000 35.230 ;
        RECT 18.670 34.610 19.185 34.615 ;
        RECT 12.300 34.070 12.530 34.590 ;
        RECT 12.780 34.070 13.010 34.590 ;
        RECT 13.260 34.070 13.490 34.590 ;
        RECT 13.740 34.070 13.970 34.590 ;
        RECT 14.220 34.070 14.450 34.590 ;
        RECT 14.700 34.070 14.930 34.590 ;
        RECT 15.180 34.070 15.410 34.590 ;
        RECT 15.660 34.070 15.890 34.590 ;
        RECT 16.140 34.070 16.370 34.590 ;
        RECT 16.620 34.070 16.850 34.590 ;
        RECT 17.100 34.070 17.330 34.590 ;
        RECT 18.645 34.115 19.185 34.610 ;
        RECT 18.645 34.110 18.875 34.115 ;
        RECT 12.250 33.915 12.580 33.930 ;
        RECT 12.235 33.655 12.595 33.915 ;
        RECT 12.250 33.630 12.580 33.655 ;
        RECT 12.810 33.370 12.980 34.070 ;
        RECT 13.210 33.915 13.540 33.930 ;
        RECT 13.190 33.655 13.550 33.915 ;
        RECT 13.210 33.630 13.540 33.655 ;
        RECT 13.770 33.370 13.940 34.070 ;
        RECT 14.170 33.915 14.500 33.930 ;
        RECT 14.150 33.655 14.510 33.915 ;
        RECT 14.170 33.630 14.500 33.655 ;
        RECT 14.730 33.370 14.900 34.070 ;
        RECT 15.130 33.915 15.460 33.930 ;
        RECT 15.110 33.655 15.470 33.915 ;
        RECT 15.130 33.630 15.460 33.655 ;
        RECT 15.690 33.370 15.860 34.070 ;
        RECT 16.090 33.910 16.420 33.930 ;
        RECT 16.075 33.650 16.435 33.910 ;
        RECT 16.090 33.630 16.420 33.650 ;
        RECT 16.650 33.370 16.820 34.070 ;
        RECT 17.050 33.910 17.380 33.930 ;
        RECT 17.035 33.650 17.395 33.910 ;
        RECT 17.050 33.630 17.380 33.650 ;
        RECT 11.410 33.200 16.820 33.370 ;
        RECT 19.015 33.370 19.185 34.115 ;
        RECT 20.385 34.070 20.615 34.590 ;
        RECT 21.345 34.070 21.575 34.590 ;
        RECT 22.305 34.070 22.535 34.590 ;
        RECT 23.265 34.070 23.495 34.590 ;
        RECT 24.225 34.070 24.455 34.590 ;
        RECT 19.855 33.915 20.185 33.930 ;
        RECT 19.840 33.655 20.200 33.915 ;
        RECT 19.855 33.630 20.185 33.655 ;
        RECT 20.415 33.370 20.585 34.070 ;
        RECT 20.815 33.915 21.145 33.930 ;
        RECT 20.795 33.655 21.155 33.915 ;
        RECT 20.815 33.630 21.145 33.655 ;
        RECT 21.375 33.370 21.545 34.070 ;
        RECT 21.775 33.915 22.105 33.930 ;
        RECT 21.755 33.655 22.115 33.915 ;
        RECT 21.775 33.630 22.105 33.655 ;
        RECT 22.335 33.370 22.505 34.070 ;
        RECT 22.735 33.915 23.065 33.930 ;
        RECT 22.715 33.655 23.075 33.915 ;
        RECT 22.735 33.630 23.065 33.655 ;
        RECT 23.295 33.370 23.465 34.070 ;
        RECT 23.695 33.910 24.025 33.930 ;
        RECT 23.680 33.650 24.040 33.910 ;
        RECT 23.695 33.630 24.025 33.650 ;
        RECT 24.255 33.370 24.425 34.070 ;
        RECT 24.655 33.910 24.985 33.930 ;
        RECT 24.640 33.650 25.000 33.910 ;
        RECT 24.655 33.630 24.985 33.650 ;
        RECT 19.015 33.200 24.425 33.370 ;
        RECT 11.410 31.805 16.820 31.975 ;
        RECT 1.535 29.675 1.765 31.035 ;
        RECT 2.495 29.675 2.725 31.035 ;
        RECT 3.455 29.675 3.685 31.035 ;
        RECT 4.415 29.675 4.645 31.035 ;
        RECT 5.375 29.675 5.605 31.035 ;
        RECT 6.335 29.675 6.565 31.035 ;
        RECT 1.565 28.970 1.735 29.675 ;
        RECT 2.525 28.970 2.695 29.675 ;
        RECT 3.485 28.970 3.655 29.675 ;
        RECT 4.445 28.970 4.615 29.675 ;
        RECT 5.405 28.970 5.575 29.675 ;
        RECT 6.365 28.970 6.535 29.675 ;
        RECT 11.410 28.990 11.580 31.805 ;
        RECT 12.810 31.055 12.980 31.805 ;
        RECT 13.770 31.055 13.940 31.805 ;
        RECT 14.730 31.055 14.900 31.805 ;
        RECT 15.690 31.055 15.860 31.805 ;
        RECT 16.650 31.055 16.820 31.805 ;
        RECT 19.015 31.805 24.425 31.975 ;
        RECT 12.300 29.695 12.530 31.055 ;
        RECT 12.780 29.695 13.010 31.055 ;
        RECT 13.260 29.695 13.490 31.055 ;
        RECT 13.740 29.695 13.970 31.055 ;
        RECT 14.220 29.695 14.450 31.055 ;
        RECT 14.700 29.695 14.930 31.055 ;
        RECT 15.180 29.695 15.410 31.055 ;
        RECT 15.660 29.695 15.890 31.055 ;
        RECT 16.140 29.695 16.370 31.055 ;
        RECT 16.620 29.695 16.850 31.055 ;
        RECT 17.100 29.695 17.330 31.055 ;
        RECT 10.505 28.970 11.580 28.990 ;
        RECT 1.565 28.820 11.580 28.970 ;
        RECT 1.565 28.800 10.705 28.820 ;
        RECT 1.565 28.135 1.735 28.800 ;
        RECT 2.525 28.135 2.695 28.800 ;
        RECT 3.485 28.135 3.655 28.800 ;
        RECT 4.445 28.135 4.615 28.800 ;
        RECT 5.405 28.135 5.575 28.800 ;
        RECT 6.365 28.135 6.535 28.800 ;
        RECT 1.535 27.615 1.765 28.135 ;
        RECT 2.495 27.615 2.725 28.135 ;
        RECT 3.455 27.615 3.685 28.135 ;
        RECT 4.415 27.615 4.645 28.135 ;
        RECT 5.375 27.615 5.605 28.135 ;
        RECT 6.335 27.615 6.565 28.135 ;
        RECT 11.410 26.935 11.580 28.820 ;
        RECT 12.330 28.990 12.500 29.695 ;
        RECT 13.290 28.990 13.460 29.695 ;
        RECT 14.250 28.990 14.420 29.695 ;
        RECT 15.210 28.990 15.380 29.695 ;
        RECT 16.170 28.990 16.340 29.695 ;
        RECT 17.130 28.990 17.300 29.695 ;
        RECT 19.015 28.990 19.185 31.805 ;
        RECT 20.415 31.055 20.585 31.805 ;
        RECT 21.375 31.055 21.545 31.805 ;
        RECT 22.335 31.055 22.505 31.805 ;
        RECT 23.295 31.055 23.465 31.805 ;
        RECT 24.255 31.055 24.425 31.805 ;
        RECT 20.385 29.695 20.615 31.055 ;
        RECT 21.345 29.695 21.575 31.055 ;
        RECT 22.305 29.695 22.535 31.055 ;
        RECT 23.265 29.695 23.495 31.055 ;
        RECT 24.225 29.695 24.455 31.055 ;
        RECT 12.330 28.820 19.185 28.990 ;
        RECT 12.330 28.155 12.500 28.820 ;
        RECT 13.290 28.155 13.460 28.820 ;
        RECT 14.250 28.155 14.420 28.820 ;
        RECT 15.210 28.155 15.380 28.820 ;
        RECT 16.170 28.155 16.340 28.820 ;
        RECT 17.130 28.155 17.300 28.820 ;
        RECT 19.015 28.180 19.185 28.820 ;
        RECT 26.630 28.525 27.000 28.795 ;
        RECT 18.670 28.175 19.185 28.180 ;
        RECT 12.300 27.635 12.530 28.155 ;
        RECT 12.780 27.635 13.010 28.155 ;
        RECT 13.260 27.635 13.490 28.155 ;
        RECT 13.740 27.635 13.970 28.155 ;
        RECT 14.220 27.635 14.450 28.155 ;
        RECT 14.700 27.635 14.930 28.155 ;
        RECT 15.180 27.635 15.410 28.155 ;
        RECT 15.660 27.635 15.890 28.155 ;
        RECT 16.140 27.635 16.370 28.155 ;
        RECT 16.620 27.635 16.850 28.155 ;
        RECT 17.100 27.635 17.330 28.155 ;
        RECT 18.645 27.680 19.185 28.175 ;
        RECT 18.645 27.675 18.875 27.680 ;
        RECT 12.250 27.480 12.580 27.495 ;
        RECT 12.235 27.220 12.595 27.480 ;
        RECT 12.250 27.195 12.580 27.220 ;
        RECT 12.810 26.935 12.980 27.635 ;
        RECT 13.210 27.480 13.540 27.495 ;
        RECT 13.190 27.220 13.550 27.480 ;
        RECT 13.210 27.195 13.540 27.220 ;
        RECT 13.770 26.935 13.940 27.635 ;
        RECT 14.170 27.480 14.500 27.495 ;
        RECT 14.150 27.220 14.510 27.480 ;
        RECT 14.170 27.195 14.500 27.220 ;
        RECT 14.730 26.935 14.900 27.635 ;
        RECT 15.130 27.480 15.460 27.495 ;
        RECT 15.110 27.220 15.470 27.480 ;
        RECT 15.130 27.195 15.460 27.220 ;
        RECT 15.690 26.935 15.860 27.635 ;
        RECT 16.090 27.475 16.420 27.495 ;
        RECT 16.075 27.215 16.435 27.475 ;
        RECT 16.090 27.195 16.420 27.215 ;
        RECT 16.650 26.935 16.820 27.635 ;
        RECT 17.050 27.475 17.380 27.495 ;
        RECT 17.035 27.215 17.395 27.475 ;
        RECT 17.050 27.195 17.380 27.215 ;
        RECT 11.410 26.765 16.820 26.935 ;
        RECT 19.015 26.935 19.185 27.680 ;
        RECT 20.385 27.635 20.615 28.155 ;
        RECT 21.345 27.635 21.575 28.155 ;
        RECT 22.305 27.635 22.535 28.155 ;
        RECT 23.265 27.635 23.495 28.155 ;
        RECT 24.225 27.635 24.455 28.155 ;
        RECT 19.855 27.480 20.185 27.495 ;
        RECT 19.840 27.220 20.200 27.480 ;
        RECT 19.855 27.195 20.185 27.220 ;
        RECT 20.415 26.935 20.585 27.635 ;
        RECT 20.815 27.480 21.145 27.495 ;
        RECT 20.795 27.220 21.155 27.480 ;
        RECT 20.815 27.195 21.145 27.220 ;
        RECT 21.375 26.935 21.545 27.635 ;
        RECT 21.775 27.480 22.105 27.495 ;
        RECT 21.755 27.220 22.115 27.480 ;
        RECT 21.775 27.195 22.105 27.220 ;
        RECT 22.335 26.935 22.505 27.635 ;
        RECT 22.735 27.480 23.065 27.495 ;
        RECT 22.715 27.220 23.075 27.480 ;
        RECT 22.735 27.195 23.065 27.220 ;
        RECT 23.295 26.935 23.465 27.635 ;
        RECT 23.695 27.475 24.025 27.495 ;
        RECT 23.680 27.215 24.040 27.475 ;
        RECT 23.695 27.195 24.025 27.215 ;
        RECT 24.255 26.935 24.425 27.635 ;
        RECT 24.655 27.475 24.985 27.495 ;
        RECT 24.640 27.215 25.000 27.475 ;
        RECT 24.655 27.195 24.985 27.215 ;
        RECT 19.015 26.765 24.425 26.935 ;
        RECT 11.410 25.370 16.820 25.540 ;
        RECT 1.535 23.240 1.765 24.600 ;
        RECT 2.495 23.240 2.725 24.600 ;
        RECT 3.455 23.240 3.685 24.600 ;
        RECT 4.415 23.240 4.645 24.600 ;
        RECT 5.375 23.240 5.605 24.600 ;
        RECT 6.335 23.240 6.565 24.600 ;
        RECT 1.565 22.535 1.735 23.240 ;
        RECT 2.525 22.535 2.695 23.240 ;
        RECT 3.485 22.535 3.655 23.240 ;
        RECT 4.445 22.535 4.615 23.240 ;
        RECT 5.405 22.535 5.575 23.240 ;
        RECT 6.365 22.535 6.535 23.240 ;
        RECT 11.410 22.555 11.580 25.370 ;
        RECT 12.810 24.620 12.980 25.370 ;
        RECT 13.770 24.620 13.940 25.370 ;
        RECT 14.730 24.620 14.900 25.370 ;
        RECT 15.690 24.620 15.860 25.370 ;
        RECT 16.650 24.620 16.820 25.370 ;
        RECT 19.015 25.370 24.425 25.540 ;
        RECT 12.300 23.260 12.530 24.620 ;
        RECT 12.780 23.260 13.010 24.620 ;
        RECT 13.260 23.260 13.490 24.620 ;
        RECT 13.740 23.260 13.970 24.620 ;
        RECT 14.220 23.260 14.450 24.620 ;
        RECT 14.700 23.260 14.930 24.620 ;
        RECT 15.180 23.260 15.410 24.620 ;
        RECT 15.660 23.260 15.890 24.620 ;
        RECT 16.140 23.260 16.370 24.620 ;
        RECT 16.620 23.260 16.850 24.620 ;
        RECT 17.100 23.260 17.330 24.620 ;
        RECT 10.505 22.535 11.580 22.555 ;
        RECT 1.565 22.385 11.580 22.535 ;
        RECT 1.565 22.365 10.705 22.385 ;
        RECT 1.565 21.700 1.735 22.365 ;
        RECT 2.525 21.700 2.695 22.365 ;
        RECT 3.485 21.700 3.655 22.365 ;
        RECT 4.445 21.700 4.615 22.365 ;
        RECT 5.405 21.700 5.575 22.365 ;
        RECT 6.365 21.700 6.535 22.365 ;
        RECT 1.535 21.180 1.765 21.700 ;
        RECT 2.495 21.180 2.725 21.700 ;
        RECT 3.455 21.180 3.685 21.700 ;
        RECT 4.415 21.180 4.645 21.700 ;
        RECT 5.375 21.180 5.605 21.700 ;
        RECT 6.335 21.180 6.565 21.700 ;
        RECT 11.410 20.500 11.580 22.385 ;
        RECT 12.330 22.555 12.500 23.260 ;
        RECT 13.290 22.555 13.460 23.260 ;
        RECT 14.250 22.555 14.420 23.260 ;
        RECT 15.210 22.555 15.380 23.260 ;
        RECT 16.170 22.555 16.340 23.260 ;
        RECT 17.130 22.555 17.300 23.260 ;
        RECT 19.015 22.555 19.185 25.370 ;
        RECT 20.415 24.620 20.585 25.370 ;
        RECT 21.375 24.620 21.545 25.370 ;
        RECT 22.335 24.620 22.505 25.370 ;
        RECT 23.295 24.620 23.465 25.370 ;
        RECT 24.255 24.620 24.425 25.370 ;
        RECT 20.385 23.260 20.615 24.620 ;
        RECT 21.345 23.260 21.575 24.620 ;
        RECT 22.305 23.260 22.535 24.620 ;
        RECT 23.265 23.260 23.495 24.620 ;
        RECT 24.225 23.260 24.455 24.620 ;
        RECT 12.330 22.385 19.185 22.555 ;
        RECT 12.330 21.720 12.500 22.385 ;
        RECT 13.290 21.720 13.460 22.385 ;
        RECT 14.250 21.720 14.420 22.385 ;
        RECT 15.210 21.720 15.380 22.385 ;
        RECT 16.170 21.720 16.340 22.385 ;
        RECT 17.130 21.720 17.300 22.385 ;
        RECT 19.015 21.745 19.185 22.385 ;
        RECT 26.630 22.090 27.000 22.360 ;
        RECT 18.670 21.740 19.185 21.745 ;
        RECT 12.300 21.200 12.530 21.720 ;
        RECT 12.780 21.200 13.010 21.720 ;
        RECT 13.260 21.200 13.490 21.720 ;
        RECT 13.740 21.200 13.970 21.720 ;
        RECT 14.220 21.200 14.450 21.720 ;
        RECT 14.700 21.200 14.930 21.720 ;
        RECT 15.180 21.200 15.410 21.720 ;
        RECT 15.660 21.200 15.890 21.720 ;
        RECT 16.140 21.200 16.370 21.720 ;
        RECT 16.620 21.200 16.850 21.720 ;
        RECT 17.100 21.200 17.330 21.720 ;
        RECT 18.645 21.245 19.185 21.740 ;
        RECT 18.645 21.240 18.875 21.245 ;
        RECT 12.250 21.045 12.580 21.060 ;
        RECT 12.235 20.785 12.595 21.045 ;
        RECT 12.250 20.760 12.580 20.785 ;
        RECT 12.810 20.500 12.980 21.200 ;
        RECT 13.210 21.045 13.540 21.060 ;
        RECT 13.190 20.785 13.550 21.045 ;
        RECT 13.210 20.760 13.540 20.785 ;
        RECT 13.770 20.500 13.940 21.200 ;
        RECT 14.170 21.045 14.500 21.060 ;
        RECT 14.150 20.785 14.510 21.045 ;
        RECT 14.170 20.760 14.500 20.785 ;
        RECT 14.730 20.500 14.900 21.200 ;
        RECT 15.130 21.045 15.460 21.060 ;
        RECT 15.110 20.785 15.470 21.045 ;
        RECT 15.130 20.760 15.460 20.785 ;
        RECT 15.690 20.500 15.860 21.200 ;
        RECT 16.090 21.040 16.420 21.060 ;
        RECT 16.075 20.780 16.435 21.040 ;
        RECT 16.090 20.760 16.420 20.780 ;
        RECT 16.650 20.500 16.820 21.200 ;
        RECT 17.050 21.040 17.380 21.060 ;
        RECT 17.035 20.780 17.395 21.040 ;
        RECT 17.050 20.760 17.380 20.780 ;
        RECT 11.410 20.330 16.820 20.500 ;
        RECT 19.015 20.500 19.185 21.245 ;
        RECT 20.385 21.200 20.615 21.720 ;
        RECT 21.345 21.200 21.575 21.720 ;
        RECT 22.305 21.200 22.535 21.720 ;
        RECT 23.265 21.200 23.495 21.720 ;
        RECT 24.225 21.200 24.455 21.720 ;
        RECT 19.855 21.045 20.185 21.060 ;
        RECT 19.840 20.785 20.200 21.045 ;
        RECT 19.855 20.760 20.185 20.785 ;
        RECT 20.415 20.500 20.585 21.200 ;
        RECT 20.815 21.045 21.145 21.060 ;
        RECT 20.795 20.785 21.155 21.045 ;
        RECT 20.815 20.760 21.145 20.785 ;
        RECT 21.375 20.500 21.545 21.200 ;
        RECT 21.775 21.045 22.105 21.060 ;
        RECT 21.755 20.785 22.115 21.045 ;
        RECT 21.775 20.760 22.105 20.785 ;
        RECT 22.335 20.500 22.505 21.200 ;
        RECT 22.735 21.045 23.065 21.060 ;
        RECT 22.715 20.785 23.075 21.045 ;
        RECT 22.735 20.760 23.065 20.785 ;
        RECT 23.295 20.500 23.465 21.200 ;
        RECT 23.695 21.040 24.025 21.060 ;
        RECT 23.680 20.780 24.040 21.040 ;
        RECT 23.695 20.760 24.025 20.780 ;
        RECT 24.255 20.500 24.425 21.200 ;
        RECT 24.655 21.040 24.985 21.060 ;
        RECT 24.640 20.780 25.000 21.040 ;
        RECT 24.655 20.760 24.985 20.780 ;
        RECT 19.015 20.330 24.425 20.500 ;
        RECT 11.410 18.935 16.820 19.105 ;
        RECT 1.535 16.805 1.765 18.165 ;
        RECT 2.495 16.805 2.725 18.165 ;
        RECT 3.455 16.805 3.685 18.165 ;
        RECT 4.415 16.805 4.645 18.165 ;
        RECT 5.375 16.805 5.605 18.165 ;
        RECT 6.335 16.805 6.565 18.165 ;
        RECT 1.565 16.100 1.735 16.805 ;
        RECT 2.525 16.100 2.695 16.805 ;
        RECT 3.485 16.100 3.655 16.805 ;
        RECT 4.445 16.100 4.615 16.805 ;
        RECT 5.405 16.100 5.575 16.805 ;
        RECT 6.365 16.100 6.535 16.805 ;
        RECT 11.410 16.120 11.580 18.935 ;
        RECT 12.810 18.185 12.980 18.935 ;
        RECT 13.770 18.185 13.940 18.935 ;
        RECT 14.730 18.185 14.900 18.935 ;
        RECT 15.690 18.185 15.860 18.935 ;
        RECT 16.650 18.185 16.820 18.935 ;
        RECT 19.015 18.935 24.425 19.105 ;
        RECT 12.300 16.825 12.530 18.185 ;
        RECT 12.780 16.825 13.010 18.185 ;
        RECT 13.260 16.825 13.490 18.185 ;
        RECT 13.740 16.825 13.970 18.185 ;
        RECT 14.220 16.825 14.450 18.185 ;
        RECT 14.700 16.825 14.930 18.185 ;
        RECT 15.180 16.825 15.410 18.185 ;
        RECT 15.660 16.825 15.890 18.185 ;
        RECT 16.140 16.825 16.370 18.185 ;
        RECT 16.620 16.825 16.850 18.185 ;
        RECT 17.100 16.825 17.330 18.185 ;
        RECT 10.505 16.100 11.580 16.120 ;
        RECT 1.565 15.950 11.580 16.100 ;
        RECT 1.565 15.930 10.705 15.950 ;
        RECT 1.565 15.265 1.735 15.930 ;
        RECT 2.525 15.265 2.695 15.930 ;
        RECT 3.485 15.265 3.655 15.930 ;
        RECT 4.445 15.265 4.615 15.930 ;
        RECT 5.405 15.265 5.575 15.930 ;
        RECT 6.365 15.265 6.535 15.930 ;
        RECT 1.535 14.745 1.765 15.265 ;
        RECT 2.495 14.745 2.725 15.265 ;
        RECT 3.455 14.745 3.685 15.265 ;
        RECT 4.415 14.745 4.645 15.265 ;
        RECT 5.375 14.745 5.605 15.265 ;
        RECT 6.335 14.745 6.565 15.265 ;
        RECT 11.410 14.065 11.580 15.950 ;
        RECT 12.330 16.120 12.500 16.825 ;
        RECT 13.290 16.120 13.460 16.825 ;
        RECT 14.250 16.120 14.420 16.825 ;
        RECT 15.210 16.120 15.380 16.825 ;
        RECT 16.170 16.120 16.340 16.825 ;
        RECT 17.130 16.120 17.300 16.825 ;
        RECT 19.015 16.120 19.185 18.935 ;
        RECT 20.415 18.185 20.585 18.935 ;
        RECT 21.375 18.185 21.545 18.935 ;
        RECT 22.335 18.185 22.505 18.935 ;
        RECT 23.295 18.185 23.465 18.935 ;
        RECT 24.255 18.185 24.425 18.935 ;
        RECT 20.385 16.825 20.615 18.185 ;
        RECT 21.345 16.825 21.575 18.185 ;
        RECT 22.305 16.825 22.535 18.185 ;
        RECT 23.265 16.825 23.495 18.185 ;
        RECT 24.225 16.825 24.455 18.185 ;
        RECT 12.330 15.950 19.185 16.120 ;
        RECT 12.330 15.285 12.500 15.950 ;
        RECT 13.290 15.285 13.460 15.950 ;
        RECT 14.250 15.285 14.420 15.950 ;
        RECT 15.210 15.285 15.380 15.950 ;
        RECT 16.170 15.285 16.340 15.950 ;
        RECT 17.130 15.285 17.300 15.950 ;
        RECT 19.015 15.310 19.185 15.950 ;
        RECT 26.630 15.655 27.000 15.925 ;
        RECT 18.670 15.305 19.185 15.310 ;
        RECT 12.300 14.765 12.530 15.285 ;
        RECT 12.780 14.765 13.010 15.285 ;
        RECT 13.260 14.765 13.490 15.285 ;
        RECT 13.740 14.765 13.970 15.285 ;
        RECT 14.220 14.765 14.450 15.285 ;
        RECT 14.700 14.765 14.930 15.285 ;
        RECT 15.180 14.765 15.410 15.285 ;
        RECT 15.660 14.765 15.890 15.285 ;
        RECT 16.140 14.765 16.370 15.285 ;
        RECT 16.620 14.765 16.850 15.285 ;
        RECT 17.100 14.765 17.330 15.285 ;
        RECT 18.645 14.810 19.185 15.305 ;
        RECT 18.645 14.805 18.875 14.810 ;
        RECT 12.250 14.610 12.580 14.625 ;
        RECT 12.235 14.350 12.595 14.610 ;
        RECT 12.250 14.325 12.580 14.350 ;
        RECT 12.810 14.065 12.980 14.765 ;
        RECT 13.210 14.610 13.540 14.625 ;
        RECT 13.190 14.350 13.550 14.610 ;
        RECT 13.210 14.325 13.540 14.350 ;
        RECT 13.770 14.065 13.940 14.765 ;
        RECT 14.170 14.610 14.500 14.625 ;
        RECT 14.150 14.350 14.510 14.610 ;
        RECT 14.170 14.325 14.500 14.350 ;
        RECT 14.730 14.065 14.900 14.765 ;
        RECT 15.130 14.610 15.460 14.625 ;
        RECT 15.110 14.350 15.470 14.610 ;
        RECT 15.130 14.325 15.460 14.350 ;
        RECT 15.690 14.065 15.860 14.765 ;
        RECT 16.090 14.605 16.420 14.625 ;
        RECT 16.075 14.345 16.435 14.605 ;
        RECT 16.090 14.325 16.420 14.345 ;
        RECT 16.650 14.065 16.820 14.765 ;
        RECT 17.050 14.605 17.380 14.625 ;
        RECT 17.035 14.345 17.395 14.605 ;
        RECT 17.050 14.325 17.380 14.345 ;
        RECT 11.410 13.895 16.820 14.065 ;
        RECT 19.015 14.065 19.185 14.810 ;
        RECT 20.385 14.765 20.615 15.285 ;
        RECT 21.345 14.765 21.575 15.285 ;
        RECT 22.305 14.765 22.535 15.285 ;
        RECT 23.265 14.765 23.495 15.285 ;
        RECT 24.225 14.765 24.455 15.285 ;
        RECT 19.855 14.610 20.185 14.625 ;
        RECT 19.840 14.350 20.200 14.610 ;
        RECT 19.855 14.325 20.185 14.350 ;
        RECT 20.415 14.065 20.585 14.765 ;
        RECT 20.815 14.610 21.145 14.625 ;
        RECT 20.795 14.350 21.155 14.610 ;
        RECT 20.815 14.325 21.145 14.350 ;
        RECT 21.375 14.065 21.545 14.765 ;
        RECT 21.775 14.610 22.105 14.625 ;
        RECT 21.755 14.350 22.115 14.610 ;
        RECT 21.775 14.325 22.105 14.350 ;
        RECT 22.335 14.065 22.505 14.765 ;
        RECT 22.735 14.610 23.065 14.625 ;
        RECT 22.715 14.350 23.075 14.610 ;
        RECT 22.735 14.325 23.065 14.350 ;
        RECT 23.295 14.065 23.465 14.765 ;
        RECT 23.695 14.605 24.025 14.625 ;
        RECT 23.680 14.345 24.040 14.605 ;
        RECT 23.695 14.325 24.025 14.345 ;
        RECT 24.255 14.065 24.425 14.765 ;
        RECT 24.655 14.605 24.985 14.625 ;
        RECT 24.640 14.345 25.000 14.605 ;
        RECT 24.655 14.325 24.985 14.345 ;
        RECT 19.015 13.895 24.425 14.065 ;
        RECT 11.410 12.500 16.820 12.670 ;
        RECT 1.535 10.370 1.765 11.730 ;
        RECT 2.495 10.370 2.725 11.730 ;
        RECT 3.455 10.370 3.685 11.730 ;
        RECT 4.415 10.370 4.645 11.730 ;
        RECT 5.375 10.370 5.605 11.730 ;
        RECT 6.335 10.370 6.565 11.730 ;
        RECT 1.565 9.665 1.735 10.370 ;
        RECT 2.525 9.665 2.695 10.370 ;
        RECT 3.485 9.665 3.655 10.370 ;
        RECT 4.445 9.665 4.615 10.370 ;
        RECT 5.405 9.665 5.575 10.370 ;
        RECT 6.365 9.665 6.535 10.370 ;
        RECT 11.410 9.685 11.580 12.500 ;
        RECT 12.810 11.750 12.980 12.500 ;
        RECT 13.770 11.750 13.940 12.500 ;
        RECT 14.730 11.750 14.900 12.500 ;
        RECT 15.690 11.750 15.860 12.500 ;
        RECT 16.650 11.750 16.820 12.500 ;
        RECT 19.015 12.500 24.425 12.670 ;
        RECT 12.300 10.390 12.530 11.750 ;
        RECT 12.780 10.390 13.010 11.750 ;
        RECT 13.260 10.390 13.490 11.750 ;
        RECT 13.740 10.390 13.970 11.750 ;
        RECT 14.220 10.390 14.450 11.750 ;
        RECT 14.700 10.390 14.930 11.750 ;
        RECT 15.180 10.390 15.410 11.750 ;
        RECT 15.660 10.390 15.890 11.750 ;
        RECT 16.140 10.390 16.370 11.750 ;
        RECT 16.620 10.390 16.850 11.750 ;
        RECT 17.100 10.390 17.330 11.750 ;
        RECT 10.505 9.665 11.580 9.685 ;
        RECT 1.565 9.515 11.580 9.665 ;
        RECT 1.565 9.495 10.705 9.515 ;
        RECT 1.565 8.830 1.735 9.495 ;
        RECT 2.525 8.830 2.695 9.495 ;
        RECT 3.485 8.830 3.655 9.495 ;
        RECT 4.445 8.830 4.615 9.495 ;
        RECT 5.405 8.830 5.575 9.495 ;
        RECT 6.365 8.830 6.535 9.495 ;
        RECT 1.535 8.310 1.765 8.830 ;
        RECT 2.495 8.310 2.725 8.830 ;
        RECT 3.455 8.310 3.685 8.830 ;
        RECT 4.415 8.310 4.645 8.830 ;
        RECT 5.375 8.310 5.605 8.830 ;
        RECT 6.335 8.310 6.565 8.830 ;
        RECT 11.410 7.630 11.580 9.515 ;
        RECT 12.330 9.685 12.500 10.390 ;
        RECT 13.290 9.685 13.460 10.390 ;
        RECT 14.250 9.685 14.420 10.390 ;
        RECT 15.210 9.685 15.380 10.390 ;
        RECT 16.170 9.685 16.340 10.390 ;
        RECT 17.130 9.685 17.300 10.390 ;
        RECT 19.015 9.685 19.185 12.500 ;
        RECT 20.415 11.750 20.585 12.500 ;
        RECT 21.375 11.750 21.545 12.500 ;
        RECT 22.335 11.750 22.505 12.500 ;
        RECT 23.295 11.750 23.465 12.500 ;
        RECT 24.255 11.750 24.425 12.500 ;
        RECT 20.385 10.390 20.615 11.750 ;
        RECT 21.345 10.390 21.575 11.750 ;
        RECT 22.305 10.390 22.535 11.750 ;
        RECT 23.265 10.390 23.495 11.750 ;
        RECT 24.225 10.390 24.455 11.750 ;
        RECT 12.330 9.515 19.185 9.685 ;
        RECT 12.330 8.850 12.500 9.515 ;
        RECT 13.290 8.850 13.460 9.515 ;
        RECT 14.250 8.850 14.420 9.515 ;
        RECT 15.210 8.850 15.380 9.515 ;
        RECT 16.170 8.850 16.340 9.515 ;
        RECT 17.130 8.850 17.300 9.515 ;
        RECT 19.015 8.875 19.185 9.515 ;
        RECT 26.630 9.220 27.000 9.490 ;
        RECT 18.670 8.870 19.185 8.875 ;
        RECT 12.300 8.330 12.530 8.850 ;
        RECT 12.780 8.330 13.010 8.850 ;
        RECT 13.260 8.330 13.490 8.850 ;
        RECT 13.740 8.330 13.970 8.850 ;
        RECT 14.220 8.330 14.450 8.850 ;
        RECT 14.700 8.330 14.930 8.850 ;
        RECT 15.180 8.330 15.410 8.850 ;
        RECT 15.660 8.330 15.890 8.850 ;
        RECT 16.140 8.330 16.370 8.850 ;
        RECT 16.620 8.330 16.850 8.850 ;
        RECT 17.100 8.330 17.330 8.850 ;
        RECT 18.645 8.375 19.185 8.870 ;
        RECT 18.645 8.370 18.875 8.375 ;
        RECT 12.250 8.175 12.580 8.190 ;
        RECT 12.235 7.915 12.595 8.175 ;
        RECT 12.250 7.890 12.580 7.915 ;
        RECT 12.810 7.630 12.980 8.330 ;
        RECT 13.210 8.175 13.540 8.190 ;
        RECT 13.190 7.915 13.550 8.175 ;
        RECT 13.210 7.890 13.540 7.915 ;
        RECT 13.770 7.630 13.940 8.330 ;
        RECT 14.170 8.175 14.500 8.190 ;
        RECT 14.150 7.915 14.510 8.175 ;
        RECT 14.170 7.890 14.500 7.915 ;
        RECT 14.730 7.630 14.900 8.330 ;
        RECT 15.130 8.175 15.460 8.190 ;
        RECT 15.110 7.915 15.470 8.175 ;
        RECT 15.130 7.890 15.460 7.915 ;
        RECT 15.690 7.630 15.860 8.330 ;
        RECT 16.090 8.170 16.420 8.190 ;
        RECT 16.075 7.910 16.435 8.170 ;
        RECT 16.090 7.890 16.420 7.910 ;
        RECT 16.650 7.630 16.820 8.330 ;
        RECT 17.050 8.170 17.380 8.190 ;
        RECT 17.035 7.910 17.395 8.170 ;
        RECT 17.050 7.890 17.380 7.910 ;
        RECT 11.410 7.460 16.820 7.630 ;
        RECT 19.015 7.630 19.185 8.375 ;
        RECT 20.385 8.330 20.615 8.850 ;
        RECT 21.345 8.330 21.575 8.850 ;
        RECT 22.305 8.330 22.535 8.850 ;
        RECT 23.265 8.330 23.495 8.850 ;
        RECT 24.225 8.330 24.455 8.850 ;
        RECT 19.855 8.175 20.185 8.190 ;
        RECT 19.840 7.915 20.200 8.175 ;
        RECT 19.855 7.890 20.185 7.915 ;
        RECT 20.415 7.630 20.585 8.330 ;
        RECT 20.815 8.175 21.145 8.190 ;
        RECT 20.795 7.915 21.155 8.175 ;
        RECT 20.815 7.890 21.145 7.915 ;
        RECT 21.375 7.630 21.545 8.330 ;
        RECT 21.775 8.175 22.105 8.190 ;
        RECT 21.755 7.915 22.115 8.175 ;
        RECT 21.775 7.890 22.105 7.915 ;
        RECT 22.335 7.630 22.505 8.330 ;
        RECT 22.735 8.175 23.065 8.190 ;
        RECT 22.715 7.915 23.075 8.175 ;
        RECT 22.735 7.890 23.065 7.915 ;
        RECT 23.295 7.630 23.465 8.330 ;
        RECT 23.695 8.170 24.025 8.190 ;
        RECT 23.680 7.910 24.040 8.170 ;
        RECT 23.695 7.890 24.025 7.910 ;
        RECT 24.255 7.630 24.425 8.330 ;
        RECT 24.655 8.170 24.985 8.190 ;
        RECT 24.640 7.910 25.000 8.170 ;
        RECT 24.655 7.890 24.985 7.910 ;
        RECT 19.015 7.460 24.425 7.630 ;
        RECT 11.410 6.065 16.820 6.235 ;
        RECT 1.535 3.935 1.765 5.295 ;
        RECT 2.495 3.935 2.725 5.295 ;
        RECT 3.455 3.935 3.685 5.295 ;
        RECT 4.415 3.935 4.645 5.295 ;
        RECT 5.375 3.935 5.605 5.295 ;
        RECT 6.335 3.935 6.565 5.295 ;
        RECT 1.565 3.230 1.735 3.935 ;
        RECT 2.525 3.230 2.695 3.935 ;
        RECT 3.485 3.230 3.655 3.935 ;
        RECT 4.445 3.230 4.615 3.935 ;
        RECT 5.405 3.230 5.575 3.935 ;
        RECT 6.365 3.230 6.535 3.935 ;
        RECT 11.410 3.250 11.580 6.065 ;
        RECT 12.810 5.315 12.980 6.065 ;
        RECT 13.770 5.315 13.940 6.065 ;
        RECT 14.730 5.315 14.900 6.065 ;
        RECT 15.690 5.315 15.860 6.065 ;
        RECT 16.650 5.315 16.820 6.065 ;
        RECT 19.015 6.065 24.425 6.235 ;
        RECT 12.300 3.955 12.530 5.315 ;
        RECT 12.780 3.955 13.010 5.315 ;
        RECT 13.260 3.955 13.490 5.315 ;
        RECT 13.740 3.955 13.970 5.315 ;
        RECT 14.220 3.955 14.450 5.315 ;
        RECT 14.700 3.955 14.930 5.315 ;
        RECT 15.180 3.955 15.410 5.315 ;
        RECT 15.660 3.955 15.890 5.315 ;
        RECT 16.140 3.955 16.370 5.315 ;
        RECT 16.620 3.955 16.850 5.315 ;
        RECT 17.100 3.955 17.330 5.315 ;
        RECT 10.505 3.230 11.580 3.250 ;
        RECT 1.565 3.080 11.580 3.230 ;
        RECT 1.565 3.060 10.705 3.080 ;
        RECT 1.565 2.395 1.735 3.060 ;
        RECT 2.525 2.395 2.695 3.060 ;
        RECT 3.485 2.395 3.655 3.060 ;
        RECT 4.445 2.395 4.615 3.060 ;
        RECT 5.405 2.395 5.575 3.060 ;
        RECT 6.365 2.395 6.535 3.060 ;
        RECT 1.535 1.875 1.765 2.395 ;
        RECT 2.495 1.875 2.725 2.395 ;
        RECT 3.455 1.875 3.685 2.395 ;
        RECT 4.415 1.875 4.645 2.395 ;
        RECT 5.375 1.875 5.605 2.395 ;
        RECT 6.335 1.875 6.565 2.395 ;
        RECT 11.410 1.195 11.580 3.080 ;
        RECT 12.330 3.250 12.500 3.955 ;
        RECT 13.290 3.250 13.460 3.955 ;
        RECT 14.250 3.250 14.420 3.955 ;
        RECT 15.210 3.250 15.380 3.955 ;
        RECT 16.170 3.250 16.340 3.955 ;
        RECT 17.130 3.250 17.300 3.955 ;
        RECT 19.015 3.250 19.185 6.065 ;
        RECT 20.415 5.315 20.585 6.065 ;
        RECT 21.375 5.315 21.545 6.065 ;
        RECT 22.335 5.315 22.505 6.065 ;
        RECT 23.295 5.315 23.465 6.065 ;
        RECT 24.255 5.315 24.425 6.065 ;
        RECT 20.385 3.955 20.615 5.315 ;
        RECT 21.345 3.955 21.575 5.315 ;
        RECT 22.305 3.955 22.535 5.315 ;
        RECT 23.265 3.955 23.495 5.315 ;
        RECT 24.225 3.955 24.455 5.315 ;
        RECT 12.330 3.080 19.185 3.250 ;
        RECT 12.330 2.415 12.500 3.080 ;
        RECT 13.290 2.415 13.460 3.080 ;
        RECT 14.250 2.415 14.420 3.080 ;
        RECT 15.210 2.415 15.380 3.080 ;
        RECT 16.170 2.415 16.340 3.080 ;
        RECT 17.130 2.415 17.300 3.080 ;
        RECT 19.015 2.440 19.185 3.080 ;
        RECT 26.630 2.785 27.000 3.055 ;
        RECT 18.670 2.435 19.185 2.440 ;
        RECT 12.300 1.895 12.530 2.415 ;
        RECT 12.780 1.895 13.010 2.415 ;
        RECT 13.260 1.895 13.490 2.415 ;
        RECT 13.740 1.895 13.970 2.415 ;
        RECT 14.220 1.895 14.450 2.415 ;
        RECT 14.700 1.895 14.930 2.415 ;
        RECT 15.180 1.895 15.410 2.415 ;
        RECT 15.660 1.895 15.890 2.415 ;
        RECT 16.140 1.895 16.370 2.415 ;
        RECT 16.620 1.895 16.850 2.415 ;
        RECT 17.100 1.895 17.330 2.415 ;
        RECT 18.645 1.940 19.185 2.435 ;
        RECT 18.645 1.935 18.875 1.940 ;
        RECT 12.250 1.740 12.580 1.755 ;
        RECT 12.235 1.480 12.595 1.740 ;
        RECT 12.250 1.455 12.580 1.480 ;
        RECT 12.810 1.195 12.980 1.895 ;
        RECT 13.210 1.740 13.540 1.755 ;
        RECT 13.190 1.480 13.550 1.740 ;
        RECT 13.210 1.455 13.540 1.480 ;
        RECT 13.770 1.195 13.940 1.895 ;
        RECT 14.170 1.740 14.500 1.755 ;
        RECT 14.150 1.480 14.510 1.740 ;
        RECT 14.170 1.455 14.500 1.480 ;
        RECT 14.730 1.195 14.900 1.895 ;
        RECT 15.130 1.740 15.460 1.755 ;
        RECT 15.110 1.480 15.470 1.740 ;
        RECT 15.130 1.455 15.460 1.480 ;
        RECT 15.690 1.195 15.860 1.895 ;
        RECT 16.090 1.735 16.420 1.755 ;
        RECT 16.075 1.475 16.435 1.735 ;
        RECT 16.090 1.455 16.420 1.475 ;
        RECT 16.650 1.195 16.820 1.895 ;
        RECT 17.050 1.735 17.380 1.755 ;
        RECT 17.035 1.475 17.395 1.735 ;
        RECT 17.050 1.455 17.380 1.475 ;
        RECT 11.410 1.025 16.820 1.195 ;
        RECT 19.015 1.195 19.185 1.940 ;
        RECT 20.385 1.895 20.615 2.415 ;
        RECT 21.345 1.895 21.575 2.415 ;
        RECT 22.305 1.895 22.535 2.415 ;
        RECT 23.265 1.895 23.495 2.415 ;
        RECT 24.225 1.895 24.455 2.415 ;
        RECT 19.855 1.740 20.185 1.755 ;
        RECT 19.840 1.480 20.200 1.740 ;
        RECT 19.855 1.455 20.185 1.480 ;
        RECT 20.415 1.195 20.585 1.895 ;
        RECT 20.815 1.740 21.145 1.755 ;
        RECT 20.795 1.480 21.155 1.740 ;
        RECT 20.815 1.455 21.145 1.480 ;
        RECT 21.375 1.195 21.545 1.895 ;
        RECT 21.775 1.740 22.105 1.755 ;
        RECT 21.755 1.480 22.115 1.740 ;
        RECT 21.775 1.455 22.105 1.480 ;
        RECT 22.335 1.195 22.505 1.895 ;
        RECT 22.735 1.740 23.065 1.755 ;
        RECT 22.715 1.480 23.075 1.740 ;
        RECT 22.735 1.455 23.065 1.480 ;
        RECT 23.295 1.195 23.465 1.895 ;
        RECT 23.695 1.735 24.025 1.755 ;
        RECT 23.680 1.475 24.040 1.735 ;
        RECT 23.695 1.455 24.025 1.475 ;
        RECT 24.255 1.195 24.425 1.895 ;
        RECT 24.655 1.735 24.985 1.755 ;
        RECT 24.640 1.475 25.000 1.735 ;
        RECT 24.655 1.455 24.985 1.475 ;
        RECT 19.015 1.025 24.425 1.195 ;
      LAYER via ;
        RECT 26.685 202.275 26.945 202.535 ;
        RECT 12.285 200.965 12.545 201.225 ;
        RECT 13.240 200.965 13.500 201.225 ;
        RECT 14.200 200.965 14.460 201.225 ;
        RECT 15.160 200.965 15.420 201.225 ;
        RECT 16.125 200.960 16.385 201.220 ;
        RECT 17.085 200.960 17.345 201.220 ;
        RECT 19.890 200.965 20.150 201.225 ;
        RECT 20.845 200.965 21.105 201.225 ;
        RECT 21.805 200.965 22.065 201.225 ;
        RECT 22.765 200.965 23.025 201.225 ;
        RECT 23.730 200.960 23.990 201.220 ;
        RECT 24.690 200.960 24.950 201.220 ;
        RECT 26.685 195.840 26.945 196.100 ;
        RECT 12.285 194.530 12.545 194.790 ;
        RECT 13.240 194.530 13.500 194.790 ;
        RECT 14.200 194.530 14.460 194.790 ;
        RECT 15.160 194.530 15.420 194.790 ;
        RECT 16.125 194.525 16.385 194.785 ;
        RECT 17.085 194.525 17.345 194.785 ;
        RECT 19.890 194.530 20.150 194.790 ;
        RECT 20.845 194.530 21.105 194.790 ;
        RECT 21.805 194.530 22.065 194.790 ;
        RECT 22.765 194.530 23.025 194.790 ;
        RECT 23.730 194.525 23.990 194.785 ;
        RECT 24.690 194.525 24.950 194.785 ;
        RECT 26.685 189.405 26.945 189.665 ;
        RECT 12.285 188.095 12.545 188.355 ;
        RECT 13.240 188.095 13.500 188.355 ;
        RECT 14.200 188.095 14.460 188.355 ;
        RECT 15.160 188.095 15.420 188.355 ;
        RECT 16.125 188.090 16.385 188.350 ;
        RECT 17.085 188.090 17.345 188.350 ;
        RECT 19.890 188.095 20.150 188.355 ;
        RECT 20.845 188.095 21.105 188.355 ;
        RECT 21.805 188.095 22.065 188.355 ;
        RECT 22.765 188.095 23.025 188.355 ;
        RECT 23.730 188.090 23.990 188.350 ;
        RECT 24.690 188.090 24.950 188.350 ;
        RECT 26.685 182.970 26.945 183.230 ;
        RECT 12.285 181.660 12.545 181.920 ;
        RECT 13.240 181.660 13.500 181.920 ;
        RECT 14.200 181.660 14.460 181.920 ;
        RECT 15.160 181.660 15.420 181.920 ;
        RECT 16.125 181.655 16.385 181.915 ;
        RECT 17.085 181.655 17.345 181.915 ;
        RECT 19.890 181.660 20.150 181.920 ;
        RECT 20.845 181.660 21.105 181.920 ;
        RECT 21.805 181.660 22.065 181.920 ;
        RECT 22.765 181.660 23.025 181.920 ;
        RECT 23.730 181.655 23.990 181.915 ;
        RECT 24.690 181.655 24.950 181.915 ;
        RECT 26.685 176.535 26.945 176.795 ;
        RECT 12.285 175.225 12.545 175.485 ;
        RECT 13.240 175.225 13.500 175.485 ;
        RECT 14.200 175.225 14.460 175.485 ;
        RECT 15.160 175.225 15.420 175.485 ;
        RECT 16.125 175.220 16.385 175.480 ;
        RECT 17.085 175.220 17.345 175.480 ;
        RECT 19.890 175.225 20.150 175.485 ;
        RECT 20.845 175.225 21.105 175.485 ;
        RECT 21.805 175.225 22.065 175.485 ;
        RECT 22.765 175.225 23.025 175.485 ;
        RECT 23.730 175.220 23.990 175.480 ;
        RECT 24.690 175.220 24.950 175.480 ;
        RECT 26.685 170.100 26.945 170.360 ;
        RECT 12.285 168.790 12.545 169.050 ;
        RECT 13.240 168.790 13.500 169.050 ;
        RECT 14.200 168.790 14.460 169.050 ;
        RECT 15.160 168.790 15.420 169.050 ;
        RECT 16.125 168.785 16.385 169.045 ;
        RECT 17.085 168.785 17.345 169.045 ;
        RECT 19.890 168.790 20.150 169.050 ;
        RECT 20.845 168.790 21.105 169.050 ;
        RECT 21.805 168.790 22.065 169.050 ;
        RECT 22.765 168.790 23.025 169.050 ;
        RECT 23.730 168.785 23.990 169.045 ;
        RECT 24.690 168.785 24.950 169.045 ;
        RECT 26.685 163.665 26.945 163.925 ;
        RECT 12.285 162.355 12.545 162.615 ;
        RECT 13.240 162.355 13.500 162.615 ;
        RECT 14.200 162.355 14.460 162.615 ;
        RECT 15.160 162.355 15.420 162.615 ;
        RECT 16.125 162.350 16.385 162.610 ;
        RECT 17.085 162.350 17.345 162.610 ;
        RECT 19.890 162.355 20.150 162.615 ;
        RECT 20.845 162.355 21.105 162.615 ;
        RECT 21.805 162.355 22.065 162.615 ;
        RECT 22.765 162.355 23.025 162.615 ;
        RECT 23.730 162.350 23.990 162.610 ;
        RECT 24.690 162.350 24.950 162.610 ;
        RECT 26.685 157.230 26.945 157.490 ;
        RECT 12.285 155.920 12.545 156.180 ;
        RECT 13.240 155.920 13.500 156.180 ;
        RECT 14.200 155.920 14.460 156.180 ;
        RECT 15.160 155.920 15.420 156.180 ;
        RECT 16.125 155.915 16.385 156.175 ;
        RECT 17.085 155.915 17.345 156.175 ;
        RECT 19.890 155.920 20.150 156.180 ;
        RECT 20.845 155.920 21.105 156.180 ;
        RECT 21.805 155.920 22.065 156.180 ;
        RECT 22.765 155.920 23.025 156.180 ;
        RECT 23.730 155.915 23.990 156.175 ;
        RECT 24.690 155.915 24.950 156.175 ;
        RECT 26.685 150.795 26.945 151.055 ;
        RECT 12.285 149.485 12.545 149.745 ;
        RECT 13.240 149.485 13.500 149.745 ;
        RECT 14.200 149.485 14.460 149.745 ;
        RECT 15.160 149.485 15.420 149.745 ;
        RECT 16.125 149.480 16.385 149.740 ;
        RECT 17.085 149.480 17.345 149.740 ;
        RECT 19.890 149.485 20.150 149.745 ;
        RECT 20.845 149.485 21.105 149.745 ;
        RECT 21.805 149.485 22.065 149.745 ;
        RECT 22.765 149.485 23.025 149.745 ;
        RECT 23.730 149.480 23.990 149.740 ;
        RECT 24.690 149.480 24.950 149.740 ;
        RECT 26.685 144.360 26.945 144.620 ;
        RECT 12.285 143.050 12.545 143.310 ;
        RECT 13.240 143.050 13.500 143.310 ;
        RECT 14.200 143.050 14.460 143.310 ;
        RECT 15.160 143.050 15.420 143.310 ;
        RECT 16.125 143.045 16.385 143.305 ;
        RECT 17.085 143.045 17.345 143.305 ;
        RECT 19.890 143.050 20.150 143.310 ;
        RECT 20.845 143.050 21.105 143.310 ;
        RECT 21.805 143.050 22.065 143.310 ;
        RECT 22.765 143.050 23.025 143.310 ;
        RECT 23.730 143.045 23.990 143.305 ;
        RECT 24.690 143.045 24.950 143.305 ;
        RECT 26.685 137.925 26.945 138.185 ;
        RECT 12.285 136.615 12.545 136.875 ;
        RECT 13.240 136.615 13.500 136.875 ;
        RECT 14.200 136.615 14.460 136.875 ;
        RECT 15.160 136.615 15.420 136.875 ;
        RECT 16.125 136.610 16.385 136.870 ;
        RECT 17.085 136.610 17.345 136.870 ;
        RECT 19.890 136.615 20.150 136.875 ;
        RECT 20.845 136.615 21.105 136.875 ;
        RECT 21.805 136.615 22.065 136.875 ;
        RECT 22.765 136.615 23.025 136.875 ;
        RECT 23.730 136.610 23.990 136.870 ;
        RECT 24.690 136.610 24.950 136.870 ;
        RECT 26.685 131.490 26.945 131.750 ;
        RECT 12.285 130.180 12.545 130.440 ;
        RECT 13.240 130.180 13.500 130.440 ;
        RECT 14.200 130.180 14.460 130.440 ;
        RECT 15.160 130.180 15.420 130.440 ;
        RECT 16.125 130.175 16.385 130.435 ;
        RECT 17.085 130.175 17.345 130.435 ;
        RECT 19.890 130.180 20.150 130.440 ;
        RECT 20.845 130.180 21.105 130.440 ;
        RECT 21.805 130.180 22.065 130.440 ;
        RECT 22.765 130.180 23.025 130.440 ;
        RECT 23.730 130.175 23.990 130.435 ;
        RECT 24.690 130.175 24.950 130.435 ;
        RECT 26.685 125.055 26.945 125.315 ;
        RECT 12.285 123.745 12.545 124.005 ;
        RECT 13.240 123.745 13.500 124.005 ;
        RECT 14.200 123.745 14.460 124.005 ;
        RECT 15.160 123.745 15.420 124.005 ;
        RECT 16.125 123.740 16.385 124.000 ;
        RECT 17.085 123.740 17.345 124.000 ;
        RECT 19.890 123.745 20.150 124.005 ;
        RECT 20.845 123.745 21.105 124.005 ;
        RECT 21.805 123.745 22.065 124.005 ;
        RECT 22.765 123.745 23.025 124.005 ;
        RECT 23.730 123.740 23.990 124.000 ;
        RECT 24.690 123.740 24.950 124.000 ;
        RECT 26.685 118.620 26.945 118.880 ;
        RECT 12.285 117.310 12.545 117.570 ;
        RECT 13.240 117.310 13.500 117.570 ;
        RECT 14.200 117.310 14.460 117.570 ;
        RECT 15.160 117.310 15.420 117.570 ;
        RECT 16.125 117.305 16.385 117.565 ;
        RECT 17.085 117.305 17.345 117.565 ;
        RECT 19.890 117.310 20.150 117.570 ;
        RECT 20.845 117.310 21.105 117.570 ;
        RECT 21.805 117.310 22.065 117.570 ;
        RECT 22.765 117.310 23.025 117.570 ;
        RECT 23.730 117.305 23.990 117.565 ;
        RECT 24.690 117.305 24.950 117.565 ;
        RECT 26.685 112.185 26.945 112.445 ;
        RECT 12.285 110.875 12.545 111.135 ;
        RECT 13.240 110.875 13.500 111.135 ;
        RECT 14.200 110.875 14.460 111.135 ;
        RECT 15.160 110.875 15.420 111.135 ;
        RECT 16.125 110.870 16.385 111.130 ;
        RECT 17.085 110.870 17.345 111.130 ;
        RECT 19.890 110.875 20.150 111.135 ;
        RECT 20.845 110.875 21.105 111.135 ;
        RECT 21.805 110.875 22.065 111.135 ;
        RECT 22.765 110.875 23.025 111.135 ;
        RECT 23.730 110.870 23.990 111.130 ;
        RECT 24.690 110.870 24.950 111.130 ;
        RECT 26.685 105.750 26.945 106.010 ;
        RECT 12.285 104.440 12.545 104.700 ;
        RECT 13.240 104.440 13.500 104.700 ;
        RECT 14.200 104.440 14.460 104.700 ;
        RECT 15.160 104.440 15.420 104.700 ;
        RECT 16.125 104.435 16.385 104.695 ;
        RECT 17.085 104.435 17.345 104.695 ;
        RECT 19.890 104.440 20.150 104.700 ;
        RECT 20.845 104.440 21.105 104.700 ;
        RECT 21.805 104.440 22.065 104.700 ;
        RECT 22.765 104.440 23.025 104.700 ;
        RECT 23.730 104.435 23.990 104.695 ;
        RECT 24.690 104.435 24.950 104.695 ;
        RECT 26.685 99.315 26.945 99.575 ;
        RECT 12.285 98.005 12.545 98.265 ;
        RECT 13.240 98.005 13.500 98.265 ;
        RECT 14.200 98.005 14.460 98.265 ;
        RECT 15.160 98.005 15.420 98.265 ;
        RECT 16.125 98.000 16.385 98.260 ;
        RECT 17.085 98.000 17.345 98.260 ;
        RECT 19.890 98.005 20.150 98.265 ;
        RECT 20.845 98.005 21.105 98.265 ;
        RECT 21.805 98.005 22.065 98.265 ;
        RECT 22.765 98.005 23.025 98.265 ;
        RECT 23.730 98.000 23.990 98.260 ;
        RECT 24.690 98.000 24.950 98.260 ;
        RECT 26.685 92.880 26.945 93.140 ;
        RECT 12.285 91.570 12.545 91.830 ;
        RECT 13.240 91.570 13.500 91.830 ;
        RECT 14.200 91.570 14.460 91.830 ;
        RECT 15.160 91.570 15.420 91.830 ;
        RECT 16.125 91.565 16.385 91.825 ;
        RECT 17.085 91.565 17.345 91.825 ;
        RECT 19.890 91.570 20.150 91.830 ;
        RECT 20.845 91.570 21.105 91.830 ;
        RECT 21.805 91.570 22.065 91.830 ;
        RECT 22.765 91.570 23.025 91.830 ;
        RECT 23.730 91.565 23.990 91.825 ;
        RECT 24.690 91.565 24.950 91.825 ;
        RECT 26.685 86.445 26.945 86.705 ;
        RECT 12.285 85.135 12.545 85.395 ;
        RECT 13.240 85.135 13.500 85.395 ;
        RECT 14.200 85.135 14.460 85.395 ;
        RECT 15.160 85.135 15.420 85.395 ;
        RECT 16.125 85.130 16.385 85.390 ;
        RECT 17.085 85.130 17.345 85.390 ;
        RECT 19.890 85.135 20.150 85.395 ;
        RECT 20.845 85.135 21.105 85.395 ;
        RECT 21.805 85.135 22.065 85.395 ;
        RECT 22.765 85.135 23.025 85.395 ;
        RECT 23.730 85.130 23.990 85.390 ;
        RECT 24.690 85.130 24.950 85.390 ;
        RECT 26.685 80.010 26.945 80.270 ;
        RECT 12.285 78.700 12.545 78.960 ;
        RECT 13.240 78.700 13.500 78.960 ;
        RECT 14.200 78.700 14.460 78.960 ;
        RECT 15.160 78.700 15.420 78.960 ;
        RECT 16.125 78.695 16.385 78.955 ;
        RECT 17.085 78.695 17.345 78.955 ;
        RECT 19.890 78.700 20.150 78.960 ;
        RECT 20.845 78.700 21.105 78.960 ;
        RECT 21.805 78.700 22.065 78.960 ;
        RECT 22.765 78.700 23.025 78.960 ;
        RECT 23.730 78.695 23.990 78.955 ;
        RECT 24.690 78.695 24.950 78.955 ;
        RECT 26.685 73.575 26.945 73.835 ;
        RECT 12.285 72.265 12.545 72.525 ;
        RECT 13.240 72.265 13.500 72.525 ;
        RECT 14.200 72.265 14.460 72.525 ;
        RECT 15.160 72.265 15.420 72.525 ;
        RECT 16.125 72.260 16.385 72.520 ;
        RECT 17.085 72.260 17.345 72.520 ;
        RECT 19.890 72.265 20.150 72.525 ;
        RECT 20.845 72.265 21.105 72.525 ;
        RECT 21.805 72.265 22.065 72.525 ;
        RECT 22.765 72.265 23.025 72.525 ;
        RECT 23.730 72.260 23.990 72.520 ;
        RECT 24.690 72.260 24.950 72.520 ;
        RECT 26.685 67.140 26.945 67.400 ;
        RECT 12.285 65.830 12.545 66.090 ;
        RECT 13.240 65.830 13.500 66.090 ;
        RECT 14.200 65.830 14.460 66.090 ;
        RECT 15.160 65.830 15.420 66.090 ;
        RECT 16.125 65.825 16.385 66.085 ;
        RECT 17.085 65.825 17.345 66.085 ;
        RECT 19.890 65.830 20.150 66.090 ;
        RECT 20.845 65.830 21.105 66.090 ;
        RECT 21.805 65.830 22.065 66.090 ;
        RECT 22.765 65.830 23.025 66.090 ;
        RECT 23.730 65.825 23.990 66.085 ;
        RECT 24.690 65.825 24.950 66.085 ;
        RECT 26.685 60.705 26.945 60.965 ;
        RECT 12.285 59.395 12.545 59.655 ;
        RECT 13.240 59.395 13.500 59.655 ;
        RECT 14.200 59.395 14.460 59.655 ;
        RECT 15.160 59.395 15.420 59.655 ;
        RECT 16.125 59.390 16.385 59.650 ;
        RECT 17.085 59.390 17.345 59.650 ;
        RECT 19.890 59.395 20.150 59.655 ;
        RECT 20.845 59.395 21.105 59.655 ;
        RECT 21.805 59.395 22.065 59.655 ;
        RECT 22.765 59.395 23.025 59.655 ;
        RECT 23.730 59.390 23.990 59.650 ;
        RECT 24.690 59.390 24.950 59.650 ;
        RECT 26.685 54.270 26.945 54.530 ;
        RECT 12.285 52.960 12.545 53.220 ;
        RECT 13.240 52.960 13.500 53.220 ;
        RECT 14.200 52.960 14.460 53.220 ;
        RECT 15.160 52.960 15.420 53.220 ;
        RECT 16.125 52.955 16.385 53.215 ;
        RECT 17.085 52.955 17.345 53.215 ;
        RECT 19.890 52.960 20.150 53.220 ;
        RECT 20.845 52.960 21.105 53.220 ;
        RECT 21.805 52.960 22.065 53.220 ;
        RECT 22.765 52.960 23.025 53.220 ;
        RECT 23.730 52.955 23.990 53.215 ;
        RECT 24.690 52.955 24.950 53.215 ;
        RECT 26.685 47.835 26.945 48.095 ;
        RECT 12.285 46.525 12.545 46.785 ;
        RECT 13.240 46.525 13.500 46.785 ;
        RECT 14.200 46.525 14.460 46.785 ;
        RECT 15.160 46.525 15.420 46.785 ;
        RECT 16.125 46.520 16.385 46.780 ;
        RECT 17.085 46.520 17.345 46.780 ;
        RECT 19.890 46.525 20.150 46.785 ;
        RECT 20.845 46.525 21.105 46.785 ;
        RECT 21.805 46.525 22.065 46.785 ;
        RECT 22.765 46.525 23.025 46.785 ;
        RECT 23.730 46.520 23.990 46.780 ;
        RECT 24.690 46.520 24.950 46.780 ;
        RECT 26.685 41.400 26.945 41.660 ;
        RECT 12.285 40.090 12.545 40.350 ;
        RECT 13.240 40.090 13.500 40.350 ;
        RECT 14.200 40.090 14.460 40.350 ;
        RECT 15.160 40.090 15.420 40.350 ;
        RECT 16.125 40.085 16.385 40.345 ;
        RECT 17.085 40.085 17.345 40.345 ;
        RECT 19.890 40.090 20.150 40.350 ;
        RECT 20.845 40.090 21.105 40.350 ;
        RECT 21.805 40.090 22.065 40.350 ;
        RECT 22.765 40.090 23.025 40.350 ;
        RECT 23.730 40.085 23.990 40.345 ;
        RECT 24.690 40.085 24.950 40.345 ;
        RECT 26.685 34.965 26.945 35.225 ;
        RECT 12.285 33.655 12.545 33.915 ;
        RECT 13.240 33.655 13.500 33.915 ;
        RECT 14.200 33.655 14.460 33.915 ;
        RECT 15.160 33.655 15.420 33.915 ;
        RECT 16.125 33.650 16.385 33.910 ;
        RECT 17.085 33.650 17.345 33.910 ;
        RECT 19.890 33.655 20.150 33.915 ;
        RECT 20.845 33.655 21.105 33.915 ;
        RECT 21.805 33.655 22.065 33.915 ;
        RECT 22.765 33.655 23.025 33.915 ;
        RECT 23.730 33.650 23.990 33.910 ;
        RECT 24.690 33.650 24.950 33.910 ;
        RECT 26.685 28.530 26.945 28.790 ;
        RECT 12.285 27.220 12.545 27.480 ;
        RECT 13.240 27.220 13.500 27.480 ;
        RECT 14.200 27.220 14.460 27.480 ;
        RECT 15.160 27.220 15.420 27.480 ;
        RECT 16.125 27.215 16.385 27.475 ;
        RECT 17.085 27.215 17.345 27.475 ;
        RECT 19.890 27.220 20.150 27.480 ;
        RECT 20.845 27.220 21.105 27.480 ;
        RECT 21.805 27.220 22.065 27.480 ;
        RECT 22.765 27.220 23.025 27.480 ;
        RECT 23.730 27.215 23.990 27.475 ;
        RECT 24.690 27.215 24.950 27.475 ;
        RECT 26.685 22.095 26.945 22.355 ;
        RECT 12.285 20.785 12.545 21.045 ;
        RECT 13.240 20.785 13.500 21.045 ;
        RECT 14.200 20.785 14.460 21.045 ;
        RECT 15.160 20.785 15.420 21.045 ;
        RECT 16.125 20.780 16.385 21.040 ;
        RECT 17.085 20.780 17.345 21.040 ;
        RECT 19.890 20.785 20.150 21.045 ;
        RECT 20.845 20.785 21.105 21.045 ;
        RECT 21.805 20.785 22.065 21.045 ;
        RECT 22.765 20.785 23.025 21.045 ;
        RECT 23.730 20.780 23.990 21.040 ;
        RECT 24.690 20.780 24.950 21.040 ;
        RECT 26.685 15.660 26.945 15.920 ;
        RECT 12.285 14.350 12.545 14.610 ;
        RECT 13.240 14.350 13.500 14.610 ;
        RECT 14.200 14.350 14.460 14.610 ;
        RECT 15.160 14.350 15.420 14.610 ;
        RECT 16.125 14.345 16.385 14.605 ;
        RECT 17.085 14.345 17.345 14.605 ;
        RECT 19.890 14.350 20.150 14.610 ;
        RECT 20.845 14.350 21.105 14.610 ;
        RECT 21.805 14.350 22.065 14.610 ;
        RECT 22.765 14.350 23.025 14.610 ;
        RECT 23.730 14.345 23.990 14.605 ;
        RECT 24.690 14.345 24.950 14.605 ;
        RECT 26.685 9.225 26.945 9.485 ;
        RECT 12.285 7.915 12.545 8.175 ;
        RECT 13.240 7.915 13.500 8.175 ;
        RECT 14.200 7.915 14.460 8.175 ;
        RECT 15.160 7.915 15.420 8.175 ;
        RECT 16.125 7.910 16.385 8.170 ;
        RECT 17.085 7.910 17.345 8.170 ;
        RECT 19.890 7.915 20.150 8.175 ;
        RECT 20.845 7.915 21.105 8.175 ;
        RECT 21.805 7.915 22.065 8.175 ;
        RECT 22.765 7.915 23.025 8.175 ;
        RECT 23.730 7.910 23.990 8.170 ;
        RECT 24.690 7.910 24.950 8.170 ;
        RECT 26.685 2.790 26.945 3.050 ;
        RECT 12.285 1.480 12.545 1.740 ;
        RECT 13.240 1.480 13.500 1.740 ;
        RECT 14.200 1.480 14.460 1.740 ;
        RECT 15.160 1.480 15.420 1.740 ;
        RECT 16.125 1.475 16.385 1.735 ;
        RECT 17.085 1.475 17.345 1.735 ;
        RECT 19.890 1.480 20.150 1.740 ;
        RECT 20.845 1.480 21.105 1.740 ;
        RECT 21.805 1.480 22.065 1.740 ;
        RECT 22.765 1.480 23.025 1.740 ;
        RECT 23.730 1.475 23.990 1.735 ;
        RECT 24.690 1.475 24.950 1.735 ;
      LAYER met2 ;
        RECT 18 146 26 149 ;
        RECT 26.680 202.500 26.950 202.590 ;
        RECT 25.890 202.240 26.950 202.500 ;
        RECT 12.285 201.225 12.545 201.275 ;
        RECT 13.240 201.225 13.500 201.275 ;
        RECT 14.200 201.225 14.460 201.275 ;
        RECT 15.160 201.225 15.420 201.275 ;
        RECT 16.125 201.225 16.385 201.270 ;
        RECT 17.085 201.225 17.345 201.270 ;
        RECT 19.890 201.225 20.150 201.275 ;
        RECT 20.845 201.225 21.105 201.275 ;
        RECT 21.805 201.225 22.065 201.275 ;
        RECT 22.765 201.225 23.025 201.275 ;
        RECT 23.730 201.225 23.990 201.270 ;
        RECT 24.690 201.225 24.950 201.270 ;
        RECT 25.890 201.225 26.150 202.240 ;
        RECT 26.680 202.220 26.950 202.240 ;
        RECT 11.145 200.965 26.150 201.225 ;
        RECT 12.285 200.915 12.545 200.965 ;
        RECT 13.240 200.915 13.500 200.965 ;
        RECT 14.200 200.915 14.460 200.965 ;
        RECT 15.160 200.915 15.420 200.965 ;
        RECT 16.125 200.910 16.385 200.965 ;
        RECT 17.085 200.910 17.345 200.965 ;
        RECT 19.890 200.915 20.150 200.965 ;
        RECT 20.845 200.915 21.105 200.965 ;
        RECT 21.805 200.915 22.065 200.965 ;
        RECT 22.765 200.915 23.025 200.965 ;
        RECT 23.730 200.910 23.990 200.965 ;
        RECT 24.690 200.910 24.950 200.965 ;
        RECT 26.680 196.065 26.950 196.155 ;
        RECT 25.890 195.805 26.950 196.065 ;
        RECT 12.285 194.790 12.545 194.840 ;
        RECT 13.240 194.790 13.500 194.840 ;
        RECT 14.200 194.790 14.460 194.840 ;
        RECT 15.160 194.790 15.420 194.840 ;
        RECT 16.125 194.790 16.385 194.835 ;
        RECT 17.085 194.790 17.345 194.835 ;
        RECT 19.890 194.790 20.150 194.840 ;
        RECT 20.845 194.790 21.105 194.840 ;
        RECT 21.805 194.790 22.065 194.840 ;
        RECT 22.765 194.790 23.025 194.840 ;
        RECT 23.730 194.790 23.990 194.835 ;
        RECT 24.690 194.790 24.950 194.835 ;
        RECT 25.890 194.790 26.150 195.805 ;
        RECT 26.680 195.785 26.950 195.805 ;
        RECT 11.145 194.530 26.150 194.790 ;
        RECT 12.285 194.480 12.545 194.530 ;
        RECT 13.240 194.480 13.500 194.530 ;
        RECT 14.200 194.480 14.460 194.530 ;
        RECT 15.160 194.480 15.420 194.530 ;
        RECT 16.125 194.475 16.385 194.530 ;
        RECT 17.085 194.475 17.345 194.530 ;
        RECT 19.890 194.480 20.150 194.530 ;
        RECT 20.845 194.480 21.105 194.530 ;
        RECT 21.805 194.480 22.065 194.530 ;
        RECT 22.765 194.480 23.025 194.530 ;
        RECT 23.730 194.475 23.990 194.530 ;
        RECT 24.690 194.475 24.950 194.530 ;
        RECT 26.680 189.630 26.950 189.720 ;
        RECT 25.890 189.370 26.950 189.630 ;
        RECT 12.285 188.355 12.545 188.405 ;
        RECT 13.240 188.355 13.500 188.405 ;
        RECT 14.200 188.355 14.460 188.405 ;
        RECT 15.160 188.355 15.420 188.405 ;
        RECT 16.125 188.355 16.385 188.400 ;
        RECT 17.085 188.355 17.345 188.400 ;
        RECT 19.890 188.355 20.150 188.405 ;
        RECT 20.845 188.355 21.105 188.405 ;
        RECT 21.805 188.355 22.065 188.405 ;
        RECT 22.765 188.355 23.025 188.405 ;
        RECT 23.730 188.355 23.990 188.400 ;
        RECT 24.690 188.355 24.950 188.400 ;
        RECT 25.890 188.355 26.150 189.370 ;
        RECT 26.680 189.350 26.950 189.370 ;
        RECT 11.145 188.095 26.150 188.355 ;
        RECT 12.285 188.045 12.545 188.095 ;
        RECT 13.240 188.045 13.500 188.095 ;
        RECT 14.200 188.045 14.460 188.095 ;
        RECT 15.160 188.045 15.420 188.095 ;
        RECT 16.125 188.040 16.385 188.095 ;
        RECT 17.085 188.040 17.345 188.095 ;
        RECT 19.890 188.045 20.150 188.095 ;
        RECT 20.845 188.045 21.105 188.095 ;
        RECT 21.805 188.045 22.065 188.095 ;
        RECT 22.765 188.045 23.025 188.095 ;
        RECT 23.730 188.040 23.990 188.095 ;
        RECT 24.690 188.040 24.950 188.095 ;
        RECT 26.680 183.195 26.950 183.285 ;
        RECT 25.890 182.935 26.950 183.195 ;
        RECT 12.285 181.920 12.545 181.970 ;
        RECT 13.240 181.920 13.500 181.970 ;
        RECT 14.200 181.920 14.460 181.970 ;
        RECT 15.160 181.920 15.420 181.970 ;
        RECT 16.125 181.920 16.385 181.965 ;
        RECT 17.085 181.920 17.345 181.965 ;
        RECT 19.890 181.920 20.150 181.970 ;
        RECT 20.845 181.920 21.105 181.970 ;
        RECT 21.805 181.920 22.065 181.970 ;
        RECT 22.765 181.920 23.025 181.970 ;
        RECT 23.730 181.920 23.990 181.965 ;
        RECT 24.690 181.920 24.950 181.965 ;
        RECT 25.890 181.920 26.150 182.935 ;
        RECT 26.680 182.915 26.950 182.935 ;
        RECT 11.145 181.660 26.150 181.920 ;
        RECT 12.285 181.610 12.545 181.660 ;
        RECT 13.240 181.610 13.500 181.660 ;
        RECT 14.200 181.610 14.460 181.660 ;
        RECT 15.160 181.610 15.420 181.660 ;
        RECT 16.125 181.605 16.385 181.660 ;
        RECT 17.085 181.605 17.345 181.660 ;
        RECT 19.890 181.610 20.150 181.660 ;
        RECT 20.845 181.610 21.105 181.660 ;
        RECT 21.805 181.610 22.065 181.660 ;
        RECT 22.765 181.610 23.025 181.660 ;
        RECT 23.730 181.605 23.990 181.660 ;
        RECT 24.690 181.605 24.950 181.660 ;
        RECT 26.680 176.760 26.950 176.850 ;
        RECT 25.890 176.500 26.950 176.760 ;
        RECT 12.285 175.485 12.545 175.535 ;
        RECT 13.240 175.485 13.500 175.535 ;
        RECT 14.200 175.485 14.460 175.535 ;
        RECT 15.160 175.485 15.420 175.535 ;
        RECT 16.125 175.485 16.385 175.530 ;
        RECT 17.085 175.485 17.345 175.530 ;
        RECT 19.890 175.485 20.150 175.535 ;
        RECT 20.845 175.485 21.105 175.535 ;
        RECT 21.805 175.485 22.065 175.535 ;
        RECT 22.765 175.485 23.025 175.535 ;
        RECT 23.730 175.485 23.990 175.530 ;
        RECT 24.690 175.485 24.950 175.530 ;
        RECT 25.890 175.485 26.150 176.500 ;
        RECT 26.680 176.480 26.950 176.500 ;
        RECT 11.145 175.225 26.150 175.485 ;
        RECT 12.285 175.175 12.545 175.225 ;
        RECT 13.240 175.175 13.500 175.225 ;
        RECT 14.200 175.175 14.460 175.225 ;
        RECT 15.160 175.175 15.420 175.225 ;
        RECT 16.125 175.170 16.385 175.225 ;
        RECT 17.085 175.170 17.345 175.225 ;
        RECT 19.890 175.175 20.150 175.225 ;
        RECT 20.845 175.175 21.105 175.225 ;
        RECT 21.805 175.175 22.065 175.225 ;
        RECT 22.765 175.175 23.025 175.225 ;
        RECT 23.730 175.170 23.990 175.225 ;
        RECT 24.690 175.170 24.950 175.225 ;
        RECT 26.680 170.325 26.950 170.415 ;
        RECT 25.890 170.065 26.950 170.325 ;
        RECT 12.285 169.050 12.545 169.100 ;
        RECT 13.240 169.050 13.500 169.100 ;
        RECT 14.200 169.050 14.460 169.100 ;
        RECT 15.160 169.050 15.420 169.100 ;
        RECT 16.125 169.050 16.385 169.095 ;
        RECT 17.085 169.050 17.345 169.095 ;
        RECT 19.890 169.050 20.150 169.100 ;
        RECT 20.845 169.050 21.105 169.100 ;
        RECT 21.805 169.050 22.065 169.100 ;
        RECT 22.765 169.050 23.025 169.100 ;
        RECT 23.730 169.050 23.990 169.095 ;
        RECT 24.690 169.050 24.950 169.095 ;
        RECT 25.890 169.050 26.150 170.065 ;
        RECT 26.680 170.045 26.950 170.065 ;
        RECT 11.145 168.790 26.150 169.050 ;
        RECT 12.285 168.740 12.545 168.790 ;
        RECT 13.240 168.740 13.500 168.790 ;
        RECT 14.200 168.740 14.460 168.790 ;
        RECT 15.160 168.740 15.420 168.790 ;
        RECT 16.125 168.735 16.385 168.790 ;
        RECT 17.085 168.735 17.345 168.790 ;
        RECT 19.890 168.740 20.150 168.790 ;
        RECT 20.845 168.740 21.105 168.790 ;
        RECT 21.805 168.740 22.065 168.790 ;
        RECT 22.765 168.740 23.025 168.790 ;
        RECT 23.730 168.735 23.990 168.790 ;
        RECT 24.690 168.735 24.950 168.790 ;
        RECT 26.680 163.890 26.950 163.980 ;
        RECT 25.890 163.630 26.950 163.890 ;
        RECT 12.285 162.615 12.545 162.665 ;
        RECT 13.240 162.615 13.500 162.665 ;
        RECT 14.200 162.615 14.460 162.665 ;
        RECT 15.160 162.615 15.420 162.665 ;
        RECT 16.125 162.615 16.385 162.660 ;
        RECT 17.085 162.615 17.345 162.660 ;
        RECT 19.890 162.615 20.150 162.665 ;
        RECT 20.845 162.615 21.105 162.665 ;
        RECT 21.805 162.615 22.065 162.665 ;
        RECT 22.765 162.615 23.025 162.665 ;
        RECT 23.730 162.615 23.990 162.660 ;
        RECT 24.690 162.615 24.950 162.660 ;
        RECT 25.890 162.615 26.150 163.630 ;
        RECT 26.680 163.610 26.950 163.630 ;
        RECT 11.145 162.355 26.150 162.615 ;
        RECT 12.285 162.305 12.545 162.355 ;
        RECT 13.240 162.305 13.500 162.355 ;
        RECT 14.200 162.305 14.460 162.355 ;
        RECT 15.160 162.305 15.420 162.355 ;
        RECT 16.125 162.300 16.385 162.355 ;
        RECT 17.085 162.300 17.345 162.355 ;
        RECT 19.890 162.305 20.150 162.355 ;
        RECT 20.845 162.305 21.105 162.355 ;
        RECT 21.805 162.305 22.065 162.355 ;
        RECT 22.765 162.305 23.025 162.355 ;
        RECT 23.730 162.300 23.990 162.355 ;
        RECT 24.690 162.300 24.950 162.355 ;
        RECT 26.680 157.455 26.950 157.545 ;
        RECT 25.890 157.195 26.950 157.455 ;
        RECT 12.285 156.180 12.545 156.230 ;
        RECT 13.240 156.180 13.500 156.230 ;
        RECT 14.200 156.180 14.460 156.230 ;
        RECT 15.160 156.180 15.420 156.230 ;
        RECT 16.125 156.180 16.385 156.225 ;
        RECT 17.085 156.180 17.345 156.225 ;
        RECT 19.890 156.180 20.150 156.230 ;
        RECT 20.845 156.180 21.105 156.230 ;
        RECT 21.805 156.180 22.065 156.230 ;
        RECT 22.765 156.180 23.025 156.230 ;
        RECT 23.730 156.180 23.990 156.225 ;
        RECT 24.690 156.180 24.950 156.225 ;
        RECT 25.890 156.180 26.150 157.195 ;
        RECT 26.680 157.175 26.950 157.195 ;
        RECT 11.145 155.920 26.150 156.180 ;
        RECT 12.285 155.870 12.545 155.920 ;
        RECT 13.240 155.870 13.500 155.920 ;
        RECT 14.200 155.870 14.460 155.920 ;
        RECT 15.160 155.870 15.420 155.920 ;
        RECT 16.125 155.865 16.385 155.920 ;
        RECT 17.085 155.865 17.345 155.920 ;
        RECT 19.890 155.870 20.150 155.920 ;
        RECT 20.845 155.870 21.105 155.920 ;
        RECT 21.805 155.870 22.065 155.920 ;
        RECT 22.765 155.870 23.025 155.920 ;
        RECT 23.730 155.865 23.990 155.920 ;
        RECT 24.690 155.865 24.950 155.920 ;
        RECT 26.680 151.020 26.950 151.110 ;
        RECT 25.890 150.760 26.950 151.020 ;
        RECT 12.285 149.745 12.545 149.795 ;
        RECT 13.240 149.745 13.500 149.795 ;
        RECT 14.200 149.745 14.460 149.795 ;
        RECT 15.160 149.745 15.420 149.795 ;
        RECT 16.125 149.745 16.385 149.790 ;
        RECT 17.085 149.745 17.345 149.790 ;
        RECT 19.890 149.745 20.150 149.795 ;
        RECT 20.845 149.745 21.105 149.795 ;
        RECT 21.805 149.745 22.065 149.795 ;
        RECT 22.765 149.745 23.025 149.795 ;
        RECT 23.730 149.745 23.990 149.790 ;
        RECT 24.690 149.745 24.950 149.790 ;
        RECT 25.890 149.745 26.150 150.760 ;
        RECT 26.680 150.740 26.950 150.760 ;
        RECT 11.145 149.485 26.150 149.745 ;
        RECT 12.285 149.435 12.545 149.485 ;
        RECT 13.240 149.435 13.500 149.485 ;
        RECT 14.200 149.435 14.460 149.485 ;
        RECT 15.160 149.435 15.420 149.485 ;
        RECT 16.125 149.430 16.385 149.485 ;
        RECT 17.085 149.430 17.345 149.485 ;
        RECT 19.890 149.435 20.150 149.485 ;
        RECT 20.845 149.435 21.105 149.485 ;
        RECT 21.805 149.435 22.065 149.485 ;
        RECT 22.765 149.435 23.025 149.485 ;
        RECT 23.730 149.430 23.990 149.485 ;
        RECT 24.690 149.430 24.950 149.485 ;
        RECT 26.680 144.585 26.950 144.675 ;
        RECT 25.890 144.325 26.950 144.585 ;
        RECT 12.285 143.310 12.545 143.360 ;
        RECT 13.240 143.310 13.500 143.360 ;
        RECT 14.200 143.310 14.460 143.360 ;
        RECT 15.160 143.310 15.420 143.360 ;
        RECT 16.125 143.310 16.385 143.355 ;
        RECT 17.085 143.310 17.345 143.355 ;
        RECT 19.890 143.310 20.150 143.360 ;
        RECT 20.845 143.310 21.105 143.360 ;
        RECT 21.805 143.310 22.065 143.360 ;
        RECT 22.765 143.310 23.025 143.360 ;
        RECT 23.730 143.310 23.990 143.355 ;
        RECT 24.690 143.310 24.950 143.355 ;
        RECT 25.890 143.310 26.150 144.325 ;
        RECT 26.680 144.305 26.950 144.325 ;
        RECT 11.145 143.050 26.150 143.310 ;
        RECT 12.285 143.000 12.545 143.050 ;
        RECT 13.240 143.000 13.500 143.050 ;
        RECT 14.200 143.000 14.460 143.050 ;
        RECT 15.160 143.000 15.420 143.050 ;
        RECT 16.125 142.995 16.385 143.050 ;
        RECT 17.085 142.995 17.345 143.050 ;
        RECT 19.890 143.000 20.150 143.050 ;
        RECT 20.845 143.000 21.105 143.050 ;
        RECT 21.805 143.000 22.065 143.050 ;
        RECT 22.765 143.000 23.025 143.050 ;
        RECT 23.730 142.995 23.990 143.050 ;
        RECT 24.690 142.995 24.950 143.050 ;
        RECT 26.680 138.150 26.950 138.240 ;
        RECT 25.890 137.890 26.950 138.150 ;
        RECT 12.285 136.875 12.545 136.925 ;
        RECT 13.240 136.875 13.500 136.925 ;
        RECT 14.200 136.875 14.460 136.925 ;
        RECT 15.160 136.875 15.420 136.925 ;
        RECT 16.125 136.875 16.385 136.920 ;
        RECT 17.085 136.875 17.345 136.920 ;
        RECT 19.890 136.875 20.150 136.925 ;
        RECT 20.845 136.875 21.105 136.925 ;
        RECT 21.805 136.875 22.065 136.925 ;
        RECT 22.765 136.875 23.025 136.925 ;
        RECT 23.730 136.875 23.990 136.920 ;
        RECT 24.690 136.875 24.950 136.920 ;
        RECT 25.890 136.875 26.150 137.890 ;
        RECT 26.680 137.870 26.950 137.890 ;
        RECT 11.145 136.615 26.150 136.875 ;
        RECT 12.285 136.565 12.545 136.615 ;
        RECT 13.240 136.565 13.500 136.615 ;
        RECT 14.200 136.565 14.460 136.615 ;
        RECT 15.160 136.565 15.420 136.615 ;
        RECT 16.125 136.560 16.385 136.615 ;
        RECT 17.085 136.560 17.345 136.615 ;
        RECT 19.890 136.565 20.150 136.615 ;
        RECT 20.845 136.565 21.105 136.615 ;
        RECT 21.805 136.565 22.065 136.615 ;
        RECT 22.765 136.565 23.025 136.615 ;
        RECT 23.730 136.560 23.990 136.615 ;
        RECT 24.690 136.560 24.950 136.615 ;
        RECT 26.680 131.715 26.950 131.805 ;
        RECT 25.890 131.455 26.950 131.715 ;
        RECT 12.285 130.440 12.545 130.490 ;
        RECT 13.240 130.440 13.500 130.490 ;
        RECT 14.200 130.440 14.460 130.490 ;
        RECT 15.160 130.440 15.420 130.490 ;
        RECT 16.125 130.440 16.385 130.485 ;
        RECT 17.085 130.440 17.345 130.485 ;
        RECT 19.890 130.440 20.150 130.490 ;
        RECT 20.845 130.440 21.105 130.490 ;
        RECT 21.805 130.440 22.065 130.490 ;
        RECT 22.765 130.440 23.025 130.490 ;
        RECT 23.730 130.440 23.990 130.485 ;
        RECT 24.690 130.440 24.950 130.485 ;
        RECT 25.890 130.440 26.150 131.455 ;
        RECT 26.680 131.435 26.950 131.455 ;
        RECT 11.145 130.180 26.150 130.440 ;
        RECT 12.285 130.130 12.545 130.180 ;
        RECT 13.240 130.130 13.500 130.180 ;
        RECT 14.200 130.130 14.460 130.180 ;
        RECT 15.160 130.130 15.420 130.180 ;
        RECT 16.125 130.125 16.385 130.180 ;
        RECT 17.085 130.125 17.345 130.180 ;
        RECT 19.890 130.130 20.150 130.180 ;
        RECT 20.845 130.130 21.105 130.180 ;
        RECT 21.805 130.130 22.065 130.180 ;
        RECT 22.765 130.130 23.025 130.180 ;
        RECT 23.730 130.125 23.990 130.180 ;
        RECT 24.690 130.125 24.950 130.180 ;
        RECT 26.680 125.280 26.950 125.370 ;
        RECT 25.890 125.020 26.950 125.280 ;
        RECT 12.285 124.005 12.545 124.055 ;
        RECT 13.240 124.005 13.500 124.055 ;
        RECT 14.200 124.005 14.460 124.055 ;
        RECT 15.160 124.005 15.420 124.055 ;
        RECT 16.125 124.005 16.385 124.050 ;
        RECT 17.085 124.005 17.345 124.050 ;
        RECT 19.890 124.005 20.150 124.055 ;
        RECT 20.845 124.005 21.105 124.055 ;
        RECT 21.805 124.005 22.065 124.055 ;
        RECT 22.765 124.005 23.025 124.055 ;
        RECT 23.730 124.005 23.990 124.050 ;
        RECT 24.690 124.005 24.950 124.050 ;
        RECT 25.890 124.005 26.150 125.020 ;
        RECT 26.680 125.000 26.950 125.020 ;
        RECT 11.145 123.745 26.150 124.005 ;
        RECT 12.285 123.695 12.545 123.745 ;
        RECT 13.240 123.695 13.500 123.745 ;
        RECT 14.200 123.695 14.460 123.745 ;
        RECT 15.160 123.695 15.420 123.745 ;
        RECT 16.125 123.690 16.385 123.745 ;
        RECT 17.085 123.690 17.345 123.745 ;
        RECT 19.890 123.695 20.150 123.745 ;
        RECT 20.845 123.695 21.105 123.745 ;
        RECT 21.805 123.695 22.065 123.745 ;
        RECT 22.765 123.695 23.025 123.745 ;
        RECT 23.730 123.690 23.990 123.745 ;
        RECT 24.690 123.690 24.950 123.745 ;
        RECT 26.680 118.845 26.950 118.935 ;
        RECT 25.890 118.585 26.950 118.845 ;
        RECT 12.285 117.570 12.545 117.620 ;
        RECT 13.240 117.570 13.500 117.620 ;
        RECT 14.200 117.570 14.460 117.620 ;
        RECT 15.160 117.570 15.420 117.620 ;
        RECT 16.125 117.570 16.385 117.615 ;
        RECT 17.085 117.570 17.345 117.615 ;
        RECT 19.890 117.570 20.150 117.620 ;
        RECT 20.845 117.570 21.105 117.620 ;
        RECT 21.805 117.570 22.065 117.620 ;
        RECT 22.765 117.570 23.025 117.620 ;
        RECT 23.730 117.570 23.990 117.615 ;
        RECT 24.690 117.570 24.950 117.615 ;
        RECT 25.890 117.570 26.150 118.585 ;
        RECT 26.680 118.565 26.950 118.585 ;
        RECT 11.145 117.310 26.150 117.570 ;
        RECT 12.285 117.260 12.545 117.310 ;
        RECT 13.240 117.260 13.500 117.310 ;
        RECT 14.200 117.260 14.460 117.310 ;
        RECT 15.160 117.260 15.420 117.310 ;
        RECT 16.125 117.255 16.385 117.310 ;
        RECT 17.085 117.255 17.345 117.310 ;
        RECT 19.890 117.260 20.150 117.310 ;
        RECT 20.845 117.260 21.105 117.310 ;
        RECT 21.805 117.260 22.065 117.310 ;
        RECT 22.765 117.260 23.025 117.310 ;
        RECT 23.730 117.255 23.990 117.310 ;
        RECT 24.690 117.255 24.950 117.310 ;
        RECT 26.680 112.410 26.950 112.500 ;
        RECT 25.890 112.150 26.950 112.410 ;
        RECT 12.285 111.135 12.545 111.185 ;
        RECT 13.240 111.135 13.500 111.185 ;
        RECT 14.200 111.135 14.460 111.185 ;
        RECT 15.160 111.135 15.420 111.185 ;
        RECT 16.125 111.135 16.385 111.180 ;
        RECT 17.085 111.135 17.345 111.180 ;
        RECT 19.890 111.135 20.150 111.185 ;
        RECT 20.845 111.135 21.105 111.185 ;
        RECT 21.805 111.135 22.065 111.185 ;
        RECT 22.765 111.135 23.025 111.185 ;
        RECT 23.730 111.135 23.990 111.180 ;
        RECT 24.690 111.135 24.950 111.180 ;
        RECT 25.890 111.135 26.150 112.150 ;
        RECT 26.680 112.130 26.950 112.150 ;
        RECT 11.145 110.875 26.150 111.135 ;
        RECT 12.285 110.825 12.545 110.875 ;
        RECT 13.240 110.825 13.500 110.875 ;
        RECT 14.200 110.825 14.460 110.875 ;
        RECT 15.160 110.825 15.420 110.875 ;
        RECT 16.125 110.820 16.385 110.875 ;
        RECT 17.085 110.820 17.345 110.875 ;
        RECT 19.890 110.825 20.150 110.875 ;
        RECT 20.845 110.825 21.105 110.875 ;
        RECT 21.805 110.825 22.065 110.875 ;
        RECT 22.765 110.825 23.025 110.875 ;
        RECT 23.730 110.820 23.990 110.875 ;
        RECT 24.690 110.820 24.950 110.875 ;
        RECT 26.680 105.975 26.950 106.065 ;
        RECT 25.890 105.715 26.950 105.975 ;
        RECT 12.285 104.700 12.545 104.750 ;
        RECT 13.240 104.700 13.500 104.750 ;
        RECT 14.200 104.700 14.460 104.750 ;
        RECT 15.160 104.700 15.420 104.750 ;
        RECT 16.125 104.700 16.385 104.745 ;
        RECT 17.085 104.700 17.345 104.745 ;
        RECT 19.890 104.700 20.150 104.750 ;
        RECT 20.845 104.700 21.105 104.750 ;
        RECT 21.805 104.700 22.065 104.750 ;
        RECT 22.765 104.700 23.025 104.750 ;
        RECT 23.730 104.700 23.990 104.745 ;
        RECT 24.690 104.700 24.950 104.745 ;
        RECT 25.890 104.700 26.150 105.715 ;
        RECT 26.680 105.695 26.950 105.715 ;
        RECT 11.145 104.440 26.150 104.700 ;
        RECT 12.285 104.390 12.545 104.440 ;
        RECT 13.240 104.390 13.500 104.440 ;
        RECT 14.200 104.390 14.460 104.440 ;
        RECT 15.160 104.390 15.420 104.440 ;
        RECT 16.125 104.385 16.385 104.440 ;
        RECT 17.085 104.385 17.345 104.440 ;
        RECT 19.890 104.390 20.150 104.440 ;
        RECT 20.845 104.390 21.105 104.440 ;
        RECT 21.805 104.390 22.065 104.440 ;
        RECT 22.765 104.390 23.025 104.440 ;
        RECT 23.730 104.385 23.990 104.440 ;
        RECT 24.690 104.385 24.950 104.440 ;
        RECT 26.680 99.540 26.950 99.630 ;
        RECT 25.890 99.280 26.950 99.540 ;
        RECT 12.285 98.265 12.545 98.315 ;
        RECT 13.240 98.265 13.500 98.315 ;
        RECT 14.200 98.265 14.460 98.315 ;
        RECT 15.160 98.265 15.420 98.315 ;
        RECT 16.125 98.265 16.385 98.310 ;
        RECT 17.085 98.265 17.345 98.310 ;
        RECT 19.890 98.265 20.150 98.315 ;
        RECT 20.845 98.265 21.105 98.315 ;
        RECT 21.805 98.265 22.065 98.315 ;
        RECT 22.765 98.265 23.025 98.315 ;
        RECT 23.730 98.265 23.990 98.310 ;
        RECT 24.690 98.265 24.950 98.310 ;
        RECT 25.890 98.265 26.150 99.280 ;
        RECT 26.680 99.260 26.950 99.280 ;
        RECT 11.145 98.005 26.150 98.265 ;
        RECT 12.285 97.955 12.545 98.005 ;
        RECT 13.240 97.955 13.500 98.005 ;
        RECT 14.200 97.955 14.460 98.005 ;
        RECT 15.160 97.955 15.420 98.005 ;
        RECT 16.125 97.950 16.385 98.005 ;
        RECT 17.085 97.950 17.345 98.005 ;
        RECT 19.890 97.955 20.150 98.005 ;
        RECT 20.845 97.955 21.105 98.005 ;
        RECT 21.805 97.955 22.065 98.005 ;
        RECT 22.765 97.955 23.025 98.005 ;
        RECT 23.730 97.950 23.990 98.005 ;
        RECT 24.690 97.950 24.950 98.005 ;
        RECT 26.680 93.105 26.950 93.195 ;
        RECT 25.890 92.845 26.950 93.105 ;
        RECT 12.285 91.830 12.545 91.880 ;
        RECT 13.240 91.830 13.500 91.880 ;
        RECT 14.200 91.830 14.460 91.880 ;
        RECT 15.160 91.830 15.420 91.880 ;
        RECT 16.125 91.830 16.385 91.875 ;
        RECT 17.085 91.830 17.345 91.875 ;
        RECT 19.890 91.830 20.150 91.880 ;
        RECT 20.845 91.830 21.105 91.880 ;
        RECT 21.805 91.830 22.065 91.880 ;
        RECT 22.765 91.830 23.025 91.880 ;
        RECT 23.730 91.830 23.990 91.875 ;
        RECT 24.690 91.830 24.950 91.875 ;
        RECT 25.890 91.830 26.150 92.845 ;
        RECT 26.680 92.825 26.950 92.845 ;
        RECT 11.145 91.570 26.150 91.830 ;
        RECT 12.285 91.520 12.545 91.570 ;
        RECT 13.240 91.520 13.500 91.570 ;
        RECT 14.200 91.520 14.460 91.570 ;
        RECT 15.160 91.520 15.420 91.570 ;
        RECT 16.125 91.515 16.385 91.570 ;
        RECT 17.085 91.515 17.345 91.570 ;
        RECT 19.890 91.520 20.150 91.570 ;
        RECT 20.845 91.520 21.105 91.570 ;
        RECT 21.805 91.520 22.065 91.570 ;
        RECT 22.765 91.520 23.025 91.570 ;
        RECT 23.730 91.515 23.990 91.570 ;
        RECT 24.690 91.515 24.950 91.570 ;
        RECT 26.680 86.670 26.950 86.760 ;
        RECT 25.890 86.410 26.950 86.670 ;
        RECT 12.285 85.395 12.545 85.445 ;
        RECT 13.240 85.395 13.500 85.445 ;
        RECT 14.200 85.395 14.460 85.445 ;
        RECT 15.160 85.395 15.420 85.445 ;
        RECT 16.125 85.395 16.385 85.440 ;
        RECT 17.085 85.395 17.345 85.440 ;
        RECT 19.890 85.395 20.150 85.445 ;
        RECT 20.845 85.395 21.105 85.445 ;
        RECT 21.805 85.395 22.065 85.445 ;
        RECT 22.765 85.395 23.025 85.445 ;
        RECT 23.730 85.395 23.990 85.440 ;
        RECT 24.690 85.395 24.950 85.440 ;
        RECT 25.890 85.395 26.150 86.410 ;
        RECT 26.680 86.390 26.950 86.410 ;
        RECT 11.145 85.135 26.150 85.395 ;
        RECT 12.285 85.085 12.545 85.135 ;
        RECT 13.240 85.085 13.500 85.135 ;
        RECT 14.200 85.085 14.460 85.135 ;
        RECT 15.160 85.085 15.420 85.135 ;
        RECT 16.125 85.080 16.385 85.135 ;
        RECT 17.085 85.080 17.345 85.135 ;
        RECT 19.890 85.085 20.150 85.135 ;
        RECT 20.845 85.085 21.105 85.135 ;
        RECT 21.805 85.085 22.065 85.135 ;
        RECT 22.765 85.085 23.025 85.135 ;
        RECT 23.730 85.080 23.990 85.135 ;
        RECT 24.690 85.080 24.950 85.135 ;
        RECT 26.680 80.235 26.950 80.325 ;
        RECT 25.890 79.975 26.950 80.235 ;
        RECT 12.285 78.960 12.545 79.010 ;
        RECT 13.240 78.960 13.500 79.010 ;
        RECT 14.200 78.960 14.460 79.010 ;
        RECT 15.160 78.960 15.420 79.010 ;
        RECT 16.125 78.960 16.385 79.005 ;
        RECT 17.085 78.960 17.345 79.005 ;
        RECT 19.890 78.960 20.150 79.010 ;
        RECT 20.845 78.960 21.105 79.010 ;
        RECT 21.805 78.960 22.065 79.010 ;
        RECT 22.765 78.960 23.025 79.010 ;
        RECT 23.730 78.960 23.990 79.005 ;
        RECT 24.690 78.960 24.950 79.005 ;
        RECT 25.890 78.960 26.150 79.975 ;
        RECT 26.680 79.955 26.950 79.975 ;
        RECT 11.145 78.700 26.150 78.960 ;
        RECT 12.285 78.650 12.545 78.700 ;
        RECT 13.240 78.650 13.500 78.700 ;
        RECT 14.200 78.650 14.460 78.700 ;
        RECT 15.160 78.650 15.420 78.700 ;
        RECT 16.125 78.645 16.385 78.700 ;
        RECT 17.085 78.645 17.345 78.700 ;
        RECT 19.890 78.650 20.150 78.700 ;
        RECT 20.845 78.650 21.105 78.700 ;
        RECT 21.805 78.650 22.065 78.700 ;
        RECT 22.765 78.650 23.025 78.700 ;
        RECT 23.730 78.645 23.990 78.700 ;
        RECT 24.690 78.645 24.950 78.700 ;
        RECT 26.680 73.800 26.950 73.890 ;
        RECT 25.890 73.540 26.950 73.800 ;
        RECT 12.285 72.525 12.545 72.575 ;
        RECT 13.240 72.525 13.500 72.575 ;
        RECT 14.200 72.525 14.460 72.575 ;
        RECT 15.160 72.525 15.420 72.575 ;
        RECT 16.125 72.525 16.385 72.570 ;
        RECT 17.085 72.525 17.345 72.570 ;
        RECT 19.890 72.525 20.150 72.575 ;
        RECT 20.845 72.525 21.105 72.575 ;
        RECT 21.805 72.525 22.065 72.575 ;
        RECT 22.765 72.525 23.025 72.575 ;
        RECT 23.730 72.525 23.990 72.570 ;
        RECT 24.690 72.525 24.950 72.570 ;
        RECT 25.890 72.525 26.150 73.540 ;
        RECT 26.680 73.520 26.950 73.540 ;
        RECT 11.145 72.265 26.150 72.525 ;
        RECT 12.285 72.215 12.545 72.265 ;
        RECT 13.240 72.215 13.500 72.265 ;
        RECT 14.200 72.215 14.460 72.265 ;
        RECT 15.160 72.215 15.420 72.265 ;
        RECT 16.125 72.210 16.385 72.265 ;
        RECT 17.085 72.210 17.345 72.265 ;
        RECT 19.890 72.215 20.150 72.265 ;
        RECT 20.845 72.215 21.105 72.265 ;
        RECT 21.805 72.215 22.065 72.265 ;
        RECT 22.765 72.215 23.025 72.265 ;
        RECT 23.730 72.210 23.990 72.265 ;
        RECT 24.690 72.210 24.950 72.265 ;
        RECT 26.680 67.365 26.950 67.455 ;
        RECT 25.890 67.105 26.950 67.365 ;
        RECT 12.285 66.090 12.545 66.140 ;
        RECT 13.240 66.090 13.500 66.140 ;
        RECT 14.200 66.090 14.460 66.140 ;
        RECT 15.160 66.090 15.420 66.140 ;
        RECT 16.125 66.090 16.385 66.135 ;
        RECT 17.085 66.090 17.345 66.135 ;
        RECT 19.890 66.090 20.150 66.140 ;
        RECT 20.845 66.090 21.105 66.140 ;
        RECT 21.805 66.090 22.065 66.140 ;
        RECT 22.765 66.090 23.025 66.140 ;
        RECT 23.730 66.090 23.990 66.135 ;
        RECT 24.690 66.090 24.950 66.135 ;
        RECT 25.890 66.090 26.150 67.105 ;
        RECT 26.680 67.085 26.950 67.105 ;
        RECT 11.145 65.830 26.150 66.090 ;
        RECT 12.285 65.780 12.545 65.830 ;
        RECT 13.240 65.780 13.500 65.830 ;
        RECT 14.200 65.780 14.460 65.830 ;
        RECT 15.160 65.780 15.420 65.830 ;
        RECT 16.125 65.775 16.385 65.830 ;
        RECT 17.085 65.775 17.345 65.830 ;
        RECT 19.890 65.780 20.150 65.830 ;
        RECT 20.845 65.780 21.105 65.830 ;
        RECT 21.805 65.780 22.065 65.830 ;
        RECT 22.765 65.780 23.025 65.830 ;
        RECT 23.730 65.775 23.990 65.830 ;
        RECT 24.690 65.775 24.950 65.830 ;
        RECT 26.680 60.930 26.950 61.020 ;
        RECT 25.890 60.670 26.950 60.930 ;
        RECT 12.285 59.655 12.545 59.705 ;
        RECT 13.240 59.655 13.500 59.705 ;
        RECT 14.200 59.655 14.460 59.705 ;
        RECT 15.160 59.655 15.420 59.705 ;
        RECT 16.125 59.655 16.385 59.700 ;
        RECT 17.085 59.655 17.345 59.700 ;
        RECT 19.890 59.655 20.150 59.705 ;
        RECT 20.845 59.655 21.105 59.705 ;
        RECT 21.805 59.655 22.065 59.705 ;
        RECT 22.765 59.655 23.025 59.705 ;
        RECT 23.730 59.655 23.990 59.700 ;
        RECT 24.690 59.655 24.950 59.700 ;
        RECT 25.890 59.655 26.150 60.670 ;
        RECT 26.680 60.650 26.950 60.670 ;
        RECT 11.145 59.395 26.150 59.655 ;
        RECT 12.285 59.345 12.545 59.395 ;
        RECT 13.240 59.345 13.500 59.395 ;
        RECT 14.200 59.345 14.460 59.395 ;
        RECT 15.160 59.345 15.420 59.395 ;
        RECT 16.125 59.340 16.385 59.395 ;
        RECT 17.085 59.340 17.345 59.395 ;
        RECT 19.890 59.345 20.150 59.395 ;
        RECT 20.845 59.345 21.105 59.395 ;
        RECT 21.805 59.345 22.065 59.395 ;
        RECT 22.765 59.345 23.025 59.395 ;
        RECT 23.730 59.340 23.990 59.395 ;
        RECT 24.690 59.340 24.950 59.395 ;
        RECT 26.680 54.495 26.950 54.585 ;
        RECT 25.890 54.235 26.950 54.495 ;
        RECT 12.285 53.220 12.545 53.270 ;
        RECT 13.240 53.220 13.500 53.270 ;
        RECT 14.200 53.220 14.460 53.270 ;
        RECT 15.160 53.220 15.420 53.270 ;
        RECT 16.125 53.220 16.385 53.265 ;
        RECT 17.085 53.220 17.345 53.265 ;
        RECT 19.890 53.220 20.150 53.270 ;
        RECT 20.845 53.220 21.105 53.270 ;
        RECT 21.805 53.220 22.065 53.270 ;
        RECT 22.765 53.220 23.025 53.270 ;
        RECT 23.730 53.220 23.990 53.265 ;
        RECT 24.690 53.220 24.950 53.265 ;
        RECT 25.890 53.220 26.150 54.235 ;
        RECT 26.680 54.215 26.950 54.235 ;
        RECT 11.145 52.960 26.150 53.220 ;
        RECT 12.285 52.910 12.545 52.960 ;
        RECT 13.240 52.910 13.500 52.960 ;
        RECT 14.200 52.910 14.460 52.960 ;
        RECT 15.160 52.910 15.420 52.960 ;
        RECT 16.125 52.905 16.385 52.960 ;
        RECT 17.085 52.905 17.345 52.960 ;
        RECT 19.890 52.910 20.150 52.960 ;
        RECT 20.845 52.910 21.105 52.960 ;
        RECT 21.805 52.910 22.065 52.960 ;
        RECT 22.765 52.910 23.025 52.960 ;
        RECT 23.730 52.905 23.990 52.960 ;
        RECT 24.690 52.905 24.950 52.960 ;
        RECT 26.680 48.060 26.950 48.150 ;
        RECT 25.890 47.800 26.950 48.060 ;
        RECT 12.285 46.785 12.545 46.835 ;
        RECT 13.240 46.785 13.500 46.835 ;
        RECT 14.200 46.785 14.460 46.835 ;
        RECT 15.160 46.785 15.420 46.835 ;
        RECT 16.125 46.785 16.385 46.830 ;
        RECT 17.085 46.785 17.345 46.830 ;
        RECT 19.890 46.785 20.150 46.835 ;
        RECT 20.845 46.785 21.105 46.835 ;
        RECT 21.805 46.785 22.065 46.835 ;
        RECT 22.765 46.785 23.025 46.835 ;
        RECT 23.730 46.785 23.990 46.830 ;
        RECT 24.690 46.785 24.950 46.830 ;
        RECT 25.890 46.785 26.150 47.800 ;
        RECT 26.680 47.780 26.950 47.800 ;
        RECT 11.145 46.525 26.150 46.785 ;
        RECT 12.285 46.475 12.545 46.525 ;
        RECT 13.240 46.475 13.500 46.525 ;
        RECT 14.200 46.475 14.460 46.525 ;
        RECT 15.160 46.475 15.420 46.525 ;
        RECT 16.125 46.470 16.385 46.525 ;
        RECT 17.085 46.470 17.345 46.525 ;
        RECT 19.890 46.475 20.150 46.525 ;
        RECT 20.845 46.475 21.105 46.525 ;
        RECT 21.805 46.475 22.065 46.525 ;
        RECT 22.765 46.475 23.025 46.525 ;
        RECT 23.730 46.470 23.990 46.525 ;
        RECT 24.690 46.470 24.950 46.525 ;
        RECT 26.680 41.625 26.950 41.715 ;
        RECT 25.890 41.365 26.950 41.625 ;
        RECT 12.285 40.350 12.545 40.400 ;
        RECT 13.240 40.350 13.500 40.400 ;
        RECT 14.200 40.350 14.460 40.400 ;
        RECT 15.160 40.350 15.420 40.400 ;
        RECT 16.125 40.350 16.385 40.395 ;
        RECT 17.085 40.350 17.345 40.395 ;
        RECT 19.890 40.350 20.150 40.400 ;
        RECT 20.845 40.350 21.105 40.400 ;
        RECT 21.805 40.350 22.065 40.400 ;
        RECT 22.765 40.350 23.025 40.400 ;
        RECT 23.730 40.350 23.990 40.395 ;
        RECT 24.690 40.350 24.950 40.395 ;
        RECT 25.890 40.350 26.150 41.365 ;
        RECT 26.680 41.345 26.950 41.365 ;
        RECT 11.145 40.090 26.150 40.350 ;
        RECT 12.285 40.040 12.545 40.090 ;
        RECT 13.240 40.040 13.500 40.090 ;
        RECT 14.200 40.040 14.460 40.090 ;
        RECT 15.160 40.040 15.420 40.090 ;
        RECT 16.125 40.035 16.385 40.090 ;
        RECT 17.085 40.035 17.345 40.090 ;
        RECT 19.890 40.040 20.150 40.090 ;
        RECT 20.845 40.040 21.105 40.090 ;
        RECT 21.805 40.040 22.065 40.090 ;
        RECT 22.765 40.040 23.025 40.090 ;
        RECT 23.730 40.035 23.990 40.090 ;
        RECT 24.690 40.035 24.950 40.090 ;
        RECT 26.680 35.190 26.950 35.280 ;
        RECT 25.890 34.930 26.950 35.190 ;
        RECT 12.285 33.915 12.545 33.965 ;
        RECT 13.240 33.915 13.500 33.965 ;
        RECT 14.200 33.915 14.460 33.965 ;
        RECT 15.160 33.915 15.420 33.965 ;
        RECT 16.125 33.915 16.385 33.960 ;
        RECT 17.085 33.915 17.345 33.960 ;
        RECT 19.890 33.915 20.150 33.965 ;
        RECT 20.845 33.915 21.105 33.965 ;
        RECT 21.805 33.915 22.065 33.965 ;
        RECT 22.765 33.915 23.025 33.965 ;
        RECT 23.730 33.915 23.990 33.960 ;
        RECT 24.690 33.915 24.950 33.960 ;
        RECT 25.890 33.915 26.150 34.930 ;
        RECT 26.680 34.910 26.950 34.930 ;
        RECT 11.145 33.655 26.150 33.915 ;
        RECT 12.285 33.605 12.545 33.655 ;
        RECT 13.240 33.605 13.500 33.655 ;
        RECT 14.200 33.605 14.460 33.655 ;
        RECT 15.160 33.605 15.420 33.655 ;
        RECT 16.125 33.600 16.385 33.655 ;
        RECT 17.085 33.600 17.345 33.655 ;
        RECT 19.890 33.605 20.150 33.655 ;
        RECT 20.845 33.605 21.105 33.655 ;
        RECT 21.805 33.605 22.065 33.655 ;
        RECT 22.765 33.605 23.025 33.655 ;
        RECT 23.730 33.600 23.990 33.655 ;
        RECT 24.690 33.600 24.950 33.655 ;
        RECT 26.680 28.755 26.950 28.845 ;
        RECT 25.890 28.495 26.950 28.755 ;
        RECT 12.285 27.480 12.545 27.530 ;
        RECT 13.240 27.480 13.500 27.530 ;
        RECT 14.200 27.480 14.460 27.530 ;
        RECT 15.160 27.480 15.420 27.530 ;
        RECT 16.125 27.480 16.385 27.525 ;
        RECT 17.085 27.480 17.345 27.525 ;
        RECT 19.890 27.480 20.150 27.530 ;
        RECT 20.845 27.480 21.105 27.530 ;
        RECT 21.805 27.480 22.065 27.530 ;
        RECT 22.765 27.480 23.025 27.530 ;
        RECT 23.730 27.480 23.990 27.525 ;
        RECT 24.690 27.480 24.950 27.525 ;
        RECT 25.890 27.480 26.150 28.495 ;
        RECT 26.680 28.475 26.950 28.495 ;
        RECT 11.145 27.220 26.150 27.480 ;
        RECT 12.285 27.170 12.545 27.220 ;
        RECT 13.240 27.170 13.500 27.220 ;
        RECT 14.200 27.170 14.460 27.220 ;
        RECT 15.160 27.170 15.420 27.220 ;
        RECT 16.125 27.165 16.385 27.220 ;
        RECT 17.085 27.165 17.345 27.220 ;
        RECT 19.890 27.170 20.150 27.220 ;
        RECT 20.845 27.170 21.105 27.220 ;
        RECT 21.805 27.170 22.065 27.220 ;
        RECT 22.765 27.170 23.025 27.220 ;
        RECT 23.730 27.165 23.990 27.220 ;
        RECT 24.690 27.165 24.950 27.220 ;
        RECT 26.680 22.320 26.950 22.410 ;
        RECT 25.890 22.060 26.950 22.320 ;
        RECT 12.285 21.045 12.545 21.095 ;
        RECT 13.240 21.045 13.500 21.095 ;
        RECT 14.200 21.045 14.460 21.095 ;
        RECT 15.160 21.045 15.420 21.095 ;
        RECT 16.125 21.045 16.385 21.090 ;
        RECT 17.085 21.045 17.345 21.090 ;
        RECT 19.890 21.045 20.150 21.095 ;
        RECT 20.845 21.045 21.105 21.095 ;
        RECT 21.805 21.045 22.065 21.095 ;
        RECT 22.765 21.045 23.025 21.095 ;
        RECT 23.730 21.045 23.990 21.090 ;
        RECT 24.690 21.045 24.950 21.090 ;
        RECT 25.890 21.045 26.150 22.060 ;
        RECT 26.680 22.040 26.950 22.060 ;
        RECT 11.145 20.785 26.150 21.045 ;
        RECT 12.285 20.735 12.545 20.785 ;
        RECT 13.240 20.735 13.500 20.785 ;
        RECT 14.200 20.735 14.460 20.785 ;
        RECT 15.160 20.735 15.420 20.785 ;
        RECT 16.125 20.730 16.385 20.785 ;
        RECT 17.085 20.730 17.345 20.785 ;
        RECT 19.890 20.735 20.150 20.785 ;
        RECT 20.845 20.735 21.105 20.785 ;
        RECT 21.805 20.735 22.065 20.785 ;
        RECT 22.765 20.735 23.025 20.785 ;
        RECT 23.730 20.730 23.990 20.785 ;
        RECT 24.690 20.730 24.950 20.785 ;
        RECT 26.680 15.885 26.950 15.975 ;
        RECT 25.890 15.625 26.950 15.885 ;
        RECT 12.285 14.610 12.545 14.660 ;
        RECT 13.240 14.610 13.500 14.660 ;
        RECT 14.200 14.610 14.460 14.660 ;
        RECT 15.160 14.610 15.420 14.660 ;
        RECT 16.125 14.610 16.385 14.655 ;
        RECT 17.085 14.610 17.345 14.655 ;
        RECT 19.890 14.610 20.150 14.660 ;
        RECT 20.845 14.610 21.105 14.660 ;
        RECT 21.805 14.610 22.065 14.660 ;
        RECT 22.765 14.610 23.025 14.660 ;
        RECT 23.730 14.610 23.990 14.655 ;
        RECT 24.690 14.610 24.950 14.655 ;
        RECT 25.890 14.610 26.150 15.625 ;
        RECT 26.680 15.605 26.950 15.625 ;
        RECT 11.145 14.350 26.150 14.610 ;
        RECT 12.285 14.300 12.545 14.350 ;
        RECT 13.240 14.300 13.500 14.350 ;
        RECT 14.200 14.300 14.460 14.350 ;
        RECT 15.160 14.300 15.420 14.350 ;
        RECT 16.125 14.295 16.385 14.350 ;
        RECT 17.085 14.295 17.345 14.350 ;
        RECT 19.890 14.300 20.150 14.350 ;
        RECT 20.845 14.300 21.105 14.350 ;
        RECT 21.805 14.300 22.065 14.350 ;
        RECT 22.765 14.300 23.025 14.350 ;
        RECT 23.730 14.295 23.990 14.350 ;
        RECT 24.690 14.295 24.950 14.350 ;
        RECT 26.680 9.450 26.950 9.540 ;
        RECT 25.890 9.190 26.950 9.450 ;
        RECT 12.285 8.175 12.545 8.225 ;
        RECT 13.240 8.175 13.500 8.225 ;
        RECT 14.200 8.175 14.460 8.225 ;
        RECT 15.160 8.175 15.420 8.225 ;
        RECT 16.125 8.175 16.385 8.220 ;
        RECT 17.085 8.175 17.345 8.220 ;
        RECT 19.890 8.175 20.150 8.225 ;
        RECT 20.845 8.175 21.105 8.225 ;
        RECT 21.805 8.175 22.065 8.225 ;
        RECT 22.765 8.175 23.025 8.225 ;
        RECT 23.730 8.175 23.990 8.220 ;
        RECT 24.690 8.175 24.950 8.220 ;
        RECT 25.890 8.175 26.150 9.190 ;
        RECT 26.680 9.170 26.950 9.190 ;
        RECT 11.145 7.915 26.150 8.175 ;
        RECT 12.285 7.865 12.545 7.915 ;
        RECT 13.240 7.865 13.500 7.915 ;
        RECT 14.200 7.865 14.460 7.915 ;
        RECT 15.160 7.865 15.420 7.915 ;
        RECT 16.125 7.860 16.385 7.915 ;
        RECT 17.085 7.860 17.345 7.915 ;
        RECT 19.890 7.865 20.150 7.915 ;
        RECT 20.845 7.865 21.105 7.915 ;
        RECT 21.805 7.865 22.065 7.915 ;
        RECT 22.765 7.865 23.025 7.915 ;
        RECT 23.730 7.860 23.990 7.915 ;
        RECT 24.690 7.860 24.950 7.915 ;
        RECT 26.680 3.015 26.950 3.105 ;
        RECT 25.890 2.755 26.950 3.015 ;
        RECT 12.285 1.740 12.545 1.790 ;
        RECT 13.240 1.740 13.500 1.790 ;
        RECT 14.200 1.740 14.460 1.790 ;
        RECT 15.160 1.740 15.420 1.790 ;
        RECT 16.125 1.740 16.385 1.785 ;
        RECT 17.085 1.740 17.345 1.785 ;
        RECT 19.890 1.740 20.150 1.790 ;
        RECT 20.845 1.740 21.105 1.790 ;
        RECT 21.805 1.740 22.065 1.790 ;
        RECT 22.765 1.740 23.025 1.790 ;
        RECT 23.730 1.740 23.990 1.785 ;
        RECT 24.690 1.740 24.950 1.785 ;
        RECT 25.890 1.740 26.150 2.755 ;
        RECT 26.680 2.735 26.950 2.755 ;
        RECT 11.145 1.480 26.150 1.740 ;
        RECT 12.285 1.430 12.545 1.480 ;
        RECT 13.240 1.430 13.500 1.480 ;
        RECT 14.200 1.430 14.460 1.480 ;
        RECT 15.160 1.430 15.420 1.480 ;
        RECT 16.125 1.425 16.385 1.480 ;
        RECT 17.085 1.425 17.345 1.480 ;
        RECT 19.890 1.430 20.150 1.480 ;
        RECT 20.845 1.430 21.105 1.480 ;
        RECT 21.805 1.430 22.065 1.480 ;
        RECT 22.765 1.430 23.025 1.480 ;
        RECT 23.730 1.425 23.990 1.480 ;
        RECT 24.690 1.425 24.950 1.480 ;
  END
END switch
END LIBRARY

