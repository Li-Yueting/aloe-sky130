magic
tech sky130A
magscale 1 2
timestamp 1622522911
<< pwell >>
rect -2747 -679 2747 679
<< nmoslvt >>
rect -2551 -531 -2351 469
rect -2293 -531 -2093 469
rect -2035 -531 -1835 469
rect -1777 -531 -1577 469
rect -1519 -531 -1319 469
rect -1261 -531 -1061 469
rect -1003 -531 -803 469
rect -745 -531 -545 469
rect -487 -531 -287 469
rect -229 -531 -29 469
rect 29 -531 229 469
rect 287 -531 487 469
rect 545 -531 745 469
rect 803 -531 1003 469
rect 1061 -531 1261 469
rect 1319 -531 1519 469
rect 1577 -531 1777 469
rect 1835 -531 2035 469
rect 2093 -531 2293 469
rect 2351 -531 2551 469
<< ndiff >>
rect -2609 457 -2551 469
rect -2609 -519 -2597 457
rect -2563 -519 -2551 457
rect -2609 -531 -2551 -519
rect -2351 457 -2293 469
rect -2351 -519 -2339 457
rect -2305 -519 -2293 457
rect -2351 -531 -2293 -519
rect -2093 457 -2035 469
rect -2093 -519 -2081 457
rect -2047 -519 -2035 457
rect -2093 -531 -2035 -519
rect -1835 457 -1777 469
rect -1835 -519 -1823 457
rect -1789 -519 -1777 457
rect -1835 -531 -1777 -519
rect -1577 457 -1519 469
rect -1577 -519 -1565 457
rect -1531 -519 -1519 457
rect -1577 -531 -1519 -519
rect -1319 457 -1261 469
rect -1319 -519 -1307 457
rect -1273 -519 -1261 457
rect -1319 -531 -1261 -519
rect -1061 457 -1003 469
rect -1061 -519 -1049 457
rect -1015 -519 -1003 457
rect -1061 -531 -1003 -519
rect -803 457 -745 469
rect -803 -519 -791 457
rect -757 -519 -745 457
rect -803 -531 -745 -519
rect -545 457 -487 469
rect -545 -519 -533 457
rect -499 -519 -487 457
rect -545 -531 -487 -519
rect -287 457 -229 469
rect -287 -519 -275 457
rect -241 -519 -229 457
rect -287 -531 -229 -519
rect -29 457 29 469
rect -29 -519 -17 457
rect 17 -519 29 457
rect -29 -531 29 -519
rect 229 457 287 469
rect 229 -519 241 457
rect 275 -519 287 457
rect 229 -531 287 -519
rect 487 457 545 469
rect 487 -519 499 457
rect 533 -519 545 457
rect 487 -531 545 -519
rect 745 457 803 469
rect 745 -519 757 457
rect 791 -519 803 457
rect 745 -531 803 -519
rect 1003 457 1061 469
rect 1003 -519 1015 457
rect 1049 -519 1061 457
rect 1003 -531 1061 -519
rect 1261 457 1319 469
rect 1261 -519 1273 457
rect 1307 -519 1319 457
rect 1261 -531 1319 -519
rect 1519 457 1577 469
rect 1519 -519 1531 457
rect 1565 -519 1577 457
rect 1519 -531 1577 -519
rect 1777 457 1835 469
rect 1777 -519 1789 457
rect 1823 -519 1835 457
rect 1777 -531 1835 -519
rect 2035 457 2093 469
rect 2035 -519 2047 457
rect 2081 -519 2093 457
rect 2035 -531 2093 -519
rect 2293 457 2351 469
rect 2293 -519 2305 457
rect 2339 -519 2351 457
rect 2293 -531 2351 -519
rect 2551 457 2609 469
rect 2551 -519 2563 457
rect 2597 -519 2609 457
rect 2551 -531 2609 -519
<< ndiffc >>
rect -2597 -519 -2563 457
rect -2339 -519 -2305 457
rect -2081 -519 -2047 457
rect -1823 -519 -1789 457
rect -1565 -519 -1531 457
rect -1307 -519 -1273 457
rect -1049 -519 -1015 457
rect -791 -519 -757 457
rect -533 -519 -499 457
rect -275 -519 -241 457
rect -17 -519 17 457
rect 241 -519 275 457
rect 499 -519 533 457
rect 757 -519 791 457
rect 1015 -519 1049 457
rect 1273 -519 1307 457
rect 1531 -519 1565 457
rect 1789 -519 1823 457
rect 2047 -519 2081 457
rect 2305 -519 2339 457
rect 2563 -519 2597 457
<< psubdiff >>
rect -2711 609 -2615 643
rect 2615 609 2711 643
rect -2711 547 -2677 609
rect 2677 547 2711 609
rect -2711 -609 -2677 -547
rect 2677 -609 2711 -547
rect -2711 -643 -2615 -609
rect 2615 -643 2711 -609
<< psubdiffcont >>
rect -2615 609 2615 643
rect -2711 -547 -2677 547
rect 2677 -547 2711 547
rect -2615 -643 2615 -609
<< poly >>
rect -2551 541 -2351 557
rect -2551 507 -2535 541
rect -2367 507 -2351 541
rect -2551 469 -2351 507
rect -2293 541 -2093 557
rect -2293 507 -2277 541
rect -2109 507 -2093 541
rect -2293 469 -2093 507
rect -2035 541 -1835 557
rect -2035 507 -2019 541
rect -1851 507 -1835 541
rect -2035 469 -1835 507
rect -1777 541 -1577 557
rect -1777 507 -1761 541
rect -1593 507 -1577 541
rect -1777 469 -1577 507
rect -1519 541 -1319 557
rect -1519 507 -1503 541
rect -1335 507 -1319 541
rect -1519 469 -1319 507
rect -1261 541 -1061 557
rect -1261 507 -1245 541
rect -1077 507 -1061 541
rect -1261 469 -1061 507
rect -1003 541 -803 557
rect -1003 507 -987 541
rect -819 507 -803 541
rect -1003 469 -803 507
rect -745 541 -545 557
rect -745 507 -729 541
rect -561 507 -545 541
rect -745 469 -545 507
rect -487 541 -287 557
rect -487 507 -471 541
rect -303 507 -287 541
rect -487 469 -287 507
rect -229 541 -29 557
rect -229 507 -213 541
rect -45 507 -29 541
rect -229 469 -29 507
rect 29 541 229 557
rect 29 507 45 541
rect 213 507 229 541
rect 29 469 229 507
rect 287 541 487 557
rect 287 507 303 541
rect 471 507 487 541
rect 287 469 487 507
rect 545 541 745 557
rect 545 507 561 541
rect 729 507 745 541
rect 545 469 745 507
rect 803 541 1003 557
rect 803 507 819 541
rect 987 507 1003 541
rect 803 469 1003 507
rect 1061 541 1261 557
rect 1061 507 1077 541
rect 1245 507 1261 541
rect 1061 469 1261 507
rect 1319 541 1519 557
rect 1319 507 1335 541
rect 1503 507 1519 541
rect 1319 469 1519 507
rect 1577 541 1777 557
rect 1577 507 1593 541
rect 1761 507 1777 541
rect 1577 469 1777 507
rect 1835 541 2035 557
rect 1835 507 1851 541
rect 2019 507 2035 541
rect 1835 469 2035 507
rect 2093 541 2293 557
rect 2093 507 2109 541
rect 2277 507 2293 541
rect 2093 469 2293 507
rect 2351 541 2551 557
rect 2351 507 2367 541
rect 2535 507 2551 541
rect 2351 469 2551 507
rect -2551 -557 -2351 -531
rect -2293 -557 -2093 -531
rect -2035 -557 -1835 -531
rect -1777 -557 -1577 -531
rect -1519 -557 -1319 -531
rect -1261 -557 -1061 -531
rect -1003 -557 -803 -531
rect -745 -557 -545 -531
rect -487 -557 -287 -531
rect -229 -557 -29 -531
rect 29 -557 229 -531
rect 287 -557 487 -531
rect 545 -557 745 -531
rect 803 -557 1003 -531
rect 1061 -557 1261 -531
rect 1319 -557 1519 -531
rect 1577 -557 1777 -531
rect 1835 -557 2035 -531
rect 2093 -557 2293 -531
rect 2351 -557 2551 -531
<< polycont >>
rect -2535 507 -2367 541
rect -2277 507 -2109 541
rect -2019 507 -1851 541
rect -1761 507 -1593 541
rect -1503 507 -1335 541
rect -1245 507 -1077 541
rect -987 507 -819 541
rect -729 507 -561 541
rect -471 507 -303 541
rect -213 507 -45 541
rect 45 507 213 541
rect 303 507 471 541
rect 561 507 729 541
rect 819 507 987 541
rect 1077 507 1245 541
rect 1335 507 1503 541
rect 1593 507 1761 541
rect 1851 507 2019 541
rect 2109 507 2277 541
rect 2367 507 2535 541
<< locali >>
rect -2711 609 -2615 643
rect 2615 609 2711 643
rect -2711 547 -2677 609
rect 2677 547 2711 609
rect -2551 507 -2535 541
rect -2367 507 -2351 541
rect -2293 507 -2277 541
rect -2109 507 -2093 541
rect -2035 507 -2019 541
rect -1851 507 -1835 541
rect -1777 507 -1761 541
rect -1593 507 -1577 541
rect -1519 507 -1503 541
rect -1335 507 -1319 541
rect -1261 507 -1245 541
rect -1077 507 -1061 541
rect -1003 507 -987 541
rect -819 507 -803 541
rect -745 507 -729 541
rect -561 507 -545 541
rect -487 507 -471 541
rect -303 507 -287 541
rect -229 507 -213 541
rect -45 507 -29 541
rect 29 507 45 541
rect 213 507 229 541
rect 287 507 303 541
rect 471 507 487 541
rect 545 507 561 541
rect 729 507 745 541
rect 803 507 819 541
rect 987 507 1003 541
rect 1061 507 1077 541
rect 1245 507 1261 541
rect 1319 507 1335 541
rect 1503 507 1519 541
rect 1577 507 1593 541
rect 1761 507 1777 541
rect 1835 507 1851 541
rect 2019 507 2035 541
rect 2093 507 2109 541
rect 2277 507 2293 541
rect 2351 507 2367 541
rect 2535 507 2551 541
rect -2597 457 -2563 473
rect -2597 -535 -2563 -519
rect -2339 457 -2305 473
rect -2339 -535 -2305 -519
rect -2081 457 -2047 473
rect -2081 -535 -2047 -519
rect -1823 457 -1789 473
rect -1823 -535 -1789 -519
rect -1565 457 -1531 473
rect -1565 -535 -1531 -519
rect -1307 457 -1273 473
rect -1307 -535 -1273 -519
rect -1049 457 -1015 473
rect -1049 -535 -1015 -519
rect -791 457 -757 473
rect -791 -535 -757 -519
rect -533 457 -499 473
rect -533 -535 -499 -519
rect -275 457 -241 473
rect -275 -535 -241 -519
rect -17 457 17 473
rect -17 -535 17 -519
rect 241 457 275 473
rect 241 -535 275 -519
rect 499 457 533 473
rect 499 -535 533 -519
rect 757 457 791 473
rect 757 -535 791 -519
rect 1015 457 1049 473
rect 1015 -535 1049 -519
rect 1273 457 1307 473
rect 1273 -535 1307 -519
rect 1531 457 1565 473
rect 1531 -535 1565 -519
rect 1789 457 1823 473
rect 1789 -535 1823 -519
rect 2047 457 2081 473
rect 2047 -535 2081 -519
rect 2305 457 2339 473
rect 2305 -535 2339 -519
rect 2563 457 2597 473
rect 2563 -535 2597 -519
rect -2711 -643 -2677 -547
rect 2677 -643 2711 -547
<< viali >>
rect -2493 507 -2409 541
rect -2235 507 -2151 541
rect -1977 507 -1893 541
rect -1719 507 -1635 541
rect -1461 507 -1377 541
rect -1203 507 -1119 541
rect -945 507 -861 541
rect -687 507 -603 541
rect -429 507 -345 541
rect -171 507 -87 541
rect 87 507 171 541
rect 345 507 429 541
rect 603 507 687 541
rect 861 507 945 541
rect 1119 507 1203 541
rect 1377 507 1461 541
rect 1635 507 1719 541
rect 1893 507 1977 541
rect 2151 507 2235 541
rect 2409 507 2493 541
rect -2711 -487 -2677 487
rect -2597 -519 -2563 457
rect -2339 -519 -2305 457
rect -2081 -519 -2047 457
rect -1823 -519 -1789 457
rect -1565 -519 -1531 457
rect -1307 -519 -1273 457
rect -1049 -519 -1015 457
rect -791 -519 -757 457
rect -533 -519 -499 457
rect -275 -519 -241 457
rect -17 -519 17 457
rect 241 -519 275 457
rect 499 -519 533 457
rect 757 -519 791 457
rect 1015 -519 1049 457
rect 1273 -519 1307 457
rect 1531 -519 1565 457
rect 1789 -519 1823 457
rect 2047 -519 2081 457
rect 2305 -519 2339 457
rect 2563 -519 2597 457
rect 2677 -487 2711 487
rect -2677 -643 -2615 -609
rect -2615 -643 2615 -609
rect 2615 -643 2677 -609
<< metal1 >>
rect -2505 541 -2397 547
rect -2505 507 -2493 541
rect -2409 507 -2397 541
rect -2505 501 -2397 507
rect -2247 541 -2139 547
rect -2247 507 -2235 541
rect -2151 507 -2139 541
rect -2247 501 -2139 507
rect -1989 541 -1881 547
rect -1989 507 -1977 541
rect -1893 507 -1881 541
rect -1989 501 -1881 507
rect -1731 541 -1623 547
rect -1731 507 -1719 541
rect -1635 507 -1623 541
rect -1731 501 -1623 507
rect -1473 541 -1365 547
rect -1473 507 -1461 541
rect -1377 507 -1365 541
rect -1473 501 -1365 507
rect -1215 541 -1107 547
rect -1215 507 -1203 541
rect -1119 507 -1107 541
rect -1215 501 -1107 507
rect -957 541 -849 547
rect -957 507 -945 541
rect -861 507 -849 541
rect -957 501 -849 507
rect -699 541 -591 547
rect -699 507 -687 541
rect -603 507 -591 541
rect -699 501 -591 507
rect -441 541 -333 547
rect -441 507 -429 541
rect -345 507 -333 541
rect -441 501 -333 507
rect -183 541 -75 547
rect -183 507 -171 541
rect -87 507 -75 541
rect -183 501 -75 507
rect 75 541 183 547
rect 75 507 87 541
rect 171 507 183 541
rect 75 501 183 507
rect 333 541 441 547
rect 333 507 345 541
rect 429 507 441 541
rect 333 501 441 507
rect 591 541 699 547
rect 591 507 603 541
rect 687 507 699 541
rect 591 501 699 507
rect 849 541 957 547
rect 849 507 861 541
rect 945 507 957 541
rect 849 501 957 507
rect 1107 541 1215 547
rect 1107 507 1119 541
rect 1203 507 1215 541
rect 1107 501 1215 507
rect 1365 541 1473 547
rect 1365 507 1377 541
rect 1461 507 1473 541
rect 1365 501 1473 507
rect 1623 541 1731 547
rect 1623 507 1635 541
rect 1719 507 1731 541
rect 1623 501 1731 507
rect 1881 541 1989 547
rect 1881 507 1893 541
rect 1977 507 1989 541
rect 1881 501 1989 507
rect 2139 541 2247 547
rect 2139 507 2151 541
rect 2235 507 2247 541
rect 2139 501 2247 507
rect 2397 541 2505 547
rect 2397 507 2409 541
rect 2493 507 2505 541
rect 2397 501 2505 507
rect -2717 487 -2671 499
rect -2717 -487 -2711 487
rect -2677 -487 -2671 487
rect 2671 487 2717 499
rect -2717 -499 -2671 -487
rect -2603 457 -2557 469
rect -2603 -519 -2597 457
rect -2563 -519 -2557 457
rect -2603 -531 -2557 -519
rect -2345 457 -2299 469
rect -2345 -519 -2339 457
rect -2305 -519 -2299 457
rect -2345 -531 -2299 -519
rect -2087 457 -2041 469
rect -2087 -519 -2081 457
rect -2047 -519 -2041 457
rect -2087 -531 -2041 -519
rect -1829 457 -1783 469
rect -1829 -519 -1823 457
rect -1789 -519 -1783 457
rect -1829 -531 -1783 -519
rect -1571 457 -1525 469
rect -1571 -519 -1565 457
rect -1531 -519 -1525 457
rect -1571 -531 -1525 -519
rect -1313 457 -1267 469
rect -1313 -519 -1307 457
rect -1273 -519 -1267 457
rect -1313 -531 -1267 -519
rect -1055 457 -1009 469
rect -1055 -519 -1049 457
rect -1015 -519 -1009 457
rect -1055 -531 -1009 -519
rect -797 457 -751 469
rect -797 -519 -791 457
rect -757 -519 -751 457
rect -797 -531 -751 -519
rect -539 457 -493 469
rect -539 -519 -533 457
rect -499 -519 -493 457
rect -539 -531 -493 -519
rect -281 457 -235 469
rect -281 -519 -275 457
rect -241 -519 -235 457
rect -281 -531 -235 -519
rect -23 457 23 469
rect -23 -519 -17 457
rect 17 -519 23 457
rect -23 -531 23 -519
rect 235 457 281 469
rect 235 -519 241 457
rect 275 -519 281 457
rect 235 -531 281 -519
rect 493 457 539 469
rect 493 -519 499 457
rect 533 -519 539 457
rect 493 -531 539 -519
rect 751 457 797 469
rect 751 -519 757 457
rect 791 -519 797 457
rect 751 -531 797 -519
rect 1009 457 1055 469
rect 1009 -519 1015 457
rect 1049 -519 1055 457
rect 1009 -531 1055 -519
rect 1267 457 1313 469
rect 1267 -519 1273 457
rect 1307 -519 1313 457
rect 1267 -531 1313 -519
rect 1525 457 1571 469
rect 1525 -519 1531 457
rect 1565 -519 1571 457
rect 1525 -531 1571 -519
rect 1783 457 1829 469
rect 1783 -519 1789 457
rect 1823 -519 1829 457
rect 1783 -531 1829 -519
rect 2041 457 2087 469
rect 2041 -519 2047 457
rect 2081 -519 2087 457
rect 2041 -531 2087 -519
rect 2299 457 2345 469
rect 2299 -519 2305 457
rect 2339 -519 2345 457
rect 2299 -531 2345 -519
rect 2557 457 2603 469
rect 2557 -519 2563 457
rect 2597 -519 2603 457
rect 2671 -487 2677 487
rect 2711 -487 2717 487
rect 2671 -499 2717 -487
rect 2557 -531 2603 -519
rect -2689 -609 2689 -603
rect -2689 -643 -2677 -609
rect 2677 -643 2689 -609
rect -2689 -649 2689 -643
<< properties >>
string gencell sky130_fd_pr__nfet_01v8_lvt
string FIXED_BBOX -2694 -626 2694 626
string parameters w 5 l 1 m 1 nf 20 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 0 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__nfet_01v8 sky130_fd_pr__nfet_01v8_lvt  sky130_fd_bs_flash__special_sonosfet_star  sky130_fd_pr__nfet_g5v0d10v5 sky130_fd_pr__nfet_05v0_nvt  sky130_fd_pr__nfet_03v3_nvt} full_metal 1 viasrc 100 viadrn 100 viagate 50 viagb 100 viagr 80 viagl 80 viagt 0
string library sky130
<< end >>
