** sch_path:
*+ /home/users/xingyuni/ee372/bandgapReferenceCircuit/schematics/tsmc_bandgap_real_tempsweep.sch
**.subckt tsmc_bandgap_real_tempsweep
V1 VDD GND 'VDD' pwl 0us 0 5us 'VDD'
XQ2 GND GND Veb GND sky130_fd_pr__pnp_05v5_W3p40L3p40 nf=1 mult=1
Vr4 Vb net2 0
.save  i(vr4)
Vr2 Vb net1 0
.save  i(vr2)
Vm1 net5 Va 0
.save  i(vm1)
Vm2 net4 Vb 0
.save  i(vm2)
Vm3 net6 vbg 0
.save  i(vm3)
Vr1 Va net3 0
.save  i(vr1)
Vq2 Va Veb 0
.save  i(vq2)
XQ1 GND GND vbneg GND sky130_fd_pr__pnp_05v5_W3p40L3p40 m=39 nf=1 mult=1
XM5 vgate Va Vq GND sky130_fd_pr__nfet_01v8_lvt L='2' W='1' nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=26.95 m=26.95
XM6 Vq Vx GND GND sky130_fd_pr__nfet_01v8_lvt L=2 W=1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=3.65 m=3.65
XM9 vg Vb Vq GND sky130_fd_pr__nfet_01v8_lvt L='2' W='1' nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=26.95 m=26.95
XM7 Vx Vx GND GND sky130_fd_pr__nfet_01v8_lvt L=2 W=1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=3.65 m=3.65
XM13 Vx vgate VDD VDD sky130_fd_pr__pfet_01v8_lvt L=2 W=1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=77.32 m=77.32
XM1 net5 vgate VDD VDD sky130_fd_pr__pfet_01v8_lvt L=2 W=1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=386.6 m=386.6
XM2 net4 vgate VDD VDD sky130_fd_pr__pfet_01v8_lvt L=2 W=1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=386.6 m=386.6
XM3 net6 vgate VDD VDD sky130_fd_pr__pfet_01v8_lvt L=2 W=1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=386.6 m=386.6
XR1 GND net3 GND sky130_fd_pr__res_xhigh_po_0p35 L=21.839 mult=1 m=1
XR2 GND net2 GND sky130_fd_pr__res_xhigh_po_0p35 L=21.839 mult=1 m=1
XR3 vbneg net1 GND sky130_fd_pr__res_xhigh_po_0p35 L=3.763 mult=1 m=1
XR4 GND vbg GND sky130_fd_pr__res_xhigh_po_0p35 L=17.38 mult=1 m=1
XM4 vg vg VDD VDD sky130_fd_pr__pfet_01v8_lvt L=2 W=1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=38.66 m=38.66
XM8 vgate vg VDD VDD sky130_fd_pr__pfet_01v8_lvt L=2 W=1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=38.66 m=38.66
XM10 vgate porst GND GND sky130_fd_pr__nfet_01v8_lvt L='2' W='1' nf=1 ad='int((nf+1)/2) * W/nf * 0.29'
+ as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)'
+ nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=34 m=34
V2 porst GND 0 pulse(0V 1.8V 10us 0us 0us 5us)
C1 VDD vgate 20p m=1
C2 Va GND 20p m=1
**** begin user architecture code

.include /home/users/xingyuni/ee372/skywater-pdk/libraries/sky130_fd_pr_ngspice/latest/cells/nfet_01v8/sky130_fd_pr__nfet_01v8__tt.corner.spice
.include /home/users/xingyuni/ee372/skywater-pdk/libraries/sky130_fd_pr_ngspice/latest/cells/nfet_01v8_lvt/sky130_fd_pr__nfet_01v8_lvt__tt.corner.spice
.include /home/users/xingyuni/ee372/skywater-pdk/libraries/sky130_fd_pr_ngspice/latest/cells/pfet_01v8/sky130_fd_pr__pfet_01v8__tt.corner.spice
.include /home/users/xingyuni/ee372/skywater-pdk/libraries/sky130_fd_pr_ngspice/latest/cells/nfet_03v3_nvt/sky130_fd_pr__nfet_03v3_nvt__tt.corner.spice
.include /home/users/xingyuni/ee372/skywater-pdk/libraries/sky130_fd_pr_ngspice/latest/cells/nfet_05v0_nvt/sky130_fd_pr__nfet_05v0_nvt__tt.corner.spice
.include /home/users/xingyuni/ee372/skywater-pdk/libraries/sky130_fd_pr_ngspice/latest/cells/esd_nfet_01v8/sky130_fd_pr__esd_nfet_01v8__tt.corner.spice
.include /home/users/xingyuni/ee372/skywater-pdk/libraries/sky130_fd_pr_ngspice/latest/cells/pfet_01v8_lvt/sky130_fd_pr__pfet_01v8_lvt__tt.corner.spice
.include /home/users/xingyuni/ee372/skywater-pdk/libraries/sky130_fd_pr_ngspice/latest/cells/pfet_01v8_hvt/sky130_fd_pr__pfet_01v8_hvt__tt.corner.spice
.include /home/users/xingyuni/ee372/skywater-pdk/libraries/sky130_fd_pr_ngspice/latest/cells/esd_pfet_g5v0d10v5/sky130_fd_pr__esd_pfet_g5v0d10v5__tt.corner.spice
.include /home/users/xingyuni/ee372/skywater-pdk/libraries/sky130_fd_pr_ngspice/latest/cells/pfet_g5v0d10v5/sky130_fd_pr__pfet_g5v0d10v5__tt.corner.spice
.include /home/users/xingyuni/ee372/skywater-pdk/libraries/sky130_fd_pr_ngspice/latest/cells/pfet_g5v0d16v0/sky130_fd_pr__pfet_g5v0d16v0__tt.corner.spice
.include /home/users/xingyuni/ee372/skywater-pdk/libraries/sky130_fd_pr_ngspice/latest/cells/nfet_g5v0d10v5/sky130_fd_pr__nfet_g5v0d10v5__tt.corner.spice
.include /home/users/xingyuni/ee372/skywater-pdk/libraries/sky130_fd_pr_ngspice/latest/cells/nfet_g5v0d16v0/sky130_fd_pr__nfet_g5v0d16v0__tt_discrete.corner.spice
.include /home/users/xingyuni/ee372/skywater-pdk/libraries/sky130_fd_pr_ngspice/latest/cells/esd_nfet_g5v0d10v5/sky130_fd_pr__esd_nfet_g5v0d10v5__tt.corner.spice
.include /home/users/xingyuni/ee372/skywater-pdk/libraries/sky130_fd_pr_ngspice/latest/models/corners/tt/nonfet.spice
* Mismatch parameters
.include /home/users/xingyuni/ee372/skywater-pdk/libraries/sky130_fd_pr_ngspice/latest/cells/nfet_01v8/sky130_fd_pr__nfet_01v8__mismatch.corner.spice
.include /home/users/xingyuni/ee372/skywater-pdk/libraries/sky130_fd_pr_ngspice/latest/cells/pfet_01v8/sky130_fd_pr__pfet_01v8__mismatch.corner.spice
.include /home/users/xingyuni/ee372/skywater-pdk/libraries/sky130_fd_pr_ngspice/latest/cells/nfet_01v8_lvt/sky130_fd_pr__nfet_01v8_lvt__mismatch.corner.spice
.include /home/users/xingyuni/ee372/skywater-pdk/libraries/sky130_fd_pr_ngspice/latest/cells/pfet_01v8_lvt/sky130_fd_pr__pfet_01v8_lvt__mismatch.corner.spice
.include /home/users/xingyuni/ee372/skywater-pdk/libraries/sky130_fd_pr_ngspice/latest/cells/pfet_01v8_hvt/sky130_fd_pr__pfet_01v8_hvt__mismatch.corner.spice
.include /home/users/xingyuni/ee372/skywater-pdk/libraries/sky130_fd_pr_ngspice/latest/cells/nfet_g5v0d10v5/sky130_fd_pr__nfet_g5v0d10v5__mismatch.corner.spice
.include /home/users/xingyuni/ee372/skywater-pdk/libraries/sky130_fd_pr_ngspice/latest/cells/pfet_g5v0d10v5/sky130_fd_pr__pfet_g5v0d10v5__mismatch.corner.spice
.include /home/users/xingyuni/ee372/skywater-pdk/libraries/sky130_fd_pr_ngspice/latest/cells/nfet_05v0_nvt/sky130_fd_pr__nfet_05v0_nvt__mismatch.corner.spice
.include /home/users/xingyuni/ee372/skywater-pdk/libraries/sky130_fd_pr_ngspice/latest/cells/nfet_03v3_nvt/sky130_fd_pr__nfet_03v3_nvt__mismatch.corner.spice
* Resistor/home/users/xingyuni/ee372/skywater-pdk/libraries/sky130_fd_pr_ngspice/latest/Capacitor
.include /home/users/xingyuni/ee372/skywater-pdk/libraries/sky130_fd_pr_ngspice/latest/models/r+c/res_typical__cap_typical.spice
.include /home/users/xingyuni/ee372/skywater-pdk/libraries/sky130_fd_pr_ngspice/latest/models/r+c/res_typical__cap_typical__lin.spice
* Special cells
.include /home/users/xingyuni/ee372/skywater-pdk/libraries/sky130_fd_pr_ngspice/latest/models/corners/tt/specialized_cells.spice
* All models
.include /home/users/xingyuni/ee372/skywater-pdk/libraries/sky130_fd_pr_ngspice/latest/models/all.spice
.include /home/users/xingyuni/ee372/skywater-pdk/libraries/sky130_fd_pr_ngspice/latest/cells/pnp_05v5/sky130_fd_pr__pnp_05v5_W3p40L3p40.model.spice
* Corner
.include /home/users/xingyuni/ee372/skywater-pdk/libraries/sky130_fd_pr_ngspice/latest/models/corners/tt/rf.spice



.option savecurrents
.option warn=1
.param VDD=1.8
.param R3val='22.187k'
.param alpha='1'
.param R2R3ratio='5.6555038*alpha'
.param R2val='R3val*R2R3ratio'
.param R4R2ratio=0.79694273
.param R4val='R2val*R4R2ratio'
.nodeset v(vgate)=1.3
.option temp=0
.dc temp -10 80 10m
.control
save all  @m.xm13.msky130_fd_pr__pfet_01v8_lvt[gm]  @m.xm3.msky130_fd_pr__pfet_01v8_lvt[gm]
+  @m.xm4.msky130_fd_pr__pfet_01v8_lvt[gm]  @m.xm5.msky130_fd_pr__nfet_01v8_lvt[gm]  @m.xm6.msky130_fd_pr__nfet_01v8_lvt[gm]
+  @m.xm7.msky130_fd_pr__nfet_01v8_lvt[gm]  @m.xm8.msky130_fd_pr__pfet_01v8_lvt[gm]  @m.xm9.msky130_fd_pr__nfet_01v8_lvt[gm]
run
*plot Vbg
*plot deriv(Vbg)
save vbg deriv(vbg)
let i = vm3#branch
let indx27 = 3700
let indx0 = 1000
let indx70 = 8000
*indx is the index of temperature sweep for 27degC
echo 'Vbg @ 27degC'
let vbg27c = vbg[indx27]
print vbg27c
echo 'dVbe/degC & ppm @ 27degC'
print deriv(vbg)[indx27] deriv(vbg)[indx27]/vbg27c
echo 'ppm real'
print (vbg[indx70]-vbg[indx0])/vbg[indx27]/(70-0)*1e6
*plot deriv(vbg)/vbg27c
*plot v(va, vb) vs i
*plot vm1#branch vm2#branch vm3#branch
save deriv(vbg)/vbg27c
let vsg = vdd - vgate
let vsd1 = vdd - va
let vsd2 = vdd - vb
let vsd3 = vdd - vbg
let vthp = @m.xm1.msky130_fd_pr__pfet_01v8_lvt['vth']
let vov = vsg - vthp
*plot vov vsd1 vsd2 vsd3
let deltav = vb - vbneg
let r4 =vbg/vm3#branch
let r1 =va/vr1#branch
let r2 =vb/vr4#branch
let r3 =deltav/vr2#branch
let vptat =(r2/r3*deltav)
let sum = veb+vptat
*plot veb vptat sum
*plot deriv(veb) deriv(vptat)
save veb vptat sum deriv(veb) deriv(vptat)
let gm1=@m.xm1.msky130_fd_pr__pfet_01v8_lvt[gm]
let gm2=@m.xm2.msky130_fd_pr__pfet_01v8_lvt[gm]
let Av2=gm2 * ((r3 + r3/ln(39)) * r2 / (r3 + r3/ln(39) + r2) )
let Av1=gm1 * (r1 * r3/ln(39))/(r1 + r3/ln(39))
*plot Av1 Av2 Av2/Av1
let gm13=@m.xm13.msky130_fd_pr__pfet_01v8_lvt[gm]
let gm3=@m.xm3.msky130_fd_pr__pfet_01v8_lvt[gm]
let gm4=@m.xm4.msky130_fd_pr__pfet_01v8_lvt[gm]
let gm5=@m.xm5.msky130_fd_pr__nfet_01v8_lvt[gm]
let gm6=@m.xm6.msky130_fd_pr__nfet_01v8_lvt[gm]
let gm7=@m.xm7.msky130_fd_pr__nfet_01v8_lvt[gm]
let gm8=@m.xm8.msky130_fd_pr__pfet_01v8_lvt[gm]
let gm9=@m.xm9.msky130_fd_pr__nfet_01v8_lvt[gm]
let vdsat1=2/(gm1/vm1#branch)
let vdsat2=2/(gm2/vm2#branch)
let vdsat3=2/(gm3/vm3#branch)
let vdsat4=2/(gm4/@m.xm4.msky130_fd_pr__pfet_01v8_lvt[id])
let vdsat5=2/(gm5/@m.xm5.msky130_fd_pr__nfet_01v8_lvt[id])
let vdsat6=2/(gm6/@m.xm6.msky130_fd_pr__nfet_01v8_lvt[id])
let vdsat7=2/(gm7/@m.xm7.msky130_fd_pr__nfet_01v8_lvt[id])
let vdsat8=2/(gm8/@m.xm8.msky130_fd_pr__pfet_01v8_lvt[id])
let vdsat9=2/(gm9/@m.xm9.msky130_fd_pr__nfet_01v8_lvt[id])
let vdsat13=2/(gm13/@m.xm13.msky130_fd_pr__pfet_01v8_lvt[id])
save (vdd-va-vdsat1) (vdd-vb-vdsat2) (vdd-vbg-vdsat3)  (vdd-vgate-vdsat4) (vgate-vq-vdsat5)
+ (vq-0-vdsat6)  (vx-0-vdsat7) (vdd-vg-vdsat8) (vg-vq-vdsat9) (vdd-vx-vdsat13)

write
unset askquit
quit
.endc


**** end user architecture code
**.ends
.GLOBAL VDD
.GLOBAL GND
.end
