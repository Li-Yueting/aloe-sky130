VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO sky130_asc_cap_mim_m3_1
  CLASS CORE ;
  FOREIGN sky130_asc_cap_mim_m3_1 ;
  ORIGIN 0.000 0.000 ;
  SIZE 36.855 BY 9.400 ;
  SITE unitasc ;
  PIN Cin
    DIRECTION INOUT ;
    PORT
      LAYER met4 ;
        RECT 3.450 5.310 3.930 8.190 ;
        RECT 7.045 5.310 7.525 8.190 ;
        RECT 10.640 5.310 11.120 8.190 ;
        RECT 14.235 5.310 14.715 8.190 ;
        RECT 17.830 5.310 18.310 8.190 ;
        RECT 21.425 5.310 21.905 8.190 ;
        RECT 25.020 5.310 25.500 8.190 ;
        RECT 28.615 5.310 29.095 8.190 ;
        RECT 32.210 5.310 32.690 8.190 ;
        RECT 35.805 5.310 36.285 8.190 ;
        RECT 3.450 1.810 3.930 4.690 ;
        RECT 7.045 1.810 7.525 4.690 ;
        RECT 10.640 1.810 11.120 4.690 ;
        RECT 14.235 1.810 14.715 4.690 ;
        RECT 17.830 1.810 18.310 4.690 ;
        RECT 21.425 1.810 21.905 4.690 ;
        RECT 25.020 1.810 25.500 4.690 ;
        RECT 28.615 1.810 29.095 4.690 ;
        RECT 32.210 1.810 32.690 4.690 ;
        RECT 35.805 1.810 36.285 4.690 ;
    END
  END Cin
  PIN Cout
    DIRECTION INOUT ;
    PORT
      LAYER met4 ;
        RECT 1.150 7.555 2.750 7.650 ;
        RECT 4.750 7.555 6.350 7.650 ;
        RECT 8.350 7.555 9.950 7.650 ;
        RECT 11.950 7.555 13.550 7.650 ;
        RECT 15.550 7.555 17.150 7.650 ;
        RECT 19.150 7.555 20.750 7.650 ;
        RECT 22.750 7.555 24.350 7.650 ;
        RECT 26.350 7.555 27.950 7.650 ;
        RECT 29.950 7.555 31.550 7.650 ;
        RECT 33.550 7.555 35.150 7.650 ;
        RECT 1.150 5.945 2.760 7.555 ;
        RECT 4.745 5.945 6.355 7.555 ;
        RECT 8.340 5.945 9.950 7.555 ;
        RECT 11.935 5.945 13.550 7.555 ;
        RECT 15.530 5.945 17.150 7.555 ;
        RECT 19.125 5.945 20.750 7.555 ;
        RECT 22.720 5.945 24.350 7.555 ;
        RECT 26.315 5.945 27.950 7.555 ;
        RECT 29.910 5.945 31.550 7.555 ;
        RECT 33.505 5.945 35.150 7.555 ;
        RECT 1.150 4.055 2.750 5.945 ;
        RECT 4.750 4.055 6.350 5.945 ;
        RECT 8.350 4.055 9.950 5.945 ;
        RECT 11.950 4.055 13.550 5.945 ;
        RECT 15.550 4.055 17.150 5.945 ;
        RECT 19.150 4.055 20.750 5.945 ;
        RECT 22.750 4.055 24.350 5.945 ;
        RECT 26.350 4.055 27.950 5.945 ;
        RECT 29.950 4.055 31.550 5.945 ;
        RECT 33.550 4.055 35.150 5.945 ;
        RECT 1.150 2.445 2.760 4.055 ;
        RECT 4.745 2.445 6.355 4.055 ;
        RECT 8.340 2.445 9.950 4.055 ;
        RECT 11.935 2.445 13.550 4.055 ;
        RECT 15.530 2.445 17.150 4.055 ;
        RECT 19.125 2.445 20.750 4.055 ;
        RECT 22.720 2.445 24.350 4.055 ;
        RECT 26.315 2.445 27.950 4.055 ;
        RECT 29.910 2.445 31.550 4.055 ;
        RECT 33.505 2.445 35.150 4.055 ;
        RECT 1.150 1.450 2.750 2.445 ;
        RECT 4.750 1.450 6.350 2.445 ;
        RECT 8.350 1.450 9.950 2.445 ;
        RECT 11.950 1.450 13.550 2.445 ;
        RECT 15.550 1.450 17.150 2.445 ;
        RECT 19.150 1.450 20.750 2.445 ;
        RECT 22.750 1.450 24.350 2.445 ;
        RECT 26.350 1.450 27.950 2.445 ;
        RECT 29.950 1.450 31.550 2.445 ;
        RECT 33.550 1.450 35.150 2.445 ;
        RECT 0.460 0.750 36.300 1.450 ;
    END
  END Cout
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.460 9.100 36.300 9.700 ;
    END
  END VPWR
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.460 -0.300 36.300 0.300 ;
    END
  END VGND
  OBS
      LAYER li1 ;
        RECT 0.460 9.250 36.300 9.550 ;
        RECT 0.460 -0.150 36.300 0.150 ;
      LAYER mcon ;
        RECT 1.310 9.250 1.610 9.550 ;
        RECT 3.310 9.250 3.610 9.550 ;
        RECT 5.310 9.250 5.610 9.550 ;
        RECT 7.310 9.250 7.610 9.550 ;
        RECT 9.310 9.250 9.610 9.550 ;
        RECT 11.310 9.250 11.610 9.550 ;
        RECT 13.310 9.250 13.610 9.550 ;
        RECT 15.310 9.250 15.610 9.550 ;
        RECT 17.310 9.250 17.610 9.550 ;
        RECT 19.310 9.250 19.610 9.550 ;
        RECT 21.310 9.250 21.610 9.550 ;
        RECT 23.310 9.250 23.610 9.550 ;
        RECT 25.310 9.250 25.610 9.550 ;
        RECT 27.310 9.250 27.610 9.550 ;
        RECT 29.310 9.250 29.610 9.550 ;
        RECT 31.310 9.250 31.610 9.550 ;
        RECT 33.310 9.250 33.610 9.550 ;
        RECT 35.310 9.250 35.610 9.550 ;
        RECT 1.310 -0.150 1.610 0.150 ;
        RECT 3.310 -0.150 3.610 0.150 ;
        RECT 5.310 -0.150 5.610 0.150 ;
        RECT 7.310 -0.150 7.610 0.150 ;
        RECT 9.310 -0.150 9.610 0.150 ;
        RECT 11.310 -0.150 11.610 0.150 ;
        RECT 13.310 -0.150 13.610 0.150 ;
        RECT 15.310 -0.150 15.610 0.150 ;
        RECT 17.310 -0.150 17.610 0.150 ;
        RECT 19.310 -0.150 19.610 0.150 ;
        RECT 21.310 -0.150 21.610 0.150 ;
        RECT 23.310 -0.150 23.610 0.150 ;
        RECT 25.310 -0.150 25.610 0.150 ;
        RECT 27.310 -0.150 27.610 0.150 ;
        RECT 29.310 -0.150 29.610 0.150 ;
        RECT 31.310 -0.150 31.610 0.150 ;
        RECT 33.310 -0.150 33.610 0.150 ;
        RECT 35.310 -0.150 35.610 0.150 ;
      LAYER met2 ;
        RECT 0.450 7.850 1.450 8.250 ;
        RECT 0.560 0.800 1.360 1.300 ;
      LAYER via2 ;
        RECT 0.550 7.900 1.350 8.200 ;
        RECT 0.660 0.850 1.260 1.250 ;
      LAYER met3 ;
        RECT 0.450 1.750 36.310 8.250 ;
        RECT 0.460 0.750 1.460 1.350 ;
      LAYER via3 ;
        RECT 3.530 5.390 3.850 8.110 ;
        RECT 7.125 5.390 7.445 8.110 ;
        RECT 10.720 5.390 11.040 8.110 ;
        RECT 14.315 5.390 14.635 8.110 ;
        RECT 17.910 5.390 18.230 8.110 ;
        RECT 21.505 5.390 21.825 8.110 ;
        RECT 25.100 5.390 25.420 8.110 ;
        RECT 28.695 5.390 29.015 8.110 ;
        RECT 32.290 5.390 32.610 8.110 ;
        RECT 35.885 5.390 36.205 8.110 ;
        RECT 3.530 1.890 3.850 4.610 ;
        RECT 7.125 1.890 7.445 4.610 ;
        RECT 10.720 1.890 11.040 4.610 ;
        RECT 14.315 1.890 14.635 4.610 ;
        RECT 17.910 1.890 18.230 4.610 ;
        RECT 21.505 1.890 21.825 4.610 ;
        RECT 25.100 1.890 25.420 4.610 ;
        RECT 28.695 1.890 29.015 4.610 ;
        RECT 32.290 1.890 32.610 4.610 ;
        RECT 35.885 1.890 36.205 4.610 ;
        RECT 0.560 0.800 1.360 1.300 ;
  END
END sky130_asc_cap_mim_m3_1
END LIBRARY

