* NGSPICE file created from bgr_top.ext - technology: sky130A

.subckt sky130_asc_res_xhigh_po_2p85_1 Rin Rout VPWR VGND a_2148_115#
X0 Rin a_2148_115# VGND sky130_fd_pr__res_xhigh_po w=2.85e+06u l=7.88e+06u
X1 Rout a_2148_115# VGND sky130_fd_pr__res_xhigh_po w=2.85e+06u l=7.88e+06u
C0 a_2148_115# VPWR 0.17fF
C1 Rin VPWR 0.17fF
C2 Rin Rout 0.12fF
C3 VPWR VGND 2.31fF
C4 Rout VGND 1.26fF
C5 Rin VGND 0.78fF
C6 a_2148_115# VGND 2.70fF
.ends

.subckt sky130_asc_pfet_01v8_lvt_60 GATE SOURCE DRAIN VGND VPWR VSUBS
X0 DRAIN GATE SOURCE VPWR sky130_fd_pr__pfet_01v8_lvt ad=5.79855e+13p pd=4.1788e+08u as=5.6115e+13p ps=4.044e+08u w=6.45e+06u l=2e+06u
X1 SOURCE GATE DRAIN VPWR sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=6.45e+06u l=2e+06u
X2 DRAIN GATE SOURCE VPWR sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=6.45e+06u l=2e+06u
X3 SOURCE GATE DRAIN VPWR sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=6.45e+06u l=2e+06u
X4 DRAIN GATE SOURCE VPWR sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=6.45e+06u l=2e+06u
X5 DRAIN GATE SOURCE VPWR sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=6.45e+06u l=2e+06u
X6 DRAIN GATE SOURCE VPWR sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=6.45e+06u l=2e+06u
X7 DRAIN GATE SOURCE VPWR sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=6.45e+06u l=2e+06u
X8 DRAIN GATE SOURCE VPWR sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=6.45e+06u l=2e+06u
X9 SOURCE GATE DRAIN VPWR sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=6.45e+06u l=2e+06u
X10 DRAIN GATE SOURCE VPWR sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=6.45e+06u l=2e+06u
X11 SOURCE GATE DRAIN VPWR sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=6.45e+06u l=2e+06u
X12 SOURCE GATE DRAIN VPWR sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=6.45e+06u l=2e+06u
X13 DRAIN GATE SOURCE VPWR sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=6.45e+06u l=2e+06u
X14 DRAIN GATE SOURCE VPWR sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=6.45e+06u l=2e+06u
X15 SOURCE GATE DRAIN VPWR sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=6.45e+06u l=2e+06u
X16 SOURCE GATE DRAIN VPWR sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=6.45e+06u l=2e+06u
X17 DRAIN GATE SOURCE VPWR sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=6.45e+06u l=2e+06u
X18 SOURCE GATE DRAIN VPWR sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=6.45e+06u l=2e+06u
X19 DRAIN GATE SOURCE VPWR sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=6.45e+06u l=2e+06u
X20 SOURCE GATE DRAIN VPWR sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=6.45e+06u l=2e+06u
X21 DRAIN GATE SOURCE VPWR sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=6.45e+06u l=2e+06u
X22 SOURCE GATE DRAIN VPWR sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=6.45e+06u l=2e+06u
X23 DRAIN GATE SOURCE VPWR sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=6.45e+06u l=2e+06u
X24 SOURCE GATE DRAIN VPWR sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=6.45e+06u l=2e+06u
X25 DRAIN GATE SOURCE VPWR sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=6.45e+06u l=2e+06u
X26 SOURCE GATE DRAIN VPWR sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=6.45e+06u l=2e+06u
X27 SOURCE GATE DRAIN VPWR sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=6.45e+06u l=2e+06u
X28 DRAIN GATE SOURCE VPWR sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=6.45e+06u l=2e+06u
X29 SOURCE GATE DRAIN VPWR sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=6.45e+06u l=2e+06u
X30 DRAIN GATE SOURCE VPWR sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=6.45e+06u l=2e+06u
X31 SOURCE GATE DRAIN VPWR sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=6.45e+06u l=2e+06u
X32 DRAIN GATE SOURCE VPWR sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=6.45e+06u l=2e+06u
X33 SOURCE GATE DRAIN VPWR sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=6.45e+06u l=2e+06u
X34 DRAIN GATE SOURCE VPWR sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=6.45e+06u l=2e+06u
X35 SOURCE GATE DRAIN VPWR sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=6.45e+06u l=2e+06u
X36 DRAIN GATE SOURCE VPWR sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=6.45e+06u l=2e+06u
X37 SOURCE GATE DRAIN VPWR sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=6.45e+06u l=2e+06u
X38 DRAIN GATE SOURCE VPWR sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=6.45e+06u l=2e+06u
X39 SOURCE GATE DRAIN VPWR sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=6.45e+06u l=2e+06u
X40 SOURCE GATE DRAIN VPWR sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=6.45e+06u l=2e+06u
X41 DRAIN GATE SOURCE VPWR sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=6.45e+06u l=2e+06u
X42 DRAIN GATE SOURCE VPWR sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=6.45e+06u l=2e+06u
X43 DRAIN GATE SOURCE VPWR sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=6.45e+06u l=2e+06u
X44 SOURCE GATE DRAIN VPWR sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=6.45e+06u l=2e+06u
X45 SOURCE GATE DRAIN VPWR sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=6.45e+06u l=2e+06u
X46 DRAIN GATE SOURCE VPWR sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=6.45e+06u l=2e+06u
X47 SOURCE GATE DRAIN VPWR sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=6.45e+06u l=2e+06u
X48 SOURCE GATE DRAIN VPWR sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=6.45e+06u l=2e+06u
X49 SOURCE GATE DRAIN VPWR sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=6.45e+06u l=2e+06u
X50 DRAIN GATE SOURCE VPWR sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=6.45e+06u l=2e+06u
X51 SOURCE GATE DRAIN VPWR sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=6.45e+06u l=2e+06u
X52 SOURCE GATE DRAIN VPWR sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=6.45e+06u l=2e+06u
X53 SOURCE GATE DRAIN VPWR sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=6.45e+06u l=2e+06u
X54 DRAIN GATE SOURCE VPWR sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=6.45e+06u l=2e+06u
X55 SOURCE GATE DRAIN VPWR sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=6.45e+06u l=2e+06u
X56 DRAIN GATE SOURCE VPWR sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=6.45e+06u l=2e+06u
X57 DRAIN GATE SOURCE VPWR sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=6.45e+06u l=2e+06u
X58 SOURCE GATE DRAIN VPWR sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=6.45e+06u l=2e+06u
X59 DRAIN GATE SOURCE VPWR sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=6.45e+06u l=2e+06u
C0 VGND DRAIN 5.28fF
C1 VGND GATE 12.31fF
C2 SOURCE DRAIN 1.25fF
C3 SOURCE VPWR 22.83fF
C4 SOURCE GATE 0.18fF
C5 VGND SOURCE 0.32fF
C6 DRAIN VPWR 1.83fF
C7 DRAIN GATE 25.46fF
C8 GATE VPWR 27.32fF
C9 VGND VSUBS 25.41fF
C10 SOURCE VSUBS 0.00fF
C11 DRAIN VSUBS 9.62fF
C12 GATE VSUBS 30.27fF
C13 VPWR VSUBS 142.65fF
.ends

.subckt sky130_asc_pnp_05v5_W3p40L3p40_7 Emitter Base Collector VPWR VGND
X0 Collector Base Emitter sky130_fd_pr__pnp_05v5 area=0p
X1 Collector Base Emitter sky130_fd_pr__pnp_05v5 area=0p
X2 Collector Base Emitter sky130_fd_pr__pnp_05v5 area=0p
X3 Collector Base Emitter sky130_fd_pr__pnp_05v5 area=0p
X4 Collector Base Emitter sky130_fd_pr__pnp_05v5 area=0p
X5 Collector Base Emitter sky130_fd_pr__pnp_05v5 area=0p
X6 Collector Base Emitter sky130_fd_pr__pnp_05v5 area=0p
C0 Base Emitter 18.67fF
C1 VGND Collector 9.81fF
C2 VPWR Collector 11.49fF
C3 Emitter Collector 9.06fF
C4 Base Collector 28.86fF
.ends

.subckt sky130_asc_res_xhigh_po_2p85_2 Rin Rout VPWR a_2723_115# VGND
X0 Rout a_2723_115# VGND sky130_fd_pr__res_xhigh_po w=2.85e+06u l=1.075e+07u
X1 Rin a_2723_115# VGND sky130_fd_pr__res_xhigh_po w=2.85e+06u l=1.075e+07u
C0 Rin VPWR 0.17fF
C1 Rout Rin 0.12fF
C2 a_2723_115# VPWR 0.17fF
C3 VPWR VGND 2.83fF
C4 Rout VGND 1.26fF
C5 Rin VGND 0.78fF
C6 a_2723_115# VGND 2.70fF
.ends

.subckt sky130_asc_pfet_01v8_lvt_12 GATE SOURCE DRAIN VGND VPWR VSUBS
X0 SOURCE GATE DRAIN VPWR sky130_fd_pr__pfet_01v8_lvt ad=1.1223e+13p pd=8.088e+07u as=1.30935e+13p ps=9.436e+07u w=6.45e+06u l=2e+06u
X1 DRAIN GATE SOURCE VPWR sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=6.45e+06u l=2e+06u
X2 DRAIN GATE SOURCE VPWR sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=6.45e+06u l=2e+06u
X3 SOURCE GATE DRAIN VPWR sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=6.45e+06u l=2e+06u
X4 SOURCE GATE DRAIN VPWR sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=6.45e+06u l=2e+06u
X5 DRAIN GATE SOURCE VPWR sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=6.45e+06u l=2e+06u
X6 SOURCE GATE DRAIN VPWR sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=6.45e+06u l=2e+06u
X7 DRAIN GATE SOURCE VPWR sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=6.45e+06u l=2e+06u
X8 DRAIN GATE SOURCE VPWR sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=6.45e+06u l=2e+06u
X9 SOURCE GATE DRAIN VPWR sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=6.45e+06u l=2e+06u
X10 SOURCE GATE DRAIN VPWR sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=6.45e+06u l=2e+06u
X11 DRAIN GATE SOURCE VPWR sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=6.45e+06u l=2e+06u
C0 SOURCE VGND 0.06fF
C1 VGND DRAIN 1.08fF
C2 VGND GATE 2.51fF
C3 SOURCE DRAIN 0.26fF
C4 SOURCE GATE 0.04fF
C5 SOURCE VPWR 4.54fF
C6 GATE DRAIN 5.17fF
C7 VPWR DRAIN 0.42fF
C8 VPWR GATE 5.46fF
C9 VGND VSUBS 5.31fF
C10 SOURCE VSUBS 0.00fF
C11 DRAIN VSUBS 1.99fF
C12 GATE VSUBS 6.20fF
C13 VPWR VSUBS 29.52fF
.ends

.subckt sky130_asc_nfet_01v8_lvt_9 GATE SOURCE DRAIN VPWR VGND
X0 SOURCE GATE DRAIN VGND sky130_fd_pr__nfet_01v8_lvt ad=5.8e+12p pd=4.29e+07u as=5.8e+12p ps=4.29e+07u w=4e+06u l=2e+06u
X1 SOURCE GATE DRAIN VGND sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=2e+06u
X2 DRAIN GATE SOURCE VGND sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=2e+06u
X3 SOURCE GATE DRAIN VGND sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=2e+06u
X4 DRAIN GATE SOURCE VGND sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=2e+06u
X5 SOURCE GATE DRAIN VGND sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=2e+06u
X6 DRAIN GATE SOURCE VGND sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=2e+06u
X7 SOURCE GATE DRAIN VGND sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=2e+06u
X8 DRAIN GATE SOURCE VGND sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=2e+06u
C0 SOURCE DRAIN 0.05fF
C1 SOURCE GATE 0.01fF
C2 DRAIN GATE 1.66fF
C3 SOURCE VPWR 1.38fF
C4 VPWR VGND 3.99fF
C5 SOURCE VGND 2.64fF
C6 DRAIN VGND 2.28fF
C7 GATE VGND 11.48fF
.ends

.subckt sky130_asc_pfet_01v8_lvt_6 GATE SOURCE DRAIN VGND VPWR VSUBS
X0 SOURCE GATE DRAIN VPWR sky130_fd_pr__pfet_01v8_lvt ad=5.6115e+12p pd=4.044e+07u as=7.482e+12p ps=5.392e+07u w=6.45e+06u l=2e+06u
X1 SOURCE GATE DRAIN VPWR sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=6.45e+06u l=2e+06u
X2 DRAIN GATE SOURCE VPWR sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=6.45e+06u l=2e+06u
X3 DRAIN GATE SOURCE VPWR sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=6.45e+06u l=2e+06u
X4 SOURCE GATE DRAIN VPWR sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=6.45e+06u l=2e+06u
X5 DRAIN GATE SOURCE VPWR sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=6.45e+06u l=2e+06u
C0 VPWR GATE 2.73fF
C1 DRAIN GATE 2.63fF
C2 SOURCE GATE 0.02fF
C3 VGND GATE 1.28fF
C4 DRAIN VPWR 0.24fF
C5 VPWR SOURCE 2.27fF
C6 DRAIN SOURCE 0.14fF
C7 DRAIN VGND 0.56fF
C8 VGND SOURCE 0.03fF
C9 VGND VSUBS 2.79fF
C10 SOURCE VSUBS 0.00fF
C11 DRAIN VSUBS 1.04fF
C12 GATE VSUBS 3.19fF
C13 VPWR VSUBS 15.38fF
.ends

.subckt sky130_asc_pnp_05v5_W3p40L3p40_1 Emitter Base Collector VPWR VGND
X0 Collector Base Emitter sky130_fd_pr__pnp_05v5 area=0p
C0 Emitter Base 1.55fF
C1 VGND Collector 1.50fF
C2 VPWR Collector 1.46fF
C3 Emitter Collector 0.40fF
C4 Base Collector 3.33fF
.ends

.subckt sky130_asc_cap_mim_m3_1 Cin Cout VPWR VGND VSUBS
X0 Cout Cin sky130_fd_pr__cap_mim_m3_1 l=2e+06u w=2e+06u
X1 Cout Cin sky130_fd_pr__cap_mim_m3_1 l=2e+06u w=2e+06u
X2 Cout Cin sky130_fd_pr__cap_mim_m3_1 l=2e+06u w=2e+06u
X3 Cout Cin sky130_fd_pr__cap_mim_m3_1 l=2e+06u w=2e+06u
X4 Cout Cin sky130_fd_pr__cap_mim_m3_1 l=2e+06u w=2e+06u
X5 Cout Cin sky130_fd_pr__cap_mim_m3_1 l=2e+06u w=2e+06u
X6 Cout Cin sky130_fd_pr__cap_mim_m3_1 l=2e+06u w=2e+06u
X7 Cout Cin sky130_fd_pr__cap_mim_m3_1 l=2e+06u w=2e+06u
X8 Cout Cin sky130_fd_pr__cap_mim_m3_1 l=2e+06u w=2e+06u
X9 Cout Cin sky130_fd_pr__cap_mim_m3_1 l=2e+06u w=2e+06u
X10 Cout Cin sky130_fd_pr__cap_mim_m3_1 l=2e+06u w=2e+06u
X11 Cout Cin sky130_fd_pr__cap_mim_m3_1 l=2e+06u w=2e+06u
X12 Cout Cin sky130_fd_pr__cap_mim_m3_1 l=2e+06u w=2e+06u
X13 Cout Cin sky130_fd_pr__cap_mim_m3_1 l=2e+06u w=2e+06u
X14 Cout Cin sky130_fd_pr__cap_mim_m3_1 l=2e+06u w=2e+06u
X15 Cout Cin sky130_fd_pr__cap_mim_m3_1 l=2e+06u w=2e+06u
X16 Cout Cin sky130_fd_pr__cap_mim_m3_1 l=2e+06u w=2e+06u
X17 Cout Cin sky130_fd_pr__cap_mim_m3_1 l=2e+06u w=2e+06u
X18 Cout Cin sky130_fd_pr__cap_mim_m3_1 l=2e+06u w=2e+06u
X19 Cout Cin sky130_fd_pr__cap_mim_m3_1 l=2e+06u w=2e+06u
C0 Cin Cout 28.31fF
C1 Cout VSUBS 2.81fF
C2 Cin VSUBS 6.38fF
C3 VGND VSUBS 6.63fF
C4 VPWR VSUBS 6.63fF
.ends

.subckt sky130_asc_pnp_05v5_W3p40L3p40_8 Emitter Base Collector VPWR VGND
X0 Collector Base Emitter sky130_fd_pr__pnp_05v5 area=0p
X1 Collector Base Emitter sky130_fd_pr__pnp_05v5 area=0p
X2 Collector Base Emitter sky130_fd_pr__pnp_05v5 area=0p
X3 Collector Base Emitter sky130_fd_pr__pnp_05v5 area=0p
X4 Collector Base Emitter sky130_fd_pr__pnp_05v5 area=0p
X5 Collector Base Emitter sky130_fd_pr__pnp_05v5 area=0p
X6 Collector Base Emitter sky130_fd_pr__pnp_05v5 area=0p
X7 Collector Base Emitter sky130_fd_pr__pnp_05v5 area=0p
C0 Emitter Base 21.50fF
C1 VGND Collector 11.20fF
C2 VPWR Collector 13.12fF
C3 Emitter Collector 10.49fF
C4 Base Collector 33.06fF
.ends

.subckt sky130_asc_nfet_01v8_lvt_1 GATE SOURCE DRAIN VPWR VGND
X0 SOURCE GATE DRAIN VGND sky130_fd_pr__nfet_01v8_lvt ad=1.16e+12p pd=8.58e+06u as=1.16e+12p ps=8.58e+06u w=4e+06u l=2e+06u
C0 GATE DRAIN 0.18fF
C1 VPWR SOURCE 0.17fF
C2 GATE SOURCE 0.00fF
C3 DRAIN SOURCE 0.01fF
C4 VPWR VGND 0.64fF
C5 SOURCE VGND 0.40fF
C6 DRAIN VGND 0.34fF
C7 GATE VGND 1.34fF
.ends

.subckt bgr_top porst va vb vbg VSS VDD
Xsky130_asc_res_xhigh_po_2p85_1_7 sky130_asc_res_xhigh_po_2p85_1_7/Rin sky130_asc_res_xhigh_po_2p85_1_6/Rin
+ VDD VSS sky130_asc_res_xhigh_po_2p85_1_7/a_2148_115# sky130_asc_res_xhigh_po_2p85_1
Xsky130_asc_res_xhigh_po_2p85_1_8 vbg sky130_asc_res_xhigh_po_2p85_1_7/Rin VDD VSS
+ sky130_asc_res_xhigh_po_2p85_1_8/a_2148_115# sky130_asc_res_xhigh_po_2p85_1
Xsky130_asc_res_xhigh_po_2p85_1_9 sky130_asc_res_xhigh_po_2p85_1_9/Rin sky130_asc_res_xhigh_po_2p85_2_0/Rin
+ VDD VSS sky130_asc_res_xhigh_po_2p85_1_9/a_2148_115# sky130_asc_res_xhigh_po_2p85_1
Xsky130_asc_pfet_01v8_lvt_60_0 sky130_asc_cap_mim_m3_1_4/Cout VDD vbg VSS VDD VSS
+ sky130_asc_pfet_01v8_lvt_60
Xsky130_asc_pfet_01v8_lvt_60_1 sky130_asc_cap_mim_m3_1_4/Cout VDD vb VSS VDD VSS sky130_asc_pfet_01v8_lvt_60
Xsky130_asc_pfet_01v8_lvt_60_2 sky130_asc_cap_mim_m3_1_4/Cout VDD va VSS VDD VSS sky130_asc_pfet_01v8_lvt_60
Xsky130_asc_res_xhigh_po_2p85_1_30 va sky130_asc_res_xhigh_po_2p85_1_29/Rin VDD VSS
+ sky130_asc_res_xhigh_po_2p85_1_30/a_2148_115# sky130_asc_res_xhigh_po_2p85_1
Xsky130_asc_res_xhigh_po_2p85_1_20 vb sky130_asc_res_xhigh_po_2p85_1_19/Rin VDD VSS
+ sky130_asc_res_xhigh_po_2p85_1_20/a_2148_115# sky130_asc_res_xhigh_po_2p85_1
Xsky130_asc_pnp_05v5_W3p40L3p40_7_0 sky130_asc_res_xhigh_po_2p85_1_19/Rout VSS VSS
+ VDD VSS sky130_asc_pnp_05v5_W3p40L3p40_7
Xsky130_asc_res_xhigh_po_2p85_1_21 sky130_asc_res_xhigh_po_2p85_1_21/Rin sky130_asc_res_xhigh_po_2p85_2_1/Rin
+ VDD VSS sky130_asc_res_xhigh_po_2p85_1_21/a_2148_115# sky130_asc_res_xhigh_po_2p85_1
Xsky130_asc_res_xhigh_po_2p85_1_10 sky130_asc_res_xhigh_po_2p85_1_10/Rin sky130_asc_res_xhigh_po_2p85_1_9/Rin
+ VDD VSS sky130_asc_res_xhigh_po_2p85_1_10/a_2148_115# sky130_asc_res_xhigh_po_2p85_1
Xsky130_asc_res_xhigh_po_2p85_2_0 sky130_asc_res_xhigh_po_2p85_2_0/Rin VSS VDD sky130_asc_res_xhigh_po_2p85_2_0/a_2723_115#
+ VSS sky130_asc_res_xhigh_po_2p85_2
Xsky130_asc_res_xhigh_po_2p85_1_22 sky130_asc_res_xhigh_po_2p85_1_22/Rin sky130_asc_res_xhigh_po_2p85_1_21/Rin
+ VDD VSS sky130_asc_res_xhigh_po_2p85_1_22/a_2148_115# sky130_asc_res_xhigh_po_2p85_1
Xsky130_asc_res_xhigh_po_2p85_1_11 sky130_asc_res_xhigh_po_2p85_1_11/Rin sky130_asc_res_xhigh_po_2p85_1_10/Rin
+ VDD VSS sky130_asc_res_xhigh_po_2p85_1_11/a_2148_115# sky130_asc_res_xhigh_po_2p85_1
Xsky130_asc_res_xhigh_po_2p85_2_1 sky130_asc_res_xhigh_po_2p85_2_1/Rin VSS VDD sky130_asc_res_xhigh_po_2p85_2_1/a_2723_115#
+ VSS sky130_asc_res_xhigh_po_2p85_2
Xsky130_asc_res_xhigh_po_2p85_1_12 sky130_asc_res_xhigh_po_2p85_1_12/Rin sky130_asc_res_xhigh_po_2p85_1_11/Rin
+ VDD VSS sky130_asc_res_xhigh_po_2p85_1_12/a_2148_115# sky130_asc_res_xhigh_po_2p85_1
Xsky130_asc_res_xhigh_po_2p85_1_23 sky130_asc_res_xhigh_po_2p85_1_23/Rin sky130_asc_res_xhigh_po_2p85_1_22/Rin
+ VDD VSS sky130_asc_res_xhigh_po_2p85_1_23/a_2148_115# sky130_asc_res_xhigh_po_2p85_1
Xsky130_asc_res_xhigh_po_2p85_1_13 sky130_asc_res_xhigh_po_2p85_1_13/Rin sky130_asc_res_xhigh_po_2p85_1_12/Rin
+ VDD VSS sky130_asc_res_xhigh_po_2p85_1_13/a_2148_115# sky130_asc_res_xhigh_po_2p85_1
Xsky130_asc_res_xhigh_po_2p85_1_24 sky130_asc_res_xhigh_po_2p85_1_24/Rin sky130_asc_res_xhigh_po_2p85_1_23/Rin
+ VDD VSS sky130_asc_res_xhigh_po_2p85_1_24/a_2148_115# sky130_asc_res_xhigh_po_2p85_1
Xsky130_asc_pfet_01v8_lvt_12_0 VDD VDD va VSS VDD VSS sky130_asc_pfet_01v8_lvt_12
Xsky130_asc_res_xhigh_po_2p85_1_25 sky130_asc_res_xhigh_po_2p85_1_25/Rin sky130_asc_res_xhigh_po_2p85_1_24/Rin
+ VDD VSS sky130_asc_res_xhigh_po_2p85_1_25/a_2148_115# sky130_asc_res_xhigh_po_2p85_1
Xsky130_asc_res_xhigh_po_2p85_1_14 sky130_asc_res_xhigh_po_2p85_1_14/Rin sky130_asc_res_xhigh_po_2p85_1_13/Rin
+ VDD VSS sky130_asc_res_xhigh_po_2p85_1_14/a_2148_115# sky130_asc_res_xhigh_po_2p85_1
Xsky130_asc_pfet_01v8_lvt_12_1 sky130_asc_cap_mim_m3_1_4/Cout VDD sky130_asc_nfet_01v8_lvt_1_1/GATE
+ VSS VDD VSS sky130_asc_pfet_01v8_lvt_12
Xsky130_asc_res_xhigh_po_2p85_1_15 sky130_asc_res_xhigh_po_2p85_1_15/Rin sky130_asc_res_xhigh_po_2p85_1_14/Rin
+ VDD VSS sky130_asc_res_xhigh_po_2p85_1_15/a_2148_115# sky130_asc_res_xhigh_po_2p85_1
Xsky130_asc_res_xhigh_po_2p85_1_26 sky130_asc_res_xhigh_po_2p85_1_26/Rin sky130_asc_res_xhigh_po_2p85_1_25/Rin
+ VDD VSS sky130_asc_res_xhigh_po_2p85_1_26/a_2148_115# sky130_asc_res_xhigh_po_2p85_1
Xsky130_asc_res_xhigh_po_2p85_1_16 sky130_asc_res_xhigh_po_2p85_1_18/Rin sky130_asc_res_xhigh_po_2p85_1_15/Rin
+ VDD VSS sky130_asc_res_xhigh_po_2p85_1_16/a_2148_115# sky130_asc_res_xhigh_po_2p85_1
Xsky130_asc_res_xhigh_po_2p85_1_27 sky130_asc_res_xhigh_po_2p85_1_27/Rin sky130_asc_res_xhigh_po_2p85_1_26/Rin
+ VDD VSS sky130_asc_res_xhigh_po_2p85_1_27/a_2148_115# sky130_asc_res_xhigh_po_2p85_1
Xsky130_asc_res_xhigh_po_2p85_1_28 sky130_asc_res_xhigh_po_2p85_1_28/Rin sky130_asc_res_xhigh_po_2p85_1_27/Rin
+ VDD VSS sky130_asc_res_xhigh_po_2p85_1_28/a_2148_115# sky130_asc_res_xhigh_po_2p85_1
Xsky130_asc_res_xhigh_po_2p85_1_17 sky130_asc_res_xhigh_po_2p85_1_17/Rin vb VDD VSS
+ sky130_asc_res_xhigh_po_2p85_1_17/a_2148_115# sky130_asc_res_xhigh_po_2p85_1
Xsky130_asc_nfet_01v8_lvt_9_0 porst VSS sky130_asc_cap_mim_m3_1_4/Cout VDD VSS sky130_asc_nfet_01v8_lvt_9
Xsky130_asc_res_xhigh_po_2p85_1_18 sky130_asc_res_xhigh_po_2p85_1_18/Rin sky130_asc_res_xhigh_po_2p85_1_17/Rin
+ VDD VSS sky130_asc_res_xhigh_po_2p85_1_18/a_2148_115# sky130_asc_res_xhigh_po_2p85_1
Xsky130_asc_res_xhigh_po_2p85_1_29 sky130_asc_res_xhigh_po_2p85_1_29/Rin sky130_asc_res_xhigh_po_2p85_1_28/Rin
+ VDD VSS sky130_asc_res_xhigh_po_2p85_1_29/a_2148_115# sky130_asc_res_xhigh_po_2p85_1
Xsky130_asc_pfet_01v8_lvt_6_0 sky130_asc_pfet_01v8_lvt_6_1/GATE VDD sky130_asc_cap_mim_m3_1_4/Cout
+ VSS VDD VSS sky130_asc_pfet_01v8_lvt_6
Xsky130_asc_nfet_01v8_lvt_9_1 va sky130_asc_nfet_01v8_lvt_1_1/DRAIN sky130_asc_cap_mim_m3_1_4/Cout
+ VDD VSS sky130_asc_nfet_01v8_lvt_9
Xsky130_asc_res_xhigh_po_2p85_1_19 sky130_asc_res_xhigh_po_2p85_1_19/Rin sky130_asc_res_xhigh_po_2p85_1_19/Rout
+ VDD VSS sky130_asc_res_xhigh_po_2p85_1_19/a_2148_115# sky130_asc_res_xhigh_po_2p85_1
Xsky130_asc_pfet_01v8_lvt_6_1 sky130_asc_pfet_01v8_lvt_6_1/GATE VDD sky130_asc_pfet_01v8_lvt_6_1/GATE
+ VSS VDD VSS sky130_asc_pfet_01v8_lvt_6
Xsky130_asc_pnp_05v5_W3p40L3p40_1_0 va VSS VSS VDD VSS sky130_asc_pnp_05v5_W3p40L3p40_1
Xsky130_asc_nfet_01v8_lvt_9_2 vb sky130_asc_nfet_01v8_lvt_1_1/DRAIN sky130_asc_pfet_01v8_lvt_6_1/GATE
+ VDD VSS sky130_asc_nfet_01v8_lvt_9
Xsky130_asc_cap_mim_m3_1_0 VDD sky130_asc_cap_mim_m3_1_4/Cout VDD VSS VSS sky130_asc_cap_mim_m3_1
Xsky130_asc_cap_mim_m3_1_1 VDD sky130_asc_cap_mim_m3_1_4/Cout VDD VSS VSS sky130_asc_cap_mim_m3_1
Xsky130_asc_pnp_05v5_W3p40L3p40_8_0 sky130_asc_res_xhigh_po_2p85_1_19/Rout VSS VSS
+ VDD VSS sky130_asc_pnp_05v5_W3p40L3p40_8
Xsky130_asc_cap_mim_m3_1_2 VDD sky130_asc_cap_mim_m3_1_4/Cout VDD VSS VSS sky130_asc_cap_mim_m3_1
Xsky130_asc_pnp_05v5_W3p40L3p40_8_1 sky130_asc_res_xhigh_po_2p85_1_19/Rout VSS VSS
+ VDD VSS sky130_asc_pnp_05v5_W3p40L3p40_8
Xsky130_asc_cap_mim_m3_1_3 VDD sky130_asc_cap_mim_m3_1_4/Cout VDD VSS VSS sky130_asc_cap_mim_m3_1
Xsky130_asc_pnp_05v5_W3p40L3p40_8_2 sky130_asc_res_xhigh_po_2p85_1_19/Rout VSS VSS
+ VDD VSS sky130_asc_pnp_05v5_W3p40L3p40_8
Xsky130_asc_cap_mim_m3_1_4 VDD sky130_asc_cap_mim_m3_1_4/Cout VDD VSS VSS sky130_asc_cap_mim_m3_1
Xsky130_asc_pnp_05v5_W3p40L3p40_8_3 sky130_asc_res_xhigh_po_2p85_1_19/Rout VSS VSS
+ VDD VSS sky130_asc_pnp_05v5_W3p40L3p40_8
Xsky130_asc_cap_mim_m3_1_5 va VSS VDD VSS VSS sky130_asc_cap_mim_m3_1
Xsky130_asc_cap_mim_m3_1_6 va VSS VDD VSS VSS sky130_asc_cap_mim_m3_1
Xsky130_asc_res_xhigh_po_2p85_1_0 sky130_asc_res_xhigh_po_2p85_1_0/Rin VSS VDD VSS
+ sky130_asc_res_xhigh_po_2p85_1_0/a_2148_115# sky130_asc_res_xhigh_po_2p85_1
Xsky130_asc_nfet_01v8_lvt_1_0 sky130_asc_nfet_01v8_lvt_1_1/GATE VSS sky130_asc_nfet_01v8_lvt_1_1/GATE
+ VDD VSS sky130_asc_nfet_01v8_lvt_1
Xsky130_asc_res_xhigh_po_2p85_1_1 sky130_asc_res_xhigh_po_2p85_1_1/Rin sky130_asc_res_xhigh_po_2p85_1_0/Rin
+ VDD VSS sky130_asc_res_xhigh_po_2p85_1_1/a_2148_115# sky130_asc_res_xhigh_po_2p85_1
Xsky130_asc_cap_mim_m3_1_7 va VSS VDD VSS VSS sky130_asc_cap_mim_m3_1
Xsky130_asc_nfet_01v8_lvt_1_1 sky130_asc_nfet_01v8_lvt_1_1/GATE VSS sky130_asc_nfet_01v8_lvt_1_1/DRAIN
+ VDD VSS sky130_asc_nfet_01v8_lvt_1
Xsky130_asc_cap_mim_m3_1_8 va VSS VDD VSS VSS sky130_asc_cap_mim_m3_1
Xsky130_asc_res_xhigh_po_2p85_1_2 sky130_asc_res_xhigh_po_2p85_1_2/Rin sky130_asc_res_xhigh_po_2p85_1_1/Rin
+ VDD VSS sky130_asc_res_xhigh_po_2p85_1_2/a_2148_115# sky130_asc_res_xhigh_po_2p85_1
Xsky130_asc_res_xhigh_po_2p85_1_3 sky130_asc_res_xhigh_po_2p85_1_3/Rin sky130_asc_res_xhigh_po_2p85_1_2/Rin
+ VDD VSS sky130_asc_res_xhigh_po_2p85_1_3/a_2148_115# sky130_asc_res_xhigh_po_2p85_1
Xsky130_asc_cap_mim_m3_1_9 va VSS VDD VSS VSS sky130_asc_cap_mim_m3_1
Xsky130_asc_res_xhigh_po_2p85_1_4 sky130_asc_res_xhigh_po_2p85_1_4/Rin sky130_asc_res_xhigh_po_2p85_1_3/Rin
+ VDD VSS sky130_asc_res_xhigh_po_2p85_1_4/a_2148_115# sky130_asc_res_xhigh_po_2p85_1
Xsky130_asc_res_xhigh_po_2p85_1_5 sky130_asc_res_xhigh_po_2p85_1_5/Rin sky130_asc_res_xhigh_po_2p85_1_4/Rin
+ VDD VSS sky130_asc_res_xhigh_po_2p85_1_5/a_2148_115# sky130_asc_res_xhigh_po_2p85_1
Xsky130_asc_res_xhigh_po_2p85_1_6 sky130_asc_res_xhigh_po_2p85_1_6/Rin sky130_asc_res_xhigh_po_2p85_1_5/Rin
+ VDD VSS sky130_asc_res_xhigh_po_2p85_1_6/a_2148_115# sky130_asc_res_xhigh_po_2p85_1
C0 sky130_asc_res_xhigh_po_2p85_1_6/Rin sky130_asc_res_xhigh_po_2p85_1_8/a_2148_115# 0.21fF
C1 vb sky130_asc_pfet_01v8_lvt_6_1/GATE 0.10fF
C2 sky130_asc_res_xhigh_po_2p85_1_22/Rin sky130_asc_res_xhigh_po_2p85_1_23/Rin 0.48fF
C3 sky130_asc_res_xhigh_po_2p85_1_28/Rin sky130_asc_res_xhigh_po_2p85_2_1/Rin 0.88fF
C4 VDD sky130_asc_res_xhigh_po_2p85_1_19/Rin 0.63fF
C5 sky130_asc_res_xhigh_po_2p85_1_11/Rin sky130_asc_res_xhigh_po_2p85_1_18/Rin 0.45fF
C6 sky130_asc_res_xhigh_po_2p85_1_23/Rin sky130_asc_pfet_01v8_lvt_6_1/GATE 0.09fF
C7 sky130_asc_res_xhigh_po_2p85_1_28/a_2148_115# sky130_asc_res_xhigh_po_2p85_1_25/Rin 0.23fF
C8 sky130_asc_cap_mim_m3_1_4/Cout VDD 2.34fF
C9 va sky130_asc_res_xhigh_po_2p85_1_24/Rin 0.67fF
C10 VDD sky130_asc_res_xhigh_po_2p85_1_2/Rin 0.11fF
C11 sky130_asc_res_xhigh_po_2p85_1_0/a_2148_115# sky130_asc_res_xhigh_po_2p85_1_1/Rin 0.20fF
C12 VDD sky130_asc_res_xhigh_po_2p85_1_15/Rin 0.11fF
C13 sky130_asc_res_xhigh_po_2p85_1_22/Rin sky130_asc_res_xhigh_po_2p85_1_21/Rin 0.45fF
C14 sky130_asc_res_xhigh_po_2p85_1_26/a_2148_115# sky130_asc_res_xhigh_po_2p85_1_22/Rin 0.20fF
C15 sky130_asc_res_xhigh_po_2p85_2_1/a_2723_115# sky130_asc_res_xhigh_po_2p85_1_28/Rin 0.20fF
C16 VDD sky130_asc_nfet_01v8_lvt_1_1/DRAIN 0.63fF
C17 sky130_asc_res_xhigh_po_2p85_1_22/a_2148_115# sky130_asc_res_xhigh_po_2p85_1_23/Rin 0.30fF
C18 sky130_asc_cap_mim_m3_1_4/Cout sky130_asc_nfet_01v8_lvt_1_1/DRAIN 0.30fF
C19 sky130_asc_res_xhigh_po_2p85_1_28/Rin sky130_asc_res_xhigh_po_2p85_1_28/a_2148_115# 0.01fF
C20 sky130_asc_res_xhigh_po_2p85_1_28/Rin sky130_asc_res_xhigh_po_2p85_1_29/Rin 0.45fF
C21 sky130_asc_res_xhigh_po_2p85_1_19/Rout sky130_asc_res_xhigh_po_2p85_1_25/Rin 1.60fF
C22 sky130_asc_res_xhigh_po_2p85_1_5/Rin sky130_asc_res_xhigh_po_2p85_1_4/a_2148_115# 0.49fF
C23 sky130_asc_res_xhigh_po_2p85_1_26/Rin sky130_asc_res_xhigh_po_2p85_1_29/a_2148_115# 0.20fF
C24 sky130_asc_res_xhigh_po_2p85_1_27/Rin sky130_asc_res_xhigh_po_2p85_1_19/Rout 0.04fF
C25 sky130_asc_res_xhigh_po_2p85_1_29/Rin sky130_asc_nfet_01v8_lvt_1_1/GATE 0.03fF
C26 sky130_asc_res_xhigh_po_2p85_2_0/Rin sky130_asc_res_xhigh_po_2p85_1_17/a_2148_115# 0.21fF
C27 sky130_asc_res_xhigh_po_2p85_1_1/a_2148_115# sky130_asc_res_xhigh_po_2p85_1_1/Rin 0.66fF
C28 VDD sky130_asc_pfet_01v8_lvt_6_1/GATE 0.09fF
C29 sky130_asc_res_xhigh_po_2p85_1_24/Rin sky130_asc_res_xhigh_po_2p85_1_25/Rin 0.03fF
C30 sky130_asc_res_xhigh_po_2p85_1_0/a_2148_115# sky130_asc_res_xhigh_po_2p85_1_0/Rin 0.53fF
C31 sky130_asc_res_xhigh_po_2p85_1_24/a_2148_115# sky130_asc_res_xhigh_po_2p85_1_23/Rin 0.05fF
C32 VDD sky130_asc_res_xhigh_po_2p85_2_1/Rin 1.27fF
C33 sky130_asc_cap_mim_m3_1_4/Cout sky130_asc_pfet_01v8_lvt_6_1/GATE 0.50fF
C34 sky130_asc_res_xhigh_po_2p85_1_17/a_2148_115# sky130_asc_res_xhigh_po_2p85_1_17/Rin 0.04fF
C35 sky130_asc_res_xhigh_po_2p85_1_27/Rin sky130_asc_res_xhigh_po_2p85_1_24/Rin 0.07fF
C36 sky130_asc_res_xhigh_po_2p85_1_14/Rin sky130_asc_res_xhigh_po_2p85_1_12/Rin -0.01fF
C37 vb sky130_asc_res_xhigh_po_2p85_1_19/Rout 0.03fF
C38 sky130_asc_res_xhigh_po_2p85_1_14/Rin sky130_asc_res_xhigh_po_2p85_1_13/a_2148_115# 0.50fF
C39 sky130_asc_res_xhigh_po_2p85_1_9/Rin sky130_asc_res_xhigh_po_2p85_1_17/a_2148_115# 0.20fF
C40 va sky130_asc_res_xhigh_po_2p85_1_27/Rin 2.09fF
C41 sky130_asc_res_xhigh_po_2p85_1_27/a_2148_115# sky130_asc_res_xhigh_po_2p85_1_26/Rin 0.86fF
C42 VDD sky130_asc_res_xhigh_po_2p85_1_1/Rin 0.61fF
C43 sky130_asc_res_xhigh_po_2p85_1_19/a_2148_115# vb 0.20fF
C44 sky130_asc_res_xhigh_po_2p85_1_11/Rin sky130_asc_res_xhigh_po_2p85_1_14/Rin 0.05fF
C45 sky130_asc_nfet_01v8_lvt_1_1/DRAIN sky130_asc_pfet_01v8_lvt_6_1/GATE 0.19fF
C46 sky130_asc_res_xhigh_po_2p85_1_1/Rin sky130_asc_res_xhigh_po_2p85_1_2/Rin 0.04fF
C47 sky130_asc_res_xhigh_po_2p85_1_4/a_2148_115# sky130_asc_res_xhigh_po_2p85_1_4/Rin 0.70fF
C48 sky130_asc_res_xhigh_po_2p85_1_28/Rin sky130_asc_res_xhigh_po_2p85_1_24/Rin 0.03fF
C49 sky130_asc_res_xhigh_po_2p85_1_18/Rin sky130_asc_res_xhigh_po_2p85_2_0/a_2723_115# 0.19fF
C50 vbg sky130_asc_res_xhigh_po_2p85_1_7/Rin 0.45fF
C51 sky130_asc_res_xhigh_po_2p85_1_18/Rin VDD 1.77fF
C52 va vb 0.04fF
C53 sky130_asc_res_xhigh_po_2p85_1_28/Rin va 0.02fF
C54 sky130_asc_res_xhigh_po_2p85_1_11/Rin sky130_asc_res_xhigh_po_2p85_1_10/Rin 1.93fF
C55 sky130_asc_res_xhigh_po_2p85_1_19/Rout sky130_asc_res_xhigh_po_2p85_1_21/Rin 1.01fF
C56 va sky130_asc_nfet_01v8_lvt_1_1/GATE 0.46fF
C57 sky130_asc_res_xhigh_po_2p85_1_14/Rin sky130_asc_res_xhigh_po_2p85_1_14/a_2148_115# 0.97fF
C58 sky130_asc_res_xhigh_po_2p85_1_5/Rin sky130_asc_res_xhigh_po_2p85_1_4/Rin 0.38fF
C59 vbg VDD 0.64fF
C60 sky130_asc_cap_mim_m3_1_4/Cout vbg -0.15fF
C61 sky130_asc_res_xhigh_po_2p85_1_5/Rin sky130_asc_res_xhigh_po_2p85_1_6/a_2148_115# 0.36fF
C62 sky130_asc_res_xhigh_po_2p85_1_14/Rin sky130_asc_res_xhigh_po_2p85_1_13/Rin 0.05fF
C63 sky130_asc_res_xhigh_po_2p85_1_6/Rin VDD 0.13fF
C64 VDD sky130_asc_res_xhigh_po_2p85_1_0/Rin 1.11fF
C65 sky130_asc_res_xhigh_po_2p85_1_22/Rin sky130_asc_res_xhigh_po_2p85_1_22/a_2148_115# 1.26fF
C66 sky130_asc_res_xhigh_po_2p85_1_21/Rin sky130_asc_res_xhigh_po_2p85_1_24/Rin 1.69fF
C67 sky130_asc_res_xhigh_po_2p85_1_29/Rin sky130_asc_nfet_01v8_lvt_1_1/DRAIN 0.25fF
C68 sky130_asc_res_xhigh_po_2p85_1_19/a_2148_115# sky130_asc_res_xhigh_po_2p85_1_19/Rin 0.77fF
C69 sky130_asc_res_xhigh_po_2p85_1_25/a_2148_115# sky130_asc_res_xhigh_po_2p85_1_25/Rin 0.37fF
C70 VDD sky130_asc_res_xhigh_po_2p85_1_19/Rout 0.32fF
C71 sky130_asc_res_xhigh_po_2p85_2_1/a_2723_115# sky130_asc_res_xhigh_po_2p85_2_1/Rin 0.26fF
C72 sky130_asc_res_xhigh_po_2p85_1_12/Rin sky130_asc_res_xhigh_po_2p85_1_14/a_2148_115# 0.20fF
C73 sky130_asc_res_xhigh_po_2p85_1_9/a_2148_115# sky130_asc_res_xhigh_po_2p85_1_10/Rin 0.20fF
C74 sky130_asc_res_xhigh_po_2p85_1_12/Rin sky130_asc_res_xhigh_po_2p85_1_13/Rin 0.52fF
C75 sky130_asc_res_xhigh_po_2p85_1_28/Rin sky130_asc_res_xhigh_po_2p85_1_25/Rin 0.22fF
C76 VDD sky130_asc_res_xhigh_po_2p85_1_24/Rin 2.81fF
C77 VDD sky130_asc_res_xhigh_po_2p85_1_3/Rin 0.21fF
C78 sky130_asc_res_xhigh_po_2p85_1_28/Rin sky130_asc_res_xhigh_po_2p85_1_27/Rin 0.03fF
C79 sky130_asc_res_xhigh_po_2p85_1_6/a_2148_115# sky130_asc_res_xhigh_po_2p85_1_4/Rin 0.20fF
C80 va VDD 3.77fF
C81 sky130_asc_res_xhigh_po_2p85_1_18/a_2148_115# sky130_asc_res_xhigh_po_2p85_1_15/Rin 0.20fF
C82 sky130_asc_res_xhigh_po_2p85_1_21/a_2148_115# sky130_asc_res_xhigh_po_2p85_1_25/Rin 0.34fF
C83 sky130_asc_cap_mim_m3_1_4/Cout va 0.93fF
C84 sky130_asc_res_xhigh_po_2p85_1_7/a_2148_115# sky130_asc_res_xhigh_po_2p85_1_0/Rin 0.20fF
C85 sky130_asc_res_xhigh_po_2p85_1_9/Rin sky130_asc_res_xhigh_po_2p85_1_10/Rin 0.63fF
C86 porst sky130_asc_nfet_01v8_lvt_1_1/GATE 3.36fF
C87 sky130_asc_res_xhigh_po_2p85_2_1/a_2723_115# sky130_asc_res_xhigh_po_2p85_1_29/Rin -0.37fF
C88 sky130_asc_res_xhigh_po_2p85_1_14/Rin sky130_asc_res_xhigh_po_2p85_1_15/Rin 0.58fF
C89 sky130_asc_res_xhigh_po_2p85_1_21/Rin sky130_asc_res_xhigh_po_2p85_1_25/Rin 0.39fF
C90 sky130_asc_res_xhigh_po_2p85_1_22/Rin sky130_asc_res_xhigh_po_2p85_1_24/Rin 0.45fF
C91 sky130_asc_res_xhigh_po_2p85_1_11/Rin sky130_asc_res_xhigh_po_2p85_1_9/Rin 0.62fF
C92 sky130_asc_res_xhigh_po_2p85_1_5/Rin sky130_asc_res_xhigh_po_2p85_1_3/Rin 0.28fF
C93 vb sky130_asc_nfet_01v8_lvt_1_1/GATE 0.04fF
C94 sky130_asc_res_xhigh_po_2p85_1_13/Rin sky130_asc_res_xhigh_po_2p85_1_14/a_2148_115# 0.29fF
C95 VDD sky130_asc_res_xhigh_po_2p85_1_10/Rin 0.11fF
C96 VDD sky130_asc_res_xhigh_po_2p85_1_12/Rin 0.11fF
C97 sky130_asc_pfet_01v8_lvt_6_1/GATE sky130_asc_res_xhigh_po_2p85_1_24/Rin 0.12fF
C98 sky130_asc_res_xhigh_po_2p85_1_24/Rin sky130_asc_res_xhigh_po_2p85_2_1/Rin 0.12fF
C99 sky130_asc_res_xhigh_po_2p85_1_27/Rin sky130_asc_res_xhigh_po_2p85_1_29/a_2148_115# 0.23fF
C100 sky130_asc_res_xhigh_po_2p85_1_25/a_2148_115# sky130_asc_res_xhigh_po_2p85_1_21/Rin 0.30fF
C101 sky130_asc_res_xhigh_po_2p85_1_5/Rin sky130_asc_res_xhigh_po_2p85_1_8/a_2148_115# 0.20fF
C102 VDD sky130_asc_res_xhigh_po_2p85_1_25/Rin 3.79fF
C103 va sky130_asc_res_xhigh_po_2p85_2_1/Rin 0.67fF
C104 sky130_asc_res_xhigh_po_2p85_2_0/Rin sky130_asc_res_xhigh_po_2p85_1_17/Rin 0.10fF
C105 sky130_asc_res_xhigh_po_2p85_1_11/Rin VDD 0.45fF
C106 sky130_asc_res_xhigh_po_2p85_1_13/a_2148_115# sky130_asc_res_xhigh_po_2p85_1_15/Rin 0.20fF
C107 VDD sky130_asc_res_xhigh_po_2p85_1_27/Rin 0.27fF
C108 sky130_asc_res_xhigh_po_2p85_1_28/Rin sky130_asc_res_xhigh_po_2p85_1_21/Rin 0.52fF
C109 sky130_asc_res_xhigh_po_2p85_1_9/a_2148_115# sky130_asc_res_xhigh_po_2p85_1_9/Rin 0.61fF
C110 sky130_asc_res_xhigh_po_2p85_1_27/a_2148_115# sky130_asc_res_xhigh_po_2p85_1_25/Rin 0.20fF
C111 sky130_asc_res_xhigh_po_2p85_1_11/Rin sky130_asc_res_xhigh_po_2p85_1_15/Rin 0.45fF
C112 vb sky130_asc_res_xhigh_po_2p85_1_19/Rin 0.62fF
C113 sky130_asc_res_xhigh_po_2p85_1_3/Rin sky130_asc_res_xhigh_po_2p85_1_4/Rin 0.45fF
C114 VDD porst 0.50fF
C115 sky130_asc_cap_mim_m3_1_4/Cout porst 2.06fF
C116 sky130_asc_res_xhigh_po_2p85_1_6/a_2148_115# sky130_asc_res_xhigh_po_2p85_1_3/Rin 0.20fF
C117 sky130_asc_res_xhigh_po_2p85_1_18/Rin sky130_asc_res_xhigh_po_2p85_1_18/a_2148_115# 0.43fF
C118 VDD vb 2.46fF
C119 sky130_asc_cap_mim_m3_1_4/Cout vb 0.77fF
C120 sky130_asc_res_xhigh_po_2p85_1_28/Rin VDD 1.92fF
C121 sky130_asc_res_xhigh_po_2p85_1_24/Rin sky130_asc_res_xhigh_po_2p85_1_28/a_2148_115# 0.23fF
C122 VDD sky130_asc_res_xhigh_po_2p85_1_23/Rin 0.11fF
C123 VDD sky130_asc_nfet_01v8_lvt_1_1/GATE 4.11fF
C124 sky130_asc_res_xhigh_po_2p85_2_0/Rin sky130_asc_res_xhigh_po_2p85_2_0/a_2723_115# 0.22fF
C125 sky130_asc_cap_mim_m3_1_4/Cout sky130_asc_nfet_01v8_lvt_1_1/GATE 1.56fF
C126 sky130_asc_res_xhigh_po_2p85_2_0/Rin VDD 1.23fF
C127 sky130_asc_res_xhigh_po_2p85_1_26/a_2148_115# sky130_asc_res_xhigh_po_2p85_1_21/Rin 0.20fF
C128 sky130_asc_res_xhigh_po_2p85_1_17/Rin sky130_asc_res_xhigh_po_2p85_2_0/a_2723_115# 0.56fF
C129 VDD sky130_asc_res_xhigh_po_2p85_1_17/Rin 0.39fF
C130 sky130_asc_res_xhigh_po_2p85_1_29/Rin sky130_asc_res_xhigh_po_2p85_1_30/a_2148_115# -0.28fF
C131 sky130_asc_res_xhigh_po_2p85_1_26/Rin sky130_asc_res_xhigh_po_2p85_1_25/Rin 0.45fF
C132 sky130_asc_res_xhigh_po_2p85_1_27/Rin sky130_asc_res_xhigh_po_2p85_2_1/Rin 0.03fF
C133 sky130_asc_res_xhigh_po_2p85_1_3/Rin sky130_asc_res_xhigh_po_2p85_1_0/Rin 0.03fF
C134 sky130_asc_res_xhigh_po_2p85_1_7/Rin VDD 0.11fF
C135 sky130_asc_res_xhigh_po_2p85_1_9/Rin VDD 0.97fF
C136 VDD sky130_asc_res_xhigh_po_2p85_1_21/Rin 2.08fF
C137 sky130_asc_res_xhigh_po_2p85_1_25/a_2148_115# sky130_asc_res_xhigh_po_2p85_2_1/Rin 0.30fF
C138 sky130_asc_res_xhigh_po_2p85_1_1/a_2148_115# sky130_asc_res_xhigh_po_2p85_1_2/Rin 0.20fF
C139 sky130_asc_nfet_01v8_lvt_1_1/DRAIN sky130_asc_nfet_01v8_lvt_1_1/GATE 0.83fF
C140 VDD VSS 1041.96fF
C141 porst VSS 30.18fF
C142 sky130_asc_res_xhigh_po_2p85_1_5/Rin VSS 3.87fF
C143 sky130_asc_res_xhigh_po_2p85_1_29/Rin VSS 4.95fF
C144 sky130_asc_res_xhigh_po_2p85_1_2/Rin VSS 3.89fF
C145 sky130_asc_res_xhigh_po_2p85_1_3/Rin VSS 5.31fF
C146 sky130_asc_res_xhigh_po_2p85_1_7/Rin VSS 3.68fF
C147 vbg VSS 22.69fF
C148 sky130_asc_res_xhigh_po_2p85_1_10/Rin VSS 2.72fF
C149 sky130_asc_res_xhigh_po_2p85_1_13/Rin VSS 5.09fF
C150 sky130_asc_res_xhigh_po_2p85_1_25/Rin VSS 8.60fF
C151 sky130_asc_nfet_01v8_lvt_1_1/DRAIN VSS 6.15fF
C152 sky130_asc_res_xhigh_po_2p85_1_24/Rin VSS 7.75fF
C153 sky130_asc_res_xhigh_po_2p85_1_19/Rout VSS 56.79fF
C154 sky130_asc_nfet_01v8_lvt_1_1/GATE VSS 9.55fF
C155 sky130_asc_pfet_01v8_lvt_6_1/GATE VSS 10.49fF
C156 sky130_asc_res_xhigh_po_2p85_1_6/Rin VSS 4.12fF
C157 sky130_asc_res_xhigh_po_2p85_1_6/a_2148_115# VSS 2.70fF
C158 sky130_asc_res_xhigh_po_2p85_1_5/a_2148_115# VSS 2.70fF
C159 sky130_asc_res_xhigh_po_2p85_1_4/Rin VSS 3.13fF
C160 sky130_asc_res_xhigh_po_2p85_1_4/a_2148_115# VSS 2.70fF
C161 sky130_asc_res_xhigh_po_2p85_1_3/a_2148_115# VSS 2.70fF
C162 sky130_asc_res_xhigh_po_2p85_1_1/Rin VSS 3.62fF
C163 sky130_asc_res_xhigh_po_2p85_1_2/a_2148_115# VSS 2.70fF
C164 sky130_asc_res_xhigh_po_2p85_1_0/Rin VSS 3.61fF
C165 sky130_asc_res_xhigh_po_2p85_1_1/a_2148_115# VSS 2.70fF
C166 sky130_asc_res_xhigh_po_2p85_1_0/a_2148_115# VSS 2.70fF
C167 sky130_asc_cap_mim_m3_1_4/Cout VSS 124.81fF
C168 sky130_asc_res_xhigh_po_2p85_1_19/a_2148_115# VSS 2.70fF
C169 sky130_asc_res_xhigh_po_2p85_1_29/a_2148_115# VSS 2.70fF
C170 sky130_asc_res_xhigh_po_2p85_1_18/Rin VSS 2.69fF
C171 sky130_asc_res_xhigh_po_2p85_1_18/a_2148_115# VSS 2.70fF
C172 sky130_asc_res_xhigh_po_2p85_1_17/Rin VSS 3.69fF
C173 sky130_asc_res_xhigh_po_2p85_1_17/a_2148_115# VSS 2.70fF
C174 sky130_asc_res_xhigh_po_2p85_1_28/Rin VSS 7.24fF
C175 sky130_asc_res_xhigh_po_2p85_1_28/a_2148_115# VSS 2.70fF
C176 sky130_asc_res_xhigh_po_2p85_1_26/Rin VSS 3.05fF
C177 sky130_asc_res_xhigh_po_2p85_1_27/Rin VSS 4.90fF
C178 sky130_asc_res_xhigh_po_2p85_1_27/a_2148_115# VSS 2.70fF
C179 sky130_asc_res_xhigh_po_2p85_1_15/Rin VSS 3.59fF
C180 sky130_asc_res_xhigh_po_2p85_1_16/a_2148_115# VSS 2.70fF
C181 sky130_asc_res_xhigh_po_2p85_1_26/a_2148_115# VSS 2.70fF
C182 sky130_asc_res_xhigh_po_2p85_1_14/Rin VSS 3.69fF
C183 sky130_asc_res_xhigh_po_2p85_1_15/a_2148_115# VSS 2.70fF
C184 sky130_asc_res_xhigh_po_2p85_1_14/a_2148_115# VSS 2.70fF
C185 sky130_asc_res_xhigh_po_2p85_1_25/a_2148_115# VSS 2.70fF
C186 sky130_asc_res_xhigh_po_2p85_1_23/Rin VSS 4.57fF
C187 sky130_asc_res_xhigh_po_2p85_1_24/a_2148_115# VSS 2.70fF
C188 sky130_asc_res_xhigh_po_2p85_1_12/Rin VSS 4.20fF
C189 sky130_asc_res_xhigh_po_2p85_1_13/a_2148_115# VSS 2.70fF
C190 sky130_asc_res_xhigh_po_2p85_1_23/a_2148_115# VSS 2.70fF
C191 sky130_asc_res_xhigh_po_2p85_1_12/a_2148_115# VSS 2.70fF
C192 sky130_asc_res_xhigh_po_2p85_2_1/Rin VSS 3.58fF
C193 sky130_asc_res_xhigh_po_2p85_2_1/a_2723_115# VSS 2.70fF
C194 sky130_asc_res_xhigh_po_2p85_1_11/Rin VSS 3.68fF
C195 sky130_asc_res_xhigh_po_2p85_1_11/a_2148_115# VSS 2.70fF
C196 sky130_asc_res_xhigh_po_2p85_1_22/Rin VSS 2.60fF
C197 sky130_asc_res_xhigh_po_2p85_1_22/a_2148_115# VSS 2.70fF
C198 sky130_asc_res_xhigh_po_2p85_2_0/a_2723_115# VSS 2.70fF
C199 sky130_asc_res_xhigh_po_2p85_1_9/Rin VSS 3.68fF
C200 sky130_asc_res_xhigh_po_2p85_1_10/a_2148_115# VSS 2.70fF
C201 sky130_asc_res_xhigh_po_2p85_1_21/Rin VSS 7.17fF
C202 sky130_asc_res_xhigh_po_2p85_1_21/a_2148_115# VSS 2.70fF
C203 sky130_asc_res_xhigh_po_2p85_1_19/Rin VSS 3.83fF
C204 sky130_asc_res_xhigh_po_2p85_1_20/a_2148_115# VSS 2.70fF
C205 sky130_asc_res_xhigh_po_2p85_1_30/a_2148_115# VSS 2.70fF
C206 va VSS 75.00fF
C207 vb VSS 43.67fF
C208 sky130_asc_res_xhigh_po_2p85_2_0/Rin VSS 4.68fF
C209 sky130_asc_res_xhigh_po_2p85_1_9/a_2148_115# VSS 2.70fF
C210 sky130_asc_res_xhigh_po_2p85_1_8/a_2148_115# VSS 2.70fF
C211 sky130_asc_res_xhigh_po_2p85_1_7/a_2148_115# VSS 2.90fF
.ends

