magic
tech sky130A
magscale 1 2
timestamp 1652011718
<< locali >>
rect -18 1850 152 1910
rect 212 1850 552 1910
rect 612 1850 952 1910
rect 1012 1850 1352 1910
rect 1412 1850 1752 1910
rect 1812 1850 2152 1910
rect 2212 1850 2552 1910
rect 2612 1850 2952 1910
rect 3012 1850 3352 1910
rect 3412 1850 3752 1910
rect 3812 1850 4152 1910
rect 4212 1850 4552 1910
rect 4612 1850 4952 1910
rect 5012 1850 5352 1910
rect 5412 1850 5752 1910
rect 5812 1850 6152 1910
rect 6212 1850 6552 1910
rect 6612 1850 6952 1910
rect 7012 1850 7150 1910
rect -18 -30 152 30
rect 212 -30 552 30
rect 612 -30 952 30
rect 1012 -30 1352 30
rect 1412 -30 1752 30
rect 1812 -30 2152 30
rect 2212 -30 2552 30
rect 2612 -30 2952 30
rect 3012 -30 3352 30
rect 3412 -30 3752 30
rect 3812 -30 4152 30
rect 4212 -30 4552 30
rect 4612 -30 4952 30
rect 5012 -30 5352 30
rect 5412 -30 5752 30
rect 5812 -30 6152 30
rect 6212 -30 6552 30
rect 6612 -30 6952 30
rect 7012 -30 7150 30
<< viali >>
rect 152 1850 212 1910
rect 552 1850 612 1910
rect 952 1850 1012 1910
rect 1352 1850 1412 1910
rect 1752 1850 1812 1910
rect 2152 1850 2212 1910
rect 2552 1850 2612 1910
rect 2952 1850 3012 1910
rect 3352 1850 3412 1910
rect 3752 1850 3812 1910
rect 4152 1850 4212 1910
rect 4552 1850 4612 1910
rect 4952 1850 5012 1910
rect 5352 1850 5412 1910
rect 5752 1850 5812 1910
rect 6152 1850 6212 1910
rect 6552 1850 6612 1910
rect 6952 1850 7012 1910
rect 152 -30 212 30
rect 552 -30 612 30
rect 952 -30 1012 30
rect 1352 -30 1412 30
rect 1752 -30 1812 30
rect 2152 -30 2212 30
rect 2552 -30 2612 30
rect 2952 -30 3012 30
rect 3352 -30 3412 30
rect 3752 -30 3812 30
rect 4152 -30 4212 30
rect 4552 -30 4612 30
rect 4952 -30 5012 30
rect 5352 -30 5412 30
rect 5752 -30 5812 30
rect 6152 -30 6212 30
rect 6552 -30 6612 30
rect 6952 -30 7012 30
<< metal1 >>
rect -18 1910 7150 1940
rect -18 1850 152 1910
rect 212 1850 552 1910
rect 612 1850 952 1910
rect 1012 1850 1352 1910
rect 1412 1850 1752 1910
rect 1812 1850 2152 1910
rect 2212 1850 2552 1910
rect 2612 1850 2952 1910
rect 3012 1850 3352 1910
rect 3412 1850 3752 1910
rect 3812 1850 4152 1910
rect 4212 1850 4552 1910
rect 4612 1850 4952 1910
rect 5012 1850 5352 1910
rect 5412 1850 5752 1910
rect 5812 1850 6152 1910
rect 6212 1850 6552 1910
rect 6612 1850 6952 1910
rect 7012 1850 7150 1910
rect -18 1820 7150 1850
rect -18 30 7150 60
rect -18 -30 152 30
rect 212 -30 552 30
rect 612 -30 952 30
rect 1012 -30 1352 30
rect 1412 -30 1752 30
rect 1812 -30 2152 30
rect 2212 -30 2552 30
rect 2612 -30 2952 30
rect 3012 -30 3352 30
rect 3412 -30 3752 30
rect 3812 -30 4152 30
rect 4212 -30 4552 30
rect 4612 -30 4952 30
rect 5012 -30 5352 30
rect 5412 -30 5752 30
rect 5812 -30 6152 30
rect 6212 -30 6552 30
rect 6612 -30 6952 30
rect 7012 -30 7150 30
rect -18 -60 7150 -30
<< metal3 >>
rect -20 1650 7150 1690
rect -20 1622 7151 1650
rect -20 1078 596 1622
rect 660 1078 1315 1622
rect 1379 1078 2034 1622
rect 2098 1078 2753 1622
rect 2817 1078 3472 1622
rect 3536 1078 4191 1622
rect 4255 1078 4910 1622
rect 4974 1078 5629 1622
rect 5693 1078 6348 1622
rect 6412 1078 7067 1622
rect 7131 1078 7151 1622
rect -20 1050 7151 1078
rect -20 950 7150 1050
rect -20 922 7151 950
rect -20 378 596 922
rect 660 378 1315 922
rect 1379 378 2034 922
rect 2098 378 2753 922
rect 2817 378 3472 922
rect 3536 378 4191 922
rect 4255 378 4910 922
rect 4974 378 5629 922
rect 5693 378 6348 922
rect 6412 378 7067 922
rect 7131 378 7151 922
rect -20 350 7151 378
<< via3 >>
rect 596 1078 660 1622
rect 1315 1078 1379 1622
rect 2034 1078 2098 1622
rect 2753 1078 2817 1622
rect 3472 1078 3536 1622
rect 4191 1078 4255 1622
rect 4910 1078 4974 1622
rect 5629 1078 5693 1622
rect 6348 1078 6412 1622
rect 7067 1078 7131 1622
rect 596 378 660 922
rect 1315 378 1379 922
rect 2034 378 2098 922
rect 2753 378 2817 922
rect 3472 378 3536 922
rect 4191 378 4255 922
rect 4910 378 4974 922
rect 5629 378 5693 922
rect 6348 378 6412 922
rect 7067 378 7131 922
<< mimcap >>
rect 81 1510 481 1550
rect 81 1190 121 1510
rect 441 1190 481 1510
rect 81 1150 481 1190
rect 800 1510 1200 1550
rect 800 1190 840 1510
rect 1160 1190 1200 1510
rect 800 1150 1200 1190
rect 1519 1510 1919 1550
rect 1519 1190 1559 1510
rect 1879 1190 1919 1510
rect 1519 1150 1919 1190
rect 2238 1510 2638 1550
rect 2238 1190 2278 1510
rect 2598 1190 2638 1510
rect 2238 1150 2638 1190
rect 2957 1510 3357 1550
rect 2957 1190 2997 1510
rect 3317 1190 3357 1510
rect 2957 1150 3357 1190
rect 3676 1510 4076 1550
rect 3676 1190 3716 1510
rect 4036 1190 4076 1510
rect 3676 1150 4076 1190
rect 4395 1510 4795 1550
rect 4395 1190 4435 1510
rect 4755 1190 4795 1510
rect 4395 1150 4795 1190
rect 5114 1510 5514 1550
rect 5114 1190 5154 1510
rect 5474 1190 5514 1510
rect 5114 1150 5514 1190
rect 5833 1510 6233 1550
rect 5833 1190 5873 1510
rect 6193 1190 6233 1510
rect 5833 1150 6233 1190
rect 6552 1510 6952 1550
rect 6552 1190 6592 1510
rect 6912 1190 6952 1510
rect 6552 1150 6952 1190
rect 81 810 481 850
rect 81 490 121 810
rect 441 490 481 810
rect 81 450 481 490
rect 800 810 1200 850
rect 800 490 840 810
rect 1160 490 1200 810
rect 800 450 1200 490
rect 1519 810 1919 850
rect 1519 490 1559 810
rect 1879 490 1919 810
rect 1519 450 1919 490
rect 2238 810 2638 850
rect 2238 490 2278 810
rect 2598 490 2638 810
rect 2238 450 2638 490
rect 2957 810 3357 850
rect 2957 490 2997 810
rect 3317 490 3357 810
rect 2957 450 3357 490
rect 3676 810 4076 850
rect 3676 490 3716 810
rect 4036 490 4076 810
rect 3676 450 4076 490
rect 4395 810 4795 850
rect 4395 490 4435 810
rect 4755 490 4795 810
rect 4395 450 4795 490
rect 5114 810 5514 850
rect 5114 490 5154 810
rect 5474 490 5514 810
rect 5114 450 5514 490
rect 5833 810 6233 850
rect 5833 490 5873 810
rect 6193 490 6233 810
rect 5833 450 6233 490
rect 6552 810 6952 850
rect 6552 490 6592 810
rect 6912 490 6952 810
rect 6552 450 6952 490
<< mimcapcontact >>
rect 121 1190 441 1510
rect 840 1190 1160 1510
rect 1559 1190 1879 1510
rect 2278 1190 2598 1510
rect 2997 1190 3317 1510
rect 3716 1190 4036 1510
rect 4435 1190 4755 1510
rect 5154 1190 5474 1510
rect 5873 1190 6193 1510
rect 6592 1190 6912 1510
rect 121 490 441 810
rect 840 490 1160 810
rect 1559 490 1879 810
rect 2278 490 2598 810
rect 2997 490 3317 810
rect 3716 490 4036 810
rect 4435 490 4755 810
rect 5154 490 5474 810
rect 5873 490 6193 810
rect 6592 490 6912 810
<< metal4 >>
rect 580 1622 676 1638
rect 120 1511 440 1530
rect 120 1510 442 1511
rect 120 1190 121 1510
rect 441 1190 442 1510
rect 120 1189 442 1190
rect 120 811 440 1189
rect 580 1078 596 1622
rect 660 1078 676 1622
rect 1299 1622 1395 1638
rect 840 1511 1160 1530
rect 839 1510 1161 1511
rect 839 1190 840 1510
rect 1160 1190 1161 1510
rect 839 1189 1161 1190
rect 580 1062 676 1078
rect 580 922 676 938
rect 120 810 442 811
rect 120 490 121 810
rect 441 490 442 810
rect 120 489 442 490
rect 120 290 440 489
rect 580 378 596 922
rect 660 378 676 922
rect 840 811 1160 1189
rect 1299 1078 1315 1622
rect 1379 1078 1395 1622
rect 2018 1622 2114 1638
rect 1560 1511 1880 1530
rect 1558 1510 1880 1511
rect 1558 1190 1559 1510
rect 1879 1190 1880 1510
rect 1558 1189 1880 1190
rect 1299 1062 1395 1078
rect 1299 922 1395 938
rect 839 810 1161 811
rect 839 490 840 810
rect 1160 490 1161 810
rect 839 489 1161 490
rect 580 362 676 378
rect 840 290 1160 489
rect 1299 378 1315 922
rect 1379 378 1395 922
rect 1560 811 1880 1189
rect 2018 1078 2034 1622
rect 2098 1078 2114 1622
rect 2737 1622 2833 1638
rect 2280 1511 2600 1530
rect 2277 1510 2600 1511
rect 2277 1190 2278 1510
rect 2598 1190 2600 1510
rect 2277 1189 2600 1190
rect 2018 1062 2114 1078
rect 1558 810 1880 811
rect 1558 490 1559 810
rect 1879 490 1880 810
rect 1558 489 1880 490
rect 1299 362 1395 378
rect 1560 290 1880 489
rect 2018 922 2114 938
rect 2018 378 2034 922
rect 2098 378 2114 922
rect 2280 811 2600 1189
rect 2737 1078 2753 1622
rect 2817 1078 2833 1622
rect 3456 1622 3552 1638
rect 3000 1511 3320 1530
rect 2996 1510 3320 1511
rect 2996 1190 2997 1510
rect 3317 1190 3320 1510
rect 2996 1189 3320 1190
rect 2737 1062 2833 1078
rect 2277 810 2600 811
rect 2277 490 2278 810
rect 2598 490 2600 810
rect 2277 489 2600 490
rect 2018 362 2114 378
rect 2280 290 2600 489
rect 2737 922 2833 938
rect 2737 378 2753 922
rect 2817 378 2833 922
rect 3000 811 3320 1189
rect 3456 1078 3472 1622
rect 3536 1078 3552 1622
rect 4175 1622 4271 1638
rect 3720 1511 4040 1530
rect 3715 1510 4040 1511
rect 3715 1190 3716 1510
rect 4036 1190 4040 1510
rect 3715 1189 4040 1190
rect 3456 1062 3552 1078
rect 2996 810 3320 811
rect 2996 490 2997 810
rect 3317 490 3320 810
rect 2996 489 3320 490
rect 2737 362 2833 378
rect 3000 290 3320 489
rect 3456 922 3552 938
rect 3456 378 3472 922
rect 3536 378 3552 922
rect 3720 811 4040 1189
rect 4175 1078 4191 1622
rect 4255 1078 4271 1622
rect 4894 1622 4990 1638
rect 4440 1511 4760 1530
rect 4434 1510 4760 1511
rect 4434 1190 4435 1510
rect 4755 1190 4760 1510
rect 4434 1189 4760 1190
rect 4175 1062 4271 1078
rect 3715 810 4040 811
rect 3715 490 3716 810
rect 4036 490 4040 810
rect 3715 489 4040 490
rect 3456 362 3552 378
rect 3720 290 4040 489
rect 4175 922 4271 938
rect 4175 378 4191 922
rect 4255 378 4271 922
rect 4440 811 4760 1189
rect 4894 1078 4910 1622
rect 4974 1078 4990 1622
rect 5613 1622 5709 1638
rect 5160 1511 5480 1530
rect 5153 1510 5480 1511
rect 5153 1190 5154 1510
rect 5474 1190 5480 1510
rect 5153 1189 5480 1190
rect 4894 1062 4990 1078
rect 4434 810 4760 811
rect 4434 490 4435 810
rect 4755 490 4760 810
rect 4434 489 4760 490
rect 4175 362 4271 378
rect 4440 290 4760 489
rect 4894 922 4990 938
rect 4894 378 4910 922
rect 4974 378 4990 922
rect 5160 811 5480 1189
rect 5613 1078 5629 1622
rect 5693 1078 5709 1622
rect 6332 1622 6428 1638
rect 5880 1511 6200 1530
rect 5872 1510 6200 1511
rect 5872 1190 5873 1510
rect 6193 1190 6200 1510
rect 5872 1189 6200 1190
rect 5613 1062 5709 1078
rect 5153 810 5480 811
rect 5153 490 5154 810
rect 5474 490 5480 810
rect 5153 489 5480 490
rect 4894 362 4990 378
rect 5160 290 5480 489
rect 5613 922 5709 938
rect 5613 378 5629 922
rect 5693 378 5709 922
rect 5880 811 6200 1189
rect 6332 1078 6348 1622
rect 6412 1078 6428 1622
rect 7051 1622 7147 1638
rect 6600 1511 6920 1530
rect 6591 1510 6920 1511
rect 6591 1190 6592 1510
rect 6912 1190 6920 1510
rect 6591 1189 6920 1190
rect 6332 1062 6428 1078
rect 5872 810 6200 811
rect 5872 490 5873 810
rect 6193 490 6200 810
rect 5872 489 6200 490
rect 5613 362 5709 378
rect 5880 290 6200 489
rect 6332 922 6428 938
rect 6332 378 6348 922
rect 6412 378 6428 922
rect 6600 811 6920 1189
rect 7051 1078 7067 1622
rect 7131 1078 7147 1622
rect 7051 1062 7147 1078
rect 6591 810 6920 811
rect 6591 490 6592 810
rect 6912 490 6920 810
rect 6591 489 6920 490
rect 6332 362 6428 378
rect 6600 290 6920 489
rect 7051 922 7147 938
rect 7051 378 7067 922
rect 7131 378 7147 922
rect 7051 362 7147 378
rect -18 190 7150 290
<< labels >>
flabel metal3 -20 1630 40 1690 1 FreeSans 800 0 0 0 c0
port 1 n default bidirectional
flabel metal4 -18 210 42 270 1 FreeSans 800 0 0 0 c1
port 2 n default bidirectional
flabel metal1 -18 1850 42 1910 1 FreeSans 800 0 0 0 VPWR
port 3 n power bidirectional
flabel metal1 -18 -30 42 30 1 FreeSans 800 0 0 0 VGND
port 4 n ground bidirectional
<< properties >>
string FIXED_BBOX 0 0 7171 1880
string LEFclass CORE
string LEFsite unitasc
<< end >>
