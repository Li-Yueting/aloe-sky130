magic
tech sky130A
magscale 1 2
timestamp 1652146752
<< pwell >>
rect 0 1457 9380 1610
rect 0 423 153 1457
rect 1187 423 1493 1457
rect 2527 423 2833 1457
rect 3867 423 4173 1457
rect 5207 423 5513 1457
rect 6547 423 6853 1457
rect 7887 423 8193 1457
rect 9227 423 9380 1457
rect 0 270 9380 423
<< nbase >>
rect 153 423 1187 1457
rect 1493 423 2527 1457
rect 2833 423 3867 1457
rect 4173 423 5207 1457
rect 5513 423 6547 1457
rect 6853 423 7887 1457
rect 8193 423 9227 1457
<< pdiff >>
rect 330 1228 1010 1280
rect 330 1194 384 1228
rect 418 1194 474 1228
rect 508 1194 564 1228
rect 598 1194 654 1228
rect 688 1194 744 1228
rect 778 1194 834 1228
rect 868 1194 924 1228
rect 958 1194 1010 1228
rect 330 1138 1010 1194
rect 330 1104 384 1138
rect 418 1104 474 1138
rect 508 1104 564 1138
rect 598 1104 654 1138
rect 688 1104 744 1138
rect 778 1104 834 1138
rect 868 1104 924 1138
rect 958 1104 1010 1138
rect 330 1048 1010 1104
rect 330 1014 384 1048
rect 418 1014 474 1048
rect 508 1014 564 1048
rect 598 1014 654 1048
rect 688 1014 744 1048
rect 778 1014 834 1048
rect 868 1014 924 1048
rect 958 1014 1010 1048
rect 330 958 1010 1014
rect 330 924 384 958
rect 418 924 474 958
rect 508 924 564 958
rect 598 924 654 958
rect 688 924 744 958
rect 778 924 834 958
rect 868 924 924 958
rect 958 924 1010 958
rect 330 868 1010 924
rect 330 834 384 868
rect 418 834 474 868
rect 508 834 564 868
rect 598 834 654 868
rect 688 834 744 868
rect 778 834 834 868
rect 868 834 924 868
rect 958 834 1010 868
rect 330 778 1010 834
rect 330 744 384 778
rect 418 744 474 778
rect 508 744 564 778
rect 598 744 654 778
rect 688 744 744 778
rect 778 744 834 778
rect 868 744 924 778
rect 958 744 1010 778
rect 330 688 1010 744
rect 330 654 384 688
rect 418 654 474 688
rect 508 654 564 688
rect 598 654 654 688
rect 688 654 744 688
rect 778 654 834 688
rect 868 654 924 688
rect 958 654 1010 688
rect 330 600 1010 654
rect 1670 1228 2350 1280
rect 1670 1194 1724 1228
rect 1758 1194 1814 1228
rect 1848 1194 1904 1228
rect 1938 1194 1994 1228
rect 2028 1194 2084 1228
rect 2118 1194 2174 1228
rect 2208 1194 2264 1228
rect 2298 1194 2350 1228
rect 1670 1138 2350 1194
rect 1670 1104 1724 1138
rect 1758 1104 1814 1138
rect 1848 1104 1904 1138
rect 1938 1104 1994 1138
rect 2028 1104 2084 1138
rect 2118 1104 2174 1138
rect 2208 1104 2264 1138
rect 2298 1104 2350 1138
rect 1670 1048 2350 1104
rect 1670 1014 1724 1048
rect 1758 1014 1814 1048
rect 1848 1014 1904 1048
rect 1938 1014 1994 1048
rect 2028 1014 2084 1048
rect 2118 1014 2174 1048
rect 2208 1014 2264 1048
rect 2298 1014 2350 1048
rect 1670 958 2350 1014
rect 1670 924 1724 958
rect 1758 924 1814 958
rect 1848 924 1904 958
rect 1938 924 1994 958
rect 2028 924 2084 958
rect 2118 924 2174 958
rect 2208 924 2264 958
rect 2298 924 2350 958
rect 1670 868 2350 924
rect 1670 834 1724 868
rect 1758 834 1814 868
rect 1848 834 1904 868
rect 1938 834 1994 868
rect 2028 834 2084 868
rect 2118 834 2174 868
rect 2208 834 2264 868
rect 2298 834 2350 868
rect 1670 778 2350 834
rect 1670 744 1724 778
rect 1758 744 1814 778
rect 1848 744 1904 778
rect 1938 744 1994 778
rect 2028 744 2084 778
rect 2118 744 2174 778
rect 2208 744 2264 778
rect 2298 744 2350 778
rect 1670 688 2350 744
rect 1670 654 1724 688
rect 1758 654 1814 688
rect 1848 654 1904 688
rect 1938 654 1994 688
rect 2028 654 2084 688
rect 2118 654 2174 688
rect 2208 654 2264 688
rect 2298 654 2350 688
rect 1670 600 2350 654
rect 3010 1228 3690 1280
rect 3010 1194 3064 1228
rect 3098 1194 3154 1228
rect 3188 1194 3244 1228
rect 3278 1194 3334 1228
rect 3368 1194 3424 1228
rect 3458 1194 3514 1228
rect 3548 1194 3604 1228
rect 3638 1194 3690 1228
rect 3010 1138 3690 1194
rect 3010 1104 3064 1138
rect 3098 1104 3154 1138
rect 3188 1104 3244 1138
rect 3278 1104 3334 1138
rect 3368 1104 3424 1138
rect 3458 1104 3514 1138
rect 3548 1104 3604 1138
rect 3638 1104 3690 1138
rect 3010 1048 3690 1104
rect 3010 1014 3064 1048
rect 3098 1014 3154 1048
rect 3188 1014 3244 1048
rect 3278 1014 3334 1048
rect 3368 1014 3424 1048
rect 3458 1014 3514 1048
rect 3548 1014 3604 1048
rect 3638 1014 3690 1048
rect 3010 958 3690 1014
rect 3010 924 3064 958
rect 3098 924 3154 958
rect 3188 924 3244 958
rect 3278 924 3334 958
rect 3368 924 3424 958
rect 3458 924 3514 958
rect 3548 924 3604 958
rect 3638 924 3690 958
rect 3010 868 3690 924
rect 3010 834 3064 868
rect 3098 834 3154 868
rect 3188 834 3244 868
rect 3278 834 3334 868
rect 3368 834 3424 868
rect 3458 834 3514 868
rect 3548 834 3604 868
rect 3638 834 3690 868
rect 3010 778 3690 834
rect 3010 744 3064 778
rect 3098 744 3154 778
rect 3188 744 3244 778
rect 3278 744 3334 778
rect 3368 744 3424 778
rect 3458 744 3514 778
rect 3548 744 3604 778
rect 3638 744 3690 778
rect 3010 688 3690 744
rect 3010 654 3064 688
rect 3098 654 3154 688
rect 3188 654 3244 688
rect 3278 654 3334 688
rect 3368 654 3424 688
rect 3458 654 3514 688
rect 3548 654 3604 688
rect 3638 654 3690 688
rect 3010 600 3690 654
rect 4350 1228 5030 1280
rect 4350 1194 4404 1228
rect 4438 1194 4494 1228
rect 4528 1194 4584 1228
rect 4618 1194 4674 1228
rect 4708 1194 4764 1228
rect 4798 1194 4854 1228
rect 4888 1194 4944 1228
rect 4978 1194 5030 1228
rect 4350 1138 5030 1194
rect 4350 1104 4404 1138
rect 4438 1104 4494 1138
rect 4528 1104 4584 1138
rect 4618 1104 4674 1138
rect 4708 1104 4764 1138
rect 4798 1104 4854 1138
rect 4888 1104 4944 1138
rect 4978 1104 5030 1138
rect 4350 1048 5030 1104
rect 4350 1014 4404 1048
rect 4438 1014 4494 1048
rect 4528 1014 4584 1048
rect 4618 1014 4674 1048
rect 4708 1014 4764 1048
rect 4798 1014 4854 1048
rect 4888 1014 4944 1048
rect 4978 1014 5030 1048
rect 4350 958 5030 1014
rect 4350 924 4404 958
rect 4438 924 4494 958
rect 4528 924 4584 958
rect 4618 924 4674 958
rect 4708 924 4764 958
rect 4798 924 4854 958
rect 4888 924 4944 958
rect 4978 924 5030 958
rect 4350 868 5030 924
rect 4350 834 4404 868
rect 4438 834 4494 868
rect 4528 834 4584 868
rect 4618 834 4674 868
rect 4708 834 4764 868
rect 4798 834 4854 868
rect 4888 834 4944 868
rect 4978 834 5030 868
rect 4350 778 5030 834
rect 4350 744 4404 778
rect 4438 744 4494 778
rect 4528 744 4584 778
rect 4618 744 4674 778
rect 4708 744 4764 778
rect 4798 744 4854 778
rect 4888 744 4944 778
rect 4978 744 5030 778
rect 4350 688 5030 744
rect 4350 654 4404 688
rect 4438 654 4494 688
rect 4528 654 4584 688
rect 4618 654 4674 688
rect 4708 654 4764 688
rect 4798 654 4854 688
rect 4888 654 4944 688
rect 4978 654 5030 688
rect 4350 600 5030 654
rect 5690 1228 6370 1280
rect 5690 1194 5744 1228
rect 5778 1194 5834 1228
rect 5868 1194 5924 1228
rect 5958 1194 6014 1228
rect 6048 1194 6104 1228
rect 6138 1194 6194 1228
rect 6228 1194 6284 1228
rect 6318 1194 6370 1228
rect 5690 1138 6370 1194
rect 5690 1104 5744 1138
rect 5778 1104 5834 1138
rect 5868 1104 5924 1138
rect 5958 1104 6014 1138
rect 6048 1104 6104 1138
rect 6138 1104 6194 1138
rect 6228 1104 6284 1138
rect 6318 1104 6370 1138
rect 5690 1048 6370 1104
rect 5690 1014 5744 1048
rect 5778 1014 5834 1048
rect 5868 1014 5924 1048
rect 5958 1014 6014 1048
rect 6048 1014 6104 1048
rect 6138 1014 6194 1048
rect 6228 1014 6284 1048
rect 6318 1014 6370 1048
rect 5690 958 6370 1014
rect 5690 924 5744 958
rect 5778 924 5834 958
rect 5868 924 5924 958
rect 5958 924 6014 958
rect 6048 924 6104 958
rect 6138 924 6194 958
rect 6228 924 6284 958
rect 6318 924 6370 958
rect 5690 868 6370 924
rect 5690 834 5744 868
rect 5778 834 5834 868
rect 5868 834 5924 868
rect 5958 834 6014 868
rect 6048 834 6104 868
rect 6138 834 6194 868
rect 6228 834 6284 868
rect 6318 834 6370 868
rect 5690 778 6370 834
rect 5690 744 5744 778
rect 5778 744 5834 778
rect 5868 744 5924 778
rect 5958 744 6014 778
rect 6048 744 6104 778
rect 6138 744 6194 778
rect 6228 744 6284 778
rect 6318 744 6370 778
rect 5690 688 6370 744
rect 5690 654 5744 688
rect 5778 654 5834 688
rect 5868 654 5924 688
rect 5958 654 6014 688
rect 6048 654 6104 688
rect 6138 654 6194 688
rect 6228 654 6284 688
rect 6318 654 6370 688
rect 5690 600 6370 654
rect 7030 1228 7710 1280
rect 7030 1194 7084 1228
rect 7118 1194 7174 1228
rect 7208 1194 7264 1228
rect 7298 1194 7354 1228
rect 7388 1194 7444 1228
rect 7478 1194 7534 1228
rect 7568 1194 7624 1228
rect 7658 1194 7710 1228
rect 7030 1138 7710 1194
rect 7030 1104 7084 1138
rect 7118 1104 7174 1138
rect 7208 1104 7264 1138
rect 7298 1104 7354 1138
rect 7388 1104 7444 1138
rect 7478 1104 7534 1138
rect 7568 1104 7624 1138
rect 7658 1104 7710 1138
rect 7030 1048 7710 1104
rect 7030 1014 7084 1048
rect 7118 1014 7174 1048
rect 7208 1014 7264 1048
rect 7298 1014 7354 1048
rect 7388 1014 7444 1048
rect 7478 1014 7534 1048
rect 7568 1014 7624 1048
rect 7658 1014 7710 1048
rect 7030 958 7710 1014
rect 7030 924 7084 958
rect 7118 924 7174 958
rect 7208 924 7264 958
rect 7298 924 7354 958
rect 7388 924 7444 958
rect 7478 924 7534 958
rect 7568 924 7624 958
rect 7658 924 7710 958
rect 7030 868 7710 924
rect 7030 834 7084 868
rect 7118 834 7174 868
rect 7208 834 7264 868
rect 7298 834 7354 868
rect 7388 834 7444 868
rect 7478 834 7534 868
rect 7568 834 7624 868
rect 7658 834 7710 868
rect 7030 778 7710 834
rect 7030 744 7084 778
rect 7118 744 7174 778
rect 7208 744 7264 778
rect 7298 744 7354 778
rect 7388 744 7444 778
rect 7478 744 7534 778
rect 7568 744 7624 778
rect 7658 744 7710 778
rect 7030 688 7710 744
rect 7030 654 7084 688
rect 7118 654 7174 688
rect 7208 654 7264 688
rect 7298 654 7354 688
rect 7388 654 7444 688
rect 7478 654 7534 688
rect 7568 654 7624 688
rect 7658 654 7710 688
rect 7030 600 7710 654
rect 8370 1228 9050 1280
rect 8370 1194 8424 1228
rect 8458 1194 8514 1228
rect 8548 1194 8604 1228
rect 8638 1194 8694 1228
rect 8728 1194 8784 1228
rect 8818 1194 8874 1228
rect 8908 1194 8964 1228
rect 8998 1194 9050 1228
rect 8370 1138 9050 1194
rect 8370 1104 8424 1138
rect 8458 1104 8514 1138
rect 8548 1104 8604 1138
rect 8638 1104 8694 1138
rect 8728 1104 8784 1138
rect 8818 1104 8874 1138
rect 8908 1104 8964 1138
rect 8998 1104 9050 1138
rect 8370 1048 9050 1104
rect 8370 1014 8424 1048
rect 8458 1014 8514 1048
rect 8548 1014 8604 1048
rect 8638 1014 8694 1048
rect 8728 1014 8784 1048
rect 8818 1014 8874 1048
rect 8908 1014 8964 1048
rect 8998 1014 9050 1048
rect 8370 958 9050 1014
rect 8370 924 8424 958
rect 8458 924 8514 958
rect 8548 924 8604 958
rect 8638 924 8694 958
rect 8728 924 8784 958
rect 8818 924 8874 958
rect 8908 924 8964 958
rect 8998 924 9050 958
rect 8370 868 9050 924
rect 8370 834 8424 868
rect 8458 834 8514 868
rect 8548 834 8604 868
rect 8638 834 8694 868
rect 8728 834 8784 868
rect 8818 834 8874 868
rect 8908 834 8964 868
rect 8998 834 9050 868
rect 8370 778 9050 834
rect 8370 744 8424 778
rect 8458 744 8514 778
rect 8548 744 8604 778
rect 8638 744 8694 778
rect 8728 744 8784 778
rect 8818 744 8874 778
rect 8908 744 8964 778
rect 8998 744 9050 778
rect 8370 688 9050 744
rect 8370 654 8424 688
rect 8458 654 8514 688
rect 8548 654 8604 688
rect 8638 654 8694 688
rect 8728 654 8784 688
rect 8818 654 8874 688
rect 8908 654 8964 688
rect 8998 654 9050 688
rect 8370 600 9050 654
<< pdiffc >>
rect 384 1194 418 1228
rect 474 1194 508 1228
rect 564 1194 598 1228
rect 654 1194 688 1228
rect 744 1194 778 1228
rect 834 1194 868 1228
rect 924 1194 958 1228
rect 384 1104 418 1138
rect 474 1104 508 1138
rect 564 1104 598 1138
rect 654 1104 688 1138
rect 744 1104 778 1138
rect 834 1104 868 1138
rect 924 1104 958 1138
rect 384 1014 418 1048
rect 474 1014 508 1048
rect 564 1014 598 1048
rect 654 1014 688 1048
rect 744 1014 778 1048
rect 834 1014 868 1048
rect 924 1014 958 1048
rect 384 924 418 958
rect 474 924 508 958
rect 564 924 598 958
rect 654 924 688 958
rect 744 924 778 958
rect 834 924 868 958
rect 924 924 958 958
rect 384 834 418 868
rect 474 834 508 868
rect 564 834 598 868
rect 654 834 688 868
rect 744 834 778 868
rect 834 834 868 868
rect 924 834 958 868
rect 384 744 418 778
rect 474 744 508 778
rect 564 744 598 778
rect 654 744 688 778
rect 744 744 778 778
rect 834 744 868 778
rect 924 744 958 778
rect 384 654 418 688
rect 474 654 508 688
rect 564 654 598 688
rect 654 654 688 688
rect 744 654 778 688
rect 834 654 868 688
rect 924 654 958 688
rect 1724 1194 1758 1228
rect 1814 1194 1848 1228
rect 1904 1194 1938 1228
rect 1994 1194 2028 1228
rect 2084 1194 2118 1228
rect 2174 1194 2208 1228
rect 2264 1194 2298 1228
rect 1724 1104 1758 1138
rect 1814 1104 1848 1138
rect 1904 1104 1938 1138
rect 1994 1104 2028 1138
rect 2084 1104 2118 1138
rect 2174 1104 2208 1138
rect 2264 1104 2298 1138
rect 1724 1014 1758 1048
rect 1814 1014 1848 1048
rect 1904 1014 1938 1048
rect 1994 1014 2028 1048
rect 2084 1014 2118 1048
rect 2174 1014 2208 1048
rect 2264 1014 2298 1048
rect 1724 924 1758 958
rect 1814 924 1848 958
rect 1904 924 1938 958
rect 1994 924 2028 958
rect 2084 924 2118 958
rect 2174 924 2208 958
rect 2264 924 2298 958
rect 1724 834 1758 868
rect 1814 834 1848 868
rect 1904 834 1938 868
rect 1994 834 2028 868
rect 2084 834 2118 868
rect 2174 834 2208 868
rect 2264 834 2298 868
rect 1724 744 1758 778
rect 1814 744 1848 778
rect 1904 744 1938 778
rect 1994 744 2028 778
rect 2084 744 2118 778
rect 2174 744 2208 778
rect 2264 744 2298 778
rect 1724 654 1758 688
rect 1814 654 1848 688
rect 1904 654 1938 688
rect 1994 654 2028 688
rect 2084 654 2118 688
rect 2174 654 2208 688
rect 2264 654 2298 688
rect 3064 1194 3098 1228
rect 3154 1194 3188 1228
rect 3244 1194 3278 1228
rect 3334 1194 3368 1228
rect 3424 1194 3458 1228
rect 3514 1194 3548 1228
rect 3604 1194 3638 1228
rect 3064 1104 3098 1138
rect 3154 1104 3188 1138
rect 3244 1104 3278 1138
rect 3334 1104 3368 1138
rect 3424 1104 3458 1138
rect 3514 1104 3548 1138
rect 3604 1104 3638 1138
rect 3064 1014 3098 1048
rect 3154 1014 3188 1048
rect 3244 1014 3278 1048
rect 3334 1014 3368 1048
rect 3424 1014 3458 1048
rect 3514 1014 3548 1048
rect 3604 1014 3638 1048
rect 3064 924 3098 958
rect 3154 924 3188 958
rect 3244 924 3278 958
rect 3334 924 3368 958
rect 3424 924 3458 958
rect 3514 924 3548 958
rect 3604 924 3638 958
rect 3064 834 3098 868
rect 3154 834 3188 868
rect 3244 834 3278 868
rect 3334 834 3368 868
rect 3424 834 3458 868
rect 3514 834 3548 868
rect 3604 834 3638 868
rect 3064 744 3098 778
rect 3154 744 3188 778
rect 3244 744 3278 778
rect 3334 744 3368 778
rect 3424 744 3458 778
rect 3514 744 3548 778
rect 3604 744 3638 778
rect 3064 654 3098 688
rect 3154 654 3188 688
rect 3244 654 3278 688
rect 3334 654 3368 688
rect 3424 654 3458 688
rect 3514 654 3548 688
rect 3604 654 3638 688
rect 4404 1194 4438 1228
rect 4494 1194 4528 1228
rect 4584 1194 4618 1228
rect 4674 1194 4708 1228
rect 4764 1194 4798 1228
rect 4854 1194 4888 1228
rect 4944 1194 4978 1228
rect 4404 1104 4438 1138
rect 4494 1104 4528 1138
rect 4584 1104 4618 1138
rect 4674 1104 4708 1138
rect 4764 1104 4798 1138
rect 4854 1104 4888 1138
rect 4944 1104 4978 1138
rect 4404 1014 4438 1048
rect 4494 1014 4528 1048
rect 4584 1014 4618 1048
rect 4674 1014 4708 1048
rect 4764 1014 4798 1048
rect 4854 1014 4888 1048
rect 4944 1014 4978 1048
rect 4404 924 4438 958
rect 4494 924 4528 958
rect 4584 924 4618 958
rect 4674 924 4708 958
rect 4764 924 4798 958
rect 4854 924 4888 958
rect 4944 924 4978 958
rect 4404 834 4438 868
rect 4494 834 4528 868
rect 4584 834 4618 868
rect 4674 834 4708 868
rect 4764 834 4798 868
rect 4854 834 4888 868
rect 4944 834 4978 868
rect 4404 744 4438 778
rect 4494 744 4528 778
rect 4584 744 4618 778
rect 4674 744 4708 778
rect 4764 744 4798 778
rect 4854 744 4888 778
rect 4944 744 4978 778
rect 4404 654 4438 688
rect 4494 654 4528 688
rect 4584 654 4618 688
rect 4674 654 4708 688
rect 4764 654 4798 688
rect 4854 654 4888 688
rect 4944 654 4978 688
rect 5744 1194 5778 1228
rect 5834 1194 5868 1228
rect 5924 1194 5958 1228
rect 6014 1194 6048 1228
rect 6104 1194 6138 1228
rect 6194 1194 6228 1228
rect 6284 1194 6318 1228
rect 5744 1104 5778 1138
rect 5834 1104 5868 1138
rect 5924 1104 5958 1138
rect 6014 1104 6048 1138
rect 6104 1104 6138 1138
rect 6194 1104 6228 1138
rect 6284 1104 6318 1138
rect 5744 1014 5778 1048
rect 5834 1014 5868 1048
rect 5924 1014 5958 1048
rect 6014 1014 6048 1048
rect 6104 1014 6138 1048
rect 6194 1014 6228 1048
rect 6284 1014 6318 1048
rect 5744 924 5778 958
rect 5834 924 5868 958
rect 5924 924 5958 958
rect 6014 924 6048 958
rect 6104 924 6138 958
rect 6194 924 6228 958
rect 6284 924 6318 958
rect 5744 834 5778 868
rect 5834 834 5868 868
rect 5924 834 5958 868
rect 6014 834 6048 868
rect 6104 834 6138 868
rect 6194 834 6228 868
rect 6284 834 6318 868
rect 5744 744 5778 778
rect 5834 744 5868 778
rect 5924 744 5958 778
rect 6014 744 6048 778
rect 6104 744 6138 778
rect 6194 744 6228 778
rect 6284 744 6318 778
rect 5744 654 5778 688
rect 5834 654 5868 688
rect 5924 654 5958 688
rect 6014 654 6048 688
rect 6104 654 6138 688
rect 6194 654 6228 688
rect 6284 654 6318 688
rect 7084 1194 7118 1228
rect 7174 1194 7208 1228
rect 7264 1194 7298 1228
rect 7354 1194 7388 1228
rect 7444 1194 7478 1228
rect 7534 1194 7568 1228
rect 7624 1194 7658 1228
rect 7084 1104 7118 1138
rect 7174 1104 7208 1138
rect 7264 1104 7298 1138
rect 7354 1104 7388 1138
rect 7444 1104 7478 1138
rect 7534 1104 7568 1138
rect 7624 1104 7658 1138
rect 7084 1014 7118 1048
rect 7174 1014 7208 1048
rect 7264 1014 7298 1048
rect 7354 1014 7388 1048
rect 7444 1014 7478 1048
rect 7534 1014 7568 1048
rect 7624 1014 7658 1048
rect 7084 924 7118 958
rect 7174 924 7208 958
rect 7264 924 7298 958
rect 7354 924 7388 958
rect 7444 924 7478 958
rect 7534 924 7568 958
rect 7624 924 7658 958
rect 7084 834 7118 868
rect 7174 834 7208 868
rect 7264 834 7298 868
rect 7354 834 7388 868
rect 7444 834 7478 868
rect 7534 834 7568 868
rect 7624 834 7658 868
rect 7084 744 7118 778
rect 7174 744 7208 778
rect 7264 744 7298 778
rect 7354 744 7388 778
rect 7444 744 7478 778
rect 7534 744 7568 778
rect 7624 744 7658 778
rect 7084 654 7118 688
rect 7174 654 7208 688
rect 7264 654 7298 688
rect 7354 654 7388 688
rect 7444 654 7478 688
rect 7534 654 7568 688
rect 7624 654 7658 688
rect 8424 1194 8458 1228
rect 8514 1194 8548 1228
rect 8604 1194 8638 1228
rect 8694 1194 8728 1228
rect 8784 1194 8818 1228
rect 8874 1194 8908 1228
rect 8964 1194 8998 1228
rect 8424 1104 8458 1138
rect 8514 1104 8548 1138
rect 8604 1104 8638 1138
rect 8694 1104 8728 1138
rect 8784 1104 8818 1138
rect 8874 1104 8908 1138
rect 8964 1104 8998 1138
rect 8424 1014 8458 1048
rect 8514 1014 8548 1048
rect 8604 1014 8638 1048
rect 8694 1014 8728 1048
rect 8784 1014 8818 1048
rect 8874 1014 8908 1048
rect 8964 1014 8998 1048
rect 8424 924 8458 958
rect 8514 924 8548 958
rect 8604 924 8638 958
rect 8694 924 8728 958
rect 8784 924 8818 958
rect 8874 924 8908 958
rect 8964 924 8998 958
rect 8424 834 8458 868
rect 8514 834 8548 868
rect 8604 834 8638 868
rect 8694 834 8728 868
rect 8784 834 8818 868
rect 8874 834 8908 868
rect 8964 834 8998 868
rect 8424 744 8458 778
rect 8514 744 8548 778
rect 8604 744 8638 778
rect 8694 744 8728 778
rect 8784 744 8818 778
rect 8874 744 8908 778
rect 8964 744 8998 778
rect 8424 654 8458 688
rect 8514 654 8548 688
rect 8604 654 8638 688
rect 8694 654 8728 688
rect 8784 654 8818 688
rect 8874 654 8908 688
rect 8964 654 8998 688
<< psubdiff >>
rect 26 1549 9354 1584
rect 26 1526 156 1549
rect 26 1492 60 1526
rect 94 1515 156 1526
rect 190 1515 246 1549
rect 280 1515 336 1549
rect 370 1515 426 1549
rect 460 1515 516 1549
rect 550 1515 606 1549
rect 640 1515 696 1549
rect 730 1515 786 1549
rect 820 1515 876 1549
rect 910 1515 966 1549
rect 1000 1515 1056 1549
rect 1090 1515 1146 1549
rect 1180 1526 1496 1549
rect 1180 1515 1247 1526
rect 94 1492 1247 1515
rect 1281 1492 1400 1526
rect 1434 1515 1496 1526
rect 1530 1515 1586 1549
rect 1620 1515 1676 1549
rect 1710 1515 1766 1549
rect 1800 1515 1856 1549
rect 1890 1515 1946 1549
rect 1980 1515 2036 1549
rect 2070 1515 2126 1549
rect 2160 1515 2216 1549
rect 2250 1515 2306 1549
rect 2340 1515 2396 1549
rect 2430 1515 2486 1549
rect 2520 1526 2836 1549
rect 2520 1515 2587 1526
rect 1434 1492 2587 1515
rect 2621 1492 2740 1526
rect 2774 1515 2836 1526
rect 2870 1515 2926 1549
rect 2960 1515 3016 1549
rect 3050 1515 3106 1549
rect 3140 1515 3196 1549
rect 3230 1515 3286 1549
rect 3320 1515 3376 1549
rect 3410 1515 3466 1549
rect 3500 1515 3556 1549
rect 3590 1515 3646 1549
rect 3680 1515 3736 1549
rect 3770 1515 3826 1549
rect 3860 1526 4176 1549
rect 3860 1515 3927 1526
rect 2774 1492 3927 1515
rect 3961 1492 4080 1526
rect 4114 1515 4176 1526
rect 4210 1515 4266 1549
rect 4300 1515 4356 1549
rect 4390 1515 4446 1549
rect 4480 1515 4536 1549
rect 4570 1515 4626 1549
rect 4660 1515 4716 1549
rect 4750 1515 4806 1549
rect 4840 1515 4896 1549
rect 4930 1515 4986 1549
rect 5020 1515 5076 1549
rect 5110 1515 5166 1549
rect 5200 1526 5516 1549
rect 5200 1515 5267 1526
rect 4114 1492 5267 1515
rect 5301 1492 5420 1526
rect 5454 1515 5516 1526
rect 5550 1515 5606 1549
rect 5640 1515 5696 1549
rect 5730 1515 5786 1549
rect 5820 1515 5876 1549
rect 5910 1515 5966 1549
rect 6000 1515 6056 1549
rect 6090 1515 6146 1549
rect 6180 1515 6236 1549
rect 6270 1515 6326 1549
rect 6360 1515 6416 1549
rect 6450 1515 6506 1549
rect 6540 1526 6856 1549
rect 6540 1515 6607 1526
rect 5454 1492 6607 1515
rect 6641 1492 6760 1526
rect 6794 1515 6856 1526
rect 6890 1515 6946 1549
rect 6980 1515 7036 1549
rect 7070 1515 7126 1549
rect 7160 1515 7216 1549
rect 7250 1515 7306 1549
rect 7340 1515 7396 1549
rect 7430 1515 7486 1549
rect 7520 1515 7576 1549
rect 7610 1515 7666 1549
rect 7700 1515 7756 1549
rect 7790 1515 7846 1549
rect 7880 1526 8196 1549
rect 7880 1515 7947 1526
rect 6794 1492 7947 1515
rect 7981 1492 8100 1526
rect 8134 1515 8196 1526
rect 8230 1515 8286 1549
rect 8320 1515 8376 1549
rect 8410 1515 8466 1549
rect 8500 1515 8556 1549
rect 8590 1515 8646 1549
rect 8680 1515 8736 1549
rect 8770 1515 8826 1549
rect 8860 1515 8916 1549
rect 8950 1515 9006 1549
rect 9040 1515 9096 1549
rect 9130 1515 9186 1549
rect 9220 1526 9354 1549
rect 9220 1515 9287 1526
rect 8134 1492 9287 1515
rect 9321 1492 9354 1526
rect 26 1483 9354 1492
rect 26 1436 127 1483
rect 26 1402 60 1436
rect 94 1402 127 1436
rect 1213 1436 1467 1483
rect 26 1346 127 1402
rect 26 1312 60 1346
rect 94 1312 127 1346
rect 26 1256 127 1312
rect 26 1222 60 1256
rect 94 1222 127 1256
rect 26 1166 127 1222
rect 26 1132 60 1166
rect 94 1132 127 1166
rect 26 1076 127 1132
rect 26 1042 60 1076
rect 94 1042 127 1076
rect 26 986 127 1042
rect 26 952 60 986
rect 94 952 127 986
rect 26 896 127 952
rect 26 862 60 896
rect 94 862 127 896
rect 26 806 127 862
rect 26 772 60 806
rect 94 772 127 806
rect 26 716 127 772
rect 26 682 60 716
rect 94 682 127 716
rect 26 626 127 682
rect 26 592 60 626
rect 94 592 127 626
rect 26 536 127 592
rect 26 502 60 536
rect 94 502 127 536
rect 26 446 127 502
rect 1213 1402 1247 1436
rect 1281 1402 1400 1436
rect 1434 1402 1467 1436
rect 2553 1436 2807 1483
rect 1213 1346 1467 1402
rect 1213 1312 1247 1346
rect 1281 1312 1400 1346
rect 1434 1312 1467 1346
rect 1213 1256 1467 1312
rect 1213 1222 1247 1256
rect 1281 1222 1400 1256
rect 1434 1222 1467 1256
rect 1213 1166 1467 1222
rect 1213 1132 1247 1166
rect 1281 1132 1400 1166
rect 1434 1132 1467 1166
rect 1213 1076 1467 1132
rect 1213 1042 1247 1076
rect 1281 1042 1400 1076
rect 1434 1042 1467 1076
rect 1213 986 1467 1042
rect 1213 952 1247 986
rect 1281 952 1400 986
rect 1434 952 1467 986
rect 1213 896 1467 952
rect 1213 862 1247 896
rect 1281 862 1400 896
rect 1434 862 1467 896
rect 1213 806 1467 862
rect 1213 772 1247 806
rect 1281 772 1400 806
rect 1434 772 1467 806
rect 1213 716 1467 772
rect 1213 682 1247 716
rect 1281 682 1400 716
rect 1434 682 1467 716
rect 1213 626 1467 682
rect 1213 592 1247 626
rect 1281 592 1400 626
rect 1434 592 1467 626
rect 1213 536 1467 592
rect 1213 502 1247 536
rect 1281 502 1400 536
rect 1434 502 1467 536
rect 26 412 60 446
rect 94 412 127 446
rect 26 397 127 412
rect 1213 446 1467 502
rect 2553 1402 2587 1436
rect 2621 1402 2740 1436
rect 2774 1402 2807 1436
rect 3893 1436 4147 1483
rect 2553 1346 2807 1402
rect 2553 1312 2587 1346
rect 2621 1312 2740 1346
rect 2774 1312 2807 1346
rect 2553 1256 2807 1312
rect 2553 1222 2587 1256
rect 2621 1222 2740 1256
rect 2774 1222 2807 1256
rect 2553 1166 2807 1222
rect 2553 1132 2587 1166
rect 2621 1132 2740 1166
rect 2774 1132 2807 1166
rect 2553 1076 2807 1132
rect 2553 1042 2587 1076
rect 2621 1042 2740 1076
rect 2774 1042 2807 1076
rect 2553 986 2807 1042
rect 2553 952 2587 986
rect 2621 952 2740 986
rect 2774 952 2807 986
rect 2553 896 2807 952
rect 2553 862 2587 896
rect 2621 862 2740 896
rect 2774 862 2807 896
rect 2553 806 2807 862
rect 2553 772 2587 806
rect 2621 772 2740 806
rect 2774 772 2807 806
rect 2553 716 2807 772
rect 2553 682 2587 716
rect 2621 682 2740 716
rect 2774 682 2807 716
rect 2553 626 2807 682
rect 2553 592 2587 626
rect 2621 592 2740 626
rect 2774 592 2807 626
rect 2553 536 2807 592
rect 2553 502 2587 536
rect 2621 502 2740 536
rect 2774 502 2807 536
rect 1213 412 1247 446
rect 1281 412 1400 446
rect 1434 412 1467 446
rect 1213 397 1467 412
rect 2553 446 2807 502
rect 3893 1402 3927 1436
rect 3961 1402 4080 1436
rect 4114 1402 4147 1436
rect 5233 1436 5487 1483
rect 3893 1346 4147 1402
rect 3893 1312 3927 1346
rect 3961 1312 4080 1346
rect 4114 1312 4147 1346
rect 3893 1256 4147 1312
rect 3893 1222 3927 1256
rect 3961 1222 4080 1256
rect 4114 1222 4147 1256
rect 3893 1166 4147 1222
rect 3893 1132 3927 1166
rect 3961 1132 4080 1166
rect 4114 1132 4147 1166
rect 3893 1076 4147 1132
rect 3893 1042 3927 1076
rect 3961 1042 4080 1076
rect 4114 1042 4147 1076
rect 3893 986 4147 1042
rect 3893 952 3927 986
rect 3961 952 4080 986
rect 4114 952 4147 986
rect 3893 896 4147 952
rect 3893 862 3927 896
rect 3961 862 4080 896
rect 4114 862 4147 896
rect 3893 806 4147 862
rect 3893 772 3927 806
rect 3961 772 4080 806
rect 4114 772 4147 806
rect 3893 716 4147 772
rect 3893 682 3927 716
rect 3961 682 4080 716
rect 4114 682 4147 716
rect 3893 626 4147 682
rect 3893 592 3927 626
rect 3961 592 4080 626
rect 4114 592 4147 626
rect 3893 536 4147 592
rect 3893 502 3927 536
rect 3961 502 4080 536
rect 4114 502 4147 536
rect 2553 412 2587 446
rect 2621 412 2740 446
rect 2774 412 2807 446
rect 2553 397 2807 412
rect 3893 446 4147 502
rect 5233 1402 5267 1436
rect 5301 1402 5420 1436
rect 5454 1402 5487 1436
rect 6573 1436 6827 1483
rect 5233 1346 5487 1402
rect 5233 1312 5267 1346
rect 5301 1312 5420 1346
rect 5454 1312 5487 1346
rect 5233 1256 5487 1312
rect 5233 1222 5267 1256
rect 5301 1222 5420 1256
rect 5454 1222 5487 1256
rect 5233 1166 5487 1222
rect 5233 1132 5267 1166
rect 5301 1132 5420 1166
rect 5454 1132 5487 1166
rect 5233 1076 5487 1132
rect 5233 1042 5267 1076
rect 5301 1042 5420 1076
rect 5454 1042 5487 1076
rect 5233 986 5487 1042
rect 5233 952 5267 986
rect 5301 952 5420 986
rect 5454 952 5487 986
rect 5233 896 5487 952
rect 5233 862 5267 896
rect 5301 862 5420 896
rect 5454 862 5487 896
rect 5233 806 5487 862
rect 5233 772 5267 806
rect 5301 772 5420 806
rect 5454 772 5487 806
rect 5233 716 5487 772
rect 5233 682 5267 716
rect 5301 682 5420 716
rect 5454 682 5487 716
rect 5233 626 5487 682
rect 5233 592 5267 626
rect 5301 592 5420 626
rect 5454 592 5487 626
rect 5233 536 5487 592
rect 5233 502 5267 536
rect 5301 502 5420 536
rect 5454 502 5487 536
rect 3893 412 3927 446
rect 3961 412 4080 446
rect 4114 412 4147 446
rect 3893 397 4147 412
rect 5233 446 5487 502
rect 6573 1402 6607 1436
rect 6641 1402 6760 1436
rect 6794 1402 6827 1436
rect 7913 1436 8167 1483
rect 6573 1346 6827 1402
rect 6573 1312 6607 1346
rect 6641 1312 6760 1346
rect 6794 1312 6827 1346
rect 6573 1256 6827 1312
rect 6573 1222 6607 1256
rect 6641 1222 6760 1256
rect 6794 1222 6827 1256
rect 6573 1166 6827 1222
rect 6573 1132 6607 1166
rect 6641 1132 6760 1166
rect 6794 1132 6827 1166
rect 6573 1076 6827 1132
rect 6573 1042 6607 1076
rect 6641 1042 6760 1076
rect 6794 1042 6827 1076
rect 6573 986 6827 1042
rect 6573 952 6607 986
rect 6641 952 6760 986
rect 6794 952 6827 986
rect 6573 896 6827 952
rect 6573 862 6607 896
rect 6641 862 6760 896
rect 6794 862 6827 896
rect 6573 806 6827 862
rect 6573 772 6607 806
rect 6641 772 6760 806
rect 6794 772 6827 806
rect 6573 716 6827 772
rect 6573 682 6607 716
rect 6641 682 6760 716
rect 6794 682 6827 716
rect 6573 626 6827 682
rect 6573 592 6607 626
rect 6641 592 6760 626
rect 6794 592 6827 626
rect 6573 536 6827 592
rect 6573 502 6607 536
rect 6641 502 6760 536
rect 6794 502 6827 536
rect 5233 412 5267 446
rect 5301 412 5420 446
rect 5454 412 5487 446
rect 5233 397 5487 412
rect 6573 446 6827 502
rect 7913 1402 7947 1436
rect 7981 1402 8100 1436
rect 8134 1402 8167 1436
rect 9253 1436 9354 1483
rect 7913 1346 8167 1402
rect 7913 1312 7947 1346
rect 7981 1312 8100 1346
rect 8134 1312 8167 1346
rect 7913 1256 8167 1312
rect 7913 1222 7947 1256
rect 7981 1222 8100 1256
rect 8134 1222 8167 1256
rect 7913 1166 8167 1222
rect 7913 1132 7947 1166
rect 7981 1132 8100 1166
rect 8134 1132 8167 1166
rect 7913 1076 8167 1132
rect 7913 1042 7947 1076
rect 7981 1042 8100 1076
rect 8134 1042 8167 1076
rect 7913 986 8167 1042
rect 7913 952 7947 986
rect 7981 952 8100 986
rect 8134 952 8167 986
rect 7913 896 8167 952
rect 7913 862 7947 896
rect 7981 862 8100 896
rect 8134 862 8167 896
rect 7913 806 8167 862
rect 7913 772 7947 806
rect 7981 772 8100 806
rect 8134 772 8167 806
rect 7913 716 8167 772
rect 7913 682 7947 716
rect 7981 682 8100 716
rect 8134 682 8167 716
rect 7913 626 8167 682
rect 7913 592 7947 626
rect 7981 592 8100 626
rect 8134 592 8167 626
rect 7913 536 8167 592
rect 7913 502 7947 536
rect 7981 502 8100 536
rect 8134 502 8167 536
rect 6573 412 6607 446
rect 6641 412 6760 446
rect 6794 412 6827 446
rect 6573 397 6827 412
rect 7913 446 8167 502
rect 9253 1402 9287 1436
rect 9321 1402 9354 1436
rect 9253 1346 9354 1402
rect 9253 1312 9287 1346
rect 9321 1312 9354 1346
rect 9253 1256 9354 1312
rect 9253 1222 9287 1256
rect 9321 1222 9354 1256
rect 9253 1166 9354 1222
rect 9253 1132 9287 1166
rect 9321 1132 9354 1166
rect 9253 1076 9354 1132
rect 9253 1042 9287 1076
rect 9321 1042 9354 1076
rect 9253 986 9354 1042
rect 9253 952 9287 986
rect 9321 952 9354 986
rect 9253 896 9354 952
rect 9253 862 9287 896
rect 9321 862 9354 896
rect 9253 806 9354 862
rect 9253 772 9287 806
rect 9321 772 9354 806
rect 9253 716 9354 772
rect 9253 682 9287 716
rect 9321 682 9354 716
rect 9253 626 9354 682
rect 9253 592 9287 626
rect 9321 592 9354 626
rect 9253 536 9354 592
rect 9253 502 9287 536
rect 9321 502 9354 536
rect 7913 412 7947 446
rect 7981 412 8100 446
rect 8134 412 8167 446
rect 7913 397 8167 412
rect 9253 446 9354 502
rect 9253 412 9287 446
rect 9321 412 9354 446
rect 9253 397 9354 412
rect 26 362 9354 397
rect 26 328 156 362
rect 190 328 246 362
rect 280 328 336 362
rect 370 328 426 362
rect 460 328 516 362
rect 550 328 606 362
rect 640 328 696 362
rect 730 328 786 362
rect 820 328 876 362
rect 910 328 966 362
rect 1000 328 1056 362
rect 1090 328 1146 362
rect 1180 328 1496 362
rect 1530 328 1586 362
rect 1620 328 1676 362
rect 1710 328 1766 362
rect 1800 328 1856 362
rect 1890 328 1946 362
rect 1980 328 2036 362
rect 2070 328 2126 362
rect 2160 328 2216 362
rect 2250 328 2306 362
rect 2340 328 2396 362
rect 2430 328 2486 362
rect 2520 328 2836 362
rect 2870 328 2926 362
rect 2960 328 3016 362
rect 3050 328 3106 362
rect 3140 328 3196 362
rect 3230 328 3286 362
rect 3320 328 3376 362
rect 3410 328 3466 362
rect 3500 328 3556 362
rect 3590 328 3646 362
rect 3680 328 3736 362
rect 3770 328 3826 362
rect 3860 328 4176 362
rect 4210 328 4266 362
rect 4300 328 4356 362
rect 4390 328 4446 362
rect 4480 328 4536 362
rect 4570 328 4626 362
rect 4660 328 4716 362
rect 4750 328 4806 362
rect 4840 328 4896 362
rect 4930 328 4986 362
rect 5020 328 5076 362
rect 5110 328 5166 362
rect 5200 328 5516 362
rect 5550 328 5606 362
rect 5640 328 5696 362
rect 5730 328 5786 362
rect 5820 328 5876 362
rect 5910 328 5966 362
rect 6000 328 6056 362
rect 6090 328 6146 362
rect 6180 328 6236 362
rect 6270 328 6326 362
rect 6360 328 6416 362
rect 6450 328 6506 362
rect 6540 328 6856 362
rect 6890 328 6946 362
rect 6980 328 7036 362
rect 7070 328 7126 362
rect 7160 328 7216 362
rect 7250 328 7306 362
rect 7340 328 7396 362
rect 7430 328 7486 362
rect 7520 328 7576 362
rect 7610 328 7666 362
rect 7700 328 7756 362
rect 7790 328 7846 362
rect 7880 328 8196 362
rect 8230 328 8286 362
rect 8320 328 8376 362
rect 8410 328 8466 362
rect 8500 328 8556 362
rect 8590 328 8646 362
rect 8680 328 8736 362
rect 8770 328 8826 362
rect 8860 328 8916 362
rect 8950 328 9006 362
rect 9040 328 9096 362
rect 9130 328 9186 362
rect 9220 328 9354 362
rect 26 296 9354 328
<< nsubdiff >>
rect 189 1402 1151 1421
rect 189 1368 320 1402
rect 354 1368 410 1402
rect 444 1368 500 1402
rect 534 1368 590 1402
rect 624 1368 680 1402
rect 714 1368 770 1402
rect 804 1368 860 1402
rect 894 1368 950 1402
rect 984 1368 1040 1402
rect 1074 1368 1151 1402
rect 189 1349 1151 1368
rect 189 1345 261 1349
rect 189 1311 208 1345
rect 242 1311 261 1345
rect 189 1255 261 1311
rect 1079 1326 1151 1349
rect 1079 1292 1098 1326
rect 1132 1292 1151 1326
rect 189 1221 208 1255
rect 242 1221 261 1255
rect 189 1165 261 1221
rect 189 1131 208 1165
rect 242 1131 261 1165
rect 189 1075 261 1131
rect 189 1041 208 1075
rect 242 1041 261 1075
rect 189 985 261 1041
rect 189 951 208 985
rect 242 951 261 985
rect 189 895 261 951
rect 189 861 208 895
rect 242 861 261 895
rect 189 805 261 861
rect 189 771 208 805
rect 242 771 261 805
rect 189 715 261 771
rect 189 681 208 715
rect 242 681 261 715
rect 189 625 261 681
rect 189 591 208 625
rect 242 591 261 625
rect 1079 1236 1151 1292
rect 1079 1202 1098 1236
rect 1132 1202 1151 1236
rect 1079 1146 1151 1202
rect 1079 1112 1098 1146
rect 1132 1112 1151 1146
rect 1079 1056 1151 1112
rect 1079 1022 1098 1056
rect 1132 1022 1151 1056
rect 1079 966 1151 1022
rect 1079 932 1098 966
rect 1132 932 1151 966
rect 1079 876 1151 932
rect 1079 842 1098 876
rect 1132 842 1151 876
rect 1079 786 1151 842
rect 1079 752 1098 786
rect 1132 752 1151 786
rect 1079 696 1151 752
rect 1079 662 1098 696
rect 1132 662 1151 696
rect 1079 606 1151 662
rect 189 531 261 591
rect 1079 572 1098 606
rect 1132 572 1151 606
rect 1079 531 1151 572
rect 189 512 1151 531
rect 189 478 286 512
rect 320 478 376 512
rect 410 478 466 512
rect 500 478 556 512
rect 590 478 646 512
rect 680 478 736 512
rect 770 478 826 512
rect 860 478 916 512
rect 950 478 1006 512
rect 1040 478 1151 512
rect 189 459 1151 478
rect 1529 1402 2491 1421
rect 1529 1368 1660 1402
rect 1694 1368 1750 1402
rect 1784 1368 1840 1402
rect 1874 1368 1930 1402
rect 1964 1368 2020 1402
rect 2054 1368 2110 1402
rect 2144 1368 2200 1402
rect 2234 1368 2290 1402
rect 2324 1368 2380 1402
rect 2414 1368 2491 1402
rect 1529 1349 2491 1368
rect 1529 1345 1601 1349
rect 1529 1311 1548 1345
rect 1582 1311 1601 1345
rect 1529 1255 1601 1311
rect 2419 1326 2491 1349
rect 2419 1292 2438 1326
rect 2472 1292 2491 1326
rect 1529 1221 1548 1255
rect 1582 1221 1601 1255
rect 1529 1165 1601 1221
rect 1529 1131 1548 1165
rect 1582 1131 1601 1165
rect 1529 1075 1601 1131
rect 1529 1041 1548 1075
rect 1582 1041 1601 1075
rect 1529 985 1601 1041
rect 1529 951 1548 985
rect 1582 951 1601 985
rect 1529 895 1601 951
rect 1529 861 1548 895
rect 1582 861 1601 895
rect 1529 805 1601 861
rect 1529 771 1548 805
rect 1582 771 1601 805
rect 1529 715 1601 771
rect 1529 681 1548 715
rect 1582 681 1601 715
rect 1529 625 1601 681
rect 1529 591 1548 625
rect 1582 591 1601 625
rect 2419 1236 2491 1292
rect 2419 1202 2438 1236
rect 2472 1202 2491 1236
rect 2419 1146 2491 1202
rect 2419 1112 2438 1146
rect 2472 1112 2491 1146
rect 2419 1056 2491 1112
rect 2419 1022 2438 1056
rect 2472 1022 2491 1056
rect 2419 966 2491 1022
rect 2419 932 2438 966
rect 2472 932 2491 966
rect 2419 876 2491 932
rect 2419 842 2438 876
rect 2472 842 2491 876
rect 2419 786 2491 842
rect 2419 752 2438 786
rect 2472 752 2491 786
rect 2419 696 2491 752
rect 2419 662 2438 696
rect 2472 662 2491 696
rect 2419 606 2491 662
rect 1529 531 1601 591
rect 2419 572 2438 606
rect 2472 572 2491 606
rect 2419 531 2491 572
rect 1529 512 2491 531
rect 1529 478 1626 512
rect 1660 478 1716 512
rect 1750 478 1806 512
rect 1840 478 1896 512
rect 1930 478 1986 512
rect 2020 478 2076 512
rect 2110 478 2166 512
rect 2200 478 2256 512
rect 2290 478 2346 512
rect 2380 478 2491 512
rect 1529 459 2491 478
rect 2869 1402 3831 1421
rect 2869 1368 3000 1402
rect 3034 1368 3090 1402
rect 3124 1368 3180 1402
rect 3214 1368 3270 1402
rect 3304 1368 3360 1402
rect 3394 1368 3450 1402
rect 3484 1368 3540 1402
rect 3574 1368 3630 1402
rect 3664 1368 3720 1402
rect 3754 1368 3831 1402
rect 2869 1349 3831 1368
rect 2869 1345 2941 1349
rect 2869 1311 2888 1345
rect 2922 1311 2941 1345
rect 2869 1255 2941 1311
rect 3759 1326 3831 1349
rect 3759 1292 3778 1326
rect 3812 1292 3831 1326
rect 2869 1221 2888 1255
rect 2922 1221 2941 1255
rect 2869 1165 2941 1221
rect 2869 1131 2888 1165
rect 2922 1131 2941 1165
rect 2869 1075 2941 1131
rect 2869 1041 2888 1075
rect 2922 1041 2941 1075
rect 2869 985 2941 1041
rect 2869 951 2888 985
rect 2922 951 2941 985
rect 2869 895 2941 951
rect 2869 861 2888 895
rect 2922 861 2941 895
rect 2869 805 2941 861
rect 2869 771 2888 805
rect 2922 771 2941 805
rect 2869 715 2941 771
rect 2869 681 2888 715
rect 2922 681 2941 715
rect 2869 625 2941 681
rect 2869 591 2888 625
rect 2922 591 2941 625
rect 3759 1236 3831 1292
rect 3759 1202 3778 1236
rect 3812 1202 3831 1236
rect 3759 1146 3831 1202
rect 3759 1112 3778 1146
rect 3812 1112 3831 1146
rect 3759 1056 3831 1112
rect 3759 1022 3778 1056
rect 3812 1022 3831 1056
rect 3759 966 3831 1022
rect 3759 932 3778 966
rect 3812 932 3831 966
rect 3759 876 3831 932
rect 3759 842 3778 876
rect 3812 842 3831 876
rect 3759 786 3831 842
rect 3759 752 3778 786
rect 3812 752 3831 786
rect 3759 696 3831 752
rect 3759 662 3778 696
rect 3812 662 3831 696
rect 3759 606 3831 662
rect 2869 531 2941 591
rect 3759 572 3778 606
rect 3812 572 3831 606
rect 3759 531 3831 572
rect 2869 512 3831 531
rect 2869 478 2966 512
rect 3000 478 3056 512
rect 3090 478 3146 512
rect 3180 478 3236 512
rect 3270 478 3326 512
rect 3360 478 3416 512
rect 3450 478 3506 512
rect 3540 478 3596 512
rect 3630 478 3686 512
rect 3720 478 3831 512
rect 2869 459 3831 478
rect 4209 1402 5171 1421
rect 4209 1368 4340 1402
rect 4374 1368 4430 1402
rect 4464 1368 4520 1402
rect 4554 1368 4610 1402
rect 4644 1368 4700 1402
rect 4734 1368 4790 1402
rect 4824 1368 4880 1402
rect 4914 1368 4970 1402
rect 5004 1368 5060 1402
rect 5094 1368 5171 1402
rect 4209 1349 5171 1368
rect 4209 1345 4281 1349
rect 4209 1311 4228 1345
rect 4262 1311 4281 1345
rect 4209 1255 4281 1311
rect 5099 1326 5171 1349
rect 5099 1292 5118 1326
rect 5152 1292 5171 1326
rect 4209 1221 4228 1255
rect 4262 1221 4281 1255
rect 4209 1165 4281 1221
rect 4209 1131 4228 1165
rect 4262 1131 4281 1165
rect 4209 1075 4281 1131
rect 4209 1041 4228 1075
rect 4262 1041 4281 1075
rect 4209 985 4281 1041
rect 4209 951 4228 985
rect 4262 951 4281 985
rect 4209 895 4281 951
rect 4209 861 4228 895
rect 4262 861 4281 895
rect 4209 805 4281 861
rect 4209 771 4228 805
rect 4262 771 4281 805
rect 4209 715 4281 771
rect 4209 681 4228 715
rect 4262 681 4281 715
rect 4209 625 4281 681
rect 4209 591 4228 625
rect 4262 591 4281 625
rect 5099 1236 5171 1292
rect 5099 1202 5118 1236
rect 5152 1202 5171 1236
rect 5099 1146 5171 1202
rect 5099 1112 5118 1146
rect 5152 1112 5171 1146
rect 5099 1056 5171 1112
rect 5099 1022 5118 1056
rect 5152 1022 5171 1056
rect 5099 966 5171 1022
rect 5099 932 5118 966
rect 5152 932 5171 966
rect 5099 876 5171 932
rect 5099 842 5118 876
rect 5152 842 5171 876
rect 5099 786 5171 842
rect 5099 752 5118 786
rect 5152 752 5171 786
rect 5099 696 5171 752
rect 5099 662 5118 696
rect 5152 662 5171 696
rect 5099 606 5171 662
rect 4209 531 4281 591
rect 5099 572 5118 606
rect 5152 572 5171 606
rect 5099 531 5171 572
rect 4209 512 5171 531
rect 4209 478 4306 512
rect 4340 478 4396 512
rect 4430 478 4486 512
rect 4520 478 4576 512
rect 4610 478 4666 512
rect 4700 478 4756 512
rect 4790 478 4846 512
rect 4880 478 4936 512
rect 4970 478 5026 512
rect 5060 478 5171 512
rect 4209 459 5171 478
rect 5549 1402 6511 1421
rect 5549 1368 5680 1402
rect 5714 1368 5770 1402
rect 5804 1368 5860 1402
rect 5894 1368 5950 1402
rect 5984 1368 6040 1402
rect 6074 1368 6130 1402
rect 6164 1368 6220 1402
rect 6254 1368 6310 1402
rect 6344 1368 6400 1402
rect 6434 1368 6511 1402
rect 5549 1349 6511 1368
rect 5549 1345 5621 1349
rect 5549 1311 5568 1345
rect 5602 1311 5621 1345
rect 5549 1255 5621 1311
rect 6439 1326 6511 1349
rect 6439 1292 6458 1326
rect 6492 1292 6511 1326
rect 5549 1221 5568 1255
rect 5602 1221 5621 1255
rect 5549 1165 5621 1221
rect 5549 1131 5568 1165
rect 5602 1131 5621 1165
rect 5549 1075 5621 1131
rect 5549 1041 5568 1075
rect 5602 1041 5621 1075
rect 5549 985 5621 1041
rect 5549 951 5568 985
rect 5602 951 5621 985
rect 5549 895 5621 951
rect 5549 861 5568 895
rect 5602 861 5621 895
rect 5549 805 5621 861
rect 5549 771 5568 805
rect 5602 771 5621 805
rect 5549 715 5621 771
rect 5549 681 5568 715
rect 5602 681 5621 715
rect 5549 625 5621 681
rect 5549 591 5568 625
rect 5602 591 5621 625
rect 6439 1236 6511 1292
rect 6439 1202 6458 1236
rect 6492 1202 6511 1236
rect 6439 1146 6511 1202
rect 6439 1112 6458 1146
rect 6492 1112 6511 1146
rect 6439 1056 6511 1112
rect 6439 1022 6458 1056
rect 6492 1022 6511 1056
rect 6439 966 6511 1022
rect 6439 932 6458 966
rect 6492 932 6511 966
rect 6439 876 6511 932
rect 6439 842 6458 876
rect 6492 842 6511 876
rect 6439 786 6511 842
rect 6439 752 6458 786
rect 6492 752 6511 786
rect 6439 696 6511 752
rect 6439 662 6458 696
rect 6492 662 6511 696
rect 6439 606 6511 662
rect 5549 531 5621 591
rect 6439 572 6458 606
rect 6492 572 6511 606
rect 6439 531 6511 572
rect 5549 512 6511 531
rect 5549 478 5646 512
rect 5680 478 5736 512
rect 5770 478 5826 512
rect 5860 478 5916 512
rect 5950 478 6006 512
rect 6040 478 6096 512
rect 6130 478 6186 512
rect 6220 478 6276 512
rect 6310 478 6366 512
rect 6400 478 6511 512
rect 5549 459 6511 478
rect 6889 1402 7851 1421
rect 6889 1368 7020 1402
rect 7054 1368 7110 1402
rect 7144 1368 7200 1402
rect 7234 1368 7290 1402
rect 7324 1368 7380 1402
rect 7414 1368 7470 1402
rect 7504 1368 7560 1402
rect 7594 1368 7650 1402
rect 7684 1368 7740 1402
rect 7774 1368 7851 1402
rect 6889 1349 7851 1368
rect 6889 1345 6961 1349
rect 6889 1311 6908 1345
rect 6942 1311 6961 1345
rect 6889 1255 6961 1311
rect 7779 1326 7851 1349
rect 7779 1292 7798 1326
rect 7832 1292 7851 1326
rect 6889 1221 6908 1255
rect 6942 1221 6961 1255
rect 6889 1165 6961 1221
rect 6889 1131 6908 1165
rect 6942 1131 6961 1165
rect 6889 1075 6961 1131
rect 6889 1041 6908 1075
rect 6942 1041 6961 1075
rect 6889 985 6961 1041
rect 6889 951 6908 985
rect 6942 951 6961 985
rect 6889 895 6961 951
rect 6889 861 6908 895
rect 6942 861 6961 895
rect 6889 805 6961 861
rect 6889 771 6908 805
rect 6942 771 6961 805
rect 6889 715 6961 771
rect 6889 681 6908 715
rect 6942 681 6961 715
rect 6889 625 6961 681
rect 6889 591 6908 625
rect 6942 591 6961 625
rect 7779 1236 7851 1292
rect 7779 1202 7798 1236
rect 7832 1202 7851 1236
rect 7779 1146 7851 1202
rect 7779 1112 7798 1146
rect 7832 1112 7851 1146
rect 7779 1056 7851 1112
rect 7779 1022 7798 1056
rect 7832 1022 7851 1056
rect 7779 966 7851 1022
rect 7779 932 7798 966
rect 7832 932 7851 966
rect 7779 876 7851 932
rect 7779 842 7798 876
rect 7832 842 7851 876
rect 7779 786 7851 842
rect 7779 752 7798 786
rect 7832 752 7851 786
rect 7779 696 7851 752
rect 7779 662 7798 696
rect 7832 662 7851 696
rect 7779 606 7851 662
rect 6889 531 6961 591
rect 7779 572 7798 606
rect 7832 572 7851 606
rect 7779 531 7851 572
rect 6889 512 7851 531
rect 6889 478 6986 512
rect 7020 478 7076 512
rect 7110 478 7166 512
rect 7200 478 7256 512
rect 7290 478 7346 512
rect 7380 478 7436 512
rect 7470 478 7526 512
rect 7560 478 7616 512
rect 7650 478 7706 512
rect 7740 478 7851 512
rect 6889 459 7851 478
rect 8229 1402 9191 1421
rect 8229 1368 8360 1402
rect 8394 1368 8450 1402
rect 8484 1368 8540 1402
rect 8574 1368 8630 1402
rect 8664 1368 8720 1402
rect 8754 1368 8810 1402
rect 8844 1368 8900 1402
rect 8934 1368 8990 1402
rect 9024 1368 9080 1402
rect 9114 1368 9191 1402
rect 8229 1349 9191 1368
rect 8229 1345 8301 1349
rect 8229 1311 8248 1345
rect 8282 1311 8301 1345
rect 8229 1255 8301 1311
rect 9119 1326 9191 1349
rect 9119 1292 9138 1326
rect 9172 1292 9191 1326
rect 8229 1221 8248 1255
rect 8282 1221 8301 1255
rect 8229 1165 8301 1221
rect 8229 1131 8248 1165
rect 8282 1131 8301 1165
rect 8229 1075 8301 1131
rect 8229 1041 8248 1075
rect 8282 1041 8301 1075
rect 8229 985 8301 1041
rect 8229 951 8248 985
rect 8282 951 8301 985
rect 8229 895 8301 951
rect 8229 861 8248 895
rect 8282 861 8301 895
rect 8229 805 8301 861
rect 8229 771 8248 805
rect 8282 771 8301 805
rect 8229 715 8301 771
rect 8229 681 8248 715
rect 8282 681 8301 715
rect 8229 625 8301 681
rect 8229 591 8248 625
rect 8282 591 8301 625
rect 9119 1236 9191 1292
rect 9119 1202 9138 1236
rect 9172 1202 9191 1236
rect 9119 1146 9191 1202
rect 9119 1112 9138 1146
rect 9172 1112 9191 1146
rect 9119 1056 9191 1112
rect 9119 1022 9138 1056
rect 9172 1022 9191 1056
rect 9119 966 9191 1022
rect 9119 932 9138 966
rect 9172 932 9191 966
rect 9119 876 9191 932
rect 9119 842 9138 876
rect 9172 842 9191 876
rect 9119 786 9191 842
rect 9119 752 9138 786
rect 9172 752 9191 786
rect 9119 696 9191 752
rect 9119 662 9138 696
rect 9172 662 9191 696
rect 9119 606 9191 662
rect 8229 531 8301 591
rect 9119 572 9138 606
rect 9172 572 9191 606
rect 9119 531 9191 572
rect 8229 512 9191 531
rect 8229 478 8326 512
rect 8360 478 8416 512
rect 8450 478 8506 512
rect 8540 478 8596 512
rect 8630 478 8686 512
rect 8720 478 8776 512
rect 8810 478 8866 512
rect 8900 478 8956 512
rect 8990 478 9046 512
rect 9080 478 9191 512
rect 8229 459 9191 478
<< psubdiffcont >>
rect 60 1492 94 1526
rect 156 1515 190 1549
rect 246 1515 280 1549
rect 336 1515 370 1549
rect 426 1515 460 1549
rect 516 1515 550 1549
rect 606 1515 640 1549
rect 696 1515 730 1549
rect 786 1515 820 1549
rect 876 1515 910 1549
rect 966 1515 1000 1549
rect 1056 1515 1090 1549
rect 1146 1515 1180 1549
rect 1247 1492 1281 1526
rect 1400 1492 1434 1526
rect 1496 1515 1530 1549
rect 1586 1515 1620 1549
rect 1676 1515 1710 1549
rect 1766 1515 1800 1549
rect 1856 1515 1890 1549
rect 1946 1515 1980 1549
rect 2036 1515 2070 1549
rect 2126 1515 2160 1549
rect 2216 1515 2250 1549
rect 2306 1515 2340 1549
rect 2396 1515 2430 1549
rect 2486 1515 2520 1549
rect 2587 1492 2621 1526
rect 2740 1492 2774 1526
rect 2836 1515 2870 1549
rect 2926 1515 2960 1549
rect 3016 1515 3050 1549
rect 3106 1515 3140 1549
rect 3196 1515 3230 1549
rect 3286 1515 3320 1549
rect 3376 1515 3410 1549
rect 3466 1515 3500 1549
rect 3556 1515 3590 1549
rect 3646 1515 3680 1549
rect 3736 1515 3770 1549
rect 3826 1515 3860 1549
rect 3927 1492 3961 1526
rect 4080 1492 4114 1526
rect 4176 1515 4210 1549
rect 4266 1515 4300 1549
rect 4356 1515 4390 1549
rect 4446 1515 4480 1549
rect 4536 1515 4570 1549
rect 4626 1515 4660 1549
rect 4716 1515 4750 1549
rect 4806 1515 4840 1549
rect 4896 1515 4930 1549
rect 4986 1515 5020 1549
rect 5076 1515 5110 1549
rect 5166 1515 5200 1549
rect 5267 1492 5301 1526
rect 5420 1492 5454 1526
rect 5516 1515 5550 1549
rect 5606 1515 5640 1549
rect 5696 1515 5730 1549
rect 5786 1515 5820 1549
rect 5876 1515 5910 1549
rect 5966 1515 6000 1549
rect 6056 1515 6090 1549
rect 6146 1515 6180 1549
rect 6236 1515 6270 1549
rect 6326 1515 6360 1549
rect 6416 1515 6450 1549
rect 6506 1515 6540 1549
rect 6607 1492 6641 1526
rect 6760 1492 6794 1526
rect 6856 1515 6890 1549
rect 6946 1515 6980 1549
rect 7036 1515 7070 1549
rect 7126 1515 7160 1549
rect 7216 1515 7250 1549
rect 7306 1515 7340 1549
rect 7396 1515 7430 1549
rect 7486 1515 7520 1549
rect 7576 1515 7610 1549
rect 7666 1515 7700 1549
rect 7756 1515 7790 1549
rect 7846 1515 7880 1549
rect 7947 1492 7981 1526
rect 8100 1492 8134 1526
rect 8196 1515 8230 1549
rect 8286 1515 8320 1549
rect 8376 1515 8410 1549
rect 8466 1515 8500 1549
rect 8556 1515 8590 1549
rect 8646 1515 8680 1549
rect 8736 1515 8770 1549
rect 8826 1515 8860 1549
rect 8916 1515 8950 1549
rect 9006 1515 9040 1549
rect 9096 1515 9130 1549
rect 9186 1515 9220 1549
rect 9287 1492 9321 1526
rect 60 1402 94 1436
rect 60 1312 94 1346
rect 60 1222 94 1256
rect 60 1132 94 1166
rect 60 1042 94 1076
rect 60 952 94 986
rect 60 862 94 896
rect 60 772 94 806
rect 60 682 94 716
rect 60 592 94 626
rect 60 502 94 536
rect 1247 1402 1281 1436
rect 1400 1402 1434 1436
rect 1247 1312 1281 1346
rect 1400 1312 1434 1346
rect 1247 1222 1281 1256
rect 1400 1222 1434 1256
rect 1247 1132 1281 1166
rect 1400 1132 1434 1166
rect 1247 1042 1281 1076
rect 1400 1042 1434 1076
rect 1247 952 1281 986
rect 1400 952 1434 986
rect 1247 862 1281 896
rect 1400 862 1434 896
rect 1247 772 1281 806
rect 1400 772 1434 806
rect 1247 682 1281 716
rect 1400 682 1434 716
rect 1247 592 1281 626
rect 1400 592 1434 626
rect 1247 502 1281 536
rect 1400 502 1434 536
rect 60 412 94 446
rect 2587 1402 2621 1436
rect 2740 1402 2774 1436
rect 2587 1312 2621 1346
rect 2740 1312 2774 1346
rect 2587 1222 2621 1256
rect 2740 1222 2774 1256
rect 2587 1132 2621 1166
rect 2740 1132 2774 1166
rect 2587 1042 2621 1076
rect 2740 1042 2774 1076
rect 2587 952 2621 986
rect 2740 952 2774 986
rect 2587 862 2621 896
rect 2740 862 2774 896
rect 2587 772 2621 806
rect 2740 772 2774 806
rect 2587 682 2621 716
rect 2740 682 2774 716
rect 2587 592 2621 626
rect 2740 592 2774 626
rect 2587 502 2621 536
rect 2740 502 2774 536
rect 1247 412 1281 446
rect 1400 412 1434 446
rect 3927 1402 3961 1436
rect 4080 1402 4114 1436
rect 3927 1312 3961 1346
rect 4080 1312 4114 1346
rect 3927 1222 3961 1256
rect 4080 1222 4114 1256
rect 3927 1132 3961 1166
rect 4080 1132 4114 1166
rect 3927 1042 3961 1076
rect 4080 1042 4114 1076
rect 3927 952 3961 986
rect 4080 952 4114 986
rect 3927 862 3961 896
rect 4080 862 4114 896
rect 3927 772 3961 806
rect 4080 772 4114 806
rect 3927 682 3961 716
rect 4080 682 4114 716
rect 3927 592 3961 626
rect 4080 592 4114 626
rect 3927 502 3961 536
rect 4080 502 4114 536
rect 2587 412 2621 446
rect 2740 412 2774 446
rect 5267 1402 5301 1436
rect 5420 1402 5454 1436
rect 5267 1312 5301 1346
rect 5420 1312 5454 1346
rect 5267 1222 5301 1256
rect 5420 1222 5454 1256
rect 5267 1132 5301 1166
rect 5420 1132 5454 1166
rect 5267 1042 5301 1076
rect 5420 1042 5454 1076
rect 5267 952 5301 986
rect 5420 952 5454 986
rect 5267 862 5301 896
rect 5420 862 5454 896
rect 5267 772 5301 806
rect 5420 772 5454 806
rect 5267 682 5301 716
rect 5420 682 5454 716
rect 5267 592 5301 626
rect 5420 592 5454 626
rect 5267 502 5301 536
rect 5420 502 5454 536
rect 3927 412 3961 446
rect 4080 412 4114 446
rect 6607 1402 6641 1436
rect 6760 1402 6794 1436
rect 6607 1312 6641 1346
rect 6760 1312 6794 1346
rect 6607 1222 6641 1256
rect 6760 1222 6794 1256
rect 6607 1132 6641 1166
rect 6760 1132 6794 1166
rect 6607 1042 6641 1076
rect 6760 1042 6794 1076
rect 6607 952 6641 986
rect 6760 952 6794 986
rect 6607 862 6641 896
rect 6760 862 6794 896
rect 6607 772 6641 806
rect 6760 772 6794 806
rect 6607 682 6641 716
rect 6760 682 6794 716
rect 6607 592 6641 626
rect 6760 592 6794 626
rect 6607 502 6641 536
rect 6760 502 6794 536
rect 5267 412 5301 446
rect 5420 412 5454 446
rect 7947 1402 7981 1436
rect 8100 1402 8134 1436
rect 7947 1312 7981 1346
rect 8100 1312 8134 1346
rect 7947 1222 7981 1256
rect 8100 1222 8134 1256
rect 7947 1132 7981 1166
rect 8100 1132 8134 1166
rect 7947 1042 7981 1076
rect 8100 1042 8134 1076
rect 7947 952 7981 986
rect 8100 952 8134 986
rect 7947 862 7981 896
rect 8100 862 8134 896
rect 7947 772 7981 806
rect 8100 772 8134 806
rect 7947 682 7981 716
rect 8100 682 8134 716
rect 7947 592 7981 626
rect 8100 592 8134 626
rect 7947 502 7981 536
rect 8100 502 8134 536
rect 6607 412 6641 446
rect 6760 412 6794 446
rect 9287 1402 9321 1436
rect 9287 1312 9321 1346
rect 9287 1222 9321 1256
rect 9287 1132 9321 1166
rect 9287 1042 9321 1076
rect 9287 952 9321 986
rect 9287 862 9321 896
rect 9287 772 9321 806
rect 9287 682 9321 716
rect 9287 592 9321 626
rect 9287 502 9321 536
rect 7947 412 7981 446
rect 8100 412 8134 446
rect 9287 412 9321 446
rect 156 328 190 362
rect 246 328 280 362
rect 336 328 370 362
rect 426 328 460 362
rect 516 328 550 362
rect 606 328 640 362
rect 696 328 730 362
rect 786 328 820 362
rect 876 328 910 362
rect 966 328 1000 362
rect 1056 328 1090 362
rect 1146 328 1180 362
rect 1496 328 1530 362
rect 1586 328 1620 362
rect 1676 328 1710 362
rect 1766 328 1800 362
rect 1856 328 1890 362
rect 1946 328 1980 362
rect 2036 328 2070 362
rect 2126 328 2160 362
rect 2216 328 2250 362
rect 2306 328 2340 362
rect 2396 328 2430 362
rect 2486 328 2520 362
rect 2836 328 2870 362
rect 2926 328 2960 362
rect 3016 328 3050 362
rect 3106 328 3140 362
rect 3196 328 3230 362
rect 3286 328 3320 362
rect 3376 328 3410 362
rect 3466 328 3500 362
rect 3556 328 3590 362
rect 3646 328 3680 362
rect 3736 328 3770 362
rect 3826 328 3860 362
rect 4176 328 4210 362
rect 4266 328 4300 362
rect 4356 328 4390 362
rect 4446 328 4480 362
rect 4536 328 4570 362
rect 4626 328 4660 362
rect 4716 328 4750 362
rect 4806 328 4840 362
rect 4896 328 4930 362
rect 4986 328 5020 362
rect 5076 328 5110 362
rect 5166 328 5200 362
rect 5516 328 5550 362
rect 5606 328 5640 362
rect 5696 328 5730 362
rect 5786 328 5820 362
rect 5876 328 5910 362
rect 5966 328 6000 362
rect 6056 328 6090 362
rect 6146 328 6180 362
rect 6236 328 6270 362
rect 6326 328 6360 362
rect 6416 328 6450 362
rect 6506 328 6540 362
rect 6856 328 6890 362
rect 6946 328 6980 362
rect 7036 328 7070 362
rect 7126 328 7160 362
rect 7216 328 7250 362
rect 7306 328 7340 362
rect 7396 328 7430 362
rect 7486 328 7520 362
rect 7576 328 7610 362
rect 7666 328 7700 362
rect 7756 328 7790 362
rect 7846 328 7880 362
rect 8196 328 8230 362
rect 8286 328 8320 362
rect 8376 328 8410 362
rect 8466 328 8500 362
rect 8556 328 8590 362
rect 8646 328 8680 362
rect 8736 328 8770 362
rect 8826 328 8860 362
rect 8916 328 8950 362
rect 9006 328 9040 362
rect 9096 328 9130 362
rect 9186 328 9220 362
<< nsubdiffcont >>
rect 320 1368 354 1402
rect 410 1368 444 1402
rect 500 1368 534 1402
rect 590 1368 624 1402
rect 680 1368 714 1402
rect 770 1368 804 1402
rect 860 1368 894 1402
rect 950 1368 984 1402
rect 1040 1368 1074 1402
rect 208 1311 242 1345
rect 1098 1292 1132 1326
rect 208 1221 242 1255
rect 208 1131 242 1165
rect 208 1041 242 1075
rect 208 951 242 985
rect 208 861 242 895
rect 208 771 242 805
rect 208 681 242 715
rect 208 591 242 625
rect 1098 1202 1132 1236
rect 1098 1112 1132 1146
rect 1098 1022 1132 1056
rect 1098 932 1132 966
rect 1098 842 1132 876
rect 1098 752 1132 786
rect 1098 662 1132 696
rect 1098 572 1132 606
rect 286 478 320 512
rect 376 478 410 512
rect 466 478 500 512
rect 556 478 590 512
rect 646 478 680 512
rect 736 478 770 512
rect 826 478 860 512
rect 916 478 950 512
rect 1006 478 1040 512
rect 1660 1368 1694 1402
rect 1750 1368 1784 1402
rect 1840 1368 1874 1402
rect 1930 1368 1964 1402
rect 2020 1368 2054 1402
rect 2110 1368 2144 1402
rect 2200 1368 2234 1402
rect 2290 1368 2324 1402
rect 2380 1368 2414 1402
rect 1548 1311 1582 1345
rect 2438 1292 2472 1326
rect 1548 1221 1582 1255
rect 1548 1131 1582 1165
rect 1548 1041 1582 1075
rect 1548 951 1582 985
rect 1548 861 1582 895
rect 1548 771 1582 805
rect 1548 681 1582 715
rect 1548 591 1582 625
rect 2438 1202 2472 1236
rect 2438 1112 2472 1146
rect 2438 1022 2472 1056
rect 2438 932 2472 966
rect 2438 842 2472 876
rect 2438 752 2472 786
rect 2438 662 2472 696
rect 2438 572 2472 606
rect 1626 478 1660 512
rect 1716 478 1750 512
rect 1806 478 1840 512
rect 1896 478 1930 512
rect 1986 478 2020 512
rect 2076 478 2110 512
rect 2166 478 2200 512
rect 2256 478 2290 512
rect 2346 478 2380 512
rect 3000 1368 3034 1402
rect 3090 1368 3124 1402
rect 3180 1368 3214 1402
rect 3270 1368 3304 1402
rect 3360 1368 3394 1402
rect 3450 1368 3484 1402
rect 3540 1368 3574 1402
rect 3630 1368 3664 1402
rect 3720 1368 3754 1402
rect 2888 1311 2922 1345
rect 3778 1292 3812 1326
rect 2888 1221 2922 1255
rect 2888 1131 2922 1165
rect 2888 1041 2922 1075
rect 2888 951 2922 985
rect 2888 861 2922 895
rect 2888 771 2922 805
rect 2888 681 2922 715
rect 2888 591 2922 625
rect 3778 1202 3812 1236
rect 3778 1112 3812 1146
rect 3778 1022 3812 1056
rect 3778 932 3812 966
rect 3778 842 3812 876
rect 3778 752 3812 786
rect 3778 662 3812 696
rect 3778 572 3812 606
rect 2966 478 3000 512
rect 3056 478 3090 512
rect 3146 478 3180 512
rect 3236 478 3270 512
rect 3326 478 3360 512
rect 3416 478 3450 512
rect 3506 478 3540 512
rect 3596 478 3630 512
rect 3686 478 3720 512
rect 4340 1368 4374 1402
rect 4430 1368 4464 1402
rect 4520 1368 4554 1402
rect 4610 1368 4644 1402
rect 4700 1368 4734 1402
rect 4790 1368 4824 1402
rect 4880 1368 4914 1402
rect 4970 1368 5004 1402
rect 5060 1368 5094 1402
rect 4228 1311 4262 1345
rect 5118 1292 5152 1326
rect 4228 1221 4262 1255
rect 4228 1131 4262 1165
rect 4228 1041 4262 1075
rect 4228 951 4262 985
rect 4228 861 4262 895
rect 4228 771 4262 805
rect 4228 681 4262 715
rect 4228 591 4262 625
rect 5118 1202 5152 1236
rect 5118 1112 5152 1146
rect 5118 1022 5152 1056
rect 5118 932 5152 966
rect 5118 842 5152 876
rect 5118 752 5152 786
rect 5118 662 5152 696
rect 5118 572 5152 606
rect 4306 478 4340 512
rect 4396 478 4430 512
rect 4486 478 4520 512
rect 4576 478 4610 512
rect 4666 478 4700 512
rect 4756 478 4790 512
rect 4846 478 4880 512
rect 4936 478 4970 512
rect 5026 478 5060 512
rect 5680 1368 5714 1402
rect 5770 1368 5804 1402
rect 5860 1368 5894 1402
rect 5950 1368 5984 1402
rect 6040 1368 6074 1402
rect 6130 1368 6164 1402
rect 6220 1368 6254 1402
rect 6310 1368 6344 1402
rect 6400 1368 6434 1402
rect 5568 1311 5602 1345
rect 6458 1292 6492 1326
rect 5568 1221 5602 1255
rect 5568 1131 5602 1165
rect 5568 1041 5602 1075
rect 5568 951 5602 985
rect 5568 861 5602 895
rect 5568 771 5602 805
rect 5568 681 5602 715
rect 5568 591 5602 625
rect 6458 1202 6492 1236
rect 6458 1112 6492 1146
rect 6458 1022 6492 1056
rect 6458 932 6492 966
rect 6458 842 6492 876
rect 6458 752 6492 786
rect 6458 662 6492 696
rect 6458 572 6492 606
rect 5646 478 5680 512
rect 5736 478 5770 512
rect 5826 478 5860 512
rect 5916 478 5950 512
rect 6006 478 6040 512
rect 6096 478 6130 512
rect 6186 478 6220 512
rect 6276 478 6310 512
rect 6366 478 6400 512
rect 7020 1368 7054 1402
rect 7110 1368 7144 1402
rect 7200 1368 7234 1402
rect 7290 1368 7324 1402
rect 7380 1368 7414 1402
rect 7470 1368 7504 1402
rect 7560 1368 7594 1402
rect 7650 1368 7684 1402
rect 7740 1368 7774 1402
rect 6908 1311 6942 1345
rect 7798 1292 7832 1326
rect 6908 1221 6942 1255
rect 6908 1131 6942 1165
rect 6908 1041 6942 1075
rect 6908 951 6942 985
rect 6908 861 6942 895
rect 6908 771 6942 805
rect 6908 681 6942 715
rect 6908 591 6942 625
rect 7798 1202 7832 1236
rect 7798 1112 7832 1146
rect 7798 1022 7832 1056
rect 7798 932 7832 966
rect 7798 842 7832 876
rect 7798 752 7832 786
rect 7798 662 7832 696
rect 7798 572 7832 606
rect 6986 478 7020 512
rect 7076 478 7110 512
rect 7166 478 7200 512
rect 7256 478 7290 512
rect 7346 478 7380 512
rect 7436 478 7470 512
rect 7526 478 7560 512
rect 7616 478 7650 512
rect 7706 478 7740 512
rect 8360 1368 8394 1402
rect 8450 1368 8484 1402
rect 8540 1368 8574 1402
rect 8630 1368 8664 1402
rect 8720 1368 8754 1402
rect 8810 1368 8844 1402
rect 8900 1368 8934 1402
rect 8990 1368 9024 1402
rect 9080 1368 9114 1402
rect 8248 1311 8282 1345
rect 9138 1292 9172 1326
rect 8248 1221 8282 1255
rect 8248 1131 8282 1165
rect 8248 1041 8282 1075
rect 8248 951 8282 985
rect 8248 861 8282 895
rect 8248 771 8282 805
rect 8248 681 8282 715
rect 8248 591 8282 625
rect 9138 1202 9172 1236
rect 9138 1112 9172 1146
rect 9138 1022 9172 1056
rect 9138 932 9172 966
rect 9138 842 9172 876
rect 9138 752 9172 786
rect 9138 662 9172 696
rect 9138 572 9172 606
rect 8326 478 8360 512
rect 8416 478 8450 512
rect 8506 478 8540 512
rect 8596 478 8630 512
rect 8686 478 8720 512
rect 8776 478 8810 512
rect 8866 478 8900 512
rect 8956 478 8990 512
rect 9046 478 9080 512
<< locali >>
rect 0 1850 170 1910
rect 230 1850 370 1910
rect 430 1850 570 1910
rect 630 1850 770 1910
rect 830 1850 970 1910
rect 1030 1850 1170 1910
rect 1230 1850 1370 1910
rect 1430 1850 1570 1910
rect 1630 1850 1770 1910
rect 1830 1850 1970 1910
rect 2030 1850 2170 1910
rect 2230 1850 2370 1910
rect 2430 1850 2570 1910
rect 2630 1850 2770 1910
rect 2830 1850 2970 1910
rect 3030 1850 3170 1910
rect 3230 1850 3370 1910
rect 3430 1850 3570 1910
rect 3630 1850 3770 1910
rect 3830 1850 3970 1910
rect 4030 1850 4170 1910
rect 4230 1850 4370 1910
rect 4430 1850 4570 1910
rect 4630 1850 4770 1910
rect 4830 1850 4970 1910
rect 5030 1850 5170 1910
rect 5230 1850 5370 1910
rect 5430 1850 5570 1910
rect 5630 1850 5770 1910
rect 5830 1850 5970 1910
rect 6030 1850 6170 1910
rect 6230 1850 6370 1910
rect 6430 1850 6570 1910
rect 6630 1850 6770 1910
rect 6830 1850 6970 1910
rect 7030 1850 7170 1910
rect 7230 1850 7370 1910
rect 7430 1850 7570 1910
rect 7630 1850 7770 1910
rect 7830 1850 7970 1910
rect 8030 1850 8170 1910
rect 8230 1850 8370 1910
rect 8430 1850 8570 1910
rect 8630 1850 8770 1910
rect 8830 1850 8970 1910
rect 9030 1850 9170 1910
rect 9230 1850 9380 1910
rect 26 1549 9357 1584
rect 26 1526 156 1549
rect 26 1492 60 1526
rect 94 1515 156 1526
rect 190 1515 246 1549
rect 280 1515 336 1549
rect 370 1515 426 1549
rect 460 1515 516 1549
rect 550 1515 606 1549
rect 640 1515 696 1549
rect 730 1515 786 1549
rect 820 1515 876 1549
rect 910 1515 966 1549
rect 1000 1515 1056 1549
rect 1090 1515 1146 1549
rect 1180 1526 1496 1549
rect 1180 1515 1247 1526
rect 94 1492 1247 1515
rect 1281 1492 1400 1526
rect 1434 1515 1496 1526
rect 1530 1515 1586 1549
rect 1620 1515 1676 1549
rect 1710 1515 1766 1549
rect 1800 1515 1856 1549
rect 1890 1515 1946 1549
rect 1980 1515 2036 1549
rect 2070 1515 2126 1549
rect 2160 1515 2216 1549
rect 2250 1515 2306 1549
rect 2340 1515 2396 1549
rect 2430 1515 2486 1549
rect 2520 1526 2836 1549
rect 2520 1515 2587 1526
rect 1434 1492 2587 1515
rect 2621 1492 2740 1526
rect 2774 1515 2836 1526
rect 2870 1515 2926 1549
rect 2960 1515 3016 1549
rect 3050 1515 3106 1549
rect 3140 1515 3196 1549
rect 3230 1515 3286 1549
rect 3320 1515 3376 1549
rect 3410 1515 3466 1549
rect 3500 1515 3556 1549
rect 3590 1515 3646 1549
rect 3680 1515 3736 1549
rect 3770 1515 3826 1549
rect 3860 1526 4176 1549
rect 3860 1515 3927 1526
rect 2774 1492 3927 1515
rect 3961 1492 4080 1526
rect 4114 1515 4176 1526
rect 4210 1515 4266 1549
rect 4300 1515 4356 1549
rect 4390 1515 4446 1549
rect 4480 1515 4536 1549
rect 4570 1515 4626 1549
rect 4660 1515 4716 1549
rect 4750 1515 4806 1549
rect 4840 1515 4896 1549
rect 4930 1515 4986 1549
rect 5020 1515 5076 1549
rect 5110 1515 5166 1549
rect 5200 1526 5516 1549
rect 5200 1515 5267 1526
rect 4114 1492 5267 1515
rect 5301 1492 5420 1526
rect 5454 1515 5516 1526
rect 5550 1515 5606 1549
rect 5640 1515 5696 1549
rect 5730 1515 5786 1549
rect 5820 1515 5876 1549
rect 5910 1515 5966 1549
rect 6000 1515 6056 1549
rect 6090 1515 6146 1549
rect 6180 1515 6236 1549
rect 6270 1515 6326 1549
rect 6360 1515 6416 1549
rect 6450 1515 6506 1549
rect 6540 1526 6856 1549
rect 6540 1515 6607 1526
rect 5454 1492 6607 1515
rect 6641 1492 6760 1526
rect 6794 1515 6856 1526
rect 6890 1515 6946 1549
rect 6980 1515 7036 1549
rect 7070 1515 7126 1549
rect 7160 1515 7216 1549
rect 7250 1515 7306 1549
rect 7340 1515 7396 1549
rect 7430 1515 7486 1549
rect 7520 1515 7576 1549
rect 7610 1515 7666 1549
rect 7700 1515 7756 1549
rect 7790 1515 7846 1549
rect 7880 1526 8196 1549
rect 7880 1515 7947 1526
rect 6794 1492 7947 1515
rect 7981 1492 8100 1526
rect 8134 1515 8196 1526
rect 8230 1515 8286 1549
rect 8320 1515 8376 1549
rect 8410 1515 8466 1549
rect 8500 1515 8556 1549
rect 8590 1515 8646 1549
rect 8680 1515 8736 1549
rect 8770 1515 8826 1549
rect 8860 1515 8916 1549
rect 8950 1515 9006 1549
rect 9040 1515 9096 1549
rect 9130 1515 9186 1549
rect 9220 1526 9357 1549
rect 9220 1515 9287 1526
rect 8134 1492 9287 1515
rect 9321 1492 9357 1526
rect 26 1436 9357 1492
rect 26 1402 60 1436
rect 94 1410 1247 1436
rect 94 1402 125 1410
rect 26 1346 125 1402
rect 26 1312 60 1346
rect 94 1312 125 1346
rect 26 1256 125 1312
rect 26 1222 60 1256
rect 94 1222 125 1256
rect 26 1166 125 1222
rect 26 1132 60 1166
rect 94 1132 125 1166
rect 26 1076 125 1132
rect 26 1042 60 1076
rect 94 1042 125 1076
rect 26 986 125 1042
rect 26 952 60 986
rect 94 952 125 986
rect 26 896 125 952
rect 26 862 60 896
rect 94 862 125 896
rect 26 806 125 862
rect 26 772 60 806
rect 94 772 125 806
rect 26 716 125 772
rect 26 682 60 716
rect 94 682 125 716
rect 26 626 125 682
rect 26 592 60 626
rect 94 592 125 626
rect 26 536 125 592
rect 26 502 60 536
rect 94 502 125 536
rect 26 470 125 502
rect 189 1402 1151 1410
rect 189 1368 320 1402
rect 354 1368 410 1402
rect 444 1368 500 1402
rect 534 1368 590 1402
rect 624 1368 680 1402
rect 714 1368 770 1402
rect 804 1368 860 1402
rect 894 1368 950 1402
rect 984 1368 1040 1402
rect 1074 1368 1151 1402
rect 189 1349 1151 1368
rect 189 1345 261 1349
rect 189 1311 208 1345
rect 242 1311 261 1345
rect 189 1255 261 1311
rect 1079 1326 1151 1349
rect 1079 1292 1098 1326
rect 1132 1292 1151 1326
rect 189 1221 208 1255
rect 242 1221 261 1255
rect 189 1165 261 1221
rect 189 1131 208 1165
rect 242 1131 261 1165
rect 189 1075 261 1131
rect 189 1041 208 1075
rect 242 1041 261 1075
rect 189 985 261 1041
rect 189 951 208 985
rect 242 951 261 985
rect 189 895 261 951
rect 189 861 208 895
rect 242 861 261 895
rect 189 805 261 861
rect 189 771 208 805
rect 242 771 261 805
rect 189 715 261 771
rect 189 681 208 715
rect 242 681 261 715
rect 189 625 261 681
rect 189 591 208 625
rect 242 591 261 625
rect 323 1228 1017 1287
rect 323 1194 384 1228
rect 418 1200 474 1228
rect 508 1200 564 1228
rect 598 1200 654 1228
rect 430 1194 474 1200
rect 530 1194 564 1200
rect 630 1194 654 1200
rect 688 1200 744 1228
rect 688 1194 696 1200
rect 323 1166 396 1194
rect 430 1166 496 1194
rect 530 1166 596 1194
rect 630 1166 696 1194
rect 730 1194 744 1200
rect 778 1200 834 1228
rect 778 1194 796 1200
rect 730 1166 796 1194
rect 830 1194 834 1200
rect 868 1200 924 1228
rect 868 1194 896 1200
rect 958 1194 1017 1228
rect 830 1166 896 1194
rect 930 1166 1017 1194
rect 323 1138 1017 1166
rect 323 1104 384 1138
rect 418 1104 474 1138
rect 508 1104 564 1138
rect 598 1104 654 1138
rect 688 1104 744 1138
rect 778 1104 834 1138
rect 868 1104 924 1138
rect 958 1104 1017 1138
rect 323 1100 1017 1104
rect 323 1066 396 1100
rect 430 1066 496 1100
rect 530 1066 596 1100
rect 630 1066 696 1100
rect 730 1066 796 1100
rect 830 1066 896 1100
rect 930 1066 1017 1100
rect 323 1048 1017 1066
rect 323 1014 384 1048
rect 418 1014 474 1048
rect 508 1014 564 1048
rect 598 1014 654 1048
rect 688 1014 744 1048
rect 778 1014 834 1048
rect 868 1014 924 1048
rect 958 1014 1017 1048
rect 323 1000 1017 1014
rect 323 966 396 1000
rect 430 966 496 1000
rect 530 966 596 1000
rect 630 966 696 1000
rect 730 966 796 1000
rect 830 966 896 1000
rect 930 966 1017 1000
rect 323 958 1017 966
rect 323 924 384 958
rect 418 924 474 958
rect 508 924 564 958
rect 598 924 654 958
rect 688 924 744 958
rect 778 924 834 958
rect 868 924 924 958
rect 958 924 1017 958
rect 323 900 1017 924
rect 323 868 396 900
rect 430 868 496 900
rect 530 868 596 900
rect 630 868 696 900
rect 323 834 384 868
rect 430 866 474 868
rect 530 866 564 868
rect 630 866 654 868
rect 418 834 474 866
rect 508 834 564 866
rect 598 834 654 866
rect 688 866 696 868
rect 730 868 796 900
rect 730 866 744 868
rect 688 834 744 866
rect 778 866 796 868
rect 830 868 896 900
rect 930 868 1017 900
rect 830 866 834 868
rect 778 834 834 866
rect 868 866 896 868
rect 868 834 924 866
rect 958 834 1017 868
rect 323 800 1017 834
rect 323 778 396 800
rect 430 778 496 800
rect 530 778 596 800
rect 630 778 696 800
rect 323 744 384 778
rect 430 766 474 778
rect 530 766 564 778
rect 630 766 654 778
rect 418 744 474 766
rect 508 744 564 766
rect 598 744 654 766
rect 688 766 696 778
rect 730 778 796 800
rect 730 766 744 778
rect 688 744 744 766
rect 778 766 796 778
rect 830 778 896 800
rect 930 778 1017 800
rect 830 766 834 778
rect 778 744 834 766
rect 868 766 896 778
rect 868 744 924 766
rect 958 744 1017 778
rect 323 700 1017 744
rect 323 688 396 700
rect 430 688 496 700
rect 530 688 596 700
rect 630 688 696 700
rect 323 654 384 688
rect 430 666 474 688
rect 530 666 564 688
rect 630 666 654 688
rect 418 654 474 666
rect 508 654 564 666
rect 598 654 654 666
rect 688 666 696 688
rect 730 688 796 700
rect 730 666 744 688
rect 688 654 744 666
rect 778 666 796 688
rect 830 688 896 700
rect 930 688 1017 700
rect 830 666 834 688
rect 778 654 834 666
rect 868 666 896 688
rect 868 654 924 666
rect 958 654 1017 688
rect 323 593 1017 654
rect 1079 1236 1151 1292
rect 1079 1202 1098 1236
rect 1132 1202 1151 1236
rect 1079 1146 1151 1202
rect 1079 1112 1098 1146
rect 1132 1112 1151 1146
rect 1079 1056 1151 1112
rect 1079 1022 1098 1056
rect 1132 1022 1151 1056
rect 1079 966 1151 1022
rect 1079 932 1098 966
rect 1132 932 1151 966
rect 1079 876 1151 932
rect 1079 842 1098 876
rect 1132 842 1151 876
rect 1079 786 1151 842
rect 1079 752 1098 786
rect 1132 752 1151 786
rect 1079 696 1151 752
rect 1079 662 1098 696
rect 1132 662 1151 696
rect 1079 606 1151 662
rect 189 531 261 591
rect 1079 572 1098 606
rect 1132 572 1151 606
rect 1079 531 1151 572
rect 189 512 1151 531
rect 189 478 286 512
rect 320 478 376 512
rect 410 478 466 512
rect 500 478 556 512
rect 590 478 646 512
rect 680 478 736 512
rect 770 478 826 512
rect 860 478 916 512
rect 950 478 1006 512
rect 1040 478 1151 512
rect 189 470 1151 478
rect 1215 1402 1247 1410
rect 1281 1402 1400 1436
rect 1434 1410 2587 1436
rect 1434 1402 1465 1410
rect 1215 1346 1465 1402
rect 1215 1312 1247 1346
rect 1281 1312 1400 1346
rect 1434 1312 1465 1346
rect 1215 1256 1465 1312
rect 1215 1222 1247 1256
rect 1281 1222 1400 1256
rect 1434 1222 1465 1256
rect 1215 1166 1465 1222
rect 1215 1132 1247 1166
rect 1281 1132 1400 1166
rect 1434 1132 1465 1166
rect 1215 1076 1465 1132
rect 1215 1042 1247 1076
rect 1281 1042 1400 1076
rect 1434 1042 1465 1076
rect 1215 986 1465 1042
rect 1215 952 1247 986
rect 1281 952 1400 986
rect 1434 952 1465 986
rect 1215 896 1465 952
rect 1215 862 1247 896
rect 1281 862 1400 896
rect 1434 862 1465 896
rect 1215 806 1465 862
rect 1215 772 1247 806
rect 1281 772 1400 806
rect 1434 772 1465 806
rect 1215 716 1465 772
rect 1215 682 1247 716
rect 1281 682 1400 716
rect 1434 682 1465 716
rect 1215 626 1465 682
rect 1215 592 1247 626
rect 1281 592 1400 626
rect 1434 592 1465 626
rect 1215 536 1465 592
rect 1215 502 1247 536
rect 1281 502 1400 536
rect 1434 502 1465 536
rect 1215 470 1465 502
rect 1529 1402 2491 1410
rect 1529 1368 1660 1402
rect 1694 1368 1750 1402
rect 1784 1368 1840 1402
rect 1874 1368 1930 1402
rect 1964 1368 2020 1402
rect 2054 1368 2110 1402
rect 2144 1368 2200 1402
rect 2234 1368 2290 1402
rect 2324 1368 2380 1402
rect 2414 1368 2491 1402
rect 1529 1349 2491 1368
rect 1529 1345 1601 1349
rect 1529 1311 1548 1345
rect 1582 1311 1601 1345
rect 1529 1255 1601 1311
rect 2419 1326 2491 1349
rect 2419 1292 2438 1326
rect 2472 1292 2491 1326
rect 1529 1221 1548 1255
rect 1582 1221 1601 1255
rect 1529 1165 1601 1221
rect 1529 1131 1548 1165
rect 1582 1131 1601 1165
rect 1529 1075 1601 1131
rect 1529 1041 1548 1075
rect 1582 1041 1601 1075
rect 1529 985 1601 1041
rect 1529 951 1548 985
rect 1582 951 1601 985
rect 1529 895 1601 951
rect 1529 861 1548 895
rect 1582 861 1601 895
rect 1529 805 1601 861
rect 1529 771 1548 805
rect 1582 771 1601 805
rect 1529 715 1601 771
rect 1529 681 1548 715
rect 1582 681 1601 715
rect 1529 625 1601 681
rect 1529 591 1548 625
rect 1582 591 1601 625
rect 1663 1228 2357 1287
rect 1663 1194 1724 1228
rect 1758 1200 1814 1228
rect 1848 1200 1904 1228
rect 1938 1200 1994 1228
rect 1770 1194 1814 1200
rect 1870 1194 1904 1200
rect 1970 1194 1994 1200
rect 2028 1200 2084 1228
rect 2028 1194 2036 1200
rect 1663 1166 1736 1194
rect 1770 1166 1836 1194
rect 1870 1166 1936 1194
rect 1970 1166 2036 1194
rect 2070 1194 2084 1200
rect 2118 1200 2174 1228
rect 2118 1194 2136 1200
rect 2070 1166 2136 1194
rect 2170 1194 2174 1200
rect 2208 1200 2264 1228
rect 2208 1194 2236 1200
rect 2298 1194 2357 1228
rect 2170 1166 2236 1194
rect 2270 1166 2357 1194
rect 1663 1138 2357 1166
rect 1663 1104 1724 1138
rect 1758 1104 1814 1138
rect 1848 1104 1904 1138
rect 1938 1104 1994 1138
rect 2028 1104 2084 1138
rect 2118 1104 2174 1138
rect 2208 1104 2264 1138
rect 2298 1104 2357 1138
rect 1663 1100 2357 1104
rect 1663 1066 1736 1100
rect 1770 1066 1836 1100
rect 1870 1066 1936 1100
rect 1970 1066 2036 1100
rect 2070 1066 2136 1100
rect 2170 1066 2236 1100
rect 2270 1066 2357 1100
rect 1663 1048 2357 1066
rect 1663 1014 1724 1048
rect 1758 1014 1814 1048
rect 1848 1014 1904 1048
rect 1938 1014 1994 1048
rect 2028 1014 2084 1048
rect 2118 1014 2174 1048
rect 2208 1014 2264 1048
rect 2298 1014 2357 1048
rect 1663 1000 2357 1014
rect 1663 966 1736 1000
rect 1770 966 1836 1000
rect 1870 966 1936 1000
rect 1970 966 2036 1000
rect 2070 966 2136 1000
rect 2170 966 2236 1000
rect 2270 966 2357 1000
rect 1663 958 2357 966
rect 1663 924 1724 958
rect 1758 924 1814 958
rect 1848 924 1904 958
rect 1938 924 1994 958
rect 2028 924 2084 958
rect 2118 924 2174 958
rect 2208 924 2264 958
rect 2298 924 2357 958
rect 1663 900 2357 924
rect 1663 868 1736 900
rect 1770 868 1836 900
rect 1870 868 1936 900
rect 1970 868 2036 900
rect 1663 834 1724 868
rect 1770 866 1814 868
rect 1870 866 1904 868
rect 1970 866 1994 868
rect 1758 834 1814 866
rect 1848 834 1904 866
rect 1938 834 1994 866
rect 2028 866 2036 868
rect 2070 868 2136 900
rect 2070 866 2084 868
rect 2028 834 2084 866
rect 2118 866 2136 868
rect 2170 868 2236 900
rect 2270 868 2357 900
rect 2170 866 2174 868
rect 2118 834 2174 866
rect 2208 866 2236 868
rect 2208 834 2264 866
rect 2298 834 2357 868
rect 1663 800 2357 834
rect 1663 778 1736 800
rect 1770 778 1836 800
rect 1870 778 1936 800
rect 1970 778 2036 800
rect 1663 744 1724 778
rect 1770 766 1814 778
rect 1870 766 1904 778
rect 1970 766 1994 778
rect 1758 744 1814 766
rect 1848 744 1904 766
rect 1938 744 1994 766
rect 2028 766 2036 778
rect 2070 778 2136 800
rect 2070 766 2084 778
rect 2028 744 2084 766
rect 2118 766 2136 778
rect 2170 778 2236 800
rect 2270 778 2357 800
rect 2170 766 2174 778
rect 2118 744 2174 766
rect 2208 766 2236 778
rect 2208 744 2264 766
rect 2298 744 2357 778
rect 1663 700 2357 744
rect 1663 688 1736 700
rect 1770 688 1836 700
rect 1870 688 1936 700
rect 1970 688 2036 700
rect 1663 654 1724 688
rect 1770 666 1814 688
rect 1870 666 1904 688
rect 1970 666 1994 688
rect 1758 654 1814 666
rect 1848 654 1904 666
rect 1938 654 1994 666
rect 2028 666 2036 688
rect 2070 688 2136 700
rect 2070 666 2084 688
rect 2028 654 2084 666
rect 2118 666 2136 688
rect 2170 688 2236 700
rect 2270 688 2357 700
rect 2170 666 2174 688
rect 2118 654 2174 666
rect 2208 666 2236 688
rect 2208 654 2264 666
rect 2298 654 2357 688
rect 1663 593 2357 654
rect 2419 1236 2491 1292
rect 2419 1202 2438 1236
rect 2472 1202 2491 1236
rect 2419 1146 2491 1202
rect 2419 1112 2438 1146
rect 2472 1112 2491 1146
rect 2419 1056 2491 1112
rect 2419 1022 2438 1056
rect 2472 1022 2491 1056
rect 2419 966 2491 1022
rect 2419 932 2438 966
rect 2472 932 2491 966
rect 2419 876 2491 932
rect 2419 842 2438 876
rect 2472 842 2491 876
rect 2419 786 2491 842
rect 2419 752 2438 786
rect 2472 752 2491 786
rect 2419 696 2491 752
rect 2419 662 2438 696
rect 2472 662 2491 696
rect 2419 606 2491 662
rect 1529 531 1601 591
rect 2419 572 2438 606
rect 2472 572 2491 606
rect 2419 531 2491 572
rect 1529 512 2491 531
rect 1529 478 1626 512
rect 1660 478 1716 512
rect 1750 478 1806 512
rect 1840 478 1896 512
rect 1930 478 1986 512
rect 2020 478 2076 512
rect 2110 478 2166 512
rect 2200 478 2256 512
rect 2290 478 2346 512
rect 2380 478 2491 512
rect 1529 470 2491 478
rect 2555 1402 2587 1410
rect 2621 1402 2740 1436
rect 2774 1410 3927 1436
rect 2774 1402 2805 1410
rect 2555 1346 2805 1402
rect 2555 1312 2587 1346
rect 2621 1312 2740 1346
rect 2774 1312 2805 1346
rect 2555 1256 2805 1312
rect 2555 1222 2587 1256
rect 2621 1222 2740 1256
rect 2774 1222 2805 1256
rect 2555 1166 2805 1222
rect 2555 1132 2587 1166
rect 2621 1132 2740 1166
rect 2774 1132 2805 1166
rect 2555 1076 2805 1132
rect 2555 1042 2587 1076
rect 2621 1042 2740 1076
rect 2774 1042 2805 1076
rect 2555 986 2805 1042
rect 2555 952 2587 986
rect 2621 952 2740 986
rect 2774 952 2805 986
rect 2555 896 2805 952
rect 2555 862 2587 896
rect 2621 862 2740 896
rect 2774 862 2805 896
rect 2555 806 2805 862
rect 2555 772 2587 806
rect 2621 772 2740 806
rect 2774 772 2805 806
rect 2555 716 2805 772
rect 2555 682 2587 716
rect 2621 682 2740 716
rect 2774 682 2805 716
rect 2555 626 2805 682
rect 2555 592 2587 626
rect 2621 592 2740 626
rect 2774 592 2805 626
rect 2555 536 2805 592
rect 2555 502 2587 536
rect 2621 502 2740 536
rect 2774 502 2805 536
rect 2555 470 2805 502
rect 2869 1402 3831 1410
rect 2869 1368 3000 1402
rect 3034 1368 3090 1402
rect 3124 1368 3180 1402
rect 3214 1368 3270 1402
rect 3304 1368 3360 1402
rect 3394 1368 3450 1402
rect 3484 1368 3540 1402
rect 3574 1368 3630 1402
rect 3664 1368 3720 1402
rect 3754 1368 3831 1402
rect 2869 1349 3831 1368
rect 2869 1345 2941 1349
rect 2869 1311 2888 1345
rect 2922 1311 2941 1345
rect 2869 1255 2941 1311
rect 3759 1326 3831 1349
rect 3759 1292 3778 1326
rect 3812 1292 3831 1326
rect 2869 1221 2888 1255
rect 2922 1221 2941 1255
rect 2869 1165 2941 1221
rect 2869 1131 2888 1165
rect 2922 1131 2941 1165
rect 2869 1075 2941 1131
rect 2869 1041 2888 1075
rect 2922 1041 2941 1075
rect 2869 985 2941 1041
rect 2869 951 2888 985
rect 2922 951 2941 985
rect 2869 895 2941 951
rect 2869 861 2888 895
rect 2922 861 2941 895
rect 2869 805 2941 861
rect 2869 771 2888 805
rect 2922 771 2941 805
rect 2869 715 2941 771
rect 2869 681 2888 715
rect 2922 681 2941 715
rect 2869 625 2941 681
rect 2869 591 2888 625
rect 2922 591 2941 625
rect 3003 1228 3697 1287
rect 3003 1194 3064 1228
rect 3098 1200 3154 1228
rect 3188 1200 3244 1228
rect 3278 1200 3334 1228
rect 3110 1194 3154 1200
rect 3210 1194 3244 1200
rect 3310 1194 3334 1200
rect 3368 1200 3424 1228
rect 3368 1194 3376 1200
rect 3003 1166 3076 1194
rect 3110 1166 3176 1194
rect 3210 1166 3276 1194
rect 3310 1166 3376 1194
rect 3410 1194 3424 1200
rect 3458 1200 3514 1228
rect 3458 1194 3476 1200
rect 3410 1166 3476 1194
rect 3510 1194 3514 1200
rect 3548 1200 3604 1228
rect 3548 1194 3576 1200
rect 3638 1194 3697 1228
rect 3510 1166 3576 1194
rect 3610 1166 3697 1194
rect 3003 1138 3697 1166
rect 3003 1104 3064 1138
rect 3098 1104 3154 1138
rect 3188 1104 3244 1138
rect 3278 1104 3334 1138
rect 3368 1104 3424 1138
rect 3458 1104 3514 1138
rect 3548 1104 3604 1138
rect 3638 1104 3697 1138
rect 3003 1100 3697 1104
rect 3003 1066 3076 1100
rect 3110 1066 3176 1100
rect 3210 1066 3276 1100
rect 3310 1066 3376 1100
rect 3410 1066 3476 1100
rect 3510 1066 3576 1100
rect 3610 1066 3697 1100
rect 3003 1048 3697 1066
rect 3003 1014 3064 1048
rect 3098 1014 3154 1048
rect 3188 1014 3244 1048
rect 3278 1014 3334 1048
rect 3368 1014 3424 1048
rect 3458 1014 3514 1048
rect 3548 1014 3604 1048
rect 3638 1014 3697 1048
rect 3003 1000 3697 1014
rect 3003 966 3076 1000
rect 3110 966 3176 1000
rect 3210 966 3276 1000
rect 3310 966 3376 1000
rect 3410 966 3476 1000
rect 3510 966 3576 1000
rect 3610 966 3697 1000
rect 3003 958 3697 966
rect 3003 924 3064 958
rect 3098 924 3154 958
rect 3188 924 3244 958
rect 3278 924 3334 958
rect 3368 924 3424 958
rect 3458 924 3514 958
rect 3548 924 3604 958
rect 3638 924 3697 958
rect 3003 900 3697 924
rect 3003 868 3076 900
rect 3110 868 3176 900
rect 3210 868 3276 900
rect 3310 868 3376 900
rect 3003 834 3064 868
rect 3110 866 3154 868
rect 3210 866 3244 868
rect 3310 866 3334 868
rect 3098 834 3154 866
rect 3188 834 3244 866
rect 3278 834 3334 866
rect 3368 866 3376 868
rect 3410 868 3476 900
rect 3410 866 3424 868
rect 3368 834 3424 866
rect 3458 866 3476 868
rect 3510 868 3576 900
rect 3610 868 3697 900
rect 3510 866 3514 868
rect 3458 834 3514 866
rect 3548 866 3576 868
rect 3548 834 3604 866
rect 3638 834 3697 868
rect 3003 800 3697 834
rect 3003 778 3076 800
rect 3110 778 3176 800
rect 3210 778 3276 800
rect 3310 778 3376 800
rect 3003 744 3064 778
rect 3110 766 3154 778
rect 3210 766 3244 778
rect 3310 766 3334 778
rect 3098 744 3154 766
rect 3188 744 3244 766
rect 3278 744 3334 766
rect 3368 766 3376 778
rect 3410 778 3476 800
rect 3410 766 3424 778
rect 3368 744 3424 766
rect 3458 766 3476 778
rect 3510 778 3576 800
rect 3610 778 3697 800
rect 3510 766 3514 778
rect 3458 744 3514 766
rect 3548 766 3576 778
rect 3548 744 3604 766
rect 3638 744 3697 778
rect 3003 700 3697 744
rect 3003 688 3076 700
rect 3110 688 3176 700
rect 3210 688 3276 700
rect 3310 688 3376 700
rect 3003 654 3064 688
rect 3110 666 3154 688
rect 3210 666 3244 688
rect 3310 666 3334 688
rect 3098 654 3154 666
rect 3188 654 3244 666
rect 3278 654 3334 666
rect 3368 666 3376 688
rect 3410 688 3476 700
rect 3410 666 3424 688
rect 3368 654 3424 666
rect 3458 666 3476 688
rect 3510 688 3576 700
rect 3610 688 3697 700
rect 3510 666 3514 688
rect 3458 654 3514 666
rect 3548 666 3576 688
rect 3548 654 3604 666
rect 3638 654 3697 688
rect 3003 593 3697 654
rect 3759 1236 3831 1292
rect 3759 1202 3778 1236
rect 3812 1202 3831 1236
rect 3759 1146 3831 1202
rect 3759 1112 3778 1146
rect 3812 1112 3831 1146
rect 3759 1056 3831 1112
rect 3759 1022 3778 1056
rect 3812 1022 3831 1056
rect 3759 966 3831 1022
rect 3759 932 3778 966
rect 3812 932 3831 966
rect 3759 876 3831 932
rect 3759 842 3778 876
rect 3812 842 3831 876
rect 3759 786 3831 842
rect 3759 752 3778 786
rect 3812 752 3831 786
rect 3759 696 3831 752
rect 3759 662 3778 696
rect 3812 662 3831 696
rect 3759 606 3831 662
rect 2869 531 2941 591
rect 3759 572 3778 606
rect 3812 572 3831 606
rect 3759 531 3831 572
rect 2869 512 3831 531
rect 2869 478 2966 512
rect 3000 478 3056 512
rect 3090 478 3146 512
rect 3180 478 3236 512
rect 3270 478 3326 512
rect 3360 478 3416 512
rect 3450 478 3506 512
rect 3540 478 3596 512
rect 3630 478 3686 512
rect 3720 478 3831 512
rect 2869 470 3831 478
rect 3895 1402 3927 1410
rect 3961 1402 4080 1436
rect 4114 1410 5267 1436
rect 4114 1402 4145 1410
rect 3895 1346 4145 1402
rect 3895 1312 3927 1346
rect 3961 1312 4080 1346
rect 4114 1312 4145 1346
rect 3895 1256 4145 1312
rect 3895 1222 3927 1256
rect 3961 1222 4080 1256
rect 4114 1222 4145 1256
rect 3895 1166 4145 1222
rect 3895 1132 3927 1166
rect 3961 1132 4080 1166
rect 4114 1132 4145 1166
rect 3895 1076 4145 1132
rect 3895 1042 3927 1076
rect 3961 1042 4080 1076
rect 4114 1042 4145 1076
rect 3895 986 4145 1042
rect 3895 952 3927 986
rect 3961 952 4080 986
rect 4114 952 4145 986
rect 3895 896 4145 952
rect 3895 862 3927 896
rect 3961 862 4080 896
rect 4114 862 4145 896
rect 3895 806 4145 862
rect 3895 772 3927 806
rect 3961 772 4080 806
rect 4114 772 4145 806
rect 3895 716 4145 772
rect 3895 682 3927 716
rect 3961 682 4080 716
rect 4114 682 4145 716
rect 3895 626 4145 682
rect 3895 592 3927 626
rect 3961 592 4080 626
rect 4114 592 4145 626
rect 3895 536 4145 592
rect 3895 502 3927 536
rect 3961 502 4080 536
rect 4114 502 4145 536
rect 3895 470 4145 502
rect 4209 1402 5171 1410
rect 4209 1368 4340 1402
rect 4374 1368 4430 1402
rect 4464 1368 4520 1402
rect 4554 1368 4610 1402
rect 4644 1368 4700 1402
rect 4734 1368 4790 1402
rect 4824 1368 4880 1402
rect 4914 1368 4970 1402
rect 5004 1368 5060 1402
rect 5094 1368 5171 1402
rect 4209 1349 5171 1368
rect 4209 1345 4281 1349
rect 4209 1311 4228 1345
rect 4262 1311 4281 1345
rect 4209 1255 4281 1311
rect 5099 1326 5171 1349
rect 5099 1292 5118 1326
rect 5152 1292 5171 1326
rect 4209 1221 4228 1255
rect 4262 1221 4281 1255
rect 4209 1165 4281 1221
rect 4209 1131 4228 1165
rect 4262 1131 4281 1165
rect 4209 1075 4281 1131
rect 4209 1041 4228 1075
rect 4262 1041 4281 1075
rect 4209 985 4281 1041
rect 4209 951 4228 985
rect 4262 951 4281 985
rect 4209 895 4281 951
rect 4209 861 4228 895
rect 4262 861 4281 895
rect 4209 805 4281 861
rect 4209 771 4228 805
rect 4262 771 4281 805
rect 4209 715 4281 771
rect 4209 681 4228 715
rect 4262 681 4281 715
rect 4209 625 4281 681
rect 4209 591 4228 625
rect 4262 591 4281 625
rect 4343 1228 5037 1287
rect 4343 1194 4404 1228
rect 4438 1200 4494 1228
rect 4528 1200 4584 1228
rect 4618 1200 4674 1228
rect 4450 1194 4494 1200
rect 4550 1194 4584 1200
rect 4650 1194 4674 1200
rect 4708 1200 4764 1228
rect 4708 1194 4716 1200
rect 4343 1166 4416 1194
rect 4450 1166 4516 1194
rect 4550 1166 4616 1194
rect 4650 1166 4716 1194
rect 4750 1194 4764 1200
rect 4798 1200 4854 1228
rect 4798 1194 4816 1200
rect 4750 1166 4816 1194
rect 4850 1194 4854 1200
rect 4888 1200 4944 1228
rect 4888 1194 4916 1200
rect 4978 1194 5037 1228
rect 4850 1166 4916 1194
rect 4950 1166 5037 1194
rect 4343 1138 5037 1166
rect 4343 1104 4404 1138
rect 4438 1104 4494 1138
rect 4528 1104 4584 1138
rect 4618 1104 4674 1138
rect 4708 1104 4764 1138
rect 4798 1104 4854 1138
rect 4888 1104 4944 1138
rect 4978 1104 5037 1138
rect 4343 1100 5037 1104
rect 4343 1066 4416 1100
rect 4450 1066 4516 1100
rect 4550 1066 4616 1100
rect 4650 1066 4716 1100
rect 4750 1066 4816 1100
rect 4850 1066 4916 1100
rect 4950 1066 5037 1100
rect 4343 1048 5037 1066
rect 4343 1014 4404 1048
rect 4438 1014 4494 1048
rect 4528 1014 4584 1048
rect 4618 1014 4674 1048
rect 4708 1014 4764 1048
rect 4798 1014 4854 1048
rect 4888 1014 4944 1048
rect 4978 1014 5037 1048
rect 4343 1000 5037 1014
rect 4343 966 4416 1000
rect 4450 966 4516 1000
rect 4550 966 4616 1000
rect 4650 966 4716 1000
rect 4750 966 4816 1000
rect 4850 966 4916 1000
rect 4950 966 5037 1000
rect 4343 958 5037 966
rect 4343 924 4404 958
rect 4438 924 4494 958
rect 4528 924 4584 958
rect 4618 924 4674 958
rect 4708 924 4764 958
rect 4798 924 4854 958
rect 4888 924 4944 958
rect 4978 924 5037 958
rect 4343 900 5037 924
rect 4343 868 4416 900
rect 4450 868 4516 900
rect 4550 868 4616 900
rect 4650 868 4716 900
rect 4343 834 4404 868
rect 4450 866 4494 868
rect 4550 866 4584 868
rect 4650 866 4674 868
rect 4438 834 4494 866
rect 4528 834 4584 866
rect 4618 834 4674 866
rect 4708 866 4716 868
rect 4750 868 4816 900
rect 4750 866 4764 868
rect 4708 834 4764 866
rect 4798 866 4816 868
rect 4850 868 4916 900
rect 4950 868 5037 900
rect 4850 866 4854 868
rect 4798 834 4854 866
rect 4888 866 4916 868
rect 4888 834 4944 866
rect 4978 834 5037 868
rect 4343 800 5037 834
rect 4343 778 4416 800
rect 4450 778 4516 800
rect 4550 778 4616 800
rect 4650 778 4716 800
rect 4343 744 4404 778
rect 4450 766 4494 778
rect 4550 766 4584 778
rect 4650 766 4674 778
rect 4438 744 4494 766
rect 4528 744 4584 766
rect 4618 744 4674 766
rect 4708 766 4716 778
rect 4750 778 4816 800
rect 4750 766 4764 778
rect 4708 744 4764 766
rect 4798 766 4816 778
rect 4850 778 4916 800
rect 4950 778 5037 800
rect 4850 766 4854 778
rect 4798 744 4854 766
rect 4888 766 4916 778
rect 4888 744 4944 766
rect 4978 744 5037 778
rect 4343 700 5037 744
rect 4343 688 4416 700
rect 4450 688 4516 700
rect 4550 688 4616 700
rect 4650 688 4716 700
rect 4343 654 4404 688
rect 4450 666 4494 688
rect 4550 666 4584 688
rect 4650 666 4674 688
rect 4438 654 4494 666
rect 4528 654 4584 666
rect 4618 654 4674 666
rect 4708 666 4716 688
rect 4750 688 4816 700
rect 4750 666 4764 688
rect 4708 654 4764 666
rect 4798 666 4816 688
rect 4850 688 4916 700
rect 4950 688 5037 700
rect 4850 666 4854 688
rect 4798 654 4854 666
rect 4888 666 4916 688
rect 4888 654 4944 666
rect 4978 654 5037 688
rect 4343 593 5037 654
rect 5099 1236 5171 1292
rect 5099 1202 5118 1236
rect 5152 1202 5171 1236
rect 5099 1146 5171 1202
rect 5099 1112 5118 1146
rect 5152 1112 5171 1146
rect 5099 1056 5171 1112
rect 5099 1022 5118 1056
rect 5152 1022 5171 1056
rect 5099 966 5171 1022
rect 5099 932 5118 966
rect 5152 932 5171 966
rect 5099 876 5171 932
rect 5099 842 5118 876
rect 5152 842 5171 876
rect 5099 786 5171 842
rect 5099 752 5118 786
rect 5152 752 5171 786
rect 5099 696 5171 752
rect 5099 662 5118 696
rect 5152 662 5171 696
rect 5099 606 5171 662
rect 4209 531 4281 591
rect 5099 572 5118 606
rect 5152 572 5171 606
rect 5099 531 5171 572
rect 4209 512 5171 531
rect 4209 478 4306 512
rect 4340 478 4396 512
rect 4430 478 4486 512
rect 4520 478 4576 512
rect 4610 478 4666 512
rect 4700 478 4756 512
rect 4790 478 4846 512
rect 4880 478 4936 512
rect 4970 478 5026 512
rect 5060 478 5171 512
rect 4209 470 5171 478
rect 5235 1402 5267 1410
rect 5301 1402 5420 1436
rect 5454 1410 6607 1436
rect 5454 1402 5485 1410
rect 5235 1346 5485 1402
rect 5235 1312 5267 1346
rect 5301 1312 5420 1346
rect 5454 1312 5485 1346
rect 5235 1256 5485 1312
rect 5235 1222 5267 1256
rect 5301 1222 5420 1256
rect 5454 1222 5485 1256
rect 5235 1166 5485 1222
rect 5235 1132 5267 1166
rect 5301 1132 5420 1166
rect 5454 1132 5485 1166
rect 5235 1076 5485 1132
rect 5235 1042 5267 1076
rect 5301 1042 5420 1076
rect 5454 1042 5485 1076
rect 5235 986 5485 1042
rect 5235 952 5267 986
rect 5301 952 5420 986
rect 5454 952 5485 986
rect 5235 896 5485 952
rect 5235 862 5267 896
rect 5301 862 5420 896
rect 5454 862 5485 896
rect 5235 806 5485 862
rect 5235 772 5267 806
rect 5301 772 5420 806
rect 5454 772 5485 806
rect 5235 716 5485 772
rect 5235 682 5267 716
rect 5301 682 5420 716
rect 5454 682 5485 716
rect 5235 626 5485 682
rect 5235 592 5267 626
rect 5301 592 5420 626
rect 5454 592 5485 626
rect 5235 536 5485 592
rect 5235 502 5267 536
rect 5301 502 5420 536
rect 5454 502 5485 536
rect 5235 470 5485 502
rect 5549 1402 6511 1410
rect 5549 1368 5680 1402
rect 5714 1368 5770 1402
rect 5804 1368 5860 1402
rect 5894 1368 5950 1402
rect 5984 1368 6040 1402
rect 6074 1368 6130 1402
rect 6164 1368 6220 1402
rect 6254 1368 6310 1402
rect 6344 1368 6400 1402
rect 6434 1368 6511 1402
rect 5549 1349 6511 1368
rect 5549 1345 5621 1349
rect 5549 1311 5568 1345
rect 5602 1311 5621 1345
rect 5549 1255 5621 1311
rect 6439 1326 6511 1349
rect 6439 1292 6458 1326
rect 6492 1292 6511 1326
rect 5549 1221 5568 1255
rect 5602 1221 5621 1255
rect 5549 1165 5621 1221
rect 5549 1131 5568 1165
rect 5602 1131 5621 1165
rect 5549 1075 5621 1131
rect 5549 1041 5568 1075
rect 5602 1041 5621 1075
rect 5549 985 5621 1041
rect 5549 951 5568 985
rect 5602 951 5621 985
rect 5549 895 5621 951
rect 5549 861 5568 895
rect 5602 861 5621 895
rect 5549 805 5621 861
rect 5549 771 5568 805
rect 5602 771 5621 805
rect 5549 715 5621 771
rect 5549 681 5568 715
rect 5602 681 5621 715
rect 5549 625 5621 681
rect 5549 591 5568 625
rect 5602 591 5621 625
rect 5683 1228 6377 1287
rect 5683 1194 5744 1228
rect 5778 1200 5834 1228
rect 5868 1200 5924 1228
rect 5958 1200 6014 1228
rect 5790 1194 5834 1200
rect 5890 1194 5924 1200
rect 5990 1194 6014 1200
rect 6048 1200 6104 1228
rect 6048 1194 6056 1200
rect 5683 1166 5756 1194
rect 5790 1166 5856 1194
rect 5890 1166 5956 1194
rect 5990 1166 6056 1194
rect 6090 1194 6104 1200
rect 6138 1200 6194 1228
rect 6138 1194 6156 1200
rect 6090 1166 6156 1194
rect 6190 1194 6194 1200
rect 6228 1200 6284 1228
rect 6228 1194 6256 1200
rect 6318 1194 6377 1228
rect 6190 1166 6256 1194
rect 6290 1166 6377 1194
rect 5683 1138 6377 1166
rect 5683 1104 5744 1138
rect 5778 1104 5834 1138
rect 5868 1104 5924 1138
rect 5958 1104 6014 1138
rect 6048 1104 6104 1138
rect 6138 1104 6194 1138
rect 6228 1104 6284 1138
rect 6318 1104 6377 1138
rect 5683 1100 6377 1104
rect 5683 1066 5756 1100
rect 5790 1066 5856 1100
rect 5890 1066 5956 1100
rect 5990 1066 6056 1100
rect 6090 1066 6156 1100
rect 6190 1066 6256 1100
rect 6290 1066 6377 1100
rect 5683 1048 6377 1066
rect 5683 1014 5744 1048
rect 5778 1014 5834 1048
rect 5868 1014 5924 1048
rect 5958 1014 6014 1048
rect 6048 1014 6104 1048
rect 6138 1014 6194 1048
rect 6228 1014 6284 1048
rect 6318 1014 6377 1048
rect 5683 1000 6377 1014
rect 5683 966 5756 1000
rect 5790 966 5856 1000
rect 5890 966 5956 1000
rect 5990 966 6056 1000
rect 6090 966 6156 1000
rect 6190 966 6256 1000
rect 6290 966 6377 1000
rect 5683 958 6377 966
rect 5683 924 5744 958
rect 5778 924 5834 958
rect 5868 924 5924 958
rect 5958 924 6014 958
rect 6048 924 6104 958
rect 6138 924 6194 958
rect 6228 924 6284 958
rect 6318 924 6377 958
rect 5683 900 6377 924
rect 5683 868 5756 900
rect 5790 868 5856 900
rect 5890 868 5956 900
rect 5990 868 6056 900
rect 5683 834 5744 868
rect 5790 866 5834 868
rect 5890 866 5924 868
rect 5990 866 6014 868
rect 5778 834 5834 866
rect 5868 834 5924 866
rect 5958 834 6014 866
rect 6048 866 6056 868
rect 6090 868 6156 900
rect 6090 866 6104 868
rect 6048 834 6104 866
rect 6138 866 6156 868
rect 6190 868 6256 900
rect 6290 868 6377 900
rect 6190 866 6194 868
rect 6138 834 6194 866
rect 6228 866 6256 868
rect 6228 834 6284 866
rect 6318 834 6377 868
rect 5683 800 6377 834
rect 5683 778 5756 800
rect 5790 778 5856 800
rect 5890 778 5956 800
rect 5990 778 6056 800
rect 5683 744 5744 778
rect 5790 766 5834 778
rect 5890 766 5924 778
rect 5990 766 6014 778
rect 5778 744 5834 766
rect 5868 744 5924 766
rect 5958 744 6014 766
rect 6048 766 6056 778
rect 6090 778 6156 800
rect 6090 766 6104 778
rect 6048 744 6104 766
rect 6138 766 6156 778
rect 6190 778 6256 800
rect 6290 778 6377 800
rect 6190 766 6194 778
rect 6138 744 6194 766
rect 6228 766 6256 778
rect 6228 744 6284 766
rect 6318 744 6377 778
rect 5683 700 6377 744
rect 5683 688 5756 700
rect 5790 688 5856 700
rect 5890 688 5956 700
rect 5990 688 6056 700
rect 5683 654 5744 688
rect 5790 666 5834 688
rect 5890 666 5924 688
rect 5990 666 6014 688
rect 5778 654 5834 666
rect 5868 654 5924 666
rect 5958 654 6014 666
rect 6048 666 6056 688
rect 6090 688 6156 700
rect 6090 666 6104 688
rect 6048 654 6104 666
rect 6138 666 6156 688
rect 6190 688 6256 700
rect 6290 688 6377 700
rect 6190 666 6194 688
rect 6138 654 6194 666
rect 6228 666 6256 688
rect 6228 654 6284 666
rect 6318 654 6377 688
rect 5683 593 6377 654
rect 6439 1236 6511 1292
rect 6439 1202 6458 1236
rect 6492 1202 6511 1236
rect 6439 1146 6511 1202
rect 6439 1112 6458 1146
rect 6492 1112 6511 1146
rect 6439 1056 6511 1112
rect 6439 1022 6458 1056
rect 6492 1022 6511 1056
rect 6439 966 6511 1022
rect 6439 932 6458 966
rect 6492 932 6511 966
rect 6439 876 6511 932
rect 6439 842 6458 876
rect 6492 842 6511 876
rect 6439 786 6511 842
rect 6439 752 6458 786
rect 6492 752 6511 786
rect 6439 696 6511 752
rect 6439 662 6458 696
rect 6492 662 6511 696
rect 6439 606 6511 662
rect 5549 531 5621 591
rect 6439 572 6458 606
rect 6492 572 6511 606
rect 6439 531 6511 572
rect 5549 512 6511 531
rect 5549 478 5646 512
rect 5680 478 5736 512
rect 5770 478 5826 512
rect 5860 478 5916 512
rect 5950 478 6006 512
rect 6040 478 6096 512
rect 6130 478 6186 512
rect 6220 478 6276 512
rect 6310 478 6366 512
rect 6400 478 6511 512
rect 5549 470 6511 478
rect 6575 1402 6607 1410
rect 6641 1402 6760 1436
rect 6794 1410 7947 1436
rect 6794 1402 6825 1410
rect 6575 1346 6825 1402
rect 6575 1312 6607 1346
rect 6641 1312 6760 1346
rect 6794 1312 6825 1346
rect 6575 1256 6825 1312
rect 6575 1222 6607 1256
rect 6641 1222 6760 1256
rect 6794 1222 6825 1256
rect 6575 1166 6825 1222
rect 6575 1132 6607 1166
rect 6641 1132 6760 1166
rect 6794 1132 6825 1166
rect 6575 1076 6825 1132
rect 6575 1042 6607 1076
rect 6641 1042 6760 1076
rect 6794 1042 6825 1076
rect 6575 986 6825 1042
rect 6575 952 6607 986
rect 6641 952 6760 986
rect 6794 952 6825 986
rect 6575 896 6825 952
rect 6575 862 6607 896
rect 6641 862 6760 896
rect 6794 862 6825 896
rect 6575 806 6825 862
rect 6575 772 6607 806
rect 6641 772 6760 806
rect 6794 772 6825 806
rect 6575 716 6825 772
rect 6575 682 6607 716
rect 6641 682 6760 716
rect 6794 682 6825 716
rect 6575 626 6825 682
rect 6575 592 6607 626
rect 6641 592 6760 626
rect 6794 592 6825 626
rect 6575 536 6825 592
rect 6575 502 6607 536
rect 6641 502 6760 536
rect 6794 502 6825 536
rect 6575 470 6825 502
rect 6889 1402 7851 1410
rect 6889 1368 7020 1402
rect 7054 1368 7110 1402
rect 7144 1368 7200 1402
rect 7234 1368 7290 1402
rect 7324 1368 7380 1402
rect 7414 1368 7470 1402
rect 7504 1368 7560 1402
rect 7594 1368 7650 1402
rect 7684 1368 7740 1402
rect 7774 1368 7851 1402
rect 6889 1349 7851 1368
rect 6889 1345 6961 1349
rect 6889 1311 6908 1345
rect 6942 1311 6961 1345
rect 6889 1255 6961 1311
rect 7779 1326 7851 1349
rect 7779 1292 7798 1326
rect 7832 1292 7851 1326
rect 6889 1221 6908 1255
rect 6942 1221 6961 1255
rect 6889 1165 6961 1221
rect 6889 1131 6908 1165
rect 6942 1131 6961 1165
rect 6889 1075 6961 1131
rect 6889 1041 6908 1075
rect 6942 1041 6961 1075
rect 6889 985 6961 1041
rect 6889 951 6908 985
rect 6942 951 6961 985
rect 6889 895 6961 951
rect 6889 861 6908 895
rect 6942 861 6961 895
rect 6889 805 6961 861
rect 6889 771 6908 805
rect 6942 771 6961 805
rect 6889 715 6961 771
rect 6889 681 6908 715
rect 6942 681 6961 715
rect 6889 625 6961 681
rect 6889 591 6908 625
rect 6942 591 6961 625
rect 7023 1228 7717 1287
rect 7023 1194 7084 1228
rect 7118 1200 7174 1228
rect 7208 1200 7264 1228
rect 7298 1200 7354 1228
rect 7130 1194 7174 1200
rect 7230 1194 7264 1200
rect 7330 1194 7354 1200
rect 7388 1200 7444 1228
rect 7388 1194 7396 1200
rect 7023 1166 7096 1194
rect 7130 1166 7196 1194
rect 7230 1166 7296 1194
rect 7330 1166 7396 1194
rect 7430 1194 7444 1200
rect 7478 1200 7534 1228
rect 7478 1194 7496 1200
rect 7430 1166 7496 1194
rect 7530 1194 7534 1200
rect 7568 1200 7624 1228
rect 7568 1194 7596 1200
rect 7658 1194 7717 1228
rect 7530 1166 7596 1194
rect 7630 1166 7717 1194
rect 7023 1138 7717 1166
rect 7023 1104 7084 1138
rect 7118 1104 7174 1138
rect 7208 1104 7264 1138
rect 7298 1104 7354 1138
rect 7388 1104 7444 1138
rect 7478 1104 7534 1138
rect 7568 1104 7624 1138
rect 7658 1104 7717 1138
rect 7023 1100 7717 1104
rect 7023 1066 7096 1100
rect 7130 1066 7196 1100
rect 7230 1066 7296 1100
rect 7330 1066 7396 1100
rect 7430 1066 7496 1100
rect 7530 1066 7596 1100
rect 7630 1066 7717 1100
rect 7023 1048 7717 1066
rect 7023 1014 7084 1048
rect 7118 1014 7174 1048
rect 7208 1014 7264 1048
rect 7298 1014 7354 1048
rect 7388 1014 7444 1048
rect 7478 1014 7534 1048
rect 7568 1014 7624 1048
rect 7658 1014 7717 1048
rect 7023 1000 7717 1014
rect 7023 966 7096 1000
rect 7130 966 7196 1000
rect 7230 966 7296 1000
rect 7330 966 7396 1000
rect 7430 966 7496 1000
rect 7530 966 7596 1000
rect 7630 966 7717 1000
rect 7023 958 7717 966
rect 7023 924 7084 958
rect 7118 924 7174 958
rect 7208 924 7264 958
rect 7298 924 7354 958
rect 7388 924 7444 958
rect 7478 924 7534 958
rect 7568 924 7624 958
rect 7658 924 7717 958
rect 7023 900 7717 924
rect 7023 868 7096 900
rect 7130 868 7196 900
rect 7230 868 7296 900
rect 7330 868 7396 900
rect 7023 834 7084 868
rect 7130 866 7174 868
rect 7230 866 7264 868
rect 7330 866 7354 868
rect 7118 834 7174 866
rect 7208 834 7264 866
rect 7298 834 7354 866
rect 7388 866 7396 868
rect 7430 868 7496 900
rect 7430 866 7444 868
rect 7388 834 7444 866
rect 7478 866 7496 868
rect 7530 868 7596 900
rect 7630 868 7717 900
rect 7530 866 7534 868
rect 7478 834 7534 866
rect 7568 866 7596 868
rect 7568 834 7624 866
rect 7658 834 7717 868
rect 7023 800 7717 834
rect 7023 778 7096 800
rect 7130 778 7196 800
rect 7230 778 7296 800
rect 7330 778 7396 800
rect 7023 744 7084 778
rect 7130 766 7174 778
rect 7230 766 7264 778
rect 7330 766 7354 778
rect 7118 744 7174 766
rect 7208 744 7264 766
rect 7298 744 7354 766
rect 7388 766 7396 778
rect 7430 778 7496 800
rect 7430 766 7444 778
rect 7388 744 7444 766
rect 7478 766 7496 778
rect 7530 778 7596 800
rect 7630 778 7717 800
rect 7530 766 7534 778
rect 7478 744 7534 766
rect 7568 766 7596 778
rect 7568 744 7624 766
rect 7658 744 7717 778
rect 7023 700 7717 744
rect 7023 688 7096 700
rect 7130 688 7196 700
rect 7230 688 7296 700
rect 7330 688 7396 700
rect 7023 654 7084 688
rect 7130 666 7174 688
rect 7230 666 7264 688
rect 7330 666 7354 688
rect 7118 654 7174 666
rect 7208 654 7264 666
rect 7298 654 7354 666
rect 7388 666 7396 688
rect 7430 688 7496 700
rect 7430 666 7444 688
rect 7388 654 7444 666
rect 7478 666 7496 688
rect 7530 688 7596 700
rect 7630 688 7717 700
rect 7530 666 7534 688
rect 7478 654 7534 666
rect 7568 666 7596 688
rect 7568 654 7624 666
rect 7658 654 7717 688
rect 7023 593 7717 654
rect 7779 1236 7851 1292
rect 7779 1202 7798 1236
rect 7832 1202 7851 1236
rect 7779 1146 7851 1202
rect 7779 1112 7798 1146
rect 7832 1112 7851 1146
rect 7779 1056 7851 1112
rect 7779 1022 7798 1056
rect 7832 1022 7851 1056
rect 7779 966 7851 1022
rect 7779 932 7798 966
rect 7832 932 7851 966
rect 7779 876 7851 932
rect 7779 842 7798 876
rect 7832 842 7851 876
rect 7779 786 7851 842
rect 7779 752 7798 786
rect 7832 752 7851 786
rect 7779 696 7851 752
rect 7779 662 7798 696
rect 7832 662 7851 696
rect 7779 606 7851 662
rect 6889 531 6961 591
rect 7779 572 7798 606
rect 7832 572 7851 606
rect 7779 531 7851 572
rect 6889 512 7851 531
rect 6889 478 6986 512
rect 7020 478 7076 512
rect 7110 478 7166 512
rect 7200 478 7256 512
rect 7290 478 7346 512
rect 7380 478 7436 512
rect 7470 478 7526 512
rect 7560 478 7616 512
rect 7650 478 7706 512
rect 7740 478 7851 512
rect 6889 470 7851 478
rect 7915 1402 7947 1410
rect 7981 1402 8100 1436
rect 8134 1410 9287 1436
rect 8134 1402 8165 1410
rect 7915 1346 8165 1402
rect 7915 1312 7947 1346
rect 7981 1312 8100 1346
rect 8134 1312 8165 1346
rect 7915 1256 8165 1312
rect 7915 1222 7947 1256
rect 7981 1222 8100 1256
rect 8134 1222 8165 1256
rect 7915 1166 8165 1222
rect 7915 1132 7947 1166
rect 7981 1132 8100 1166
rect 8134 1132 8165 1166
rect 7915 1076 8165 1132
rect 7915 1042 7947 1076
rect 7981 1042 8100 1076
rect 8134 1042 8165 1076
rect 7915 986 8165 1042
rect 7915 952 7947 986
rect 7981 952 8100 986
rect 8134 952 8165 986
rect 7915 896 8165 952
rect 7915 862 7947 896
rect 7981 862 8100 896
rect 8134 862 8165 896
rect 7915 806 8165 862
rect 7915 772 7947 806
rect 7981 772 8100 806
rect 8134 772 8165 806
rect 7915 716 8165 772
rect 7915 682 7947 716
rect 7981 682 8100 716
rect 8134 682 8165 716
rect 7915 626 8165 682
rect 7915 592 7947 626
rect 7981 592 8100 626
rect 8134 592 8165 626
rect 7915 536 8165 592
rect 7915 502 7947 536
rect 7981 502 8100 536
rect 8134 502 8165 536
rect 7915 470 8165 502
rect 8229 1402 9191 1410
rect 8229 1368 8360 1402
rect 8394 1368 8450 1402
rect 8484 1368 8540 1402
rect 8574 1368 8630 1402
rect 8664 1368 8720 1402
rect 8754 1368 8810 1402
rect 8844 1368 8900 1402
rect 8934 1368 8990 1402
rect 9024 1368 9080 1402
rect 9114 1368 9191 1402
rect 8229 1349 9191 1368
rect 8229 1345 8301 1349
rect 8229 1311 8248 1345
rect 8282 1311 8301 1345
rect 8229 1255 8301 1311
rect 9119 1326 9191 1349
rect 9119 1292 9138 1326
rect 9172 1292 9191 1326
rect 8229 1221 8248 1255
rect 8282 1221 8301 1255
rect 8229 1165 8301 1221
rect 8229 1131 8248 1165
rect 8282 1131 8301 1165
rect 8229 1075 8301 1131
rect 8229 1041 8248 1075
rect 8282 1041 8301 1075
rect 8229 985 8301 1041
rect 8229 951 8248 985
rect 8282 951 8301 985
rect 8229 895 8301 951
rect 8229 861 8248 895
rect 8282 861 8301 895
rect 8229 805 8301 861
rect 8229 771 8248 805
rect 8282 771 8301 805
rect 8229 715 8301 771
rect 8229 681 8248 715
rect 8282 681 8301 715
rect 8229 625 8301 681
rect 8229 591 8248 625
rect 8282 591 8301 625
rect 8363 1228 9057 1287
rect 8363 1194 8424 1228
rect 8458 1200 8514 1228
rect 8548 1200 8604 1228
rect 8638 1200 8694 1228
rect 8470 1194 8514 1200
rect 8570 1194 8604 1200
rect 8670 1194 8694 1200
rect 8728 1200 8784 1228
rect 8728 1194 8736 1200
rect 8363 1166 8436 1194
rect 8470 1166 8536 1194
rect 8570 1166 8636 1194
rect 8670 1166 8736 1194
rect 8770 1194 8784 1200
rect 8818 1200 8874 1228
rect 8818 1194 8836 1200
rect 8770 1166 8836 1194
rect 8870 1194 8874 1200
rect 8908 1200 8964 1228
rect 8908 1194 8936 1200
rect 8998 1194 9057 1228
rect 8870 1166 8936 1194
rect 8970 1166 9057 1194
rect 8363 1138 9057 1166
rect 8363 1104 8424 1138
rect 8458 1104 8514 1138
rect 8548 1104 8604 1138
rect 8638 1104 8694 1138
rect 8728 1104 8784 1138
rect 8818 1104 8874 1138
rect 8908 1104 8964 1138
rect 8998 1104 9057 1138
rect 8363 1100 9057 1104
rect 8363 1066 8436 1100
rect 8470 1066 8536 1100
rect 8570 1066 8636 1100
rect 8670 1066 8736 1100
rect 8770 1066 8836 1100
rect 8870 1066 8936 1100
rect 8970 1066 9057 1100
rect 8363 1048 9057 1066
rect 8363 1014 8424 1048
rect 8458 1014 8514 1048
rect 8548 1014 8604 1048
rect 8638 1014 8694 1048
rect 8728 1014 8784 1048
rect 8818 1014 8874 1048
rect 8908 1014 8964 1048
rect 8998 1014 9057 1048
rect 8363 1000 9057 1014
rect 8363 966 8436 1000
rect 8470 966 8536 1000
rect 8570 966 8636 1000
rect 8670 966 8736 1000
rect 8770 966 8836 1000
rect 8870 966 8936 1000
rect 8970 966 9057 1000
rect 8363 958 9057 966
rect 8363 924 8424 958
rect 8458 924 8514 958
rect 8548 924 8604 958
rect 8638 924 8694 958
rect 8728 924 8784 958
rect 8818 924 8874 958
rect 8908 924 8964 958
rect 8998 924 9057 958
rect 8363 900 9057 924
rect 8363 868 8436 900
rect 8470 868 8536 900
rect 8570 868 8636 900
rect 8670 868 8736 900
rect 8363 834 8424 868
rect 8470 866 8514 868
rect 8570 866 8604 868
rect 8670 866 8694 868
rect 8458 834 8514 866
rect 8548 834 8604 866
rect 8638 834 8694 866
rect 8728 866 8736 868
rect 8770 868 8836 900
rect 8770 866 8784 868
rect 8728 834 8784 866
rect 8818 866 8836 868
rect 8870 868 8936 900
rect 8970 868 9057 900
rect 8870 866 8874 868
rect 8818 834 8874 866
rect 8908 866 8936 868
rect 8908 834 8964 866
rect 8998 834 9057 868
rect 8363 800 9057 834
rect 8363 778 8436 800
rect 8470 778 8536 800
rect 8570 778 8636 800
rect 8670 778 8736 800
rect 8363 744 8424 778
rect 8470 766 8514 778
rect 8570 766 8604 778
rect 8670 766 8694 778
rect 8458 744 8514 766
rect 8548 744 8604 766
rect 8638 744 8694 766
rect 8728 766 8736 778
rect 8770 778 8836 800
rect 8770 766 8784 778
rect 8728 744 8784 766
rect 8818 766 8836 778
rect 8870 778 8936 800
rect 8970 778 9057 800
rect 8870 766 8874 778
rect 8818 744 8874 766
rect 8908 766 8936 778
rect 8908 744 8964 766
rect 8998 744 9057 778
rect 8363 700 9057 744
rect 8363 688 8436 700
rect 8470 688 8536 700
rect 8570 688 8636 700
rect 8670 688 8736 700
rect 8363 654 8424 688
rect 8470 666 8514 688
rect 8570 666 8604 688
rect 8670 666 8694 688
rect 8458 654 8514 666
rect 8548 654 8604 666
rect 8638 654 8694 666
rect 8728 666 8736 688
rect 8770 688 8836 700
rect 8770 666 8784 688
rect 8728 654 8784 666
rect 8818 666 8836 688
rect 8870 688 8936 700
rect 8970 688 9057 700
rect 8870 666 8874 688
rect 8818 654 8874 666
rect 8908 666 8936 688
rect 8908 654 8964 666
rect 8998 654 9057 688
rect 8363 593 9057 654
rect 9119 1236 9191 1292
rect 9119 1202 9138 1236
rect 9172 1202 9191 1236
rect 9119 1146 9191 1202
rect 9119 1112 9138 1146
rect 9172 1112 9191 1146
rect 9119 1056 9191 1112
rect 9119 1022 9138 1056
rect 9172 1022 9191 1056
rect 9119 966 9191 1022
rect 9119 932 9138 966
rect 9172 932 9191 966
rect 9119 876 9191 932
rect 9119 842 9138 876
rect 9172 842 9191 876
rect 9119 786 9191 842
rect 9119 752 9138 786
rect 9172 752 9191 786
rect 9119 696 9191 752
rect 9119 662 9138 696
rect 9172 662 9191 696
rect 9119 606 9191 662
rect 8229 531 8301 591
rect 9119 572 9138 606
rect 9172 572 9191 606
rect 9119 531 9191 572
rect 8229 512 9191 531
rect 8229 478 8326 512
rect 8360 478 8416 512
rect 8450 478 8506 512
rect 8540 478 8596 512
rect 8630 478 8686 512
rect 8720 478 8776 512
rect 8810 478 8866 512
rect 8900 478 8956 512
rect 8990 478 9046 512
rect 9080 478 9191 512
rect 8229 470 9191 478
rect 9255 1402 9287 1410
rect 9321 1410 9357 1436
rect 9321 1402 9354 1410
rect 9255 1346 9354 1402
rect 9255 1312 9287 1346
rect 9321 1312 9354 1346
rect 9255 1256 9354 1312
rect 9255 1222 9287 1256
rect 9321 1222 9354 1256
rect 9255 1166 9354 1222
rect 9255 1132 9287 1166
rect 9321 1132 9354 1166
rect 9255 1076 9354 1132
rect 9255 1042 9287 1076
rect 9321 1042 9354 1076
rect 9255 986 9354 1042
rect 9255 952 9287 986
rect 9321 952 9354 986
rect 9255 896 9354 952
rect 9255 862 9287 896
rect 9321 862 9354 896
rect 9255 806 9354 862
rect 9255 772 9287 806
rect 9321 772 9354 806
rect 9255 716 9354 772
rect 9255 682 9287 716
rect 9321 682 9354 716
rect 9255 626 9354 682
rect 9255 592 9287 626
rect 9321 592 9354 626
rect 9255 536 9354 592
rect 9255 502 9287 536
rect 9321 502 9354 536
rect 9255 470 9354 502
rect 26 446 9357 470
rect 26 412 60 446
rect 94 412 1247 446
rect 1281 412 1400 446
rect 1434 412 2587 446
rect 2621 412 2740 446
rect 2774 412 3927 446
rect 3961 412 4080 446
rect 4114 412 5267 446
rect 5301 412 5420 446
rect 5454 412 6607 446
rect 6641 412 6760 446
rect 6794 412 7947 446
rect 7981 412 8100 446
rect 8134 412 9287 446
rect 9321 412 9357 446
rect 26 362 9357 412
rect 26 328 156 362
rect 190 328 246 362
rect 280 328 336 362
rect 370 328 426 362
rect 460 328 516 362
rect 550 328 606 362
rect 640 328 696 362
rect 730 328 786 362
rect 820 328 876 362
rect 910 328 966 362
rect 1000 328 1056 362
rect 1090 328 1146 362
rect 1180 328 1496 362
rect 1530 328 1586 362
rect 1620 328 1676 362
rect 1710 328 1766 362
rect 1800 328 1856 362
rect 1890 328 1946 362
rect 1980 328 2036 362
rect 2070 328 2126 362
rect 2160 328 2216 362
rect 2250 328 2306 362
rect 2340 328 2396 362
rect 2430 328 2486 362
rect 2520 328 2836 362
rect 2870 328 2926 362
rect 2960 328 3016 362
rect 3050 328 3106 362
rect 3140 328 3196 362
rect 3230 328 3286 362
rect 3320 328 3376 362
rect 3410 328 3466 362
rect 3500 328 3556 362
rect 3590 328 3646 362
rect 3680 328 3736 362
rect 3770 328 3826 362
rect 3860 328 4176 362
rect 4210 328 4266 362
rect 4300 328 4356 362
rect 4390 328 4446 362
rect 4480 328 4536 362
rect 4570 328 4626 362
rect 4660 328 4716 362
rect 4750 328 4806 362
rect 4840 328 4896 362
rect 4930 328 4986 362
rect 5020 328 5076 362
rect 5110 328 5166 362
rect 5200 328 5516 362
rect 5550 328 5606 362
rect 5640 328 5696 362
rect 5730 328 5786 362
rect 5820 328 5876 362
rect 5910 328 5966 362
rect 6000 328 6056 362
rect 6090 328 6146 362
rect 6180 328 6236 362
rect 6270 328 6326 362
rect 6360 328 6416 362
rect 6450 328 6506 362
rect 6540 328 6856 362
rect 6890 328 6946 362
rect 6980 328 7036 362
rect 7070 328 7126 362
rect 7160 328 7216 362
rect 7250 328 7306 362
rect 7340 328 7396 362
rect 7430 328 7486 362
rect 7520 328 7576 362
rect 7610 328 7666 362
rect 7700 328 7756 362
rect 7790 328 7846 362
rect 7880 328 8196 362
rect 8230 328 8286 362
rect 8320 328 8376 362
rect 8410 328 8466 362
rect 8500 328 8556 362
rect 8590 328 8646 362
rect 8680 328 8736 362
rect 8770 328 8826 362
rect 8860 328 8916 362
rect 8950 328 9006 362
rect 9040 328 9096 362
rect 9130 328 9186 362
rect 9220 328 9357 362
rect 26 296 9357 328
rect 0 -30 170 30
rect 230 -30 370 30
rect 430 -30 570 30
rect 630 -30 770 30
rect 830 -30 970 30
rect 1030 -30 1170 30
rect 1230 -30 1370 30
rect 1430 -30 1570 30
rect 1630 -30 1770 30
rect 1830 -30 1970 30
rect 2030 -30 2170 30
rect 2230 -30 2370 30
rect 2430 -30 2570 30
rect 2630 -30 2770 30
rect 2830 -30 2970 30
rect 3030 -30 3170 30
rect 3230 -30 3370 30
rect 3430 -30 3570 30
rect 3630 -30 3770 30
rect 3830 -30 3970 30
rect 4030 -30 4170 30
rect 4230 -30 4370 30
rect 4430 -30 4570 30
rect 4630 -30 4770 30
rect 4830 -30 4970 30
rect 5030 -30 5170 30
rect 5230 -30 5370 30
rect 5430 -30 5570 30
rect 5630 -30 5770 30
rect 5830 -30 5970 30
rect 6030 -30 6170 30
rect 6230 -30 6370 30
rect 6430 -30 6570 30
rect 6630 -30 6770 30
rect 6830 -30 6970 30
rect 7030 -30 7170 30
rect 7230 -30 7370 30
rect 7430 -30 7570 30
rect 7630 -30 7770 30
rect 7830 -30 7970 30
rect 8030 -30 8170 30
rect 8230 -30 8370 30
rect 8430 -30 8570 30
rect 8630 -30 8770 30
rect 8830 -30 8970 30
rect 9030 -30 9170 30
rect 9230 -30 9380 30
<< viali >>
rect 170 1850 230 1910
rect 370 1850 430 1910
rect 570 1850 630 1910
rect 770 1850 830 1910
rect 970 1850 1030 1910
rect 1170 1850 1230 1910
rect 1370 1850 1430 1910
rect 1570 1850 1630 1910
rect 1770 1850 1830 1910
rect 1970 1850 2030 1910
rect 2170 1850 2230 1910
rect 2370 1850 2430 1910
rect 2570 1850 2630 1910
rect 2770 1850 2830 1910
rect 2970 1850 3030 1910
rect 3170 1850 3230 1910
rect 3370 1850 3430 1910
rect 3570 1850 3630 1910
rect 3770 1850 3830 1910
rect 3970 1850 4030 1910
rect 4170 1850 4230 1910
rect 4370 1850 4430 1910
rect 4570 1850 4630 1910
rect 4770 1850 4830 1910
rect 4970 1850 5030 1910
rect 5170 1850 5230 1910
rect 5370 1850 5430 1910
rect 5570 1850 5630 1910
rect 5770 1850 5830 1910
rect 5970 1850 6030 1910
rect 6170 1850 6230 1910
rect 6370 1850 6430 1910
rect 6570 1850 6630 1910
rect 6770 1850 6830 1910
rect 6970 1850 7030 1910
rect 7170 1850 7230 1910
rect 7370 1850 7430 1910
rect 7570 1850 7630 1910
rect 7770 1850 7830 1910
rect 7970 1850 8030 1910
rect 8170 1850 8230 1910
rect 8370 1850 8430 1910
rect 8570 1850 8630 1910
rect 8770 1850 8830 1910
rect 8970 1850 9030 1910
rect 9170 1850 9230 1910
rect 396 1194 418 1200
rect 418 1194 430 1200
rect 496 1194 508 1200
rect 508 1194 530 1200
rect 596 1194 598 1200
rect 598 1194 630 1200
rect 396 1166 430 1194
rect 496 1166 530 1194
rect 596 1166 630 1194
rect 696 1166 730 1200
rect 796 1166 830 1200
rect 896 1194 924 1200
rect 924 1194 930 1200
rect 896 1166 930 1194
rect 396 1066 430 1100
rect 496 1066 530 1100
rect 596 1066 630 1100
rect 696 1066 730 1100
rect 796 1066 830 1100
rect 896 1066 930 1100
rect 396 966 430 1000
rect 496 966 530 1000
rect 596 966 630 1000
rect 696 966 730 1000
rect 796 966 830 1000
rect 896 966 930 1000
rect 396 868 430 900
rect 496 868 530 900
rect 596 868 630 900
rect 396 866 418 868
rect 418 866 430 868
rect 496 866 508 868
rect 508 866 530 868
rect 596 866 598 868
rect 598 866 630 868
rect 696 866 730 900
rect 796 866 830 900
rect 896 868 930 900
rect 896 866 924 868
rect 924 866 930 868
rect 396 778 430 800
rect 496 778 530 800
rect 596 778 630 800
rect 396 766 418 778
rect 418 766 430 778
rect 496 766 508 778
rect 508 766 530 778
rect 596 766 598 778
rect 598 766 630 778
rect 696 766 730 800
rect 796 766 830 800
rect 896 778 930 800
rect 896 766 924 778
rect 924 766 930 778
rect 396 688 430 700
rect 496 688 530 700
rect 596 688 630 700
rect 396 666 418 688
rect 418 666 430 688
rect 496 666 508 688
rect 508 666 530 688
rect 596 666 598 688
rect 598 666 630 688
rect 696 666 730 700
rect 796 666 830 700
rect 896 688 930 700
rect 896 666 924 688
rect 924 666 930 688
rect 1736 1194 1758 1200
rect 1758 1194 1770 1200
rect 1836 1194 1848 1200
rect 1848 1194 1870 1200
rect 1936 1194 1938 1200
rect 1938 1194 1970 1200
rect 1736 1166 1770 1194
rect 1836 1166 1870 1194
rect 1936 1166 1970 1194
rect 2036 1166 2070 1200
rect 2136 1166 2170 1200
rect 2236 1194 2264 1200
rect 2264 1194 2270 1200
rect 2236 1166 2270 1194
rect 1736 1066 1770 1100
rect 1836 1066 1870 1100
rect 1936 1066 1970 1100
rect 2036 1066 2070 1100
rect 2136 1066 2170 1100
rect 2236 1066 2270 1100
rect 1736 966 1770 1000
rect 1836 966 1870 1000
rect 1936 966 1970 1000
rect 2036 966 2070 1000
rect 2136 966 2170 1000
rect 2236 966 2270 1000
rect 1736 868 1770 900
rect 1836 868 1870 900
rect 1936 868 1970 900
rect 1736 866 1758 868
rect 1758 866 1770 868
rect 1836 866 1848 868
rect 1848 866 1870 868
rect 1936 866 1938 868
rect 1938 866 1970 868
rect 2036 866 2070 900
rect 2136 866 2170 900
rect 2236 868 2270 900
rect 2236 866 2264 868
rect 2264 866 2270 868
rect 1736 778 1770 800
rect 1836 778 1870 800
rect 1936 778 1970 800
rect 1736 766 1758 778
rect 1758 766 1770 778
rect 1836 766 1848 778
rect 1848 766 1870 778
rect 1936 766 1938 778
rect 1938 766 1970 778
rect 2036 766 2070 800
rect 2136 766 2170 800
rect 2236 778 2270 800
rect 2236 766 2264 778
rect 2264 766 2270 778
rect 1736 688 1770 700
rect 1836 688 1870 700
rect 1936 688 1970 700
rect 1736 666 1758 688
rect 1758 666 1770 688
rect 1836 666 1848 688
rect 1848 666 1870 688
rect 1936 666 1938 688
rect 1938 666 1970 688
rect 2036 666 2070 700
rect 2136 666 2170 700
rect 2236 688 2270 700
rect 2236 666 2264 688
rect 2264 666 2270 688
rect 3076 1194 3098 1200
rect 3098 1194 3110 1200
rect 3176 1194 3188 1200
rect 3188 1194 3210 1200
rect 3276 1194 3278 1200
rect 3278 1194 3310 1200
rect 3076 1166 3110 1194
rect 3176 1166 3210 1194
rect 3276 1166 3310 1194
rect 3376 1166 3410 1200
rect 3476 1166 3510 1200
rect 3576 1194 3604 1200
rect 3604 1194 3610 1200
rect 3576 1166 3610 1194
rect 3076 1066 3110 1100
rect 3176 1066 3210 1100
rect 3276 1066 3310 1100
rect 3376 1066 3410 1100
rect 3476 1066 3510 1100
rect 3576 1066 3610 1100
rect 3076 966 3110 1000
rect 3176 966 3210 1000
rect 3276 966 3310 1000
rect 3376 966 3410 1000
rect 3476 966 3510 1000
rect 3576 966 3610 1000
rect 3076 868 3110 900
rect 3176 868 3210 900
rect 3276 868 3310 900
rect 3076 866 3098 868
rect 3098 866 3110 868
rect 3176 866 3188 868
rect 3188 866 3210 868
rect 3276 866 3278 868
rect 3278 866 3310 868
rect 3376 866 3410 900
rect 3476 866 3510 900
rect 3576 868 3610 900
rect 3576 866 3604 868
rect 3604 866 3610 868
rect 3076 778 3110 800
rect 3176 778 3210 800
rect 3276 778 3310 800
rect 3076 766 3098 778
rect 3098 766 3110 778
rect 3176 766 3188 778
rect 3188 766 3210 778
rect 3276 766 3278 778
rect 3278 766 3310 778
rect 3376 766 3410 800
rect 3476 766 3510 800
rect 3576 778 3610 800
rect 3576 766 3604 778
rect 3604 766 3610 778
rect 3076 688 3110 700
rect 3176 688 3210 700
rect 3276 688 3310 700
rect 3076 666 3098 688
rect 3098 666 3110 688
rect 3176 666 3188 688
rect 3188 666 3210 688
rect 3276 666 3278 688
rect 3278 666 3310 688
rect 3376 666 3410 700
rect 3476 666 3510 700
rect 3576 688 3610 700
rect 3576 666 3604 688
rect 3604 666 3610 688
rect 4416 1194 4438 1200
rect 4438 1194 4450 1200
rect 4516 1194 4528 1200
rect 4528 1194 4550 1200
rect 4616 1194 4618 1200
rect 4618 1194 4650 1200
rect 4416 1166 4450 1194
rect 4516 1166 4550 1194
rect 4616 1166 4650 1194
rect 4716 1166 4750 1200
rect 4816 1166 4850 1200
rect 4916 1194 4944 1200
rect 4944 1194 4950 1200
rect 4916 1166 4950 1194
rect 4416 1066 4450 1100
rect 4516 1066 4550 1100
rect 4616 1066 4650 1100
rect 4716 1066 4750 1100
rect 4816 1066 4850 1100
rect 4916 1066 4950 1100
rect 4416 966 4450 1000
rect 4516 966 4550 1000
rect 4616 966 4650 1000
rect 4716 966 4750 1000
rect 4816 966 4850 1000
rect 4916 966 4950 1000
rect 4416 868 4450 900
rect 4516 868 4550 900
rect 4616 868 4650 900
rect 4416 866 4438 868
rect 4438 866 4450 868
rect 4516 866 4528 868
rect 4528 866 4550 868
rect 4616 866 4618 868
rect 4618 866 4650 868
rect 4716 866 4750 900
rect 4816 866 4850 900
rect 4916 868 4950 900
rect 4916 866 4944 868
rect 4944 866 4950 868
rect 4416 778 4450 800
rect 4516 778 4550 800
rect 4616 778 4650 800
rect 4416 766 4438 778
rect 4438 766 4450 778
rect 4516 766 4528 778
rect 4528 766 4550 778
rect 4616 766 4618 778
rect 4618 766 4650 778
rect 4716 766 4750 800
rect 4816 766 4850 800
rect 4916 778 4950 800
rect 4916 766 4944 778
rect 4944 766 4950 778
rect 4416 688 4450 700
rect 4516 688 4550 700
rect 4616 688 4650 700
rect 4416 666 4438 688
rect 4438 666 4450 688
rect 4516 666 4528 688
rect 4528 666 4550 688
rect 4616 666 4618 688
rect 4618 666 4650 688
rect 4716 666 4750 700
rect 4816 666 4850 700
rect 4916 688 4950 700
rect 4916 666 4944 688
rect 4944 666 4950 688
rect 5756 1194 5778 1200
rect 5778 1194 5790 1200
rect 5856 1194 5868 1200
rect 5868 1194 5890 1200
rect 5956 1194 5958 1200
rect 5958 1194 5990 1200
rect 5756 1166 5790 1194
rect 5856 1166 5890 1194
rect 5956 1166 5990 1194
rect 6056 1166 6090 1200
rect 6156 1166 6190 1200
rect 6256 1194 6284 1200
rect 6284 1194 6290 1200
rect 6256 1166 6290 1194
rect 5756 1066 5790 1100
rect 5856 1066 5890 1100
rect 5956 1066 5990 1100
rect 6056 1066 6090 1100
rect 6156 1066 6190 1100
rect 6256 1066 6290 1100
rect 5756 966 5790 1000
rect 5856 966 5890 1000
rect 5956 966 5990 1000
rect 6056 966 6090 1000
rect 6156 966 6190 1000
rect 6256 966 6290 1000
rect 5756 868 5790 900
rect 5856 868 5890 900
rect 5956 868 5990 900
rect 5756 866 5778 868
rect 5778 866 5790 868
rect 5856 866 5868 868
rect 5868 866 5890 868
rect 5956 866 5958 868
rect 5958 866 5990 868
rect 6056 866 6090 900
rect 6156 866 6190 900
rect 6256 868 6290 900
rect 6256 866 6284 868
rect 6284 866 6290 868
rect 5756 778 5790 800
rect 5856 778 5890 800
rect 5956 778 5990 800
rect 5756 766 5778 778
rect 5778 766 5790 778
rect 5856 766 5868 778
rect 5868 766 5890 778
rect 5956 766 5958 778
rect 5958 766 5990 778
rect 6056 766 6090 800
rect 6156 766 6190 800
rect 6256 778 6290 800
rect 6256 766 6284 778
rect 6284 766 6290 778
rect 5756 688 5790 700
rect 5856 688 5890 700
rect 5956 688 5990 700
rect 5756 666 5778 688
rect 5778 666 5790 688
rect 5856 666 5868 688
rect 5868 666 5890 688
rect 5956 666 5958 688
rect 5958 666 5990 688
rect 6056 666 6090 700
rect 6156 666 6190 700
rect 6256 688 6290 700
rect 6256 666 6284 688
rect 6284 666 6290 688
rect 7096 1194 7118 1200
rect 7118 1194 7130 1200
rect 7196 1194 7208 1200
rect 7208 1194 7230 1200
rect 7296 1194 7298 1200
rect 7298 1194 7330 1200
rect 7096 1166 7130 1194
rect 7196 1166 7230 1194
rect 7296 1166 7330 1194
rect 7396 1166 7430 1200
rect 7496 1166 7530 1200
rect 7596 1194 7624 1200
rect 7624 1194 7630 1200
rect 7596 1166 7630 1194
rect 7096 1066 7130 1100
rect 7196 1066 7230 1100
rect 7296 1066 7330 1100
rect 7396 1066 7430 1100
rect 7496 1066 7530 1100
rect 7596 1066 7630 1100
rect 7096 966 7130 1000
rect 7196 966 7230 1000
rect 7296 966 7330 1000
rect 7396 966 7430 1000
rect 7496 966 7530 1000
rect 7596 966 7630 1000
rect 7096 868 7130 900
rect 7196 868 7230 900
rect 7296 868 7330 900
rect 7096 866 7118 868
rect 7118 866 7130 868
rect 7196 866 7208 868
rect 7208 866 7230 868
rect 7296 866 7298 868
rect 7298 866 7330 868
rect 7396 866 7430 900
rect 7496 866 7530 900
rect 7596 868 7630 900
rect 7596 866 7624 868
rect 7624 866 7630 868
rect 7096 778 7130 800
rect 7196 778 7230 800
rect 7296 778 7330 800
rect 7096 766 7118 778
rect 7118 766 7130 778
rect 7196 766 7208 778
rect 7208 766 7230 778
rect 7296 766 7298 778
rect 7298 766 7330 778
rect 7396 766 7430 800
rect 7496 766 7530 800
rect 7596 778 7630 800
rect 7596 766 7624 778
rect 7624 766 7630 778
rect 7096 688 7130 700
rect 7196 688 7230 700
rect 7296 688 7330 700
rect 7096 666 7118 688
rect 7118 666 7130 688
rect 7196 666 7208 688
rect 7208 666 7230 688
rect 7296 666 7298 688
rect 7298 666 7330 688
rect 7396 666 7430 700
rect 7496 666 7530 700
rect 7596 688 7630 700
rect 7596 666 7624 688
rect 7624 666 7630 688
rect 8436 1194 8458 1200
rect 8458 1194 8470 1200
rect 8536 1194 8548 1200
rect 8548 1194 8570 1200
rect 8636 1194 8638 1200
rect 8638 1194 8670 1200
rect 8436 1166 8470 1194
rect 8536 1166 8570 1194
rect 8636 1166 8670 1194
rect 8736 1166 8770 1200
rect 8836 1166 8870 1200
rect 8936 1194 8964 1200
rect 8964 1194 8970 1200
rect 8936 1166 8970 1194
rect 8436 1066 8470 1100
rect 8536 1066 8570 1100
rect 8636 1066 8670 1100
rect 8736 1066 8770 1100
rect 8836 1066 8870 1100
rect 8936 1066 8970 1100
rect 8436 966 8470 1000
rect 8536 966 8570 1000
rect 8636 966 8670 1000
rect 8736 966 8770 1000
rect 8836 966 8870 1000
rect 8936 966 8970 1000
rect 8436 868 8470 900
rect 8536 868 8570 900
rect 8636 868 8670 900
rect 8436 866 8458 868
rect 8458 866 8470 868
rect 8536 866 8548 868
rect 8548 866 8570 868
rect 8636 866 8638 868
rect 8638 866 8670 868
rect 8736 866 8770 900
rect 8836 866 8870 900
rect 8936 868 8970 900
rect 8936 866 8964 868
rect 8964 866 8970 868
rect 8436 778 8470 800
rect 8536 778 8570 800
rect 8636 778 8670 800
rect 8436 766 8458 778
rect 8458 766 8470 778
rect 8536 766 8548 778
rect 8548 766 8570 778
rect 8636 766 8638 778
rect 8638 766 8670 778
rect 8736 766 8770 800
rect 8836 766 8870 800
rect 8936 778 8970 800
rect 8936 766 8964 778
rect 8964 766 8970 778
rect 8436 688 8470 700
rect 8536 688 8570 700
rect 8636 688 8670 700
rect 8436 666 8458 688
rect 8458 666 8470 688
rect 8536 666 8548 688
rect 8548 666 8570 688
rect 8636 666 8638 688
rect 8638 666 8670 688
rect 8736 666 8770 700
rect 8836 666 8870 700
rect 8936 688 8970 700
rect 8936 666 8964 688
rect 8964 666 8970 688
rect 170 -30 230 30
rect 370 -30 430 30
rect 570 -30 630 30
rect 770 -30 830 30
rect 970 -30 1030 30
rect 1170 -30 1230 30
rect 1370 -30 1430 30
rect 1570 -30 1630 30
rect 1770 -30 1830 30
rect 1970 -30 2030 30
rect 2170 -30 2230 30
rect 2370 -30 2430 30
rect 2570 -30 2630 30
rect 2770 -30 2830 30
rect 2970 -30 3030 30
rect 3170 -30 3230 30
rect 3370 -30 3430 30
rect 3570 -30 3630 30
rect 3770 -30 3830 30
rect 3970 -30 4030 30
rect 4170 -30 4230 30
rect 4370 -30 4430 30
rect 4570 -30 4630 30
rect 4770 -30 4830 30
rect 4970 -30 5030 30
rect 5170 -30 5230 30
rect 5370 -30 5430 30
rect 5570 -30 5630 30
rect 5770 -30 5830 30
rect 5970 -30 6030 30
rect 6170 -30 6230 30
rect 6370 -30 6430 30
rect 6570 -30 6630 30
rect 6770 -30 6830 30
rect 6970 -30 7030 30
rect 7170 -30 7230 30
rect 7370 -30 7430 30
rect 7570 -30 7630 30
rect 7770 -30 7830 30
rect 7970 -30 8030 30
rect 8170 -30 8230 30
rect 8370 -30 8430 30
rect 8570 -30 8630 30
rect 8770 -30 8830 30
rect 8970 -30 9030 30
rect 9170 -30 9230 30
<< metal1 >>
rect 0 1910 9380 1940
rect 0 1850 170 1910
rect 230 1850 370 1910
rect 430 1850 570 1910
rect 630 1850 770 1910
rect 830 1850 970 1910
rect 1030 1850 1170 1910
rect 1230 1850 1370 1910
rect 1430 1850 1570 1910
rect 1630 1850 1770 1910
rect 1830 1850 1970 1910
rect 2030 1850 2170 1910
rect 2230 1850 2370 1910
rect 2430 1850 2570 1910
rect 2630 1850 2770 1910
rect 2830 1850 2970 1910
rect 3030 1850 3170 1910
rect 3230 1850 3370 1910
rect 3430 1850 3570 1910
rect 3630 1850 3770 1910
rect 3830 1850 3970 1910
rect 4030 1850 4170 1910
rect 4230 1850 4370 1910
rect 4430 1850 4570 1910
rect 4630 1850 4770 1910
rect 4830 1850 4970 1910
rect 5030 1850 5170 1910
rect 5230 1850 5370 1910
rect 5430 1850 5570 1910
rect 5630 1850 5770 1910
rect 5830 1850 5970 1910
rect 6030 1850 6170 1910
rect 6230 1850 6370 1910
rect 6430 1850 6570 1910
rect 6630 1850 6770 1910
rect 6830 1850 6970 1910
rect 7030 1850 7170 1910
rect 7230 1850 7370 1910
rect 7430 1850 7570 1910
rect 7630 1850 7770 1910
rect 7830 1850 7970 1910
rect 8030 1850 8170 1910
rect 8230 1850 8370 1910
rect 8430 1850 8570 1910
rect 8630 1850 8770 1910
rect 8830 1850 8970 1910
rect 9030 1850 9170 1910
rect 9230 1850 9380 1910
rect 0 1820 9380 1850
rect 364 1200 9062 1246
rect 364 1166 396 1200
rect 430 1166 496 1200
rect 530 1166 596 1200
rect 630 1166 696 1200
rect 730 1166 796 1200
rect 830 1166 896 1200
rect 930 1166 1736 1200
rect 1770 1166 1836 1200
rect 1870 1166 1936 1200
rect 1970 1166 2036 1200
rect 2070 1166 2136 1200
rect 2170 1166 2236 1200
rect 2270 1166 3076 1200
rect 3110 1166 3176 1200
rect 3210 1166 3276 1200
rect 3310 1166 3376 1200
rect 3410 1166 3476 1200
rect 3510 1166 3576 1200
rect 3610 1166 4416 1200
rect 4450 1166 4516 1200
rect 4550 1166 4616 1200
rect 4650 1166 4716 1200
rect 4750 1166 4816 1200
rect 4850 1166 4916 1200
rect 4950 1166 5756 1200
rect 5790 1166 5856 1200
rect 5890 1166 5956 1200
rect 5990 1166 6056 1200
rect 6090 1166 6156 1200
rect 6190 1166 6256 1200
rect 6290 1166 7096 1200
rect 7130 1166 7196 1200
rect 7230 1166 7296 1200
rect 7330 1166 7396 1200
rect 7430 1166 7496 1200
rect 7530 1166 7596 1200
rect 7630 1166 8436 1200
rect 8470 1166 8536 1200
rect 8570 1166 8636 1200
rect 8670 1166 8736 1200
rect 8770 1166 8836 1200
rect 8870 1166 8936 1200
rect 8970 1166 9062 1200
rect 364 1100 9062 1166
rect 364 1066 396 1100
rect 430 1066 496 1100
rect 530 1066 596 1100
rect 630 1066 696 1100
rect 730 1066 796 1100
rect 830 1066 896 1100
rect 930 1066 1736 1100
rect 1770 1066 1836 1100
rect 1870 1066 1936 1100
rect 1970 1066 2036 1100
rect 2070 1066 2136 1100
rect 2170 1066 2236 1100
rect 2270 1066 3076 1100
rect 3110 1066 3176 1100
rect 3210 1066 3276 1100
rect 3310 1066 3376 1100
rect 3410 1066 3476 1100
rect 3510 1066 3576 1100
rect 3610 1066 4416 1100
rect 4450 1066 4516 1100
rect 4550 1066 4616 1100
rect 4650 1066 4716 1100
rect 4750 1066 4816 1100
rect 4850 1066 4916 1100
rect 4950 1066 5756 1100
rect 5790 1066 5856 1100
rect 5890 1066 5956 1100
rect 5990 1066 6056 1100
rect 6090 1066 6156 1100
rect 6190 1066 6256 1100
rect 6290 1066 7096 1100
rect 7130 1066 7196 1100
rect 7230 1066 7296 1100
rect 7330 1066 7396 1100
rect 7430 1066 7496 1100
rect 7530 1066 7596 1100
rect 7630 1066 8436 1100
rect 8470 1066 8536 1100
rect 8570 1066 8636 1100
rect 8670 1066 8736 1100
rect 8770 1066 8836 1100
rect 8870 1066 8936 1100
rect 8970 1066 9062 1100
rect 364 1000 9062 1066
rect 364 966 396 1000
rect 430 966 496 1000
rect 530 966 596 1000
rect 630 966 696 1000
rect 730 966 796 1000
rect 830 966 896 1000
rect 930 966 1736 1000
rect 1770 966 1836 1000
rect 1870 966 1936 1000
rect 1970 966 2036 1000
rect 2070 966 2136 1000
rect 2170 966 2236 1000
rect 2270 966 3076 1000
rect 3110 966 3176 1000
rect 3210 966 3276 1000
rect 3310 966 3376 1000
rect 3410 966 3476 1000
rect 3510 966 3576 1000
rect 3610 966 4416 1000
rect 4450 966 4516 1000
rect 4550 966 4616 1000
rect 4650 966 4716 1000
rect 4750 966 4816 1000
rect 4850 966 4916 1000
rect 4950 966 5756 1000
rect 5790 966 5856 1000
rect 5890 966 5956 1000
rect 5990 966 6056 1000
rect 6090 966 6156 1000
rect 6190 966 6256 1000
rect 6290 966 7096 1000
rect 7130 966 7196 1000
rect 7230 966 7296 1000
rect 7330 966 7396 1000
rect 7430 966 7496 1000
rect 7530 966 7596 1000
rect 7630 966 8436 1000
rect 8470 966 8536 1000
rect 8570 966 8636 1000
rect 8670 966 8736 1000
rect 8770 966 8836 1000
rect 8870 966 8936 1000
rect 8970 966 9062 1000
rect 364 900 9062 966
rect 364 866 396 900
rect 430 866 496 900
rect 530 866 596 900
rect 630 866 696 900
rect 730 866 796 900
rect 830 866 896 900
rect 930 866 1736 900
rect 1770 866 1836 900
rect 1870 866 1936 900
rect 1970 866 2036 900
rect 2070 866 2136 900
rect 2170 866 2236 900
rect 2270 866 3076 900
rect 3110 866 3176 900
rect 3210 866 3276 900
rect 3310 866 3376 900
rect 3410 866 3476 900
rect 3510 866 3576 900
rect 3610 866 4416 900
rect 4450 866 4516 900
rect 4550 866 4616 900
rect 4650 866 4716 900
rect 4750 866 4816 900
rect 4850 866 4916 900
rect 4950 866 5756 900
rect 5790 866 5856 900
rect 5890 866 5956 900
rect 5990 866 6056 900
rect 6090 866 6156 900
rect 6190 866 6256 900
rect 6290 866 7096 900
rect 7130 866 7196 900
rect 7230 866 7296 900
rect 7330 866 7396 900
rect 7430 866 7496 900
rect 7530 866 7596 900
rect 7630 866 8436 900
rect 8470 866 8536 900
rect 8570 866 8636 900
rect 8670 866 8736 900
rect 8770 866 8836 900
rect 8870 866 8936 900
rect 8970 866 9062 900
rect 364 800 9062 866
rect 364 766 396 800
rect 430 766 496 800
rect 530 766 596 800
rect 630 766 696 800
rect 730 766 796 800
rect 830 766 896 800
rect 930 766 1736 800
rect 1770 766 1836 800
rect 1870 766 1936 800
rect 1970 766 2036 800
rect 2070 766 2136 800
rect 2170 766 2236 800
rect 2270 766 3076 800
rect 3110 766 3176 800
rect 3210 766 3276 800
rect 3310 766 3376 800
rect 3410 766 3476 800
rect 3510 766 3576 800
rect 3610 766 4416 800
rect 4450 766 4516 800
rect 4550 766 4616 800
rect 4650 766 4716 800
rect 4750 766 4816 800
rect 4850 766 4916 800
rect 4950 766 5756 800
rect 5790 766 5856 800
rect 5890 766 5956 800
rect 5990 766 6056 800
rect 6090 766 6156 800
rect 6190 766 6256 800
rect 6290 766 7096 800
rect 7130 766 7196 800
rect 7230 766 7296 800
rect 7330 766 7396 800
rect 7430 766 7496 800
rect 7530 766 7596 800
rect 7630 766 8436 800
rect 8470 766 8536 800
rect 8570 766 8636 800
rect 8670 766 8736 800
rect 8770 766 8836 800
rect 8870 766 8936 800
rect 8970 766 9062 800
rect 364 700 9062 766
rect 364 666 396 700
rect 430 666 496 700
rect 530 666 596 700
rect 630 666 696 700
rect 730 666 796 700
rect 830 666 896 700
rect 930 666 1736 700
rect 1770 666 1836 700
rect 1870 666 1936 700
rect 1970 666 2036 700
rect 2070 666 2136 700
rect 2170 666 2236 700
rect 2270 666 3076 700
rect 3110 666 3176 700
rect 3210 666 3276 700
rect 3310 666 3376 700
rect 3410 666 3476 700
rect 3510 666 3576 700
rect 3610 666 4416 700
rect 4450 666 4516 700
rect 4550 666 4616 700
rect 4650 666 4716 700
rect 4750 666 4816 700
rect 4850 666 4916 700
rect 4950 666 5756 700
rect 5790 666 5856 700
rect 5890 666 5956 700
rect 5990 666 6056 700
rect 6090 666 6156 700
rect 6190 666 6256 700
rect 6290 666 7096 700
rect 7130 666 7196 700
rect 7230 666 7296 700
rect 7330 666 7396 700
rect 7430 666 7496 700
rect 7530 666 7596 700
rect 7630 666 8436 700
rect 8470 666 8536 700
rect 8570 666 8636 700
rect 8670 666 8736 700
rect 8770 666 8836 700
rect 8870 666 8936 700
rect 8970 666 9062 700
rect 364 634 9062 666
rect 0 30 9380 60
rect 0 -30 170 30
rect 230 -30 370 30
rect 430 -30 570 30
rect 630 -30 770 30
rect 830 -30 970 30
rect 1030 -30 1170 30
rect 1230 -30 1370 30
rect 1430 -30 1570 30
rect 1630 -30 1770 30
rect 1830 -30 1970 30
rect 2030 -30 2170 30
rect 2230 -30 2370 30
rect 2430 -30 2570 30
rect 2630 -30 2770 30
rect 2830 -30 2970 30
rect 3030 -30 3170 30
rect 3230 -30 3370 30
rect 3430 -30 3570 30
rect 3630 -30 3770 30
rect 3830 -30 3970 30
rect 4030 -30 4170 30
rect 4230 -30 4370 30
rect 4430 -30 4570 30
rect 4630 -30 4770 30
rect 4830 -30 4970 30
rect 5030 -30 5170 30
rect 5230 -30 5370 30
rect 5430 -30 5570 30
rect 5630 -30 5770 30
rect 5830 -30 5970 30
rect 6030 -30 6170 30
rect 6230 -30 6370 30
rect 6430 -30 6570 30
rect 6630 -30 6770 30
rect 6830 -30 6970 30
rect 7030 -30 7170 30
rect 7230 -30 7370 30
rect 7430 -30 7570 30
rect 7630 -30 7770 30
rect 7830 -30 7970 30
rect 8030 -30 8170 30
rect 8230 -30 8370 30
rect 8430 -30 8570 30
rect 8630 -30 8770 30
rect 8830 -30 8970 30
rect 9030 -30 9170 30
rect 9230 -30 9380 30
rect 0 -60 9380 -30
<< pnp3p40 >>
rect 153 423 1187 1457
rect 1493 423 2527 1457
rect 2833 423 3867 1457
rect 4173 423 5207 1457
rect 5513 423 6547 1457
rect 6853 423 7887 1457
rect 8193 423 9227 1457
<< labels >>
flabel locali 4830 1524 4950 1564 1 FreeSans 480 0 0 0 Collector
port 3 n default bidirectional
flabel locali 4794 1372 4914 1412 1 FreeSans 480 0 0 0 Base
port 2 n default bidirectional
flabel metal1 4582 1010 4810 1140 1 FreeSans 480 0 0 0 Emitter
port 1 n default bidirectional
flabel metal1 0 1850 60 1910 1 FreeSans 800 0 0 0 VPWR
port 4 n power bidirectional
flabel metal1 0 -30 60 30 1 FreeSans 800 0 0 0 VGND
port 5 n ground bidirectional
flabel locali 8594 896 8842 1000 0 FreeSans 400 0 0 0 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_5/Emitter
flabel locali 8653 1522 8754 1571 0 FreeSans 400 0 0 0 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_5/Collector
flabel locali 8630 1372 8748 1412 0 FreeSans 400 0 0 0 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_5/Base
flabel locali 7254 896 7502 1000 0 FreeSans 400 0 0 0 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_4/Emitter
flabel locali 7313 1522 7414 1571 0 FreeSans 400 0 0 0 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_4/Collector
flabel locali 7290 1372 7408 1412 0 FreeSans 400 0 0 0 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_4/Base
flabel locali 5914 896 6162 1000 0 FreeSans 400 0 0 0 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_3/Emitter
flabel locali 5973 1522 6074 1571 0 FreeSans 400 0 0 0 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_3/Collector
flabel locali 5950 1372 6068 1412 0 FreeSans 400 0 0 0 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_3/Base
flabel locali 4574 896 4822 1000 0 FreeSans 400 0 0 0 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_2/Emitter
flabel locali 4633 1522 4734 1571 0 FreeSans 400 0 0 0 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_2/Collector
flabel locali 4610 1372 4728 1412 0 FreeSans 400 0 0 0 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_2/Base
flabel locali 3234 896 3482 1000 0 FreeSans 400 0 0 0 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_1/Emitter
flabel locali 3293 1522 3394 1571 0 FreeSans 400 0 0 0 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_1/Collector
flabel locali 3270 1372 3388 1412 0 FreeSans 400 0 0 0 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_1/Base
flabel locali 1894 896 2142 1000 0 FreeSans 400 0 0 0 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0/Emitter
flabel locali 1953 1522 2054 1571 0 FreeSans 400 0 0 0 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0/Collector
flabel locali 1930 1372 2048 1412 0 FreeSans 400 0 0 0 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0/Base
flabel locali 554 896 802 1000 0 FreeSans 400 0 0 0 xm1/Emitter
flabel locali 613 1522 714 1571 0 FreeSans 400 0 0 0 xm1/Collector
flabel locali 590 1372 708 1412 0 FreeSans 400 0 0 0 xm1/Base
<< properties >>
string FIXED_BBOX 0 0 9380 1880
string LEFclass CORE
string LEFsite unitasc
<< end >>
