magic
tech sky130A
magscale 1 2
timestamp 1654590091
<< nwell >>
rect 2316 42091 5590 42095
rect 163 41729 5590 42091
rect 163 41445 5588 41729
rect 163 41441 2483 41445
rect 5236 41426 5588 41445
rect 2316 40804 5590 40808
rect 163 40442 5590 40804
rect 163 40158 5588 40442
rect 163 40154 2483 40158
rect 5236 40139 5588 40158
rect 2316 39517 5590 39521
rect 163 39155 5590 39517
rect 163 38871 5588 39155
rect 163 38867 2483 38871
rect 5236 38852 5588 38871
rect 2316 38230 5590 38234
rect 163 37868 5590 38230
rect 163 37584 5588 37868
rect 163 37580 2483 37584
rect 5236 37565 5588 37584
rect 2316 36943 5590 36947
rect 163 36581 5590 36943
rect 163 36297 5588 36581
rect 163 36293 2483 36297
rect 5236 36278 5588 36297
rect 2316 35656 5590 35660
rect 163 35294 5590 35656
rect 163 35010 5588 35294
rect 163 35006 2483 35010
rect 5236 34991 5588 35010
rect 2316 34369 5590 34373
rect 163 34007 5590 34369
rect 163 33723 5588 34007
rect 163 33719 2483 33723
rect 5236 33704 5588 33723
rect 2316 33082 5590 33086
rect 163 32720 5590 33082
rect 163 32436 5588 32720
rect 163 32432 2483 32436
rect 5236 32417 5588 32436
rect 2316 31795 5590 31799
rect 163 31433 5590 31795
rect 163 31149 5588 31433
rect 163 31145 2483 31149
rect 5236 31130 5588 31149
rect 2316 30508 5590 30512
rect 163 30146 5590 30508
rect 163 29862 5588 30146
rect 163 29858 2483 29862
rect 5236 29843 5588 29862
rect 2316 29221 5590 29225
rect 163 28859 5590 29221
rect 163 28575 5588 28859
rect 163 28571 2483 28575
rect 5236 28556 5588 28575
rect 2316 27934 5590 27938
rect 163 27572 5590 27934
rect 163 27288 5588 27572
rect 163 27284 2483 27288
rect 5236 27269 5588 27288
rect 2316 26647 5590 26651
rect 163 26285 5590 26647
rect 163 26001 5588 26285
rect 163 25997 2483 26001
rect 5236 25982 5588 26001
rect 2316 25360 5590 25364
rect 163 24998 5590 25360
rect 163 24714 5588 24998
rect 163 24710 2483 24714
rect 5236 24695 5588 24714
rect 2316 24073 5590 24077
rect 163 23711 5590 24073
rect 163 23427 5588 23711
rect 163 23423 2483 23427
rect 5236 23408 5588 23427
rect 2316 22786 5590 22790
rect 163 22424 5590 22786
rect 163 22140 5588 22424
rect 163 22136 2483 22140
rect 5236 22121 5588 22140
rect 2316 21499 5590 21503
rect 163 21137 5590 21499
rect 163 20853 5588 21137
rect 163 20849 2483 20853
rect 5236 20834 5588 20853
rect 2316 20212 5590 20216
rect 163 19850 5590 20212
rect 163 19566 5588 19850
rect 163 19562 2483 19566
rect 5236 19547 5588 19566
rect 2316 18925 5590 18929
rect 163 18563 5590 18925
rect 163 18279 5588 18563
rect 163 18275 2483 18279
rect 5236 18260 5588 18279
rect 2316 17638 5590 17642
rect 163 17276 5590 17638
rect 163 16992 5588 17276
rect 163 16988 2483 16992
rect 5236 16973 5588 16992
rect 2316 16351 5590 16355
rect 163 15989 5590 16351
rect 163 15705 5588 15989
rect 163 15701 2483 15705
rect 5236 15686 5588 15705
rect 2316 15064 5590 15068
rect 163 14702 5590 15064
rect 163 14418 5588 14702
rect 163 14414 2483 14418
rect 5236 14399 5588 14418
rect 2316 13777 5590 13781
rect 163 13415 5590 13777
rect 163 13131 5588 13415
rect 163 13127 2483 13131
rect 5236 13112 5588 13131
rect 2316 12490 5590 12494
rect 163 12128 5590 12490
rect 163 11844 5588 12128
rect 163 11840 2483 11844
rect 5236 11825 5588 11844
rect 2316 11203 5590 11207
rect 163 10841 5590 11203
rect 163 10557 5588 10841
rect 163 10553 2483 10557
rect 5236 10538 5588 10557
rect 2316 9916 5590 9920
rect 163 9554 5590 9916
rect 163 9270 5588 9554
rect 163 9266 2483 9270
rect 5236 9251 5588 9270
rect 2316 8629 5590 8633
rect 163 8267 5590 8629
rect 163 7983 5588 8267
rect 163 7979 2483 7983
rect 5236 7964 5588 7983
rect 2316 7342 5590 7346
rect 163 6980 5590 7342
rect 163 6696 5588 6980
rect 163 6692 2483 6696
rect 5236 6677 5588 6696
rect 2316 6055 5590 6059
rect 163 5693 5590 6055
rect 163 5409 5588 5693
rect 163 5405 2483 5409
rect 5236 5390 5588 5409
rect 2316 4768 5590 4772
rect 163 4406 5590 4768
rect 163 4122 5588 4406
rect 163 4118 2483 4122
rect 5236 4103 5588 4122
rect 2316 3481 5590 3485
rect 163 3119 5590 3481
rect 163 2835 5588 3119
rect 163 2831 2483 2835
rect 5236 2816 5588 2835
rect 2316 2194 5590 2198
rect 163 1832 5590 2194
rect 163 1548 5588 1832
rect 163 1544 2483 1548
rect 5236 1529 5588 1548
<< pwell >>
rect 3584 41433 3840 41445
rect 1153 41429 5121 41433
rect 173 41369 5121 41429
rect 173 41368 5394 41369
rect 173 41306 5508 41368
rect 173 41182 5509 41306
rect 173 41148 5521 41182
rect 173 41045 5509 41148
rect 173 41041 3840 41045
rect 173 40987 1447 41041
rect 2326 40991 3840 41041
rect 3847 40992 5509 41045
rect 3847 40991 5121 40992
rect 3584 40981 3840 40991
rect 3584 40146 3840 40158
rect 1153 40142 5121 40146
rect 173 40082 5121 40142
rect 173 40081 5394 40082
rect 173 40019 5508 40081
rect 173 39895 5509 40019
rect 173 39861 5521 39895
rect 173 39758 5509 39861
rect 173 39754 3840 39758
rect 173 39700 1447 39754
rect 2326 39704 3840 39754
rect 3847 39705 5509 39758
rect 3847 39704 5121 39705
rect 3584 39694 3840 39704
rect 3584 38859 3840 38871
rect 1153 38855 5121 38859
rect 173 38795 5121 38855
rect 173 38794 5394 38795
rect 173 38732 5508 38794
rect 173 38608 5509 38732
rect 173 38574 5521 38608
rect 173 38471 5509 38574
rect 173 38467 3840 38471
rect 173 38413 1447 38467
rect 2326 38417 3840 38467
rect 3847 38418 5509 38471
rect 3847 38417 5121 38418
rect 3584 38407 3840 38417
rect 3584 37572 3840 37584
rect 1153 37568 5121 37572
rect 173 37508 5121 37568
rect 173 37507 5394 37508
rect 173 37445 5508 37507
rect 173 37321 5509 37445
rect 173 37287 5521 37321
rect 173 37184 5509 37287
rect 173 37180 3840 37184
rect 173 37126 1447 37180
rect 2326 37130 3840 37180
rect 3847 37131 5509 37184
rect 3847 37130 5121 37131
rect 3584 37120 3840 37130
rect 3584 36285 3840 36297
rect 1153 36281 5121 36285
rect 173 36221 5121 36281
rect 173 36220 5394 36221
rect 173 36158 5508 36220
rect 173 36034 5509 36158
rect 173 36000 5521 36034
rect 173 35897 5509 36000
rect 173 35893 3840 35897
rect 173 35839 1447 35893
rect 2326 35843 3840 35893
rect 3847 35844 5509 35897
rect 3847 35843 5121 35844
rect 3584 35833 3840 35843
rect 3584 34998 3840 35010
rect 1153 34994 5121 34998
rect 173 34934 5121 34994
rect 173 34933 5394 34934
rect 173 34871 5508 34933
rect 173 34747 5509 34871
rect 173 34713 5521 34747
rect 173 34610 5509 34713
rect 173 34606 3840 34610
rect 173 34552 1447 34606
rect 2326 34556 3840 34606
rect 3847 34557 5509 34610
rect 3847 34556 5121 34557
rect 3584 34546 3840 34556
rect 3584 33711 3840 33723
rect 1153 33707 5121 33711
rect 173 33647 5121 33707
rect 173 33646 5394 33647
rect 173 33584 5508 33646
rect 173 33460 5509 33584
rect 173 33426 5521 33460
rect 173 33323 5509 33426
rect 173 33319 3840 33323
rect 173 33265 1447 33319
rect 2326 33269 3840 33319
rect 3847 33270 5509 33323
rect 3847 33269 5121 33270
rect 3584 33259 3840 33269
rect 3584 32424 3840 32436
rect 1153 32420 5121 32424
rect 173 32360 5121 32420
rect 173 32359 5394 32360
rect 173 32297 5508 32359
rect 173 32173 5509 32297
rect 173 32139 5521 32173
rect 173 32036 5509 32139
rect 173 32032 3840 32036
rect 173 31978 1447 32032
rect 2326 31982 3840 32032
rect 3847 31983 5509 32036
rect 3847 31982 5121 31983
rect 3584 31972 3840 31982
rect 3584 31137 3840 31149
rect 1153 31133 5121 31137
rect 173 31073 5121 31133
rect 173 31072 5394 31073
rect 173 31010 5508 31072
rect 173 30886 5509 31010
rect 173 30852 5521 30886
rect 173 30749 5509 30852
rect 173 30745 3840 30749
rect 173 30691 1447 30745
rect 2326 30695 3840 30745
rect 3847 30696 5509 30749
rect 3847 30695 5121 30696
rect 3584 30685 3840 30695
rect 3584 29850 3840 29862
rect 1153 29846 5121 29850
rect 173 29786 5121 29846
rect 173 29785 5394 29786
rect 173 29723 5508 29785
rect 173 29599 5509 29723
rect 173 29565 5521 29599
rect 173 29462 5509 29565
rect 173 29458 3840 29462
rect 173 29404 1447 29458
rect 2326 29408 3840 29458
rect 3847 29409 5509 29462
rect 3847 29408 5121 29409
rect 3584 29398 3840 29408
rect 3584 28563 3840 28575
rect 1153 28559 5121 28563
rect 173 28499 5121 28559
rect 173 28498 5394 28499
rect 173 28436 5508 28498
rect 173 28312 5509 28436
rect 173 28278 5521 28312
rect 173 28175 5509 28278
rect 173 28171 3840 28175
rect 173 28117 1447 28171
rect 2326 28121 3840 28171
rect 3847 28122 5509 28175
rect 3847 28121 5121 28122
rect 3584 28111 3840 28121
rect 3584 27276 3840 27288
rect 1153 27272 5121 27276
rect 173 27212 5121 27272
rect 173 27211 5394 27212
rect 173 27149 5508 27211
rect 173 27025 5509 27149
rect 173 26991 5521 27025
rect 173 26888 5509 26991
rect 173 26884 3840 26888
rect 173 26830 1447 26884
rect 2326 26834 3840 26884
rect 3847 26835 5509 26888
rect 3847 26834 5121 26835
rect 3584 26824 3840 26834
rect 3584 25989 3840 26001
rect 1153 25985 5121 25989
rect 173 25925 5121 25985
rect 173 25924 5394 25925
rect 173 25862 5508 25924
rect 173 25738 5509 25862
rect 173 25704 5521 25738
rect 173 25601 5509 25704
rect 173 25597 3840 25601
rect 173 25543 1447 25597
rect 2326 25547 3840 25597
rect 3847 25548 5509 25601
rect 3847 25547 5121 25548
rect 3584 25537 3840 25547
rect 3584 24702 3840 24714
rect 1153 24698 5121 24702
rect 173 24638 5121 24698
rect 173 24637 5394 24638
rect 173 24575 5508 24637
rect 173 24451 5509 24575
rect 173 24417 5521 24451
rect 173 24314 5509 24417
rect 173 24310 3840 24314
rect 173 24256 1447 24310
rect 2326 24260 3840 24310
rect 3847 24261 5509 24314
rect 3847 24260 5121 24261
rect 3584 24250 3840 24260
rect 3584 23415 3840 23427
rect 1153 23411 5121 23415
rect 173 23351 5121 23411
rect 173 23350 5394 23351
rect 173 23288 5508 23350
rect 173 23164 5509 23288
rect 173 23130 5521 23164
rect 173 23027 5509 23130
rect 173 23023 3840 23027
rect 173 22969 1447 23023
rect 2326 22973 3840 23023
rect 3847 22974 5509 23027
rect 3847 22973 5121 22974
rect 3584 22963 3840 22973
rect 3584 22128 3840 22140
rect 1153 22124 5121 22128
rect 173 22064 5121 22124
rect 173 22063 5394 22064
rect 173 22001 5508 22063
rect 173 21877 5509 22001
rect 173 21843 5521 21877
rect 173 21740 5509 21843
rect 173 21736 3840 21740
rect 173 21682 1447 21736
rect 2326 21686 3840 21736
rect 3847 21687 5509 21740
rect 3847 21686 5121 21687
rect 3584 21676 3840 21686
rect 3584 20841 3840 20853
rect 1153 20837 5121 20841
rect 173 20777 5121 20837
rect 173 20776 5394 20777
rect 173 20714 5508 20776
rect 173 20590 5509 20714
rect 173 20556 5521 20590
rect 173 20453 5509 20556
rect 173 20449 3840 20453
rect 173 20395 1447 20449
rect 2326 20399 3840 20449
rect 3847 20400 5509 20453
rect 3847 20399 5121 20400
rect 3584 20389 3840 20399
rect 3584 19554 3840 19566
rect 1153 19550 5121 19554
rect 173 19490 5121 19550
rect 173 19489 5394 19490
rect 173 19427 5508 19489
rect 173 19303 5509 19427
rect 173 19269 5521 19303
rect 173 19166 5509 19269
rect 173 19162 3840 19166
rect 173 19108 1447 19162
rect 2326 19112 3840 19162
rect 3847 19113 5509 19166
rect 3847 19112 5121 19113
rect 3584 19102 3840 19112
rect 3584 18267 3840 18279
rect 1153 18263 5121 18267
rect 173 18203 5121 18263
rect 173 18202 5394 18203
rect 173 18140 5508 18202
rect 173 18016 5509 18140
rect 173 17982 5521 18016
rect 173 17879 5509 17982
rect 173 17875 3840 17879
rect 173 17821 1447 17875
rect 2326 17825 3840 17875
rect 3847 17826 5509 17879
rect 3847 17825 5121 17826
rect 3584 17815 3840 17825
rect 3584 16980 3840 16992
rect 1153 16976 5121 16980
rect 173 16916 5121 16976
rect 173 16915 5394 16916
rect 173 16853 5508 16915
rect 173 16729 5509 16853
rect 173 16695 5521 16729
rect 173 16592 5509 16695
rect 173 16588 3840 16592
rect 173 16534 1447 16588
rect 2326 16538 3840 16588
rect 3847 16539 5509 16592
rect 3847 16538 5121 16539
rect 3584 16528 3840 16538
rect 3584 15693 3840 15705
rect 1153 15689 5121 15693
rect 173 15629 5121 15689
rect 173 15628 5394 15629
rect 173 15566 5508 15628
rect 173 15442 5509 15566
rect 173 15408 5521 15442
rect 173 15305 5509 15408
rect 173 15301 3840 15305
rect 173 15247 1447 15301
rect 2326 15251 3840 15301
rect 3847 15252 5509 15305
rect 3847 15251 5121 15252
rect 3584 15241 3840 15251
rect 3584 14406 3840 14418
rect 1153 14402 5121 14406
rect 173 14342 5121 14402
rect 173 14341 5394 14342
rect 173 14279 5508 14341
rect 173 14155 5509 14279
rect 173 14121 5521 14155
rect 173 14018 5509 14121
rect 173 14014 3840 14018
rect 173 13960 1447 14014
rect 2326 13964 3840 14014
rect 3847 13965 5509 14018
rect 3847 13964 5121 13965
rect 3584 13954 3840 13964
rect 3584 13119 3840 13131
rect 1153 13115 5121 13119
rect 173 13055 5121 13115
rect 173 13054 5394 13055
rect 173 12992 5508 13054
rect 173 12868 5509 12992
rect 173 12834 5521 12868
rect 173 12731 5509 12834
rect 173 12727 3840 12731
rect 173 12673 1447 12727
rect 2326 12677 3840 12727
rect 3847 12678 5509 12731
rect 3847 12677 5121 12678
rect 3584 12667 3840 12677
rect 3584 11832 3840 11844
rect 1153 11828 5121 11832
rect 173 11768 5121 11828
rect 173 11767 5394 11768
rect 173 11705 5508 11767
rect 173 11581 5509 11705
rect 173 11547 5521 11581
rect 173 11444 5509 11547
rect 173 11440 3840 11444
rect 173 11386 1447 11440
rect 2326 11390 3840 11440
rect 3847 11391 5509 11444
rect 3847 11390 5121 11391
rect 3584 11380 3840 11390
rect 3584 10545 3840 10557
rect 1153 10541 5121 10545
rect 173 10481 5121 10541
rect 173 10480 5394 10481
rect 173 10418 5508 10480
rect 173 10294 5509 10418
rect 173 10260 5521 10294
rect 173 10157 5509 10260
rect 173 10153 3840 10157
rect 173 10099 1447 10153
rect 2326 10103 3840 10153
rect 3847 10104 5509 10157
rect 3847 10103 5121 10104
rect 3584 10093 3840 10103
rect 3584 9258 3840 9270
rect 1153 9254 5121 9258
rect 173 9194 5121 9254
rect 173 9193 5394 9194
rect 173 9131 5508 9193
rect 173 9007 5509 9131
rect 173 8973 5521 9007
rect 173 8870 5509 8973
rect 173 8866 3840 8870
rect 173 8812 1447 8866
rect 2326 8816 3840 8866
rect 3847 8817 5509 8870
rect 3847 8816 5121 8817
rect 3584 8806 3840 8816
rect 3584 7971 3840 7983
rect 1153 7967 5121 7971
rect 173 7907 5121 7967
rect 173 7906 5394 7907
rect 173 7844 5508 7906
rect 173 7720 5509 7844
rect 173 7686 5521 7720
rect 173 7583 5509 7686
rect 173 7579 3840 7583
rect 173 7525 1447 7579
rect 2326 7529 3840 7579
rect 3847 7530 5509 7583
rect 3847 7529 5121 7530
rect 3584 7519 3840 7529
rect 3584 6684 3840 6696
rect 1153 6680 5121 6684
rect 173 6620 5121 6680
rect 173 6619 5394 6620
rect 173 6557 5508 6619
rect 173 6433 5509 6557
rect 173 6399 5521 6433
rect 173 6296 5509 6399
rect 173 6292 3840 6296
rect 173 6238 1447 6292
rect 2326 6242 3840 6292
rect 3847 6243 5509 6296
rect 3847 6242 5121 6243
rect 3584 6232 3840 6242
rect 3584 5397 3840 5409
rect 1153 5393 5121 5397
rect 173 5333 5121 5393
rect 173 5332 5394 5333
rect 173 5270 5508 5332
rect 173 5146 5509 5270
rect 173 5112 5521 5146
rect 173 5009 5509 5112
rect 173 5005 3840 5009
rect 173 4951 1447 5005
rect 2326 4955 3840 5005
rect 3847 4956 5509 5009
rect 3847 4955 5121 4956
rect 3584 4945 3840 4955
rect 3584 4110 3840 4122
rect 1153 4106 5121 4110
rect 173 4046 5121 4106
rect 173 4045 5394 4046
rect 173 3983 5508 4045
rect 173 3859 5509 3983
rect 173 3825 5521 3859
rect 173 3722 5509 3825
rect 173 3718 3840 3722
rect 173 3664 1447 3718
rect 2326 3668 3840 3718
rect 3847 3669 5509 3722
rect 3847 3668 5121 3669
rect 3584 3658 3840 3668
rect 3584 2823 3840 2835
rect 1153 2819 5121 2823
rect 173 2759 5121 2819
rect 173 2758 5394 2759
rect 173 2696 5508 2758
rect 173 2572 5509 2696
rect 173 2538 5521 2572
rect 173 2435 5509 2538
rect 173 2431 3840 2435
rect 173 2377 1447 2431
rect 2326 2381 3840 2431
rect 3847 2382 5509 2435
rect 3847 2381 5121 2382
rect 3584 2371 3840 2381
rect 3584 1536 3840 1548
rect 1153 1532 5121 1536
rect 173 1472 5121 1532
rect 173 1471 5394 1472
rect 173 1409 5508 1471
rect 173 1285 5509 1409
rect 173 1251 5521 1285
rect 173 1148 5509 1251
rect 173 1144 3840 1148
rect 173 1090 1447 1144
rect 2326 1094 3840 1144
rect 3847 1095 5509 1148
rect 3847 1094 5121 1095
rect 3584 1084 3840 1094
<< nmos >>
rect 363 41187 393 41291
rect 459 41187 489 41291
rect 555 41187 585 41291
rect 651 41187 681 41291
rect 747 41187 777 41291
rect 843 41187 873 41291
rect 939 41187 969 41291
rect 1035 41187 1065 41291
rect 1131 41187 1161 41291
rect 1227 41187 1257 41291
rect 2516 41191 2546 41295
rect 2612 41191 2642 41295
rect 2708 41191 2738 41295
rect 2804 41191 2834 41295
rect 2900 41191 2930 41295
rect 2996 41191 3026 41295
rect 3092 41191 3122 41295
rect 3188 41191 3218 41295
rect 3284 41191 3314 41295
rect 3380 41191 3410 41295
rect 3693 41199 3723 41299
rect 4037 41191 4067 41295
rect 4133 41191 4163 41295
rect 4229 41191 4259 41295
rect 4325 41191 4355 41295
rect 4421 41191 4451 41295
rect 4517 41191 4547 41295
rect 4613 41191 4643 41295
rect 4709 41191 4739 41295
rect 4805 41191 4835 41295
rect 4901 41191 4931 41295
rect 363 39900 393 40004
rect 459 39900 489 40004
rect 555 39900 585 40004
rect 651 39900 681 40004
rect 747 39900 777 40004
rect 843 39900 873 40004
rect 939 39900 969 40004
rect 1035 39900 1065 40004
rect 1131 39900 1161 40004
rect 1227 39900 1257 40004
rect 2516 39904 2546 40008
rect 2612 39904 2642 40008
rect 2708 39904 2738 40008
rect 2804 39904 2834 40008
rect 2900 39904 2930 40008
rect 2996 39904 3026 40008
rect 3092 39904 3122 40008
rect 3188 39904 3218 40008
rect 3284 39904 3314 40008
rect 3380 39904 3410 40008
rect 3693 39912 3723 40012
rect 4037 39904 4067 40008
rect 4133 39904 4163 40008
rect 4229 39904 4259 40008
rect 4325 39904 4355 40008
rect 4421 39904 4451 40008
rect 4517 39904 4547 40008
rect 4613 39904 4643 40008
rect 4709 39904 4739 40008
rect 4805 39904 4835 40008
rect 4901 39904 4931 40008
rect 363 38613 393 38717
rect 459 38613 489 38717
rect 555 38613 585 38717
rect 651 38613 681 38717
rect 747 38613 777 38717
rect 843 38613 873 38717
rect 939 38613 969 38717
rect 1035 38613 1065 38717
rect 1131 38613 1161 38717
rect 1227 38613 1257 38717
rect 2516 38617 2546 38721
rect 2612 38617 2642 38721
rect 2708 38617 2738 38721
rect 2804 38617 2834 38721
rect 2900 38617 2930 38721
rect 2996 38617 3026 38721
rect 3092 38617 3122 38721
rect 3188 38617 3218 38721
rect 3284 38617 3314 38721
rect 3380 38617 3410 38721
rect 3693 38625 3723 38725
rect 4037 38617 4067 38721
rect 4133 38617 4163 38721
rect 4229 38617 4259 38721
rect 4325 38617 4355 38721
rect 4421 38617 4451 38721
rect 4517 38617 4547 38721
rect 4613 38617 4643 38721
rect 4709 38617 4739 38721
rect 4805 38617 4835 38721
rect 4901 38617 4931 38721
rect 363 37326 393 37430
rect 459 37326 489 37430
rect 555 37326 585 37430
rect 651 37326 681 37430
rect 747 37326 777 37430
rect 843 37326 873 37430
rect 939 37326 969 37430
rect 1035 37326 1065 37430
rect 1131 37326 1161 37430
rect 1227 37326 1257 37430
rect 2516 37330 2546 37434
rect 2612 37330 2642 37434
rect 2708 37330 2738 37434
rect 2804 37330 2834 37434
rect 2900 37330 2930 37434
rect 2996 37330 3026 37434
rect 3092 37330 3122 37434
rect 3188 37330 3218 37434
rect 3284 37330 3314 37434
rect 3380 37330 3410 37434
rect 3693 37338 3723 37438
rect 4037 37330 4067 37434
rect 4133 37330 4163 37434
rect 4229 37330 4259 37434
rect 4325 37330 4355 37434
rect 4421 37330 4451 37434
rect 4517 37330 4547 37434
rect 4613 37330 4643 37434
rect 4709 37330 4739 37434
rect 4805 37330 4835 37434
rect 4901 37330 4931 37434
rect 363 36039 393 36143
rect 459 36039 489 36143
rect 555 36039 585 36143
rect 651 36039 681 36143
rect 747 36039 777 36143
rect 843 36039 873 36143
rect 939 36039 969 36143
rect 1035 36039 1065 36143
rect 1131 36039 1161 36143
rect 1227 36039 1257 36143
rect 2516 36043 2546 36147
rect 2612 36043 2642 36147
rect 2708 36043 2738 36147
rect 2804 36043 2834 36147
rect 2900 36043 2930 36147
rect 2996 36043 3026 36147
rect 3092 36043 3122 36147
rect 3188 36043 3218 36147
rect 3284 36043 3314 36147
rect 3380 36043 3410 36147
rect 3693 36051 3723 36151
rect 4037 36043 4067 36147
rect 4133 36043 4163 36147
rect 4229 36043 4259 36147
rect 4325 36043 4355 36147
rect 4421 36043 4451 36147
rect 4517 36043 4547 36147
rect 4613 36043 4643 36147
rect 4709 36043 4739 36147
rect 4805 36043 4835 36147
rect 4901 36043 4931 36147
rect 363 34752 393 34856
rect 459 34752 489 34856
rect 555 34752 585 34856
rect 651 34752 681 34856
rect 747 34752 777 34856
rect 843 34752 873 34856
rect 939 34752 969 34856
rect 1035 34752 1065 34856
rect 1131 34752 1161 34856
rect 1227 34752 1257 34856
rect 2516 34756 2546 34860
rect 2612 34756 2642 34860
rect 2708 34756 2738 34860
rect 2804 34756 2834 34860
rect 2900 34756 2930 34860
rect 2996 34756 3026 34860
rect 3092 34756 3122 34860
rect 3188 34756 3218 34860
rect 3284 34756 3314 34860
rect 3380 34756 3410 34860
rect 3693 34764 3723 34864
rect 4037 34756 4067 34860
rect 4133 34756 4163 34860
rect 4229 34756 4259 34860
rect 4325 34756 4355 34860
rect 4421 34756 4451 34860
rect 4517 34756 4547 34860
rect 4613 34756 4643 34860
rect 4709 34756 4739 34860
rect 4805 34756 4835 34860
rect 4901 34756 4931 34860
rect 363 33465 393 33569
rect 459 33465 489 33569
rect 555 33465 585 33569
rect 651 33465 681 33569
rect 747 33465 777 33569
rect 843 33465 873 33569
rect 939 33465 969 33569
rect 1035 33465 1065 33569
rect 1131 33465 1161 33569
rect 1227 33465 1257 33569
rect 2516 33469 2546 33573
rect 2612 33469 2642 33573
rect 2708 33469 2738 33573
rect 2804 33469 2834 33573
rect 2900 33469 2930 33573
rect 2996 33469 3026 33573
rect 3092 33469 3122 33573
rect 3188 33469 3218 33573
rect 3284 33469 3314 33573
rect 3380 33469 3410 33573
rect 3693 33477 3723 33577
rect 4037 33469 4067 33573
rect 4133 33469 4163 33573
rect 4229 33469 4259 33573
rect 4325 33469 4355 33573
rect 4421 33469 4451 33573
rect 4517 33469 4547 33573
rect 4613 33469 4643 33573
rect 4709 33469 4739 33573
rect 4805 33469 4835 33573
rect 4901 33469 4931 33573
rect 363 32178 393 32282
rect 459 32178 489 32282
rect 555 32178 585 32282
rect 651 32178 681 32282
rect 747 32178 777 32282
rect 843 32178 873 32282
rect 939 32178 969 32282
rect 1035 32178 1065 32282
rect 1131 32178 1161 32282
rect 1227 32178 1257 32282
rect 2516 32182 2546 32286
rect 2612 32182 2642 32286
rect 2708 32182 2738 32286
rect 2804 32182 2834 32286
rect 2900 32182 2930 32286
rect 2996 32182 3026 32286
rect 3092 32182 3122 32286
rect 3188 32182 3218 32286
rect 3284 32182 3314 32286
rect 3380 32182 3410 32286
rect 3693 32190 3723 32290
rect 4037 32182 4067 32286
rect 4133 32182 4163 32286
rect 4229 32182 4259 32286
rect 4325 32182 4355 32286
rect 4421 32182 4451 32286
rect 4517 32182 4547 32286
rect 4613 32182 4643 32286
rect 4709 32182 4739 32286
rect 4805 32182 4835 32286
rect 4901 32182 4931 32286
rect 363 30891 393 30995
rect 459 30891 489 30995
rect 555 30891 585 30995
rect 651 30891 681 30995
rect 747 30891 777 30995
rect 843 30891 873 30995
rect 939 30891 969 30995
rect 1035 30891 1065 30995
rect 1131 30891 1161 30995
rect 1227 30891 1257 30995
rect 2516 30895 2546 30999
rect 2612 30895 2642 30999
rect 2708 30895 2738 30999
rect 2804 30895 2834 30999
rect 2900 30895 2930 30999
rect 2996 30895 3026 30999
rect 3092 30895 3122 30999
rect 3188 30895 3218 30999
rect 3284 30895 3314 30999
rect 3380 30895 3410 30999
rect 3693 30903 3723 31003
rect 4037 30895 4067 30999
rect 4133 30895 4163 30999
rect 4229 30895 4259 30999
rect 4325 30895 4355 30999
rect 4421 30895 4451 30999
rect 4517 30895 4547 30999
rect 4613 30895 4643 30999
rect 4709 30895 4739 30999
rect 4805 30895 4835 30999
rect 4901 30895 4931 30999
rect 363 29604 393 29708
rect 459 29604 489 29708
rect 555 29604 585 29708
rect 651 29604 681 29708
rect 747 29604 777 29708
rect 843 29604 873 29708
rect 939 29604 969 29708
rect 1035 29604 1065 29708
rect 1131 29604 1161 29708
rect 1227 29604 1257 29708
rect 2516 29608 2546 29712
rect 2612 29608 2642 29712
rect 2708 29608 2738 29712
rect 2804 29608 2834 29712
rect 2900 29608 2930 29712
rect 2996 29608 3026 29712
rect 3092 29608 3122 29712
rect 3188 29608 3218 29712
rect 3284 29608 3314 29712
rect 3380 29608 3410 29712
rect 3693 29616 3723 29716
rect 4037 29608 4067 29712
rect 4133 29608 4163 29712
rect 4229 29608 4259 29712
rect 4325 29608 4355 29712
rect 4421 29608 4451 29712
rect 4517 29608 4547 29712
rect 4613 29608 4643 29712
rect 4709 29608 4739 29712
rect 4805 29608 4835 29712
rect 4901 29608 4931 29712
rect 363 28317 393 28421
rect 459 28317 489 28421
rect 555 28317 585 28421
rect 651 28317 681 28421
rect 747 28317 777 28421
rect 843 28317 873 28421
rect 939 28317 969 28421
rect 1035 28317 1065 28421
rect 1131 28317 1161 28421
rect 1227 28317 1257 28421
rect 2516 28321 2546 28425
rect 2612 28321 2642 28425
rect 2708 28321 2738 28425
rect 2804 28321 2834 28425
rect 2900 28321 2930 28425
rect 2996 28321 3026 28425
rect 3092 28321 3122 28425
rect 3188 28321 3218 28425
rect 3284 28321 3314 28425
rect 3380 28321 3410 28425
rect 3693 28329 3723 28429
rect 4037 28321 4067 28425
rect 4133 28321 4163 28425
rect 4229 28321 4259 28425
rect 4325 28321 4355 28425
rect 4421 28321 4451 28425
rect 4517 28321 4547 28425
rect 4613 28321 4643 28425
rect 4709 28321 4739 28425
rect 4805 28321 4835 28425
rect 4901 28321 4931 28425
rect 363 27030 393 27134
rect 459 27030 489 27134
rect 555 27030 585 27134
rect 651 27030 681 27134
rect 747 27030 777 27134
rect 843 27030 873 27134
rect 939 27030 969 27134
rect 1035 27030 1065 27134
rect 1131 27030 1161 27134
rect 1227 27030 1257 27134
rect 2516 27034 2546 27138
rect 2612 27034 2642 27138
rect 2708 27034 2738 27138
rect 2804 27034 2834 27138
rect 2900 27034 2930 27138
rect 2996 27034 3026 27138
rect 3092 27034 3122 27138
rect 3188 27034 3218 27138
rect 3284 27034 3314 27138
rect 3380 27034 3410 27138
rect 3693 27042 3723 27142
rect 4037 27034 4067 27138
rect 4133 27034 4163 27138
rect 4229 27034 4259 27138
rect 4325 27034 4355 27138
rect 4421 27034 4451 27138
rect 4517 27034 4547 27138
rect 4613 27034 4643 27138
rect 4709 27034 4739 27138
rect 4805 27034 4835 27138
rect 4901 27034 4931 27138
rect 363 25743 393 25847
rect 459 25743 489 25847
rect 555 25743 585 25847
rect 651 25743 681 25847
rect 747 25743 777 25847
rect 843 25743 873 25847
rect 939 25743 969 25847
rect 1035 25743 1065 25847
rect 1131 25743 1161 25847
rect 1227 25743 1257 25847
rect 2516 25747 2546 25851
rect 2612 25747 2642 25851
rect 2708 25747 2738 25851
rect 2804 25747 2834 25851
rect 2900 25747 2930 25851
rect 2996 25747 3026 25851
rect 3092 25747 3122 25851
rect 3188 25747 3218 25851
rect 3284 25747 3314 25851
rect 3380 25747 3410 25851
rect 3693 25755 3723 25855
rect 4037 25747 4067 25851
rect 4133 25747 4163 25851
rect 4229 25747 4259 25851
rect 4325 25747 4355 25851
rect 4421 25747 4451 25851
rect 4517 25747 4547 25851
rect 4613 25747 4643 25851
rect 4709 25747 4739 25851
rect 4805 25747 4835 25851
rect 4901 25747 4931 25851
rect 363 24456 393 24560
rect 459 24456 489 24560
rect 555 24456 585 24560
rect 651 24456 681 24560
rect 747 24456 777 24560
rect 843 24456 873 24560
rect 939 24456 969 24560
rect 1035 24456 1065 24560
rect 1131 24456 1161 24560
rect 1227 24456 1257 24560
rect 2516 24460 2546 24564
rect 2612 24460 2642 24564
rect 2708 24460 2738 24564
rect 2804 24460 2834 24564
rect 2900 24460 2930 24564
rect 2996 24460 3026 24564
rect 3092 24460 3122 24564
rect 3188 24460 3218 24564
rect 3284 24460 3314 24564
rect 3380 24460 3410 24564
rect 3693 24468 3723 24568
rect 4037 24460 4067 24564
rect 4133 24460 4163 24564
rect 4229 24460 4259 24564
rect 4325 24460 4355 24564
rect 4421 24460 4451 24564
rect 4517 24460 4547 24564
rect 4613 24460 4643 24564
rect 4709 24460 4739 24564
rect 4805 24460 4835 24564
rect 4901 24460 4931 24564
rect 363 23169 393 23273
rect 459 23169 489 23273
rect 555 23169 585 23273
rect 651 23169 681 23273
rect 747 23169 777 23273
rect 843 23169 873 23273
rect 939 23169 969 23273
rect 1035 23169 1065 23273
rect 1131 23169 1161 23273
rect 1227 23169 1257 23273
rect 2516 23173 2546 23277
rect 2612 23173 2642 23277
rect 2708 23173 2738 23277
rect 2804 23173 2834 23277
rect 2900 23173 2930 23277
rect 2996 23173 3026 23277
rect 3092 23173 3122 23277
rect 3188 23173 3218 23277
rect 3284 23173 3314 23277
rect 3380 23173 3410 23277
rect 3693 23181 3723 23281
rect 4037 23173 4067 23277
rect 4133 23173 4163 23277
rect 4229 23173 4259 23277
rect 4325 23173 4355 23277
rect 4421 23173 4451 23277
rect 4517 23173 4547 23277
rect 4613 23173 4643 23277
rect 4709 23173 4739 23277
rect 4805 23173 4835 23277
rect 4901 23173 4931 23277
rect 363 21882 393 21986
rect 459 21882 489 21986
rect 555 21882 585 21986
rect 651 21882 681 21986
rect 747 21882 777 21986
rect 843 21882 873 21986
rect 939 21882 969 21986
rect 1035 21882 1065 21986
rect 1131 21882 1161 21986
rect 1227 21882 1257 21986
rect 2516 21886 2546 21990
rect 2612 21886 2642 21990
rect 2708 21886 2738 21990
rect 2804 21886 2834 21990
rect 2900 21886 2930 21990
rect 2996 21886 3026 21990
rect 3092 21886 3122 21990
rect 3188 21886 3218 21990
rect 3284 21886 3314 21990
rect 3380 21886 3410 21990
rect 3693 21894 3723 21994
rect 4037 21886 4067 21990
rect 4133 21886 4163 21990
rect 4229 21886 4259 21990
rect 4325 21886 4355 21990
rect 4421 21886 4451 21990
rect 4517 21886 4547 21990
rect 4613 21886 4643 21990
rect 4709 21886 4739 21990
rect 4805 21886 4835 21990
rect 4901 21886 4931 21990
rect 363 20595 393 20699
rect 459 20595 489 20699
rect 555 20595 585 20699
rect 651 20595 681 20699
rect 747 20595 777 20699
rect 843 20595 873 20699
rect 939 20595 969 20699
rect 1035 20595 1065 20699
rect 1131 20595 1161 20699
rect 1227 20595 1257 20699
rect 2516 20599 2546 20703
rect 2612 20599 2642 20703
rect 2708 20599 2738 20703
rect 2804 20599 2834 20703
rect 2900 20599 2930 20703
rect 2996 20599 3026 20703
rect 3092 20599 3122 20703
rect 3188 20599 3218 20703
rect 3284 20599 3314 20703
rect 3380 20599 3410 20703
rect 3693 20607 3723 20707
rect 4037 20599 4067 20703
rect 4133 20599 4163 20703
rect 4229 20599 4259 20703
rect 4325 20599 4355 20703
rect 4421 20599 4451 20703
rect 4517 20599 4547 20703
rect 4613 20599 4643 20703
rect 4709 20599 4739 20703
rect 4805 20599 4835 20703
rect 4901 20599 4931 20703
rect 363 19308 393 19412
rect 459 19308 489 19412
rect 555 19308 585 19412
rect 651 19308 681 19412
rect 747 19308 777 19412
rect 843 19308 873 19412
rect 939 19308 969 19412
rect 1035 19308 1065 19412
rect 1131 19308 1161 19412
rect 1227 19308 1257 19412
rect 2516 19312 2546 19416
rect 2612 19312 2642 19416
rect 2708 19312 2738 19416
rect 2804 19312 2834 19416
rect 2900 19312 2930 19416
rect 2996 19312 3026 19416
rect 3092 19312 3122 19416
rect 3188 19312 3218 19416
rect 3284 19312 3314 19416
rect 3380 19312 3410 19416
rect 3693 19320 3723 19420
rect 4037 19312 4067 19416
rect 4133 19312 4163 19416
rect 4229 19312 4259 19416
rect 4325 19312 4355 19416
rect 4421 19312 4451 19416
rect 4517 19312 4547 19416
rect 4613 19312 4643 19416
rect 4709 19312 4739 19416
rect 4805 19312 4835 19416
rect 4901 19312 4931 19416
rect 363 18021 393 18125
rect 459 18021 489 18125
rect 555 18021 585 18125
rect 651 18021 681 18125
rect 747 18021 777 18125
rect 843 18021 873 18125
rect 939 18021 969 18125
rect 1035 18021 1065 18125
rect 1131 18021 1161 18125
rect 1227 18021 1257 18125
rect 2516 18025 2546 18129
rect 2612 18025 2642 18129
rect 2708 18025 2738 18129
rect 2804 18025 2834 18129
rect 2900 18025 2930 18129
rect 2996 18025 3026 18129
rect 3092 18025 3122 18129
rect 3188 18025 3218 18129
rect 3284 18025 3314 18129
rect 3380 18025 3410 18129
rect 3693 18033 3723 18133
rect 4037 18025 4067 18129
rect 4133 18025 4163 18129
rect 4229 18025 4259 18129
rect 4325 18025 4355 18129
rect 4421 18025 4451 18129
rect 4517 18025 4547 18129
rect 4613 18025 4643 18129
rect 4709 18025 4739 18129
rect 4805 18025 4835 18129
rect 4901 18025 4931 18129
rect 363 16734 393 16838
rect 459 16734 489 16838
rect 555 16734 585 16838
rect 651 16734 681 16838
rect 747 16734 777 16838
rect 843 16734 873 16838
rect 939 16734 969 16838
rect 1035 16734 1065 16838
rect 1131 16734 1161 16838
rect 1227 16734 1257 16838
rect 2516 16738 2546 16842
rect 2612 16738 2642 16842
rect 2708 16738 2738 16842
rect 2804 16738 2834 16842
rect 2900 16738 2930 16842
rect 2996 16738 3026 16842
rect 3092 16738 3122 16842
rect 3188 16738 3218 16842
rect 3284 16738 3314 16842
rect 3380 16738 3410 16842
rect 3693 16746 3723 16846
rect 4037 16738 4067 16842
rect 4133 16738 4163 16842
rect 4229 16738 4259 16842
rect 4325 16738 4355 16842
rect 4421 16738 4451 16842
rect 4517 16738 4547 16842
rect 4613 16738 4643 16842
rect 4709 16738 4739 16842
rect 4805 16738 4835 16842
rect 4901 16738 4931 16842
rect 363 15447 393 15551
rect 459 15447 489 15551
rect 555 15447 585 15551
rect 651 15447 681 15551
rect 747 15447 777 15551
rect 843 15447 873 15551
rect 939 15447 969 15551
rect 1035 15447 1065 15551
rect 1131 15447 1161 15551
rect 1227 15447 1257 15551
rect 2516 15451 2546 15555
rect 2612 15451 2642 15555
rect 2708 15451 2738 15555
rect 2804 15451 2834 15555
rect 2900 15451 2930 15555
rect 2996 15451 3026 15555
rect 3092 15451 3122 15555
rect 3188 15451 3218 15555
rect 3284 15451 3314 15555
rect 3380 15451 3410 15555
rect 3693 15459 3723 15559
rect 4037 15451 4067 15555
rect 4133 15451 4163 15555
rect 4229 15451 4259 15555
rect 4325 15451 4355 15555
rect 4421 15451 4451 15555
rect 4517 15451 4547 15555
rect 4613 15451 4643 15555
rect 4709 15451 4739 15555
rect 4805 15451 4835 15555
rect 4901 15451 4931 15555
rect 363 14160 393 14264
rect 459 14160 489 14264
rect 555 14160 585 14264
rect 651 14160 681 14264
rect 747 14160 777 14264
rect 843 14160 873 14264
rect 939 14160 969 14264
rect 1035 14160 1065 14264
rect 1131 14160 1161 14264
rect 1227 14160 1257 14264
rect 2516 14164 2546 14268
rect 2612 14164 2642 14268
rect 2708 14164 2738 14268
rect 2804 14164 2834 14268
rect 2900 14164 2930 14268
rect 2996 14164 3026 14268
rect 3092 14164 3122 14268
rect 3188 14164 3218 14268
rect 3284 14164 3314 14268
rect 3380 14164 3410 14268
rect 3693 14172 3723 14272
rect 4037 14164 4067 14268
rect 4133 14164 4163 14268
rect 4229 14164 4259 14268
rect 4325 14164 4355 14268
rect 4421 14164 4451 14268
rect 4517 14164 4547 14268
rect 4613 14164 4643 14268
rect 4709 14164 4739 14268
rect 4805 14164 4835 14268
rect 4901 14164 4931 14268
rect 363 12873 393 12977
rect 459 12873 489 12977
rect 555 12873 585 12977
rect 651 12873 681 12977
rect 747 12873 777 12977
rect 843 12873 873 12977
rect 939 12873 969 12977
rect 1035 12873 1065 12977
rect 1131 12873 1161 12977
rect 1227 12873 1257 12977
rect 2516 12877 2546 12981
rect 2612 12877 2642 12981
rect 2708 12877 2738 12981
rect 2804 12877 2834 12981
rect 2900 12877 2930 12981
rect 2996 12877 3026 12981
rect 3092 12877 3122 12981
rect 3188 12877 3218 12981
rect 3284 12877 3314 12981
rect 3380 12877 3410 12981
rect 3693 12885 3723 12985
rect 4037 12877 4067 12981
rect 4133 12877 4163 12981
rect 4229 12877 4259 12981
rect 4325 12877 4355 12981
rect 4421 12877 4451 12981
rect 4517 12877 4547 12981
rect 4613 12877 4643 12981
rect 4709 12877 4739 12981
rect 4805 12877 4835 12981
rect 4901 12877 4931 12981
rect 363 11586 393 11690
rect 459 11586 489 11690
rect 555 11586 585 11690
rect 651 11586 681 11690
rect 747 11586 777 11690
rect 843 11586 873 11690
rect 939 11586 969 11690
rect 1035 11586 1065 11690
rect 1131 11586 1161 11690
rect 1227 11586 1257 11690
rect 2516 11590 2546 11694
rect 2612 11590 2642 11694
rect 2708 11590 2738 11694
rect 2804 11590 2834 11694
rect 2900 11590 2930 11694
rect 2996 11590 3026 11694
rect 3092 11590 3122 11694
rect 3188 11590 3218 11694
rect 3284 11590 3314 11694
rect 3380 11590 3410 11694
rect 3693 11598 3723 11698
rect 4037 11590 4067 11694
rect 4133 11590 4163 11694
rect 4229 11590 4259 11694
rect 4325 11590 4355 11694
rect 4421 11590 4451 11694
rect 4517 11590 4547 11694
rect 4613 11590 4643 11694
rect 4709 11590 4739 11694
rect 4805 11590 4835 11694
rect 4901 11590 4931 11694
rect 363 10299 393 10403
rect 459 10299 489 10403
rect 555 10299 585 10403
rect 651 10299 681 10403
rect 747 10299 777 10403
rect 843 10299 873 10403
rect 939 10299 969 10403
rect 1035 10299 1065 10403
rect 1131 10299 1161 10403
rect 1227 10299 1257 10403
rect 2516 10303 2546 10407
rect 2612 10303 2642 10407
rect 2708 10303 2738 10407
rect 2804 10303 2834 10407
rect 2900 10303 2930 10407
rect 2996 10303 3026 10407
rect 3092 10303 3122 10407
rect 3188 10303 3218 10407
rect 3284 10303 3314 10407
rect 3380 10303 3410 10407
rect 3693 10311 3723 10411
rect 4037 10303 4067 10407
rect 4133 10303 4163 10407
rect 4229 10303 4259 10407
rect 4325 10303 4355 10407
rect 4421 10303 4451 10407
rect 4517 10303 4547 10407
rect 4613 10303 4643 10407
rect 4709 10303 4739 10407
rect 4805 10303 4835 10407
rect 4901 10303 4931 10407
rect 363 9012 393 9116
rect 459 9012 489 9116
rect 555 9012 585 9116
rect 651 9012 681 9116
rect 747 9012 777 9116
rect 843 9012 873 9116
rect 939 9012 969 9116
rect 1035 9012 1065 9116
rect 1131 9012 1161 9116
rect 1227 9012 1257 9116
rect 2516 9016 2546 9120
rect 2612 9016 2642 9120
rect 2708 9016 2738 9120
rect 2804 9016 2834 9120
rect 2900 9016 2930 9120
rect 2996 9016 3026 9120
rect 3092 9016 3122 9120
rect 3188 9016 3218 9120
rect 3284 9016 3314 9120
rect 3380 9016 3410 9120
rect 3693 9024 3723 9124
rect 4037 9016 4067 9120
rect 4133 9016 4163 9120
rect 4229 9016 4259 9120
rect 4325 9016 4355 9120
rect 4421 9016 4451 9120
rect 4517 9016 4547 9120
rect 4613 9016 4643 9120
rect 4709 9016 4739 9120
rect 4805 9016 4835 9120
rect 4901 9016 4931 9120
rect 363 7725 393 7829
rect 459 7725 489 7829
rect 555 7725 585 7829
rect 651 7725 681 7829
rect 747 7725 777 7829
rect 843 7725 873 7829
rect 939 7725 969 7829
rect 1035 7725 1065 7829
rect 1131 7725 1161 7829
rect 1227 7725 1257 7829
rect 2516 7729 2546 7833
rect 2612 7729 2642 7833
rect 2708 7729 2738 7833
rect 2804 7729 2834 7833
rect 2900 7729 2930 7833
rect 2996 7729 3026 7833
rect 3092 7729 3122 7833
rect 3188 7729 3218 7833
rect 3284 7729 3314 7833
rect 3380 7729 3410 7833
rect 3693 7737 3723 7837
rect 4037 7729 4067 7833
rect 4133 7729 4163 7833
rect 4229 7729 4259 7833
rect 4325 7729 4355 7833
rect 4421 7729 4451 7833
rect 4517 7729 4547 7833
rect 4613 7729 4643 7833
rect 4709 7729 4739 7833
rect 4805 7729 4835 7833
rect 4901 7729 4931 7833
rect 363 6438 393 6542
rect 459 6438 489 6542
rect 555 6438 585 6542
rect 651 6438 681 6542
rect 747 6438 777 6542
rect 843 6438 873 6542
rect 939 6438 969 6542
rect 1035 6438 1065 6542
rect 1131 6438 1161 6542
rect 1227 6438 1257 6542
rect 2516 6442 2546 6546
rect 2612 6442 2642 6546
rect 2708 6442 2738 6546
rect 2804 6442 2834 6546
rect 2900 6442 2930 6546
rect 2996 6442 3026 6546
rect 3092 6442 3122 6546
rect 3188 6442 3218 6546
rect 3284 6442 3314 6546
rect 3380 6442 3410 6546
rect 3693 6450 3723 6550
rect 4037 6442 4067 6546
rect 4133 6442 4163 6546
rect 4229 6442 4259 6546
rect 4325 6442 4355 6546
rect 4421 6442 4451 6546
rect 4517 6442 4547 6546
rect 4613 6442 4643 6546
rect 4709 6442 4739 6546
rect 4805 6442 4835 6546
rect 4901 6442 4931 6546
rect 363 5151 393 5255
rect 459 5151 489 5255
rect 555 5151 585 5255
rect 651 5151 681 5255
rect 747 5151 777 5255
rect 843 5151 873 5255
rect 939 5151 969 5255
rect 1035 5151 1065 5255
rect 1131 5151 1161 5255
rect 1227 5151 1257 5255
rect 2516 5155 2546 5259
rect 2612 5155 2642 5259
rect 2708 5155 2738 5259
rect 2804 5155 2834 5259
rect 2900 5155 2930 5259
rect 2996 5155 3026 5259
rect 3092 5155 3122 5259
rect 3188 5155 3218 5259
rect 3284 5155 3314 5259
rect 3380 5155 3410 5259
rect 3693 5163 3723 5263
rect 4037 5155 4067 5259
rect 4133 5155 4163 5259
rect 4229 5155 4259 5259
rect 4325 5155 4355 5259
rect 4421 5155 4451 5259
rect 4517 5155 4547 5259
rect 4613 5155 4643 5259
rect 4709 5155 4739 5259
rect 4805 5155 4835 5259
rect 4901 5155 4931 5259
rect 363 3864 393 3968
rect 459 3864 489 3968
rect 555 3864 585 3968
rect 651 3864 681 3968
rect 747 3864 777 3968
rect 843 3864 873 3968
rect 939 3864 969 3968
rect 1035 3864 1065 3968
rect 1131 3864 1161 3968
rect 1227 3864 1257 3968
rect 2516 3868 2546 3972
rect 2612 3868 2642 3972
rect 2708 3868 2738 3972
rect 2804 3868 2834 3972
rect 2900 3868 2930 3972
rect 2996 3868 3026 3972
rect 3092 3868 3122 3972
rect 3188 3868 3218 3972
rect 3284 3868 3314 3972
rect 3380 3868 3410 3972
rect 3693 3876 3723 3976
rect 4037 3868 4067 3972
rect 4133 3868 4163 3972
rect 4229 3868 4259 3972
rect 4325 3868 4355 3972
rect 4421 3868 4451 3972
rect 4517 3868 4547 3972
rect 4613 3868 4643 3972
rect 4709 3868 4739 3972
rect 4805 3868 4835 3972
rect 4901 3868 4931 3972
rect 363 2577 393 2681
rect 459 2577 489 2681
rect 555 2577 585 2681
rect 651 2577 681 2681
rect 747 2577 777 2681
rect 843 2577 873 2681
rect 939 2577 969 2681
rect 1035 2577 1065 2681
rect 1131 2577 1161 2681
rect 1227 2577 1257 2681
rect 2516 2581 2546 2685
rect 2612 2581 2642 2685
rect 2708 2581 2738 2685
rect 2804 2581 2834 2685
rect 2900 2581 2930 2685
rect 2996 2581 3026 2685
rect 3092 2581 3122 2685
rect 3188 2581 3218 2685
rect 3284 2581 3314 2685
rect 3380 2581 3410 2685
rect 3693 2589 3723 2689
rect 4037 2581 4067 2685
rect 4133 2581 4163 2685
rect 4229 2581 4259 2685
rect 4325 2581 4355 2685
rect 4421 2581 4451 2685
rect 4517 2581 4547 2685
rect 4613 2581 4643 2685
rect 4709 2581 4739 2685
rect 4805 2581 4835 2685
rect 4901 2581 4931 2685
rect 363 1290 393 1394
rect 459 1290 489 1394
rect 555 1290 585 1394
rect 651 1290 681 1394
rect 747 1290 777 1394
rect 843 1290 873 1394
rect 939 1290 969 1394
rect 1035 1290 1065 1394
rect 1131 1290 1161 1394
rect 1227 1290 1257 1394
rect 2516 1294 2546 1398
rect 2612 1294 2642 1398
rect 2708 1294 2738 1398
rect 2804 1294 2834 1398
rect 2900 1294 2930 1398
rect 2996 1294 3026 1398
rect 3092 1294 3122 1398
rect 3188 1294 3218 1398
rect 3284 1294 3314 1398
rect 3380 1294 3410 1398
rect 3693 1302 3723 1402
rect 4037 1294 4067 1398
rect 4133 1294 4163 1398
rect 4229 1294 4259 1398
rect 4325 1294 4355 1398
rect 4421 1294 4451 1398
rect 4517 1294 4547 1398
rect 4613 1294 4643 1398
rect 4709 1294 4739 1398
rect 4805 1294 4835 1398
rect 4901 1294 4931 1398
<< scnmos >>
rect 5400 41212 5430 41342
rect 5400 39925 5430 40055
rect 5400 38638 5430 38768
rect 5400 37351 5430 37481
rect 5400 36064 5430 36194
rect 5400 34777 5430 34907
rect 5400 33490 5430 33620
rect 5400 32203 5430 32333
rect 5400 30916 5430 31046
rect 5400 29629 5430 29759
rect 5400 28342 5430 28472
rect 5400 27055 5430 27185
rect 5400 25768 5430 25898
rect 5400 24481 5430 24611
rect 5400 23194 5430 23324
rect 5400 21907 5430 22037
rect 5400 20620 5430 20750
rect 5400 19333 5430 19463
rect 5400 18046 5430 18176
rect 5400 16759 5430 16889
rect 5400 15472 5430 15602
rect 5400 14185 5430 14315
rect 5400 12898 5430 13028
rect 5400 11611 5430 11741
rect 5400 10324 5430 10454
rect 5400 9037 5430 9167
rect 5400 7750 5430 7880
rect 5400 6463 5430 6593
rect 5400 5176 5430 5306
rect 5400 3889 5430 4019
rect 5400 2602 5430 2732
rect 5400 1315 5430 1445
<< pmos >>
rect 363 41599 393 41871
rect 459 41599 489 41871
rect 555 41599 585 41871
rect 651 41599 681 41871
rect 747 41599 777 41871
rect 843 41599 873 41871
rect 939 41599 969 41871
rect 1035 41599 1065 41871
rect 1131 41599 1161 41871
rect 1227 41599 1257 41871
rect 2516 41603 2546 41875
rect 2612 41603 2642 41875
rect 2708 41603 2738 41875
rect 2804 41603 2834 41875
rect 2900 41603 2930 41875
rect 2996 41603 3026 41875
rect 3092 41603 3122 41875
rect 3188 41603 3218 41875
rect 3284 41603 3314 41875
rect 3380 41603 3410 41875
rect 4037 41603 4067 41875
rect 4133 41603 4163 41875
rect 4229 41603 4259 41875
rect 4325 41603 4355 41875
rect 4421 41603 4451 41875
rect 4517 41603 4547 41875
rect 4613 41603 4643 41875
rect 4709 41603 4739 41875
rect 4805 41603 4835 41875
rect 4901 41603 4931 41875
rect 363 40312 393 40584
rect 459 40312 489 40584
rect 555 40312 585 40584
rect 651 40312 681 40584
rect 747 40312 777 40584
rect 843 40312 873 40584
rect 939 40312 969 40584
rect 1035 40312 1065 40584
rect 1131 40312 1161 40584
rect 1227 40312 1257 40584
rect 2516 40316 2546 40588
rect 2612 40316 2642 40588
rect 2708 40316 2738 40588
rect 2804 40316 2834 40588
rect 2900 40316 2930 40588
rect 2996 40316 3026 40588
rect 3092 40316 3122 40588
rect 3188 40316 3218 40588
rect 3284 40316 3314 40588
rect 3380 40316 3410 40588
rect 4037 40316 4067 40588
rect 4133 40316 4163 40588
rect 4229 40316 4259 40588
rect 4325 40316 4355 40588
rect 4421 40316 4451 40588
rect 4517 40316 4547 40588
rect 4613 40316 4643 40588
rect 4709 40316 4739 40588
rect 4805 40316 4835 40588
rect 4901 40316 4931 40588
rect 363 39025 393 39297
rect 459 39025 489 39297
rect 555 39025 585 39297
rect 651 39025 681 39297
rect 747 39025 777 39297
rect 843 39025 873 39297
rect 939 39025 969 39297
rect 1035 39025 1065 39297
rect 1131 39025 1161 39297
rect 1227 39025 1257 39297
rect 2516 39029 2546 39301
rect 2612 39029 2642 39301
rect 2708 39029 2738 39301
rect 2804 39029 2834 39301
rect 2900 39029 2930 39301
rect 2996 39029 3026 39301
rect 3092 39029 3122 39301
rect 3188 39029 3218 39301
rect 3284 39029 3314 39301
rect 3380 39029 3410 39301
rect 4037 39029 4067 39301
rect 4133 39029 4163 39301
rect 4229 39029 4259 39301
rect 4325 39029 4355 39301
rect 4421 39029 4451 39301
rect 4517 39029 4547 39301
rect 4613 39029 4643 39301
rect 4709 39029 4739 39301
rect 4805 39029 4835 39301
rect 4901 39029 4931 39301
rect 363 37738 393 38010
rect 459 37738 489 38010
rect 555 37738 585 38010
rect 651 37738 681 38010
rect 747 37738 777 38010
rect 843 37738 873 38010
rect 939 37738 969 38010
rect 1035 37738 1065 38010
rect 1131 37738 1161 38010
rect 1227 37738 1257 38010
rect 2516 37742 2546 38014
rect 2612 37742 2642 38014
rect 2708 37742 2738 38014
rect 2804 37742 2834 38014
rect 2900 37742 2930 38014
rect 2996 37742 3026 38014
rect 3092 37742 3122 38014
rect 3188 37742 3218 38014
rect 3284 37742 3314 38014
rect 3380 37742 3410 38014
rect 4037 37742 4067 38014
rect 4133 37742 4163 38014
rect 4229 37742 4259 38014
rect 4325 37742 4355 38014
rect 4421 37742 4451 38014
rect 4517 37742 4547 38014
rect 4613 37742 4643 38014
rect 4709 37742 4739 38014
rect 4805 37742 4835 38014
rect 4901 37742 4931 38014
rect 363 36451 393 36723
rect 459 36451 489 36723
rect 555 36451 585 36723
rect 651 36451 681 36723
rect 747 36451 777 36723
rect 843 36451 873 36723
rect 939 36451 969 36723
rect 1035 36451 1065 36723
rect 1131 36451 1161 36723
rect 1227 36451 1257 36723
rect 2516 36455 2546 36727
rect 2612 36455 2642 36727
rect 2708 36455 2738 36727
rect 2804 36455 2834 36727
rect 2900 36455 2930 36727
rect 2996 36455 3026 36727
rect 3092 36455 3122 36727
rect 3188 36455 3218 36727
rect 3284 36455 3314 36727
rect 3380 36455 3410 36727
rect 4037 36455 4067 36727
rect 4133 36455 4163 36727
rect 4229 36455 4259 36727
rect 4325 36455 4355 36727
rect 4421 36455 4451 36727
rect 4517 36455 4547 36727
rect 4613 36455 4643 36727
rect 4709 36455 4739 36727
rect 4805 36455 4835 36727
rect 4901 36455 4931 36727
rect 363 35164 393 35436
rect 459 35164 489 35436
rect 555 35164 585 35436
rect 651 35164 681 35436
rect 747 35164 777 35436
rect 843 35164 873 35436
rect 939 35164 969 35436
rect 1035 35164 1065 35436
rect 1131 35164 1161 35436
rect 1227 35164 1257 35436
rect 2516 35168 2546 35440
rect 2612 35168 2642 35440
rect 2708 35168 2738 35440
rect 2804 35168 2834 35440
rect 2900 35168 2930 35440
rect 2996 35168 3026 35440
rect 3092 35168 3122 35440
rect 3188 35168 3218 35440
rect 3284 35168 3314 35440
rect 3380 35168 3410 35440
rect 4037 35168 4067 35440
rect 4133 35168 4163 35440
rect 4229 35168 4259 35440
rect 4325 35168 4355 35440
rect 4421 35168 4451 35440
rect 4517 35168 4547 35440
rect 4613 35168 4643 35440
rect 4709 35168 4739 35440
rect 4805 35168 4835 35440
rect 4901 35168 4931 35440
rect 363 33877 393 34149
rect 459 33877 489 34149
rect 555 33877 585 34149
rect 651 33877 681 34149
rect 747 33877 777 34149
rect 843 33877 873 34149
rect 939 33877 969 34149
rect 1035 33877 1065 34149
rect 1131 33877 1161 34149
rect 1227 33877 1257 34149
rect 2516 33881 2546 34153
rect 2612 33881 2642 34153
rect 2708 33881 2738 34153
rect 2804 33881 2834 34153
rect 2900 33881 2930 34153
rect 2996 33881 3026 34153
rect 3092 33881 3122 34153
rect 3188 33881 3218 34153
rect 3284 33881 3314 34153
rect 3380 33881 3410 34153
rect 4037 33881 4067 34153
rect 4133 33881 4163 34153
rect 4229 33881 4259 34153
rect 4325 33881 4355 34153
rect 4421 33881 4451 34153
rect 4517 33881 4547 34153
rect 4613 33881 4643 34153
rect 4709 33881 4739 34153
rect 4805 33881 4835 34153
rect 4901 33881 4931 34153
rect 363 32590 393 32862
rect 459 32590 489 32862
rect 555 32590 585 32862
rect 651 32590 681 32862
rect 747 32590 777 32862
rect 843 32590 873 32862
rect 939 32590 969 32862
rect 1035 32590 1065 32862
rect 1131 32590 1161 32862
rect 1227 32590 1257 32862
rect 2516 32594 2546 32866
rect 2612 32594 2642 32866
rect 2708 32594 2738 32866
rect 2804 32594 2834 32866
rect 2900 32594 2930 32866
rect 2996 32594 3026 32866
rect 3092 32594 3122 32866
rect 3188 32594 3218 32866
rect 3284 32594 3314 32866
rect 3380 32594 3410 32866
rect 4037 32594 4067 32866
rect 4133 32594 4163 32866
rect 4229 32594 4259 32866
rect 4325 32594 4355 32866
rect 4421 32594 4451 32866
rect 4517 32594 4547 32866
rect 4613 32594 4643 32866
rect 4709 32594 4739 32866
rect 4805 32594 4835 32866
rect 4901 32594 4931 32866
rect 363 31303 393 31575
rect 459 31303 489 31575
rect 555 31303 585 31575
rect 651 31303 681 31575
rect 747 31303 777 31575
rect 843 31303 873 31575
rect 939 31303 969 31575
rect 1035 31303 1065 31575
rect 1131 31303 1161 31575
rect 1227 31303 1257 31575
rect 2516 31307 2546 31579
rect 2612 31307 2642 31579
rect 2708 31307 2738 31579
rect 2804 31307 2834 31579
rect 2900 31307 2930 31579
rect 2996 31307 3026 31579
rect 3092 31307 3122 31579
rect 3188 31307 3218 31579
rect 3284 31307 3314 31579
rect 3380 31307 3410 31579
rect 4037 31307 4067 31579
rect 4133 31307 4163 31579
rect 4229 31307 4259 31579
rect 4325 31307 4355 31579
rect 4421 31307 4451 31579
rect 4517 31307 4547 31579
rect 4613 31307 4643 31579
rect 4709 31307 4739 31579
rect 4805 31307 4835 31579
rect 4901 31307 4931 31579
rect 363 30016 393 30288
rect 459 30016 489 30288
rect 555 30016 585 30288
rect 651 30016 681 30288
rect 747 30016 777 30288
rect 843 30016 873 30288
rect 939 30016 969 30288
rect 1035 30016 1065 30288
rect 1131 30016 1161 30288
rect 1227 30016 1257 30288
rect 2516 30020 2546 30292
rect 2612 30020 2642 30292
rect 2708 30020 2738 30292
rect 2804 30020 2834 30292
rect 2900 30020 2930 30292
rect 2996 30020 3026 30292
rect 3092 30020 3122 30292
rect 3188 30020 3218 30292
rect 3284 30020 3314 30292
rect 3380 30020 3410 30292
rect 4037 30020 4067 30292
rect 4133 30020 4163 30292
rect 4229 30020 4259 30292
rect 4325 30020 4355 30292
rect 4421 30020 4451 30292
rect 4517 30020 4547 30292
rect 4613 30020 4643 30292
rect 4709 30020 4739 30292
rect 4805 30020 4835 30292
rect 4901 30020 4931 30292
rect 363 28729 393 29001
rect 459 28729 489 29001
rect 555 28729 585 29001
rect 651 28729 681 29001
rect 747 28729 777 29001
rect 843 28729 873 29001
rect 939 28729 969 29001
rect 1035 28729 1065 29001
rect 1131 28729 1161 29001
rect 1227 28729 1257 29001
rect 2516 28733 2546 29005
rect 2612 28733 2642 29005
rect 2708 28733 2738 29005
rect 2804 28733 2834 29005
rect 2900 28733 2930 29005
rect 2996 28733 3026 29005
rect 3092 28733 3122 29005
rect 3188 28733 3218 29005
rect 3284 28733 3314 29005
rect 3380 28733 3410 29005
rect 4037 28733 4067 29005
rect 4133 28733 4163 29005
rect 4229 28733 4259 29005
rect 4325 28733 4355 29005
rect 4421 28733 4451 29005
rect 4517 28733 4547 29005
rect 4613 28733 4643 29005
rect 4709 28733 4739 29005
rect 4805 28733 4835 29005
rect 4901 28733 4931 29005
rect 363 27442 393 27714
rect 459 27442 489 27714
rect 555 27442 585 27714
rect 651 27442 681 27714
rect 747 27442 777 27714
rect 843 27442 873 27714
rect 939 27442 969 27714
rect 1035 27442 1065 27714
rect 1131 27442 1161 27714
rect 1227 27442 1257 27714
rect 2516 27446 2546 27718
rect 2612 27446 2642 27718
rect 2708 27446 2738 27718
rect 2804 27446 2834 27718
rect 2900 27446 2930 27718
rect 2996 27446 3026 27718
rect 3092 27446 3122 27718
rect 3188 27446 3218 27718
rect 3284 27446 3314 27718
rect 3380 27446 3410 27718
rect 4037 27446 4067 27718
rect 4133 27446 4163 27718
rect 4229 27446 4259 27718
rect 4325 27446 4355 27718
rect 4421 27446 4451 27718
rect 4517 27446 4547 27718
rect 4613 27446 4643 27718
rect 4709 27446 4739 27718
rect 4805 27446 4835 27718
rect 4901 27446 4931 27718
rect 363 26155 393 26427
rect 459 26155 489 26427
rect 555 26155 585 26427
rect 651 26155 681 26427
rect 747 26155 777 26427
rect 843 26155 873 26427
rect 939 26155 969 26427
rect 1035 26155 1065 26427
rect 1131 26155 1161 26427
rect 1227 26155 1257 26427
rect 2516 26159 2546 26431
rect 2612 26159 2642 26431
rect 2708 26159 2738 26431
rect 2804 26159 2834 26431
rect 2900 26159 2930 26431
rect 2996 26159 3026 26431
rect 3092 26159 3122 26431
rect 3188 26159 3218 26431
rect 3284 26159 3314 26431
rect 3380 26159 3410 26431
rect 4037 26159 4067 26431
rect 4133 26159 4163 26431
rect 4229 26159 4259 26431
rect 4325 26159 4355 26431
rect 4421 26159 4451 26431
rect 4517 26159 4547 26431
rect 4613 26159 4643 26431
rect 4709 26159 4739 26431
rect 4805 26159 4835 26431
rect 4901 26159 4931 26431
rect 363 24868 393 25140
rect 459 24868 489 25140
rect 555 24868 585 25140
rect 651 24868 681 25140
rect 747 24868 777 25140
rect 843 24868 873 25140
rect 939 24868 969 25140
rect 1035 24868 1065 25140
rect 1131 24868 1161 25140
rect 1227 24868 1257 25140
rect 2516 24872 2546 25144
rect 2612 24872 2642 25144
rect 2708 24872 2738 25144
rect 2804 24872 2834 25144
rect 2900 24872 2930 25144
rect 2996 24872 3026 25144
rect 3092 24872 3122 25144
rect 3188 24872 3218 25144
rect 3284 24872 3314 25144
rect 3380 24872 3410 25144
rect 4037 24872 4067 25144
rect 4133 24872 4163 25144
rect 4229 24872 4259 25144
rect 4325 24872 4355 25144
rect 4421 24872 4451 25144
rect 4517 24872 4547 25144
rect 4613 24872 4643 25144
rect 4709 24872 4739 25144
rect 4805 24872 4835 25144
rect 4901 24872 4931 25144
rect 363 23581 393 23853
rect 459 23581 489 23853
rect 555 23581 585 23853
rect 651 23581 681 23853
rect 747 23581 777 23853
rect 843 23581 873 23853
rect 939 23581 969 23853
rect 1035 23581 1065 23853
rect 1131 23581 1161 23853
rect 1227 23581 1257 23853
rect 2516 23585 2546 23857
rect 2612 23585 2642 23857
rect 2708 23585 2738 23857
rect 2804 23585 2834 23857
rect 2900 23585 2930 23857
rect 2996 23585 3026 23857
rect 3092 23585 3122 23857
rect 3188 23585 3218 23857
rect 3284 23585 3314 23857
rect 3380 23585 3410 23857
rect 4037 23585 4067 23857
rect 4133 23585 4163 23857
rect 4229 23585 4259 23857
rect 4325 23585 4355 23857
rect 4421 23585 4451 23857
rect 4517 23585 4547 23857
rect 4613 23585 4643 23857
rect 4709 23585 4739 23857
rect 4805 23585 4835 23857
rect 4901 23585 4931 23857
rect 363 22294 393 22566
rect 459 22294 489 22566
rect 555 22294 585 22566
rect 651 22294 681 22566
rect 747 22294 777 22566
rect 843 22294 873 22566
rect 939 22294 969 22566
rect 1035 22294 1065 22566
rect 1131 22294 1161 22566
rect 1227 22294 1257 22566
rect 2516 22298 2546 22570
rect 2612 22298 2642 22570
rect 2708 22298 2738 22570
rect 2804 22298 2834 22570
rect 2900 22298 2930 22570
rect 2996 22298 3026 22570
rect 3092 22298 3122 22570
rect 3188 22298 3218 22570
rect 3284 22298 3314 22570
rect 3380 22298 3410 22570
rect 4037 22298 4067 22570
rect 4133 22298 4163 22570
rect 4229 22298 4259 22570
rect 4325 22298 4355 22570
rect 4421 22298 4451 22570
rect 4517 22298 4547 22570
rect 4613 22298 4643 22570
rect 4709 22298 4739 22570
rect 4805 22298 4835 22570
rect 4901 22298 4931 22570
rect 363 21007 393 21279
rect 459 21007 489 21279
rect 555 21007 585 21279
rect 651 21007 681 21279
rect 747 21007 777 21279
rect 843 21007 873 21279
rect 939 21007 969 21279
rect 1035 21007 1065 21279
rect 1131 21007 1161 21279
rect 1227 21007 1257 21279
rect 2516 21011 2546 21283
rect 2612 21011 2642 21283
rect 2708 21011 2738 21283
rect 2804 21011 2834 21283
rect 2900 21011 2930 21283
rect 2996 21011 3026 21283
rect 3092 21011 3122 21283
rect 3188 21011 3218 21283
rect 3284 21011 3314 21283
rect 3380 21011 3410 21283
rect 4037 21011 4067 21283
rect 4133 21011 4163 21283
rect 4229 21011 4259 21283
rect 4325 21011 4355 21283
rect 4421 21011 4451 21283
rect 4517 21011 4547 21283
rect 4613 21011 4643 21283
rect 4709 21011 4739 21283
rect 4805 21011 4835 21283
rect 4901 21011 4931 21283
rect 363 19720 393 19992
rect 459 19720 489 19992
rect 555 19720 585 19992
rect 651 19720 681 19992
rect 747 19720 777 19992
rect 843 19720 873 19992
rect 939 19720 969 19992
rect 1035 19720 1065 19992
rect 1131 19720 1161 19992
rect 1227 19720 1257 19992
rect 2516 19724 2546 19996
rect 2612 19724 2642 19996
rect 2708 19724 2738 19996
rect 2804 19724 2834 19996
rect 2900 19724 2930 19996
rect 2996 19724 3026 19996
rect 3092 19724 3122 19996
rect 3188 19724 3218 19996
rect 3284 19724 3314 19996
rect 3380 19724 3410 19996
rect 4037 19724 4067 19996
rect 4133 19724 4163 19996
rect 4229 19724 4259 19996
rect 4325 19724 4355 19996
rect 4421 19724 4451 19996
rect 4517 19724 4547 19996
rect 4613 19724 4643 19996
rect 4709 19724 4739 19996
rect 4805 19724 4835 19996
rect 4901 19724 4931 19996
rect 363 18433 393 18705
rect 459 18433 489 18705
rect 555 18433 585 18705
rect 651 18433 681 18705
rect 747 18433 777 18705
rect 843 18433 873 18705
rect 939 18433 969 18705
rect 1035 18433 1065 18705
rect 1131 18433 1161 18705
rect 1227 18433 1257 18705
rect 2516 18437 2546 18709
rect 2612 18437 2642 18709
rect 2708 18437 2738 18709
rect 2804 18437 2834 18709
rect 2900 18437 2930 18709
rect 2996 18437 3026 18709
rect 3092 18437 3122 18709
rect 3188 18437 3218 18709
rect 3284 18437 3314 18709
rect 3380 18437 3410 18709
rect 4037 18437 4067 18709
rect 4133 18437 4163 18709
rect 4229 18437 4259 18709
rect 4325 18437 4355 18709
rect 4421 18437 4451 18709
rect 4517 18437 4547 18709
rect 4613 18437 4643 18709
rect 4709 18437 4739 18709
rect 4805 18437 4835 18709
rect 4901 18437 4931 18709
rect 363 17146 393 17418
rect 459 17146 489 17418
rect 555 17146 585 17418
rect 651 17146 681 17418
rect 747 17146 777 17418
rect 843 17146 873 17418
rect 939 17146 969 17418
rect 1035 17146 1065 17418
rect 1131 17146 1161 17418
rect 1227 17146 1257 17418
rect 2516 17150 2546 17422
rect 2612 17150 2642 17422
rect 2708 17150 2738 17422
rect 2804 17150 2834 17422
rect 2900 17150 2930 17422
rect 2996 17150 3026 17422
rect 3092 17150 3122 17422
rect 3188 17150 3218 17422
rect 3284 17150 3314 17422
rect 3380 17150 3410 17422
rect 4037 17150 4067 17422
rect 4133 17150 4163 17422
rect 4229 17150 4259 17422
rect 4325 17150 4355 17422
rect 4421 17150 4451 17422
rect 4517 17150 4547 17422
rect 4613 17150 4643 17422
rect 4709 17150 4739 17422
rect 4805 17150 4835 17422
rect 4901 17150 4931 17422
rect 363 15859 393 16131
rect 459 15859 489 16131
rect 555 15859 585 16131
rect 651 15859 681 16131
rect 747 15859 777 16131
rect 843 15859 873 16131
rect 939 15859 969 16131
rect 1035 15859 1065 16131
rect 1131 15859 1161 16131
rect 1227 15859 1257 16131
rect 2516 15863 2546 16135
rect 2612 15863 2642 16135
rect 2708 15863 2738 16135
rect 2804 15863 2834 16135
rect 2900 15863 2930 16135
rect 2996 15863 3026 16135
rect 3092 15863 3122 16135
rect 3188 15863 3218 16135
rect 3284 15863 3314 16135
rect 3380 15863 3410 16135
rect 4037 15863 4067 16135
rect 4133 15863 4163 16135
rect 4229 15863 4259 16135
rect 4325 15863 4355 16135
rect 4421 15863 4451 16135
rect 4517 15863 4547 16135
rect 4613 15863 4643 16135
rect 4709 15863 4739 16135
rect 4805 15863 4835 16135
rect 4901 15863 4931 16135
rect 363 14572 393 14844
rect 459 14572 489 14844
rect 555 14572 585 14844
rect 651 14572 681 14844
rect 747 14572 777 14844
rect 843 14572 873 14844
rect 939 14572 969 14844
rect 1035 14572 1065 14844
rect 1131 14572 1161 14844
rect 1227 14572 1257 14844
rect 2516 14576 2546 14848
rect 2612 14576 2642 14848
rect 2708 14576 2738 14848
rect 2804 14576 2834 14848
rect 2900 14576 2930 14848
rect 2996 14576 3026 14848
rect 3092 14576 3122 14848
rect 3188 14576 3218 14848
rect 3284 14576 3314 14848
rect 3380 14576 3410 14848
rect 4037 14576 4067 14848
rect 4133 14576 4163 14848
rect 4229 14576 4259 14848
rect 4325 14576 4355 14848
rect 4421 14576 4451 14848
rect 4517 14576 4547 14848
rect 4613 14576 4643 14848
rect 4709 14576 4739 14848
rect 4805 14576 4835 14848
rect 4901 14576 4931 14848
rect 363 13285 393 13557
rect 459 13285 489 13557
rect 555 13285 585 13557
rect 651 13285 681 13557
rect 747 13285 777 13557
rect 843 13285 873 13557
rect 939 13285 969 13557
rect 1035 13285 1065 13557
rect 1131 13285 1161 13557
rect 1227 13285 1257 13557
rect 2516 13289 2546 13561
rect 2612 13289 2642 13561
rect 2708 13289 2738 13561
rect 2804 13289 2834 13561
rect 2900 13289 2930 13561
rect 2996 13289 3026 13561
rect 3092 13289 3122 13561
rect 3188 13289 3218 13561
rect 3284 13289 3314 13561
rect 3380 13289 3410 13561
rect 4037 13289 4067 13561
rect 4133 13289 4163 13561
rect 4229 13289 4259 13561
rect 4325 13289 4355 13561
rect 4421 13289 4451 13561
rect 4517 13289 4547 13561
rect 4613 13289 4643 13561
rect 4709 13289 4739 13561
rect 4805 13289 4835 13561
rect 4901 13289 4931 13561
rect 363 11998 393 12270
rect 459 11998 489 12270
rect 555 11998 585 12270
rect 651 11998 681 12270
rect 747 11998 777 12270
rect 843 11998 873 12270
rect 939 11998 969 12270
rect 1035 11998 1065 12270
rect 1131 11998 1161 12270
rect 1227 11998 1257 12270
rect 2516 12002 2546 12274
rect 2612 12002 2642 12274
rect 2708 12002 2738 12274
rect 2804 12002 2834 12274
rect 2900 12002 2930 12274
rect 2996 12002 3026 12274
rect 3092 12002 3122 12274
rect 3188 12002 3218 12274
rect 3284 12002 3314 12274
rect 3380 12002 3410 12274
rect 4037 12002 4067 12274
rect 4133 12002 4163 12274
rect 4229 12002 4259 12274
rect 4325 12002 4355 12274
rect 4421 12002 4451 12274
rect 4517 12002 4547 12274
rect 4613 12002 4643 12274
rect 4709 12002 4739 12274
rect 4805 12002 4835 12274
rect 4901 12002 4931 12274
rect 363 10711 393 10983
rect 459 10711 489 10983
rect 555 10711 585 10983
rect 651 10711 681 10983
rect 747 10711 777 10983
rect 843 10711 873 10983
rect 939 10711 969 10983
rect 1035 10711 1065 10983
rect 1131 10711 1161 10983
rect 1227 10711 1257 10983
rect 2516 10715 2546 10987
rect 2612 10715 2642 10987
rect 2708 10715 2738 10987
rect 2804 10715 2834 10987
rect 2900 10715 2930 10987
rect 2996 10715 3026 10987
rect 3092 10715 3122 10987
rect 3188 10715 3218 10987
rect 3284 10715 3314 10987
rect 3380 10715 3410 10987
rect 4037 10715 4067 10987
rect 4133 10715 4163 10987
rect 4229 10715 4259 10987
rect 4325 10715 4355 10987
rect 4421 10715 4451 10987
rect 4517 10715 4547 10987
rect 4613 10715 4643 10987
rect 4709 10715 4739 10987
rect 4805 10715 4835 10987
rect 4901 10715 4931 10987
rect 363 9424 393 9696
rect 459 9424 489 9696
rect 555 9424 585 9696
rect 651 9424 681 9696
rect 747 9424 777 9696
rect 843 9424 873 9696
rect 939 9424 969 9696
rect 1035 9424 1065 9696
rect 1131 9424 1161 9696
rect 1227 9424 1257 9696
rect 2516 9428 2546 9700
rect 2612 9428 2642 9700
rect 2708 9428 2738 9700
rect 2804 9428 2834 9700
rect 2900 9428 2930 9700
rect 2996 9428 3026 9700
rect 3092 9428 3122 9700
rect 3188 9428 3218 9700
rect 3284 9428 3314 9700
rect 3380 9428 3410 9700
rect 4037 9428 4067 9700
rect 4133 9428 4163 9700
rect 4229 9428 4259 9700
rect 4325 9428 4355 9700
rect 4421 9428 4451 9700
rect 4517 9428 4547 9700
rect 4613 9428 4643 9700
rect 4709 9428 4739 9700
rect 4805 9428 4835 9700
rect 4901 9428 4931 9700
rect 363 8137 393 8409
rect 459 8137 489 8409
rect 555 8137 585 8409
rect 651 8137 681 8409
rect 747 8137 777 8409
rect 843 8137 873 8409
rect 939 8137 969 8409
rect 1035 8137 1065 8409
rect 1131 8137 1161 8409
rect 1227 8137 1257 8409
rect 2516 8141 2546 8413
rect 2612 8141 2642 8413
rect 2708 8141 2738 8413
rect 2804 8141 2834 8413
rect 2900 8141 2930 8413
rect 2996 8141 3026 8413
rect 3092 8141 3122 8413
rect 3188 8141 3218 8413
rect 3284 8141 3314 8413
rect 3380 8141 3410 8413
rect 4037 8141 4067 8413
rect 4133 8141 4163 8413
rect 4229 8141 4259 8413
rect 4325 8141 4355 8413
rect 4421 8141 4451 8413
rect 4517 8141 4547 8413
rect 4613 8141 4643 8413
rect 4709 8141 4739 8413
rect 4805 8141 4835 8413
rect 4901 8141 4931 8413
rect 363 6850 393 7122
rect 459 6850 489 7122
rect 555 6850 585 7122
rect 651 6850 681 7122
rect 747 6850 777 7122
rect 843 6850 873 7122
rect 939 6850 969 7122
rect 1035 6850 1065 7122
rect 1131 6850 1161 7122
rect 1227 6850 1257 7122
rect 2516 6854 2546 7126
rect 2612 6854 2642 7126
rect 2708 6854 2738 7126
rect 2804 6854 2834 7126
rect 2900 6854 2930 7126
rect 2996 6854 3026 7126
rect 3092 6854 3122 7126
rect 3188 6854 3218 7126
rect 3284 6854 3314 7126
rect 3380 6854 3410 7126
rect 4037 6854 4067 7126
rect 4133 6854 4163 7126
rect 4229 6854 4259 7126
rect 4325 6854 4355 7126
rect 4421 6854 4451 7126
rect 4517 6854 4547 7126
rect 4613 6854 4643 7126
rect 4709 6854 4739 7126
rect 4805 6854 4835 7126
rect 4901 6854 4931 7126
rect 363 5563 393 5835
rect 459 5563 489 5835
rect 555 5563 585 5835
rect 651 5563 681 5835
rect 747 5563 777 5835
rect 843 5563 873 5835
rect 939 5563 969 5835
rect 1035 5563 1065 5835
rect 1131 5563 1161 5835
rect 1227 5563 1257 5835
rect 2516 5567 2546 5839
rect 2612 5567 2642 5839
rect 2708 5567 2738 5839
rect 2804 5567 2834 5839
rect 2900 5567 2930 5839
rect 2996 5567 3026 5839
rect 3092 5567 3122 5839
rect 3188 5567 3218 5839
rect 3284 5567 3314 5839
rect 3380 5567 3410 5839
rect 4037 5567 4067 5839
rect 4133 5567 4163 5839
rect 4229 5567 4259 5839
rect 4325 5567 4355 5839
rect 4421 5567 4451 5839
rect 4517 5567 4547 5839
rect 4613 5567 4643 5839
rect 4709 5567 4739 5839
rect 4805 5567 4835 5839
rect 4901 5567 4931 5839
rect 363 4276 393 4548
rect 459 4276 489 4548
rect 555 4276 585 4548
rect 651 4276 681 4548
rect 747 4276 777 4548
rect 843 4276 873 4548
rect 939 4276 969 4548
rect 1035 4276 1065 4548
rect 1131 4276 1161 4548
rect 1227 4276 1257 4548
rect 2516 4280 2546 4552
rect 2612 4280 2642 4552
rect 2708 4280 2738 4552
rect 2804 4280 2834 4552
rect 2900 4280 2930 4552
rect 2996 4280 3026 4552
rect 3092 4280 3122 4552
rect 3188 4280 3218 4552
rect 3284 4280 3314 4552
rect 3380 4280 3410 4552
rect 4037 4280 4067 4552
rect 4133 4280 4163 4552
rect 4229 4280 4259 4552
rect 4325 4280 4355 4552
rect 4421 4280 4451 4552
rect 4517 4280 4547 4552
rect 4613 4280 4643 4552
rect 4709 4280 4739 4552
rect 4805 4280 4835 4552
rect 4901 4280 4931 4552
rect 363 2989 393 3261
rect 459 2989 489 3261
rect 555 2989 585 3261
rect 651 2989 681 3261
rect 747 2989 777 3261
rect 843 2989 873 3261
rect 939 2989 969 3261
rect 1035 2989 1065 3261
rect 1131 2989 1161 3261
rect 1227 2989 1257 3261
rect 2516 2993 2546 3265
rect 2612 2993 2642 3265
rect 2708 2993 2738 3265
rect 2804 2993 2834 3265
rect 2900 2993 2930 3265
rect 2996 2993 3026 3265
rect 3092 2993 3122 3265
rect 3188 2993 3218 3265
rect 3284 2993 3314 3265
rect 3380 2993 3410 3265
rect 4037 2993 4067 3265
rect 4133 2993 4163 3265
rect 4229 2993 4259 3265
rect 4325 2993 4355 3265
rect 4421 2993 4451 3265
rect 4517 2993 4547 3265
rect 4613 2993 4643 3265
rect 4709 2993 4739 3265
rect 4805 2993 4835 3265
rect 4901 2993 4931 3265
rect 363 1702 393 1974
rect 459 1702 489 1974
rect 555 1702 585 1974
rect 651 1702 681 1974
rect 747 1702 777 1974
rect 843 1702 873 1974
rect 939 1702 969 1974
rect 1035 1702 1065 1974
rect 1131 1702 1161 1974
rect 1227 1702 1257 1974
rect 2516 1706 2546 1978
rect 2612 1706 2642 1978
rect 2708 1706 2738 1978
rect 2804 1706 2834 1978
rect 2900 1706 2930 1978
rect 2996 1706 3026 1978
rect 3092 1706 3122 1978
rect 3188 1706 3218 1978
rect 3284 1706 3314 1978
rect 3380 1706 3410 1978
rect 4037 1706 4067 1978
rect 4133 1706 4163 1978
rect 4229 1706 4259 1978
rect 4325 1706 4355 1978
rect 4421 1706 4451 1978
rect 4517 1706 4547 1978
rect 4613 1706 4643 1978
rect 4709 1706 4739 1978
rect 4805 1706 4835 1978
rect 4901 1706 4931 1978
<< scpmoshvt >>
rect 5400 41462 5430 41662
rect 5400 40175 5430 40375
rect 5400 38888 5430 39088
rect 5400 37601 5430 37801
rect 5400 36314 5430 36514
rect 5400 35027 5430 35227
rect 5400 33740 5430 33940
rect 5400 32453 5430 32653
rect 5400 31166 5430 31366
rect 5400 29879 5430 30079
rect 5400 28592 5430 28792
rect 5400 27305 5430 27505
rect 5400 26018 5430 26218
rect 5400 24731 5430 24931
rect 5400 23444 5430 23644
rect 5400 22157 5430 22357
rect 5400 20870 5430 21070
rect 5400 19583 5430 19783
rect 5400 18296 5430 18496
rect 5400 17009 5430 17209
rect 5400 15722 5430 15922
rect 5400 14435 5430 14635
rect 5400 13148 5430 13348
rect 5400 11861 5430 12061
rect 5400 10574 5430 10774
rect 5400 9287 5430 9487
rect 5400 8000 5430 8200
rect 5400 6713 5430 6913
rect 5400 5426 5430 5626
rect 5400 4139 5430 4339
rect 5400 2852 5430 3052
rect 5400 1565 5430 1765
<< ndiff >>
rect 301 41256 363 41291
rect 301 41222 313 41256
rect 347 41222 363 41256
rect 301 41187 363 41222
rect 393 41256 459 41291
rect 393 41222 409 41256
rect 443 41222 459 41256
rect 393 41187 459 41222
rect 489 41256 555 41291
rect 489 41222 505 41256
rect 539 41222 555 41256
rect 489 41187 555 41222
rect 585 41256 651 41291
rect 585 41222 601 41256
rect 635 41222 651 41256
rect 585 41187 651 41222
rect 681 41256 747 41291
rect 681 41222 697 41256
rect 731 41222 747 41256
rect 681 41187 747 41222
rect 777 41256 843 41291
rect 777 41222 793 41256
rect 827 41222 843 41256
rect 777 41187 843 41222
rect 873 41256 939 41291
rect 873 41222 889 41256
rect 923 41222 939 41256
rect 873 41187 939 41222
rect 969 41256 1035 41291
rect 969 41222 985 41256
rect 1019 41222 1035 41256
rect 969 41187 1035 41222
rect 1065 41256 1131 41291
rect 1065 41222 1081 41256
rect 1115 41222 1131 41256
rect 1065 41187 1131 41222
rect 1161 41256 1227 41291
rect 1161 41222 1177 41256
rect 1211 41222 1227 41256
rect 1161 41187 1227 41222
rect 1257 41256 1319 41291
rect 1257 41222 1273 41256
rect 1307 41222 1319 41256
rect 1257 41187 1319 41222
rect 2454 41260 2516 41295
rect 2454 41226 2466 41260
rect 2500 41226 2516 41260
rect 2454 41191 2516 41226
rect 2546 41260 2612 41295
rect 2546 41226 2562 41260
rect 2596 41226 2612 41260
rect 2546 41191 2612 41226
rect 2642 41260 2708 41295
rect 2642 41226 2658 41260
rect 2692 41226 2708 41260
rect 2642 41191 2708 41226
rect 2738 41260 2804 41295
rect 2738 41226 2754 41260
rect 2788 41226 2804 41260
rect 2738 41191 2804 41226
rect 2834 41260 2900 41295
rect 2834 41226 2850 41260
rect 2884 41226 2900 41260
rect 2834 41191 2900 41226
rect 2930 41260 2996 41295
rect 2930 41226 2946 41260
rect 2980 41226 2996 41260
rect 2930 41191 2996 41226
rect 3026 41260 3092 41295
rect 3026 41226 3042 41260
rect 3076 41226 3092 41260
rect 3026 41191 3092 41226
rect 3122 41260 3188 41295
rect 3122 41226 3138 41260
rect 3172 41226 3188 41260
rect 3122 41191 3188 41226
rect 3218 41260 3284 41295
rect 3218 41226 3234 41260
rect 3268 41226 3284 41260
rect 3218 41191 3284 41226
rect 3314 41260 3380 41295
rect 3314 41226 3330 41260
rect 3364 41226 3380 41260
rect 3314 41191 3380 41226
rect 3410 41260 3472 41295
rect 3410 41226 3426 41260
rect 3460 41226 3472 41260
rect 3410 41191 3472 41226
rect 3635 41287 3693 41299
rect 3635 41211 3647 41287
rect 3681 41211 3693 41287
rect 3635 41199 3693 41211
rect 3723 41287 3781 41299
rect 3723 41211 3735 41287
rect 3769 41211 3781 41287
rect 3723 41199 3781 41211
rect 3975 41260 4037 41295
rect 3975 41226 3987 41260
rect 4021 41226 4037 41260
rect 3975 41191 4037 41226
rect 4067 41260 4133 41295
rect 4067 41226 4083 41260
rect 4117 41226 4133 41260
rect 4067 41191 4133 41226
rect 4163 41260 4229 41295
rect 4163 41226 4179 41260
rect 4213 41226 4229 41260
rect 4163 41191 4229 41226
rect 4259 41260 4325 41295
rect 4259 41226 4275 41260
rect 4309 41226 4325 41260
rect 4259 41191 4325 41226
rect 4355 41260 4421 41295
rect 4355 41226 4371 41260
rect 4405 41226 4421 41260
rect 4355 41191 4421 41226
rect 4451 41260 4517 41295
rect 4451 41226 4467 41260
rect 4501 41226 4517 41260
rect 4451 41191 4517 41226
rect 4547 41260 4613 41295
rect 4547 41226 4563 41260
rect 4597 41226 4613 41260
rect 4547 41191 4613 41226
rect 4643 41260 4709 41295
rect 4643 41226 4659 41260
rect 4693 41226 4709 41260
rect 4643 41191 4709 41226
rect 4739 41260 4805 41295
rect 4739 41226 4755 41260
rect 4789 41226 4805 41260
rect 4739 41191 4805 41226
rect 4835 41260 4901 41295
rect 4835 41226 4851 41260
rect 4885 41226 4901 41260
rect 4835 41191 4901 41226
rect 4931 41260 4993 41295
rect 4931 41226 4947 41260
rect 4981 41226 4993 41260
rect 4931 41191 4993 41226
rect 5348 41330 5400 41342
rect 5348 41296 5356 41330
rect 5390 41296 5400 41330
rect 5348 41262 5400 41296
rect 5348 41228 5356 41262
rect 5390 41228 5400 41262
rect 5348 41212 5400 41228
rect 5430 41330 5482 41342
rect 5430 41296 5440 41330
rect 5474 41296 5482 41330
rect 5430 41262 5482 41296
rect 5430 41228 5440 41262
rect 5474 41228 5482 41262
rect 5430 41212 5482 41228
rect 301 39969 363 40004
rect 301 39935 313 39969
rect 347 39935 363 39969
rect 301 39900 363 39935
rect 393 39969 459 40004
rect 393 39935 409 39969
rect 443 39935 459 39969
rect 393 39900 459 39935
rect 489 39969 555 40004
rect 489 39935 505 39969
rect 539 39935 555 39969
rect 489 39900 555 39935
rect 585 39969 651 40004
rect 585 39935 601 39969
rect 635 39935 651 39969
rect 585 39900 651 39935
rect 681 39969 747 40004
rect 681 39935 697 39969
rect 731 39935 747 39969
rect 681 39900 747 39935
rect 777 39969 843 40004
rect 777 39935 793 39969
rect 827 39935 843 39969
rect 777 39900 843 39935
rect 873 39969 939 40004
rect 873 39935 889 39969
rect 923 39935 939 39969
rect 873 39900 939 39935
rect 969 39969 1035 40004
rect 969 39935 985 39969
rect 1019 39935 1035 39969
rect 969 39900 1035 39935
rect 1065 39969 1131 40004
rect 1065 39935 1081 39969
rect 1115 39935 1131 39969
rect 1065 39900 1131 39935
rect 1161 39969 1227 40004
rect 1161 39935 1177 39969
rect 1211 39935 1227 39969
rect 1161 39900 1227 39935
rect 1257 39969 1319 40004
rect 1257 39935 1273 39969
rect 1307 39935 1319 39969
rect 1257 39900 1319 39935
rect 2454 39973 2516 40008
rect 2454 39939 2466 39973
rect 2500 39939 2516 39973
rect 2454 39904 2516 39939
rect 2546 39973 2612 40008
rect 2546 39939 2562 39973
rect 2596 39939 2612 39973
rect 2546 39904 2612 39939
rect 2642 39973 2708 40008
rect 2642 39939 2658 39973
rect 2692 39939 2708 39973
rect 2642 39904 2708 39939
rect 2738 39973 2804 40008
rect 2738 39939 2754 39973
rect 2788 39939 2804 39973
rect 2738 39904 2804 39939
rect 2834 39973 2900 40008
rect 2834 39939 2850 39973
rect 2884 39939 2900 39973
rect 2834 39904 2900 39939
rect 2930 39973 2996 40008
rect 2930 39939 2946 39973
rect 2980 39939 2996 39973
rect 2930 39904 2996 39939
rect 3026 39973 3092 40008
rect 3026 39939 3042 39973
rect 3076 39939 3092 39973
rect 3026 39904 3092 39939
rect 3122 39973 3188 40008
rect 3122 39939 3138 39973
rect 3172 39939 3188 39973
rect 3122 39904 3188 39939
rect 3218 39973 3284 40008
rect 3218 39939 3234 39973
rect 3268 39939 3284 39973
rect 3218 39904 3284 39939
rect 3314 39973 3380 40008
rect 3314 39939 3330 39973
rect 3364 39939 3380 39973
rect 3314 39904 3380 39939
rect 3410 39973 3472 40008
rect 3410 39939 3426 39973
rect 3460 39939 3472 39973
rect 3410 39904 3472 39939
rect 3635 40000 3693 40012
rect 3635 39924 3647 40000
rect 3681 39924 3693 40000
rect 3635 39912 3693 39924
rect 3723 40000 3781 40012
rect 3723 39924 3735 40000
rect 3769 39924 3781 40000
rect 3723 39912 3781 39924
rect 3975 39973 4037 40008
rect 3975 39939 3987 39973
rect 4021 39939 4037 39973
rect 3975 39904 4037 39939
rect 4067 39973 4133 40008
rect 4067 39939 4083 39973
rect 4117 39939 4133 39973
rect 4067 39904 4133 39939
rect 4163 39973 4229 40008
rect 4163 39939 4179 39973
rect 4213 39939 4229 39973
rect 4163 39904 4229 39939
rect 4259 39973 4325 40008
rect 4259 39939 4275 39973
rect 4309 39939 4325 39973
rect 4259 39904 4325 39939
rect 4355 39973 4421 40008
rect 4355 39939 4371 39973
rect 4405 39939 4421 39973
rect 4355 39904 4421 39939
rect 4451 39973 4517 40008
rect 4451 39939 4467 39973
rect 4501 39939 4517 39973
rect 4451 39904 4517 39939
rect 4547 39973 4613 40008
rect 4547 39939 4563 39973
rect 4597 39939 4613 39973
rect 4547 39904 4613 39939
rect 4643 39973 4709 40008
rect 4643 39939 4659 39973
rect 4693 39939 4709 39973
rect 4643 39904 4709 39939
rect 4739 39973 4805 40008
rect 4739 39939 4755 39973
rect 4789 39939 4805 39973
rect 4739 39904 4805 39939
rect 4835 39973 4901 40008
rect 4835 39939 4851 39973
rect 4885 39939 4901 39973
rect 4835 39904 4901 39939
rect 4931 39973 4993 40008
rect 4931 39939 4947 39973
rect 4981 39939 4993 39973
rect 4931 39904 4993 39939
rect 5348 40043 5400 40055
rect 5348 40009 5356 40043
rect 5390 40009 5400 40043
rect 5348 39975 5400 40009
rect 5348 39941 5356 39975
rect 5390 39941 5400 39975
rect 5348 39925 5400 39941
rect 5430 40043 5482 40055
rect 5430 40009 5440 40043
rect 5474 40009 5482 40043
rect 5430 39975 5482 40009
rect 5430 39941 5440 39975
rect 5474 39941 5482 39975
rect 5430 39925 5482 39941
rect 301 38682 363 38717
rect 301 38648 313 38682
rect 347 38648 363 38682
rect 301 38613 363 38648
rect 393 38682 459 38717
rect 393 38648 409 38682
rect 443 38648 459 38682
rect 393 38613 459 38648
rect 489 38682 555 38717
rect 489 38648 505 38682
rect 539 38648 555 38682
rect 489 38613 555 38648
rect 585 38682 651 38717
rect 585 38648 601 38682
rect 635 38648 651 38682
rect 585 38613 651 38648
rect 681 38682 747 38717
rect 681 38648 697 38682
rect 731 38648 747 38682
rect 681 38613 747 38648
rect 777 38682 843 38717
rect 777 38648 793 38682
rect 827 38648 843 38682
rect 777 38613 843 38648
rect 873 38682 939 38717
rect 873 38648 889 38682
rect 923 38648 939 38682
rect 873 38613 939 38648
rect 969 38682 1035 38717
rect 969 38648 985 38682
rect 1019 38648 1035 38682
rect 969 38613 1035 38648
rect 1065 38682 1131 38717
rect 1065 38648 1081 38682
rect 1115 38648 1131 38682
rect 1065 38613 1131 38648
rect 1161 38682 1227 38717
rect 1161 38648 1177 38682
rect 1211 38648 1227 38682
rect 1161 38613 1227 38648
rect 1257 38682 1319 38717
rect 1257 38648 1273 38682
rect 1307 38648 1319 38682
rect 1257 38613 1319 38648
rect 2454 38686 2516 38721
rect 2454 38652 2466 38686
rect 2500 38652 2516 38686
rect 2454 38617 2516 38652
rect 2546 38686 2612 38721
rect 2546 38652 2562 38686
rect 2596 38652 2612 38686
rect 2546 38617 2612 38652
rect 2642 38686 2708 38721
rect 2642 38652 2658 38686
rect 2692 38652 2708 38686
rect 2642 38617 2708 38652
rect 2738 38686 2804 38721
rect 2738 38652 2754 38686
rect 2788 38652 2804 38686
rect 2738 38617 2804 38652
rect 2834 38686 2900 38721
rect 2834 38652 2850 38686
rect 2884 38652 2900 38686
rect 2834 38617 2900 38652
rect 2930 38686 2996 38721
rect 2930 38652 2946 38686
rect 2980 38652 2996 38686
rect 2930 38617 2996 38652
rect 3026 38686 3092 38721
rect 3026 38652 3042 38686
rect 3076 38652 3092 38686
rect 3026 38617 3092 38652
rect 3122 38686 3188 38721
rect 3122 38652 3138 38686
rect 3172 38652 3188 38686
rect 3122 38617 3188 38652
rect 3218 38686 3284 38721
rect 3218 38652 3234 38686
rect 3268 38652 3284 38686
rect 3218 38617 3284 38652
rect 3314 38686 3380 38721
rect 3314 38652 3330 38686
rect 3364 38652 3380 38686
rect 3314 38617 3380 38652
rect 3410 38686 3472 38721
rect 3410 38652 3426 38686
rect 3460 38652 3472 38686
rect 3410 38617 3472 38652
rect 3635 38713 3693 38725
rect 3635 38637 3647 38713
rect 3681 38637 3693 38713
rect 3635 38625 3693 38637
rect 3723 38713 3781 38725
rect 3723 38637 3735 38713
rect 3769 38637 3781 38713
rect 3723 38625 3781 38637
rect 3975 38686 4037 38721
rect 3975 38652 3987 38686
rect 4021 38652 4037 38686
rect 3975 38617 4037 38652
rect 4067 38686 4133 38721
rect 4067 38652 4083 38686
rect 4117 38652 4133 38686
rect 4067 38617 4133 38652
rect 4163 38686 4229 38721
rect 4163 38652 4179 38686
rect 4213 38652 4229 38686
rect 4163 38617 4229 38652
rect 4259 38686 4325 38721
rect 4259 38652 4275 38686
rect 4309 38652 4325 38686
rect 4259 38617 4325 38652
rect 4355 38686 4421 38721
rect 4355 38652 4371 38686
rect 4405 38652 4421 38686
rect 4355 38617 4421 38652
rect 4451 38686 4517 38721
rect 4451 38652 4467 38686
rect 4501 38652 4517 38686
rect 4451 38617 4517 38652
rect 4547 38686 4613 38721
rect 4547 38652 4563 38686
rect 4597 38652 4613 38686
rect 4547 38617 4613 38652
rect 4643 38686 4709 38721
rect 4643 38652 4659 38686
rect 4693 38652 4709 38686
rect 4643 38617 4709 38652
rect 4739 38686 4805 38721
rect 4739 38652 4755 38686
rect 4789 38652 4805 38686
rect 4739 38617 4805 38652
rect 4835 38686 4901 38721
rect 4835 38652 4851 38686
rect 4885 38652 4901 38686
rect 4835 38617 4901 38652
rect 4931 38686 4993 38721
rect 4931 38652 4947 38686
rect 4981 38652 4993 38686
rect 4931 38617 4993 38652
rect 5348 38756 5400 38768
rect 5348 38722 5356 38756
rect 5390 38722 5400 38756
rect 5348 38688 5400 38722
rect 5348 38654 5356 38688
rect 5390 38654 5400 38688
rect 5348 38638 5400 38654
rect 5430 38756 5482 38768
rect 5430 38722 5440 38756
rect 5474 38722 5482 38756
rect 5430 38688 5482 38722
rect 5430 38654 5440 38688
rect 5474 38654 5482 38688
rect 5430 38638 5482 38654
rect 301 37395 363 37430
rect 301 37361 313 37395
rect 347 37361 363 37395
rect 301 37326 363 37361
rect 393 37395 459 37430
rect 393 37361 409 37395
rect 443 37361 459 37395
rect 393 37326 459 37361
rect 489 37395 555 37430
rect 489 37361 505 37395
rect 539 37361 555 37395
rect 489 37326 555 37361
rect 585 37395 651 37430
rect 585 37361 601 37395
rect 635 37361 651 37395
rect 585 37326 651 37361
rect 681 37395 747 37430
rect 681 37361 697 37395
rect 731 37361 747 37395
rect 681 37326 747 37361
rect 777 37395 843 37430
rect 777 37361 793 37395
rect 827 37361 843 37395
rect 777 37326 843 37361
rect 873 37395 939 37430
rect 873 37361 889 37395
rect 923 37361 939 37395
rect 873 37326 939 37361
rect 969 37395 1035 37430
rect 969 37361 985 37395
rect 1019 37361 1035 37395
rect 969 37326 1035 37361
rect 1065 37395 1131 37430
rect 1065 37361 1081 37395
rect 1115 37361 1131 37395
rect 1065 37326 1131 37361
rect 1161 37395 1227 37430
rect 1161 37361 1177 37395
rect 1211 37361 1227 37395
rect 1161 37326 1227 37361
rect 1257 37395 1319 37430
rect 1257 37361 1273 37395
rect 1307 37361 1319 37395
rect 1257 37326 1319 37361
rect 2454 37399 2516 37434
rect 2454 37365 2466 37399
rect 2500 37365 2516 37399
rect 2454 37330 2516 37365
rect 2546 37399 2612 37434
rect 2546 37365 2562 37399
rect 2596 37365 2612 37399
rect 2546 37330 2612 37365
rect 2642 37399 2708 37434
rect 2642 37365 2658 37399
rect 2692 37365 2708 37399
rect 2642 37330 2708 37365
rect 2738 37399 2804 37434
rect 2738 37365 2754 37399
rect 2788 37365 2804 37399
rect 2738 37330 2804 37365
rect 2834 37399 2900 37434
rect 2834 37365 2850 37399
rect 2884 37365 2900 37399
rect 2834 37330 2900 37365
rect 2930 37399 2996 37434
rect 2930 37365 2946 37399
rect 2980 37365 2996 37399
rect 2930 37330 2996 37365
rect 3026 37399 3092 37434
rect 3026 37365 3042 37399
rect 3076 37365 3092 37399
rect 3026 37330 3092 37365
rect 3122 37399 3188 37434
rect 3122 37365 3138 37399
rect 3172 37365 3188 37399
rect 3122 37330 3188 37365
rect 3218 37399 3284 37434
rect 3218 37365 3234 37399
rect 3268 37365 3284 37399
rect 3218 37330 3284 37365
rect 3314 37399 3380 37434
rect 3314 37365 3330 37399
rect 3364 37365 3380 37399
rect 3314 37330 3380 37365
rect 3410 37399 3472 37434
rect 3410 37365 3426 37399
rect 3460 37365 3472 37399
rect 3410 37330 3472 37365
rect 3635 37426 3693 37438
rect 3635 37350 3647 37426
rect 3681 37350 3693 37426
rect 3635 37338 3693 37350
rect 3723 37426 3781 37438
rect 3723 37350 3735 37426
rect 3769 37350 3781 37426
rect 3723 37338 3781 37350
rect 3975 37399 4037 37434
rect 3975 37365 3987 37399
rect 4021 37365 4037 37399
rect 3975 37330 4037 37365
rect 4067 37399 4133 37434
rect 4067 37365 4083 37399
rect 4117 37365 4133 37399
rect 4067 37330 4133 37365
rect 4163 37399 4229 37434
rect 4163 37365 4179 37399
rect 4213 37365 4229 37399
rect 4163 37330 4229 37365
rect 4259 37399 4325 37434
rect 4259 37365 4275 37399
rect 4309 37365 4325 37399
rect 4259 37330 4325 37365
rect 4355 37399 4421 37434
rect 4355 37365 4371 37399
rect 4405 37365 4421 37399
rect 4355 37330 4421 37365
rect 4451 37399 4517 37434
rect 4451 37365 4467 37399
rect 4501 37365 4517 37399
rect 4451 37330 4517 37365
rect 4547 37399 4613 37434
rect 4547 37365 4563 37399
rect 4597 37365 4613 37399
rect 4547 37330 4613 37365
rect 4643 37399 4709 37434
rect 4643 37365 4659 37399
rect 4693 37365 4709 37399
rect 4643 37330 4709 37365
rect 4739 37399 4805 37434
rect 4739 37365 4755 37399
rect 4789 37365 4805 37399
rect 4739 37330 4805 37365
rect 4835 37399 4901 37434
rect 4835 37365 4851 37399
rect 4885 37365 4901 37399
rect 4835 37330 4901 37365
rect 4931 37399 4993 37434
rect 4931 37365 4947 37399
rect 4981 37365 4993 37399
rect 4931 37330 4993 37365
rect 5348 37469 5400 37481
rect 5348 37435 5356 37469
rect 5390 37435 5400 37469
rect 5348 37401 5400 37435
rect 5348 37367 5356 37401
rect 5390 37367 5400 37401
rect 5348 37351 5400 37367
rect 5430 37469 5482 37481
rect 5430 37435 5440 37469
rect 5474 37435 5482 37469
rect 5430 37401 5482 37435
rect 5430 37367 5440 37401
rect 5474 37367 5482 37401
rect 5430 37351 5482 37367
rect 301 36108 363 36143
rect 301 36074 313 36108
rect 347 36074 363 36108
rect 301 36039 363 36074
rect 393 36108 459 36143
rect 393 36074 409 36108
rect 443 36074 459 36108
rect 393 36039 459 36074
rect 489 36108 555 36143
rect 489 36074 505 36108
rect 539 36074 555 36108
rect 489 36039 555 36074
rect 585 36108 651 36143
rect 585 36074 601 36108
rect 635 36074 651 36108
rect 585 36039 651 36074
rect 681 36108 747 36143
rect 681 36074 697 36108
rect 731 36074 747 36108
rect 681 36039 747 36074
rect 777 36108 843 36143
rect 777 36074 793 36108
rect 827 36074 843 36108
rect 777 36039 843 36074
rect 873 36108 939 36143
rect 873 36074 889 36108
rect 923 36074 939 36108
rect 873 36039 939 36074
rect 969 36108 1035 36143
rect 969 36074 985 36108
rect 1019 36074 1035 36108
rect 969 36039 1035 36074
rect 1065 36108 1131 36143
rect 1065 36074 1081 36108
rect 1115 36074 1131 36108
rect 1065 36039 1131 36074
rect 1161 36108 1227 36143
rect 1161 36074 1177 36108
rect 1211 36074 1227 36108
rect 1161 36039 1227 36074
rect 1257 36108 1319 36143
rect 1257 36074 1273 36108
rect 1307 36074 1319 36108
rect 1257 36039 1319 36074
rect 2454 36112 2516 36147
rect 2454 36078 2466 36112
rect 2500 36078 2516 36112
rect 2454 36043 2516 36078
rect 2546 36112 2612 36147
rect 2546 36078 2562 36112
rect 2596 36078 2612 36112
rect 2546 36043 2612 36078
rect 2642 36112 2708 36147
rect 2642 36078 2658 36112
rect 2692 36078 2708 36112
rect 2642 36043 2708 36078
rect 2738 36112 2804 36147
rect 2738 36078 2754 36112
rect 2788 36078 2804 36112
rect 2738 36043 2804 36078
rect 2834 36112 2900 36147
rect 2834 36078 2850 36112
rect 2884 36078 2900 36112
rect 2834 36043 2900 36078
rect 2930 36112 2996 36147
rect 2930 36078 2946 36112
rect 2980 36078 2996 36112
rect 2930 36043 2996 36078
rect 3026 36112 3092 36147
rect 3026 36078 3042 36112
rect 3076 36078 3092 36112
rect 3026 36043 3092 36078
rect 3122 36112 3188 36147
rect 3122 36078 3138 36112
rect 3172 36078 3188 36112
rect 3122 36043 3188 36078
rect 3218 36112 3284 36147
rect 3218 36078 3234 36112
rect 3268 36078 3284 36112
rect 3218 36043 3284 36078
rect 3314 36112 3380 36147
rect 3314 36078 3330 36112
rect 3364 36078 3380 36112
rect 3314 36043 3380 36078
rect 3410 36112 3472 36147
rect 3410 36078 3426 36112
rect 3460 36078 3472 36112
rect 3410 36043 3472 36078
rect 3635 36139 3693 36151
rect 3635 36063 3647 36139
rect 3681 36063 3693 36139
rect 3635 36051 3693 36063
rect 3723 36139 3781 36151
rect 3723 36063 3735 36139
rect 3769 36063 3781 36139
rect 3723 36051 3781 36063
rect 3975 36112 4037 36147
rect 3975 36078 3987 36112
rect 4021 36078 4037 36112
rect 3975 36043 4037 36078
rect 4067 36112 4133 36147
rect 4067 36078 4083 36112
rect 4117 36078 4133 36112
rect 4067 36043 4133 36078
rect 4163 36112 4229 36147
rect 4163 36078 4179 36112
rect 4213 36078 4229 36112
rect 4163 36043 4229 36078
rect 4259 36112 4325 36147
rect 4259 36078 4275 36112
rect 4309 36078 4325 36112
rect 4259 36043 4325 36078
rect 4355 36112 4421 36147
rect 4355 36078 4371 36112
rect 4405 36078 4421 36112
rect 4355 36043 4421 36078
rect 4451 36112 4517 36147
rect 4451 36078 4467 36112
rect 4501 36078 4517 36112
rect 4451 36043 4517 36078
rect 4547 36112 4613 36147
rect 4547 36078 4563 36112
rect 4597 36078 4613 36112
rect 4547 36043 4613 36078
rect 4643 36112 4709 36147
rect 4643 36078 4659 36112
rect 4693 36078 4709 36112
rect 4643 36043 4709 36078
rect 4739 36112 4805 36147
rect 4739 36078 4755 36112
rect 4789 36078 4805 36112
rect 4739 36043 4805 36078
rect 4835 36112 4901 36147
rect 4835 36078 4851 36112
rect 4885 36078 4901 36112
rect 4835 36043 4901 36078
rect 4931 36112 4993 36147
rect 4931 36078 4947 36112
rect 4981 36078 4993 36112
rect 4931 36043 4993 36078
rect 5348 36182 5400 36194
rect 5348 36148 5356 36182
rect 5390 36148 5400 36182
rect 5348 36114 5400 36148
rect 5348 36080 5356 36114
rect 5390 36080 5400 36114
rect 5348 36064 5400 36080
rect 5430 36182 5482 36194
rect 5430 36148 5440 36182
rect 5474 36148 5482 36182
rect 5430 36114 5482 36148
rect 5430 36080 5440 36114
rect 5474 36080 5482 36114
rect 5430 36064 5482 36080
rect 301 34821 363 34856
rect 301 34787 313 34821
rect 347 34787 363 34821
rect 301 34752 363 34787
rect 393 34821 459 34856
rect 393 34787 409 34821
rect 443 34787 459 34821
rect 393 34752 459 34787
rect 489 34821 555 34856
rect 489 34787 505 34821
rect 539 34787 555 34821
rect 489 34752 555 34787
rect 585 34821 651 34856
rect 585 34787 601 34821
rect 635 34787 651 34821
rect 585 34752 651 34787
rect 681 34821 747 34856
rect 681 34787 697 34821
rect 731 34787 747 34821
rect 681 34752 747 34787
rect 777 34821 843 34856
rect 777 34787 793 34821
rect 827 34787 843 34821
rect 777 34752 843 34787
rect 873 34821 939 34856
rect 873 34787 889 34821
rect 923 34787 939 34821
rect 873 34752 939 34787
rect 969 34821 1035 34856
rect 969 34787 985 34821
rect 1019 34787 1035 34821
rect 969 34752 1035 34787
rect 1065 34821 1131 34856
rect 1065 34787 1081 34821
rect 1115 34787 1131 34821
rect 1065 34752 1131 34787
rect 1161 34821 1227 34856
rect 1161 34787 1177 34821
rect 1211 34787 1227 34821
rect 1161 34752 1227 34787
rect 1257 34821 1319 34856
rect 1257 34787 1273 34821
rect 1307 34787 1319 34821
rect 1257 34752 1319 34787
rect 2454 34825 2516 34860
rect 2454 34791 2466 34825
rect 2500 34791 2516 34825
rect 2454 34756 2516 34791
rect 2546 34825 2612 34860
rect 2546 34791 2562 34825
rect 2596 34791 2612 34825
rect 2546 34756 2612 34791
rect 2642 34825 2708 34860
rect 2642 34791 2658 34825
rect 2692 34791 2708 34825
rect 2642 34756 2708 34791
rect 2738 34825 2804 34860
rect 2738 34791 2754 34825
rect 2788 34791 2804 34825
rect 2738 34756 2804 34791
rect 2834 34825 2900 34860
rect 2834 34791 2850 34825
rect 2884 34791 2900 34825
rect 2834 34756 2900 34791
rect 2930 34825 2996 34860
rect 2930 34791 2946 34825
rect 2980 34791 2996 34825
rect 2930 34756 2996 34791
rect 3026 34825 3092 34860
rect 3026 34791 3042 34825
rect 3076 34791 3092 34825
rect 3026 34756 3092 34791
rect 3122 34825 3188 34860
rect 3122 34791 3138 34825
rect 3172 34791 3188 34825
rect 3122 34756 3188 34791
rect 3218 34825 3284 34860
rect 3218 34791 3234 34825
rect 3268 34791 3284 34825
rect 3218 34756 3284 34791
rect 3314 34825 3380 34860
rect 3314 34791 3330 34825
rect 3364 34791 3380 34825
rect 3314 34756 3380 34791
rect 3410 34825 3472 34860
rect 3410 34791 3426 34825
rect 3460 34791 3472 34825
rect 3410 34756 3472 34791
rect 3635 34852 3693 34864
rect 3635 34776 3647 34852
rect 3681 34776 3693 34852
rect 3635 34764 3693 34776
rect 3723 34852 3781 34864
rect 3723 34776 3735 34852
rect 3769 34776 3781 34852
rect 3723 34764 3781 34776
rect 3975 34825 4037 34860
rect 3975 34791 3987 34825
rect 4021 34791 4037 34825
rect 3975 34756 4037 34791
rect 4067 34825 4133 34860
rect 4067 34791 4083 34825
rect 4117 34791 4133 34825
rect 4067 34756 4133 34791
rect 4163 34825 4229 34860
rect 4163 34791 4179 34825
rect 4213 34791 4229 34825
rect 4163 34756 4229 34791
rect 4259 34825 4325 34860
rect 4259 34791 4275 34825
rect 4309 34791 4325 34825
rect 4259 34756 4325 34791
rect 4355 34825 4421 34860
rect 4355 34791 4371 34825
rect 4405 34791 4421 34825
rect 4355 34756 4421 34791
rect 4451 34825 4517 34860
rect 4451 34791 4467 34825
rect 4501 34791 4517 34825
rect 4451 34756 4517 34791
rect 4547 34825 4613 34860
rect 4547 34791 4563 34825
rect 4597 34791 4613 34825
rect 4547 34756 4613 34791
rect 4643 34825 4709 34860
rect 4643 34791 4659 34825
rect 4693 34791 4709 34825
rect 4643 34756 4709 34791
rect 4739 34825 4805 34860
rect 4739 34791 4755 34825
rect 4789 34791 4805 34825
rect 4739 34756 4805 34791
rect 4835 34825 4901 34860
rect 4835 34791 4851 34825
rect 4885 34791 4901 34825
rect 4835 34756 4901 34791
rect 4931 34825 4993 34860
rect 4931 34791 4947 34825
rect 4981 34791 4993 34825
rect 4931 34756 4993 34791
rect 5348 34895 5400 34907
rect 5348 34861 5356 34895
rect 5390 34861 5400 34895
rect 5348 34827 5400 34861
rect 5348 34793 5356 34827
rect 5390 34793 5400 34827
rect 5348 34777 5400 34793
rect 5430 34895 5482 34907
rect 5430 34861 5440 34895
rect 5474 34861 5482 34895
rect 5430 34827 5482 34861
rect 5430 34793 5440 34827
rect 5474 34793 5482 34827
rect 5430 34777 5482 34793
rect 301 33534 363 33569
rect 301 33500 313 33534
rect 347 33500 363 33534
rect 301 33465 363 33500
rect 393 33534 459 33569
rect 393 33500 409 33534
rect 443 33500 459 33534
rect 393 33465 459 33500
rect 489 33534 555 33569
rect 489 33500 505 33534
rect 539 33500 555 33534
rect 489 33465 555 33500
rect 585 33534 651 33569
rect 585 33500 601 33534
rect 635 33500 651 33534
rect 585 33465 651 33500
rect 681 33534 747 33569
rect 681 33500 697 33534
rect 731 33500 747 33534
rect 681 33465 747 33500
rect 777 33534 843 33569
rect 777 33500 793 33534
rect 827 33500 843 33534
rect 777 33465 843 33500
rect 873 33534 939 33569
rect 873 33500 889 33534
rect 923 33500 939 33534
rect 873 33465 939 33500
rect 969 33534 1035 33569
rect 969 33500 985 33534
rect 1019 33500 1035 33534
rect 969 33465 1035 33500
rect 1065 33534 1131 33569
rect 1065 33500 1081 33534
rect 1115 33500 1131 33534
rect 1065 33465 1131 33500
rect 1161 33534 1227 33569
rect 1161 33500 1177 33534
rect 1211 33500 1227 33534
rect 1161 33465 1227 33500
rect 1257 33534 1319 33569
rect 1257 33500 1273 33534
rect 1307 33500 1319 33534
rect 1257 33465 1319 33500
rect 2454 33538 2516 33573
rect 2454 33504 2466 33538
rect 2500 33504 2516 33538
rect 2454 33469 2516 33504
rect 2546 33538 2612 33573
rect 2546 33504 2562 33538
rect 2596 33504 2612 33538
rect 2546 33469 2612 33504
rect 2642 33538 2708 33573
rect 2642 33504 2658 33538
rect 2692 33504 2708 33538
rect 2642 33469 2708 33504
rect 2738 33538 2804 33573
rect 2738 33504 2754 33538
rect 2788 33504 2804 33538
rect 2738 33469 2804 33504
rect 2834 33538 2900 33573
rect 2834 33504 2850 33538
rect 2884 33504 2900 33538
rect 2834 33469 2900 33504
rect 2930 33538 2996 33573
rect 2930 33504 2946 33538
rect 2980 33504 2996 33538
rect 2930 33469 2996 33504
rect 3026 33538 3092 33573
rect 3026 33504 3042 33538
rect 3076 33504 3092 33538
rect 3026 33469 3092 33504
rect 3122 33538 3188 33573
rect 3122 33504 3138 33538
rect 3172 33504 3188 33538
rect 3122 33469 3188 33504
rect 3218 33538 3284 33573
rect 3218 33504 3234 33538
rect 3268 33504 3284 33538
rect 3218 33469 3284 33504
rect 3314 33538 3380 33573
rect 3314 33504 3330 33538
rect 3364 33504 3380 33538
rect 3314 33469 3380 33504
rect 3410 33538 3472 33573
rect 3410 33504 3426 33538
rect 3460 33504 3472 33538
rect 3410 33469 3472 33504
rect 3635 33565 3693 33577
rect 3635 33489 3647 33565
rect 3681 33489 3693 33565
rect 3635 33477 3693 33489
rect 3723 33565 3781 33577
rect 3723 33489 3735 33565
rect 3769 33489 3781 33565
rect 3723 33477 3781 33489
rect 3975 33538 4037 33573
rect 3975 33504 3987 33538
rect 4021 33504 4037 33538
rect 3975 33469 4037 33504
rect 4067 33538 4133 33573
rect 4067 33504 4083 33538
rect 4117 33504 4133 33538
rect 4067 33469 4133 33504
rect 4163 33538 4229 33573
rect 4163 33504 4179 33538
rect 4213 33504 4229 33538
rect 4163 33469 4229 33504
rect 4259 33538 4325 33573
rect 4259 33504 4275 33538
rect 4309 33504 4325 33538
rect 4259 33469 4325 33504
rect 4355 33538 4421 33573
rect 4355 33504 4371 33538
rect 4405 33504 4421 33538
rect 4355 33469 4421 33504
rect 4451 33538 4517 33573
rect 4451 33504 4467 33538
rect 4501 33504 4517 33538
rect 4451 33469 4517 33504
rect 4547 33538 4613 33573
rect 4547 33504 4563 33538
rect 4597 33504 4613 33538
rect 4547 33469 4613 33504
rect 4643 33538 4709 33573
rect 4643 33504 4659 33538
rect 4693 33504 4709 33538
rect 4643 33469 4709 33504
rect 4739 33538 4805 33573
rect 4739 33504 4755 33538
rect 4789 33504 4805 33538
rect 4739 33469 4805 33504
rect 4835 33538 4901 33573
rect 4835 33504 4851 33538
rect 4885 33504 4901 33538
rect 4835 33469 4901 33504
rect 4931 33538 4993 33573
rect 4931 33504 4947 33538
rect 4981 33504 4993 33538
rect 4931 33469 4993 33504
rect 5348 33608 5400 33620
rect 5348 33574 5356 33608
rect 5390 33574 5400 33608
rect 5348 33540 5400 33574
rect 5348 33506 5356 33540
rect 5390 33506 5400 33540
rect 5348 33490 5400 33506
rect 5430 33608 5482 33620
rect 5430 33574 5440 33608
rect 5474 33574 5482 33608
rect 5430 33540 5482 33574
rect 5430 33506 5440 33540
rect 5474 33506 5482 33540
rect 5430 33490 5482 33506
rect 301 32247 363 32282
rect 301 32213 313 32247
rect 347 32213 363 32247
rect 301 32178 363 32213
rect 393 32247 459 32282
rect 393 32213 409 32247
rect 443 32213 459 32247
rect 393 32178 459 32213
rect 489 32247 555 32282
rect 489 32213 505 32247
rect 539 32213 555 32247
rect 489 32178 555 32213
rect 585 32247 651 32282
rect 585 32213 601 32247
rect 635 32213 651 32247
rect 585 32178 651 32213
rect 681 32247 747 32282
rect 681 32213 697 32247
rect 731 32213 747 32247
rect 681 32178 747 32213
rect 777 32247 843 32282
rect 777 32213 793 32247
rect 827 32213 843 32247
rect 777 32178 843 32213
rect 873 32247 939 32282
rect 873 32213 889 32247
rect 923 32213 939 32247
rect 873 32178 939 32213
rect 969 32247 1035 32282
rect 969 32213 985 32247
rect 1019 32213 1035 32247
rect 969 32178 1035 32213
rect 1065 32247 1131 32282
rect 1065 32213 1081 32247
rect 1115 32213 1131 32247
rect 1065 32178 1131 32213
rect 1161 32247 1227 32282
rect 1161 32213 1177 32247
rect 1211 32213 1227 32247
rect 1161 32178 1227 32213
rect 1257 32247 1319 32282
rect 1257 32213 1273 32247
rect 1307 32213 1319 32247
rect 1257 32178 1319 32213
rect 2454 32251 2516 32286
rect 2454 32217 2466 32251
rect 2500 32217 2516 32251
rect 2454 32182 2516 32217
rect 2546 32251 2612 32286
rect 2546 32217 2562 32251
rect 2596 32217 2612 32251
rect 2546 32182 2612 32217
rect 2642 32251 2708 32286
rect 2642 32217 2658 32251
rect 2692 32217 2708 32251
rect 2642 32182 2708 32217
rect 2738 32251 2804 32286
rect 2738 32217 2754 32251
rect 2788 32217 2804 32251
rect 2738 32182 2804 32217
rect 2834 32251 2900 32286
rect 2834 32217 2850 32251
rect 2884 32217 2900 32251
rect 2834 32182 2900 32217
rect 2930 32251 2996 32286
rect 2930 32217 2946 32251
rect 2980 32217 2996 32251
rect 2930 32182 2996 32217
rect 3026 32251 3092 32286
rect 3026 32217 3042 32251
rect 3076 32217 3092 32251
rect 3026 32182 3092 32217
rect 3122 32251 3188 32286
rect 3122 32217 3138 32251
rect 3172 32217 3188 32251
rect 3122 32182 3188 32217
rect 3218 32251 3284 32286
rect 3218 32217 3234 32251
rect 3268 32217 3284 32251
rect 3218 32182 3284 32217
rect 3314 32251 3380 32286
rect 3314 32217 3330 32251
rect 3364 32217 3380 32251
rect 3314 32182 3380 32217
rect 3410 32251 3472 32286
rect 3410 32217 3426 32251
rect 3460 32217 3472 32251
rect 3410 32182 3472 32217
rect 3635 32278 3693 32290
rect 3635 32202 3647 32278
rect 3681 32202 3693 32278
rect 3635 32190 3693 32202
rect 3723 32278 3781 32290
rect 3723 32202 3735 32278
rect 3769 32202 3781 32278
rect 3723 32190 3781 32202
rect 3975 32251 4037 32286
rect 3975 32217 3987 32251
rect 4021 32217 4037 32251
rect 3975 32182 4037 32217
rect 4067 32251 4133 32286
rect 4067 32217 4083 32251
rect 4117 32217 4133 32251
rect 4067 32182 4133 32217
rect 4163 32251 4229 32286
rect 4163 32217 4179 32251
rect 4213 32217 4229 32251
rect 4163 32182 4229 32217
rect 4259 32251 4325 32286
rect 4259 32217 4275 32251
rect 4309 32217 4325 32251
rect 4259 32182 4325 32217
rect 4355 32251 4421 32286
rect 4355 32217 4371 32251
rect 4405 32217 4421 32251
rect 4355 32182 4421 32217
rect 4451 32251 4517 32286
rect 4451 32217 4467 32251
rect 4501 32217 4517 32251
rect 4451 32182 4517 32217
rect 4547 32251 4613 32286
rect 4547 32217 4563 32251
rect 4597 32217 4613 32251
rect 4547 32182 4613 32217
rect 4643 32251 4709 32286
rect 4643 32217 4659 32251
rect 4693 32217 4709 32251
rect 4643 32182 4709 32217
rect 4739 32251 4805 32286
rect 4739 32217 4755 32251
rect 4789 32217 4805 32251
rect 4739 32182 4805 32217
rect 4835 32251 4901 32286
rect 4835 32217 4851 32251
rect 4885 32217 4901 32251
rect 4835 32182 4901 32217
rect 4931 32251 4993 32286
rect 4931 32217 4947 32251
rect 4981 32217 4993 32251
rect 4931 32182 4993 32217
rect 5348 32321 5400 32333
rect 5348 32287 5356 32321
rect 5390 32287 5400 32321
rect 5348 32253 5400 32287
rect 5348 32219 5356 32253
rect 5390 32219 5400 32253
rect 5348 32203 5400 32219
rect 5430 32321 5482 32333
rect 5430 32287 5440 32321
rect 5474 32287 5482 32321
rect 5430 32253 5482 32287
rect 5430 32219 5440 32253
rect 5474 32219 5482 32253
rect 5430 32203 5482 32219
rect 301 30960 363 30995
rect 301 30926 313 30960
rect 347 30926 363 30960
rect 301 30891 363 30926
rect 393 30960 459 30995
rect 393 30926 409 30960
rect 443 30926 459 30960
rect 393 30891 459 30926
rect 489 30960 555 30995
rect 489 30926 505 30960
rect 539 30926 555 30960
rect 489 30891 555 30926
rect 585 30960 651 30995
rect 585 30926 601 30960
rect 635 30926 651 30960
rect 585 30891 651 30926
rect 681 30960 747 30995
rect 681 30926 697 30960
rect 731 30926 747 30960
rect 681 30891 747 30926
rect 777 30960 843 30995
rect 777 30926 793 30960
rect 827 30926 843 30960
rect 777 30891 843 30926
rect 873 30960 939 30995
rect 873 30926 889 30960
rect 923 30926 939 30960
rect 873 30891 939 30926
rect 969 30960 1035 30995
rect 969 30926 985 30960
rect 1019 30926 1035 30960
rect 969 30891 1035 30926
rect 1065 30960 1131 30995
rect 1065 30926 1081 30960
rect 1115 30926 1131 30960
rect 1065 30891 1131 30926
rect 1161 30960 1227 30995
rect 1161 30926 1177 30960
rect 1211 30926 1227 30960
rect 1161 30891 1227 30926
rect 1257 30960 1319 30995
rect 1257 30926 1273 30960
rect 1307 30926 1319 30960
rect 1257 30891 1319 30926
rect 2454 30964 2516 30999
rect 2454 30930 2466 30964
rect 2500 30930 2516 30964
rect 2454 30895 2516 30930
rect 2546 30964 2612 30999
rect 2546 30930 2562 30964
rect 2596 30930 2612 30964
rect 2546 30895 2612 30930
rect 2642 30964 2708 30999
rect 2642 30930 2658 30964
rect 2692 30930 2708 30964
rect 2642 30895 2708 30930
rect 2738 30964 2804 30999
rect 2738 30930 2754 30964
rect 2788 30930 2804 30964
rect 2738 30895 2804 30930
rect 2834 30964 2900 30999
rect 2834 30930 2850 30964
rect 2884 30930 2900 30964
rect 2834 30895 2900 30930
rect 2930 30964 2996 30999
rect 2930 30930 2946 30964
rect 2980 30930 2996 30964
rect 2930 30895 2996 30930
rect 3026 30964 3092 30999
rect 3026 30930 3042 30964
rect 3076 30930 3092 30964
rect 3026 30895 3092 30930
rect 3122 30964 3188 30999
rect 3122 30930 3138 30964
rect 3172 30930 3188 30964
rect 3122 30895 3188 30930
rect 3218 30964 3284 30999
rect 3218 30930 3234 30964
rect 3268 30930 3284 30964
rect 3218 30895 3284 30930
rect 3314 30964 3380 30999
rect 3314 30930 3330 30964
rect 3364 30930 3380 30964
rect 3314 30895 3380 30930
rect 3410 30964 3472 30999
rect 3410 30930 3426 30964
rect 3460 30930 3472 30964
rect 3410 30895 3472 30930
rect 3635 30991 3693 31003
rect 3635 30915 3647 30991
rect 3681 30915 3693 30991
rect 3635 30903 3693 30915
rect 3723 30991 3781 31003
rect 3723 30915 3735 30991
rect 3769 30915 3781 30991
rect 3723 30903 3781 30915
rect 3975 30964 4037 30999
rect 3975 30930 3987 30964
rect 4021 30930 4037 30964
rect 3975 30895 4037 30930
rect 4067 30964 4133 30999
rect 4067 30930 4083 30964
rect 4117 30930 4133 30964
rect 4067 30895 4133 30930
rect 4163 30964 4229 30999
rect 4163 30930 4179 30964
rect 4213 30930 4229 30964
rect 4163 30895 4229 30930
rect 4259 30964 4325 30999
rect 4259 30930 4275 30964
rect 4309 30930 4325 30964
rect 4259 30895 4325 30930
rect 4355 30964 4421 30999
rect 4355 30930 4371 30964
rect 4405 30930 4421 30964
rect 4355 30895 4421 30930
rect 4451 30964 4517 30999
rect 4451 30930 4467 30964
rect 4501 30930 4517 30964
rect 4451 30895 4517 30930
rect 4547 30964 4613 30999
rect 4547 30930 4563 30964
rect 4597 30930 4613 30964
rect 4547 30895 4613 30930
rect 4643 30964 4709 30999
rect 4643 30930 4659 30964
rect 4693 30930 4709 30964
rect 4643 30895 4709 30930
rect 4739 30964 4805 30999
rect 4739 30930 4755 30964
rect 4789 30930 4805 30964
rect 4739 30895 4805 30930
rect 4835 30964 4901 30999
rect 4835 30930 4851 30964
rect 4885 30930 4901 30964
rect 4835 30895 4901 30930
rect 4931 30964 4993 30999
rect 4931 30930 4947 30964
rect 4981 30930 4993 30964
rect 4931 30895 4993 30930
rect 5348 31034 5400 31046
rect 5348 31000 5356 31034
rect 5390 31000 5400 31034
rect 5348 30966 5400 31000
rect 5348 30932 5356 30966
rect 5390 30932 5400 30966
rect 5348 30916 5400 30932
rect 5430 31034 5482 31046
rect 5430 31000 5440 31034
rect 5474 31000 5482 31034
rect 5430 30966 5482 31000
rect 5430 30932 5440 30966
rect 5474 30932 5482 30966
rect 5430 30916 5482 30932
rect 301 29673 363 29708
rect 301 29639 313 29673
rect 347 29639 363 29673
rect 301 29604 363 29639
rect 393 29673 459 29708
rect 393 29639 409 29673
rect 443 29639 459 29673
rect 393 29604 459 29639
rect 489 29673 555 29708
rect 489 29639 505 29673
rect 539 29639 555 29673
rect 489 29604 555 29639
rect 585 29673 651 29708
rect 585 29639 601 29673
rect 635 29639 651 29673
rect 585 29604 651 29639
rect 681 29673 747 29708
rect 681 29639 697 29673
rect 731 29639 747 29673
rect 681 29604 747 29639
rect 777 29673 843 29708
rect 777 29639 793 29673
rect 827 29639 843 29673
rect 777 29604 843 29639
rect 873 29673 939 29708
rect 873 29639 889 29673
rect 923 29639 939 29673
rect 873 29604 939 29639
rect 969 29673 1035 29708
rect 969 29639 985 29673
rect 1019 29639 1035 29673
rect 969 29604 1035 29639
rect 1065 29673 1131 29708
rect 1065 29639 1081 29673
rect 1115 29639 1131 29673
rect 1065 29604 1131 29639
rect 1161 29673 1227 29708
rect 1161 29639 1177 29673
rect 1211 29639 1227 29673
rect 1161 29604 1227 29639
rect 1257 29673 1319 29708
rect 1257 29639 1273 29673
rect 1307 29639 1319 29673
rect 1257 29604 1319 29639
rect 2454 29677 2516 29712
rect 2454 29643 2466 29677
rect 2500 29643 2516 29677
rect 2454 29608 2516 29643
rect 2546 29677 2612 29712
rect 2546 29643 2562 29677
rect 2596 29643 2612 29677
rect 2546 29608 2612 29643
rect 2642 29677 2708 29712
rect 2642 29643 2658 29677
rect 2692 29643 2708 29677
rect 2642 29608 2708 29643
rect 2738 29677 2804 29712
rect 2738 29643 2754 29677
rect 2788 29643 2804 29677
rect 2738 29608 2804 29643
rect 2834 29677 2900 29712
rect 2834 29643 2850 29677
rect 2884 29643 2900 29677
rect 2834 29608 2900 29643
rect 2930 29677 2996 29712
rect 2930 29643 2946 29677
rect 2980 29643 2996 29677
rect 2930 29608 2996 29643
rect 3026 29677 3092 29712
rect 3026 29643 3042 29677
rect 3076 29643 3092 29677
rect 3026 29608 3092 29643
rect 3122 29677 3188 29712
rect 3122 29643 3138 29677
rect 3172 29643 3188 29677
rect 3122 29608 3188 29643
rect 3218 29677 3284 29712
rect 3218 29643 3234 29677
rect 3268 29643 3284 29677
rect 3218 29608 3284 29643
rect 3314 29677 3380 29712
rect 3314 29643 3330 29677
rect 3364 29643 3380 29677
rect 3314 29608 3380 29643
rect 3410 29677 3472 29712
rect 3410 29643 3426 29677
rect 3460 29643 3472 29677
rect 3410 29608 3472 29643
rect 3635 29704 3693 29716
rect 3635 29628 3647 29704
rect 3681 29628 3693 29704
rect 3635 29616 3693 29628
rect 3723 29704 3781 29716
rect 3723 29628 3735 29704
rect 3769 29628 3781 29704
rect 3723 29616 3781 29628
rect 3975 29677 4037 29712
rect 3975 29643 3987 29677
rect 4021 29643 4037 29677
rect 3975 29608 4037 29643
rect 4067 29677 4133 29712
rect 4067 29643 4083 29677
rect 4117 29643 4133 29677
rect 4067 29608 4133 29643
rect 4163 29677 4229 29712
rect 4163 29643 4179 29677
rect 4213 29643 4229 29677
rect 4163 29608 4229 29643
rect 4259 29677 4325 29712
rect 4259 29643 4275 29677
rect 4309 29643 4325 29677
rect 4259 29608 4325 29643
rect 4355 29677 4421 29712
rect 4355 29643 4371 29677
rect 4405 29643 4421 29677
rect 4355 29608 4421 29643
rect 4451 29677 4517 29712
rect 4451 29643 4467 29677
rect 4501 29643 4517 29677
rect 4451 29608 4517 29643
rect 4547 29677 4613 29712
rect 4547 29643 4563 29677
rect 4597 29643 4613 29677
rect 4547 29608 4613 29643
rect 4643 29677 4709 29712
rect 4643 29643 4659 29677
rect 4693 29643 4709 29677
rect 4643 29608 4709 29643
rect 4739 29677 4805 29712
rect 4739 29643 4755 29677
rect 4789 29643 4805 29677
rect 4739 29608 4805 29643
rect 4835 29677 4901 29712
rect 4835 29643 4851 29677
rect 4885 29643 4901 29677
rect 4835 29608 4901 29643
rect 4931 29677 4993 29712
rect 4931 29643 4947 29677
rect 4981 29643 4993 29677
rect 4931 29608 4993 29643
rect 5348 29747 5400 29759
rect 5348 29713 5356 29747
rect 5390 29713 5400 29747
rect 5348 29679 5400 29713
rect 5348 29645 5356 29679
rect 5390 29645 5400 29679
rect 5348 29629 5400 29645
rect 5430 29747 5482 29759
rect 5430 29713 5440 29747
rect 5474 29713 5482 29747
rect 5430 29679 5482 29713
rect 5430 29645 5440 29679
rect 5474 29645 5482 29679
rect 5430 29629 5482 29645
rect 301 28386 363 28421
rect 301 28352 313 28386
rect 347 28352 363 28386
rect 301 28317 363 28352
rect 393 28386 459 28421
rect 393 28352 409 28386
rect 443 28352 459 28386
rect 393 28317 459 28352
rect 489 28386 555 28421
rect 489 28352 505 28386
rect 539 28352 555 28386
rect 489 28317 555 28352
rect 585 28386 651 28421
rect 585 28352 601 28386
rect 635 28352 651 28386
rect 585 28317 651 28352
rect 681 28386 747 28421
rect 681 28352 697 28386
rect 731 28352 747 28386
rect 681 28317 747 28352
rect 777 28386 843 28421
rect 777 28352 793 28386
rect 827 28352 843 28386
rect 777 28317 843 28352
rect 873 28386 939 28421
rect 873 28352 889 28386
rect 923 28352 939 28386
rect 873 28317 939 28352
rect 969 28386 1035 28421
rect 969 28352 985 28386
rect 1019 28352 1035 28386
rect 969 28317 1035 28352
rect 1065 28386 1131 28421
rect 1065 28352 1081 28386
rect 1115 28352 1131 28386
rect 1065 28317 1131 28352
rect 1161 28386 1227 28421
rect 1161 28352 1177 28386
rect 1211 28352 1227 28386
rect 1161 28317 1227 28352
rect 1257 28386 1319 28421
rect 1257 28352 1273 28386
rect 1307 28352 1319 28386
rect 1257 28317 1319 28352
rect 2454 28390 2516 28425
rect 2454 28356 2466 28390
rect 2500 28356 2516 28390
rect 2454 28321 2516 28356
rect 2546 28390 2612 28425
rect 2546 28356 2562 28390
rect 2596 28356 2612 28390
rect 2546 28321 2612 28356
rect 2642 28390 2708 28425
rect 2642 28356 2658 28390
rect 2692 28356 2708 28390
rect 2642 28321 2708 28356
rect 2738 28390 2804 28425
rect 2738 28356 2754 28390
rect 2788 28356 2804 28390
rect 2738 28321 2804 28356
rect 2834 28390 2900 28425
rect 2834 28356 2850 28390
rect 2884 28356 2900 28390
rect 2834 28321 2900 28356
rect 2930 28390 2996 28425
rect 2930 28356 2946 28390
rect 2980 28356 2996 28390
rect 2930 28321 2996 28356
rect 3026 28390 3092 28425
rect 3026 28356 3042 28390
rect 3076 28356 3092 28390
rect 3026 28321 3092 28356
rect 3122 28390 3188 28425
rect 3122 28356 3138 28390
rect 3172 28356 3188 28390
rect 3122 28321 3188 28356
rect 3218 28390 3284 28425
rect 3218 28356 3234 28390
rect 3268 28356 3284 28390
rect 3218 28321 3284 28356
rect 3314 28390 3380 28425
rect 3314 28356 3330 28390
rect 3364 28356 3380 28390
rect 3314 28321 3380 28356
rect 3410 28390 3472 28425
rect 3410 28356 3426 28390
rect 3460 28356 3472 28390
rect 3410 28321 3472 28356
rect 3635 28417 3693 28429
rect 3635 28341 3647 28417
rect 3681 28341 3693 28417
rect 3635 28329 3693 28341
rect 3723 28417 3781 28429
rect 3723 28341 3735 28417
rect 3769 28341 3781 28417
rect 3723 28329 3781 28341
rect 3975 28390 4037 28425
rect 3975 28356 3987 28390
rect 4021 28356 4037 28390
rect 3975 28321 4037 28356
rect 4067 28390 4133 28425
rect 4067 28356 4083 28390
rect 4117 28356 4133 28390
rect 4067 28321 4133 28356
rect 4163 28390 4229 28425
rect 4163 28356 4179 28390
rect 4213 28356 4229 28390
rect 4163 28321 4229 28356
rect 4259 28390 4325 28425
rect 4259 28356 4275 28390
rect 4309 28356 4325 28390
rect 4259 28321 4325 28356
rect 4355 28390 4421 28425
rect 4355 28356 4371 28390
rect 4405 28356 4421 28390
rect 4355 28321 4421 28356
rect 4451 28390 4517 28425
rect 4451 28356 4467 28390
rect 4501 28356 4517 28390
rect 4451 28321 4517 28356
rect 4547 28390 4613 28425
rect 4547 28356 4563 28390
rect 4597 28356 4613 28390
rect 4547 28321 4613 28356
rect 4643 28390 4709 28425
rect 4643 28356 4659 28390
rect 4693 28356 4709 28390
rect 4643 28321 4709 28356
rect 4739 28390 4805 28425
rect 4739 28356 4755 28390
rect 4789 28356 4805 28390
rect 4739 28321 4805 28356
rect 4835 28390 4901 28425
rect 4835 28356 4851 28390
rect 4885 28356 4901 28390
rect 4835 28321 4901 28356
rect 4931 28390 4993 28425
rect 4931 28356 4947 28390
rect 4981 28356 4993 28390
rect 4931 28321 4993 28356
rect 5348 28460 5400 28472
rect 5348 28426 5356 28460
rect 5390 28426 5400 28460
rect 5348 28392 5400 28426
rect 5348 28358 5356 28392
rect 5390 28358 5400 28392
rect 5348 28342 5400 28358
rect 5430 28460 5482 28472
rect 5430 28426 5440 28460
rect 5474 28426 5482 28460
rect 5430 28392 5482 28426
rect 5430 28358 5440 28392
rect 5474 28358 5482 28392
rect 5430 28342 5482 28358
rect 301 27099 363 27134
rect 301 27065 313 27099
rect 347 27065 363 27099
rect 301 27030 363 27065
rect 393 27099 459 27134
rect 393 27065 409 27099
rect 443 27065 459 27099
rect 393 27030 459 27065
rect 489 27099 555 27134
rect 489 27065 505 27099
rect 539 27065 555 27099
rect 489 27030 555 27065
rect 585 27099 651 27134
rect 585 27065 601 27099
rect 635 27065 651 27099
rect 585 27030 651 27065
rect 681 27099 747 27134
rect 681 27065 697 27099
rect 731 27065 747 27099
rect 681 27030 747 27065
rect 777 27099 843 27134
rect 777 27065 793 27099
rect 827 27065 843 27099
rect 777 27030 843 27065
rect 873 27099 939 27134
rect 873 27065 889 27099
rect 923 27065 939 27099
rect 873 27030 939 27065
rect 969 27099 1035 27134
rect 969 27065 985 27099
rect 1019 27065 1035 27099
rect 969 27030 1035 27065
rect 1065 27099 1131 27134
rect 1065 27065 1081 27099
rect 1115 27065 1131 27099
rect 1065 27030 1131 27065
rect 1161 27099 1227 27134
rect 1161 27065 1177 27099
rect 1211 27065 1227 27099
rect 1161 27030 1227 27065
rect 1257 27099 1319 27134
rect 1257 27065 1273 27099
rect 1307 27065 1319 27099
rect 1257 27030 1319 27065
rect 2454 27103 2516 27138
rect 2454 27069 2466 27103
rect 2500 27069 2516 27103
rect 2454 27034 2516 27069
rect 2546 27103 2612 27138
rect 2546 27069 2562 27103
rect 2596 27069 2612 27103
rect 2546 27034 2612 27069
rect 2642 27103 2708 27138
rect 2642 27069 2658 27103
rect 2692 27069 2708 27103
rect 2642 27034 2708 27069
rect 2738 27103 2804 27138
rect 2738 27069 2754 27103
rect 2788 27069 2804 27103
rect 2738 27034 2804 27069
rect 2834 27103 2900 27138
rect 2834 27069 2850 27103
rect 2884 27069 2900 27103
rect 2834 27034 2900 27069
rect 2930 27103 2996 27138
rect 2930 27069 2946 27103
rect 2980 27069 2996 27103
rect 2930 27034 2996 27069
rect 3026 27103 3092 27138
rect 3026 27069 3042 27103
rect 3076 27069 3092 27103
rect 3026 27034 3092 27069
rect 3122 27103 3188 27138
rect 3122 27069 3138 27103
rect 3172 27069 3188 27103
rect 3122 27034 3188 27069
rect 3218 27103 3284 27138
rect 3218 27069 3234 27103
rect 3268 27069 3284 27103
rect 3218 27034 3284 27069
rect 3314 27103 3380 27138
rect 3314 27069 3330 27103
rect 3364 27069 3380 27103
rect 3314 27034 3380 27069
rect 3410 27103 3472 27138
rect 3410 27069 3426 27103
rect 3460 27069 3472 27103
rect 3410 27034 3472 27069
rect 3635 27130 3693 27142
rect 3635 27054 3647 27130
rect 3681 27054 3693 27130
rect 3635 27042 3693 27054
rect 3723 27130 3781 27142
rect 3723 27054 3735 27130
rect 3769 27054 3781 27130
rect 3723 27042 3781 27054
rect 3975 27103 4037 27138
rect 3975 27069 3987 27103
rect 4021 27069 4037 27103
rect 3975 27034 4037 27069
rect 4067 27103 4133 27138
rect 4067 27069 4083 27103
rect 4117 27069 4133 27103
rect 4067 27034 4133 27069
rect 4163 27103 4229 27138
rect 4163 27069 4179 27103
rect 4213 27069 4229 27103
rect 4163 27034 4229 27069
rect 4259 27103 4325 27138
rect 4259 27069 4275 27103
rect 4309 27069 4325 27103
rect 4259 27034 4325 27069
rect 4355 27103 4421 27138
rect 4355 27069 4371 27103
rect 4405 27069 4421 27103
rect 4355 27034 4421 27069
rect 4451 27103 4517 27138
rect 4451 27069 4467 27103
rect 4501 27069 4517 27103
rect 4451 27034 4517 27069
rect 4547 27103 4613 27138
rect 4547 27069 4563 27103
rect 4597 27069 4613 27103
rect 4547 27034 4613 27069
rect 4643 27103 4709 27138
rect 4643 27069 4659 27103
rect 4693 27069 4709 27103
rect 4643 27034 4709 27069
rect 4739 27103 4805 27138
rect 4739 27069 4755 27103
rect 4789 27069 4805 27103
rect 4739 27034 4805 27069
rect 4835 27103 4901 27138
rect 4835 27069 4851 27103
rect 4885 27069 4901 27103
rect 4835 27034 4901 27069
rect 4931 27103 4993 27138
rect 4931 27069 4947 27103
rect 4981 27069 4993 27103
rect 4931 27034 4993 27069
rect 5348 27173 5400 27185
rect 5348 27139 5356 27173
rect 5390 27139 5400 27173
rect 5348 27105 5400 27139
rect 5348 27071 5356 27105
rect 5390 27071 5400 27105
rect 5348 27055 5400 27071
rect 5430 27173 5482 27185
rect 5430 27139 5440 27173
rect 5474 27139 5482 27173
rect 5430 27105 5482 27139
rect 5430 27071 5440 27105
rect 5474 27071 5482 27105
rect 5430 27055 5482 27071
rect 301 25812 363 25847
rect 301 25778 313 25812
rect 347 25778 363 25812
rect 301 25743 363 25778
rect 393 25812 459 25847
rect 393 25778 409 25812
rect 443 25778 459 25812
rect 393 25743 459 25778
rect 489 25812 555 25847
rect 489 25778 505 25812
rect 539 25778 555 25812
rect 489 25743 555 25778
rect 585 25812 651 25847
rect 585 25778 601 25812
rect 635 25778 651 25812
rect 585 25743 651 25778
rect 681 25812 747 25847
rect 681 25778 697 25812
rect 731 25778 747 25812
rect 681 25743 747 25778
rect 777 25812 843 25847
rect 777 25778 793 25812
rect 827 25778 843 25812
rect 777 25743 843 25778
rect 873 25812 939 25847
rect 873 25778 889 25812
rect 923 25778 939 25812
rect 873 25743 939 25778
rect 969 25812 1035 25847
rect 969 25778 985 25812
rect 1019 25778 1035 25812
rect 969 25743 1035 25778
rect 1065 25812 1131 25847
rect 1065 25778 1081 25812
rect 1115 25778 1131 25812
rect 1065 25743 1131 25778
rect 1161 25812 1227 25847
rect 1161 25778 1177 25812
rect 1211 25778 1227 25812
rect 1161 25743 1227 25778
rect 1257 25812 1319 25847
rect 1257 25778 1273 25812
rect 1307 25778 1319 25812
rect 1257 25743 1319 25778
rect 2454 25816 2516 25851
rect 2454 25782 2466 25816
rect 2500 25782 2516 25816
rect 2454 25747 2516 25782
rect 2546 25816 2612 25851
rect 2546 25782 2562 25816
rect 2596 25782 2612 25816
rect 2546 25747 2612 25782
rect 2642 25816 2708 25851
rect 2642 25782 2658 25816
rect 2692 25782 2708 25816
rect 2642 25747 2708 25782
rect 2738 25816 2804 25851
rect 2738 25782 2754 25816
rect 2788 25782 2804 25816
rect 2738 25747 2804 25782
rect 2834 25816 2900 25851
rect 2834 25782 2850 25816
rect 2884 25782 2900 25816
rect 2834 25747 2900 25782
rect 2930 25816 2996 25851
rect 2930 25782 2946 25816
rect 2980 25782 2996 25816
rect 2930 25747 2996 25782
rect 3026 25816 3092 25851
rect 3026 25782 3042 25816
rect 3076 25782 3092 25816
rect 3026 25747 3092 25782
rect 3122 25816 3188 25851
rect 3122 25782 3138 25816
rect 3172 25782 3188 25816
rect 3122 25747 3188 25782
rect 3218 25816 3284 25851
rect 3218 25782 3234 25816
rect 3268 25782 3284 25816
rect 3218 25747 3284 25782
rect 3314 25816 3380 25851
rect 3314 25782 3330 25816
rect 3364 25782 3380 25816
rect 3314 25747 3380 25782
rect 3410 25816 3472 25851
rect 3410 25782 3426 25816
rect 3460 25782 3472 25816
rect 3410 25747 3472 25782
rect 3635 25843 3693 25855
rect 3635 25767 3647 25843
rect 3681 25767 3693 25843
rect 3635 25755 3693 25767
rect 3723 25843 3781 25855
rect 3723 25767 3735 25843
rect 3769 25767 3781 25843
rect 3723 25755 3781 25767
rect 3975 25816 4037 25851
rect 3975 25782 3987 25816
rect 4021 25782 4037 25816
rect 3975 25747 4037 25782
rect 4067 25816 4133 25851
rect 4067 25782 4083 25816
rect 4117 25782 4133 25816
rect 4067 25747 4133 25782
rect 4163 25816 4229 25851
rect 4163 25782 4179 25816
rect 4213 25782 4229 25816
rect 4163 25747 4229 25782
rect 4259 25816 4325 25851
rect 4259 25782 4275 25816
rect 4309 25782 4325 25816
rect 4259 25747 4325 25782
rect 4355 25816 4421 25851
rect 4355 25782 4371 25816
rect 4405 25782 4421 25816
rect 4355 25747 4421 25782
rect 4451 25816 4517 25851
rect 4451 25782 4467 25816
rect 4501 25782 4517 25816
rect 4451 25747 4517 25782
rect 4547 25816 4613 25851
rect 4547 25782 4563 25816
rect 4597 25782 4613 25816
rect 4547 25747 4613 25782
rect 4643 25816 4709 25851
rect 4643 25782 4659 25816
rect 4693 25782 4709 25816
rect 4643 25747 4709 25782
rect 4739 25816 4805 25851
rect 4739 25782 4755 25816
rect 4789 25782 4805 25816
rect 4739 25747 4805 25782
rect 4835 25816 4901 25851
rect 4835 25782 4851 25816
rect 4885 25782 4901 25816
rect 4835 25747 4901 25782
rect 4931 25816 4993 25851
rect 4931 25782 4947 25816
rect 4981 25782 4993 25816
rect 4931 25747 4993 25782
rect 5348 25886 5400 25898
rect 5348 25852 5356 25886
rect 5390 25852 5400 25886
rect 5348 25818 5400 25852
rect 5348 25784 5356 25818
rect 5390 25784 5400 25818
rect 5348 25768 5400 25784
rect 5430 25886 5482 25898
rect 5430 25852 5440 25886
rect 5474 25852 5482 25886
rect 5430 25818 5482 25852
rect 5430 25784 5440 25818
rect 5474 25784 5482 25818
rect 5430 25768 5482 25784
rect 301 24525 363 24560
rect 301 24491 313 24525
rect 347 24491 363 24525
rect 301 24456 363 24491
rect 393 24525 459 24560
rect 393 24491 409 24525
rect 443 24491 459 24525
rect 393 24456 459 24491
rect 489 24525 555 24560
rect 489 24491 505 24525
rect 539 24491 555 24525
rect 489 24456 555 24491
rect 585 24525 651 24560
rect 585 24491 601 24525
rect 635 24491 651 24525
rect 585 24456 651 24491
rect 681 24525 747 24560
rect 681 24491 697 24525
rect 731 24491 747 24525
rect 681 24456 747 24491
rect 777 24525 843 24560
rect 777 24491 793 24525
rect 827 24491 843 24525
rect 777 24456 843 24491
rect 873 24525 939 24560
rect 873 24491 889 24525
rect 923 24491 939 24525
rect 873 24456 939 24491
rect 969 24525 1035 24560
rect 969 24491 985 24525
rect 1019 24491 1035 24525
rect 969 24456 1035 24491
rect 1065 24525 1131 24560
rect 1065 24491 1081 24525
rect 1115 24491 1131 24525
rect 1065 24456 1131 24491
rect 1161 24525 1227 24560
rect 1161 24491 1177 24525
rect 1211 24491 1227 24525
rect 1161 24456 1227 24491
rect 1257 24525 1319 24560
rect 1257 24491 1273 24525
rect 1307 24491 1319 24525
rect 1257 24456 1319 24491
rect 2454 24529 2516 24564
rect 2454 24495 2466 24529
rect 2500 24495 2516 24529
rect 2454 24460 2516 24495
rect 2546 24529 2612 24564
rect 2546 24495 2562 24529
rect 2596 24495 2612 24529
rect 2546 24460 2612 24495
rect 2642 24529 2708 24564
rect 2642 24495 2658 24529
rect 2692 24495 2708 24529
rect 2642 24460 2708 24495
rect 2738 24529 2804 24564
rect 2738 24495 2754 24529
rect 2788 24495 2804 24529
rect 2738 24460 2804 24495
rect 2834 24529 2900 24564
rect 2834 24495 2850 24529
rect 2884 24495 2900 24529
rect 2834 24460 2900 24495
rect 2930 24529 2996 24564
rect 2930 24495 2946 24529
rect 2980 24495 2996 24529
rect 2930 24460 2996 24495
rect 3026 24529 3092 24564
rect 3026 24495 3042 24529
rect 3076 24495 3092 24529
rect 3026 24460 3092 24495
rect 3122 24529 3188 24564
rect 3122 24495 3138 24529
rect 3172 24495 3188 24529
rect 3122 24460 3188 24495
rect 3218 24529 3284 24564
rect 3218 24495 3234 24529
rect 3268 24495 3284 24529
rect 3218 24460 3284 24495
rect 3314 24529 3380 24564
rect 3314 24495 3330 24529
rect 3364 24495 3380 24529
rect 3314 24460 3380 24495
rect 3410 24529 3472 24564
rect 3410 24495 3426 24529
rect 3460 24495 3472 24529
rect 3410 24460 3472 24495
rect 3635 24556 3693 24568
rect 3635 24480 3647 24556
rect 3681 24480 3693 24556
rect 3635 24468 3693 24480
rect 3723 24556 3781 24568
rect 3723 24480 3735 24556
rect 3769 24480 3781 24556
rect 3723 24468 3781 24480
rect 3975 24529 4037 24564
rect 3975 24495 3987 24529
rect 4021 24495 4037 24529
rect 3975 24460 4037 24495
rect 4067 24529 4133 24564
rect 4067 24495 4083 24529
rect 4117 24495 4133 24529
rect 4067 24460 4133 24495
rect 4163 24529 4229 24564
rect 4163 24495 4179 24529
rect 4213 24495 4229 24529
rect 4163 24460 4229 24495
rect 4259 24529 4325 24564
rect 4259 24495 4275 24529
rect 4309 24495 4325 24529
rect 4259 24460 4325 24495
rect 4355 24529 4421 24564
rect 4355 24495 4371 24529
rect 4405 24495 4421 24529
rect 4355 24460 4421 24495
rect 4451 24529 4517 24564
rect 4451 24495 4467 24529
rect 4501 24495 4517 24529
rect 4451 24460 4517 24495
rect 4547 24529 4613 24564
rect 4547 24495 4563 24529
rect 4597 24495 4613 24529
rect 4547 24460 4613 24495
rect 4643 24529 4709 24564
rect 4643 24495 4659 24529
rect 4693 24495 4709 24529
rect 4643 24460 4709 24495
rect 4739 24529 4805 24564
rect 4739 24495 4755 24529
rect 4789 24495 4805 24529
rect 4739 24460 4805 24495
rect 4835 24529 4901 24564
rect 4835 24495 4851 24529
rect 4885 24495 4901 24529
rect 4835 24460 4901 24495
rect 4931 24529 4993 24564
rect 4931 24495 4947 24529
rect 4981 24495 4993 24529
rect 4931 24460 4993 24495
rect 5348 24599 5400 24611
rect 5348 24565 5356 24599
rect 5390 24565 5400 24599
rect 5348 24531 5400 24565
rect 5348 24497 5356 24531
rect 5390 24497 5400 24531
rect 5348 24481 5400 24497
rect 5430 24599 5482 24611
rect 5430 24565 5440 24599
rect 5474 24565 5482 24599
rect 5430 24531 5482 24565
rect 5430 24497 5440 24531
rect 5474 24497 5482 24531
rect 5430 24481 5482 24497
rect 301 23238 363 23273
rect 301 23204 313 23238
rect 347 23204 363 23238
rect 301 23169 363 23204
rect 393 23238 459 23273
rect 393 23204 409 23238
rect 443 23204 459 23238
rect 393 23169 459 23204
rect 489 23238 555 23273
rect 489 23204 505 23238
rect 539 23204 555 23238
rect 489 23169 555 23204
rect 585 23238 651 23273
rect 585 23204 601 23238
rect 635 23204 651 23238
rect 585 23169 651 23204
rect 681 23238 747 23273
rect 681 23204 697 23238
rect 731 23204 747 23238
rect 681 23169 747 23204
rect 777 23238 843 23273
rect 777 23204 793 23238
rect 827 23204 843 23238
rect 777 23169 843 23204
rect 873 23238 939 23273
rect 873 23204 889 23238
rect 923 23204 939 23238
rect 873 23169 939 23204
rect 969 23238 1035 23273
rect 969 23204 985 23238
rect 1019 23204 1035 23238
rect 969 23169 1035 23204
rect 1065 23238 1131 23273
rect 1065 23204 1081 23238
rect 1115 23204 1131 23238
rect 1065 23169 1131 23204
rect 1161 23238 1227 23273
rect 1161 23204 1177 23238
rect 1211 23204 1227 23238
rect 1161 23169 1227 23204
rect 1257 23238 1319 23273
rect 1257 23204 1273 23238
rect 1307 23204 1319 23238
rect 1257 23169 1319 23204
rect 2454 23242 2516 23277
rect 2454 23208 2466 23242
rect 2500 23208 2516 23242
rect 2454 23173 2516 23208
rect 2546 23242 2612 23277
rect 2546 23208 2562 23242
rect 2596 23208 2612 23242
rect 2546 23173 2612 23208
rect 2642 23242 2708 23277
rect 2642 23208 2658 23242
rect 2692 23208 2708 23242
rect 2642 23173 2708 23208
rect 2738 23242 2804 23277
rect 2738 23208 2754 23242
rect 2788 23208 2804 23242
rect 2738 23173 2804 23208
rect 2834 23242 2900 23277
rect 2834 23208 2850 23242
rect 2884 23208 2900 23242
rect 2834 23173 2900 23208
rect 2930 23242 2996 23277
rect 2930 23208 2946 23242
rect 2980 23208 2996 23242
rect 2930 23173 2996 23208
rect 3026 23242 3092 23277
rect 3026 23208 3042 23242
rect 3076 23208 3092 23242
rect 3026 23173 3092 23208
rect 3122 23242 3188 23277
rect 3122 23208 3138 23242
rect 3172 23208 3188 23242
rect 3122 23173 3188 23208
rect 3218 23242 3284 23277
rect 3218 23208 3234 23242
rect 3268 23208 3284 23242
rect 3218 23173 3284 23208
rect 3314 23242 3380 23277
rect 3314 23208 3330 23242
rect 3364 23208 3380 23242
rect 3314 23173 3380 23208
rect 3410 23242 3472 23277
rect 3410 23208 3426 23242
rect 3460 23208 3472 23242
rect 3410 23173 3472 23208
rect 3635 23269 3693 23281
rect 3635 23193 3647 23269
rect 3681 23193 3693 23269
rect 3635 23181 3693 23193
rect 3723 23269 3781 23281
rect 3723 23193 3735 23269
rect 3769 23193 3781 23269
rect 3723 23181 3781 23193
rect 3975 23242 4037 23277
rect 3975 23208 3987 23242
rect 4021 23208 4037 23242
rect 3975 23173 4037 23208
rect 4067 23242 4133 23277
rect 4067 23208 4083 23242
rect 4117 23208 4133 23242
rect 4067 23173 4133 23208
rect 4163 23242 4229 23277
rect 4163 23208 4179 23242
rect 4213 23208 4229 23242
rect 4163 23173 4229 23208
rect 4259 23242 4325 23277
rect 4259 23208 4275 23242
rect 4309 23208 4325 23242
rect 4259 23173 4325 23208
rect 4355 23242 4421 23277
rect 4355 23208 4371 23242
rect 4405 23208 4421 23242
rect 4355 23173 4421 23208
rect 4451 23242 4517 23277
rect 4451 23208 4467 23242
rect 4501 23208 4517 23242
rect 4451 23173 4517 23208
rect 4547 23242 4613 23277
rect 4547 23208 4563 23242
rect 4597 23208 4613 23242
rect 4547 23173 4613 23208
rect 4643 23242 4709 23277
rect 4643 23208 4659 23242
rect 4693 23208 4709 23242
rect 4643 23173 4709 23208
rect 4739 23242 4805 23277
rect 4739 23208 4755 23242
rect 4789 23208 4805 23242
rect 4739 23173 4805 23208
rect 4835 23242 4901 23277
rect 4835 23208 4851 23242
rect 4885 23208 4901 23242
rect 4835 23173 4901 23208
rect 4931 23242 4993 23277
rect 4931 23208 4947 23242
rect 4981 23208 4993 23242
rect 4931 23173 4993 23208
rect 5348 23312 5400 23324
rect 5348 23278 5356 23312
rect 5390 23278 5400 23312
rect 5348 23244 5400 23278
rect 5348 23210 5356 23244
rect 5390 23210 5400 23244
rect 5348 23194 5400 23210
rect 5430 23312 5482 23324
rect 5430 23278 5440 23312
rect 5474 23278 5482 23312
rect 5430 23244 5482 23278
rect 5430 23210 5440 23244
rect 5474 23210 5482 23244
rect 5430 23194 5482 23210
rect 301 21951 363 21986
rect 301 21917 313 21951
rect 347 21917 363 21951
rect 301 21882 363 21917
rect 393 21951 459 21986
rect 393 21917 409 21951
rect 443 21917 459 21951
rect 393 21882 459 21917
rect 489 21951 555 21986
rect 489 21917 505 21951
rect 539 21917 555 21951
rect 489 21882 555 21917
rect 585 21951 651 21986
rect 585 21917 601 21951
rect 635 21917 651 21951
rect 585 21882 651 21917
rect 681 21951 747 21986
rect 681 21917 697 21951
rect 731 21917 747 21951
rect 681 21882 747 21917
rect 777 21951 843 21986
rect 777 21917 793 21951
rect 827 21917 843 21951
rect 777 21882 843 21917
rect 873 21951 939 21986
rect 873 21917 889 21951
rect 923 21917 939 21951
rect 873 21882 939 21917
rect 969 21951 1035 21986
rect 969 21917 985 21951
rect 1019 21917 1035 21951
rect 969 21882 1035 21917
rect 1065 21951 1131 21986
rect 1065 21917 1081 21951
rect 1115 21917 1131 21951
rect 1065 21882 1131 21917
rect 1161 21951 1227 21986
rect 1161 21917 1177 21951
rect 1211 21917 1227 21951
rect 1161 21882 1227 21917
rect 1257 21951 1319 21986
rect 1257 21917 1273 21951
rect 1307 21917 1319 21951
rect 1257 21882 1319 21917
rect 2454 21955 2516 21990
rect 2454 21921 2466 21955
rect 2500 21921 2516 21955
rect 2454 21886 2516 21921
rect 2546 21955 2612 21990
rect 2546 21921 2562 21955
rect 2596 21921 2612 21955
rect 2546 21886 2612 21921
rect 2642 21955 2708 21990
rect 2642 21921 2658 21955
rect 2692 21921 2708 21955
rect 2642 21886 2708 21921
rect 2738 21955 2804 21990
rect 2738 21921 2754 21955
rect 2788 21921 2804 21955
rect 2738 21886 2804 21921
rect 2834 21955 2900 21990
rect 2834 21921 2850 21955
rect 2884 21921 2900 21955
rect 2834 21886 2900 21921
rect 2930 21955 2996 21990
rect 2930 21921 2946 21955
rect 2980 21921 2996 21955
rect 2930 21886 2996 21921
rect 3026 21955 3092 21990
rect 3026 21921 3042 21955
rect 3076 21921 3092 21955
rect 3026 21886 3092 21921
rect 3122 21955 3188 21990
rect 3122 21921 3138 21955
rect 3172 21921 3188 21955
rect 3122 21886 3188 21921
rect 3218 21955 3284 21990
rect 3218 21921 3234 21955
rect 3268 21921 3284 21955
rect 3218 21886 3284 21921
rect 3314 21955 3380 21990
rect 3314 21921 3330 21955
rect 3364 21921 3380 21955
rect 3314 21886 3380 21921
rect 3410 21955 3472 21990
rect 3410 21921 3426 21955
rect 3460 21921 3472 21955
rect 3410 21886 3472 21921
rect 3635 21982 3693 21994
rect 3635 21906 3647 21982
rect 3681 21906 3693 21982
rect 3635 21894 3693 21906
rect 3723 21982 3781 21994
rect 3723 21906 3735 21982
rect 3769 21906 3781 21982
rect 3723 21894 3781 21906
rect 3975 21955 4037 21990
rect 3975 21921 3987 21955
rect 4021 21921 4037 21955
rect 3975 21886 4037 21921
rect 4067 21955 4133 21990
rect 4067 21921 4083 21955
rect 4117 21921 4133 21955
rect 4067 21886 4133 21921
rect 4163 21955 4229 21990
rect 4163 21921 4179 21955
rect 4213 21921 4229 21955
rect 4163 21886 4229 21921
rect 4259 21955 4325 21990
rect 4259 21921 4275 21955
rect 4309 21921 4325 21955
rect 4259 21886 4325 21921
rect 4355 21955 4421 21990
rect 4355 21921 4371 21955
rect 4405 21921 4421 21955
rect 4355 21886 4421 21921
rect 4451 21955 4517 21990
rect 4451 21921 4467 21955
rect 4501 21921 4517 21955
rect 4451 21886 4517 21921
rect 4547 21955 4613 21990
rect 4547 21921 4563 21955
rect 4597 21921 4613 21955
rect 4547 21886 4613 21921
rect 4643 21955 4709 21990
rect 4643 21921 4659 21955
rect 4693 21921 4709 21955
rect 4643 21886 4709 21921
rect 4739 21955 4805 21990
rect 4739 21921 4755 21955
rect 4789 21921 4805 21955
rect 4739 21886 4805 21921
rect 4835 21955 4901 21990
rect 4835 21921 4851 21955
rect 4885 21921 4901 21955
rect 4835 21886 4901 21921
rect 4931 21955 4993 21990
rect 4931 21921 4947 21955
rect 4981 21921 4993 21955
rect 4931 21886 4993 21921
rect 5348 22025 5400 22037
rect 5348 21991 5356 22025
rect 5390 21991 5400 22025
rect 5348 21957 5400 21991
rect 5348 21923 5356 21957
rect 5390 21923 5400 21957
rect 5348 21907 5400 21923
rect 5430 22025 5482 22037
rect 5430 21991 5440 22025
rect 5474 21991 5482 22025
rect 5430 21957 5482 21991
rect 5430 21923 5440 21957
rect 5474 21923 5482 21957
rect 5430 21907 5482 21923
rect 301 20664 363 20699
rect 301 20630 313 20664
rect 347 20630 363 20664
rect 301 20595 363 20630
rect 393 20664 459 20699
rect 393 20630 409 20664
rect 443 20630 459 20664
rect 393 20595 459 20630
rect 489 20664 555 20699
rect 489 20630 505 20664
rect 539 20630 555 20664
rect 489 20595 555 20630
rect 585 20664 651 20699
rect 585 20630 601 20664
rect 635 20630 651 20664
rect 585 20595 651 20630
rect 681 20664 747 20699
rect 681 20630 697 20664
rect 731 20630 747 20664
rect 681 20595 747 20630
rect 777 20664 843 20699
rect 777 20630 793 20664
rect 827 20630 843 20664
rect 777 20595 843 20630
rect 873 20664 939 20699
rect 873 20630 889 20664
rect 923 20630 939 20664
rect 873 20595 939 20630
rect 969 20664 1035 20699
rect 969 20630 985 20664
rect 1019 20630 1035 20664
rect 969 20595 1035 20630
rect 1065 20664 1131 20699
rect 1065 20630 1081 20664
rect 1115 20630 1131 20664
rect 1065 20595 1131 20630
rect 1161 20664 1227 20699
rect 1161 20630 1177 20664
rect 1211 20630 1227 20664
rect 1161 20595 1227 20630
rect 1257 20664 1319 20699
rect 1257 20630 1273 20664
rect 1307 20630 1319 20664
rect 1257 20595 1319 20630
rect 2454 20668 2516 20703
rect 2454 20634 2466 20668
rect 2500 20634 2516 20668
rect 2454 20599 2516 20634
rect 2546 20668 2612 20703
rect 2546 20634 2562 20668
rect 2596 20634 2612 20668
rect 2546 20599 2612 20634
rect 2642 20668 2708 20703
rect 2642 20634 2658 20668
rect 2692 20634 2708 20668
rect 2642 20599 2708 20634
rect 2738 20668 2804 20703
rect 2738 20634 2754 20668
rect 2788 20634 2804 20668
rect 2738 20599 2804 20634
rect 2834 20668 2900 20703
rect 2834 20634 2850 20668
rect 2884 20634 2900 20668
rect 2834 20599 2900 20634
rect 2930 20668 2996 20703
rect 2930 20634 2946 20668
rect 2980 20634 2996 20668
rect 2930 20599 2996 20634
rect 3026 20668 3092 20703
rect 3026 20634 3042 20668
rect 3076 20634 3092 20668
rect 3026 20599 3092 20634
rect 3122 20668 3188 20703
rect 3122 20634 3138 20668
rect 3172 20634 3188 20668
rect 3122 20599 3188 20634
rect 3218 20668 3284 20703
rect 3218 20634 3234 20668
rect 3268 20634 3284 20668
rect 3218 20599 3284 20634
rect 3314 20668 3380 20703
rect 3314 20634 3330 20668
rect 3364 20634 3380 20668
rect 3314 20599 3380 20634
rect 3410 20668 3472 20703
rect 3410 20634 3426 20668
rect 3460 20634 3472 20668
rect 3410 20599 3472 20634
rect 3635 20695 3693 20707
rect 3635 20619 3647 20695
rect 3681 20619 3693 20695
rect 3635 20607 3693 20619
rect 3723 20695 3781 20707
rect 3723 20619 3735 20695
rect 3769 20619 3781 20695
rect 3723 20607 3781 20619
rect 3975 20668 4037 20703
rect 3975 20634 3987 20668
rect 4021 20634 4037 20668
rect 3975 20599 4037 20634
rect 4067 20668 4133 20703
rect 4067 20634 4083 20668
rect 4117 20634 4133 20668
rect 4067 20599 4133 20634
rect 4163 20668 4229 20703
rect 4163 20634 4179 20668
rect 4213 20634 4229 20668
rect 4163 20599 4229 20634
rect 4259 20668 4325 20703
rect 4259 20634 4275 20668
rect 4309 20634 4325 20668
rect 4259 20599 4325 20634
rect 4355 20668 4421 20703
rect 4355 20634 4371 20668
rect 4405 20634 4421 20668
rect 4355 20599 4421 20634
rect 4451 20668 4517 20703
rect 4451 20634 4467 20668
rect 4501 20634 4517 20668
rect 4451 20599 4517 20634
rect 4547 20668 4613 20703
rect 4547 20634 4563 20668
rect 4597 20634 4613 20668
rect 4547 20599 4613 20634
rect 4643 20668 4709 20703
rect 4643 20634 4659 20668
rect 4693 20634 4709 20668
rect 4643 20599 4709 20634
rect 4739 20668 4805 20703
rect 4739 20634 4755 20668
rect 4789 20634 4805 20668
rect 4739 20599 4805 20634
rect 4835 20668 4901 20703
rect 4835 20634 4851 20668
rect 4885 20634 4901 20668
rect 4835 20599 4901 20634
rect 4931 20668 4993 20703
rect 4931 20634 4947 20668
rect 4981 20634 4993 20668
rect 4931 20599 4993 20634
rect 5348 20738 5400 20750
rect 5348 20704 5356 20738
rect 5390 20704 5400 20738
rect 5348 20670 5400 20704
rect 5348 20636 5356 20670
rect 5390 20636 5400 20670
rect 5348 20620 5400 20636
rect 5430 20738 5482 20750
rect 5430 20704 5440 20738
rect 5474 20704 5482 20738
rect 5430 20670 5482 20704
rect 5430 20636 5440 20670
rect 5474 20636 5482 20670
rect 5430 20620 5482 20636
rect 301 19377 363 19412
rect 301 19343 313 19377
rect 347 19343 363 19377
rect 301 19308 363 19343
rect 393 19377 459 19412
rect 393 19343 409 19377
rect 443 19343 459 19377
rect 393 19308 459 19343
rect 489 19377 555 19412
rect 489 19343 505 19377
rect 539 19343 555 19377
rect 489 19308 555 19343
rect 585 19377 651 19412
rect 585 19343 601 19377
rect 635 19343 651 19377
rect 585 19308 651 19343
rect 681 19377 747 19412
rect 681 19343 697 19377
rect 731 19343 747 19377
rect 681 19308 747 19343
rect 777 19377 843 19412
rect 777 19343 793 19377
rect 827 19343 843 19377
rect 777 19308 843 19343
rect 873 19377 939 19412
rect 873 19343 889 19377
rect 923 19343 939 19377
rect 873 19308 939 19343
rect 969 19377 1035 19412
rect 969 19343 985 19377
rect 1019 19343 1035 19377
rect 969 19308 1035 19343
rect 1065 19377 1131 19412
rect 1065 19343 1081 19377
rect 1115 19343 1131 19377
rect 1065 19308 1131 19343
rect 1161 19377 1227 19412
rect 1161 19343 1177 19377
rect 1211 19343 1227 19377
rect 1161 19308 1227 19343
rect 1257 19377 1319 19412
rect 1257 19343 1273 19377
rect 1307 19343 1319 19377
rect 1257 19308 1319 19343
rect 2454 19381 2516 19416
rect 2454 19347 2466 19381
rect 2500 19347 2516 19381
rect 2454 19312 2516 19347
rect 2546 19381 2612 19416
rect 2546 19347 2562 19381
rect 2596 19347 2612 19381
rect 2546 19312 2612 19347
rect 2642 19381 2708 19416
rect 2642 19347 2658 19381
rect 2692 19347 2708 19381
rect 2642 19312 2708 19347
rect 2738 19381 2804 19416
rect 2738 19347 2754 19381
rect 2788 19347 2804 19381
rect 2738 19312 2804 19347
rect 2834 19381 2900 19416
rect 2834 19347 2850 19381
rect 2884 19347 2900 19381
rect 2834 19312 2900 19347
rect 2930 19381 2996 19416
rect 2930 19347 2946 19381
rect 2980 19347 2996 19381
rect 2930 19312 2996 19347
rect 3026 19381 3092 19416
rect 3026 19347 3042 19381
rect 3076 19347 3092 19381
rect 3026 19312 3092 19347
rect 3122 19381 3188 19416
rect 3122 19347 3138 19381
rect 3172 19347 3188 19381
rect 3122 19312 3188 19347
rect 3218 19381 3284 19416
rect 3218 19347 3234 19381
rect 3268 19347 3284 19381
rect 3218 19312 3284 19347
rect 3314 19381 3380 19416
rect 3314 19347 3330 19381
rect 3364 19347 3380 19381
rect 3314 19312 3380 19347
rect 3410 19381 3472 19416
rect 3410 19347 3426 19381
rect 3460 19347 3472 19381
rect 3410 19312 3472 19347
rect 3635 19408 3693 19420
rect 3635 19332 3647 19408
rect 3681 19332 3693 19408
rect 3635 19320 3693 19332
rect 3723 19408 3781 19420
rect 3723 19332 3735 19408
rect 3769 19332 3781 19408
rect 3723 19320 3781 19332
rect 3975 19381 4037 19416
rect 3975 19347 3987 19381
rect 4021 19347 4037 19381
rect 3975 19312 4037 19347
rect 4067 19381 4133 19416
rect 4067 19347 4083 19381
rect 4117 19347 4133 19381
rect 4067 19312 4133 19347
rect 4163 19381 4229 19416
rect 4163 19347 4179 19381
rect 4213 19347 4229 19381
rect 4163 19312 4229 19347
rect 4259 19381 4325 19416
rect 4259 19347 4275 19381
rect 4309 19347 4325 19381
rect 4259 19312 4325 19347
rect 4355 19381 4421 19416
rect 4355 19347 4371 19381
rect 4405 19347 4421 19381
rect 4355 19312 4421 19347
rect 4451 19381 4517 19416
rect 4451 19347 4467 19381
rect 4501 19347 4517 19381
rect 4451 19312 4517 19347
rect 4547 19381 4613 19416
rect 4547 19347 4563 19381
rect 4597 19347 4613 19381
rect 4547 19312 4613 19347
rect 4643 19381 4709 19416
rect 4643 19347 4659 19381
rect 4693 19347 4709 19381
rect 4643 19312 4709 19347
rect 4739 19381 4805 19416
rect 4739 19347 4755 19381
rect 4789 19347 4805 19381
rect 4739 19312 4805 19347
rect 4835 19381 4901 19416
rect 4835 19347 4851 19381
rect 4885 19347 4901 19381
rect 4835 19312 4901 19347
rect 4931 19381 4993 19416
rect 4931 19347 4947 19381
rect 4981 19347 4993 19381
rect 4931 19312 4993 19347
rect 5348 19451 5400 19463
rect 5348 19417 5356 19451
rect 5390 19417 5400 19451
rect 5348 19383 5400 19417
rect 5348 19349 5356 19383
rect 5390 19349 5400 19383
rect 5348 19333 5400 19349
rect 5430 19451 5482 19463
rect 5430 19417 5440 19451
rect 5474 19417 5482 19451
rect 5430 19383 5482 19417
rect 5430 19349 5440 19383
rect 5474 19349 5482 19383
rect 5430 19333 5482 19349
rect 301 18090 363 18125
rect 301 18056 313 18090
rect 347 18056 363 18090
rect 301 18021 363 18056
rect 393 18090 459 18125
rect 393 18056 409 18090
rect 443 18056 459 18090
rect 393 18021 459 18056
rect 489 18090 555 18125
rect 489 18056 505 18090
rect 539 18056 555 18090
rect 489 18021 555 18056
rect 585 18090 651 18125
rect 585 18056 601 18090
rect 635 18056 651 18090
rect 585 18021 651 18056
rect 681 18090 747 18125
rect 681 18056 697 18090
rect 731 18056 747 18090
rect 681 18021 747 18056
rect 777 18090 843 18125
rect 777 18056 793 18090
rect 827 18056 843 18090
rect 777 18021 843 18056
rect 873 18090 939 18125
rect 873 18056 889 18090
rect 923 18056 939 18090
rect 873 18021 939 18056
rect 969 18090 1035 18125
rect 969 18056 985 18090
rect 1019 18056 1035 18090
rect 969 18021 1035 18056
rect 1065 18090 1131 18125
rect 1065 18056 1081 18090
rect 1115 18056 1131 18090
rect 1065 18021 1131 18056
rect 1161 18090 1227 18125
rect 1161 18056 1177 18090
rect 1211 18056 1227 18090
rect 1161 18021 1227 18056
rect 1257 18090 1319 18125
rect 1257 18056 1273 18090
rect 1307 18056 1319 18090
rect 1257 18021 1319 18056
rect 2454 18094 2516 18129
rect 2454 18060 2466 18094
rect 2500 18060 2516 18094
rect 2454 18025 2516 18060
rect 2546 18094 2612 18129
rect 2546 18060 2562 18094
rect 2596 18060 2612 18094
rect 2546 18025 2612 18060
rect 2642 18094 2708 18129
rect 2642 18060 2658 18094
rect 2692 18060 2708 18094
rect 2642 18025 2708 18060
rect 2738 18094 2804 18129
rect 2738 18060 2754 18094
rect 2788 18060 2804 18094
rect 2738 18025 2804 18060
rect 2834 18094 2900 18129
rect 2834 18060 2850 18094
rect 2884 18060 2900 18094
rect 2834 18025 2900 18060
rect 2930 18094 2996 18129
rect 2930 18060 2946 18094
rect 2980 18060 2996 18094
rect 2930 18025 2996 18060
rect 3026 18094 3092 18129
rect 3026 18060 3042 18094
rect 3076 18060 3092 18094
rect 3026 18025 3092 18060
rect 3122 18094 3188 18129
rect 3122 18060 3138 18094
rect 3172 18060 3188 18094
rect 3122 18025 3188 18060
rect 3218 18094 3284 18129
rect 3218 18060 3234 18094
rect 3268 18060 3284 18094
rect 3218 18025 3284 18060
rect 3314 18094 3380 18129
rect 3314 18060 3330 18094
rect 3364 18060 3380 18094
rect 3314 18025 3380 18060
rect 3410 18094 3472 18129
rect 3410 18060 3426 18094
rect 3460 18060 3472 18094
rect 3410 18025 3472 18060
rect 3635 18121 3693 18133
rect 3635 18045 3647 18121
rect 3681 18045 3693 18121
rect 3635 18033 3693 18045
rect 3723 18121 3781 18133
rect 3723 18045 3735 18121
rect 3769 18045 3781 18121
rect 3723 18033 3781 18045
rect 3975 18094 4037 18129
rect 3975 18060 3987 18094
rect 4021 18060 4037 18094
rect 3975 18025 4037 18060
rect 4067 18094 4133 18129
rect 4067 18060 4083 18094
rect 4117 18060 4133 18094
rect 4067 18025 4133 18060
rect 4163 18094 4229 18129
rect 4163 18060 4179 18094
rect 4213 18060 4229 18094
rect 4163 18025 4229 18060
rect 4259 18094 4325 18129
rect 4259 18060 4275 18094
rect 4309 18060 4325 18094
rect 4259 18025 4325 18060
rect 4355 18094 4421 18129
rect 4355 18060 4371 18094
rect 4405 18060 4421 18094
rect 4355 18025 4421 18060
rect 4451 18094 4517 18129
rect 4451 18060 4467 18094
rect 4501 18060 4517 18094
rect 4451 18025 4517 18060
rect 4547 18094 4613 18129
rect 4547 18060 4563 18094
rect 4597 18060 4613 18094
rect 4547 18025 4613 18060
rect 4643 18094 4709 18129
rect 4643 18060 4659 18094
rect 4693 18060 4709 18094
rect 4643 18025 4709 18060
rect 4739 18094 4805 18129
rect 4739 18060 4755 18094
rect 4789 18060 4805 18094
rect 4739 18025 4805 18060
rect 4835 18094 4901 18129
rect 4835 18060 4851 18094
rect 4885 18060 4901 18094
rect 4835 18025 4901 18060
rect 4931 18094 4993 18129
rect 4931 18060 4947 18094
rect 4981 18060 4993 18094
rect 4931 18025 4993 18060
rect 5348 18164 5400 18176
rect 5348 18130 5356 18164
rect 5390 18130 5400 18164
rect 5348 18096 5400 18130
rect 5348 18062 5356 18096
rect 5390 18062 5400 18096
rect 5348 18046 5400 18062
rect 5430 18164 5482 18176
rect 5430 18130 5440 18164
rect 5474 18130 5482 18164
rect 5430 18096 5482 18130
rect 5430 18062 5440 18096
rect 5474 18062 5482 18096
rect 5430 18046 5482 18062
rect 301 16803 363 16838
rect 301 16769 313 16803
rect 347 16769 363 16803
rect 301 16734 363 16769
rect 393 16803 459 16838
rect 393 16769 409 16803
rect 443 16769 459 16803
rect 393 16734 459 16769
rect 489 16803 555 16838
rect 489 16769 505 16803
rect 539 16769 555 16803
rect 489 16734 555 16769
rect 585 16803 651 16838
rect 585 16769 601 16803
rect 635 16769 651 16803
rect 585 16734 651 16769
rect 681 16803 747 16838
rect 681 16769 697 16803
rect 731 16769 747 16803
rect 681 16734 747 16769
rect 777 16803 843 16838
rect 777 16769 793 16803
rect 827 16769 843 16803
rect 777 16734 843 16769
rect 873 16803 939 16838
rect 873 16769 889 16803
rect 923 16769 939 16803
rect 873 16734 939 16769
rect 969 16803 1035 16838
rect 969 16769 985 16803
rect 1019 16769 1035 16803
rect 969 16734 1035 16769
rect 1065 16803 1131 16838
rect 1065 16769 1081 16803
rect 1115 16769 1131 16803
rect 1065 16734 1131 16769
rect 1161 16803 1227 16838
rect 1161 16769 1177 16803
rect 1211 16769 1227 16803
rect 1161 16734 1227 16769
rect 1257 16803 1319 16838
rect 1257 16769 1273 16803
rect 1307 16769 1319 16803
rect 1257 16734 1319 16769
rect 2454 16807 2516 16842
rect 2454 16773 2466 16807
rect 2500 16773 2516 16807
rect 2454 16738 2516 16773
rect 2546 16807 2612 16842
rect 2546 16773 2562 16807
rect 2596 16773 2612 16807
rect 2546 16738 2612 16773
rect 2642 16807 2708 16842
rect 2642 16773 2658 16807
rect 2692 16773 2708 16807
rect 2642 16738 2708 16773
rect 2738 16807 2804 16842
rect 2738 16773 2754 16807
rect 2788 16773 2804 16807
rect 2738 16738 2804 16773
rect 2834 16807 2900 16842
rect 2834 16773 2850 16807
rect 2884 16773 2900 16807
rect 2834 16738 2900 16773
rect 2930 16807 2996 16842
rect 2930 16773 2946 16807
rect 2980 16773 2996 16807
rect 2930 16738 2996 16773
rect 3026 16807 3092 16842
rect 3026 16773 3042 16807
rect 3076 16773 3092 16807
rect 3026 16738 3092 16773
rect 3122 16807 3188 16842
rect 3122 16773 3138 16807
rect 3172 16773 3188 16807
rect 3122 16738 3188 16773
rect 3218 16807 3284 16842
rect 3218 16773 3234 16807
rect 3268 16773 3284 16807
rect 3218 16738 3284 16773
rect 3314 16807 3380 16842
rect 3314 16773 3330 16807
rect 3364 16773 3380 16807
rect 3314 16738 3380 16773
rect 3410 16807 3472 16842
rect 3410 16773 3426 16807
rect 3460 16773 3472 16807
rect 3410 16738 3472 16773
rect 3635 16834 3693 16846
rect 3635 16758 3647 16834
rect 3681 16758 3693 16834
rect 3635 16746 3693 16758
rect 3723 16834 3781 16846
rect 3723 16758 3735 16834
rect 3769 16758 3781 16834
rect 3723 16746 3781 16758
rect 3975 16807 4037 16842
rect 3975 16773 3987 16807
rect 4021 16773 4037 16807
rect 3975 16738 4037 16773
rect 4067 16807 4133 16842
rect 4067 16773 4083 16807
rect 4117 16773 4133 16807
rect 4067 16738 4133 16773
rect 4163 16807 4229 16842
rect 4163 16773 4179 16807
rect 4213 16773 4229 16807
rect 4163 16738 4229 16773
rect 4259 16807 4325 16842
rect 4259 16773 4275 16807
rect 4309 16773 4325 16807
rect 4259 16738 4325 16773
rect 4355 16807 4421 16842
rect 4355 16773 4371 16807
rect 4405 16773 4421 16807
rect 4355 16738 4421 16773
rect 4451 16807 4517 16842
rect 4451 16773 4467 16807
rect 4501 16773 4517 16807
rect 4451 16738 4517 16773
rect 4547 16807 4613 16842
rect 4547 16773 4563 16807
rect 4597 16773 4613 16807
rect 4547 16738 4613 16773
rect 4643 16807 4709 16842
rect 4643 16773 4659 16807
rect 4693 16773 4709 16807
rect 4643 16738 4709 16773
rect 4739 16807 4805 16842
rect 4739 16773 4755 16807
rect 4789 16773 4805 16807
rect 4739 16738 4805 16773
rect 4835 16807 4901 16842
rect 4835 16773 4851 16807
rect 4885 16773 4901 16807
rect 4835 16738 4901 16773
rect 4931 16807 4993 16842
rect 4931 16773 4947 16807
rect 4981 16773 4993 16807
rect 4931 16738 4993 16773
rect 5348 16877 5400 16889
rect 5348 16843 5356 16877
rect 5390 16843 5400 16877
rect 5348 16809 5400 16843
rect 5348 16775 5356 16809
rect 5390 16775 5400 16809
rect 5348 16759 5400 16775
rect 5430 16877 5482 16889
rect 5430 16843 5440 16877
rect 5474 16843 5482 16877
rect 5430 16809 5482 16843
rect 5430 16775 5440 16809
rect 5474 16775 5482 16809
rect 5430 16759 5482 16775
rect 301 15516 363 15551
rect 301 15482 313 15516
rect 347 15482 363 15516
rect 301 15447 363 15482
rect 393 15516 459 15551
rect 393 15482 409 15516
rect 443 15482 459 15516
rect 393 15447 459 15482
rect 489 15516 555 15551
rect 489 15482 505 15516
rect 539 15482 555 15516
rect 489 15447 555 15482
rect 585 15516 651 15551
rect 585 15482 601 15516
rect 635 15482 651 15516
rect 585 15447 651 15482
rect 681 15516 747 15551
rect 681 15482 697 15516
rect 731 15482 747 15516
rect 681 15447 747 15482
rect 777 15516 843 15551
rect 777 15482 793 15516
rect 827 15482 843 15516
rect 777 15447 843 15482
rect 873 15516 939 15551
rect 873 15482 889 15516
rect 923 15482 939 15516
rect 873 15447 939 15482
rect 969 15516 1035 15551
rect 969 15482 985 15516
rect 1019 15482 1035 15516
rect 969 15447 1035 15482
rect 1065 15516 1131 15551
rect 1065 15482 1081 15516
rect 1115 15482 1131 15516
rect 1065 15447 1131 15482
rect 1161 15516 1227 15551
rect 1161 15482 1177 15516
rect 1211 15482 1227 15516
rect 1161 15447 1227 15482
rect 1257 15516 1319 15551
rect 1257 15482 1273 15516
rect 1307 15482 1319 15516
rect 1257 15447 1319 15482
rect 2454 15520 2516 15555
rect 2454 15486 2466 15520
rect 2500 15486 2516 15520
rect 2454 15451 2516 15486
rect 2546 15520 2612 15555
rect 2546 15486 2562 15520
rect 2596 15486 2612 15520
rect 2546 15451 2612 15486
rect 2642 15520 2708 15555
rect 2642 15486 2658 15520
rect 2692 15486 2708 15520
rect 2642 15451 2708 15486
rect 2738 15520 2804 15555
rect 2738 15486 2754 15520
rect 2788 15486 2804 15520
rect 2738 15451 2804 15486
rect 2834 15520 2900 15555
rect 2834 15486 2850 15520
rect 2884 15486 2900 15520
rect 2834 15451 2900 15486
rect 2930 15520 2996 15555
rect 2930 15486 2946 15520
rect 2980 15486 2996 15520
rect 2930 15451 2996 15486
rect 3026 15520 3092 15555
rect 3026 15486 3042 15520
rect 3076 15486 3092 15520
rect 3026 15451 3092 15486
rect 3122 15520 3188 15555
rect 3122 15486 3138 15520
rect 3172 15486 3188 15520
rect 3122 15451 3188 15486
rect 3218 15520 3284 15555
rect 3218 15486 3234 15520
rect 3268 15486 3284 15520
rect 3218 15451 3284 15486
rect 3314 15520 3380 15555
rect 3314 15486 3330 15520
rect 3364 15486 3380 15520
rect 3314 15451 3380 15486
rect 3410 15520 3472 15555
rect 3410 15486 3426 15520
rect 3460 15486 3472 15520
rect 3410 15451 3472 15486
rect 3635 15547 3693 15559
rect 3635 15471 3647 15547
rect 3681 15471 3693 15547
rect 3635 15459 3693 15471
rect 3723 15547 3781 15559
rect 3723 15471 3735 15547
rect 3769 15471 3781 15547
rect 3723 15459 3781 15471
rect 3975 15520 4037 15555
rect 3975 15486 3987 15520
rect 4021 15486 4037 15520
rect 3975 15451 4037 15486
rect 4067 15520 4133 15555
rect 4067 15486 4083 15520
rect 4117 15486 4133 15520
rect 4067 15451 4133 15486
rect 4163 15520 4229 15555
rect 4163 15486 4179 15520
rect 4213 15486 4229 15520
rect 4163 15451 4229 15486
rect 4259 15520 4325 15555
rect 4259 15486 4275 15520
rect 4309 15486 4325 15520
rect 4259 15451 4325 15486
rect 4355 15520 4421 15555
rect 4355 15486 4371 15520
rect 4405 15486 4421 15520
rect 4355 15451 4421 15486
rect 4451 15520 4517 15555
rect 4451 15486 4467 15520
rect 4501 15486 4517 15520
rect 4451 15451 4517 15486
rect 4547 15520 4613 15555
rect 4547 15486 4563 15520
rect 4597 15486 4613 15520
rect 4547 15451 4613 15486
rect 4643 15520 4709 15555
rect 4643 15486 4659 15520
rect 4693 15486 4709 15520
rect 4643 15451 4709 15486
rect 4739 15520 4805 15555
rect 4739 15486 4755 15520
rect 4789 15486 4805 15520
rect 4739 15451 4805 15486
rect 4835 15520 4901 15555
rect 4835 15486 4851 15520
rect 4885 15486 4901 15520
rect 4835 15451 4901 15486
rect 4931 15520 4993 15555
rect 4931 15486 4947 15520
rect 4981 15486 4993 15520
rect 4931 15451 4993 15486
rect 5348 15590 5400 15602
rect 5348 15556 5356 15590
rect 5390 15556 5400 15590
rect 5348 15522 5400 15556
rect 5348 15488 5356 15522
rect 5390 15488 5400 15522
rect 5348 15472 5400 15488
rect 5430 15590 5482 15602
rect 5430 15556 5440 15590
rect 5474 15556 5482 15590
rect 5430 15522 5482 15556
rect 5430 15488 5440 15522
rect 5474 15488 5482 15522
rect 5430 15472 5482 15488
rect 301 14229 363 14264
rect 301 14195 313 14229
rect 347 14195 363 14229
rect 301 14160 363 14195
rect 393 14229 459 14264
rect 393 14195 409 14229
rect 443 14195 459 14229
rect 393 14160 459 14195
rect 489 14229 555 14264
rect 489 14195 505 14229
rect 539 14195 555 14229
rect 489 14160 555 14195
rect 585 14229 651 14264
rect 585 14195 601 14229
rect 635 14195 651 14229
rect 585 14160 651 14195
rect 681 14229 747 14264
rect 681 14195 697 14229
rect 731 14195 747 14229
rect 681 14160 747 14195
rect 777 14229 843 14264
rect 777 14195 793 14229
rect 827 14195 843 14229
rect 777 14160 843 14195
rect 873 14229 939 14264
rect 873 14195 889 14229
rect 923 14195 939 14229
rect 873 14160 939 14195
rect 969 14229 1035 14264
rect 969 14195 985 14229
rect 1019 14195 1035 14229
rect 969 14160 1035 14195
rect 1065 14229 1131 14264
rect 1065 14195 1081 14229
rect 1115 14195 1131 14229
rect 1065 14160 1131 14195
rect 1161 14229 1227 14264
rect 1161 14195 1177 14229
rect 1211 14195 1227 14229
rect 1161 14160 1227 14195
rect 1257 14229 1319 14264
rect 1257 14195 1273 14229
rect 1307 14195 1319 14229
rect 1257 14160 1319 14195
rect 2454 14233 2516 14268
rect 2454 14199 2466 14233
rect 2500 14199 2516 14233
rect 2454 14164 2516 14199
rect 2546 14233 2612 14268
rect 2546 14199 2562 14233
rect 2596 14199 2612 14233
rect 2546 14164 2612 14199
rect 2642 14233 2708 14268
rect 2642 14199 2658 14233
rect 2692 14199 2708 14233
rect 2642 14164 2708 14199
rect 2738 14233 2804 14268
rect 2738 14199 2754 14233
rect 2788 14199 2804 14233
rect 2738 14164 2804 14199
rect 2834 14233 2900 14268
rect 2834 14199 2850 14233
rect 2884 14199 2900 14233
rect 2834 14164 2900 14199
rect 2930 14233 2996 14268
rect 2930 14199 2946 14233
rect 2980 14199 2996 14233
rect 2930 14164 2996 14199
rect 3026 14233 3092 14268
rect 3026 14199 3042 14233
rect 3076 14199 3092 14233
rect 3026 14164 3092 14199
rect 3122 14233 3188 14268
rect 3122 14199 3138 14233
rect 3172 14199 3188 14233
rect 3122 14164 3188 14199
rect 3218 14233 3284 14268
rect 3218 14199 3234 14233
rect 3268 14199 3284 14233
rect 3218 14164 3284 14199
rect 3314 14233 3380 14268
rect 3314 14199 3330 14233
rect 3364 14199 3380 14233
rect 3314 14164 3380 14199
rect 3410 14233 3472 14268
rect 3410 14199 3426 14233
rect 3460 14199 3472 14233
rect 3410 14164 3472 14199
rect 3635 14260 3693 14272
rect 3635 14184 3647 14260
rect 3681 14184 3693 14260
rect 3635 14172 3693 14184
rect 3723 14260 3781 14272
rect 3723 14184 3735 14260
rect 3769 14184 3781 14260
rect 3723 14172 3781 14184
rect 3975 14233 4037 14268
rect 3975 14199 3987 14233
rect 4021 14199 4037 14233
rect 3975 14164 4037 14199
rect 4067 14233 4133 14268
rect 4067 14199 4083 14233
rect 4117 14199 4133 14233
rect 4067 14164 4133 14199
rect 4163 14233 4229 14268
rect 4163 14199 4179 14233
rect 4213 14199 4229 14233
rect 4163 14164 4229 14199
rect 4259 14233 4325 14268
rect 4259 14199 4275 14233
rect 4309 14199 4325 14233
rect 4259 14164 4325 14199
rect 4355 14233 4421 14268
rect 4355 14199 4371 14233
rect 4405 14199 4421 14233
rect 4355 14164 4421 14199
rect 4451 14233 4517 14268
rect 4451 14199 4467 14233
rect 4501 14199 4517 14233
rect 4451 14164 4517 14199
rect 4547 14233 4613 14268
rect 4547 14199 4563 14233
rect 4597 14199 4613 14233
rect 4547 14164 4613 14199
rect 4643 14233 4709 14268
rect 4643 14199 4659 14233
rect 4693 14199 4709 14233
rect 4643 14164 4709 14199
rect 4739 14233 4805 14268
rect 4739 14199 4755 14233
rect 4789 14199 4805 14233
rect 4739 14164 4805 14199
rect 4835 14233 4901 14268
rect 4835 14199 4851 14233
rect 4885 14199 4901 14233
rect 4835 14164 4901 14199
rect 4931 14233 4993 14268
rect 4931 14199 4947 14233
rect 4981 14199 4993 14233
rect 4931 14164 4993 14199
rect 5348 14303 5400 14315
rect 5348 14269 5356 14303
rect 5390 14269 5400 14303
rect 5348 14235 5400 14269
rect 5348 14201 5356 14235
rect 5390 14201 5400 14235
rect 5348 14185 5400 14201
rect 5430 14303 5482 14315
rect 5430 14269 5440 14303
rect 5474 14269 5482 14303
rect 5430 14235 5482 14269
rect 5430 14201 5440 14235
rect 5474 14201 5482 14235
rect 5430 14185 5482 14201
rect 301 12942 363 12977
rect 301 12908 313 12942
rect 347 12908 363 12942
rect 301 12873 363 12908
rect 393 12942 459 12977
rect 393 12908 409 12942
rect 443 12908 459 12942
rect 393 12873 459 12908
rect 489 12942 555 12977
rect 489 12908 505 12942
rect 539 12908 555 12942
rect 489 12873 555 12908
rect 585 12942 651 12977
rect 585 12908 601 12942
rect 635 12908 651 12942
rect 585 12873 651 12908
rect 681 12942 747 12977
rect 681 12908 697 12942
rect 731 12908 747 12942
rect 681 12873 747 12908
rect 777 12942 843 12977
rect 777 12908 793 12942
rect 827 12908 843 12942
rect 777 12873 843 12908
rect 873 12942 939 12977
rect 873 12908 889 12942
rect 923 12908 939 12942
rect 873 12873 939 12908
rect 969 12942 1035 12977
rect 969 12908 985 12942
rect 1019 12908 1035 12942
rect 969 12873 1035 12908
rect 1065 12942 1131 12977
rect 1065 12908 1081 12942
rect 1115 12908 1131 12942
rect 1065 12873 1131 12908
rect 1161 12942 1227 12977
rect 1161 12908 1177 12942
rect 1211 12908 1227 12942
rect 1161 12873 1227 12908
rect 1257 12942 1319 12977
rect 1257 12908 1273 12942
rect 1307 12908 1319 12942
rect 1257 12873 1319 12908
rect 2454 12946 2516 12981
rect 2454 12912 2466 12946
rect 2500 12912 2516 12946
rect 2454 12877 2516 12912
rect 2546 12946 2612 12981
rect 2546 12912 2562 12946
rect 2596 12912 2612 12946
rect 2546 12877 2612 12912
rect 2642 12946 2708 12981
rect 2642 12912 2658 12946
rect 2692 12912 2708 12946
rect 2642 12877 2708 12912
rect 2738 12946 2804 12981
rect 2738 12912 2754 12946
rect 2788 12912 2804 12946
rect 2738 12877 2804 12912
rect 2834 12946 2900 12981
rect 2834 12912 2850 12946
rect 2884 12912 2900 12946
rect 2834 12877 2900 12912
rect 2930 12946 2996 12981
rect 2930 12912 2946 12946
rect 2980 12912 2996 12946
rect 2930 12877 2996 12912
rect 3026 12946 3092 12981
rect 3026 12912 3042 12946
rect 3076 12912 3092 12946
rect 3026 12877 3092 12912
rect 3122 12946 3188 12981
rect 3122 12912 3138 12946
rect 3172 12912 3188 12946
rect 3122 12877 3188 12912
rect 3218 12946 3284 12981
rect 3218 12912 3234 12946
rect 3268 12912 3284 12946
rect 3218 12877 3284 12912
rect 3314 12946 3380 12981
rect 3314 12912 3330 12946
rect 3364 12912 3380 12946
rect 3314 12877 3380 12912
rect 3410 12946 3472 12981
rect 3410 12912 3426 12946
rect 3460 12912 3472 12946
rect 3410 12877 3472 12912
rect 3635 12973 3693 12985
rect 3635 12897 3647 12973
rect 3681 12897 3693 12973
rect 3635 12885 3693 12897
rect 3723 12973 3781 12985
rect 3723 12897 3735 12973
rect 3769 12897 3781 12973
rect 3723 12885 3781 12897
rect 3975 12946 4037 12981
rect 3975 12912 3987 12946
rect 4021 12912 4037 12946
rect 3975 12877 4037 12912
rect 4067 12946 4133 12981
rect 4067 12912 4083 12946
rect 4117 12912 4133 12946
rect 4067 12877 4133 12912
rect 4163 12946 4229 12981
rect 4163 12912 4179 12946
rect 4213 12912 4229 12946
rect 4163 12877 4229 12912
rect 4259 12946 4325 12981
rect 4259 12912 4275 12946
rect 4309 12912 4325 12946
rect 4259 12877 4325 12912
rect 4355 12946 4421 12981
rect 4355 12912 4371 12946
rect 4405 12912 4421 12946
rect 4355 12877 4421 12912
rect 4451 12946 4517 12981
rect 4451 12912 4467 12946
rect 4501 12912 4517 12946
rect 4451 12877 4517 12912
rect 4547 12946 4613 12981
rect 4547 12912 4563 12946
rect 4597 12912 4613 12946
rect 4547 12877 4613 12912
rect 4643 12946 4709 12981
rect 4643 12912 4659 12946
rect 4693 12912 4709 12946
rect 4643 12877 4709 12912
rect 4739 12946 4805 12981
rect 4739 12912 4755 12946
rect 4789 12912 4805 12946
rect 4739 12877 4805 12912
rect 4835 12946 4901 12981
rect 4835 12912 4851 12946
rect 4885 12912 4901 12946
rect 4835 12877 4901 12912
rect 4931 12946 4993 12981
rect 4931 12912 4947 12946
rect 4981 12912 4993 12946
rect 4931 12877 4993 12912
rect 5348 13016 5400 13028
rect 5348 12982 5356 13016
rect 5390 12982 5400 13016
rect 5348 12948 5400 12982
rect 5348 12914 5356 12948
rect 5390 12914 5400 12948
rect 5348 12898 5400 12914
rect 5430 13016 5482 13028
rect 5430 12982 5440 13016
rect 5474 12982 5482 13016
rect 5430 12948 5482 12982
rect 5430 12914 5440 12948
rect 5474 12914 5482 12948
rect 5430 12898 5482 12914
rect 301 11655 363 11690
rect 301 11621 313 11655
rect 347 11621 363 11655
rect 301 11586 363 11621
rect 393 11655 459 11690
rect 393 11621 409 11655
rect 443 11621 459 11655
rect 393 11586 459 11621
rect 489 11655 555 11690
rect 489 11621 505 11655
rect 539 11621 555 11655
rect 489 11586 555 11621
rect 585 11655 651 11690
rect 585 11621 601 11655
rect 635 11621 651 11655
rect 585 11586 651 11621
rect 681 11655 747 11690
rect 681 11621 697 11655
rect 731 11621 747 11655
rect 681 11586 747 11621
rect 777 11655 843 11690
rect 777 11621 793 11655
rect 827 11621 843 11655
rect 777 11586 843 11621
rect 873 11655 939 11690
rect 873 11621 889 11655
rect 923 11621 939 11655
rect 873 11586 939 11621
rect 969 11655 1035 11690
rect 969 11621 985 11655
rect 1019 11621 1035 11655
rect 969 11586 1035 11621
rect 1065 11655 1131 11690
rect 1065 11621 1081 11655
rect 1115 11621 1131 11655
rect 1065 11586 1131 11621
rect 1161 11655 1227 11690
rect 1161 11621 1177 11655
rect 1211 11621 1227 11655
rect 1161 11586 1227 11621
rect 1257 11655 1319 11690
rect 1257 11621 1273 11655
rect 1307 11621 1319 11655
rect 1257 11586 1319 11621
rect 2454 11659 2516 11694
rect 2454 11625 2466 11659
rect 2500 11625 2516 11659
rect 2454 11590 2516 11625
rect 2546 11659 2612 11694
rect 2546 11625 2562 11659
rect 2596 11625 2612 11659
rect 2546 11590 2612 11625
rect 2642 11659 2708 11694
rect 2642 11625 2658 11659
rect 2692 11625 2708 11659
rect 2642 11590 2708 11625
rect 2738 11659 2804 11694
rect 2738 11625 2754 11659
rect 2788 11625 2804 11659
rect 2738 11590 2804 11625
rect 2834 11659 2900 11694
rect 2834 11625 2850 11659
rect 2884 11625 2900 11659
rect 2834 11590 2900 11625
rect 2930 11659 2996 11694
rect 2930 11625 2946 11659
rect 2980 11625 2996 11659
rect 2930 11590 2996 11625
rect 3026 11659 3092 11694
rect 3026 11625 3042 11659
rect 3076 11625 3092 11659
rect 3026 11590 3092 11625
rect 3122 11659 3188 11694
rect 3122 11625 3138 11659
rect 3172 11625 3188 11659
rect 3122 11590 3188 11625
rect 3218 11659 3284 11694
rect 3218 11625 3234 11659
rect 3268 11625 3284 11659
rect 3218 11590 3284 11625
rect 3314 11659 3380 11694
rect 3314 11625 3330 11659
rect 3364 11625 3380 11659
rect 3314 11590 3380 11625
rect 3410 11659 3472 11694
rect 3410 11625 3426 11659
rect 3460 11625 3472 11659
rect 3410 11590 3472 11625
rect 3635 11686 3693 11698
rect 3635 11610 3647 11686
rect 3681 11610 3693 11686
rect 3635 11598 3693 11610
rect 3723 11686 3781 11698
rect 3723 11610 3735 11686
rect 3769 11610 3781 11686
rect 3723 11598 3781 11610
rect 3975 11659 4037 11694
rect 3975 11625 3987 11659
rect 4021 11625 4037 11659
rect 3975 11590 4037 11625
rect 4067 11659 4133 11694
rect 4067 11625 4083 11659
rect 4117 11625 4133 11659
rect 4067 11590 4133 11625
rect 4163 11659 4229 11694
rect 4163 11625 4179 11659
rect 4213 11625 4229 11659
rect 4163 11590 4229 11625
rect 4259 11659 4325 11694
rect 4259 11625 4275 11659
rect 4309 11625 4325 11659
rect 4259 11590 4325 11625
rect 4355 11659 4421 11694
rect 4355 11625 4371 11659
rect 4405 11625 4421 11659
rect 4355 11590 4421 11625
rect 4451 11659 4517 11694
rect 4451 11625 4467 11659
rect 4501 11625 4517 11659
rect 4451 11590 4517 11625
rect 4547 11659 4613 11694
rect 4547 11625 4563 11659
rect 4597 11625 4613 11659
rect 4547 11590 4613 11625
rect 4643 11659 4709 11694
rect 4643 11625 4659 11659
rect 4693 11625 4709 11659
rect 4643 11590 4709 11625
rect 4739 11659 4805 11694
rect 4739 11625 4755 11659
rect 4789 11625 4805 11659
rect 4739 11590 4805 11625
rect 4835 11659 4901 11694
rect 4835 11625 4851 11659
rect 4885 11625 4901 11659
rect 4835 11590 4901 11625
rect 4931 11659 4993 11694
rect 4931 11625 4947 11659
rect 4981 11625 4993 11659
rect 4931 11590 4993 11625
rect 5348 11729 5400 11741
rect 5348 11695 5356 11729
rect 5390 11695 5400 11729
rect 5348 11661 5400 11695
rect 5348 11627 5356 11661
rect 5390 11627 5400 11661
rect 5348 11611 5400 11627
rect 5430 11729 5482 11741
rect 5430 11695 5440 11729
rect 5474 11695 5482 11729
rect 5430 11661 5482 11695
rect 5430 11627 5440 11661
rect 5474 11627 5482 11661
rect 5430 11611 5482 11627
rect 301 10368 363 10403
rect 301 10334 313 10368
rect 347 10334 363 10368
rect 301 10299 363 10334
rect 393 10368 459 10403
rect 393 10334 409 10368
rect 443 10334 459 10368
rect 393 10299 459 10334
rect 489 10368 555 10403
rect 489 10334 505 10368
rect 539 10334 555 10368
rect 489 10299 555 10334
rect 585 10368 651 10403
rect 585 10334 601 10368
rect 635 10334 651 10368
rect 585 10299 651 10334
rect 681 10368 747 10403
rect 681 10334 697 10368
rect 731 10334 747 10368
rect 681 10299 747 10334
rect 777 10368 843 10403
rect 777 10334 793 10368
rect 827 10334 843 10368
rect 777 10299 843 10334
rect 873 10368 939 10403
rect 873 10334 889 10368
rect 923 10334 939 10368
rect 873 10299 939 10334
rect 969 10368 1035 10403
rect 969 10334 985 10368
rect 1019 10334 1035 10368
rect 969 10299 1035 10334
rect 1065 10368 1131 10403
rect 1065 10334 1081 10368
rect 1115 10334 1131 10368
rect 1065 10299 1131 10334
rect 1161 10368 1227 10403
rect 1161 10334 1177 10368
rect 1211 10334 1227 10368
rect 1161 10299 1227 10334
rect 1257 10368 1319 10403
rect 1257 10334 1273 10368
rect 1307 10334 1319 10368
rect 1257 10299 1319 10334
rect 2454 10372 2516 10407
rect 2454 10338 2466 10372
rect 2500 10338 2516 10372
rect 2454 10303 2516 10338
rect 2546 10372 2612 10407
rect 2546 10338 2562 10372
rect 2596 10338 2612 10372
rect 2546 10303 2612 10338
rect 2642 10372 2708 10407
rect 2642 10338 2658 10372
rect 2692 10338 2708 10372
rect 2642 10303 2708 10338
rect 2738 10372 2804 10407
rect 2738 10338 2754 10372
rect 2788 10338 2804 10372
rect 2738 10303 2804 10338
rect 2834 10372 2900 10407
rect 2834 10338 2850 10372
rect 2884 10338 2900 10372
rect 2834 10303 2900 10338
rect 2930 10372 2996 10407
rect 2930 10338 2946 10372
rect 2980 10338 2996 10372
rect 2930 10303 2996 10338
rect 3026 10372 3092 10407
rect 3026 10338 3042 10372
rect 3076 10338 3092 10372
rect 3026 10303 3092 10338
rect 3122 10372 3188 10407
rect 3122 10338 3138 10372
rect 3172 10338 3188 10372
rect 3122 10303 3188 10338
rect 3218 10372 3284 10407
rect 3218 10338 3234 10372
rect 3268 10338 3284 10372
rect 3218 10303 3284 10338
rect 3314 10372 3380 10407
rect 3314 10338 3330 10372
rect 3364 10338 3380 10372
rect 3314 10303 3380 10338
rect 3410 10372 3472 10407
rect 3410 10338 3426 10372
rect 3460 10338 3472 10372
rect 3410 10303 3472 10338
rect 3635 10399 3693 10411
rect 3635 10323 3647 10399
rect 3681 10323 3693 10399
rect 3635 10311 3693 10323
rect 3723 10399 3781 10411
rect 3723 10323 3735 10399
rect 3769 10323 3781 10399
rect 3723 10311 3781 10323
rect 3975 10372 4037 10407
rect 3975 10338 3987 10372
rect 4021 10338 4037 10372
rect 3975 10303 4037 10338
rect 4067 10372 4133 10407
rect 4067 10338 4083 10372
rect 4117 10338 4133 10372
rect 4067 10303 4133 10338
rect 4163 10372 4229 10407
rect 4163 10338 4179 10372
rect 4213 10338 4229 10372
rect 4163 10303 4229 10338
rect 4259 10372 4325 10407
rect 4259 10338 4275 10372
rect 4309 10338 4325 10372
rect 4259 10303 4325 10338
rect 4355 10372 4421 10407
rect 4355 10338 4371 10372
rect 4405 10338 4421 10372
rect 4355 10303 4421 10338
rect 4451 10372 4517 10407
rect 4451 10338 4467 10372
rect 4501 10338 4517 10372
rect 4451 10303 4517 10338
rect 4547 10372 4613 10407
rect 4547 10338 4563 10372
rect 4597 10338 4613 10372
rect 4547 10303 4613 10338
rect 4643 10372 4709 10407
rect 4643 10338 4659 10372
rect 4693 10338 4709 10372
rect 4643 10303 4709 10338
rect 4739 10372 4805 10407
rect 4739 10338 4755 10372
rect 4789 10338 4805 10372
rect 4739 10303 4805 10338
rect 4835 10372 4901 10407
rect 4835 10338 4851 10372
rect 4885 10338 4901 10372
rect 4835 10303 4901 10338
rect 4931 10372 4993 10407
rect 4931 10338 4947 10372
rect 4981 10338 4993 10372
rect 4931 10303 4993 10338
rect 5348 10442 5400 10454
rect 5348 10408 5356 10442
rect 5390 10408 5400 10442
rect 5348 10374 5400 10408
rect 5348 10340 5356 10374
rect 5390 10340 5400 10374
rect 5348 10324 5400 10340
rect 5430 10442 5482 10454
rect 5430 10408 5440 10442
rect 5474 10408 5482 10442
rect 5430 10374 5482 10408
rect 5430 10340 5440 10374
rect 5474 10340 5482 10374
rect 5430 10324 5482 10340
rect 301 9081 363 9116
rect 301 9047 313 9081
rect 347 9047 363 9081
rect 301 9012 363 9047
rect 393 9081 459 9116
rect 393 9047 409 9081
rect 443 9047 459 9081
rect 393 9012 459 9047
rect 489 9081 555 9116
rect 489 9047 505 9081
rect 539 9047 555 9081
rect 489 9012 555 9047
rect 585 9081 651 9116
rect 585 9047 601 9081
rect 635 9047 651 9081
rect 585 9012 651 9047
rect 681 9081 747 9116
rect 681 9047 697 9081
rect 731 9047 747 9081
rect 681 9012 747 9047
rect 777 9081 843 9116
rect 777 9047 793 9081
rect 827 9047 843 9081
rect 777 9012 843 9047
rect 873 9081 939 9116
rect 873 9047 889 9081
rect 923 9047 939 9081
rect 873 9012 939 9047
rect 969 9081 1035 9116
rect 969 9047 985 9081
rect 1019 9047 1035 9081
rect 969 9012 1035 9047
rect 1065 9081 1131 9116
rect 1065 9047 1081 9081
rect 1115 9047 1131 9081
rect 1065 9012 1131 9047
rect 1161 9081 1227 9116
rect 1161 9047 1177 9081
rect 1211 9047 1227 9081
rect 1161 9012 1227 9047
rect 1257 9081 1319 9116
rect 1257 9047 1273 9081
rect 1307 9047 1319 9081
rect 1257 9012 1319 9047
rect 2454 9085 2516 9120
rect 2454 9051 2466 9085
rect 2500 9051 2516 9085
rect 2454 9016 2516 9051
rect 2546 9085 2612 9120
rect 2546 9051 2562 9085
rect 2596 9051 2612 9085
rect 2546 9016 2612 9051
rect 2642 9085 2708 9120
rect 2642 9051 2658 9085
rect 2692 9051 2708 9085
rect 2642 9016 2708 9051
rect 2738 9085 2804 9120
rect 2738 9051 2754 9085
rect 2788 9051 2804 9085
rect 2738 9016 2804 9051
rect 2834 9085 2900 9120
rect 2834 9051 2850 9085
rect 2884 9051 2900 9085
rect 2834 9016 2900 9051
rect 2930 9085 2996 9120
rect 2930 9051 2946 9085
rect 2980 9051 2996 9085
rect 2930 9016 2996 9051
rect 3026 9085 3092 9120
rect 3026 9051 3042 9085
rect 3076 9051 3092 9085
rect 3026 9016 3092 9051
rect 3122 9085 3188 9120
rect 3122 9051 3138 9085
rect 3172 9051 3188 9085
rect 3122 9016 3188 9051
rect 3218 9085 3284 9120
rect 3218 9051 3234 9085
rect 3268 9051 3284 9085
rect 3218 9016 3284 9051
rect 3314 9085 3380 9120
rect 3314 9051 3330 9085
rect 3364 9051 3380 9085
rect 3314 9016 3380 9051
rect 3410 9085 3472 9120
rect 3410 9051 3426 9085
rect 3460 9051 3472 9085
rect 3410 9016 3472 9051
rect 3635 9112 3693 9124
rect 3635 9036 3647 9112
rect 3681 9036 3693 9112
rect 3635 9024 3693 9036
rect 3723 9112 3781 9124
rect 3723 9036 3735 9112
rect 3769 9036 3781 9112
rect 3723 9024 3781 9036
rect 3975 9085 4037 9120
rect 3975 9051 3987 9085
rect 4021 9051 4037 9085
rect 3975 9016 4037 9051
rect 4067 9085 4133 9120
rect 4067 9051 4083 9085
rect 4117 9051 4133 9085
rect 4067 9016 4133 9051
rect 4163 9085 4229 9120
rect 4163 9051 4179 9085
rect 4213 9051 4229 9085
rect 4163 9016 4229 9051
rect 4259 9085 4325 9120
rect 4259 9051 4275 9085
rect 4309 9051 4325 9085
rect 4259 9016 4325 9051
rect 4355 9085 4421 9120
rect 4355 9051 4371 9085
rect 4405 9051 4421 9085
rect 4355 9016 4421 9051
rect 4451 9085 4517 9120
rect 4451 9051 4467 9085
rect 4501 9051 4517 9085
rect 4451 9016 4517 9051
rect 4547 9085 4613 9120
rect 4547 9051 4563 9085
rect 4597 9051 4613 9085
rect 4547 9016 4613 9051
rect 4643 9085 4709 9120
rect 4643 9051 4659 9085
rect 4693 9051 4709 9085
rect 4643 9016 4709 9051
rect 4739 9085 4805 9120
rect 4739 9051 4755 9085
rect 4789 9051 4805 9085
rect 4739 9016 4805 9051
rect 4835 9085 4901 9120
rect 4835 9051 4851 9085
rect 4885 9051 4901 9085
rect 4835 9016 4901 9051
rect 4931 9085 4993 9120
rect 4931 9051 4947 9085
rect 4981 9051 4993 9085
rect 4931 9016 4993 9051
rect 5348 9155 5400 9167
rect 5348 9121 5356 9155
rect 5390 9121 5400 9155
rect 5348 9087 5400 9121
rect 5348 9053 5356 9087
rect 5390 9053 5400 9087
rect 5348 9037 5400 9053
rect 5430 9155 5482 9167
rect 5430 9121 5440 9155
rect 5474 9121 5482 9155
rect 5430 9087 5482 9121
rect 5430 9053 5440 9087
rect 5474 9053 5482 9087
rect 5430 9037 5482 9053
rect 301 7794 363 7829
rect 301 7760 313 7794
rect 347 7760 363 7794
rect 301 7725 363 7760
rect 393 7794 459 7829
rect 393 7760 409 7794
rect 443 7760 459 7794
rect 393 7725 459 7760
rect 489 7794 555 7829
rect 489 7760 505 7794
rect 539 7760 555 7794
rect 489 7725 555 7760
rect 585 7794 651 7829
rect 585 7760 601 7794
rect 635 7760 651 7794
rect 585 7725 651 7760
rect 681 7794 747 7829
rect 681 7760 697 7794
rect 731 7760 747 7794
rect 681 7725 747 7760
rect 777 7794 843 7829
rect 777 7760 793 7794
rect 827 7760 843 7794
rect 777 7725 843 7760
rect 873 7794 939 7829
rect 873 7760 889 7794
rect 923 7760 939 7794
rect 873 7725 939 7760
rect 969 7794 1035 7829
rect 969 7760 985 7794
rect 1019 7760 1035 7794
rect 969 7725 1035 7760
rect 1065 7794 1131 7829
rect 1065 7760 1081 7794
rect 1115 7760 1131 7794
rect 1065 7725 1131 7760
rect 1161 7794 1227 7829
rect 1161 7760 1177 7794
rect 1211 7760 1227 7794
rect 1161 7725 1227 7760
rect 1257 7794 1319 7829
rect 1257 7760 1273 7794
rect 1307 7760 1319 7794
rect 1257 7725 1319 7760
rect 2454 7798 2516 7833
rect 2454 7764 2466 7798
rect 2500 7764 2516 7798
rect 2454 7729 2516 7764
rect 2546 7798 2612 7833
rect 2546 7764 2562 7798
rect 2596 7764 2612 7798
rect 2546 7729 2612 7764
rect 2642 7798 2708 7833
rect 2642 7764 2658 7798
rect 2692 7764 2708 7798
rect 2642 7729 2708 7764
rect 2738 7798 2804 7833
rect 2738 7764 2754 7798
rect 2788 7764 2804 7798
rect 2738 7729 2804 7764
rect 2834 7798 2900 7833
rect 2834 7764 2850 7798
rect 2884 7764 2900 7798
rect 2834 7729 2900 7764
rect 2930 7798 2996 7833
rect 2930 7764 2946 7798
rect 2980 7764 2996 7798
rect 2930 7729 2996 7764
rect 3026 7798 3092 7833
rect 3026 7764 3042 7798
rect 3076 7764 3092 7798
rect 3026 7729 3092 7764
rect 3122 7798 3188 7833
rect 3122 7764 3138 7798
rect 3172 7764 3188 7798
rect 3122 7729 3188 7764
rect 3218 7798 3284 7833
rect 3218 7764 3234 7798
rect 3268 7764 3284 7798
rect 3218 7729 3284 7764
rect 3314 7798 3380 7833
rect 3314 7764 3330 7798
rect 3364 7764 3380 7798
rect 3314 7729 3380 7764
rect 3410 7798 3472 7833
rect 3410 7764 3426 7798
rect 3460 7764 3472 7798
rect 3410 7729 3472 7764
rect 3635 7825 3693 7837
rect 3635 7749 3647 7825
rect 3681 7749 3693 7825
rect 3635 7737 3693 7749
rect 3723 7825 3781 7837
rect 3723 7749 3735 7825
rect 3769 7749 3781 7825
rect 3723 7737 3781 7749
rect 3975 7798 4037 7833
rect 3975 7764 3987 7798
rect 4021 7764 4037 7798
rect 3975 7729 4037 7764
rect 4067 7798 4133 7833
rect 4067 7764 4083 7798
rect 4117 7764 4133 7798
rect 4067 7729 4133 7764
rect 4163 7798 4229 7833
rect 4163 7764 4179 7798
rect 4213 7764 4229 7798
rect 4163 7729 4229 7764
rect 4259 7798 4325 7833
rect 4259 7764 4275 7798
rect 4309 7764 4325 7798
rect 4259 7729 4325 7764
rect 4355 7798 4421 7833
rect 4355 7764 4371 7798
rect 4405 7764 4421 7798
rect 4355 7729 4421 7764
rect 4451 7798 4517 7833
rect 4451 7764 4467 7798
rect 4501 7764 4517 7798
rect 4451 7729 4517 7764
rect 4547 7798 4613 7833
rect 4547 7764 4563 7798
rect 4597 7764 4613 7798
rect 4547 7729 4613 7764
rect 4643 7798 4709 7833
rect 4643 7764 4659 7798
rect 4693 7764 4709 7798
rect 4643 7729 4709 7764
rect 4739 7798 4805 7833
rect 4739 7764 4755 7798
rect 4789 7764 4805 7798
rect 4739 7729 4805 7764
rect 4835 7798 4901 7833
rect 4835 7764 4851 7798
rect 4885 7764 4901 7798
rect 4835 7729 4901 7764
rect 4931 7798 4993 7833
rect 4931 7764 4947 7798
rect 4981 7764 4993 7798
rect 4931 7729 4993 7764
rect 5348 7868 5400 7880
rect 5348 7834 5356 7868
rect 5390 7834 5400 7868
rect 5348 7800 5400 7834
rect 5348 7766 5356 7800
rect 5390 7766 5400 7800
rect 5348 7750 5400 7766
rect 5430 7868 5482 7880
rect 5430 7834 5440 7868
rect 5474 7834 5482 7868
rect 5430 7800 5482 7834
rect 5430 7766 5440 7800
rect 5474 7766 5482 7800
rect 5430 7750 5482 7766
rect 301 6507 363 6542
rect 301 6473 313 6507
rect 347 6473 363 6507
rect 301 6438 363 6473
rect 393 6507 459 6542
rect 393 6473 409 6507
rect 443 6473 459 6507
rect 393 6438 459 6473
rect 489 6507 555 6542
rect 489 6473 505 6507
rect 539 6473 555 6507
rect 489 6438 555 6473
rect 585 6507 651 6542
rect 585 6473 601 6507
rect 635 6473 651 6507
rect 585 6438 651 6473
rect 681 6507 747 6542
rect 681 6473 697 6507
rect 731 6473 747 6507
rect 681 6438 747 6473
rect 777 6507 843 6542
rect 777 6473 793 6507
rect 827 6473 843 6507
rect 777 6438 843 6473
rect 873 6507 939 6542
rect 873 6473 889 6507
rect 923 6473 939 6507
rect 873 6438 939 6473
rect 969 6507 1035 6542
rect 969 6473 985 6507
rect 1019 6473 1035 6507
rect 969 6438 1035 6473
rect 1065 6507 1131 6542
rect 1065 6473 1081 6507
rect 1115 6473 1131 6507
rect 1065 6438 1131 6473
rect 1161 6507 1227 6542
rect 1161 6473 1177 6507
rect 1211 6473 1227 6507
rect 1161 6438 1227 6473
rect 1257 6507 1319 6542
rect 1257 6473 1273 6507
rect 1307 6473 1319 6507
rect 1257 6438 1319 6473
rect 2454 6511 2516 6546
rect 2454 6477 2466 6511
rect 2500 6477 2516 6511
rect 2454 6442 2516 6477
rect 2546 6511 2612 6546
rect 2546 6477 2562 6511
rect 2596 6477 2612 6511
rect 2546 6442 2612 6477
rect 2642 6511 2708 6546
rect 2642 6477 2658 6511
rect 2692 6477 2708 6511
rect 2642 6442 2708 6477
rect 2738 6511 2804 6546
rect 2738 6477 2754 6511
rect 2788 6477 2804 6511
rect 2738 6442 2804 6477
rect 2834 6511 2900 6546
rect 2834 6477 2850 6511
rect 2884 6477 2900 6511
rect 2834 6442 2900 6477
rect 2930 6511 2996 6546
rect 2930 6477 2946 6511
rect 2980 6477 2996 6511
rect 2930 6442 2996 6477
rect 3026 6511 3092 6546
rect 3026 6477 3042 6511
rect 3076 6477 3092 6511
rect 3026 6442 3092 6477
rect 3122 6511 3188 6546
rect 3122 6477 3138 6511
rect 3172 6477 3188 6511
rect 3122 6442 3188 6477
rect 3218 6511 3284 6546
rect 3218 6477 3234 6511
rect 3268 6477 3284 6511
rect 3218 6442 3284 6477
rect 3314 6511 3380 6546
rect 3314 6477 3330 6511
rect 3364 6477 3380 6511
rect 3314 6442 3380 6477
rect 3410 6511 3472 6546
rect 3410 6477 3426 6511
rect 3460 6477 3472 6511
rect 3410 6442 3472 6477
rect 3635 6538 3693 6550
rect 3635 6462 3647 6538
rect 3681 6462 3693 6538
rect 3635 6450 3693 6462
rect 3723 6538 3781 6550
rect 3723 6462 3735 6538
rect 3769 6462 3781 6538
rect 3723 6450 3781 6462
rect 3975 6511 4037 6546
rect 3975 6477 3987 6511
rect 4021 6477 4037 6511
rect 3975 6442 4037 6477
rect 4067 6511 4133 6546
rect 4067 6477 4083 6511
rect 4117 6477 4133 6511
rect 4067 6442 4133 6477
rect 4163 6511 4229 6546
rect 4163 6477 4179 6511
rect 4213 6477 4229 6511
rect 4163 6442 4229 6477
rect 4259 6511 4325 6546
rect 4259 6477 4275 6511
rect 4309 6477 4325 6511
rect 4259 6442 4325 6477
rect 4355 6511 4421 6546
rect 4355 6477 4371 6511
rect 4405 6477 4421 6511
rect 4355 6442 4421 6477
rect 4451 6511 4517 6546
rect 4451 6477 4467 6511
rect 4501 6477 4517 6511
rect 4451 6442 4517 6477
rect 4547 6511 4613 6546
rect 4547 6477 4563 6511
rect 4597 6477 4613 6511
rect 4547 6442 4613 6477
rect 4643 6511 4709 6546
rect 4643 6477 4659 6511
rect 4693 6477 4709 6511
rect 4643 6442 4709 6477
rect 4739 6511 4805 6546
rect 4739 6477 4755 6511
rect 4789 6477 4805 6511
rect 4739 6442 4805 6477
rect 4835 6511 4901 6546
rect 4835 6477 4851 6511
rect 4885 6477 4901 6511
rect 4835 6442 4901 6477
rect 4931 6511 4993 6546
rect 4931 6477 4947 6511
rect 4981 6477 4993 6511
rect 4931 6442 4993 6477
rect 5348 6581 5400 6593
rect 5348 6547 5356 6581
rect 5390 6547 5400 6581
rect 5348 6513 5400 6547
rect 5348 6479 5356 6513
rect 5390 6479 5400 6513
rect 5348 6463 5400 6479
rect 5430 6581 5482 6593
rect 5430 6547 5440 6581
rect 5474 6547 5482 6581
rect 5430 6513 5482 6547
rect 5430 6479 5440 6513
rect 5474 6479 5482 6513
rect 5430 6463 5482 6479
rect 301 5220 363 5255
rect 301 5186 313 5220
rect 347 5186 363 5220
rect 301 5151 363 5186
rect 393 5220 459 5255
rect 393 5186 409 5220
rect 443 5186 459 5220
rect 393 5151 459 5186
rect 489 5220 555 5255
rect 489 5186 505 5220
rect 539 5186 555 5220
rect 489 5151 555 5186
rect 585 5220 651 5255
rect 585 5186 601 5220
rect 635 5186 651 5220
rect 585 5151 651 5186
rect 681 5220 747 5255
rect 681 5186 697 5220
rect 731 5186 747 5220
rect 681 5151 747 5186
rect 777 5220 843 5255
rect 777 5186 793 5220
rect 827 5186 843 5220
rect 777 5151 843 5186
rect 873 5220 939 5255
rect 873 5186 889 5220
rect 923 5186 939 5220
rect 873 5151 939 5186
rect 969 5220 1035 5255
rect 969 5186 985 5220
rect 1019 5186 1035 5220
rect 969 5151 1035 5186
rect 1065 5220 1131 5255
rect 1065 5186 1081 5220
rect 1115 5186 1131 5220
rect 1065 5151 1131 5186
rect 1161 5220 1227 5255
rect 1161 5186 1177 5220
rect 1211 5186 1227 5220
rect 1161 5151 1227 5186
rect 1257 5220 1319 5255
rect 1257 5186 1273 5220
rect 1307 5186 1319 5220
rect 1257 5151 1319 5186
rect 2454 5224 2516 5259
rect 2454 5190 2466 5224
rect 2500 5190 2516 5224
rect 2454 5155 2516 5190
rect 2546 5224 2612 5259
rect 2546 5190 2562 5224
rect 2596 5190 2612 5224
rect 2546 5155 2612 5190
rect 2642 5224 2708 5259
rect 2642 5190 2658 5224
rect 2692 5190 2708 5224
rect 2642 5155 2708 5190
rect 2738 5224 2804 5259
rect 2738 5190 2754 5224
rect 2788 5190 2804 5224
rect 2738 5155 2804 5190
rect 2834 5224 2900 5259
rect 2834 5190 2850 5224
rect 2884 5190 2900 5224
rect 2834 5155 2900 5190
rect 2930 5224 2996 5259
rect 2930 5190 2946 5224
rect 2980 5190 2996 5224
rect 2930 5155 2996 5190
rect 3026 5224 3092 5259
rect 3026 5190 3042 5224
rect 3076 5190 3092 5224
rect 3026 5155 3092 5190
rect 3122 5224 3188 5259
rect 3122 5190 3138 5224
rect 3172 5190 3188 5224
rect 3122 5155 3188 5190
rect 3218 5224 3284 5259
rect 3218 5190 3234 5224
rect 3268 5190 3284 5224
rect 3218 5155 3284 5190
rect 3314 5224 3380 5259
rect 3314 5190 3330 5224
rect 3364 5190 3380 5224
rect 3314 5155 3380 5190
rect 3410 5224 3472 5259
rect 3410 5190 3426 5224
rect 3460 5190 3472 5224
rect 3410 5155 3472 5190
rect 3635 5251 3693 5263
rect 3635 5175 3647 5251
rect 3681 5175 3693 5251
rect 3635 5163 3693 5175
rect 3723 5251 3781 5263
rect 3723 5175 3735 5251
rect 3769 5175 3781 5251
rect 3723 5163 3781 5175
rect 3975 5224 4037 5259
rect 3975 5190 3987 5224
rect 4021 5190 4037 5224
rect 3975 5155 4037 5190
rect 4067 5224 4133 5259
rect 4067 5190 4083 5224
rect 4117 5190 4133 5224
rect 4067 5155 4133 5190
rect 4163 5224 4229 5259
rect 4163 5190 4179 5224
rect 4213 5190 4229 5224
rect 4163 5155 4229 5190
rect 4259 5224 4325 5259
rect 4259 5190 4275 5224
rect 4309 5190 4325 5224
rect 4259 5155 4325 5190
rect 4355 5224 4421 5259
rect 4355 5190 4371 5224
rect 4405 5190 4421 5224
rect 4355 5155 4421 5190
rect 4451 5224 4517 5259
rect 4451 5190 4467 5224
rect 4501 5190 4517 5224
rect 4451 5155 4517 5190
rect 4547 5224 4613 5259
rect 4547 5190 4563 5224
rect 4597 5190 4613 5224
rect 4547 5155 4613 5190
rect 4643 5224 4709 5259
rect 4643 5190 4659 5224
rect 4693 5190 4709 5224
rect 4643 5155 4709 5190
rect 4739 5224 4805 5259
rect 4739 5190 4755 5224
rect 4789 5190 4805 5224
rect 4739 5155 4805 5190
rect 4835 5224 4901 5259
rect 4835 5190 4851 5224
rect 4885 5190 4901 5224
rect 4835 5155 4901 5190
rect 4931 5224 4993 5259
rect 4931 5190 4947 5224
rect 4981 5190 4993 5224
rect 4931 5155 4993 5190
rect 5348 5294 5400 5306
rect 5348 5260 5356 5294
rect 5390 5260 5400 5294
rect 5348 5226 5400 5260
rect 5348 5192 5356 5226
rect 5390 5192 5400 5226
rect 5348 5176 5400 5192
rect 5430 5294 5482 5306
rect 5430 5260 5440 5294
rect 5474 5260 5482 5294
rect 5430 5226 5482 5260
rect 5430 5192 5440 5226
rect 5474 5192 5482 5226
rect 5430 5176 5482 5192
rect 301 3933 363 3968
rect 301 3899 313 3933
rect 347 3899 363 3933
rect 301 3864 363 3899
rect 393 3933 459 3968
rect 393 3899 409 3933
rect 443 3899 459 3933
rect 393 3864 459 3899
rect 489 3933 555 3968
rect 489 3899 505 3933
rect 539 3899 555 3933
rect 489 3864 555 3899
rect 585 3933 651 3968
rect 585 3899 601 3933
rect 635 3899 651 3933
rect 585 3864 651 3899
rect 681 3933 747 3968
rect 681 3899 697 3933
rect 731 3899 747 3933
rect 681 3864 747 3899
rect 777 3933 843 3968
rect 777 3899 793 3933
rect 827 3899 843 3933
rect 777 3864 843 3899
rect 873 3933 939 3968
rect 873 3899 889 3933
rect 923 3899 939 3933
rect 873 3864 939 3899
rect 969 3933 1035 3968
rect 969 3899 985 3933
rect 1019 3899 1035 3933
rect 969 3864 1035 3899
rect 1065 3933 1131 3968
rect 1065 3899 1081 3933
rect 1115 3899 1131 3933
rect 1065 3864 1131 3899
rect 1161 3933 1227 3968
rect 1161 3899 1177 3933
rect 1211 3899 1227 3933
rect 1161 3864 1227 3899
rect 1257 3933 1319 3968
rect 1257 3899 1273 3933
rect 1307 3899 1319 3933
rect 1257 3864 1319 3899
rect 2454 3937 2516 3972
rect 2454 3903 2466 3937
rect 2500 3903 2516 3937
rect 2454 3868 2516 3903
rect 2546 3937 2612 3972
rect 2546 3903 2562 3937
rect 2596 3903 2612 3937
rect 2546 3868 2612 3903
rect 2642 3937 2708 3972
rect 2642 3903 2658 3937
rect 2692 3903 2708 3937
rect 2642 3868 2708 3903
rect 2738 3937 2804 3972
rect 2738 3903 2754 3937
rect 2788 3903 2804 3937
rect 2738 3868 2804 3903
rect 2834 3937 2900 3972
rect 2834 3903 2850 3937
rect 2884 3903 2900 3937
rect 2834 3868 2900 3903
rect 2930 3937 2996 3972
rect 2930 3903 2946 3937
rect 2980 3903 2996 3937
rect 2930 3868 2996 3903
rect 3026 3937 3092 3972
rect 3026 3903 3042 3937
rect 3076 3903 3092 3937
rect 3026 3868 3092 3903
rect 3122 3937 3188 3972
rect 3122 3903 3138 3937
rect 3172 3903 3188 3937
rect 3122 3868 3188 3903
rect 3218 3937 3284 3972
rect 3218 3903 3234 3937
rect 3268 3903 3284 3937
rect 3218 3868 3284 3903
rect 3314 3937 3380 3972
rect 3314 3903 3330 3937
rect 3364 3903 3380 3937
rect 3314 3868 3380 3903
rect 3410 3937 3472 3972
rect 3410 3903 3426 3937
rect 3460 3903 3472 3937
rect 3410 3868 3472 3903
rect 3635 3964 3693 3976
rect 3635 3888 3647 3964
rect 3681 3888 3693 3964
rect 3635 3876 3693 3888
rect 3723 3964 3781 3976
rect 3723 3888 3735 3964
rect 3769 3888 3781 3964
rect 3723 3876 3781 3888
rect 3975 3937 4037 3972
rect 3975 3903 3987 3937
rect 4021 3903 4037 3937
rect 3975 3868 4037 3903
rect 4067 3937 4133 3972
rect 4067 3903 4083 3937
rect 4117 3903 4133 3937
rect 4067 3868 4133 3903
rect 4163 3937 4229 3972
rect 4163 3903 4179 3937
rect 4213 3903 4229 3937
rect 4163 3868 4229 3903
rect 4259 3937 4325 3972
rect 4259 3903 4275 3937
rect 4309 3903 4325 3937
rect 4259 3868 4325 3903
rect 4355 3937 4421 3972
rect 4355 3903 4371 3937
rect 4405 3903 4421 3937
rect 4355 3868 4421 3903
rect 4451 3937 4517 3972
rect 4451 3903 4467 3937
rect 4501 3903 4517 3937
rect 4451 3868 4517 3903
rect 4547 3937 4613 3972
rect 4547 3903 4563 3937
rect 4597 3903 4613 3937
rect 4547 3868 4613 3903
rect 4643 3937 4709 3972
rect 4643 3903 4659 3937
rect 4693 3903 4709 3937
rect 4643 3868 4709 3903
rect 4739 3937 4805 3972
rect 4739 3903 4755 3937
rect 4789 3903 4805 3937
rect 4739 3868 4805 3903
rect 4835 3937 4901 3972
rect 4835 3903 4851 3937
rect 4885 3903 4901 3937
rect 4835 3868 4901 3903
rect 4931 3937 4993 3972
rect 4931 3903 4947 3937
rect 4981 3903 4993 3937
rect 4931 3868 4993 3903
rect 5348 4007 5400 4019
rect 5348 3973 5356 4007
rect 5390 3973 5400 4007
rect 5348 3939 5400 3973
rect 5348 3905 5356 3939
rect 5390 3905 5400 3939
rect 5348 3889 5400 3905
rect 5430 4007 5482 4019
rect 5430 3973 5440 4007
rect 5474 3973 5482 4007
rect 5430 3939 5482 3973
rect 5430 3905 5440 3939
rect 5474 3905 5482 3939
rect 5430 3889 5482 3905
rect 301 2646 363 2681
rect 301 2612 313 2646
rect 347 2612 363 2646
rect 301 2577 363 2612
rect 393 2646 459 2681
rect 393 2612 409 2646
rect 443 2612 459 2646
rect 393 2577 459 2612
rect 489 2646 555 2681
rect 489 2612 505 2646
rect 539 2612 555 2646
rect 489 2577 555 2612
rect 585 2646 651 2681
rect 585 2612 601 2646
rect 635 2612 651 2646
rect 585 2577 651 2612
rect 681 2646 747 2681
rect 681 2612 697 2646
rect 731 2612 747 2646
rect 681 2577 747 2612
rect 777 2646 843 2681
rect 777 2612 793 2646
rect 827 2612 843 2646
rect 777 2577 843 2612
rect 873 2646 939 2681
rect 873 2612 889 2646
rect 923 2612 939 2646
rect 873 2577 939 2612
rect 969 2646 1035 2681
rect 969 2612 985 2646
rect 1019 2612 1035 2646
rect 969 2577 1035 2612
rect 1065 2646 1131 2681
rect 1065 2612 1081 2646
rect 1115 2612 1131 2646
rect 1065 2577 1131 2612
rect 1161 2646 1227 2681
rect 1161 2612 1177 2646
rect 1211 2612 1227 2646
rect 1161 2577 1227 2612
rect 1257 2646 1319 2681
rect 1257 2612 1273 2646
rect 1307 2612 1319 2646
rect 1257 2577 1319 2612
rect 2454 2650 2516 2685
rect 2454 2616 2466 2650
rect 2500 2616 2516 2650
rect 2454 2581 2516 2616
rect 2546 2650 2612 2685
rect 2546 2616 2562 2650
rect 2596 2616 2612 2650
rect 2546 2581 2612 2616
rect 2642 2650 2708 2685
rect 2642 2616 2658 2650
rect 2692 2616 2708 2650
rect 2642 2581 2708 2616
rect 2738 2650 2804 2685
rect 2738 2616 2754 2650
rect 2788 2616 2804 2650
rect 2738 2581 2804 2616
rect 2834 2650 2900 2685
rect 2834 2616 2850 2650
rect 2884 2616 2900 2650
rect 2834 2581 2900 2616
rect 2930 2650 2996 2685
rect 2930 2616 2946 2650
rect 2980 2616 2996 2650
rect 2930 2581 2996 2616
rect 3026 2650 3092 2685
rect 3026 2616 3042 2650
rect 3076 2616 3092 2650
rect 3026 2581 3092 2616
rect 3122 2650 3188 2685
rect 3122 2616 3138 2650
rect 3172 2616 3188 2650
rect 3122 2581 3188 2616
rect 3218 2650 3284 2685
rect 3218 2616 3234 2650
rect 3268 2616 3284 2650
rect 3218 2581 3284 2616
rect 3314 2650 3380 2685
rect 3314 2616 3330 2650
rect 3364 2616 3380 2650
rect 3314 2581 3380 2616
rect 3410 2650 3472 2685
rect 3410 2616 3426 2650
rect 3460 2616 3472 2650
rect 3410 2581 3472 2616
rect 3635 2677 3693 2689
rect 3635 2601 3647 2677
rect 3681 2601 3693 2677
rect 3635 2589 3693 2601
rect 3723 2677 3781 2689
rect 3723 2601 3735 2677
rect 3769 2601 3781 2677
rect 3723 2589 3781 2601
rect 3975 2650 4037 2685
rect 3975 2616 3987 2650
rect 4021 2616 4037 2650
rect 3975 2581 4037 2616
rect 4067 2650 4133 2685
rect 4067 2616 4083 2650
rect 4117 2616 4133 2650
rect 4067 2581 4133 2616
rect 4163 2650 4229 2685
rect 4163 2616 4179 2650
rect 4213 2616 4229 2650
rect 4163 2581 4229 2616
rect 4259 2650 4325 2685
rect 4259 2616 4275 2650
rect 4309 2616 4325 2650
rect 4259 2581 4325 2616
rect 4355 2650 4421 2685
rect 4355 2616 4371 2650
rect 4405 2616 4421 2650
rect 4355 2581 4421 2616
rect 4451 2650 4517 2685
rect 4451 2616 4467 2650
rect 4501 2616 4517 2650
rect 4451 2581 4517 2616
rect 4547 2650 4613 2685
rect 4547 2616 4563 2650
rect 4597 2616 4613 2650
rect 4547 2581 4613 2616
rect 4643 2650 4709 2685
rect 4643 2616 4659 2650
rect 4693 2616 4709 2650
rect 4643 2581 4709 2616
rect 4739 2650 4805 2685
rect 4739 2616 4755 2650
rect 4789 2616 4805 2650
rect 4739 2581 4805 2616
rect 4835 2650 4901 2685
rect 4835 2616 4851 2650
rect 4885 2616 4901 2650
rect 4835 2581 4901 2616
rect 4931 2650 4993 2685
rect 4931 2616 4947 2650
rect 4981 2616 4993 2650
rect 4931 2581 4993 2616
rect 5348 2720 5400 2732
rect 5348 2686 5356 2720
rect 5390 2686 5400 2720
rect 5348 2652 5400 2686
rect 5348 2618 5356 2652
rect 5390 2618 5400 2652
rect 5348 2602 5400 2618
rect 5430 2720 5482 2732
rect 5430 2686 5440 2720
rect 5474 2686 5482 2720
rect 5430 2652 5482 2686
rect 5430 2618 5440 2652
rect 5474 2618 5482 2652
rect 5430 2602 5482 2618
rect 301 1359 363 1394
rect 301 1325 313 1359
rect 347 1325 363 1359
rect 301 1290 363 1325
rect 393 1359 459 1394
rect 393 1325 409 1359
rect 443 1325 459 1359
rect 393 1290 459 1325
rect 489 1359 555 1394
rect 489 1325 505 1359
rect 539 1325 555 1359
rect 489 1290 555 1325
rect 585 1359 651 1394
rect 585 1325 601 1359
rect 635 1325 651 1359
rect 585 1290 651 1325
rect 681 1359 747 1394
rect 681 1325 697 1359
rect 731 1325 747 1359
rect 681 1290 747 1325
rect 777 1359 843 1394
rect 777 1325 793 1359
rect 827 1325 843 1359
rect 777 1290 843 1325
rect 873 1359 939 1394
rect 873 1325 889 1359
rect 923 1325 939 1359
rect 873 1290 939 1325
rect 969 1359 1035 1394
rect 969 1325 985 1359
rect 1019 1325 1035 1359
rect 969 1290 1035 1325
rect 1065 1359 1131 1394
rect 1065 1325 1081 1359
rect 1115 1325 1131 1359
rect 1065 1290 1131 1325
rect 1161 1359 1227 1394
rect 1161 1325 1177 1359
rect 1211 1325 1227 1359
rect 1161 1290 1227 1325
rect 1257 1359 1319 1394
rect 1257 1325 1273 1359
rect 1307 1325 1319 1359
rect 1257 1290 1319 1325
rect 2454 1363 2516 1398
rect 2454 1329 2466 1363
rect 2500 1329 2516 1363
rect 2454 1294 2516 1329
rect 2546 1363 2612 1398
rect 2546 1329 2562 1363
rect 2596 1329 2612 1363
rect 2546 1294 2612 1329
rect 2642 1363 2708 1398
rect 2642 1329 2658 1363
rect 2692 1329 2708 1363
rect 2642 1294 2708 1329
rect 2738 1363 2804 1398
rect 2738 1329 2754 1363
rect 2788 1329 2804 1363
rect 2738 1294 2804 1329
rect 2834 1363 2900 1398
rect 2834 1329 2850 1363
rect 2884 1329 2900 1363
rect 2834 1294 2900 1329
rect 2930 1363 2996 1398
rect 2930 1329 2946 1363
rect 2980 1329 2996 1363
rect 2930 1294 2996 1329
rect 3026 1363 3092 1398
rect 3026 1329 3042 1363
rect 3076 1329 3092 1363
rect 3026 1294 3092 1329
rect 3122 1363 3188 1398
rect 3122 1329 3138 1363
rect 3172 1329 3188 1363
rect 3122 1294 3188 1329
rect 3218 1363 3284 1398
rect 3218 1329 3234 1363
rect 3268 1329 3284 1363
rect 3218 1294 3284 1329
rect 3314 1363 3380 1398
rect 3314 1329 3330 1363
rect 3364 1329 3380 1363
rect 3314 1294 3380 1329
rect 3410 1363 3472 1398
rect 3410 1329 3426 1363
rect 3460 1329 3472 1363
rect 3410 1294 3472 1329
rect 3635 1390 3693 1402
rect 3635 1314 3647 1390
rect 3681 1314 3693 1390
rect 3635 1302 3693 1314
rect 3723 1390 3781 1402
rect 3723 1314 3735 1390
rect 3769 1314 3781 1390
rect 3723 1302 3781 1314
rect 3975 1363 4037 1398
rect 3975 1329 3987 1363
rect 4021 1329 4037 1363
rect 3975 1294 4037 1329
rect 4067 1363 4133 1398
rect 4067 1329 4083 1363
rect 4117 1329 4133 1363
rect 4067 1294 4133 1329
rect 4163 1363 4229 1398
rect 4163 1329 4179 1363
rect 4213 1329 4229 1363
rect 4163 1294 4229 1329
rect 4259 1363 4325 1398
rect 4259 1329 4275 1363
rect 4309 1329 4325 1363
rect 4259 1294 4325 1329
rect 4355 1363 4421 1398
rect 4355 1329 4371 1363
rect 4405 1329 4421 1363
rect 4355 1294 4421 1329
rect 4451 1363 4517 1398
rect 4451 1329 4467 1363
rect 4501 1329 4517 1363
rect 4451 1294 4517 1329
rect 4547 1363 4613 1398
rect 4547 1329 4563 1363
rect 4597 1329 4613 1363
rect 4547 1294 4613 1329
rect 4643 1363 4709 1398
rect 4643 1329 4659 1363
rect 4693 1329 4709 1363
rect 4643 1294 4709 1329
rect 4739 1363 4805 1398
rect 4739 1329 4755 1363
rect 4789 1329 4805 1363
rect 4739 1294 4805 1329
rect 4835 1363 4901 1398
rect 4835 1329 4851 1363
rect 4885 1329 4901 1363
rect 4835 1294 4901 1329
rect 4931 1363 4993 1398
rect 4931 1329 4947 1363
rect 4981 1329 4993 1363
rect 4931 1294 4993 1329
rect 5348 1433 5400 1445
rect 5348 1399 5356 1433
rect 5390 1399 5400 1433
rect 5348 1365 5400 1399
rect 5348 1331 5356 1365
rect 5390 1331 5400 1365
rect 5348 1315 5400 1331
rect 5430 1433 5482 1445
rect 5430 1399 5440 1433
rect 5474 1399 5482 1433
rect 5430 1365 5482 1399
rect 5430 1331 5440 1365
rect 5474 1331 5482 1365
rect 5430 1315 5482 1331
<< pdiff >>
rect 301 41854 363 41871
rect 301 41820 313 41854
rect 347 41820 363 41854
rect 301 41786 363 41820
rect 301 41752 313 41786
rect 347 41752 363 41786
rect 301 41718 363 41752
rect 301 41684 313 41718
rect 347 41684 363 41718
rect 301 41650 363 41684
rect 301 41616 313 41650
rect 347 41616 363 41650
rect 301 41599 363 41616
rect 393 41854 459 41871
rect 393 41820 409 41854
rect 443 41820 459 41854
rect 393 41786 459 41820
rect 393 41752 409 41786
rect 443 41752 459 41786
rect 393 41718 459 41752
rect 393 41684 409 41718
rect 443 41684 459 41718
rect 393 41650 459 41684
rect 393 41616 409 41650
rect 443 41616 459 41650
rect 393 41599 459 41616
rect 489 41854 555 41871
rect 489 41820 505 41854
rect 539 41820 555 41854
rect 489 41786 555 41820
rect 489 41752 505 41786
rect 539 41752 555 41786
rect 489 41718 555 41752
rect 489 41684 505 41718
rect 539 41684 555 41718
rect 489 41650 555 41684
rect 489 41616 505 41650
rect 539 41616 555 41650
rect 489 41599 555 41616
rect 585 41854 651 41871
rect 585 41820 601 41854
rect 635 41820 651 41854
rect 585 41786 651 41820
rect 585 41752 601 41786
rect 635 41752 651 41786
rect 585 41718 651 41752
rect 585 41684 601 41718
rect 635 41684 651 41718
rect 585 41650 651 41684
rect 585 41616 601 41650
rect 635 41616 651 41650
rect 585 41599 651 41616
rect 681 41854 747 41871
rect 681 41820 697 41854
rect 731 41820 747 41854
rect 681 41786 747 41820
rect 681 41752 697 41786
rect 731 41752 747 41786
rect 681 41718 747 41752
rect 681 41684 697 41718
rect 731 41684 747 41718
rect 681 41650 747 41684
rect 681 41616 697 41650
rect 731 41616 747 41650
rect 681 41599 747 41616
rect 777 41854 843 41871
rect 777 41820 793 41854
rect 827 41820 843 41854
rect 777 41786 843 41820
rect 777 41752 793 41786
rect 827 41752 843 41786
rect 777 41718 843 41752
rect 777 41684 793 41718
rect 827 41684 843 41718
rect 777 41650 843 41684
rect 777 41616 793 41650
rect 827 41616 843 41650
rect 777 41599 843 41616
rect 873 41854 939 41871
rect 873 41820 889 41854
rect 923 41820 939 41854
rect 873 41786 939 41820
rect 873 41752 889 41786
rect 923 41752 939 41786
rect 873 41718 939 41752
rect 873 41684 889 41718
rect 923 41684 939 41718
rect 873 41650 939 41684
rect 873 41616 889 41650
rect 923 41616 939 41650
rect 873 41599 939 41616
rect 969 41854 1035 41871
rect 969 41820 985 41854
rect 1019 41820 1035 41854
rect 969 41786 1035 41820
rect 969 41752 985 41786
rect 1019 41752 1035 41786
rect 969 41718 1035 41752
rect 969 41684 985 41718
rect 1019 41684 1035 41718
rect 969 41650 1035 41684
rect 969 41616 985 41650
rect 1019 41616 1035 41650
rect 969 41599 1035 41616
rect 1065 41854 1131 41871
rect 1065 41820 1081 41854
rect 1115 41820 1131 41854
rect 1065 41786 1131 41820
rect 1065 41752 1081 41786
rect 1115 41752 1131 41786
rect 1065 41718 1131 41752
rect 1065 41684 1081 41718
rect 1115 41684 1131 41718
rect 1065 41650 1131 41684
rect 1065 41616 1081 41650
rect 1115 41616 1131 41650
rect 1065 41599 1131 41616
rect 1161 41854 1227 41871
rect 1161 41820 1177 41854
rect 1211 41820 1227 41854
rect 1161 41786 1227 41820
rect 1161 41752 1177 41786
rect 1211 41752 1227 41786
rect 1161 41718 1227 41752
rect 1161 41684 1177 41718
rect 1211 41684 1227 41718
rect 1161 41650 1227 41684
rect 1161 41616 1177 41650
rect 1211 41616 1227 41650
rect 1161 41599 1227 41616
rect 1257 41854 1319 41871
rect 1257 41820 1273 41854
rect 1307 41820 1319 41854
rect 1257 41786 1319 41820
rect 1257 41752 1273 41786
rect 1307 41752 1319 41786
rect 1257 41718 1319 41752
rect 1257 41684 1273 41718
rect 1307 41684 1319 41718
rect 1257 41650 1319 41684
rect 1257 41616 1273 41650
rect 1307 41616 1319 41650
rect 1257 41599 1319 41616
rect 2454 41858 2516 41875
rect 2454 41824 2466 41858
rect 2500 41824 2516 41858
rect 2454 41790 2516 41824
rect 2454 41756 2466 41790
rect 2500 41756 2516 41790
rect 2454 41722 2516 41756
rect 2454 41688 2466 41722
rect 2500 41688 2516 41722
rect 2454 41654 2516 41688
rect 2454 41620 2466 41654
rect 2500 41620 2516 41654
rect 2454 41603 2516 41620
rect 2546 41858 2612 41875
rect 2546 41824 2562 41858
rect 2596 41824 2612 41858
rect 2546 41790 2612 41824
rect 2546 41756 2562 41790
rect 2596 41756 2612 41790
rect 2546 41722 2612 41756
rect 2546 41688 2562 41722
rect 2596 41688 2612 41722
rect 2546 41654 2612 41688
rect 2546 41620 2562 41654
rect 2596 41620 2612 41654
rect 2546 41603 2612 41620
rect 2642 41858 2708 41875
rect 2642 41824 2658 41858
rect 2692 41824 2708 41858
rect 2642 41790 2708 41824
rect 2642 41756 2658 41790
rect 2692 41756 2708 41790
rect 2642 41722 2708 41756
rect 2642 41688 2658 41722
rect 2692 41688 2708 41722
rect 2642 41654 2708 41688
rect 2642 41620 2658 41654
rect 2692 41620 2708 41654
rect 2642 41603 2708 41620
rect 2738 41858 2804 41875
rect 2738 41824 2754 41858
rect 2788 41824 2804 41858
rect 2738 41790 2804 41824
rect 2738 41756 2754 41790
rect 2788 41756 2804 41790
rect 2738 41722 2804 41756
rect 2738 41688 2754 41722
rect 2788 41688 2804 41722
rect 2738 41654 2804 41688
rect 2738 41620 2754 41654
rect 2788 41620 2804 41654
rect 2738 41603 2804 41620
rect 2834 41858 2900 41875
rect 2834 41824 2850 41858
rect 2884 41824 2900 41858
rect 2834 41790 2900 41824
rect 2834 41756 2850 41790
rect 2884 41756 2900 41790
rect 2834 41722 2900 41756
rect 2834 41688 2850 41722
rect 2884 41688 2900 41722
rect 2834 41654 2900 41688
rect 2834 41620 2850 41654
rect 2884 41620 2900 41654
rect 2834 41603 2900 41620
rect 2930 41858 2996 41875
rect 2930 41824 2946 41858
rect 2980 41824 2996 41858
rect 2930 41790 2996 41824
rect 2930 41756 2946 41790
rect 2980 41756 2996 41790
rect 2930 41722 2996 41756
rect 2930 41688 2946 41722
rect 2980 41688 2996 41722
rect 2930 41654 2996 41688
rect 2930 41620 2946 41654
rect 2980 41620 2996 41654
rect 2930 41603 2996 41620
rect 3026 41858 3092 41875
rect 3026 41824 3042 41858
rect 3076 41824 3092 41858
rect 3026 41790 3092 41824
rect 3026 41756 3042 41790
rect 3076 41756 3092 41790
rect 3026 41722 3092 41756
rect 3026 41688 3042 41722
rect 3076 41688 3092 41722
rect 3026 41654 3092 41688
rect 3026 41620 3042 41654
rect 3076 41620 3092 41654
rect 3026 41603 3092 41620
rect 3122 41858 3188 41875
rect 3122 41824 3138 41858
rect 3172 41824 3188 41858
rect 3122 41790 3188 41824
rect 3122 41756 3138 41790
rect 3172 41756 3188 41790
rect 3122 41722 3188 41756
rect 3122 41688 3138 41722
rect 3172 41688 3188 41722
rect 3122 41654 3188 41688
rect 3122 41620 3138 41654
rect 3172 41620 3188 41654
rect 3122 41603 3188 41620
rect 3218 41858 3284 41875
rect 3218 41824 3234 41858
rect 3268 41824 3284 41858
rect 3218 41790 3284 41824
rect 3218 41756 3234 41790
rect 3268 41756 3284 41790
rect 3218 41722 3284 41756
rect 3218 41688 3234 41722
rect 3268 41688 3284 41722
rect 3218 41654 3284 41688
rect 3218 41620 3234 41654
rect 3268 41620 3284 41654
rect 3218 41603 3284 41620
rect 3314 41858 3380 41875
rect 3314 41824 3330 41858
rect 3364 41824 3380 41858
rect 3314 41790 3380 41824
rect 3314 41756 3330 41790
rect 3364 41756 3380 41790
rect 3314 41722 3380 41756
rect 3314 41688 3330 41722
rect 3364 41688 3380 41722
rect 3314 41654 3380 41688
rect 3314 41620 3330 41654
rect 3364 41620 3380 41654
rect 3314 41603 3380 41620
rect 3410 41858 3472 41875
rect 3410 41824 3426 41858
rect 3460 41824 3472 41858
rect 3410 41790 3472 41824
rect 3410 41756 3426 41790
rect 3460 41756 3472 41790
rect 3410 41722 3472 41756
rect 3410 41688 3426 41722
rect 3460 41688 3472 41722
rect 3410 41654 3472 41688
rect 3410 41620 3426 41654
rect 3460 41620 3472 41654
rect 3410 41603 3472 41620
rect 3975 41858 4037 41875
rect 3975 41824 3987 41858
rect 4021 41824 4037 41858
rect 3975 41790 4037 41824
rect 3975 41756 3987 41790
rect 4021 41756 4037 41790
rect 3975 41722 4037 41756
rect 3975 41688 3987 41722
rect 4021 41688 4037 41722
rect 3975 41654 4037 41688
rect 3975 41620 3987 41654
rect 4021 41620 4037 41654
rect 3975 41603 4037 41620
rect 4067 41858 4133 41875
rect 4067 41824 4083 41858
rect 4117 41824 4133 41858
rect 4067 41790 4133 41824
rect 4067 41756 4083 41790
rect 4117 41756 4133 41790
rect 4067 41722 4133 41756
rect 4067 41688 4083 41722
rect 4117 41688 4133 41722
rect 4067 41654 4133 41688
rect 4067 41620 4083 41654
rect 4117 41620 4133 41654
rect 4067 41603 4133 41620
rect 4163 41858 4229 41875
rect 4163 41824 4179 41858
rect 4213 41824 4229 41858
rect 4163 41790 4229 41824
rect 4163 41756 4179 41790
rect 4213 41756 4229 41790
rect 4163 41722 4229 41756
rect 4163 41688 4179 41722
rect 4213 41688 4229 41722
rect 4163 41654 4229 41688
rect 4163 41620 4179 41654
rect 4213 41620 4229 41654
rect 4163 41603 4229 41620
rect 4259 41858 4325 41875
rect 4259 41824 4275 41858
rect 4309 41824 4325 41858
rect 4259 41790 4325 41824
rect 4259 41756 4275 41790
rect 4309 41756 4325 41790
rect 4259 41722 4325 41756
rect 4259 41688 4275 41722
rect 4309 41688 4325 41722
rect 4259 41654 4325 41688
rect 4259 41620 4275 41654
rect 4309 41620 4325 41654
rect 4259 41603 4325 41620
rect 4355 41858 4421 41875
rect 4355 41824 4371 41858
rect 4405 41824 4421 41858
rect 4355 41790 4421 41824
rect 4355 41756 4371 41790
rect 4405 41756 4421 41790
rect 4355 41722 4421 41756
rect 4355 41688 4371 41722
rect 4405 41688 4421 41722
rect 4355 41654 4421 41688
rect 4355 41620 4371 41654
rect 4405 41620 4421 41654
rect 4355 41603 4421 41620
rect 4451 41858 4517 41875
rect 4451 41824 4467 41858
rect 4501 41824 4517 41858
rect 4451 41790 4517 41824
rect 4451 41756 4467 41790
rect 4501 41756 4517 41790
rect 4451 41722 4517 41756
rect 4451 41688 4467 41722
rect 4501 41688 4517 41722
rect 4451 41654 4517 41688
rect 4451 41620 4467 41654
rect 4501 41620 4517 41654
rect 4451 41603 4517 41620
rect 4547 41858 4613 41875
rect 4547 41824 4563 41858
rect 4597 41824 4613 41858
rect 4547 41790 4613 41824
rect 4547 41756 4563 41790
rect 4597 41756 4613 41790
rect 4547 41722 4613 41756
rect 4547 41688 4563 41722
rect 4597 41688 4613 41722
rect 4547 41654 4613 41688
rect 4547 41620 4563 41654
rect 4597 41620 4613 41654
rect 4547 41603 4613 41620
rect 4643 41858 4709 41875
rect 4643 41824 4659 41858
rect 4693 41824 4709 41858
rect 4643 41790 4709 41824
rect 4643 41756 4659 41790
rect 4693 41756 4709 41790
rect 4643 41722 4709 41756
rect 4643 41688 4659 41722
rect 4693 41688 4709 41722
rect 4643 41654 4709 41688
rect 4643 41620 4659 41654
rect 4693 41620 4709 41654
rect 4643 41603 4709 41620
rect 4739 41858 4805 41875
rect 4739 41824 4755 41858
rect 4789 41824 4805 41858
rect 4739 41790 4805 41824
rect 4739 41756 4755 41790
rect 4789 41756 4805 41790
rect 4739 41722 4805 41756
rect 4739 41688 4755 41722
rect 4789 41688 4805 41722
rect 4739 41654 4805 41688
rect 4739 41620 4755 41654
rect 4789 41620 4805 41654
rect 4739 41603 4805 41620
rect 4835 41858 4901 41875
rect 4835 41824 4851 41858
rect 4885 41824 4901 41858
rect 4835 41790 4901 41824
rect 4835 41756 4851 41790
rect 4885 41756 4901 41790
rect 4835 41722 4901 41756
rect 4835 41688 4851 41722
rect 4885 41688 4901 41722
rect 4835 41654 4901 41688
rect 4835 41620 4851 41654
rect 4885 41620 4901 41654
rect 4835 41603 4901 41620
rect 4931 41858 4993 41875
rect 4931 41824 4947 41858
rect 4981 41824 4993 41858
rect 4931 41790 4993 41824
rect 4931 41756 4947 41790
rect 4981 41756 4993 41790
rect 4931 41722 4993 41756
rect 4931 41688 4947 41722
rect 4981 41688 4993 41722
rect 4931 41654 4993 41688
rect 4931 41620 4947 41654
rect 4981 41620 4993 41654
rect 4931 41603 4993 41620
rect 5348 41650 5400 41662
rect 5348 41616 5356 41650
rect 5390 41616 5400 41650
rect 5348 41582 5400 41616
rect 5348 41548 5356 41582
rect 5390 41548 5400 41582
rect 5348 41514 5400 41548
rect 5348 41480 5356 41514
rect 5390 41480 5400 41514
rect 5348 41462 5400 41480
rect 5430 41650 5482 41662
rect 5430 41616 5440 41650
rect 5474 41616 5482 41650
rect 5430 41582 5482 41616
rect 5430 41548 5440 41582
rect 5474 41548 5482 41582
rect 5430 41514 5482 41548
rect 5430 41480 5440 41514
rect 5474 41480 5482 41514
rect 5430 41462 5482 41480
rect 301 40567 363 40584
rect 301 40533 313 40567
rect 347 40533 363 40567
rect 301 40499 363 40533
rect 301 40465 313 40499
rect 347 40465 363 40499
rect 301 40431 363 40465
rect 301 40397 313 40431
rect 347 40397 363 40431
rect 301 40363 363 40397
rect 301 40329 313 40363
rect 347 40329 363 40363
rect 301 40312 363 40329
rect 393 40567 459 40584
rect 393 40533 409 40567
rect 443 40533 459 40567
rect 393 40499 459 40533
rect 393 40465 409 40499
rect 443 40465 459 40499
rect 393 40431 459 40465
rect 393 40397 409 40431
rect 443 40397 459 40431
rect 393 40363 459 40397
rect 393 40329 409 40363
rect 443 40329 459 40363
rect 393 40312 459 40329
rect 489 40567 555 40584
rect 489 40533 505 40567
rect 539 40533 555 40567
rect 489 40499 555 40533
rect 489 40465 505 40499
rect 539 40465 555 40499
rect 489 40431 555 40465
rect 489 40397 505 40431
rect 539 40397 555 40431
rect 489 40363 555 40397
rect 489 40329 505 40363
rect 539 40329 555 40363
rect 489 40312 555 40329
rect 585 40567 651 40584
rect 585 40533 601 40567
rect 635 40533 651 40567
rect 585 40499 651 40533
rect 585 40465 601 40499
rect 635 40465 651 40499
rect 585 40431 651 40465
rect 585 40397 601 40431
rect 635 40397 651 40431
rect 585 40363 651 40397
rect 585 40329 601 40363
rect 635 40329 651 40363
rect 585 40312 651 40329
rect 681 40567 747 40584
rect 681 40533 697 40567
rect 731 40533 747 40567
rect 681 40499 747 40533
rect 681 40465 697 40499
rect 731 40465 747 40499
rect 681 40431 747 40465
rect 681 40397 697 40431
rect 731 40397 747 40431
rect 681 40363 747 40397
rect 681 40329 697 40363
rect 731 40329 747 40363
rect 681 40312 747 40329
rect 777 40567 843 40584
rect 777 40533 793 40567
rect 827 40533 843 40567
rect 777 40499 843 40533
rect 777 40465 793 40499
rect 827 40465 843 40499
rect 777 40431 843 40465
rect 777 40397 793 40431
rect 827 40397 843 40431
rect 777 40363 843 40397
rect 777 40329 793 40363
rect 827 40329 843 40363
rect 777 40312 843 40329
rect 873 40567 939 40584
rect 873 40533 889 40567
rect 923 40533 939 40567
rect 873 40499 939 40533
rect 873 40465 889 40499
rect 923 40465 939 40499
rect 873 40431 939 40465
rect 873 40397 889 40431
rect 923 40397 939 40431
rect 873 40363 939 40397
rect 873 40329 889 40363
rect 923 40329 939 40363
rect 873 40312 939 40329
rect 969 40567 1035 40584
rect 969 40533 985 40567
rect 1019 40533 1035 40567
rect 969 40499 1035 40533
rect 969 40465 985 40499
rect 1019 40465 1035 40499
rect 969 40431 1035 40465
rect 969 40397 985 40431
rect 1019 40397 1035 40431
rect 969 40363 1035 40397
rect 969 40329 985 40363
rect 1019 40329 1035 40363
rect 969 40312 1035 40329
rect 1065 40567 1131 40584
rect 1065 40533 1081 40567
rect 1115 40533 1131 40567
rect 1065 40499 1131 40533
rect 1065 40465 1081 40499
rect 1115 40465 1131 40499
rect 1065 40431 1131 40465
rect 1065 40397 1081 40431
rect 1115 40397 1131 40431
rect 1065 40363 1131 40397
rect 1065 40329 1081 40363
rect 1115 40329 1131 40363
rect 1065 40312 1131 40329
rect 1161 40567 1227 40584
rect 1161 40533 1177 40567
rect 1211 40533 1227 40567
rect 1161 40499 1227 40533
rect 1161 40465 1177 40499
rect 1211 40465 1227 40499
rect 1161 40431 1227 40465
rect 1161 40397 1177 40431
rect 1211 40397 1227 40431
rect 1161 40363 1227 40397
rect 1161 40329 1177 40363
rect 1211 40329 1227 40363
rect 1161 40312 1227 40329
rect 1257 40567 1319 40584
rect 1257 40533 1273 40567
rect 1307 40533 1319 40567
rect 1257 40499 1319 40533
rect 1257 40465 1273 40499
rect 1307 40465 1319 40499
rect 1257 40431 1319 40465
rect 1257 40397 1273 40431
rect 1307 40397 1319 40431
rect 1257 40363 1319 40397
rect 1257 40329 1273 40363
rect 1307 40329 1319 40363
rect 1257 40312 1319 40329
rect 2454 40571 2516 40588
rect 2454 40537 2466 40571
rect 2500 40537 2516 40571
rect 2454 40503 2516 40537
rect 2454 40469 2466 40503
rect 2500 40469 2516 40503
rect 2454 40435 2516 40469
rect 2454 40401 2466 40435
rect 2500 40401 2516 40435
rect 2454 40367 2516 40401
rect 2454 40333 2466 40367
rect 2500 40333 2516 40367
rect 2454 40316 2516 40333
rect 2546 40571 2612 40588
rect 2546 40537 2562 40571
rect 2596 40537 2612 40571
rect 2546 40503 2612 40537
rect 2546 40469 2562 40503
rect 2596 40469 2612 40503
rect 2546 40435 2612 40469
rect 2546 40401 2562 40435
rect 2596 40401 2612 40435
rect 2546 40367 2612 40401
rect 2546 40333 2562 40367
rect 2596 40333 2612 40367
rect 2546 40316 2612 40333
rect 2642 40571 2708 40588
rect 2642 40537 2658 40571
rect 2692 40537 2708 40571
rect 2642 40503 2708 40537
rect 2642 40469 2658 40503
rect 2692 40469 2708 40503
rect 2642 40435 2708 40469
rect 2642 40401 2658 40435
rect 2692 40401 2708 40435
rect 2642 40367 2708 40401
rect 2642 40333 2658 40367
rect 2692 40333 2708 40367
rect 2642 40316 2708 40333
rect 2738 40571 2804 40588
rect 2738 40537 2754 40571
rect 2788 40537 2804 40571
rect 2738 40503 2804 40537
rect 2738 40469 2754 40503
rect 2788 40469 2804 40503
rect 2738 40435 2804 40469
rect 2738 40401 2754 40435
rect 2788 40401 2804 40435
rect 2738 40367 2804 40401
rect 2738 40333 2754 40367
rect 2788 40333 2804 40367
rect 2738 40316 2804 40333
rect 2834 40571 2900 40588
rect 2834 40537 2850 40571
rect 2884 40537 2900 40571
rect 2834 40503 2900 40537
rect 2834 40469 2850 40503
rect 2884 40469 2900 40503
rect 2834 40435 2900 40469
rect 2834 40401 2850 40435
rect 2884 40401 2900 40435
rect 2834 40367 2900 40401
rect 2834 40333 2850 40367
rect 2884 40333 2900 40367
rect 2834 40316 2900 40333
rect 2930 40571 2996 40588
rect 2930 40537 2946 40571
rect 2980 40537 2996 40571
rect 2930 40503 2996 40537
rect 2930 40469 2946 40503
rect 2980 40469 2996 40503
rect 2930 40435 2996 40469
rect 2930 40401 2946 40435
rect 2980 40401 2996 40435
rect 2930 40367 2996 40401
rect 2930 40333 2946 40367
rect 2980 40333 2996 40367
rect 2930 40316 2996 40333
rect 3026 40571 3092 40588
rect 3026 40537 3042 40571
rect 3076 40537 3092 40571
rect 3026 40503 3092 40537
rect 3026 40469 3042 40503
rect 3076 40469 3092 40503
rect 3026 40435 3092 40469
rect 3026 40401 3042 40435
rect 3076 40401 3092 40435
rect 3026 40367 3092 40401
rect 3026 40333 3042 40367
rect 3076 40333 3092 40367
rect 3026 40316 3092 40333
rect 3122 40571 3188 40588
rect 3122 40537 3138 40571
rect 3172 40537 3188 40571
rect 3122 40503 3188 40537
rect 3122 40469 3138 40503
rect 3172 40469 3188 40503
rect 3122 40435 3188 40469
rect 3122 40401 3138 40435
rect 3172 40401 3188 40435
rect 3122 40367 3188 40401
rect 3122 40333 3138 40367
rect 3172 40333 3188 40367
rect 3122 40316 3188 40333
rect 3218 40571 3284 40588
rect 3218 40537 3234 40571
rect 3268 40537 3284 40571
rect 3218 40503 3284 40537
rect 3218 40469 3234 40503
rect 3268 40469 3284 40503
rect 3218 40435 3284 40469
rect 3218 40401 3234 40435
rect 3268 40401 3284 40435
rect 3218 40367 3284 40401
rect 3218 40333 3234 40367
rect 3268 40333 3284 40367
rect 3218 40316 3284 40333
rect 3314 40571 3380 40588
rect 3314 40537 3330 40571
rect 3364 40537 3380 40571
rect 3314 40503 3380 40537
rect 3314 40469 3330 40503
rect 3364 40469 3380 40503
rect 3314 40435 3380 40469
rect 3314 40401 3330 40435
rect 3364 40401 3380 40435
rect 3314 40367 3380 40401
rect 3314 40333 3330 40367
rect 3364 40333 3380 40367
rect 3314 40316 3380 40333
rect 3410 40571 3472 40588
rect 3410 40537 3426 40571
rect 3460 40537 3472 40571
rect 3410 40503 3472 40537
rect 3410 40469 3426 40503
rect 3460 40469 3472 40503
rect 3410 40435 3472 40469
rect 3410 40401 3426 40435
rect 3460 40401 3472 40435
rect 3410 40367 3472 40401
rect 3410 40333 3426 40367
rect 3460 40333 3472 40367
rect 3410 40316 3472 40333
rect 3975 40571 4037 40588
rect 3975 40537 3987 40571
rect 4021 40537 4037 40571
rect 3975 40503 4037 40537
rect 3975 40469 3987 40503
rect 4021 40469 4037 40503
rect 3975 40435 4037 40469
rect 3975 40401 3987 40435
rect 4021 40401 4037 40435
rect 3975 40367 4037 40401
rect 3975 40333 3987 40367
rect 4021 40333 4037 40367
rect 3975 40316 4037 40333
rect 4067 40571 4133 40588
rect 4067 40537 4083 40571
rect 4117 40537 4133 40571
rect 4067 40503 4133 40537
rect 4067 40469 4083 40503
rect 4117 40469 4133 40503
rect 4067 40435 4133 40469
rect 4067 40401 4083 40435
rect 4117 40401 4133 40435
rect 4067 40367 4133 40401
rect 4067 40333 4083 40367
rect 4117 40333 4133 40367
rect 4067 40316 4133 40333
rect 4163 40571 4229 40588
rect 4163 40537 4179 40571
rect 4213 40537 4229 40571
rect 4163 40503 4229 40537
rect 4163 40469 4179 40503
rect 4213 40469 4229 40503
rect 4163 40435 4229 40469
rect 4163 40401 4179 40435
rect 4213 40401 4229 40435
rect 4163 40367 4229 40401
rect 4163 40333 4179 40367
rect 4213 40333 4229 40367
rect 4163 40316 4229 40333
rect 4259 40571 4325 40588
rect 4259 40537 4275 40571
rect 4309 40537 4325 40571
rect 4259 40503 4325 40537
rect 4259 40469 4275 40503
rect 4309 40469 4325 40503
rect 4259 40435 4325 40469
rect 4259 40401 4275 40435
rect 4309 40401 4325 40435
rect 4259 40367 4325 40401
rect 4259 40333 4275 40367
rect 4309 40333 4325 40367
rect 4259 40316 4325 40333
rect 4355 40571 4421 40588
rect 4355 40537 4371 40571
rect 4405 40537 4421 40571
rect 4355 40503 4421 40537
rect 4355 40469 4371 40503
rect 4405 40469 4421 40503
rect 4355 40435 4421 40469
rect 4355 40401 4371 40435
rect 4405 40401 4421 40435
rect 4355 40367 4421 40401
rect 4355 40333 4371 40367
rect 4405 40333 4421 40367
rect 4355 40316 4421 40333
rect 4451 40571 4517 40588
rect 4451 40537 4467 40571
rect 4501 40537 4517 40571
rect 4451 40503 4517 40537
rect 4451 40469 4467 40503
rect 4501 40469 4517 40503
rect 4451 40435 4517 40469
rect 4451 40401 4467 40435
rect 4501 40401 4517 40435
rect 4451 40367 4517 40401
rect 4451 40333 4467 40367
rect 4501 40333 4517 40367
rect 4451 40316 4517 40333
rect 4547 40571 4613 40588
rect 4547 40537 4563 40571
rect 4597 40537 4613 40571
rect 4547 40503 4613 40537
rect 4547 40469 4563 40503
rect 4597 40469 4613 40503
rect 4547 40435 4613 40469
rect 4547 40401 4563 40435
rect 4597 40401 4613 40435
rect 4547 40367 4613 40401
rect 4547 40333 4563 40367
rect 4597 40333 4613 40367
rect 4547 40316 4613 40333
rect 4643 40571 4709 40588
rect 4643 40537 4659 40571
rect 4693 40537 4709 40571
rect 4643 40503 4709 40537
rect 4643 40469 4659 40503
rect 4693 40469 4709 40503
rect 4643 40435 4709 40469
rect 4643 40401 4659 40435
rect 4693 40401 4709 40435
rect 4643 40367 4709 40401
rect 4643 40333 4659 40367
rect 4693 40333 4709 40367
rect 4643 40316 4709 40333
rect 4739 40571 4805 40588
rect 4739 40537 4755 40571
rect 4789 40537 4805 40571
rect 4739 40503 4805 40537
rect 4739 40469 4755 40503
rect 4789 40469 4805 40503
rect 4739 40435 4805 40469
rect 4739 40401 4755 40435
rect 4789 40401 4805 40435
rect 4739 40367 4805 40401
rect 4739 40333 4755 40367
rect 4789 40333 4805 40367
rect 4739 40316 4805 40333
rect 4835 40571 4901 40588
rect 4835 40537 4851 40571
rect 4885 40537 4901 40571
rect 4835 40503 4901 40537
rect 4835 40469 4851 40503
rect 4885 40469 4901 40503
rect 4835 40435 4901 40469
rect 4835 40401 4851 40435
rect 4885 40401 4901 40435
rect 4835 40367 4901 40401
rect 4835 40333 4851 40367
rect 4885 40333 4901 40367
rect 4835 40316 4901 40333
rect 4931 40571 4993 40588
rect 4931 40537 4947 40571
rect 4981 40537 4993 40571
rect 4931 40503 4993 40537
rect 4931 40469 4947 40503
rect 4981 40469 4993 40503
rect 4931 40435 4993 40469
rect 4931 40401 4947 40435
rect 4981 40401 4993 40435
rect 4931 40367 4993 40401
rect 4931 40333 4947 40367
rect 4981 40333 4993 40367
rect 4931 40316 4993 40333
rect 5348 40363 5400 40375
rect 5348 40329 5356 40363
rect 5390 40329 5400 40363
rect 5348 40295 5400 40329
rect 5348 40261 5356 40295
rect 5390 40261 5400 40295
rect 5348 40227 5400 40261
rect 5348 40193 5356 40227
rect 5390 40193 5400 40227
rect 5348 40175 5400 40193
rect 5430 40363 5482 40375
rect 5430 40329 5440 40363
rect 5474 40329 5482 40363
rect 5430 40295 5482 40329
rect 5430 40261 5440 40295
rect 5474 40261 5482 40295
rect 5430 40227 5482 40261
rect 5430 40193 5440 40227
rect 5474 40193 5482 40227
rect 5430 40175 5482 40193
rect 301 39280 363 39297
rect 301 39246 313 39280
rect 347 39246 363 39280
rect 301 39212 363 39246
rect 301 39178 313 39212
rect 347 39178 363 39212
rect 301 39144 363 39178
rect 301 39110 313 39144
rect 347 39110 363 39144
rect 301 39076 363 39110
rect 301 39042 313 39076
rect 347 39042 363 39076
rect 301 39025 363 39042
rect 393 39280 459 39297
rect 393 39246 409 39280
rect 443 39246 459 39280
rect 393 39212 459 39246
rect 393 39178 409 39212
rect 443 39178 459 39212
rect 393 39144 459 39178
rect 393 39110 409 39144
rect 443 39110 459 39144
rect 393 39076 459 39110
rect 393 39042 409 39076
rect 443 39042 459 39076
rect 393 39025 459 39042
rect 489 39280 555 39297
rect 489 39246 505 39280
rect 539 39246 555 39280
rect 489 39212 555 39246
rect 489 39178 505 39212
rect 539 39178 555 39212
rect 489 39144 555 39178
rect 489 39110 505 39144
rect 539 39110 555 39144
rect 489 39076 555 39110
rect 489 39042 505 39076
rect 539 39042 555 39076
rect 489 39025 555 39042
rect 585 39280 651 39297
rect 585 39246 601 39280
rect 635 39246 651 39280
rect 585 39212 651 39246
rect 585 39178 601 39212
rect 635 39178 651 39212
rect 585 39144 651 39178
rect 585 39110 601 39144
rect 635 39110 651 39144
rect 585 39076 651 39110
rect 585 39042 601 39076
rect 635 39042 651 39076
rect 585 39025 651 39042
rect 681 39280 747 39297
rect 681 39246 697 39280
rect 731 39246 747 39280
rect 681 39212 747 39246
rect 681 39178 697 39212
rect 731 39178 747 39212
rect 681 39144 747 39178
rect 681 39110 697 39144
rect 731 39110 747 39144
rect 681 39076 747 39110
rect 681 39042 697 39076
rect 731 39042 747 39076
rect 681 39025 747 39042
rect 777 39280 843 39297
rect 777 39246 793 39280
rect 827 39246 843 39280
rect 777 39212 843 39246
rect 777 39178 793 39212
rect 827 39178 843 39212
rect 777 39144 843 39178
rect 777 39110 793 39144
rect 827 39110 843 39144
rect 777 39076 843 39110
rect 777 39042 793 39076
rect 827 39042 843 39076
rect 777 39025 843 39042
rect 873 39280 939 39297
rect 873 39246 889 39280
rect 923 39246 939 39280
rect 873 39212 939 39246
rect 873 39178 889 39212
rect 923 39178 939 39212
rect 873 39144 939 39178
rect 873 39110 889 39144
rect 923 39110 939 39144
rect 873 39076 939 39110
rect 873 39042 889 39076
rect 923 39042 939 39076
rect 873 39025 939 39042
rect 969 39280 1035 39297
rect 969 39246 985 39280
rect 1019 39246 1035 39280
rect 969 39212 1035 39246
rect 969 39178 985 39212
rect 1019 39178 1035 39212
rect 969 39144 1035 39178
rect 969 39110 985 39144
rect 1019 39110 1035 39144
rect 969 39076 1035 39110
rect 969 39042 985 39076
rect 1019 39042 1035 39076
rect 969 39025 1035 39042
rect 1065 39280 1131 39297
rect 1065 39246 1081 39280
rect 1115 39246 1131 39280
rect 1065 39212 1131 39246
rect 1065 39178 1081 39212
rect 1115 39178 1131 39212
rect 1065 39144 1131 39178
rect 1065 39110 1081 39144
rect 1115 39110 1131 39144
rect 1065 39076 1131 39110
rect 1065 39042 1081 39076
rect 1115 39042 1131 39076
rect 1065 39025 1131 39042
rect 1161 39280 1227 39297
rect 1161 39246 1177 39280
rect 1211 39246 1227 39280
rect 1161 39212 1227 39246
rect 1161 39178 1177 39212
rect 1211 39178 1227 39212
rect 1161 39144 1227 39178
rect 1161 39110 1177 39144
rect 1211 39110 1227 39144
rect 1161 39076 1227 39110
rect 1161 39042 1177 39076
rect 1211 39042 1227 39076
rect 1161 39025 1227 39042
rect 1257 39280 1319 39297
rect 1257 39246 1273 39280
rect 1307 39246 1319 39280
rect 1257 39212 1319 39246
rect 1257 39178 1273 39212
rect 1307 39178 1319 39212
rect 1257 39144 1319 39178
rect 1257 39110 1273 39144
rect 1307 39110 1319 39144
rect 1257 39076 1319 39110
rect 1257 39042 1273 39076
rect 1307 39042 1319 39076
rect 1257 39025 1319 39042
rect 2454 39284 2516 39301
rect 2454 39250 2466 39284
rect 2500 39250 2516 39284
rect 2454 39216 2516 39250
rect 2454 39182 2466 39216
rect 2500 39182 2516 39216
rect 2454 39148 2516 39182
rect 2454 39114 2466 39148
rect 2500 39114 2516 39148
rect 2454 39080 2516 39114
rect 2454 39046 2466 39080
rect 2500 39046 2516 39080
rect 2454 39029 2516 39046
rect 2546 39284 2612 39301
rect 2546 39250 2562 39284
rect 2596 39250 2612 39284
rect 2546 39216 2612 39250
rect 2546 39182 2562 39216
rect 2596 39182 2612 39216
rect 2546 39148 2612 39182
rect 2546 39114 2562 39148
rect 2596 39114 2612 39148
rect 2546 39080 2612 39114
rect 2546 39046 2562 39080
rect 2596 39046 2612 39080
rect 2546 39029 2612 39046
rect 2642 39284 2708 39301
rect 2642 39250 2658 39284
rect 2692 39250 2708 39284
rect 2642 39216 2708 39250
rect 2642 39182 2658 39216
rect 2692 39182 2708 39216
rect 2642 39148 2708 39182
rect 2642 39114 2658 39148
rect 2692 39114 2708 39148
rect 2642 39080 2708 39114
rect 2642 39046 2658 39080
rect 2692 39046 2708 39080
rect 2642 39029 2708 39046
rect 2738 39284 2804 39301
rect 2738 39250 2754 39284
rect 2788 39250 2804 39284
rect 2738 39216 2804 39250
rect 2738 39182 2754 39216
rect 2788 39182 2804 39216
rect 2738 39148 2804 39182
rect 2738 39114 2754 39148
rect 2788 39114 2804 39148
rect 2738 39080 2804 39114
rect 2738 39046 2754 39080
rect 2788 39046 2804 39080
rect 2738 39029 2804 39046
rect 2834 39284 2900 39301
rect 2834 39250 2850 39284
rect 2884 39250 2900 39284
rect 2834 39216 2900 39250
rect 2834 39182 2850 39216
rect 2884 39182 2900 39216
rect 2834 39148 2900 39182
rect 2834 39114 2850 39148
rect 2884 39114 2900 39148
rect 2834 39080 2900 39114
rect 2834 39046 2850 39080
rect 2884 39046 2900 39080
rect 2834 39029 2900 39046
rect 2930 39284 2996 39301
rect 2930 39250 2946 39284
rect 2980 39250 2996 39284
rect 2930 39216 2996 39250
rect 2930 39182 2946 39216
rect 2980 39182 2996 39216
rect 2930 39148 2996 39182
rect 2930 39114 2946 39148
rect 2980 39114 2996 39148
rect 2930 39080 2996 39114
rect 2930 39046 2946 39080
rect 2980 39046 2996 39080
rect 2930 39029 2996 39046
rect 3026 39284 3092 39301
rect 3026 39250 3042 39284
rect 3076 39250 3092 39284
rect 3026 39216 3092 39250
rect 3026 39182 3042 39216
rect 3076 39182 3092 39216
rect 3026 39148 3092 39182
rect 3026 39114 3042 39148
rect 3076 39114 3092 39148
rect 3026 39080 3092 39114
rect 3026 39046 3042 39080
rect 3076 39046 3092 39080
rect 3026 39029 3092 39046
rect 3122 39284 3188 39301
rect 3122 39250 3138 39284
rect 3172 39250 3188 39284
rect 3122 39216 3188 39250
rect 3122 39182 3138 39216
rect 3172 39182 3188 39216
rect 3122 39148 3188 39182
rect 3122 39114 3138 39148
rect 3172 39114 3188 39148
rect 3122 39080 3188 39114
rect 3122 39046 3138 39080
rect 3172 39046 3188 39080
rect 3122 39029 3188 39046
rect 3218 39284 3284 39301
rect 3218 39250 3234 39284
rect 3268 39250 3284 39284
rect 3218 39216 3284 39250
rect 3218 39182 3234 39216
rect 3268 39182 3284 39216
rect 3218 39148 3284 39182
rect 3218 39114 3234 39148
rect 3268 39114 3284 39148
rect 3218 39080 3284 39114
rect 3218 39046 3234 39080
rect 3268 39046 3284 39080
rect 3218 39029 3284 39046
rect 3314 39284 3380 39301
rect 3314 39250 3330 39284
rect 3364 39250 3380 39284
rect 3314 39216 3380 39250
rect 3314 39182 3330 39216
rect 3364 39182 3380 39216
rect 3314 39148 3380 39182
rect 3314 39114 3330 39148
rect 3364 39114 3380 39148
rect 3314 39080 3380 39114
rect 3314 39046 3330 39080
rect 3364 39046 3380 39080
rect 3314 39029 3380 39046
rect 3410 39284 3472 39301
rect 3410 39250 3426 39284
rect 3460 39250 3472 39284
rect 3410 39216 3472 39250
rect 3410 39182 3426 39216
rect 3460 39182 3472 39216
rect 3410 39148 3472 39182
rect 3410 39114 3426 39148
rect 3460 39114 3472 39148
rect 3410 39080 3472 39114
rect 3410 39046 3426 39080
rect 3460 39046 3472 39080
rect 3410 39029 3472 39046
rect 3975 39284 4037 39301
rect 3975 39250 3987 39284
rect 4021 39250 4037 39284
rect 3975 39216 4037 39250
rect 3975 39182 3987 39216
rect 4021 39182 4037 39216
rect 3975 39148 4037 39182
rect 3975 39114 3987 39148
rect 4021 39114 4037 39148
rect 3975 39080 4037 39114
rect 3975 39046 3987 39080
rect 4021 39046 4037 39080
rect 3975 39029 4037 39046
rect 4067 39284 4133 39301
rect 4067 39250 4083 39284
rect 4117 39250 4133 39284
rect 4067 39216 4133 39250
rect 4067 39182 4083 39216
rect 4117 39182 4133 39216
rect 4067 39148 4133 39182
rect 4067 39114 4083 39148
rect 4117 39114 4133 39148
rect 4067 39080 4133 39114
rect 4067 39046 4083 39080
rect 4117 39046 4133 39080
rect 4067 39029 4133 39046
rect 4163 39284 4229 39301
rect 4163 39250 4179 39284
rect 4213 39250 4229 39284
rect 4163 39216 4229 39250
rect 4163 39182 4179 39216
rect 4213 39182 4229 39216
rect 4163 39148 4229 39182
rect 4163 39114 4179 39148
rect 4213 39114 4229 39148
rect 4163 39080 4229 39114
rect 4163 39046 4179 39080
rect 4213 39046 4229 39080
rect 4163 39029 4229 39046
rect 4259 39284 4325 39301
rect 4259 39250 4275 39284
rect 4309 39250 4325 39284
rect 4259 39216 4325 39250
rect 4259 39182 4275 39216
rect 4309 39182 4325 39216
rect 4259 39148 4325 39182
rect 4259 39114 4275 39148
rect 4309 39114 4325 39148
rect 4259 39080 4325 39114
rect 4259 39046 4275 39080
rect 4309 39046 4325 39080
rect 4259 39029 4325 39046
rect 4355 39284 4421 39301
rect 4355 39250 4371 39284
rect 4405 39250 4421 39284
rect 4355 39216 4421 39250
rect 4355 39182 4371 39216
rect 4405 39182 4421 39216
rect 4355 39148 4421 39182
rect 4355 39114 4371 39148
rect 4405 39114 4421 39148
rect 4355 39080 4421 39114
rect 4355 39046 4371 39080
rect 4405 39046 4421 39080
rect 4355 39029 4421 39046
rect 4451 39284 4517 39301
rect 4451 39250 4467 39284
rect 4501 39250 4517 39284
rect 4451 39216 4517 39250
rect 4451 39182 4467 39216
rect 4501 39182 4517 39216
rect 4451 39148 4517 39182
rect 4451 39114 4467 39148
rect 4501 39114 4517 39148
rect 4451 39080 4517 39114
rect 4451 39046 4467 39080
rect 4501 39046 4517 39080
rect 4451 39029 4517 39046
rect 4547 39284 4613 39301
rect 4547 39250 4563 39284
rect 4597 39250 4613 39284
rect 4547 39216 4613 39250
rect 4547 39182 4563 39216
rect 4597 39182 4613 39216
rect 4547 39148 4613 39182
rect 4547 39114 4563 39148
rect 4597 39114 4613 39148
rect 4547 39080 4613 39114
rect 4547 39046 4563 39080
rect 4597 39046 4613 39080
rect 4547 39029 4613 39046
rect 4643 39284 4709 39301
rect 4643 39250 4659 39284
rect 4693 39250 4709 39284
rect 4643 39216 4709 39250
rect 4643 39182 4659 39216
rect 4693 39182 4709 39216
rect 4643 39148 4709 39182
rect 4643 39114 4659 39148
rect 4693 39114 4709 39148
rect 4643 39080 4709 39114
rect 4643 39046 4659 39080
rect 4693 39046 4709 39080
rect 4643 39029 4709 39046
rect 4739 39284 4805 39301
rect 4739 39250 4755 39284
rect 4789 39250 4805 39284
rect 4739 39216 4805 39250
rect 4739 39182 4755 39216
rect 4789 39182 4805 39216
rect 4739 39148 4805 39182
rect 4739 39114 4755 39148
rect 4789 39114 4805 39148
rect 4739 39080 4805 39114
rect 4739 39046 4755 39080
rect 4789 39046 4805 39080
rect 4739 39029 4805 39046
rect 4835 39284 4901 39301
rect 4835 39250 4851 39284
rect 4885 39250 4901 39284
rect 4835 39216 4901 39250
rect 4835 39182 4851 39216
rect 4885 39182 4901 39216
rect 4835 39148 4901 39182
rect 4835 39114 4851 39148
rect 4885 39114 4901 39148
rect 4835 39080 4901 39114
rect 4835 39046 4851 39080
rect 4885 39046 4901 39080
rect 4835 39029 4901 39046
rect 4931 39284 4993 39301
rect 4931 39250 4947 39284
rect 4981 39250 4993 39284
rect 4931 39216 4993 39250
rect 4931 39182 4947 39216
rect 4981 39182 4993 39216
rect 4931 39148 4993 39182
rect 4931 39114 4947 39148
rect 4981 39114 4993 39148
rect 4931 39080 4993 39114
rect 4931 39046 4947 39080
rect 4981 39046 4993 39080
rect 4931 39029 4993 39046
rect 5348 39076 5400 39088
rect 5348 39042 5356 39076
rect 5390 39042 5400 39076
rect 5348 39008 5400 39042
rect 5348 38974 5356 39008
rect 5390 38974 5400 39008
rect 5348 38940 5400 38974
rect 5348 38906 5356 38940
rect 5390 38906 5400 38940
rect 5348 38888 5400 38906
rect 5430 39076 5482 39088
rect 5430 39042 5440 39076
rect 5474 39042 5482 39076
rect 5430 39008 5482 39042
rect 5430 38974 5440 39008
rect 5474 38974 5482 39008
rect 5430 38940 5482 38974
rect 5430 38906 5440 38940
rect 5474 38906 5482 38940
rect 5430 38888 5482 38906
rect 301 37993 363 38010
rect 301 37959 313 37993
rect 347 37959 363 37993
rect 301 37925 363 37959
rect 301 37891 313 37925
rect 347 37891 363 37925
rect 301 37857 363 37891
rect 301 37823 313 37857
rect 347 37823 363 37857
rect 301 37789 363 37823
rect 301 37755 313 37789
rect 347 37755 363 37789
rect 301 37738 363 37755
rect 393 37993 459 38010
rect 393 37959 409 37993
rect 443 37959 459 37993
rect 393 37925 459 37959
rect 393 37891 409 37925
rect 443 37891 459 37925
rect 393 37857 459 37891
rect 393 37823 409 37857
rect 443 37823 459 37857
rect 393 37789 459 37823
rect 393 37755 409 37789
rect 443 37755 459 37789
rect 393 37738 459 37755
rect 489 37993 555 38010
rect 489 37959 505 37993
rect 539 37959 555 37993
rect 489 37925 555 37959
rect 489 37891 505 37925
rect 539 37891 555 37925
rect 489 37857 555 37891
rect 489 37823 505 37857
rect 539 37823 555 37857
rect 489 37789 555 37823
rect 489 37755 505 37789
rect 539 37755 555 37789
rect 489 37738 555 37755
rect 585 37993 651 38010
rect 585 37959 601 37993
rect 635 37959 651 37993
rect 585 37925 651 37959
rect 585 37891 601 37925
rect 635 37891 651 37925
rect 585 37857 651 37891
rect 585 37823 601 37857
rect 635 37823 651 37857
rect 585 37789 651 37823
rect 585 37755 601 37789
rect 635 37755 651 37789
rect 585 37738 651 37755
rect 681 37993 747 38010
rect 681 37959 697 37993
rect 731 37959 747 37993
rect 681 37925 747 37959
rect 681 37891 697 37925
rect 731 37891 747 37925
rect 681 37857 747 37891
rect 681 37823 697 37857
rect 731 37823 747 37857
rect 681 37789 747 37823
rect 681 37755 697 37789
rect 731 37755 747 37789
rect 681 37738 747 37755
rect 777 37993 843 38010
rect 777 37959 793 37993
rect 827 37959 843 37993
rect 777 37925 843 37959
rect 777 37891 793 37925
rect 827 37891 843 37925
rect 777 37857 843 37891
rect 777 37823 793 37857
rect 827 37823 843 37857
rect 777 37789 843 37823
rect 777 37755 793 37789
rect 827 37755 843 37789
rect 777 37738 843 37755
rect 873 37993 939 38010
rect 873 37959 889 37993
rect 923 37959 939 37993
rect 873 37925 939 37959
rect 873 37891 889 37925
rect 923 37891 939 37925
rect 873 37857 939 37891
rect 873 37823 889 37857
rect 923 37823 939 37857
rect 873 37789 939 37823
rect 873 37755 889 37789
rect 923 37755 939 37789
rect 873 37738 939 37755
rect 969 37993 1035 38010
rect 969 37959 985 37993
rect 1019 37959 1035 37993
rect 969 37925 1035 37959
rect 969 37891 985 37925
rect 1019 37891 1035 37925
rect 969 37857 1035 37891
rect 969 37823 985 37857
rect 1019 37823 1035 37857
rect 969 37789 1035 37823
rect 969 37755 985 37789
rect 1019 37755 1035 37789
rect 969 37738 1035 37755
rect 1065 37993 1131 38010
rect 1065 37959 1081 37993
rect 1115 37959 1131 37993
rect 1065 37925 1131 37959
rect 1065 37891 1081 37925
rect 1115 37891 1131 37925
rect 1065 37857 1131 37891
rect 1065 37823 1081 37857
rect 1115 37823 1131 37857
rect 1065 37789 1131 37823
rect 1065 37755 1081 37789
rect 1115 37755 1131 37789
rect 1065 37738 1131 37755
rect 1161 37993 1227 38010
rect 1161 37959 1177 37993
rect 1211 37959 1227 37993
rect 1161 37925 1227 37959
rect 1161 37891 1177 37925
rect 1211 37891 1227 37925
rect 1161 37857 1227 37891
rect 1161 37823 1177 37857
rect 1211 37823 1227 37857
rect 1161 37789 1227 37823
rect 1161 37755 1177 37789
rect 1211 37755 1227 37789
rect 1161 37738 1227 37755
rect 1257 37993 1319 38010
rect 1257 37959 1273 37993
rect 1307 37959 1319 37993
rect 1257 37925 1319 37959
rect 1257 37891 1273 37925
rect 1307 37891 1319 37925
rect 1257 37857 1319 37891
rect 1257 37823 1273 37857
rect 1307 37823 1319 37857
rect 1257 37789 1319 37823
rect 1257 37755 1273 37789
rect 1307 37755 1319 37789
rect 1257 37738 1319 37755
rect 2454 37997 2516 38014
rect 2454 37963 2466 37997
rect 2500 37963 2516 37997
rect 2454 37929 2516 37963
rect 2454 37895 2466 37929
rect 2500 37895 2516 37929
rect 2454 37861 2516 37895
rect 2454 37827 2466 37861
rect 2500 37827 2516 37861
rect 2454 37793 2516 37827
rect 2454 37759 2466 37793
rect 2500 37759 2516 37793
rect 2454 37742 2516 37759
rect 2546 37997 2612 38014
rect 2546 37963 2562 37997
rect 2596 37963 2612 37997
rect 2546 37929 2612 37963
rect 2546 37895 2562 37929
rect 2596 37895 2612 37929
rect 2546 37861 2612 37895
rect 2546 37827 2562 37861
rect 2596 37827 2612 37861
rect 2546 37793 2612 37827
rect 2546 37759 2562 37793
rect 2596 37759 2612 37793
rect 2546 37742 2612 37759
rect 2642 37997 2708 38014
rect 2642 37963 2658 37997
rect 2692 37963 2708 37997
rect 2642 37929 2708 37963
rect 2642 37895 2658 37929
rect 2692 37895 2708 37929
rect 2642 37861 2708 37895
rect 2642 37827 2658 37861
rect 2692 37827 2708 37861
rect 2642 37793 2708 37827
rect 2642 37759 2658 37793
rect 2692 37759 2708 37793
rect 2642 37742 2708 37759
rect 2738 37997 2804 38014
rect 2738 37963 2754 37997
rect 2788 37963 2804 37997
rect 2738 37929 2804 37963
rect 2738 37895 2754 37929
rect 2788 37895 2804 37929
rect 2738 37861 2804 37895
rect 2738 37827 2754 37861
rect 2788 37827 2804 37861
rect 2738 37793 2804 37827
rect 2738 37759 2754 37793
rect 2788 37759 2804 37793
rect 2738 37742 2804 37759
rect 2834 37997 2900 38014
rect 2834 37963 2850 37997
rect 2884 37963 2900 37997
rect 2834 37929 2900 37963
rect 2834 37895 2850 37929
rect 2884 37895 2900 37929
rect 2834 37861 2900 37895
rect 2834 37827 2850 37861
rect 2884 37827 2900 37861
rect 2834 37793 2900 37827
rect 2834 37759 2850 37793
rect 2884 37759 2900 37793
rect 2834 37742 2900 37759
rect 2930 37997 2996 38014
rect 2930 37963 2946 37997
rect 2980 37963 2996 37997
rect 2930 37929 2996 37963
rect 2930 37895 2946 37929
rect 2980 37895 2996 37929
rect 2930 37861 2996 37895
rect 2930 37827 2946 37861
rect 2980 37827 2996 37861
rect 2930 37793 2996 37827
rect 2930 37759 2946 37793
rect 2980 37759 2996 37793
rect 2930 37742 2996 37759
rect 3026 37997 3092 38014
rect 3026 37963 3042 37997
rect 3076 37963 3092 37997
rect 3026 37929 3092 37963
rect 3026 37895 3042 37929
rect 3076 37895 3092 37929
rect 3026 37861 3092 37895
rect 3026 37827 3042 37861
rect 3076 37827 3092 37861
rect 3026 37793 3092 37827
rect 3026 37759 3042 37793
rect 3076 37759 3092 37793
rect 3026 37742 3092 37759
rect 3122 37997 3188 38014
rect 3122 37963 3138 37997
rect 3172 37963 3188 37997
rect 3122 37929 3188 37963
rect 3122 37895 3138 37929
rect 3172 37895 3188 37929
rect 3122 37861 3188 37895
rect 3122 37827 3138 37861
rect 3172 37827 3188 37861
rect 3122 37793 3188 37827
rect 3122 37759 3138 37793
rect 3172 37759 3188 37793
rect 3122 37742 3188 37759
rect 3218 37997 3284 38014
rect 3218 37963 3234 37997
rect 3268 37963 3284 37997
rect 3218 37929 3284 37963
rect 3218 37895 3234 37929
rect 3268 37895 3284 37929
rect 3218 37861 3284 37895
rect 3218 37827 3234 37861
rect 3268 37827 3284 37861
rect 3218 37793 3284 37827
rect 3218 37759 3234 37793
rect 3268 37759 3284 37793
rect 3218 37742 3284 37759
rect 3314 37997 3380 38014
rect 3314 37963 3330 37997
rect 3364 37963 3380 37997
rect 3314 37929 3380 37963
rect 3314 37895 3330 37929
rect 3364 37895 3380 37929
rect 3314 37861 3380 37895
rect 3314 37827 3330 37861
rect 3364 37827 3380 37861
rect 3314 37793 3380 37827
rect 3314 37759 3330 37793
rect 3364 37759 3380 37793
rect 3314 37742 3380 37759
rect 3410 37997 3472 38014
rect 3410 37963 3426 37997
rect 3460 37963 3472 37997
rect 3410 37929 3472 37963
rect 3410 37895 3426 37929
rect 3460 37895 3472 37929
rect 3410 37861 3472 37895
rect 3410 37827 3426 37861
rect 3460 37827 3472 37861
rect 3410 37793 3472 37827
rect 3410 37759 3426 37793
rect 3460 37759 3472 37793
rect 3410 37742 3472 37759
rect 3975 37997 4037 38014
rect 3975 37963 3987 37997
rect 4021 37963 4037 37997
rect 3975 37929 4037 37963
rect 3975 37895 3987 37929
rect 4021 37895 4037 37929
rect 3975 37861 4037 37895
rect 3975 37827 3987 37861
rect 4021 37827 4037 37861
rect 3975 37793 4037 37827
rect 3975 37759 3987 37793
rect 4021 37759 4037 37793
rect 3975 37742 4037 37759
rect 4067 37997 4133 38014
rect 4067 37963 4083 37997
rect 4117 37963 4133 37997
rect 4067 37929 4133 37963
rect 4067 37895 4083 37929
rect 4117 37895 4133 37929
rect 4067 37861 4133 37895
rect 4067 37827 4083 37861
rect 4117 37827 4133 37861
rect 4067 37793 4133 37827
rect 4067 37759 4083 37793
rect 4117 37759 4133 37793
rect 4067 37742 4133 37759
rect 4163 37997 4229 38014
rect 4163 37963 4179 37997
rect 4213 37963 4229 37997
rect 4163 37929 4229 37963
rect 4163 37895 4179 37929
rect 4213 37895 4229 37929
rect 4163 37861 4229 37895
rect 4163 37827 4179 37861
rect 4213 37827 4229 37861
rect 4163 37793 4229 37827
rect 4163 37759 4179 37793
rect 4213 37759 4229 37793
rect 4163 37742 4229 37759
rect 4259 37997 4325 38014
rect 4259 37963 4275 37997
rect 4309 37963 4325 37997
rect 4259 37929 4325 37963
rect 4259 37895 4275 37929
rect 4309 37895 4325 37929
rect 4259 37861 4325 37895
rect 4259 37827 4275 37861
rect 4309 37827 4325 37861
rect 4259 37793 4325 37827
rect 4259 37759 4275 37793
rect 4309 37759 4325 37793
rect 4259 37742 4325 37759
rect 4355 37997 4421 38014
rect 4355 37963 4371 37997
rect 4405 37963 4421 37997
rect 4355 37929 4421 37963
rect 4355 37895 4371 37929
rect 4405 37895 4421 37929
rect 4355 37861 4421 37895
rect 4355 37827 4371 37861
rect 4405 37827 4421 37861
rect 4355 37793 4421 37827
rect 4355 37759 4371 37793
rect 4405 37759 4421 37793
rect 4355 37742 4421 37759
rect 4451 37997 4517 38014
rect 4451 37963 4467 37997
rect 4501 37963 4517 37997
rect 4451 37929 4517 37963
rect 4451 37895 4467 37929
rect 4501 37895 4517 37929
rect 4451 37861 4517 37895
rect 4451 37827 4467 37861
rect 4501 37827 4517 37861
rect 4451 37793 4517 37827
rect 4451 37759 4467 37793
rect 4501 37759 4517 37793
rect 4451 37742 4517 37759
rect 4547 37997 4613 38014
rect 4547 37963 4563 37997
rect 4597 37963 4613 37997
rect 4547 37929 4613 37963
rect 4547 37895 4563 37929
rect 4597 37895 4613 37929
rect 4547 37861 4613 37895
rect 4547 37827 4563 37861
rect 4597 37827 4613 37861
rect 4547 37793 4613 37827
rect 4547 37759 4563 37793
rect 4597 37759 4613 37793
rect 4547 37742 4613 37759
rect 4643 37997 4709 38014
rect 4643 37963 4659 37997
rect 4693 37963 4709 37997
rect 4643 37929 4709 37963
rect 4643 37895 4659 37929
rect 4693 37895 4709 37929
rect 4643 37861 4709 37895
rect 4643 37827 4659 37861
rect 4693 37827 4709 37861
rect 4643 37793 4709 37827
rect 4643 37759 4659 37793
rect 4693 37759 4709 37793
rect 4643 37742 4709 37759
rect 4739 37997 4805 38014
rect 4739 37963 4755 37997
rect 4789 37963 4805 37997
rect 4739 37929 4805 37963
rect 4739 37895 4755 37929
rect 4789 37895 4805 37929
rect 4739 37861 4805 37895
rect 4739 37827 4755 37861
rect 4789 37827 4805 37861
rect 4739 37793 4805 37827
rect 4739 37759 4755 37793
rect 4789 37759 4805 37793
rect 4739 37742 4805 37759
rect 4835 37997 4901 38014
rect 4835 37963 4851 37997
rect 4885 37963 4901 37997
rect 4835 37929 4901 37963
rect 4835 37895 4851 37929
rect 4885 37895 4901 37929
rect 4835 37861 4901 37895
rect 4835 37827 4851 37861
rect 4885 37827 4901 37861
rect 4835 37793 4901 37827
rect 4835 37759 4851 37793
rect 4885 37759 4901 37793
rect 4835 37742 4901 37759
rect 4931 37997 4993 38014
rect 4931 37963 4947 37997
rect 4981 37963 4993 37997
rect 4931 37929 4993 37963
rect 4931 37895 4947 37929
rect 4981 37895 4993 37929
rect 4931 37861 4993 37895
rect 4931 37827 4947 37861
rect 4981 37827 4993 37861
rect 4931 37793 4993 37827
rect 4931 37759 4947 37793
rect 4981 37759 4993 37793
rect 4931 37742 4993 37759
rect 5348 37789 5400 37801
rect 5348 37755 5356 37789
rect 5390 37755 5400 37789
rect 5348 37721 5400 37755
rect 5348 37687 5356 37721
rect 5390 37687 5400 37721
rect 5348 37653 5400 37687
rect 5348 37619 5356 37653
rect 5390 37619 5400 37653
rect 5348 37601 5400 37619
rect 5430 37789 5482 37801
rect 5430 37755 5440 37789
rect 5474 37755 5482 37789
rect 5430 37721 5482 37755
rect 5430 37687 5440 37721
rect 5474 37687 5482 37721
rect 5430 37653 5482 37687
rect 5430 37619 5440 37653
rect 5474 37619 5482 37653
rect 5430 37601 5482 37619
rect 301 36706 363 36723
rect 301 36672 313 36706
rect 347 36672 363 36706
rect 301 36638 363 36672
rect 301 36604 313 36638
rect 347 36604 363 36638
rect 301 36570 363 36604
rect 301 36536 313 36570
rect 347 36536 363 36570
rect 301 36502 363 36536
rect 301 36468 313 36502
rect 347 36468 363 36502
rect 301 36451 363 36468
rect 393 36706 459 36723
rect 393 36672 409 36706
rect 443 36672 459 36706
rect 393 36638 459 36672
rect 393 36604 409 36638
rect 443 36604 459 36638
rect 393 36570 459 36604
rect 393 36536 409 36570
rect 443 36536 459 36570
rect 393 36502 459 36536
rect 393 36468 409 36502
rect 443 36468 459 36502
rect 393 36451 459 36468
rect 489 36706 555 36723
rect 489 36672 505 36706
rect 539 36672 555 36706
rect 489 36638 555 36672
rect 489 36604 505 36638
rect 539 36604 555 36638
rect 489 36570 555 36604
rect 489 36536 505 36570
rect 539 36536 555 36570
rect 489 36502 555 36536
rect 489 36468 505 36502
rect 539 36468 555 36502
rect 489 36451 555 36468
rect 585 36706 651 36723
rect 585 36672 601 36706
rect 635 36672 651 36706
rect 585 36638 651 36672
rect 585 36604 601 36638
rect 635 36604 651 36638
rect 585 36570 651 36604
rect 585 36536 601 36570
rect 635 36536 651 36570
rect 585 36502 651 36536
rect 585 36468 601 36502
rect 635 36468 651 36502
rect 585 36451 651 36468
rect 681 36706 747 36723
rect 681 36672 697 36706
rect 731 36672 747 36706
rect 681 36638 747 36672
rect 681 36604 697 36638
rect 731 36604 747 36638
rect 681 36570 747 36604
rect 681 36536 697 36570
rect 731 36536 747 36570
rect 681 36502 747 36536
rect 681 36468 697 36502
rect 731 36468 747 36502
rect 681 36451 747 36468
rect 777 36706 843 36723
rect 777 36672 793 36706
rect 827 36672 843 36706
rect 777 36638 843 36672
rect 777 36604 793 36638
rect 827 36604 843 36638
rect 777 36570 843 36604
rect 777 36536 793 36570
rect 827 36536 843 36570
rect 777 36502 843 36536
rect 777 36468 793 36502
rect 827 36468 843 36502
rect 777 36451 843 36468
rect 873 36706 939 36723
rect 873 36672 889 36706
rect 923 36672 939 36706
rect 873 36638 939 36672
rect 873 36604 889 36638
rect 923 36604 939 36638
rect 873 36570 939 36604
rect 873 36536 889 36570
rect 923 36536 939 36570
rect 873 36502 939 36536
rect 873 36468 889 36502
rect 923 36468 939 36502
rect 873 36451 939 36468
rect 969 36706 1035 36723
rect 969 36672 985 36706
rect 1019 36672 1035 36706
rect 969 36638 1035 36672
rect 969 36604 985 36638
rect 1019 36604 1035 36638
rect 969 36570 1035 36604
rect 969 36536 985 36570
rect 1019 36536 1035 36570
rect 969 36502 1035 36536
rect 969 36468 985 36502
rect 1019 36468 1035 36502
rect 969 36451 1035 36468
rect 1065 36706 1131 36723
rect 1065 36672 1081 36706
rect 1115 36672 1131 36706
rect 1065 36638 1131 36672
rect 1065 36604 1081 36638
rect 1115 36604 1131 36638
rect 1065 36570 1131 36604
rect 1065 36536 1081 36570
rect 1115 36536 1131 36570
rect 1065 36502 1131 36536
rect 1065 36468 1081 36502
rect 1115 36468 1131 36502
rect 1065 36451 1131 36468
rect 1161 36706 1227 36723
rect 1161 36672 1177 36706
rect 1211 36672 1227 36706
rect 1161 36638 1227 36672
rect 1161 36604 1177 36638
rect 1211 36604 1227 36638
rect 1161 36570 1227 36604
rect 1161 36536 1177 36570
rect 1211 36536 1227 36570
rect 1161 36502 1227 36536
rect 1161 36468 1177 36502
rect 1211 36468 1227 36502
rect 1161 36451 1227 36468
rect 1257 36706 1319 36723
rect 1257 36672 1273 36706
rect 1307 36672 1319 36706
rect 1257 36638 1319 36672
rect 1257 36604 1273 36638
rect 1307 36604 1319 36638
rect 1257 36570 1319 36604
rect 1257 36536 1273 36570
rect 1307 36536 1319 36570
rect 1257 36502 1319 36536
rect 1257 36468 1273 36502
rect 1307 36468 1319 36502
rect 1257 36451 1319 36468
rect 2454 36710 2516 36727
rect 2454 36676 2466 36710
rect 2500 36676 2516 36710
rect 2454 36642 2516 36676
rect 2454 36608 2466 36642
rect 2500 36608 2516 36642
rect 2454 36574 2516 36608
rect 2454 36540 2466 36574
rect 2500 36540 2516 36574
rect 2454 36506 2516 36540
rect 2454 36472 2466 36506
rect 2500 36472 2516 36506
rect 2454 36455 2516 36472
rect 2546 36710 2612 36727
rect 2546 36676 2562 36710
rect 2596 36676 2612 36710
rect 2546 36642 2612 36676
rect 2546 36608 2562 36642
rect 2596 36608 2612 36642
rect 2546 36574 2612 36608
rect 2546 36540 2562 36574
rect 2596 36540 2612 36574
rect 2546 36506 2612 36540
rect 2546 36472 2562 36506
rect 2596 36472 2612 36506
rect 2546 36455 2612 36472
rect 2642 36710 2708 36727
rect 2642 36676 2658 36710
rect 2692 36676 2708 36710
rect 2642 36642 2708 36676
rect 2642 36608 2658 36642
rect 2692 36608 2708 36642
rect 2642 36574 2708 36608
rect 2642 36540 2658 36574
rect 2692 36540 2708 36574
rect 2642 36506 2708 36540
rect 2642 36472 2658 36506
rect 2692 36472 2708 36506
rect 2642 36455 2708 36472
rect 2738 36710 2804 36727
rect 2738 36676 2754 36710
rect 2788 36676 2804 36710
rect 2738 36642 2804 36676
rect 2738 36608 2754 36642
rect 2788 36608 2804 36642
rect 2738 36574 2804 36608
rect 2738 36540 2754 36574
rect 2788 36540 2804 36574
rect 2738 36506 2804 36540
rect 2738 36472 2754 36506
rect 2788 36472 2804 36506
rect 2738 36455 2804 36472
rect 2834 36710 2900 36727
rect 2834 36676 2850 36710
rect 2884 36676 2900 36710
rect 2834 36642 2900 36676
rect 2834 36608 2850 36642
rect 2884 36608 2900 36642
rect 2834 36574 2900 36608
rect 2834 36540 2850 36574
rect 2884 36540 2900 36574
rect 2834 36506 2900 36540
rect 2834 36472 2850 36506
rect 2884 36472 2900 36506
rect 2834 36455 2900 36472
rect 2930 36710 2996 36727
rect 2930 36676 2946 36710
rect 2980 36676 2996 36710
rect 2930 36642 2996 36676
rect 2930 36608 2946 36642
rect 2980 36608 2996 36642
rect 2930 36574 2996 36608
rect 2930 36540 2946 36574
rect 2980 36540 2996 36574
rect 2930 36506 2996 36540
rect 2930 36472 2946 36506
rect 2980 36472 2996 36506
rect 2930 36455 2996 36472
rect 3026 36710 3092 36727
rect 3026 36676 3042 36710
rect 3076 36676 3092 36710
rect 3026 36642 3092 36676
rect 3026 36608 3042 36642
rect 3076 36608 3092 36642
rect 3026 36574 3092 36608
rect 3026 36540 3042 36574
rect 3076 36540 3092 36574
rect 3026 36506 3092 36540
rect 3026 36472 3042 36506
rect 3076 36472 3092 36506
rect 3026 36455 3092 36472
rect 3122 36710 3188 36727
rect 3122 36676 3138 36710
rect 3172 36676 3188 36710
rect 3122 36642 3188 36676
rect 3122 36608 3138 36642
rect 3172 36608 3188 36642
rect 3122 36574 3188 36608
rect 3122 36540 3138 36574
rect 3172 36540 3188 36574
rect 3122 36506 3188 36540
rect 3122 36472 3138 36506
rect 3172 36472 3188 36506
rect 3122 36455 3188 36472
rect 3218 36710 3284 36727
rect 3218 36676 3234 36710
rect 3268 36676 3284 36710
rect 3218 36642 3284 36676
rect 3218 36608 3234 36642
rect 3268 36608 3284 36642
rect 3218 36574 3284 36608
rect 3218 36540 3234 36574
rect 3268 36540 3284 36574
rect 3218 36506 3284 36540
rect 3218 36472 3234 36506
rect 3268 36472 3284 36506
rect 3218 36455 3284 36472
rect 3314 36710 3380 36727
rect 3314 36676 3330 36710
rect 3364 36676 3380 36710
rect 3314 36642 3380 36676
rect 3314 36608 3330 36642
rect 3364 36608 3380 36642
rect 3314 36574 3380 36608
rect 3314 36540 3330 36574
rect 3364 36540 3380 36574
rect 3314 36506 3380 36540
rect 3314 36472 3330 36506
rect 3364 36472 3380 36506
rect 3314 36455 3380 36472
rect 3410 36710 3472 36727
rect 3410 36676 3426 36710
rect 3460 36676 3472 36710
rect 3410 36642 3472 36676
rect 3410 36608 3426 36642
rect 3460 36608 3472 36642
rect 3410 36574 3472 36608
rect 3410 36540 3426 36574
rect 3460 36540 3472 36574
rect 3410 36506 3472 36540
rect 3410 36472 3426 36506
rect 3460 36472 3472 36506
rect 3410 36455 3472 36472
rect 3975 36710 4037 36727
rect 3975 36676 3987 36710
rect 4021 36676 4037 36710
rect 3975 36642 4037 36676
rect 3975 36608 3987 36642
rect 4021 36608 4037 36642
rect 3975 36574 4037 36608
rect 3975 36540 3987 36574
rect 4021 36540 4037 36574
rect 3975 36506 4037 36540
rect 3975 36472 3987 36506
rect 4021 36472 4037 36506
rect 3975 36455 4037 36472
rect 4067 36710 4133 36727
rect 4067 36676 4083 36710
rect 4117 36676 4133 36710
rect 4067 36642 4133 36676
rect 4067 36608 4083 36642
rect 4117 36608 4133 36642
rect 4067 36574 4133 36608
rect 4067 36540 4083 36574
rect 4117 36540 4133 36574
rect 4067 36506 4133 36540
rect 4067 36472 4083 36506
rect 4117 36472 4133 36506
rect 4067 36455 4133 36472
rect 4163 36710 4229 36727
rect 4163 36676 4179 36710
rect 4213 36676 4229 36710
rect 4163 36642 4229 36676
rect 4163 36608 4179 36642
rect 4213 36608 4229 36642
rect 4163 36574 4229 36608
rect 4163 36540 4179 36574
rect 4213 36540 4229 36574
rect 4163 36506 4229 36540
rect 4163 36472 4179 36506
rect 4213 36472 4229 36506
rect 4163 36455 4229 36472
rect 4259 36710 4325 36727
rect 4259 36676 4275 36710
rect 4309 36676 4325 36710
rect 4259 36642 4325 36676
rect 4259 36608 4275 36642
rect 4309 36608 4325 36642
rect 4259 36574 4325 36608
rect 4259 36540 4275 36574
rect 4309 36540 4325 36574
rect 4259 36506 4325 36540
rect 4259 36472 4275 36506
rect 4309 36472 4325 36506
rect 4259 36455 4325 36472
rect 4355 36710 4421 36727
rect 4355 36676 4371 36710
rect 4405 36676 4421 36710
rect 4355 36642 4421 36676
rect 4355 36608 4371 36642
rect 4405 36608 4421 36642
rect 4355 36574 4421 36608
rect 4355 36540 4371 36574
rect 4405 36540 4421 36574
rect 4355 36506 4421 36540
rect 4355 36472 4371 36506
rect 4405 36472 4421 36506
rect 4355 36455 4421 36472
rect 4451 36710 4517 36727
rect 4451 36676 4467 36710
rect 4501 36676 4517 36710
rect 4451 36642 4517 36676
rect 4451 36608 4467 36642
rect 4501 36608 4517 36642
rect 4451 36574 4517 36608
rect 4451 36540 4467 36574
rect 4501 36540 4517 36574
rect 4451 36506 4517 36540
rect 4451 36472 4467 36506
rect 4501 36472 4517 36506
rect 4451 36455 4517 36472
rect 4547 36710 4613 36727
rect 4547 36676 4563 36710
rect 4597 36676 4613 36710
rect 4547 36642 4613 36676
rect 4547 36608 4563 36642
rect 4597 36608 4613 36642
rect 4547 36574 4613 36608
rect 4547 36540 4563 36574
rect 4597 36540 4613 36574
rect 4547 36506 4613 36540
rect 4547 36472 4563 36506
rect 4597 36472 4613 36506
rect 4547 36455 4613 36472
rect 4643 36710 4709 36727
rect 4643 36676 4659 36710
rect 4693 36676 4709 36710
rect 4643 36642 4709 36676
rect 4643 36608 4659 36642
rect 4693 36608 4709 36642
rect 4643 36574 4709 36608
rect 4643 36540 4659 36574
rect 4693 36540 4709 36574
rect 4643 36506 4709 36540
rect 4643 36472 4659 36506
rect 4693 36472 4709 36506
rect 4643 36455 4709 36472
rect 4739 36710 4805 36727
rect 4739 36676 4755 36710
rect 4789 36676 4805 36710
rect 4739 36642 4805 36676
rect 4739 36608 4755 36642
rect 4789 36608 4805 36642
rect 4739 36574 4805 36608
rect 4739 36540 4755 36574
rect 4789 36540 4805 36574
rect 4739 36506 4805 36540
rect 4739 36472 4755 36506
rect 4789 36472 4805 36506
rect 4739 36455 4805 36472
rect 4835 36710 4901 36727
rect 4835 36676 4851 36710
rect 4885 36676 4901 36710
rect 4835 36642 4901 36676
rect 4835 36608 4851 36642
rect 4885 36608 4901 36642
rect 4835 36574 4901 36608
rect 4835 36540 4851 36574
rect 4885 36540 4901 36574
rect 4835 36506 4901 36540
rect 4835 36472 4851 36506
rect 4885 36472 4901 36506
rect 4835 36455 4901 36472
rect 4931 36710 4993 36727
rect 4931 36676 4947 36710
rect 4981 36676 4993 36710
rect 4931 36642 4993 36676
rect 4931 36608 4947 36642
rect 4981 36608 4993 36642
rect 4931 36574 4993 36608
rect 4931 36540 4947 36574
rect 4981 36540 4993 36574
rect 4931 36506 4993 36540
rect 4931 36472 4947 36506
rect 4981 36472 4993 36506
rect 4931 36455 4993 36472
rect 5348 36502 5400 36514
rect 5348 36468 5356 36502
rect 5390 36468 5400 36502
rect 5348 36434 5400 36468
rect 5348 36400 5356 36434
rect 5390 36400 5400 36434
rect 5348 36366 5400 36400
rect 5348 36332 5356 36366
rect 5390 36332 5400 36366
rect 5348 36314 5400 36332
rect 5430 36502 5482 36514
rect 5430 36468 5440 36502
rect 5474 36468 5482 36502
rect 5430 36434 5482 36468
rect 5430 36400 5440 36434
rect 5474 36400 5482 36434
rect 5430 36366 5482 36400
rect 5430 36332 5440 36366
rect 5474 36332 5482 36366
rect 5430 36314 5482 36332
rect 301 35419 363 35436
rect 301 35385 313 35419
rect 347 35385 363 35419
rect 301 35351 363 35385
rect 301 35317 313 35351
rect 347 35317 363 35351
rect 301 35283 363 35317
rect 301 35249 313 35283
rect 347 35249 363 35283
rect 301 35215 363 35249
rect 301 35181 313 35215
rect 347 35181 363 35215
rect 301 35164 363 35181
rect 393 35419 459 35436
rect 393 35385 409 35419
rect 443 35385 459 35419
rect 393 35351 459 35385
rect 393 35317 409 35351
rect 443 35317 459 35351
rect 393 35283 459 35317
rect 393 35249 409 35283
rect 443 35249 459 35283
rect 393 35215 459 35249
rect 393 35181 409 35215
rect 443 35181 459 35215
rect 393 35164 459 35181
rect 489 35419 555 35436
rect 489 35385 505 35419
rect 539 35385 555 35419
rect 489 35351 555 35385
rect 489 35317 505 35351
rect 539 35317 555 35351
rect 489 35283 555 35317
rect 489 35249 505 35283
rect 539 35249 555 35283
rect 489 35215 555 35249
rect 489 35181 505 35215
rect 539 35181 555 35215
rect 489 35164 555 35181
rect 585 35419 651 35436
rect 585 35385 601 35419
rect 635 35385 651 35419
rect 585 35351 651 35385
rect 585 35317 601 35351
rect 635 35317 651 35351
rect 585 35283 651 35317
rect 585 35249 601 35283
rect 635 35249 651 35283
rect 585 35215 651 35249
rect 585 35181 601 35215
rect 635 35181 651 35215
rect 585 35164 651 35181
rect 681 35419 747 35436
rect 681 35385 697 35419
rect 731 35385 747 35419
rect 681 35351 747 35385
rect 681 35317 697 35351
rect 731 35317 747 35351
rect 681 35283 747 35317
rect 681 35249 697 35283
rect 731 35249 747 35283
rect 681 35215 747 35249
rect 681 35181 697 35215
rect 731 35181 747 35215
rect 681 35164 747 35181
rect 777 35419 843 35436
rect 777 35385 793 35419
rect 827 35385 843 35419
rect 777 35351 843 35385
rect 777 35317 793 35351
rect 827 35317 843 35351
rect 777 35283 843 35317
rect 777 35249 793 35283
rect 827 35249 843 35283
rect 777 35215 843 35249
rect 777 35181 793 35215
rect 827 35181 843 35215
rect 777 35164 843 35181
rect 873 35419 939 35436
rect 873 35385 889 35419
rect 923 35385 939 35419
rect 873 35351 939 35385
rect 873 35317 889 35351
rect 923 35317 939 35351
rect 873 35283 939 35317
rect 873 35249 889 35283
rect 923 35249 939 35283
rect 873 35215 939 35249
rect 873 35181 889 35215
rect 923 35181 939 35215
rect 873 35164 939 35181
rect 969 35419 1035 35436
rect 969 35385 985 35419
rect 1019 35385 1035 35419
rect 969 35351 1035 35385
rect 969 35317 985 35351
rect 1019 35317 1035 35351
rect 969 35283 1035 35317
rect 969 35249 985 35283
rect 1019 35249 1035 35283
rect 969 35215 1035 35249
rect 969 35181 985 35215
rect 1019 35181 1035 35215
rect 969 35164 1035 35181
rect 1065 35419 1131 35436
rect 1065 35385 1081 35419
rect 1115 35385 1131 35419
rect 1065 35351 1131 35385
rect 1065 35317 1081 35351
rect 1115 35317 1131 35351
rect 1065 35283 1131 35317
rect 1065 35249 1081 35283
rect 1115 35249 1131 35283
rect 1065 35215 1131 35249
rect 1065 35181 1081 35215
rect 1115 35181 1131 35215
rect 1065 35164 1131 35181
rect 1161 35419 1227 35436
rect 1161 35385 1177 35419
rect 1211 35385 1227 35419
rect 1161 35351 1227 35385
rect 1161 35317 1177 35351
rect 1211 35317 1227 35351
rect 1161 35283 1227 35317
rect 1161 35249 1177 35283
rect 1211 35249 1227 35283
rect 1161 35215 1227 35249
rect 1161 35181 1177 35215
rect 1211 35181 1227 35215
rect 1161 35164 1227 35181
rect 1257 35419 1319 35436
rect 1257 35385 1273 35419
rect 1307 35385 1319 35419
rect 1257 35351 1319 35385
rect 1257 35317 1273 35351
rect 1307 35317 1319 35351
rect 1257 35283 1319 35317
rect 1257 35249 1273 35283
rect 1307 35249 1319 35283
rect 1257 35215 1319 35249
rect 1257 35181 1273 35215
rect 1307 35181 1319 35215
rect 1257 35164 1319 35181
rect 2454 35423 2516 35440
rect 2454 35389 2466 35423
rect 2500 35389 2516 35423
rect 2454 35355 2516 35389
rect 2454 35321 2466 35355
rect 2500 35321 2516 35355
rect 2454 35287 2516 35321
rect 2454 35253 2466 35287
rect 2500 35253 2516 35287
rect 2454 35219 2516 35253
rect 2454 35185 2466 35219
rect 2500 35185 2516 35219
rect 2454 35168 2516 35185
rect 2546 35423 2612 35440
rect 2546 35389 2562 35423
rect 2596 35389 2612 35423
rect 2546 35355 2612 35389
rect 2546 35321 2562 35355
rect 2596 35321 2612 35355
rect 2546 35287 2612 35321
rect 2546 35253 2562 35287
rect 2596 35253 2612 35287
rect 2546 35219 2612 35253
rect 2546 35185 2562 35219
rect 2596 35185 2612 35219
rect 2546 35168 2612 35185
rect 2642 35423 2708 35440
rect 2642 35389 2658 35423
rect 2692 35389 2708 35423
rect 2642 35355 2708 35389
rect 2642 35321 2658 35355
rect 2692 35321 2708 35355
rect 2642 35287 2708 35321
rect 2642 35253 2658 35287
rect 2692 35253 2708 35287
rect 2642 35219 2708 35253
rect 2642 35185 2658 35219
rect 2692 35185 2708 35219
rect 2642 35168 2708 35185
rect 2738 35423 2804 35440
rect 2738 35389 2754 35423
rect 2788 35389 2804 35423
rect 2738 35355 2804 35389
rect 2738 35321 2754 35355
rect 2788 35321 2804 35355
rect 2738 35287 2804 35321
rect 2738 35253 2754 35287
rect 2788 35253 2804 35287
rect 2738 35219 2804 35253
rect 2738 35185 2754 35219
rect 2788 35185 2804 35219
rect 2738 35168 2804 35185
rect 2834 35423 2900 35440
rect 2834 35389 2850 35423
rect 2884 35389 2900 35423
rect 2834 35355 2900 35389
rect 2834 35321 2850 35355
rect 2884 35321 2900 35355
rect 2834 35287 2900 35321
rect 2834 35253 2850 35287
rect 2884 35253 2900 35287
rect 2834 35219 2900 35253
rect 2834 35185 2850 35219
rect 2884 35185 2900 35219
rect 2834 35168 2900 35185
rect 2930 35423 2996 35440
rect 2930 35389 2946 35423
rect 2980 35389 2996 35423
rect 2930 35355 2996 35389
rect 2930 35321 2946 35355
rect 2980 35321 2996 35355
rect 2930 35287 2996 35321
rect 2930 35253 2946 35287
rect 2980 35253 2996 35287
rect 2930 35219 2996 35253
rect 2930 35185 2946 35219
rect 2980 35185 2996 35219
rect 2930 35168 2996 35185
rect 3026 35423 3092 35440
rect 3026 35389 3042 35423
rect 3076 35389 3092 35423
rect 3026 35355 3092 35389
rect 3026 35321 3042 35355
rect 3076 35321 3092 35355
rect 3026 35287 3092 35321
rect 3026 35253 3042 35287
rect 3076 35253 3092 35287
rect 3026 35219 3092 35253
rect 3026 35185 3042 35219
rect 3076 35185 3092 35219
rect 3026 35168 3092 35185
rect 3122 35423 3188 35440
rect 3122 35389 3138 35423
rect 3172 35389 3188 35423
rect 3122 35355 3188 35389
rect 3122 35321 3138 35355
rect 3172 35321 3188 35355
rect 3122 35287 3188 35321
rect 3122 35253 3138 35287
rect 3172 35253 3188 35287
rect 3122 35219 3188 35253
rect 3122 35185 3138 35219
rect 3172 35185 3188 35219
rect 3122 35168 3188 35185
rect 3218 35423 3284 35440
rect 3218 35389 3234 35423
rect 3268 35389 3284 35423
rect 3218 35355 3284 35389
rect 3218 35321 3234 35355
rect 3268 35321 3284 35355
rect 3218 35287 3284 35321
rect 3218 35253 3234 35287
rect 3268 35253 3284 35287
rect 3218 35219 3284 35253
rect 3218 35185 3234 35219
rect 3268 35185 3284 35219
rect 3218 35168 3284 35185
rect 3314 35423 3380 35440
rect 3314 35389 3330 35423
rect 3364 35389 3380 35423
rect 3314 35355 3380 35389
rect 3314 35321 3330 35355
rect 3364 35321 3380 35355
rect 3314 35287 3380 35321
rect 3314 35253 3330 35287
rect 3364 35253 3380 35287
rect 3314 35219 3380 35253
rect 3314 35185 3330 35219
rect 3364 35185 3380 35219
rect 3314 35168 3380 35185
rect 3410 35423 3472 35440
rect 3410 35389 3426 35423
rect 3460 35389 3472 35423
rect 3410 35355 3472 35389
rect 3410 35321 3426 35355
rect 3460 35321 3472 35355
rect 3410 35287 3472 35321
rect 3410 35253 3426 35287
rect 3460 35253 3472 35287
rect 3410 35219 3472 35253
rect 3410 35185 3426 35219
rect 3460 35185 3472 35219
rect 3410 35168 3472 35185
rect 3975 35423 4037 35440
rect 3975 35389 3987 35423
rect 4021 35389 4037 35423
rect 3975 35355 4037 35389
rect 3975 35321 3987 35355
rect 4021 35321 4037 35355
rect 3975 35287 4037 35321
rect 3975 35253 3987 35287
rect 4021 35253 4037 35287
rect 3975 35219 4037 35253
rect 3975 35185 3987 35219
rect 4021 35185 4037 35219
rect 3975 35168 4037 35185
rect 4067 35423 4133 35440
rect 4067 35389 4083 35423
rect 4117 35389 4133 35423
rect 4067 35355 4133 35389
rect 4067 35321 4083 35355
rect 4117 35321 4133 35355
rect 4067 35287 4133 35321
rect 4067 35253 4083 35287
rect 4117 35253 4133 35287
rect 4067 35219 4133 35253
rect 4067 35185 4083 35219
rect 4117 35185 4133 35219
rect 4067 35168 4133 35185
rect 4163 35423 4229 35440
rect 4163 35389 4179 35423
rect 4213 35389 4229 35423
rect 4163 35355 4229 35389
rect 4163 35321 4179 35355
rect 4213 35321 4229 35355
rect 4163 35287 4229 35321
rect 4163 35253 4179 35287
rect 4213 35253 4229 35287
rect 4163 35219 4229 35253
rect 4163 35185 4179 35219
rect 4213 35185 4229 35219
rect 4163 35168 4229 35185
rect 4259 35423 4325 35440
rect 4259 35389 4275 35423
rect 4309 35389 4325 35423
rect 4259 35355 4325 35389
rect 4259 35321 4275 35355
rect 4309 35321 4325 35355
rect 4259 35287 4325 35321
rect 4259 35253 4275 35287
rect 4309 35253 4325 35287
rect 4259 35219 4325 35253
rect 4259 35185 4275 35219
rect 4309 35185 4325 35219
rect 4259 35168 4325 35185
rect 4355 35423 4421 35440
rect 4355 35389 4371 35423
rect 4405 35389 4421 35423
rect 4355 35355 4421 35389
rect 4355 35321 4371 35355
rect 4405 35321 4421 35355
rect 4355 35287 4421 35321
rect 4355 35253 4371 35287
rect 4405 35253 4421 35287
rect 4355 35219 4421 35253
rect 4355 35185 4371 35219
rect 4405 35185 4421 35219
rect 4355 35168 4421 35185
rect 4451 35423 4517 35440
rect 4451 35389 4467 35423
rect 4501 35389 4517 35423
rect 4451 35355 4517 35389
rect 4451 35321 4467 35355
rect 4501 35321 4517 35355
rect 4451 35287 4517 35321
rect 4451 35253 4467 35287
rect 4501 35253 4517 35287
rect 4451 35219 4517 35253
rect 4451 35185 4467 35219
rect 4501 35185 4517 35219
rect 4451 35168 4517 35185
rect 4547 35423 4613 35440
rect 4547 35389 4563 35423
rect 4597 35389 4613 35423
rect 4547 35355 4613 35389
rect 4547 35321 4563 35355
rect 4597 35321 4613 35355
rect 4547 35287 4613 35321
rect 4547 35253 4563 35287
rect 4597 35253 4613 35287
rect 4547 35219 4613 35253
rect 4547 35185 4563 35219
rect 4597 35185 4613 35219
rect 4547 35168 4613 35185
rect 4643 35423 4709 35440
rect 4643 35389 4659 35423
rect 4693 35389 4709 35423
rect 4643 35355 4709 35389
rect 4643 35321 4659 35355
rect 4693 35321 4709 35355
rect 4643 35287 4709 35321
rect 4643 35253 4659 35287
rect 4693 35253 4709 35287
rect 4643 35219 4709 35253
rect 4643 35185 4659 35219
rect 4693 35185 4709 35219
rect 4643 35168 4709 35185
rect 4739 35423 4805 35440
rect 4739 35389 4755 35423
rect 4789 35389 4805 35423
rect 4739 35355 4805 35389
rect 4739 35321 4755 35355
rect 4789 35321 4805 35355
rect 4739 35287 4805 35321
rect 4739 35253 4755 35287
rect 4789 35253 4805 35287
rect 4739 35219 4805 35253
rect 4739 35185 4755 35219
rect 4789 35185 4805 35219
rect 4739 35168 4805 35185
rect 4835 35423 4901 35440
rect 4835 35389 4851 35423
rect 4885 35389 4901 35423
rect 4835 35355 4901 35389
rect 4835 35321 4851 35355
rect 4885 35321 4901 35355
rect 4835 35287 4901 35321
rect 4835 35253 4851 35287
rect 4885 35253 4901 35287
rect 4835 35219 4901 35253
rect 4835 35185 4851 35219
rect 4885 35185 4901 35219
rect 4835 35168 4901 35185
rect 4931 35423 4993 35440
rect 4931 35389 4947 35423
rect 4981 35389 4993 35423
rect 4931 35355 4993 35389
rect 4931 35321 4947 35355
rect 4981 35321 4993 35355
rect 4931 35287 4993 35321
rect 4931 35253 4947 35287
rect 4981 35253 4993 35287
rect 4931 35219 4993 35253
rect 4931 35185 4947 35219
rect 4981 35185 4993 35219
rect 4931 35168 4993 35185
rect 5348 35215 5400 35227
rect 5348 35181 5356 35215
rect 5390 35181 5400 35215
rect 5348 35147 5400 35181
rect 5348 35113 5356 35147
rect 5390 35113 5400 35147
rect 5348 35079 5400 35113
rect 5348 35045 5356 35079
rect 5390 35045 5400 35079
rect 5348 35027 5400 35045
rect 5430 35215 5482 35227
rect 5430 35181 5440 35215
rect 5474 35181 5482 35215
rect 5430 35147 5482 35181
rect 5430 35113 5440 35147
rect 5474 35113 5482 35147
rect 5430 35079 5482 35113
rect 5430 35045 5440 35079
rect 5474 35045 5482 35079
rect 5430 35027 5482 35045
rect 301 34132 363 34149
rect 301 34098 313 34132
rect 347 34098 363 34132
rect 301 34064 363 34098
rect 301 34030 313 34064
rect 347 34030 363 34064
rect 301 33996 363 34030
rect 301 33962 313 33996
rect 347 33962 363 33996
rect 301 33928 363 33962
rect 301 33894 313 33928
rect 347 33894 363 33928
rect 301 33877 363 33894
rect 393 34132 459 34149
rect 393 34098 409 34132
rect 443 34098 459 34132
rect 393 34064 459 34098
rect 393 34030 409 34064
rect 443 34030 459 34064
rect 393 33996 459 34030
rect 393 33962 409 33996
rect 443 33962 459 33996
rect 393 33928 459 33962
rect 393 33894 409 33928
rect 443 33894 459 33928
rect 393 33877 459 33894
rect 489 34132 555 34149
rect 489 34098 505 34132
rect 539 34098 555 34132
rect 489 34064 555 34098
rect 489 34030 505 34064
rect 539 34030 555 34064
rect 489 33996 555 34030
rect 489 33962 505 33996
rect 539 33962 555 33996
rect 489 33928 555 33962
rect 489 33894 505 33928
rect 539 33894 555 33928
rect 489 33877 555 33894
rect 585 34132 651 34149
rect 585 34098 601 34132
rect 635 34098 651 34132
rect 585 34064 651 34098
rect 585 34030 601 34064
rect 635 34030 651 34064
rect 585 33996 651 34030
rect 585 33962 601 33996
rect 635 33962 651 33996
rect 585 33928 651 33962
rect 585 33894 601 33928
rect 635 33894 651 33928
rect 585 33877 651 33894
rect 681 34132 747 34149
rect 681 34098 697 34132
rect 731 34098 747 34132
rect 681 34064 747 34098
rect 681 34030 697 34064
rect 731 34030 747 34064
rect 681 33996 747 34030
rect 681 33962 697 33996
rect 731 33962 747 33996
rect 681 33928 747 33962
rect 681 33894 697 33928
rect 731 33894 747 33928
rect 681 33877 747 33894
rect 777 34132 843 34149
rect 777 34098 793 34132
rect 827 34098 843 34132
rect 777 34064 843 34098
rect 777 34030 793 34064
rect 827 34030 843 34064
rect 777 33996 843 34030
rect 777 33962 793 33996
rect 827 33962 843 33996
rect 777 33928 843 33962
rect 777 33894 793 33928
rect 827 33894 843 33928
rect 777 33877 843 33894
rect 873 34132 939 34149
rect 873 34098 889 34132
rect 923 34098 939 34132
rect 873 34064 939 34098
rect 873 34030 889 34064
rect 923 34030 939 34064
rect 873 33996 939 34030
rect 873 33962 889 33996
rect 923 33962 939 33996
rect 873 33928 939 33962
rect 873 33894 889 33928
rect 923 33894 939 33928
rect 873 33877 939 33894
rect 969 34132 1035 34149
rect 969 34098 985 34132
rect 1019 34098 1035 34132
rect 969 34064 1035 34098
rect 969 34030 985 34064
rect 1019 34030 1035 34064
rect 969 33996 1035 34030
rect 969 33962 985 33996
rect 1019 33962 1035 33996
rect 969 33928 1035 33962
rect 969 33894 985 33928
rect 1019 33894 1035 33928
rect 969 33877 1035 33894
rect 1065 34132 1131 34149
rect 1065 34098 1081 34132
rect 1115 34098 1131 34132
rect 1065 34064 1131 34098
rect 1065 34030 1081 34064
rect 1115 34030 1131 34064
rect 1065 33996 1131 34030
rect 1065 33962 1081 33996
rect 1115 33962 1131 33996
rect 1065 33928 1131 33962
rect 1065 33894 1081 33928
rect 1115 33894 1131 33928
rect 1065 33877 1131 33894
rect 1161 34132 1227 34149
rect 1161 34098 1177 34132
rect 1211 34098 1227 34132
rect 1161 34064 1227 34098
rect 1161 34030 1177 34064
rect 1211 34030 1227 34064
rect 1161 33996 1227 34030
rect 1161 33962 1177 33996
rect 1211 33962 1227 33996
rect 1161 33928 1227 33962
rect 1161 33894 1177 33928
rect 1211 33894 1227 33928
rect 1161 33877 1227 33894
rect 1257 34132 1319 34149
rect 1257 34098 1273 34132
rect 1307 34098 1319 34132
rect 1257 34064 1319 34098
rect 1257 34030 1273 34064
rect 1307 34030 1319 34064
rect 1257 33996 1319 34030
rect 1257 33962 1273 33996
rect 1307 33962 1319 33996
rect 1257 33928 1319 33962
rect 1257 33894 1273 33928
rect 1307 33894 1319 33928
rect 1257 33877 1319 33894
rect 2454 34136 2516 34153
rect 2454 34102 2466 34136
rect 2500 34102 2516 34136
rect 2454 34068 2516 34102
rect 2454 34034 2466 34068
rect 2500 34034 2516 34068
rect 2454 34000 2516 34034
rect 2454 33966 2466 34000
rect 2500 33966 2516 34000
rect 2454 33932 2516 33966
rect 2454 33898 2466 33932
rect 2500 33898 2516 33932
rect 2454 33881 2516 33898
rect 2546 34136 2612 34153
rect 2546 34102 2562 34136
rect 2596 34102 2612 34136
rect 2546 34068 2612 34102
rect 2546 34034 2562 34068
rect 2596 34034 2612 34068
rect 2546 34000 2612 34034
rect 2546 33966 2562 34000
rect 2596 33966 2612 34000
rect 2546 33932 2612 33966
rect 2546 33898 2562 33932
rect 2596 33898 2612 33932
rect 2546 33881 2612 33898
rect 2642 34136 2708 34153
rect 2642 34102 2658 34136
rect 2692 34102 2708 34136
rect 2642 34068 2708 34102
rect 2642 34034 2658 34068
rect 2692 34034 2708 34068
rect 2642 34000 2708 34034
rect 2642 33966 2658 34000
rect 2692 33966 2708 34000
rect 2642 33932 2708 33966
rect 2642 33898 2658 33932
rect 2692 33898 2708 33932
rect 2642 33881 2708 33898
rect 2738 34136 2804 34153
rect 2738 34102 2754 34136
rect 2788 34102 2804 34136
rect 2738 34068 2804 34102
rect 2738 34034 2754 34068
rect 2788 34034 2804 34068
rect 2738 34000 2804 34034
rect 2738 33966 2754 34000
rect 2788 33966 2804 34000
rect 2738 33932 2804 33966
rect 2738 33898 2754 33932
rect 2788 33898 2804 33932
rect 2738 33881 2804 33898
rect 2834 34136 2900 34153
rect 2834 34102 2850 34136
rect 2884 34102 2900 34136
rect 2834 34068 2900 34102
rect 2834 34034 2850 34068
rect 2884 34034 2900 34068
rect 2834 34000 2900 34034
rect 2834 33966 2850 34000
rect 2884 33966 2900 34000
rect 2834 33932 2900 33966
rect 2834 33898 2850 33932
rect 2884 33898 2900 33932
rect 2834 33881 2900 33898
rect 2930 34136 2996 34153
rect 2930 34102 2946 34136
rect 2980 34102 2996 34136
rect 2930 34068 2996 34102
rect 2930 34034 2946 34068
rect 2980 34034 2996 34068
rect 2930 34000 2996 34034
rect 2930 33966 2946 34000
rect 2980 33966 2996 34000
rect 2930 33932 2996 33966
rect 2930 33898 2946 33932
rect 2980 33898 2996 33932
rect 2930 33881 2996 33898
rect 3026 34136 3092 34153
rect 3026 34102 3042 34136
rect 3076 34102 3092 34136
rect 3026 34068 3092 34102
rect 3026 34034 3042 34068
rect 3076 34034 3092 34068
rect 3026 34000 3092 34034
rect 3026 33966 3042 34000
rect 3076 33966 3092 34000
rect 3026 33932 3092 33966
rect 3026 33898 3042 33932
rect 3076 33898 3092 33932
rect 3026 33881 3092 33898
rect 3122 34136 3188 34153
rect 3122 34102 3138 34136
rect 3172 34102 3188 34136
rect 3122 34068 3188 34102
rect 3122 34034 3138 34068
rect 3172 34034 3188 34068
rect 3122 34000 3188 34034
rect 3122 33966 3138 34000
rect 3172 33966 3188 34000
rect 3122 33932 3188 33966
rect 3122 33898 3138 33932
rect 3172 33898 3188 33932
rect 3122 33881 3188 33898
rect 3218 34136 3284 34153
rect 3218 34102 3234 34136
rect 3268 34102 3284 34136
rect 3218 34068 3284 34102
rect 3218 34034 3234 34068
rect 3268 34034 3284 34068
rect 3218 34000 3284 34034
rect 3218 33966 3234 34000
rect 3268 33966 3284 34000
rect 3218 33932 3284 33966
rect 3218 33898 3234 33932
rect 3268 33898 3284 33932
rect 3218 33881 3284 33898
rect 3314 34136 3380 34153
rect 3314 34102 3330 34136
rect 3364 34102 3380 34136
rect 3314 34068 3380 34102
rect 3314 34034 3330 34068
rect 3364 34034 3380 34068
rect 3314 34000 3380 34034
rect 3314 33966 3330 34000
rect 3364 33966 3380 34000
rect 3314 33932 3380 33966
rect 3314 33898 3330 33932
rect 3364 33898 3380 33932
rect 3314 33881 3380 33898
rect 3410 34136 3472 34153
rect 3410 34102 3426 34136
rect 3460 34102 3472 34136
rect 3410 34068 3472 34102
rect 3410 34034 3426 34068
rect 3460 34034 3472 34068
rect 3410 34000 3472 34034
rect 3410 33966 3426 34000
rect 3460 33966 3472 34000
rect 3410 33932 3472 33966
rect 3410 33898 3426 33932
rect 3460 33898 3472 33932
rect 3410 33881 3472 33898
rect 3975 34136 4037 34153
rect 3975 34102 3987 34136
rect 4021 34102 4037 34136
rect 3975 34068 4037 34102
rect 3975 34034 3987 34068
rect 4021 34034 4037 34068
rect 3975 34000 4037 34034
rect 3975 33966 3987 34000
rect 4021 33966 4037 34000
rect 3975 33932 4037 33966
rect 3975 33898 3987 33932
rect 4021 33898 4037 33932
rect 3975 33881 4037 33898
rect 4067 34136 4133 34153
rect 4067 34102 4083 34136
rect 4117 34102 4133 34136
rect 4067 34068 4133 34102
rect 4067 34034 4083 34068
rect 4117 34034 4133 34068
rect 4067 34000 4133 34034
rect 4067 33966 4083 34000
rect 4117 33966 4133 34000
rect 4067 33932 4133 33966
rect 4067 33898 4083 33932
rect 4117 33898 4133 33932
rect 4067 33881 4133 33898
rect 4163 34136 4229 34153
rect 4163 34102 4179 34136
rect 4213 34102 4229 34136
rect 4163 34068 4229 34102
rect 4163 34034 4179 34068
rect 4213 34034 4229 34068
rect 4163 34000 4229 34034
rect 4163 33966 4179 34000
rect 4213 33966 4229 34000
rect 4163 33932 4229 33966
rect 4163 33898 4179 33932
rect 4213 33898 4229 33932
rect 4163 33881 4229 33898
rect 4259 34136 4325 34153
rect 4259 34102 4275 34136
rect 4309 34102 4325 34136
rect 4259 34068 4325 34102
rect 4259 34034 4275 34068
rect 4309 34034 4325 34068
rect 4259 34000 4325 34034
rect 4259 33966 4275 34000
rect 4309 33966 4325 34000
rect 4259 33932 4325 33966
rect 4259 33898 4275 33932
rect 4309 33898 4325 33932
rect 4259 33881 4325 33898
rect 4355 34136 4421 34153
rect 4355 34102 4371 34136
rect 4405 34102 4421 34136
rect 4355 34068 4421 34102
rect 4355 34034 4371 34068
rect 4405 34034 4421 34068
rect 4355 34000 4421 34034
rect 4355 33966 4371 34000
rect 4405 33966 4421 34000
rect 4355 33932 4421 33966
rect 4355 33898 4371 33932
rect 4405 33898 4421 33932
rect 4355 33881 4421 33898
rect 4451 34136 4517 34153
rect 4451 34102 4467 34136
rect 4501 34102 4517 34136
rect 4451 34068 4517 34102
rect 4451 34034 4467 34068
rect 4501 34034 4517 34068
rect 4451 34000 4517 34034
rect 4451 33966 4467 34000
rect 4501 33966 4517 34000
rect 4451 33932 4517 33966
rect 4451 33898 4467 33932
rect 4501 33898 4517 33932
rect 4451 33881 4517 33898
rect 4547 34136 4613 34153
rect 4547 34102 4563 34136
rect 4597 34102 4613 34136
rect 4547 34068 4613 34102
rect 4547 34034 4563 34068
rect 4597 34034 4613 34068
rect 4547 34000 4613 34034
rect 4547 33966 4563 34000
rect 4597 33966 4613 34000
rect 4547 33932 4613 33966
rect 4547 33898 4563 33932
rect 4597 33898 4613 33932
rect 4547 33881 4613 33898
rect 4643 34136 4709 34153
rect 4643 34102 4659 34136
rect 4693 34102 4709 34136
rect 4643 34068 4709 34102
rect 4643 34034 4659 34068
rect 4693 34034 4709 34068
rect 4643 34000 4709 34034
rect 4643 33966 4659 34000
rect 4693 33966 4709 34000
rect 4643 33932 4709 33966
rect 4643 33898 4659 33932
rect 4693 33898 4709 33932
rect 4643 33881 4709 33898
rect 4739 34136 4805 34153
rect 4739 34102 4755 34136
rect 4789 34102 4805 34136
rect 4739 34068 4805 34102
rect 4739 34034 4755 34068
rect 4789 34034 4805 34068
rect 4739 34000 4805 34034
rect 4739 33966 4755 34000
rect 4789 33966 4805 34000
rect 4739 33932 4805 33966
rect 4739 33898 4755 33932
rect 4789 33898 4805 33932
rect 4739 33881 4805 33898
rect 4835 34136 4901 34153
rect 4835 34102 4851 34136
rect 4885 34102 4901 34136
rect 4835 34068 4901 34102
rect 4835 34034 4851 34068
rect 4885 34034 4901 34068
rect 4835 34000 4901 34034
rect 4835 33966 4851 34000
rect 4885 33966 4901 34000
rect 4835 33932 4901 33966
rect 4835 33898 4851 33932
rect 4885 33898 4901 33932
rect 4835 33881 4901 33898
rect 4931 34136 4993 34153
rect 4931 34102 4947 34136
rect 4981 34102 4993 34136
rect 4931 34068 4993 34102
rect 4931 34034 4947 34068
rect 4981 34034 4993 34068
rect 4931 34000 4993 34034
rect 4931 33966 4947 34000
rect 4981 33966 4993 34000
rect 4931 33932 4993 33966
rect 4931 33898 4947 33932
rect 4981 33898 4993 33932
rect 4931 33881 4993 33898
rect 5348 33928 5400 33940
rect 5348 33894 5356 33928
rect 5390 33894 5400 33928
rect 5348 33860 5400 33894
rect 5348 33826 5356 33860
rect 5390 33826 5400 33860
rect 5348 33792 5400 33826
rect 5348 33758 5356 33792
rect 5390 33758 5400 33792
rect 5348 33740 5400 33758
rect 5430 33928 5482 33940
rect 5430 33894 5440 33928
rect 5474 33894 5482 33928
rect 5430 33860 5482 33894
rect 5430 33826 5440 33860
rect 5474 33826 5482 33860
rect 5430 33792 5482 33826
rect 5430 33758 5440 33792
rect 5474 33758 5482 33792
rect 5430 33740 5482 33758
rect 301 32845 363 32862
rect 301 32811 313 32845
rect 347 32811 363 32845
rect 301 32777 363 32811
rect 301 32743 313 32777
rect 347 32743 363 32777
rect 301 32709 363 32743
rect 301 32675 313 32709
rect 347 32675 363 32709
rect 301 32641 363 32675
rect 301 32607 313 32641
rect 347 32607 363 32641
rect 301 32590 363 32607
rect 393 32845 459 32862
rect 393 32811 409 32845
rect 443 32811 459 32845
rect 393 32777 459 32811
rect 393 32743 409 32777
rect 443 32743 459 32777
rect 393 32709 459 32743
rect 393 32675 409 32709
rect 443 32675 459 32709
rect 393 32641 459 32675
rect 393 32607 409 32641
rect 443 32607 459 32641
rect 393 32590 459 32607
rect 489 32845 555 32862
rect 489 32811 505 32845
rect 539 32811 555 32845
rect 489 32777 555 32811
rect 489 32743 505 32777
rect 539 32743 555 32777
rect 489 32709 555 32743
rect 489 32675 505 32709
rect 539 32675 555 32709
rect 489 32641 555 32675
rect 489 32607 505 32641
rect 539 32607 555 32641
rect 489 32590 555 32607
rect 585 32845 651 32862
rect 585 32811 601 32845
rect 635 32811 651 32845
rect 585 32777 651 32811
rect 585 32743 601 32777
rect 635 32743 651 32777
rect 585 32709 651 32743
rect 585 32675 601 32709
rect 635 32675 651 32709
rect 585 32641 651 32675
rect 585 32607 601 32641
rect 635 32607 651 32641
rect 585 32590 651 32607
rect 681 32845 747 32862
rect 681 32811 697 32845
rect 731 32811 747 32845
rect 681 32777 747 32811
rect 681 32743 697 32777
rect 731 32743 747 32777
rect 681 32709 747 32743
rect 681 32675 697 32709
rect 731 32675 747 32709
rect 681 32641 747 32675
rect 681 32607 697 32641
rect 731 32607 747 32641
rect 681 32590 747 32607
rect 777 32845 843 32862
rect 777 32811 793 32845
rect 827 32811 843 32845
rect 777 32777 843 32811
rect 777 32743 793 32777
rect 827 32743 843 32777
rect 777 32709 843 32743
rect 777 32675 793 32709
rect 827 32675 843 32709
rect 777 32641 843 32675
rect 777 32607 793 32641
rect 827 32607 843 32641
rect 777 32590 843 32607
rect 873 32845 939 32862
rect 873 32811 889 32845
rect 923 32811 939 32845
rect 873 32777 939 32811
rect 873 32743 889 32777
rect 923 32743 939 32777
rect 873 32709 939 32743
rect 873 32675 889 32709
rect 923 32675 939 32709
rect 873 32641 939 32675
rect 873 32607 889 32641
rect 923 32607 939 32641
rect 873 32590 939 32607
rect 969 32845 1035 32862
rect 969 32811 985 32845
rect 1019 32811 1035 32845
rect 969 32777 1035 32811
rect 969 32743 985 32777
rect 1019 32743 1035 32777
rect 969 32709 1035 32743
rect 969 32675 985 32709
rect 1019 32675 1035 32709
rect 969 32641 1035 32675
rect 969 32607 985 32641
rect 1019 32607 1035 32641
rect 969 32590 1035 32607
rect 1065 32845 1131 32862
rect 1065 32811 1081 32845
rect 1115 32811 1131 32845
rect 1065 32777 1131 32811
rect 1065 32743 1081 32777
rect 1115 32743 1131 32777
rect 1065 32709 1131 32743
rect 1065 32675 1081 32709
rect 1115 32675 1131 32709
rect 1065 32641 1131 32675
rect 1065 32607 1081 32641
rect 1115 32607 1131 32641
rect 1065 32590 1131 32607
rect 1161 32845 1227 32862
rect 1161 32811 1177 32845
rect 1211 32811 1227 32845
rect 1161 32777 1227 32811
rect 1161 32743 1177 32777
rect 1211 32743 1227 32777
rect 1161 32709 1227 32743
rect 1161 32675 1177 32709
rect 1211 32675 1227 32709
rect 1161 32641 1227 32675
rect 1161 32607 1177 32641
rect 1211 32607 1227 32641
rect 1161 32590 1227 32607
rect 1257 32845 1319 32862
rect 1257 32811 1273 32845
rect 1307 32811 1319 32845
rect 1257 32777 1319 32811
rect 1257 32743 1273 32777
rect 1307 32743 1319 32777
rect 1257 32709 1319 32743
rect 1257 32675 1273 32709
rect 1307 32675 1319 32709
rect 1257 32641 1319 32675
rect 1257 32607 1273 32641
rect 1307 32607 1319 32641
rect 1257 32590 1319 32607
rect 2454 32849 2516 32866
rect 2454 32815 2466 32849
rect 2500 32815 2516 32849
rect 2454 32781 2516 32815
rect 2454 32747 2466 32781
rect 2500 32747 2516 32781
rect 2454 32713 2516 32747
rect 2454 32679 2466 32713
rect 2500 32679 2516 32713
rect 2454 32645 2516 32679
rect 2454 32611 2466 32645
rect 2500 32611 2516 32645
rect 2454 32594 2516 32611
rect 2546 32849 2612 32866
rect 2546 32815 2562 32849
rect 2596 32815 2612 32849
rect 2546 32781 2612 32815
rect 2546 32747 2562 32781
rect 2596 32747 2612 32781
rect 2546 32713 2612 32747
rect 2546 32679 2562 32713
rect 2596 32679 2612 32713
rect 2546 32645 2612 32679
rect 2546 32611 2562 32645
rect 2596 32611 2612 32645
rect 2546 32594 2612 32611
rect 2642 32849 2708 32866
rect 2642 32815 2658 32849
rect 2692 32815 2708 32849
rect 2642 32781 2708 32815
rect 2642 32747 2658 32781
rect 2692 32747 2708 32781
rect 2642 32713 2708 32747
rect 2642 32679 2658 32713
rect 2692 32679 2708 32713
rect 2642 32645 2708 32679
rect 2642 32611 2658 32645
rect 2692 32611 2708 32645
rect 2642 32594 2708 32611
rect 2738 32849 2804 32866
rect 2738 32815 2754 32849
rect 2788 32815 2804 32849
rect 2738 32781 2804 32815
rect 2738 32747 2754 32781
rect 2788 32747 2804 32781
rect 2738 32713 2804 32747
rect 2738 32679 2754 32713
rect 2788 32679 2804 32713
rect 2738 32645 2804 32679
rect 2738 32611 2754 32645
rect 2788 32611 2804 32645
rect 2738 32594 2804 32611
rect 2834 32849 2900 32866
rect 2834 32815 2850 32849
rect 2884 32815 2900 32849
rect 2834 32781 2900 32815
rect 2834 32747 2850 32781
rect 2884 32747 2900 32781
rect 2834 32713 2900 32747
rect 2834 32679 2850 32713
rect 2884 32679 2900 32713
rect 2834 32645 2900 32679
rect 2834 32611 2850 32645
rect 2884 32611 2900 32645
rect 2834 32594 2900 32611
rect 2930 32849 2996 32866
rect 2930 32815 2946 32849
rect 2980 32815 2996 32849
rect 2930 32781 2996 32815
rect 2930 32747 2946 32781
rect 2980 32747 2996 32781
rect 2930 32713 2996 32747
rect 2930 32679 2946 32713
rect 2980 32679 2996 32713
rect 2930 32645 2996 32679
rect 2930 32611 2946 32645
rect 2980 32611 2996 32645
rect 2930 32594 2996 32611
rect 3026 32849 3092 32866
rect 3026 32815 3042 32849
rect 3076 32815 3092 32849
rect 3026 32781 3092 32815
rect 3026 32747 3042 32781
rect 3076 32747 3092 32781
rect 3026 32713 3092 32747
rect 3026 32679 3042 32713
rect 3076 32679 3092 32713
rect 3026 32645 3092 32679
rect 3026 32611 3042 32645
rect 3076 32611 3092 32645
rect 3026 32594 3092 32611
rect 3122 32849 3188 32866
rect 3122 32815 3138 32849
rect 3172 32815 3188 32849
rect 3122 32781 3188 32815
rect 3122 32747 3138 32781
rect 3172 32747 3188 32781
rect 3122 32713 3188 32747
rect 3122 32679 3138 32713
rect 3172 32679 3188 32713
rect 3122 32645 3188 32679
rect 3122 32611 3138 32645
rect 3172 32611 3188 32645
rect 3122 32594 3188 32611
rect 3218 32849 3284 32866
rect 3218 32815 3234 32849
rect 3268 32815 3284 32849
rect 3218 32781 3284 32815
rect 3218 32747 3234 32781
rect 3268 32747 3284 32781
rect 3218 32713 3284 32747
rect 3218 32679 3234 32713
rect 3268 32679 3284 32713
rect 3218 32645 3284 32679
rect 3218 32611 3234 32645
rect 3268 32611 3284 32645
rect 3218 32594 3284 32611
rect 3314 32849 3380 32866
rect 3314 32815 3330 32849
rect 3364 32815 3380 32849
rect 3314 32781 3380 32815
rect 3314 32747 3330 32781
rect 3364 32747 3380 32781
rect 3314 32713 3380 32747
rect 3314 32679 3330 32713
rect 3364 32679 3380 32713
rect 3314 32645 3380 32679
rect 3314 32611 3330 32645
rect 3364 32611 3380 32645
rect 3314 32594 3380 32611
rect 3410 32849 3472 32866
rect 3410 32815 3426 32849
rect 3460 32815 3472 32849
rect 3410 32781 3472 32815
rect 3410 32747 3426 32781
rect 3460 32747 3472 32781
rect 3410 32713 3472 32747
rect 3410 32679 3426 32713
rect 3460 32679 3472 32713
rect 3410 32645 3472 32679
rect 3410 32611 3426 32645
rect 3460 32611 3472 32645
rect 3410 32594 3472 32611
rect 3975 32849 4037 32866
rect 3975 32815 3987 32849
rect 4021 32815 4037 32849
rect 3975 32781 4037 32815
rect 3975 32747 3987 32781
rect 4021 32747 4037 32781
rect 3975 32713 4037 32747
rect 3975 32679 3987 32713
rect 4021 32679 4037 32713
rect 3975 32645 4037 32679
rect 3975 32611 3987 32645
rect 4021 32611 4037 32645
rect 3975 32594 4037 32611
rect 4067 32849 4133 32866
rect 4067 32815 4083 32849
rect 4117 32815 4133 32849
rect 4067 32781 4133 32815
rect 4067 32747 4083 32781
rect 4117 32747 4133 32781
rect 4067 32713 4133 32747
rect 4067 32679 4083 32713
rect 4117 32679 4133 32713
rect 4067 32645 4133 32679
rect 4067 32611 4083 32645
rect 4117 32611 4133 32645
rect 4067 32594 4133 32611
rect 4163 32849 4229 32866
rect 4163 32815 4179 32849
rect 4213 32815 4229 32849
rect 4163 32781 4229 32815
rect 4163 32747 4179 32781
rect 4213 32747 4229 32781
rect 4163 32713 4229 32747
rect 4163 32679 4179 32713
rect 4213 32679 4229 32713
rect 4163 32645 4229 32679
rect 4163 32611 4179 32645
rect 4213 32611 4229 32645
rect 4163 32594 4229 32611
rect 4259 32849 4325 32866
rect 4259 32815 4275 32849
rect 4309 32815 4325 32849
rect 4259 32781 4325 32815
rect 4259 32747 4275 32781
rect 4309 32747 4325 32781
rect 4259 32713 4325 32747
rect 4259 32679 4275 32713
rect 4309 32679 4325 32713
rect 4259 32645 4325 32679
rect 4259 32611 4275 32645
rect 4309 32611 4325 32645
rect 4259 32594 4325 32611
rect 4355 32849 4421 32866
rect 4355 32815 4371 32849
rect 4405 32815 4421 32849
rect 4355 32781 4421 32815
rect 4355 32747 4371 32781
rect 4405 32747 4421 32781
rect 4355 32713 4421 32747
rect 4355 32679 4371 32713
rect 4405 32679 4421 32713
rect 4355 32645 4421 32679
rect 4355 32611 4371 32645
rect 4405 32611 4421 32645
rect 4355 32594 4421 32611
rect 4451 32849 4517 32866
rect 4451 32815 4467 32849
rect 4501 32815 4517 32849
rect 4451 32781 4517 32815
rect 4451 32747 4467 32781
rect 4501 32747 4517 32781
rect 4451 32713 4517 32747
rect 4451 32679 4467 32713
rect 4501 32679 4517 32713
rect 4451 32645 4517 32679
rect 4451 32611 4467 32645
rect 4501 32611 4517 32645
rect 4451 32594 4517 32611
rect 4547 32849 4613 32866
rect 4547 32815 4563 32849
rect 4597 32815 4613 32849
rect 4547 32781 4613 32815
rect 4547 32747 4563 32781
rect 4597 32747 4613 32781
rect 4547 32713 4613 32747
rect 4547 32679 4563 32713
rect 4597 32679 4613 32713
rect 4547 32645 4613 32679
rect 4547 32611 4563 32645
rect 4597 32611 4613 32645
rect 4547 32594 4613 32611
rect 4643 32849 4709 32866
rect 4643 32815 4659 32849
rect 4693 32815 4709 32849
rect 4643 32781 4709 32815
rect 4643 32747 4659 32781
rect 4693 32747 4709 32781
rect 4643 32713 4709 32747
rect 4643 32679 4659 32713
rect 4693 32679 4709 32713
rect 4643 32645 4709 32679
rect 4643 32611 4659 32645
rect 4693 32611 4709 32645
rect 4643 32594 4709 32611
rect 4739 32849 4805 32866
rect 4739 32815 4755 32849
rect 4789 32815 4805 32849
rect 4739 32781 4805 32815
rect 4739 32747 4755 32781
rect 4789 32747 4805 32781
rect 4739 32713 4805 32747
rect 4739 32679 4755 32713
rect 4789 32679 4805 32713
rect 4739 32645 4805 32679
rect 4739 32611 4755 32645
rect 4789 32611 4805 32645
rect 4739 32594 4805 32611
rect 4835 32849 4901 32866
rect 4835 32815 4851 32849
rect 4885 32815 4901 32849
rect 4835 32781 4901 32815
rect 4835 32747 4851 32781
rect 4885 32747 4901 32781
rect 4835 32713 4901 32747
rect 4835 32679 4851 32713
rect 4885 32679 4901 32713
rect 4835 32645 4901 32679
rect 4835 32611 4851 32645
rect 4885 32611 4901 32645
rect 4835 32594 4901 32611
rect 4931 32849 4993 32866
rect 4931 32815 4947 32849
rect 4981 32815 4993 32849
rect 4931 32781 4993 32815
rect 4931 32747 4947 32781
rect 4981 32747 4993 32781
rect 4931 32713 4993 32747
rect 4931 32679 4947 32713
rect 4981 32679 4993 32713
rect 4931 32645 4993 32679
rect 4931 32611 4947 32645
rect 4981 32611 4993 32645
rect 4931 32594 4993 32611
rect 5348 32641 5400 32653
rect 5348 32607 5356 32641
rect 5390 32607 5400 32641
rect 5348 32573 5400 32607
rect 5348 32539 5356 32573
rect 5390 32539 5400 32573
rect 5348 32505 5400 32539
rect 5348 32471 5356 32505
rect 5390 32471 5400 32505
rect 5348 32453 5400 32471
rect 5430 32641 5482 32653
rect 5430 32607 5440 32641
rect 5474 32607 5482 32641
rect 5430 32573 5482 32607
rect 5430 32539 5440 32573
rect 5474 32539 5482 32573
rect 5430 32505 5482 32539
rect 5430 32471 5440 32505
rect 5474 32471 5482 32505
rect 5430 32453 5482 32471
rect 301 31558 363 31575
rect 301 31524 313 31558
rect 347 31524 363 31558
rect 301 31490 363 31524
rect 301 31456 313 31490
rect 347 31456 363 31490
rect 301 31422 363 31456
rect 301 31388 313 31422
rect 347 31388 363 31422
rect 301 31354 363 31388
rect 301 31320 313 31354
rect 347 31320 363 31354
rect 301 31303 363 31320
rect 393 31558 459 31575
rect 393 31524 409 31558
rect 443 31524 459 31558
rect 393 31490 459 31524
rect 393 31456 409 31490
rect 443 31456 459 31490
rect 393 31422 459 31456
rect 393 31388 409 31422
rect 443 31388 459 31422
rect 393 31354 459 31388
rect 393 31320 409 31354
rect 443 31320 459 31354
rect 393 31303 459 31320
rect 489 31558 555 31575
rect 489 31524 505 31558
rect 539 31524 555 31558
rect 489 31490 555 31524
rect 489 31456 505 31490
rect 539 31456 555 31490
rect 489 31422 555 31456
rect 489 31388 505 31422
rect 539 31388 555 31422
rect 489 31354 555 31388
rect 489 31320 505 31354
rect 539 31320 555 31354
rect 489 31303 555 31320
rect 585 31558 651 31575
rect 585 31524 601 31558
rect 635 31524 651 31558
rect 585 31490 651 31524
rect 585 31456 601 31490
rect 635 31456 651 31490
rect 585 31422 651 31456
rect 585 31388 601 31422
rect 635 31388 651 31422
rect 585 31354 651 31388
rect 585 31320 601 31354
rect 635 31320 651 31354
rect 585 31303 651 31320
rect 681 31558 747 31575
rect 681 31524 697 31558
rect 731 31524 747 31558
rect 681 31490 747 31524
rect 681 31456 697 31490
rect 731 31456 747 31490
rect 681 31422 747 31456
rect 681 31388 697 31422
rect 731 31388 747 31422
rect 681 31354 747 31388
rect 681 31320 697 31354
rect 731 31320 747 31354
rect 681 31303 747 31320
rect 777 31558 843 31575
rect 777 31524 793 31558
rect 827 31524 843 31558
rect 777 31490 843 31524
rect 777 31456 793 31490
rect 827 31456 843 31490
rect 777 31422 843 31456
rect 777 31388 793 31422
rect 827 31388 843 31422
rect 777 31354 843 31388
rect 777 31320 793 31354
rect 827 31320 843 31354
rect 777 31303 843 31320
rect 873 31558 939 31575
rect 873 31524 889 31558
rect 923 31524 939 31558
rect 873 31490 939 31524
rect 873 31456 889 31490
rect 923 31456 939 31490
rect 873 31422 939 31456
rect 873 31388 889 31422
rect 923 31388 939 31422
rect 873 31354 939 31388
rect 873 31320 889 31354
rect 923 31320 939 31354
rect 873 31303 939 31320
rect 969 31558 1035 31575
rect 969 31524 985 31558
rect 1019 31524 1035 31558
rect 969 31490 1035 31524
rect 969 31456 985 31490
rect 1019 31456 1035 31490
rect 969 31422 1035 31456
rect 969 31388 985 31422
rect 1019 31388 1035 31422
rect 969 31354 1035 31388
rect 969 31320 985 31354
rect 1019 31320 1035 31354
rect 969 31303 1035 31320
rect 1065 31558 1131 31575
rect 1065 31524 1081 31558
rect 1115 31524 1131 31558
rect 1065 31490 1131 31524
rect 1065 31456 1081 31490
rect 1115 31456 1131 31490
rect 1065 31422 1131 31456
rect 1065 31388 1081 31422
rect 1115 31388 1131 31422
rect 1065 31354 1131 31388
rect 1065 31320 1081 31354
rect 1115 31320 1131 31354
rect 1065 31303 1131 31320
rect 1161 31558 1227 31575
rect 1161 31524 1177 31558
rect 1211 31524 1227 31558
rect 1161 31490 1227 31524
rect 1161 31456 1177 31490
rect 1211 31456 1227 31490
rect 1161 31422 1227 31456
rect 1161 31388 1177 31422
rect 1211 31388 1227 31422
rect 1161 31354 1227 31388
rect 1161 31320 1177 31354
rect 1211 31320 1227 31354
rect 1161 31303 1227 31320
rect 1257 31558 1319 31575
rect 1257 31524 1273 31558
rect 1307 31524 1319 31558
rect 1257 31490 1319 31524
rect 1257 31456 1273 31490
rect 1307 31456 1319 31490
rect 1257 31422 1319 31456
rect 1257 31388 1273 31422
rect 1307 31388 1319 31422
rect 1257 31354 1319 31388
rect 1257 31320 1273 31354
rect 1307 31320 1319 31354
rect 1257 31303 1319 31320
rect 2454 31562 2516 31579
rect 2454 31528 2466 31562
rect 2500 31528 2516 31562
rect 2454 31494 2516 31528
rect 2454 31460 2466 31494
rect 2500 31460 2516 31494
rect 2454 31426 2516 31460
rect 2454 31392 2466 31426
rect 2500 31392 2516 31426
rect 2454 31358 2516 31392
rect 2454 31324 2466 31358
rect 2500 31324 2516 31358
rect 2454 31307 2516 31324
rect 2546 31562 2612 31579
rect 2546 31528 2562 31562
rect 2596 31528 2612 31562
rect 2546 31494 2612 31528
rect 2546 31460 2562 31494
rect 2596 31460 2612 31494
rect 2546 31426 2612 31460
rect 2546 31392 2562 31426
rect 2596 31392 2612 31426
rect 2546 31358 2612 31392
rect 2546 31324 2562 31358
rect 2596 31324 2612 31358
rect 2546 31307 2612 31324
rect 2642 31562 2708 31579
rect 2642 31528 2658 31562
rect 2692 31528 2708 31562
rect 2642 31494 2708 31528
rect 2642 31460 2658 31494
rect 2692 31460 2708 31494
rect 2642 31426 2708 31460
rect 2642 31392 2658 31426
rect 2692 31392 2708 31426
rect 2642 31358 2708 31392
rect 2642 31324 2658 31358
rect 2692 31324 2708 31358
rect 2642 31307 2708 31324
rect 2738 31562 2804 31579
rect 2738 31528 2754 31562
rect 2788 31528 2804 31562
rect 2738 31494 2804 31528
rect 2738 31460 2754 31494
rect 2788 31460 2804 31494
rect 2738 31426 2804 31460
rect 2738 31392 2754 31426
rect 2788 31392 2804 31426
rect 2738 31358 2804 31392
rect 2738 31324 2754 31358
rect 2788 31324 2804 31358
rect 2738 31307 2804 31324
rect 2834 31562 2900 31579
rect 2834 31528 2850 31562
rect 2884 31528 2900 31562
rect 2834 31494 2900 31528
rect 2834 31460 2850 31494
rect 2884 31460 2900 31494
rect 2834 31426 2900 31460
rect 2834 31392 2850 31426
rect 2884 31392 2900 31426
rect 2834 31358 2900 31392
rect 2834 31324 2850 31358
rect 2884 31324 2900 31358
rect 2834 31307 2900 31324
rect 2930 31562 2996 31579
rect 2930 31528 2946 31562
rect 2980 31528 2996 31562
rect 2930 31494 2996 31528
rect 2930 31460 2946 31494
rect 2980 31460 2996 31494
rect 2930 31426 2996 31460
rect 2930 31392 2946 31426
rect 2980 31392 2996 31426
rect 2930 31358 2996 31392
rect 2930 31324 2946 31358
rect 2980 31324 2996 31358
rect 2930 31307 2996 31324
rect 3026 31562 3092 31579
rect 3026 31528 3042 31562
rect 3076 31528 3092 31562
rect 3026 31494 3092 31528
rect 3026 31460 3042 31494
rect 3076 31460 3092 31494
rect 3026 31426 3092 31460
rect 3026 31392 3042 31426
rect 3076 31392 3092 31426
rect 3026 31358 3092 31392
rect 3026 31324 3042 31358
rect 3076 31324 3092 31358
rect 3026 31307 3092 31324
rect 3122 31562 3188 31579
rect 3122 31528 3138 31562
rect 3172 31528 3188 31562
rect 3122 31494 3188 31528
rect 3122 31460 3138 31494
rect 3172 31460 3188 31494
rect 3122 31426 3188 31460
rect 3122 31392 3138 31426
rect 3172 31392 3188 31426
rect 3122 31358 3188 31392
rect 3122 31324 3138 31358
rect 3172 31324 3188 31358
rect 3122 31307 3188 31324
rect 3218 31562 3284 31579
rect 3218 31528 3234 31562
rect 3268 31528 3284 31562
rect 3218 31494 3284 31528
rect 3218 31460 3234 31494
rect 3268 31460 3284 31494
rect 3218 31426 3284 31460
rect 3218 31392 3234 31426
rect 3268 31392 3284 31426
rect 3218 31358 3284 31392
rect 3218 31324 3234 31358
rect 3268 31324 3284 31358
rect 3218 31307 3284 31324
rect 3314 31562 3380 31579
rect 3314 31528 3330 31562
rect 3364 31528 3380 31562
rect 3314 31494 3380 31528
rect 3314 31460 3330 31494
rect 3364 31460 3380 31494
rect 3314 31426 3380 31460
rect 3314 31392 3330 31426
rect 3364 31392 3380 31426
rect 3314 31358 3380 31392
rect 3314 31324 3330 31358
rect 3364 31324 3380 31358
rect 3314 31307 3380 31324
rect 3410 31562 3472 31579
rect 3410 31528 3426 31562
rect 3460 31528 3472 31562
rect 3410 31494 3472 31528
rect 3410 31460 3426 31494
rect 3460 31460 3472 31494
rect 3410 31426 3472 31460
rect 3410 31392 3426 31426
rect 3460 31392 3472 31426
rect 3410 31358 3472 31392
rect 3410 31324 3426 31358
rect 3460 31324 3472 31358
rect 3410 31307 3472 31324
rect 3975 31562 4037 31579
rect 3975 31528 3987 31562
rect 4021 31528 4037 31562
rect 3975 31494 4037 31528
rect 3975 31460 3987 31494
rect 4021 31460 4037 31494
rect 3975 31426 4037 31460
rect 3975 31392 3987 31426
rect 4021 31392 4037 31426
rect 3975 31358 4037 31392
rect 3975 31324 3987 31358
rect 4021 31324 4037 31358
rect 3975 31307 4037 31324
rect 4067 31562 4133 31579
rect 4067 31528 4083 31562
rect 4117 31528 4133 31562
rect 4067 31494 4133 31528
rect 4067 31460 4083 31494
rect 4117 31460 4133 31494
rect 4067 31426 4133 31460
rect 4067 31392 4083 31426
rect 4117 31392 4133 31426
rect 4067 31358 4133 31392
rect 4067 31324 4083 31358
rect 4117 31324 4133 31358
rect 4067 31307 4133 31324
rect 4163 31562 4229 31579
rect 4163 31528 4179 31562
rect 4213 31528 4229 31562
rect 4163 31494 4229 31528
rect 4163 31460 4179 31494
rect 4213 31460 4229 31494
rect 4163 31426 4229 31460
rect 4163 31392 4179 31426
rect 4213 31392 4229 31426
rect 4163 31358 4229 31392
rect 4163 31324 4179 31358
rect 4213 31324 4229 31358
rect 4163 31307 4229 31324
rect 4259 31562 4325 31579
rect 4259 31528 4275 31562
rect 4309 31528 4325 31562
rect 4259 31494 4325 31528
rect 4259 31460 4275 31494
rect 4309 31460 4325 31494
rect 4259 31426 4325 31460
rect 4259 31392 4275 31426
rect 4309 31392 4325 31426
rect 4259 31358 4325 31392
rect 4259 31324 4275 31358
rect 4309 31324 4325 31358
rect 4259 31307 4325 31324
rect 4355 31562 4421 31579
rect 4355 31528 4371 31562
rect 4405 31528 4421 31562
rect 4355 31494 4421 31528
rect 4355 31460 4371 31494
rect 4405 31460 4421 31494
rect 4355 31426 4421 31460
rect 4355 31392 4371 31426
rect 4405 31392 4421 31426
rect 4355 31358 4421 31392
rect 4355 31324 4371 31358
rect 4405 31324 4421 31358
rect 4355 31307 4421 31324
rect 4451 31562 4517 31579
rect 4451 31528 4467 31562
rect 4501 31528 4517 31562
rect 4451 31494 4517 31528
rect 4451 31460 4467 31494
rect 4501 31460 4517 31494
rect 4451 31426 4517 31460
rect 4451 31392 4467 31426
rect 4501 31392 4517 31426
rect 4451 31358 4517 31392
rect 4451 31324 4467 31358
rect 4501 31324 4517 31358
rect 4451 31307 4517 31324
rect 4547 31562 4613 31579
rect 4547 31528 4563 31562
rect 4597 31528 4613 31562
rect 4547 31494 4613 31528
rect 4547 31460 4563 31494
rect 4597 31460 4613 31494
rect 4547 31426 4613 31460
rect 4547 31392 4563 31426
rect 4597 31392 4613 31426
rect 4547 31358 4613 31392
rect 4547 31324 4563 31358
rect 4597 31324 4613 31358
rect 4547 31307 4613 31324
rect 4643 31562 4709 31579
rect 4643 31528 4659 31562
rect 4693 31528 4709 31562
rect 4643 31494 4709 31528
rect 4643 31460 4659 31494
rect 4693 31460 4709 31494
rect 4643 31426 4709 31460
rect 4643 31392 4659 31426
rect 4693 31392 4709 31426
rect 4643 31358 4709 31392
rect 4643 31324 4659 31358
rect 4693 31324 4709 31358
rect 4643 31307 4709 31324
rect 4739 31562 4805 31579
rect 4739 31528 4755 31562
rect 4789 31528 4805 31562
rect 4739 31494 4805 31528
rect 4739 31460 4755 31494
rect 4789 31460 4805 31494
rect 4739 31426 4805 31460
rect 4739 31392 4755 31426
rect 4789 31392 4805 31426
rect 4739 31358 4805 31392
rect 4739 31324 4755 31358
rect 4789 31324 4805 31358
rect 4739 31307 4805 31324
rect 4835 31562 4901 31579
rect 4835 31528 4851 31562
rect 4885 31528 4901 31562
rect 4835 31494 4901 31528
rect 4835 31460 4851 31494
rect 4885 31460 4901 31494
rect 4835 31426 4901 31460
rect 4835 31392 4851 31426
rect 4885 31392 4901 31426
rect 4835 31358 4901 31392
rect 4835 31324 4851 31358
rect 4885 31324 4901 31358
rect 4835 31307 4901 31324
rect 4931 31562 4993 31579
rect 4931 31528 4947 31562
rect 4981 31528 4993 31562
rect 4931 31494 4993 31528
rect 4931 31460 4947 31494
rect 4981 31460 4993 31494
rect 4931 31426 4993 31460
rect 4931 31392 4947 31426
rect 4981 31392 4993 31426
rect 4931 31358 4993 31392
rect 4931 31324 4947 31358
rect 4981 31324 4993 31358
rect 4931 31307 4993 31324
rect 5348 31354 5400 31366
rect 5348 31320 5356 31354
rect 5390 31320 5400 31354
rect 5348 31286 5400 31320
rect 5348 31252 5356 31286
rect 5390 31252 5400 31286
rect 5348 31218 5400 31252
rect 5348 31184 5356 31218
rect 5390 31184 5400 31218
rect 5348 31166 5400 31184
rect 5430 31354 5482 31366
rect 5430 31320 5440 31354
rect 5474 31320 5482 31354
rect 5430 31286 5482 31320
rect 5430 31252 5440 31286
rect 5474 31252 5482 31286
rect 5430 31218 5482 31252
rect 5430 31184 5440 31218
rect 5474 31184 5482 31218
rect 5430 31166 5482 31184
rect 301 30271 363 30288
rect 301 30237 313 30271
rect 347 30237 363 30271
rect 301 30203 363 30237
rect 301 30169 313 30203
rect 347 30169 363 30203
rect 301 30135 363 30169
rect 301 30101 313 30135
rect 347 30101 363 30135
rect 301 30067 363 30101
rect 301 30033 313 30067
rect 347 30033 363 30067
rect 301 30016 363 30033
rect 393 30271 459 30288
rect 393 30237 409 30271
rect 443 30237 459 30271
rect 393 30203 459 30237
rect 393 30169 409 30203
rect 443 30169 459 30203
rect 393 30135 459 30169
rect 393 30101 409 30135
rect 443 30101 459 30135
rect 393 30067 459 30101
rect 393 30033 409 30067
rect 443 30033 459 30067
rect 393 30016 459 30033
rect 489 30271 555 30288
rect 489 30237 505 30271
rect 539 30237 555 30271
rect 489 30203 555 30237
rect 489 30169 505 30203
rect 539 30169 555 30203
rect 489 30135 555 30169
rect 489 30101 505 30135
rect 539 30101 555 30135
rect 489 30067 555 30101
rect 489 30033 505 30067
rect 539 30033 555 30067
rect 489 30016 555 30033
rect 585 30271 651 30288
rect 585 30237 601 30271
rect 635 30237 651 30271
rect 585 30203 651 30237
rect 585 30169 601 30203
rect 635 30169 651 30203
rect 585 30135 651 30169
rect 585 30101 601 30135
rect 635 30101 651 30135
rect 585 30067 651 30101
rect 585 30033 601 30067
rect 635 30033 651 30067
rect 585 30016 651 30033
rect 681 30271 747 30288
rect 681 30237 697 30271
rect 731 30237 747 30271
rect 681 30203 747 30237
rect 681 30169 697 30203
rect 731 30169 747 30203
rect 681 30135 747 30169
rect 681 30101 697 30135
rect 731 30101 747 30135
rect 681 30067 747 30101
rect 681 30033 697 30067
rect 731 30033 747 30067
rect 681 30016 747 30033
rect 777 30271 843 30288
rect 777 30237 793 30271
rect 827 30237 843 30271
rect 777 30203 843 30237
rect 777 30169 793 30203
rect 827 30169 843 30203
rect 777 30135 843 30169
rect 777 30101 793 30135
rect 827 30101 843 30135
rect 777 30067 843 30101
rect 777 30033 793 30067
rect 827 30033 843 30067
rect 777 30016 843 30033
rect 873 30271 939 30288
rect 873 30237 889 30271
rect 923 30237 939 30271
rect 873 30203 939 30237
rect 873 30169 889 30203
rect 923 30169 939 30203
rect 873 30135 939 30169
rect 873 30101 889 30135
rect 923 30101 939 30135
rect 873 30067 939 30101
rect 873 30033 889 30067
rect 923 30033 939 30067
rect 873 30016 939 30033
rect 969 30271 1035 30288
rect 969 30237 985 30271
rect 1019 30237 1035 30271
rect 969 30203 1035 30237
rect 969 30169 985 30203
rect 1019 30169 1035 30203
rect 969 30135 1035 30169
rect 969 30101 985 30135
rect 1019 30101 1035 30135
rect 969 30067 1035 30101
rect 969 30033 985 30067
rect 1019 30033 1035 30067
rect 969 30016 1035 30033
rect 1065 30271 1131 30288
rect 1065 30237 1081 30271
rect 1115 30237 1131 30271
rect 1065 30203 1131 30237
rect 1065 30169 1081 30203
rect 1115 30169 1131 30203
rect 1065 30135 1131 30169
rect 1065 30101 1081 30135
rect 1115 30101 1131 30135
rect 1065 30067 1131 30101
rect 1065 30033 1081 30067
rect 1115 30033 1131 30067
rect 1065 30016 1131 30033
rect 1161 30271 1227 30288
rect 1161 30237 1177 30271
rect 1211 30237 1227 30271
rect 1161 30203 1227 30237
rect 1161 30169 1177 30203
rect 1211 30169 1227 30203
rect 1161 30135 1227 30169
rect 1161 30101 1177 30135
rect 1211 30101 1227 30135
rect 1161 30067 1227 30101
rect 1161 30033 1177 30067
rect 1211 30033 1227 30067
rect 1161 30016 1227 30033
rect 1257 30271 1319 30288
rect 1257 30237 1273 30271
rect 1307 30237 1319 30271
rect 1257 30203 1319 30237
rect 1257 30169 1273 30203
rect 1307 30169 1319 30203
rect 1257 30135 1319 30169
rect 1257 30101 1273 30135
rect 1307 30101 1319 30135
rect 1257 30067 1319 30101
rect 1257 30033 1273 30067
rect 1307 30033 1319 30067
rect 1257 30016 1319 30033
rect 2454 30275 2516 30292
rect 2454 30241 2466 30275
rect 2500 30241 2516 30275
rect 2454 30207 2516 30241
rect 2454 30173 2466 30207
rect 2500 30173 2516 30207
rect 2454 30139 2516 30173
rect 2454 30105 2466 30139
rect 2500 30105 2516 30139
rect 2454 30071 2516 30105
rect 2454 30037 2466 30071
rect 2500 30037 2516 30071
rect 2454 30020 2516 30037
rect 2546 30275 2612 30292
rect 2546 30241 2562 30275
rect 2596 30241 2612 30275
rect 2546 30207 2612 30241
rect 2546 30173 2562 30207
rect 2596 30173 2612 30207
rect 2546 30139 2612 30173
rect 2546 30105 2562 30139
rect 2596 30105 2612 30139
rect 2546 30071 2612 30105
rect 2546 30037 2562 30071
rect 2596 30037 2612 30071
rect 2546 30020 2612 30037
rect 2642 30275 2708 30292
rect 2642 30241 2658 30275
rect 2692 30241 2708 30275
rect 2642 30207 2708 30241
rect 2642 30173 2658 30207
rect 2692 30173 2708 30207
rect 2642 30139 2708 30173
rect 2642 30105 2658 30139
rect 2692 30105 2708 30139
rect 2642 30071 2708 30105
rect 2642 30037 2658 30071
rect 2692 30037 2708 30071
rect 2642 30020 2708 30037
rect 2738 30275 2804 30292
rect 2738 30241 2754 30275
rect 2788 30241 2804 30275
rect 2738 30207 2804 30241
rect 2738 30173 2754 30207
rect 2788 30173 2804 30207
rect 2738 30139 2804 30173
rect 2738 30105 2754 30139
rect 2788 30105 2804 30139
rect 2738 30071 2804 30105
rect 2738 30037 2754 30071
rect 2788 30037 2804 30071
rect 2738 30020 2804 30037
rect 2834 30275 2900 30292
rect 2834 30241 2850 30275
rect 2884 30241 2900 30275
rect 2834 30207 2900 30241
rect 2834 30173 2850 30207
rect 2884 30173 2900 30207
rect 2834 30139 2900 30173
rect 2834 30105 2850 30139
rect 2884 30105 2900 30139
rect 2834 30071 2900 30105
rect 2834 30037 2850 30071
rect 2884 30037 2900 30071
rect 2834 30020 2900 30037
rect 2930 30275 2996 30292
rect 2930 30241 2946 30275
rect 2980 30241 2996 30275
rect 2930 30207 2996 30241
rect 2930 30173 2946 30207
rect 2980 30173 2996 30207
rect 2930 30139 2996 30173
rect 2930 30105 2946 30139
rect 2980 30105 2996 30139
rect 2930 30071 2996 30105
rect 2930 30037 2946 30071
rect 2980 30037 2996 30071
rect 2930 30020 2996 30037
rect 3026 30275 3092 30292
rect 3026 30241 3042 30275
rect 3076 30241 3092 30275
rect 3026 30207 3092 30241
rect 3026 30173 3042 30207
rect 3076 30173 3092 30207
rect 3026 30139 3092 30173
rect 3026 30105 3042 30139
rect 3076 30105 3092 30139
rect 3026 30071 3092 30105
rect 3026 30037 3042 30071
rect 3076 30037 3092 30071
rect 3026 30020 3092 30037
rect 3122 30275 3188 30292
rect 3122 30241 3138 30275
rect 3172 30241 3188 30275
rect 3122 30207 3188 30241
rect 3122 30173 3138 30207
rect 3172 30173 3188 30207
rect 3122 30139 3188 30173
rect 3122 30105 3138 30139
rect 3172 30105 3188 30139
rect 3122 30071 3188 30105
rect 3122 30037 3138 30071
rect 3172 30037 3188 30071
rect 3122 30020 3188 30037
rect 3218 30275 3284 30292
rect 3218 30241 3234 30275
rect 3268 30241 3284 30275
rect 3218 30207 3284 30241
rect 3218 30173 3234 30207
rect 3268 30173 3284 30207
rect 3218 30139 3284 30173
rect 3218 30105 3234 30139
rect 3268 30105 3284 30139
rect 3218 30071 3284 30105
rect 3218 30037 3234 30071
rect 3268 30037 3284 30071
rect 3218 30020 3284 30037
rect 3314 30275 3380 30292
rect 3314 30241 3330 30275
rect 3364 30241 3380 30275
rect 3314 30207 3380 30241
rect 3314 30173 3330 30207
rect 3364 30173 3380 30207
rect 3314 30139 3380 30173
rect 3314 30105 3330 30139
rect 3364 30105 3380 30139
rect 3314 30071 3380 30105
rect 3314 30037 3330 30071
rect 3364 30037 3380 30071
rect 3314 30020 3380 30037
rect 3410 30275 3472 30292
rect 3410 30241 3426 30275
rect 3460 30241 3472 30275
rect 3410 30207 3472 30241
rect 3410 30173 3426 30207
rect 3460 30173 3472 30207
rect 3410 30139 3472 30173
rect 3410 30105 3426 30139
rect 3460 30105 3472 30139
rect 3410 30071 3472 30105
rect 3410 30037 3426 30071
rect 3460 30037 3472 30071
rect 3410 30020 3472 30037
rect 3975 30275 4037 30292
rect 3975 30241 3987 30275
rect 4021 30241 4037 30275
rect 3975 30207 4037 30241
rect 3975 30173 3987 30207
rect 4021 30173 4037 30207
rect 3975 30139 4037 30173
rect 3975 30105 3987 30139
rect 4021 30105 4037 30139
rect 3975 30071 4037 30105
rect 3975 30037 3987 30071
rect 4021 30037 4037 30071
rect 3975 30020 4037 30037
rect 4067 30275 4133 30292
rect 4067 30241 4083 30275
rect 4117 30241 4133 30275
rect 4067 30207 4133 30241
rect 4067 30173 4083 30207
rect 4117 30173 4133 30207
rect 4067 30139 4133 30173
rect 4067 30105 4083 30139
rect 4117 30105 4133 30139
rect 4067 30071 4133 30105
rect 4067 30037 4083 30071
rect 4117 30037 4133 30071
rect 4067 30020 4133 30037
rect 4163 30275 4229 30292
rect 4163 30241 4179 30275
rect 4213 30241 4229 30275
rect 4163 30207 4229 30241
rect 4163 30173 4179 30207
rect 4213 30173 4229 30207
rect 4163 30139 4229 30173
rect 4163 30105 4179 30139
rect 4213 30105 4229 30139
rect 4163 30071 4229 30105
rect 4163 30037 4179 30071
rect 4213 30037 4229 30071
rect 4163 30020 4229 30037
rect 4259 30275 4325 30292
rect 4259 30241 4275 30275
rect 4309 30241 4325 30275
rect 4259 30207 4325 30241
rect 4259 30173 4275 30207
rect 4309 30173 4325 30207
rect 4259 30139 4325 30173
rect 4259 30105 4275 30139
rect 4309 30105 4325 30139
rect 4259 30071 4325 30105
rect 4259 30037 4275 30071
rect 4309 30037 4325 30071
rect 4259 30020 4325 30037
rect 4355 30275 4421 30292
rect 4355 30241 4371 30275
rect 4405 30241 4421 30275
rect 4355 30207 4421 30241
rect 4355 30173 4371 30207
rect 4405 30173 4421 30207
rect 4355 30139 4421 30173
rect 4355 30105 4371 30139
rect 4405 30105 4421 30139
rect 4355 30071 4421 30105
rect 4355 30037 4371 30071
rect 4405 30037 4421 30071
rect 4355 30020 4421 30037
rect 4451 30275 4517 30292
rect 4451 30241 4467 30275
rect 4501 30241 4517 30275
rect 4451 30207 4517 30241
rect 4451 30173 4467 30207
rect 4501 30173 4517 30207
rect 4451 30139 4517 30173
rect 4451 30105 4467 30139
rect 4501 30105 4517 30139
rect 4451 30071 4517 30105
rect 4451 30037 4467 30071
rect 4501 30037 4517 30071
rect 4451 30020 4517 30037
rect 4547 30275 4613 30292
rect 4547 30241 4563 30275
rect 4597 30241 4613 30275
rect 4547 30207 4613 30241
rect 4547 30173 4563 30207
rect 4597 30173 4613 30207
rect 4547 30139 4613 30173
rect 4547 30105 4563 30139
rect 4597 30105 4613 30139
rect 4547 30071 4613 30105
rect 4547 30037 4563 30071
rect 4597 30037 4613 30071
rect 4547 30020 4613 30037
rect 4643 30275 4709 30292
rect 4643 30241 4659 30275
rect 4693 30241 4709 30275
rect 4643 30207 4709 30241
rect 4643 30173 4659 30207
rect 4693 30173 4709 30207
rect 4643 30139 4709 30173
rect 4643 30105 4659 30139
rect 4693 30105 4709 30139
rect 4643 30071 4709 30105
rect 4643 30037 4659 30071
rect 4693 30037 4709 30071
rect 4643 30020 4709 30037
rect 4739 30275 4805 30292
rect 4739 30241 4755 30275
rect 4789 30241 4805 30275
rect 4739 30207 4805 30241
rect 4739 30173 4755 30207
rect 4789 30173 4805 30207
rect 4739 30139 4805 30173
rect 4739 30105 4755 30139
rect 4789 30105 4805 30139
rect 4739 30071 4805 30105
rect 4739 30037 4755 30071
rect 4789 30037 4805 30071
rect 4739 30020 4805 30037
rect 4835 30275 4901 30292
rect 4835 30241 4851 30275
rect 4885 30241 4901 30275
rect 4835 30207 4901 30241
rect 4835 30173 4851 30207
rect 4885 30173 4901 30207
rect 4835 30139 4901 30173
rect 4835 30105 4851 30139
rect 4885 30105 4901 30139
rect 4835 30071 4901 30105
rect 4835 30037 4851 30071
rect 4885 30037 4901 30071
rect 4835 30020 4901 30037
rect 4931 30275 4993 30292
rect 4931 30241 4947 30275
rect 4981 30241 4993 30275
rect 4931 30207 4993 30241
rect 4931 30173 4947 30207
rect 4981 30173 4993 30207
rect 4931 30139 4993 30173
rect 4931 30105 4947 30139
rect 4981 30105 4993 30139
rect 4931 30071 4993 30105
rect 4931 30037 4947 30071
rect 4981 30037 4993 30071
rect 4931 30020 4993 30037
rect 5348 30067 5400 30079
rect 5348 30033 5356 30067
rect 5390 30033 5400 30067
rect 5348 29999 5400 30033
rect 5348 29965 5356 29999
rect 5390 29965 5400 29999
rect 5348 29931 5400 29965
rect 5348 29897 5356 29931
rect 5390 29897 5400 29931
rect 5348 29879 5400 29897
rect 5430 30067 5482 30079
rect 5430 30033 5440 30067
rect 5474 30033 5482 30067
rect 5430 29999 5482 30033
rect 5430 29965 5440 29999
rect 5474 29965 5482 29999
rect 5430 29931 5482 29965
rect 5430 29897 5440 29931
rect 5474 29897 5482 29931
rect 5430 29879 5482 29897
rect 301 28984 363 29001
rect 301 28950 313 28984
rect 347 28950 363 28984
rect 301 28916 363 28950
rect 301 28882 313 28916
rect 347 28882 363 28916
rect 301 28848 363 28882
rect 301 28814 313 28848
rect 347 28814 363 28848
rect 301 28780 363 28814
rect 301 28746 313 28780
rect 347 28746 363 28780
rect 301 28729 363 28746
rect 393 28984 459 29001
rect 393 28950 409 28984
rect 443 28950 459 28984
rect 393 28916 459 28950
rect 393 28882 409 28916
rect 443 28882 459 28916
rect 393 28848 459 28882
rect 393 28814 409 28848
rect 443 28814 459 28848
rect 393 28780 459 28814
rect 393 28746 409 28780
rect 443 28746 459 28780
rect 393 28729 459 28746
rect 489 28984 555 29001
rect 489 28950 505 28984
rect 539 28950 555 28984
rect 489 28916 555 28950
rect 489 28882 505 28916
rect 539 28882 555 28916
rect 489 28848 555 28882
rect 489 28814 505 28848
rect 539 28814 555 28848
rect 489 28780 555 28814
rect 489 28746 505 28780
rect 539 28746 555 28780
rect 489 28729 555 28746
rect 585 28984 651 29001
rect 585 28950 601 28984
rect 635 28950 651 28984
rect 585 28916 651 28950
rect 585 28882 601 28916
rect 635 28882 651 28916
rect 585 28848 651 28882
rect 585 28814 601 28848
rect 635 28814 651 28848
rect 585 28780 651 28814
rect 585 28746 601 28780
rect 635 28746 651 28780
rect 585 28729 651 28746
rect 681 28984 747 29001
rect 681 28950 697 28984
rect 731 28950 747 28984
rect 681 28916 747 28950
rect 681 28882 697 28916
rect 731 28882 747 28916
rect 681 28848 747 28882
rect 681 28814 697 28848
rect 731 28814 747 28848
rect 681 28780 747 28814
rect 681 28746 697 28780
rect 731 28746 747 28780
rect 681 28729 747 28746
rect 777 28984 843 29001
rect 777 28950 793 28984
rect 827 28950 843 28984
rect 777 28916 843 28950
rect 777 28882 793 28916
rect 827 28882 843 28916
rect 777 28848 843 28882
rect 777 28814 793 28848
rect 827 28814 843 28848
rect 777 28780 843 28814
rect 777 28746 793 28780
rect 827 28746 843 28780
rect 777 28729 843 28746
rect 873 28984 939 29001
rect 873 28950 889 28984
rect 923 28950 939 28984
rect 873 28916 939 28950
rect 873 28882 889 28916
rect 923 28882 939 28916
rect 873 28848 939 28882
rect 873 28814 889 28848
rect 923 28814 939 28848
rect 873 28780 939 28814
rect 873 28746 889 28780
rect 923 28746 939 28780
rect 873 28729 939 28746
rect 969 28984 1035 29001
rect 969 28950 985 28984
rect 1019 28950 1035 28984
rect 969 28916 1035 28950
rect 969 28882 985 28916
rect 1019 28882 1035 28916
rect 969 28848 1035 28882
rect 969 28814 985 28848
rect 1019 28814 1035 28848
rect 969 28780 1035 28814
rect 969 28746 985 28780
rect 1019 28746 1035 28780
rect 969 28729 1035 28746
rect 1065 28984 1131 29001
rect 1065 28950 1081 28984
rect 1115 28950 1131 28984
rect 1065 28916 1131 28950
rect 1065 28882 1081 28916
rect 1115 28882 1131 28916
rect 1065 28848 1131 28882
rect 1065 28814 1081 28848
rect 1115 28814 1131 28848
rect 1065 28780 1131 28814
rect 1065 28746 1081 28780
rect 1115 28746 1131 28780
rect 1065 28729 1131 28746
rect 1161 28984 1227 29001
rect 1161 28950 1177 28984
rect 1211 28950 1227 28984
rect 1161 28916 1227 28950
rect 1161 28882 1177 28916
rect 1211 28882 1227 28916
rect 1161 28848 1227 28882
rect 1161 28814 1177 28848
rect 1211 28814 1227 28848
rect 1161 28780 1227 28814
rect 1161 28746 1177 28780
rect 1211 28746 1227 28780
rect 1161 28729 1227 28746
rect 1257 28984 1319 29001
rect 1257 28950 1273 28984
rect 1307 28950 1319 28984
rect 1257 28916 1319 28950
rect 1257 28882 1273 28916
rect 1307 28882 1319 28916
rect 1257 28848 1319 28882
rect 1257 28814 1273 28848
rect 1307 28814 1319 28848
rect 1257 28780 1319 28814
rect 1257 28746 1273 28780
rect 1307 28746 1319 28780
rect 1257 28729 1319 28746
rect 2454 28988 2516 29005
rect 2454 28954 2466 28988
rect 2500 28954 2516 28988
rect 2454 28920 2516 28954
rect 2454 28886 2466 28920
rect 2500 28886 2516 28920
rect 2454 28852 2516 28886
rect 2454 28818 2466 28852
rect 2500 28818 2516 28852
rect 2454 28784 2516 28818
rect 2454 28750 2466 28784
rect 2500 28750 2516 28784
rect 2454 28733 2516 28750
rect 2546 28988 2612 29005
rect 2546 28954 2562 28988
rect 2596 28954 2612 28988
rect 2546 28920 2612 28954
rect 2546 28886 2562 28920
rect 2596 28886 2612 28920
rect 2546 28852 2612 28886
rect 2546 28818 2562 28852
rect 2596 28818 2612 28852
rect 2546 28784 2612 28818
rect 2546 28750 2562 28784
rect 2596 28750 2612 28784
rect 2546 28733 2612 28750
rect 2642 28988 2708 29005
rect 2642 28954 2658 28988
rect 2692 28954 2708 28988
rect 2642 28920 2708 28954
rect 2642 28886 2658 28920
rect 2692 28886 2708 28920
rect 2642 28852 2708 28886
rect 2642 28818 2658 28852
rect 2692 28818 2708 28852
rect 2642 28784 2708 28818
rect 2642 28750 2658 28784
rect 2692 28750 2708 28784
rect 2642 28733 2708 28750
rect 2738 28988 2804 29005
rect 2738 28954 2754 28988
rect 2788 28954 2804 28988
rect 2738 28920 2804 28954
rect 2738 28886 2754 28920
rect 2788 28886 2804 28920
rect 2738 28852 2804 28886
rect 2738 28818 2754 28852
rect 2788 28818 2804 28852
rect 2738 28784 2804 28818
rect 2738 28750 2754 28784
rect 2788 28750 2804 28784
rect 2738 28733 2804 28750
rect 2834 28988 2900 29005
rect 2834 28954 2850 28988
rect 2884 28954 2900 28988
rect 2834 28920 2900 28954
rect 2834 28886 2850 28920
rect 2884 28886 2900 28920
rect 2834 28852 2900 28886
rect 2834 28818 2850 28852
rect 2884 28818 2900 28852
rect 2834 28784 2900 28818
rect 2834 28750 2850 28784
rect 2884 28750 2900 28784
rect 2834 28733 2900 28750
rect 2930 28988 2996 29005
rect 2930 28954 2946 28988
rect 2980 28954 2996 28988
rect 2930 28920 2996 28954
rect 2930 28886 2946 28920
rect 2980 28886 2996 28920
rect 2930 28852 2996 28886
rect 2930 28818 2946 28852
rect 2980 28818 2996 28852
rect 2930 28784 2996 28818
rect 2930 28750 2946 28784
rect 2980 28750 2996 28784
rect 2930 28733 2996 28750
rect 3026 28988 3092 29005
rect 3026 28954 3042 28988
rect 3076 28954 3092 28988
rect 3026 28920 3092 28954
rect 3026 28886 3042 28920
rect 3076 28886 3092 28920
rect 3026 28852 3092 28886
rect 3026 28818 3042 28852
rect 3076 28818 3092 28852
rect 3026 28784 3092 28818
rect 3026 28750 3042 28784
rect 3076 28750 3092 28784
rect 3026 28733 3092 28750
rect 3122 28988 3188 29005
rect 3122 28954 3138 28988
rect 3172 28954 3188 28988
rect 3122 28920 3188 28954
rect 3122 28886 3138 28920
rect 3172 28886 3188 28920
rect 3122 28852 3188 28886
rect 3122 28818 3138 28852
rect 3172 28818 3188 28852
rect 3122 28784 3188 28818
rect 3122 28750 3138 28784
rect 3172 28750 3188 28784
rect 3122 28733 3188 28750
rect 3218 28988 3284 29005
rect 3218 28954 3234 28988
rect 3268 28954 3284 28988
rect 3218 28920 3284 28954
rect 3218 28886 3234 28920
rect 3268 28886 3284 28920
rect 3218 28852 3284 28886
rect 3218 28818 3234 28852
rect 3268 28818 3284 28852
rect 3218 28784 3284 28818
rect 3218 28750 3234 28784
rect 3268 28750 3284 28784
rect 3218 28733 3284 28750
rect 3314 28988 3380 29005
rect 3314 28954 3330 28988
rect 3364 28954 3380 28988
rect 3314 28920 3380 28954
rect 3314 28886 3330 28920
rect 3364 28886 3380 28920
rect 3314 28852 3380 28886
rect 3314 28818 3330 28852
rect 3364 28818 3380 28852
rect 3314 28784 3380 28818
rect 3314 28750 3330 28784
rect 3364 28750 3380 28784
rect 3314 28733 3380 28750
rect 3410 28988 3472 29005
rect 3410 28954 3426 28988
rect 3460 28954 3472 28988
rect 3410 28920 3472 28954
rect 3410 28886 3426 28920
rect 3460 28886 3472 28920
rect 3410 28852 3472 28886
rect 3410 28818 3426 28852
rect 3460 28818 3472 28852
rect 3410 28784 3472 28818
rect 3410 28750 3426 28784
rect 3460 28750 3472 28784
rect 3410 28733 3472 28750
rect 3975 28988 4037 29005
rect 3975 28954 3987 28988
rect 4021 28954 4037 28988
rect 3975 28920 4037 28954
rect 3975 28886 3987 28920
rect 4021 28886 4037 28920
rect 3975 28852 4037 28886
rect 3975 28818 3987 28852
rect 4021 28818 4037 28852
rect 3975 28784 4037 28818
rect 3975 28750 3987 28784
rect 4021 28750 4037 28784
rect 3975 28733 4037 28750
rect 4067 28988 4133 29005
rect 4067 28954 4083 28988
rect 4117 28954 4133 28988
rect 4067 28920 4133 28954
rect 4067 28886 4083 28920
rect 4117 28886 4133 28920
rect 4067 28852 4133 28886
rect 4067 28818 4083 28852
rect 4117 28818 4133 28852
rect 4067 28784 4133 28818
rect 4067 28750 4083 28784
rect 4117 28750 4133 28784
rect 4067 28733 4133 28750
rect 4163 28988 4229 29005
rect 4163 28954 4179 28988
rect 4213 28954 4229 28988
rect 4163 28920 4229 28954
rect 4163 28886 4179 28920
rect 4213 28886 4229 28920
rect 4163 28852 4229 28886
rect 4163 28818 4179 28852
rect 4213 28818 4229 28852
rect 4163 28784 4229 28818
rect 4163 28750 4179 28784
rect 4213 28750 4229 28784
rect 4163 28733 4229 28750
rect 4259 28988 4325 29005
rect 4259 28954 4275 28988
rect 4309 28954 4325 28988
rect 4259 28920 4325 28954
rect 4259 28886 4275 28920
rect 4309 28886 4325 28920
rect 4259 28852 4325 28886
rect 4259 28818 4275 28852
rect 4309 28818 4325 28852
rect 4259 28784 4325 28818
rect 4259 28750 4275 28784
rect 4309 28750 4325 28784
rect 4259 28733 4325 28750
rect 4355 28988 4421 29005
rect 4355 28954 4371 28988
rect 4405 28954 4421 28988
rect 4355 28920 4421 28954
rect 4355 28886 4371 28920
rect 4405 28886 4421 28920
rect 4355 28852 4421 28886
rect 4355 28818 4371 28852
rect 4405 28818 4421 28852
rect 4355 28784 4421 28818
rect 4355 28750 4371 28784
rect 4405 28750 4421 28784
rect 4355 28733 4421 28750
rect 4451 28988 4517 29005
rect 4451 28954 4467 28988
rect 4501 28954 4517 28988
rect 4451 28920 4517 28954
rect 4451 28886 4467 28920
rect 4501 28886 4517 28920
rect 4451 28852 4517 28886
rect 4451 28818 4467 28852
rect 4501 28818 4517 28852
rect 4451 28784 4517 28818
rect 4451 28750 4467 28784
rect 4501 28750 4517 28784
rect 4451 28733 4517 28750
rect 4547 28988 4613 29005
rect 4547 28954 4563 28988
rect 4597 28954 4613 28988
rect 4547 28920 4613 28954
rect 4547 28886 4563 28920
rect 4597 28886 4613 28920
rect 4547 28852 4613 28886
rect 4547 28818 4563 28852
rect 4597 28818 4613 28852
rect 4547 28784 4613 28818
rect 4547 28750 4563 28784
rect 4597 28750 4613 28784
rect 4547 28733 4613 28750
rect 4643 28988 4709 29005
rect 4643 28954 4659 28988
rect 4693 28954 4709 28988
rect 4643 28920 4709 28954
rect 4643 28886 4659 28920
rect 4693 28886 4709 28920
rect 4643 28852 4709 28886
rect 4643 28818 4659 28852
rect 4693 28818 4709 28852
rect 4643 28784 4709 28818
rect 4643 28750 4659 28784
rect 4693 28750 4709 28784
rect 4643 28733 4709 28750
rect 4739 28988 4805 29005
rect 4739 28954 4755 28988
rect 4789 28954 4805 28988
rect 4739 28920 4805 28954
rect 4739 28886 4755 28920
rect 4789 28886 4805 28920
rect 4739 28852 4805 28886
rect 4739 28818 4755 28852
rect 4789 28818 4805 28852
rect 4739 28784 4805 28818
rect 4739 28750 4755 28784
rect 4789 28750 4805 28784
rect 4739 28733 4805 28750
rect 4835 28988 4901 29005
rect 4835 28954 4851 28988
rect 4885 28954 4901 28988
rect 4835 28920 4901 28954
rect 4835 28886 4851 28920
rect 4885 28886 4901 28920
rect 4835 28852 4901 28886
rect 4835 28818 4851 28852
rect 4885 28818 4901 28852
rect 4835 28784 4901 28818
rect 4835 28750 4851 28784
rect 4885 28750 4901 28784
rect 4835 28733 4901 28750
rect 4931 28988 4993 29005
rect 4931 28954 4947 28988
rect 4981 28954 4993 28988
rect 4931 28920 4993 28954
rect 4931 28886 4947 28920
rect 4981 28886 4993 28920
rect 4931 28852 4993 28886
rect 4931 28818 4947 28852
rect 4981 28818 4993 28852
rect 4931 28784 4993 28818
rect 4931 28750 4947 28784
rect 4981 28750 4993 28784
rect 4931 28733 4993 28750
rect 5348 28780 5400 28792
rect 5348 28746 5356 28780
rect 5390 28746 5400 28780
rect 5348 28712 5400 28746
rect 5348 28678 5356 28712
rect 5390 28678 5400 28712
rect 5348 28644 5400 28678
rect 5348 28610 5356 28644
rect 5390 28610 5400 28644
rect 5348 28592 5400 28610
rect 5430 28780 5482 28792
rect 5430 28746 5440 28780
rect 5474 28746 5482 28780
rect 5430 28712 5482 28746
rect 5430 28678 5440 28712
rect 5474 28678 5482 28712
rect 5430 28644 5482 28678
rect 5430 28610 5440 28644
rect 5474 28610 5482 28644
rect 5430 28592 5482 28610
rect 301 27697 363 27714
rect 301 27663 313 27697
rect 347 27663 363 27697
rect 301 27629 363 27663
rect 301 27595 313 27629
rect 347 27595 363 27629
rect 301 27561 363 27595
rect 301 27527 313 27561
rect 347 27527 363 27561
rect 301 27493 363 27527
rect 301 27459 313 27493
rect 347 27459 363 27493
rect 301 27442 363 27459
rect 393 27697 459 27714
rect 393 27663 409 27697
rect 443 27663 459 27697
rect 393 27629 459 27663
rect 393 27595 409 27629
rect 443 27595 459 27629
rect 393 27561 459 27595
rect 393 27527 409 27561
rect 443 27527 459 27561
rect 393 27493 459 27527
rect 393 27459 409 27493
rect 443 27459 459 27493
rect 393 27442 459 27459
rect 489 27697 555 27714
rect 489 27663 505 27697
rect 539 27663 555 27697
rect 489 27629 555 27663
rect 489 27595 505 27629
rect 539 27595 555 27629
rect 489 27561 555 27595
rect 489 27527 505 27561
rect 539 27527 555 27561
rect 489 27493 555 27527
rect 489 27459 505 27493
rect 539 27459 555 27493
rect 489 27442 555 27459
rect 585 27697 651 27714
rect 585 27663 601 27697
rect 635 27663 651 27697
rect 585 27629 651 27663
rect 585 27595 601 27629
rect 635 27595 651 27629
rect 585 27561 651 27595
rect 585 27527 601 27561
rect 635 27527 651 27561
rect 585 27493 651 27527
rect 585 27459 601 27493
rect 635 27459 651 27493
rect 585 27442 651 27459
rect 681 27697 747 27714
rect 681 27663 697 27697
rect 731 27663 747 27697
rect 681 27629 747 27663
rect 681 27595 697 27629
rect 731 27595 747 27629
rect 681 27561 747 27595
rect 681 27527 697 27561
rect 731 27527 747 27561
rect 681 27493 747 27527
rect 681 27459 697 27493
rect 731 27459 747 27493
rect 681 27442 747 27459
rect 777 27697 843 27714
rect 777 27663 793 27697
rect 827 27663 843 27697
rect 777 27629 843 27663
rect 777 27595 793 27629
rect 827 27595 843 27629
rect 777 27561 843 27595
rect 777 27527 793 27561
rect 827 27527 843 27561
rect 777 27493 843 27527
rect 777 27459 793 27493
rect 827 27459 843 27493
rect 777 27442 843 27459
rect 873 27697 939 27714
rect 873 27663 889 27697
rect 923 27663 939 27697
rect 873 27629 939 27663
rect 873 27595 889 27629
rect 923 27595 939 27629
rect 873 27561 939 27595
rect 873 27527 889 27561
rect 923 27527 939 27561
rect 873 27493 939 27527
rect 873 27459 889 27493
rect 923 27459 939 27493
rect 873 27442 939 27459
rect 969 27697 1035 27714
rect 969 27663 985 27697
rect 1019 27663 1035 27697
rect 969 27629 1035 27663
rect 969 27595 985 27629
rect 1019 27595 1035 27629
rect 969 27561 1035 27595
rect 969 27527 985 27561
rect 1019 27527 1035 27561
rect 969 27493 1035 27527
rect 969 27459 985 27493
rect 1019 27459 1035 27493
rect 969 27442 1035 27459
rect 1065 27697 1131 27714
rect 1065 27663 1081 27697
rect 1115 27663 1131 27697
rect 1065 27629 1131 27663
rect 1065 27595 1081 27629
rect 1115 27595 1131 27629
rect 1065 27561 1131 27595
rect 1065 27527 1081 27561
rect 1115 27527 1131 27561
rect 1065 27493 1131 27527
rect 1065 27459 1081 27493
rect 1115 27459 1131 27493
rect 1065 27442 1131 27459
rect 1161 27697 1227 27714
rect 1161 27663 1177 27697
rect 1211 27663 1227 27697
rect 1161 27629 1227 27663
rect 1161 27595 1177 27629
rect 1211 27595 1227 27629
rect 1161 27561 1227 27595
rect 1161 27527 1177 27561
rect 1211 27527 1227 27561
rect 1161 27493 1227 27527
rect 1161 27459 1177 27493
rect 1211 27459 1227 27493
rect 1161 27442 1227 27459
rect 1257 27697 1319 27714
rect 1257 27663 1273 27697
rect 1307 27663 1319 27697
rect 1257 27629 1319 27663
rect 1257 27595 1273 27629
rect 1307 27595 1319 27629
rect 1257 27561 1319 27595
rect 1257 27527 1273 27561
rect 1307 27527 1319 27561
rect 1257 27493 1319 27527
rect 1257 27459 1273 27493
rect 1307 27459 1319 27493
rect 1257 27442 1319 27459
rect 2454 27701 2516 27718
rect 2454 27667 2466 27701
rect 2500 27667 2516 27701
rect 2454 27633 2516 27667
rect 2454 27599 2466 27633
rect 2500 27599 2516 27633
rect 2454 27565 2516 27599
rect 2454 27531 2466 27565
rect 2500 27531 2516 27565
rect 2454 27497 2516 27531
rect 2454 27463 2466 27497
rect 2500 27463 2516 27497
rect 2454 27446 2516 27463
rect 2546 27701 2612 27718
rect 2546 27667 2562 27701
rect 2596 27667 2612 27701
rect 2546 27633 2612 27667
rect 2546 27599 2562 27633
rect 2596 27599 2612 27633
rect 2546 27565 2612 27599
rect 2546 27531 2562 27565
rect 2596 27531 2612 27565
rect 2546 27497 2612 27531
rect 2546 27463 2562 27497
rect 2596 27463 2612 27497
rect 2546 27446 2612 27463
rect 2642 27701 2708 27718
rect 2642 27667 2658 27701
rect 2692 27667 2708 27701
rect 2642 27633 2708 27667
rect 2642 27599 2658 27633
rect 2692 27599 2708 27633
rect 2642 27565 2708 27599
rect 2642 27531 2658 27565
rect 2692 27531 2708 27565
rect 2642 27497 2708 27531
rect 2642 27463 2658 27497
rect 2692 27463 2708 27497
rect 2642 27446 2708 27463
rect 2738 27701 2804 27718
rect 2738 27667 2754 27701
rect 2788 27667 2804 27701
rect 2738 27633 2804 27667
rect 2738 27599 2754 27633
rect 2788 27599 2804 27633
rect 2738 27565 2804 27599
rect 2738 27531 2754 27565
rect 2788 27531 2804 27565
rect 2738 27497 2804 27531
rect 2738 27463 2754 27497
rect 2788 27463 2804 27497
rect 2738 27446 2804 27463
rect 2834 27701 2900 27718
rect 2834 27667 2850 27701
rect 2884 27667 2900 27701
rect 2834 27633 2900 27667
rect 2834 27599 2850 27633
rect 2884 27599 2900 27633
rect 2834 27565 2900 27599
rect 2834 27531 2850 27565
rect 2884 27531 2900 27565
rect 2834 27497 2900 27531
rect 2834 27463 2850 27497
rect 2884 27463 2900 27497
rect 2834 27446 2900 27463
rect 2930 27701 2996 27718
rect 2930 27667 2946 27701
rect 2980 27667 2996 27701
rect 2930 27633 2996 27667
rect 2930 27599 2946 27633
rect 2980 27599 2996 27633
rect 2930 27565 2996 27599
rect 2930 27531 2946 27565
rect 2980 27531 2996 27565
rect 2930 27497 2996 27531
rect 2930 27463 2946 27497
rect 2980 27463 2996 27497
rect 2930 27446 2996 27463
rect 3026 27701 3092 27718
rect 3026 27667 3042 27701
rect 3076 27667 3092 27701
rect 3026 27633 3092 27667
rect 3026 27599 3042 27633
rect 3076 27599 3092 27633
rect 3026 27565 3092 27599
rect 3026 27531 3042 27565
rect 3076 27531 3092 27565
rect 3026 27497 3092 27531
rect 3026 27463 3042 27497
rect 3076 27463 3092 27497
rect 3026 27446 3092 27463
rect 3122 27701 3188 27718
rect 3122 27667 3138 27701
rect 3172 27667 3188 27701
rect 3122 27633 3188 27667
rect 3122 27599 3138 27633
rect 3172 27599 3188 27633
rect 3122 27565 3188 27599
rect 3122 27531 3138 27565
rect 3172 27531 3188 27565
rect 3122 27497 3188 27531
rect 3122 27463 3138 27497
rect 3172 27463 3188 27497
rect 3122 27446 3188 27463
rect 3218 27701 3284 27718
rect 3218 27667 3234 27701
rect 3268 27667 3284 27701
rect 3218 27633 3284 27667
rect 3218 27599 3234 27633
rect 3268 27599 3284 27633
rect 3218 27565 3284 27599
rect 3218 27531 3234 27565
rect 3268 27531 3284 27565
rect 3218 27497 3284 27531
rect 3218 27463 3234 27497
rect 3268 27463 3284 27497
rect 3218 27446 3284 27463
rect 3314 27701 3380 27718
rect 3314 27667 3330 27701
rect 3364 27667 3380 27701
rect 3314 27633 3380 27667
rect 3314 27599 3330 27633
rect 3364 27599 3380 27633
rect 3314 27565 3380 27599
rect 3314 27531 3330 27565
rect 3364 27531 3380 27565
rect 3314 27497 3380 27531
rect 3314 27463 3330 27497
rect 3364 27463 3380 27497
rect 3314 27446 3380 27463
rect 3410 27701 3472 27718
rect 3410 27667 3426 27701
rect 3460 27667 3472 27701
rect 3410 27633 3472 27667
rect 3410 27599 3426 27633
rect 3460 27599 3472 27633
rect 3410 27565 3472 27599
rect 3410 27531 3426 27565
rect 3460 27531 3472 27565
rect 3410 27497 3472 27531
rect 3410 27463 3426 27497
rect 3460 27463 3472 27497
rect 3410 27446 3472 27463
rect 3975 27701 4037 27718
rect 3975 27667 3987 27701
rect 4021 27667 4037 27701
rect 3975 27633 4037 27667
rect 3975 27599 3987 27633
rect 4021 27599 4037 27633
rect 3975 27565 4037 27599
rect 3975 27531 3987 27565
rect 4021 27531 4037 27565
rect 3975 27497 4037 27531
rect 3975 27463 3987 27497
rect 4021 27463 4037 27497
rect 3975 27446 4037 27463
rect 4067 27701 4133 27718
rect 4067 27667 4083 27701
rect 4117 27667 4133 27701
rect 4067 27633 4133 27667
rect 4067 27599 4083 27633
rect 4117 27599 4133 27633
rect 4067 27565 4133 27599
rect 4067 27531 4083 27565
rect 4117 27531 4133 27565
rect 4067 27497 4133 27531
rect 4067 27463 4083 27497
rect 4117 27463 4133 27497
rect 4067 27446 4133 27463
rect 4163 27701 4229 27718
rect 4163 27667 4179 27701
rect 4213 27667 4229 27701
rect 4163 27633 4229 27667
rect 4163 27599 4179 27633
rect 4213 27599 4229 27633
rect 4163 27565 4229 27599
rect 4163 27531 4179 27565
rect 4213 27531 4229 27565
rect 4163 27497 4229 27531
rect 4163 27463 4179 27497
rect 4213 27463 4229 27497
rect 4163 27446 4229 27463
rect 4259 27701 4325 27718
rect 4259 27667 4275 27701
rect 4309 27667 4325 27701
rect 4259 27633 4325 27667
rect 4259 27599 4275 27633
rect 4309 27599 4325 27633
rect 4259 27565 4325 27599
rect 4259 27531 4275 27565
rect 4309 27531 4325 27565
rect 4259 27497 4325 27531
rect 4259 27463 4275 27497
rect 4309 27463 4325 27497
rect 4259 27446 4325 27463
rect 4355 27701 4421 27718
rect 4355 27667 4371 27701
rect 4405 27667 4421 27701
rect 4355 27633 4421 27667
rect 4355 27599 4371 27633
rect 4405 27599 4421 27633
rect 4355 27565 4421 27599
rect 4355 27531 4371 27565
rect 4405 27531 4421 27565
rect 4355 27497 4421 27531
rect 4355 27463 4371 27497
rect 4405 27463 4421 27497
rect 4355 27446 4421 27463
rect 4451 27701 4517 27718
rect 4451 27667 4467 27701
rect 4501 27667 4517 27701
rect 4451 27633 4517 27667
rect 4451 27599 4467 27633
rect 4501 27599 4517 27633
rect 4451 27565 4517 27599
rect 4451 27531 4467 27565
rect 4501 27531 4517 27565
rect 4451 27497 4517 27531
rect 4451 27463 4467 27497
rect 4501 27463 4517 27497
rect 4451 27446 4517 27463
rect 4547 27701 4613 27718
rect 4547 27667 4563 27701
rect 4597 27667 4613 27701
rect 4547 27633 4613 27667
rect 4547 27599 4563 27633
rect 4597 27599 4613 27633
rect 4547 27565 4613 27599
rect 4547 27531 4563 27565
rect 4597 27531 4613 27565
rect 4547 27497 4613 27531
rect 4547 27463 4563 27497
rect 4597 27463 4613 27497
rect 4547 27446 4613 27463
rect 4643 27701 4709 27718
rect 4643 27667 4659 27701
rect 4693 27667 4709 27701
rect 4643 27633 4709 27667
rect 4643 27599 4659 27633
rect 4693 27599 4709 27633
rect 4643 27565 4709 27599
rect 4643 27531 4659 27565
rect 4693 27531 4709 27565
rect 4643 27497 4709 27531
rect 4643 27463 4659 27497
rect 4693 27463 4709 27497
rect 4643 27446 4709 27463
rect 4739 27701 4805 27718
rect 4739 27667 4755 27701
rect 4789 27667 4805 27701
rect 4739 27633 4805 27667
rect 4739 27599 4755 27633
rect 4789 27599 4805 27633
rect 4739 27565 4805 27599
rect 4739 27531 4755 27565
rect 4789 27531 4805 27565
rect 4739 27497 4805 27531
rect 4739 27463 4755 27497
rect 4789 27463 4805 27497
rect 4739 27446 4805 27463
rect 4835 27701 4901 27718
rect 4835 27667 4851 27701
rect 4885 27667 4901 27701
rect 4835 27633 4901 27667
rect 4835 27599 4851 27633
rect 4885 27599 4901 27633
rect 4835 27565 4901 27599
rect 4835 27531 4851 27565
rect 4885 27531 4901 27565
rect 4835 27497 4901 27531
rect 4835 27463 4851 27497
rect 4885 27463 4901 27497
rect 4835 27446 4901 27463
rect 4931 27701 4993 27718
rect 4931 27667 4947 27701
rect 4981 27667 4993 27701
rect 4931 27633 4993 27667
rect 4931 27599 4947 27633
rect 4981 27599 4993 27633
rect 4931 27565 4993 27599
rect 4931 27531 4947 27565
rect 4981 27531 4993 27565
rect 4931 27497 4993 27531
rect 4931 27463 4947 27497
rect 4981 27463 4993 27497
rect 4931 27446 4993 27463
rect 5348 27493 5400 27505
rect 5348 27459 5356 27493
rect 5390 27459 5400 27493
rect 5348 27425 5400 27459
rect 5348 27391 5356 27425
rect 5390 27391 5400 27425
rect 5348 27357 5400 27391
rect 5348 27323 5356 27357
rect 5390 27323 5400 27357
rect 5348 27305 5400 27323
rect 5430 27493 5482 27505
rect 5430 27459 5440 27493
rect 5474 27459 5482 27493
rect 5430 27425 5482 27459
rect 5430 27391 5440 27425
rect 5474 27391 5482 27425
rect 5430 27357 5482 27391
rect 5430 27323 5440 27357
rect 5474 27323 5482 27357
rect 5430 27305 5482 27323
rect 301 26410 363 26427
rect 301 26376 313 26410
rect 347 26376 363 26410
rect 301 26342 363 26376
rect 301 26308 313 26342
rect 347 26308 363 26342
rect 301 26274 363 26308
rect 301 26240 313 26274
rect 347 26240 363 26274
rect 301 26206 363 26240
rect 301 26172 313 26206
rect 347 26172 363 26206
rect 301 26155 363 26172
rect 393 26410 459 26427
rect 393 26376 409 26410
rect 443 26376 459 26410
rect 393 26342 459 26376
rect 393 26308 409 26342
rect 443 26308 459 26342
rect 393 26274 459 26308
rect 393 26240 409 26274
rect 443 26240 459 26274
rect 393 26206 459 26240
rect 393 26172 409 26206
rect 443 26172 459 26206
rect 393 26155 459 26172
rect 489 26410 555 26427
rect 489 26376 505 26410
rect 539 26376 555 26410
rect 489 26342 555 26376
rect 489 26308 505 26342
rect 539 26308 555 26342
rect 489 26274 555 26308
rect 489 26240 505 26274
rect 539 26240 555 26274
rect 489 26206 555 26240
rect 489 26172 505 26206
rect 539 26172 555 26206
rect 489 26155 555 26172
rect 585 26410 651 26427
rect 585 26376 601 26410
rect 635 26376 651 26410
rect 585 26342 651 26376
rect 585 26308 601 26342
rect 635 26308 651 26342
rect 585 26274 651 26308
rect 585 26240 601 26274
rect 635 26240 651 26274
rect 585 26206 651 26240
rect 585 26172 601 26206
rect 635 26172 651 26206
rect 585 26155 651 26172
rect 681 26410 747 26427
rect 681 26376 697 26410
rect 731 26376 747 26410
rect 681 26342 747 26376
rect 681 26308 697 26342
rect 731 26308 747 26342
rect 681 26274 747 26308
rect 681 26240 697 26274
rect 731 26240 747 26274
rect 681 26206 747 26240
rect 681 26172 697 26206
rect 731 26172 747 26206
rect 681 26155 747 26172
rect 777 26410 843 26427
rect 777 26376 793 26410
rect 827 26376 843 26410
rect 777 26342 843 26376
rect 777 26308 793 26342
rect 827 26308 843 26342
rect 777 26274 843 26308
rect 777 26240 793 26274
rect 827 26240 843 26274
rect 777 26206 843 26240
rect 777 26172 793 26206
rect 827 26172 843 26206
rect 777 26155 843 26172
rect 873 26410 939 26427
rect 873 26376 889 26410
rect 923 26376 939 26410
rect 873 26342 939 26376
rect 873 26308 889 26342
rect 923 26308 939 26342
rect 873 26274 939 26308
rect 873 26240 889 26274
rect 923 26240 939 26274
rect 873 26206 939 26240
rect 873 26172 889 26206
rect 923 26172 939 26206
rect 873 26155 939 26172
rect 969 26410 1035 26427
rect 969 26376 985 26410
rect 1019 26376 1035 26410
rect 969 26342 1035 26376
rect 969 26308 985 26342
rect 1019 26308 1035 26342
rect 969 26274 1035 26308
rect 969 26240 985 26274
rect 1019 26240 1035 26274
rect 969 26206 1035 26240
rect 969 26172 985 26206
rect 1019 26172 1035 26206
rect 969 26155 1035 26172
rect 1065 26410 1131 26427
rect 1065 26376 1081 26410
rect 1115 26376 1131 26410
rect 1065 26342 1131 26376
rect 1065 26308 1081 26342
rect 1115 26308 1131 26342
rect 1065 26274 1131 26308
rect 1065 26240 1081 26274
rect 1115 26240 1131 26274
rect 1065 26206 1131 26240
rect 1065 26172 1081 26206
rect 1115 26172 1131 26206
rect 1065 26155 1131 26172
rect 1161 26410 1227 26427
rect 1161 26376 1177 26410
rect 1211 26376 1227 26410
rect 1161 26342 1227 26376
rect 1161 26308 1177 26342
rect 1211 26308 1227 26342
rect 1161 26274 1227 26308
rect 1161 26240 1177 26274
rect 1211 26240 1227 26274
rect 1161 26206 1227 26240
rect 1161 26172 1177 26206
rect 1211 26172 1227 26206
rect 1161 26155 1227 26172
rect 1257 26410 1319 26427
rect 1257 26376 1273 26410
rect 1307 26376 1319 26410
rect 1257 26342 1319 26376
rect 1257 26308 1273 26342
rect 1307 26308 1319 26342
rect 1257 26274 1319 26308
rect 1257 26240 1273 26274
rect 1307 26240 1319 26274
rect 1257 26206 1319 26240
rect 1257 26172 1273 26206
rect 1307 26172 1319 26206
rect 1257 26155 1319 26172
rect 2454 26414 2516 26431
rect 2454 26380 2466 26414
rect 2500 26380 2516 26414
rect 2454 26346 2516 26380
rect 2454 26312 2466 26346
rect 2500 26312 2516 26346
rect 2454 26278 2516 26312
rect 2454 26244 2466 26278
rect 2500 26244 2516 26278
rect 2454 26210 2516 26244
rect 2454 26176 2466 26210
rect 2500 26176 2516 26210
rect 2454 26159 2516 26176
rect 2546 26414 2612 26431
rect 2546 26380 2562 26414
rect 2596 26380 2612 26414
rect 2546 26346 2612 26380
rect 2546 26312 2562 26346
rect 2596 26312 2612 26346
rect 2546 26278 2612 26312
rect 2546 26244 2562 26278
rect 2596 26244 2612 26278
rect 2546 26210 2612 26244
rect 2546 26176 2562 26210
rect 2596 26176 2612 26210
rect 2546 26159 2612 26176
rect 2642 26414 2708 26431
rect 2642 26380 2658 26414
rect 2692 26380 2708 26414
rect 2642 26346 2708 26380
rect 2642 26312 2658 26346
rect 2692 26312 2708 26346
rect 2642 26278 2708 26312
rect 2642 26244 2658 26278
rect 2692 26244 2708 26278
rect 2642 26210 2708 26244
rect 2642 26176 2658 26210
rect 2692 26176 2708 26210
rect 2642 26159 2708 26176
rect 2738 26414 2804 26431
rect 2738 26380 2754 26414
rect 2788 26380 2804 26414
rect 2738 26346 2804 26380
rect 2738 26312 2754 26346
rect 2788 26312 2804 26346
rect 2738 26278 2804 26312
rect 2738 26244 2754 26278
rect 2788 26244 2804 26278
rect 2738 26210 2804 26244
rect 2738 26176 2754 26210
rect 2788 26176 2804 26210
rect 2738 26159 2804 26176
rect 2834 26414 2900 26431
rect 2834 26380 2850 26414
rect 2884 26380 2900 26414
rect 2834 26346 2900 26380
rect 2834 26312 2850 26346
rect 2884 26312 2900 26346
rect 2834 26278 2900 26312
rect 2834 26244 2850 26278
rect 2884 26244 2900 26278
rect 2834 26210 2900 26244
rect 2834 26176 2850 26210
rect 2884 26176 2900 26210
rect 2834 26159 2900 26176
rect 2930 26414 2996 26431
rect 2930 26380 2946 26414
rect 2980 26380 2996 26414
rect 2930 26346 2996 26380
rect 2930 26312 2946 26346
rect 2980 26312 2996 26346
rect 2930 26278 2996 26312
rect 2930 26244 2946 26278
rect 2980 26244 2996 26278
rect 2930 26210 2996 26244
rect 2930 26176 2946 26210
rect 2980 26176 2996 26210
rect 2930 26159 2996 26176
rect 3026 26414 3092 26431
rect 3026 26380 3042 26414
rect 3076 26380 3092 26414
rect 3026 26346 3092 26380
rect 3026 26312 3042 26346
rect 3076 26312 3092 26346
rect 3026 26278 3092 26312
rect 3026 26244 3042 26278
rect 3076 26244 3092 26278
rect 3026 26210 3092 26244
rect 3026 26176 3042 26210
rect 3076 26176 3092 26210
rect 3026 26159 3092 26176
rect 3122 26414 3188 26431
rect 3122 26380 3138 26414
rect 3172 26380 3188 26414
rect 3122 26346 3188 26380
rect 3122 26312 3138 26346
rect 3172 26312 3188 26346
rect 3122 26278 3188 26312
rect 3122 26244 3138 26278
rect 3172 26244 3188 26278
rect 3122 26210 3188 26244
rect 3122 26176 3138 26210
rect 3172 26176 3188 26210
rect 3122 26159 3188 26176
rect 3218 26414 3284 26431
rect 3218 26380 3234 26414
rect 3268 26380 3284 26414
rect 3218 26346 3284 26380
rect 3218 26312 3234 26346
rect 3268 26312 3284 26346
rect 3218 26278 3284 26312
rect 3218 26244 3234 26278
rect 3268 26244 3284 26278
rect 3218 26210 3284 26244
rect 3218 26176 3234 26210
rect 3268 26176 3284 26210
rect 3218 26159 3284 26176
rect 3314 26414 3380 26431
rect 3314 26380 3330 26414
rect 3364 26380 3380 26414
rect 3314 26346 3380 26380
rect 3314 26312 3330 26346
rect 3364 26312 3380 26346
rect 3314 26278 3380 26312
rect 3314 26244 3330 26278
rect 3364 26244 3380 26278
rect 3314 26210 3380 26244
rect 3314 26176 3330 26210
rect 3364 26176 3380 26210
rect 3314 26159 3380 26176
rect 3410 26414 3472 26431
rect 3410 26380 3426 26414
rect 3460 26380 3472 26414
rect 3410 26346 3472 26380
rect 3410 26312 3426 26346
rect 3460 26312 3472 26346
rect 3410 26278 3472 26312
rect 3410 26244 3426 26278
rect 3460 26244 3472 26278
rect 3410 26210 3472 26244
rect 3410 26176 3426 26210
rect 3460 26176 3472 26210
rect 3410 26159 3472 26176
rect 3975 26414 4037 26431
rect 3975 26380 3987 26414
rect 4021 26380 4037 26414
rect 3975 26346 4037 26380
rect 3975 26312 3987 26346
rect 4021 26312 4037 26346
rect 3975 26278 4037 26312
rect 3975 26244 3987 26278
rect 4021 26244 4037 26278
rect 3975 26210 4037 26244
rect 3975 26176 3987 26210
rect 4021 26176 4037 26210
rect 3975 26159 4037 26176
rect 4067 26414 4133 26431
rect 4067 26380 4083 26414
rect 4117 26380 4133 26414
rect 4067 26346 4133 26380
rect 4067 26312 4083 26346
rect 4117 26312 4133 26346
rect 4067 26278 4133 26312
rect 4067 26244 4083 26278
rect 4117 26244 4133 26278
rect 4067 26210 4133 26244
rect 4067 26176 4083 26210
rect 4117 26176 4133 26210
rect 4067 26159 4133 26176
rect 4163 26414 4229 26431
rect 4163 26380 4179 26414
rect 4213 26380 4229 26414
rect 4163 26346 4229 26380
rect 4163 26312 4179 26346
rect 4213 26312 4229 26346
rect 4163 26278 4229 26312
rect 4163 26244 4179 26278
rect 4213 26244 4229 26278
rect 4163 26210 4229 26244
rect 4163 26176 4179 26210
rect 4213 26176 4229 26210
rect 4163 26159 4229 26176
rect 4259 26414 4325 26431
rect 4259 26380 4275 26414
rect 4309 26380 4325 26414
rect 4259 26346 4325 26380
rect 4259 26312 4275 26346
rect 4309 26312 4325 26346
rect 4259 26278 4325 26312
rect 4259 26244 4275 26278
rect 4309 26244 4325 26278
rect 4259 26210 4325 26244
rect 4259 26176 4275 26210
rect 4309 26176 4325 26210
rect 4259 26159 4325 26176
rect 4355 26414 4421 26431
rect 4355 26380 4371 26414
rect 4405 26380 4421 26414
rect 4355 26346 4421 26380
rect 4355 26312 4371 26346
rect 4405 26312 4421 26346
rect 4355 26278 4421 26312
rect 4355 26244 4371 26278
rect 4405 26244 4421 26278
rect 4355 26210 4421 26244
rect 4355 26176 4371 26210
rect 4405 26176 4421 26210
rect 4355 26159 4421 26176
rect 4451 26414 4517 26431
rect 4451 26380 4467 26414
rect 4501 26380 4517 26414
rect 4451 26346 4517 26380
rect 4451 26312 4467 26346
rect 4501 26312 4517 26346
rect 4451 26278 4517 26312
rect 4451 26244 4467 26278
rect 4501 26244 4517 26278
rect 4451 26210 4517 26244
rect 4451 26176 4467 26210
rect 4501 26176 4517 26210
rect 4451 26159 4517 26176
rect 4547 26414 4613 26431
rect 4547 26380 4563 26414
rect 4597 26380 4613 26414
rect 4547 26346 4613 26380
rect 4547 26312 4563 26346
rect 4597 26312 4613 26346
rect 4547 26278 4613 26312
rect 4547 26244 4563 26278
rect 4597 26244 4613 26278
rect 4547 26210 4613 26244
rect 4547 26176 4563 26210
rect 4597 26176 4613 26210
rect 4547 26159 4613 26176
rect 4643 26414 4709 26431
rect 4643 26380 4659 26414
rect 4693 26380 4709 26414
rect 4643 26346 4709 26380
rect 4643 26312 4659 26346
rect 4693 26312 4709 26346
rect 4643 26278 4709 26312
rect 4643 26244 4659 26278
rect 4693 26244 4709 26278
rect 4643 26210 4709 26244
rect 4643 26176 4659 26210
rect 4693 26176 4709 26210
rect 4643 26159 4709 26176
rect 4739 26414 4805 26431
rect 4739 26380 4755 26414
rect 4789 26380 4805 26414
rect 4739 26346 4805 26380
rect 4739 26312 4755 26346
rect 4789 26312 4805 26346
rect 4739 26278 4805 26312
rect 4739 26244 4755 26278
rect 4789 26244 4805 26278
rect 4739 26210 4805 26244
rect 4739 26176 4755 26210
rect 4789 26176 4805 26210
rect 4739 26159 4805 26176
rect 4835 26414 4901 26431
rect 4835 26380 4851 26414
rect 4885 26380 4901 26414
rect 4835 26346 4901 26380
rect 4835 26312 4851 26346
rect 4885 26312 4901 26346
rect 4835 26278 4901 26312
rect 4835 26244 4851 26278
rect 4885 26244 4901 26278
rect 4835 26210 4901 26244
rect 4835 26176 4851 26210
rect 4885 26176 4901 26210
rect 4835 26159 4901 26176
rect 4931 26414 4993 26431
rect 4931 26380 4947 26414
rect 4981 26380 4993 26414
rect 4931 26346 4993 26380
rect 4931 26312 4947 26346
rect 4981 26312 4993 26346
rect 4931 26278 4993 26312
rect 4931 26244 4947 26278
rect 4981 26244 4993 26278
rect 4931 26210 4993 26244
rect 4931 26176 4947 26210
rect 4981 26176 4993 26210
rect 4931 26159 4993 26176
rect 5348 26206 5400 26218
rect 5348 26172 5356 26206
rect 5390 26172 5400 26206
rect 5348 26138 5400 26172
rect 5348 26104 5356 26138
rect 5390 26104 5400 26138
rect 5348 26070 5400 26104
rect 5348 26036 5356 26070
rect 5390 26036 5400 26070
rect 5348 26018 5400 26036
rect 5430 26206 5482 26218
rect 5430 26172 5440 26206
rect 5474 26172 5482 26206
rect 5430 26138 5482 26172
rect 5430 26104 5440 26138
rect 5474 26104 5482 26138
rect 5430 26070 5482 26104
rect 5430 26036 5440 26070
rect 5474 26036 5482 26070
rect 5430 26018 5482 26036
rect 301 25123 363 25140
rect 301 25089 313 25123
rect 347 25089 363 25123
rect 301 25055 363 25089
rect 301 25021 313 25055
rect 347 25021 363 25055
rect 301 24987 363 25021
rect 301 24953 313 24987
rect 347 24953 363 24987
rect 301 24919 363 24953
rect 301 24885 313 24919
rect 347 24885 363 24919
rect 301 24868 363 24885
rect 393 25123 459 25140
rect 393 25089 409 25123
rect 443 25089 459 25123
rect 393 25055 459 25089
rect 393 25021 409 25055
rect 443 25021 459 25055
rect 393 24987 459 25021
rect 393 24953 409 24987
rect 443 24953 459 24987
rect 393 24919 459 24953
rect 393 24885 409 24919
rect 443 24885 459 24919
rect 393 24868 459 24885
rect 489 25123 555 25140
rect 489 25089 505 25123
rect 539 25089 555 25123
rect 489 25055 555 25089
rect 489 25021 505 25055
rect 539 25021 555 25055
rect 489 24987 555 25021
rect 489 24953 505 24987
rect 539 24953 555 24987
rect 489 24919 555 24953
rect 489 24885 505 24919
rect 539 24885 555 24919
rect 489 24868 555 24885
rect 585 25123 651 25140
rect 585 25089 601 25123
rect 635 25089 651 25123
rect 585 25055 651 25089
rect 585 25021 601 25055
rect 635 25021 651 25055
rect 585 24987 651 25021
rect 585 24953 601 24987
rect 635 24953 651 24987
rect 585 24919 651 24953
rect 585 24885 601 24919
rect 635 24885 651 24919
rect 585 24868 651 24885
rect 681 25123 747 25140
rect 681 25089 697 25123
rect 731 25089 747 25123
rect 681 25055 747 25089
rect 681 25021 697 25055
rect 731 25021 747 25055
rect 681 24987 747 25021
rect 681 24953 697 24987
rect 731 24953 747 24987
rect 681 24919 747 24953
rect 681 24885 697 24919
rect 731 24885 747 24919
rect 681 24868 747 24885
rect 777 25123 843 25140
rect 777 25089 793 25123
rect 827 25089 843 25123
rect 777 25055 843 25089
rect 777 25021 793 25055
rect 827 25021 843 25055
rect 777 24987 843 25021
rect 777 24953 793 24987
rect 827 24953 843 24987
rect 777 24919 843 24953
rect 777 24885 793 24919
rect 827 24885 843 24919
rect 777 24868 843 24885
rect 873 25123 939 25140
rect 873 25089 889 25123
rect 923 25089 939 25123
rect 873 25055 939 25089
rect 873 25021 889 25055
rect 923 25021 939 25055
rect 873 24987 939 25021
rect 873 24953 889 24987
rect 923 24953 939 24987
rect 873 24919 939 24953
rect 873 24885 889 24919
rect 923 24885 939 24919
rect 873 24868 939 24885
rect 969 25123 1035 25140
rect 969 25089 985 25123
rect 1019 25089 1035 25123
rect 969 25055 1035 25089
rect 969 25021 985 25055
rect 1019 25021 1035 25055
rect 969 24987 1035 25021
rect 969 24953 985 24987
rect 1019 24953 1035 24987
rect 969 24919 1035 24953
rect 969 24885 985 24919
rect 1019 24885 1035 24919
rect 969 24868 1035 24885
rect 1065 25123 1131 25140
rect 1065 25089 1081 25123
rect 1115 25089 1131 25123
rect 1065 25055 1131 25089
rect 1065 25021 1081 25055
rect 1115 25021 1131 25055
rect 1065 24987 1131 25021
rect 1065 24953 1081 24987
rect 1115 24953 1131 24987
rect 1065 24919 1131 24953
rect 1065 24885 1081 24919
rect 1115 24885 1131 24919
rect 1065 24868 1131 24885
rect 1161 25123 1227 25140
rect 1161 25089 1177 25123
rect 1211 25089 1227 25123
rect 1161 25055 1227 25089
rect 1161 25021 1177 25055
rect 1211 25021 1227 25055
rect 1161 24987 1227 25021
rect 1161 24953 1177 24987
rect 1211 24953 1227 24987
rect 1161 24919 1227 24953
rect 1161 24885 1177 24919
rect 1211 24885 1227 24919
rect 1161 24868 1227 24885
rect 1257 25123 1319 25140
rect 1257 25089 1273 25123
rect 1307 25089 1319 25123
rect 1257 25055 1319 25089
rect 1257 25021 1273 25055
rect 1307 25021 1319 25055
rect 1257 24987 1319 25021
rect 1257 24953 1273 24987
rect 1307 24953 1319 24987
rect 1257 24919 1319 24953
rect 1257 24885 1273 24919
rect 1307 24885 1319 24919
rect 1257 24868 1319 24885
rect 2454 25127 2516 25144
rect 2454 25093 2466 25127
rect 2500 25093 2516 25127
rect 2454 25059 2516 25093
rect 2454 25025 2466 25059
rect 2500 25025 2516 25059
rect 2454 24991 2516 25025
rect 2454 24957 2466 24991
rect 2500 24957 2516 24991
rect 2454 24923 2516 24957
rect 2454 24889 2466 24923
rect 2500 24889 2516 24923
rect 2454 24872 2516 24889
rect 2546 25127 2612 25144
rect 2546 25093 2562 25127
rect 2596 25093 2612 25127
rect 2546 25059 2612 25093
rect 2546 25025 2562 25059
rect 2596 25025 2612 25059
rect 2546 24991 2612 25025
rect 2546 24957 2562 24991
rect 2596 24957 2612 24991
rect 2546 24923 2612 24957
rect 2546 24889 2562 24923
rect 2596 24889 2612 24923
rect 2546 24872 2612 24889
rect 2642 25127 2708 25144
rect 2642 25093 2658 25127
rect 2692 25093 2708 25127
rect 2642 25059 2708 25093
rect 2642 25025 2658 25059
rect 2692 25025 2708 25059
rect 2642 24991 2708 25025
rect 2642 24957 2658 24991
rect 2692 24957 2708 24991
rect 2642 24923 2708 24957
rect 2642 24889 2658 24923
rect 2692 24889 2708 24923
rect 2642 24872 2708 24889
rect 2738 25127 2804 25144
rect 2738 25093 2754 25127
rect 2788 25093 2804 25127
rect 2738 25059 2804 25093
rect 2738 25025 2754 25059
rect 2788 25025 2804 25059
rect 2738 24991 2804 25025
rect 2738 24957 2754 24991
rect 2788 24957 2804 24991
rect 2738 24923 2804 24957
rect 2738 24889 2754 24923
rect 2788 24889 2804 24923
rect 2738 24872 2804 24889
rect 2834 25127 2900 25144
rect 2834 25093 2850 25127
rect 2884 25093 2900 25127
rect 2834 25059 2900 25093
rect 2834 25025 2850 25059
rect 2884 25025 2900 25059
rect 2834 24991 2900 25025
rect 2834 24957 2850 24991
rect 2884 24957 2900 24991
rect 2834 24923 2900 24957
rect 2834 24889 2850 24923
rect 2884 24889 2900 24923
rect 2834 24872 2900 24889
rect 2930 25127 2996 25144
rect 2930 25093 2946 25127
rect 2980 25093 2996 25127
rect 2930 25059 2996 25093
rect 2930 25025 2946 25059
rect 2980 25025 2996 25059
rect 2930 24991 2996 25025
rect 2930 24957 2946 24991
rect 2980 24957 2996 24991
rect 2930 24923 2996 24957
rect 2930 24889 2946 24923
rect 2980 24889 2996 24923
rect 2930 24872 2996 24889
rect 3026 25127 3092 25144
rect 3026 25093 3042 25127
rect 3076 25093 3092 25127
rect 3026 25059 3092 25093
rect 3026 25025 3042 25059
rect 3076 25025 3092 25059
rect 3026 24991 3092 25025
rect 3026 24957 3042 24991
rect 3076 24957 3092 24991
rect 3026 24923 3092 24957
rect 3026 24889 3042 24923
rect 3076 24889 3092 24923
rect 3026 24872 3092 24889
rect 3122 25127 3188 25144
rect 3122 25093 3138 25127
rect 3172 25093 3188 25127
rect 3122 25059 3188 25093
rect 3122 25025 3138 25059
rect 3172 25025 3188 25059
rect 3122 24991 3188 25025
rect 3122 24957 3138 24991
rect 3172 24957 3188 24991
rect 3122 24923 3188 24957
rect 3122 24889 3138 24923
rect 3172 24889 3188 24923
rect 3122 24872 3188 24889
rect 3218 25127 3284 25144
rect 3218 25093 3234 25127
rect 3268 25093 3284 25127
rect 3218 25059 3284 25093
rect 3218 25025 3234 25059
rect 3268 25025 3284 25059
rect 3218 24991 3284 25025
rect 3218 24957 3234 24991
rect 3268 24957 3284 24991
rect 3218 24923 3284 24957
rect 3218 24889 3234 24923
rect 3268 24889 3284 24923
rect 3218 24872 3284 24889
rect 3314 25127 3380 25144
rect 3314 25093 3330 25127
rect 3364 25093 3380 25127
rect 3314 25059 3380 25093
rect 3314 25025 3330 25059
rect 3364 25025 3380 25059
rect 3314 24991 3380 25025
rect 3314 24957 3330 24991
rect 3364 24957 3380 24991
rect 3314 24923 3380 24957
rect 3314 24889 3330 24923
rect 3364 24889 3380 24923
rect 3314 24872 3380 24889
rect 3410 25127 3472 25144
rect 3410 25093 3426 25127
rect 3460 25093 3472 25127
rect 3410 25059 3472 25093
rect 3410 25025 3426 25059
rect 3460 25025 3472 25059
rect 3410 24991 3472 25025
rect 3410 24957 3426 24991
rect 3460 24957 3472 24991
rect 3410 24923 3472 24957
rect 3410 24889 3426 24923
rect 3460 24889 3472 24923
rect 3410 24872 3472 24889
rect 3975 25127 4037 25144
rect 3975 25093 3987 25127
rect 4021 25093 4037 25127
rect 3975 25059 4037 25093
rect 3975 25025 3987 25059
rect 4021 25025 4037 25059
rect 3975 24991 4037 25025
rect 3975 24957 3987 24991
rect 4021 24957 4037 24991
rect 3975 24923 4037 24957
rect 3975 24889 3987 24923
rect 4021 24889 4037 24923
rect 3975 24872 4037 24889
rect 4067 25127 4133 25144
rect 4067 25093 4083 25127
rect 4117 25093 4133 25127
rect 4067 25059 4133 25093
rect 4067 25025 4083 25059
rect 4117 25025 4133 25059
rect 4067 24991 4133 25025
rect 4067 24957 4083 24991
rect 4117 24957 4133 24991
rect 4067 24923 4133 24957
rect 4067 24889 4083 24923
rect 4117 24889 4133 24923
rect 4067 24872 4133 24889
rect 4163 25127 4229 25144
rect 4163 25093 4179 25127
rect 4213 25093 4229 25127
rect 4163 25059 4229 25093
rect 4163 25025 4179 25059
rect 4213 25025 4229 25059
rect 4163 24991 4229 25025
rect 4163 24957 4179 24991
rect 4213 24957 4229 24991
rect 4163 24923 4229 24957
rect 4163 24889 4179 24923
rect 4213 24889 4229 24923
rect 4163 24872 4229 24889
rect 4259 25127 4325 25144
rect 4259 25093 4275 25127
rect 4309 25093 4325 25127
rect 4259 25059 4325 25093
rect 4259 25025 4275 25059
rect 4309 25025 4325 25059
rect 4259 24991 4325 25025
rect 4259 24957 4275 24991
rect 4309 24957 4325 24991
rect 4259 24923 4325 24957
rect 4259 24889 4275 24923
rect 4309 24889 4325 24923
rect 4259 24872 4325 24889
rect 4355 25127 4421 25144
rect 4355 25093 4371 25127
rect 4405 25093 4421 25127
rect 4355 25059 4421 25093
rect 4355 25025 4371 25059
rect 4405 25025 4421 25059
rect 4355 24991 4421 25025
rect 4355 24957 4371 24991
rect 4405 24957 4421 24991
rect 4355 24923 4421 24957
rect 4355 24889 4371 24923
rect 4405 24889 4421 24923
rect 4355 24872 4421 24889
rect 4451 25127 4517 25144
rect 4451 25093 4467 25127
rect 4501 25093 4517 25127
rect 4451 25059 4517 25093
rect 4451 25025 4467 25059
rect 4501 25025 4517 25059
rect 4451 24991 4517 25025
rect 4451 24957 4467 24991
rect 4501 24957 4517 24991
rect 4451 24923 4517 24957
rect 4451 24889 4467 24923
rect 4501 24889 4517 24923
rect 4451 24872 4517 24889
rect 4547 25127 4613 25144
rect 4547 25093 4563 25127
rect 4597 25093 4613 25127
rect 4547 25059 4613 25093
rect 4547 25025 4563 25059
rect 4597 25025 4613 25059
rect 4547 24991 4613 25025
rect 4547 24957 4563 24991
rect 4597 24957 4613 24991
rect 4547 24923 4613 24957
rect 4547 24889 4563 24923
rect 4597 24889 4613 24923
rect 4547 24872 4613 24889
rect 4643 25127 4709 25144
rect 4643 25093 4659 25127
rect 4693 25093 4709 25127
rect 4643 25059 4709 25093
rect 4643 25025 4659 25059
rect 4693 25025 4709 25059
rect 4643 24991 4709 25025
rect 4643 24957 4659 24991
rect 4693 24957 4709 24991
rect 4643 24923 4709 24957
rect 4643 24889 4659 24923
rect 4693 24889 4709 24923
rect 4643 24872 4709 24889
rect 4739 25127 4805 25144
rect 4739 25093 4755 25127
rect 4789 25093 4805 25127
rect 4739 25059 4805 25093
rect 4739 25025 4755 25059
rect 4789 25025 4805 25059
rect 4739 24991 4805 25025
rect 4739 24957 4755 24991
rect 4789 24957 4805 24991
rect 4739 24923 4805 24957
rect 4739 24889 4755 24923
rect 4789 24889 4805 24923
rect 4739 24872 4805 24889
rect 4835 25127 4901 25144
rect 4835 25093 4851 25127
rect 4885 25093 4901 25127
rect 4835 25059 4901 25093
rect 4835 25025 4851 25059
rect 4885 25025 4901 25059
rect 4835 24991 4901 25025
rect 4835 24957 4851 24991
rect 4885 24957 4901 24991
rect 4835 24923 4901 24957
rect 4835 24889 4851 24923
rect 4885 24889 4901 24923
rect 4835 24872 4901 24889
rect 4931 25127 4993 25144
rect 4931 25093 4947 25127
rect 4981 25093 4993 25127
rect 4931 25059 4993 25093
rect 4931 25025 4947 25059
rect 4981 25025 4993 25059
rect 4931 24991 4993 25025
rect 4931 24957 4947 24991
rect 4981 24957 4993 24991
rect 4931 24923 4993 24957
rect 4931 24889 4947 24923
rect 4981 24889 4993 24923
rect 4931 24872 4993 24889
rect 5348 24919 5400 24931
rect 5348 24885 5356 24919
rect 5390 24885 5400 24919
rect 5348 24851 5400 24885
rect 5348 24817 5356 24851
rect 5390 24817 5400 24851
rect 5348 24783 5400 24817
rect 5348 24749 5356 24783
rect 5390 24749 5400 24783
rect 5348 24731 5400 24749
rect 5430 24919 5482 24931
rect 5430 24885 5440 24919
rect 5474 24885 5482 24919
rect 5430 24851 5482 24885
rect 5430 24817 5440 24851
rect 5474 24817 5482 24851
rect 5430 24783 5482 24817
rect 5430 24749 5440 24783
rect 5474 24749 5482 24783
rect 5430 24731 5482 24749
rect 301 23836 363 23853
rect 301 23802 313 23836
rect 347 23802 363 23836
rect 301 23768 363 23802
rect 301 23734 313 23768
rect 347 23734 363 23768
rect 301 23700 363 23734
rect 301 23666 313 23700
rect 347 23666 363 23700
rect 301 23632 363 23666
rect 301 23598 313 23632
rect 347 23598 363 23632
rect 301 23581 363 23598
rect 393 23836 459 23853
rect 393 23802 409 23836
rect 443 23802 459 23836
rect 393 23768 459 23802
rect 393 23734 409 23768
rect 443 23734 459 23768
rect 393 23700 459 23734
rect 393 23666 409 23700
rect 443 23666 459 23700
rect 393 23632 459 23666
rect 393 23598 409 23632
rect 443 23598 459 23632
rect 393 23581 459 23598
rect 489 23836 555 23853
rect 489 23802 505 23836
rect 539 23802 555 23836
rect 489 23768 555 23802
rect 489 23734 505 23768
rect 539 23734 555 23768
rect 489 23700 555 23734
rect 489 23666 505 23700
rect 539 23666 555 23700
rect 489 23632 555 23666
rect 489 23598 505 23632
rect 539 23598 555 23632
rect 489 23581 555 23598
rect 585 23836 651 23853
rect 585 23802 601 23836
rect 635 23802 651 23836
rect 585 23768 651 23802
rect 585 23734 601 23768
rect 635 23734 651 23768
rect 585 23700 651 23734
rect 585 23666 601 23700
rect 635 23666 651 23700
rect 585 23632 651 23666
rect 585 23598 601 23632
rect 635 23598 651 23632
rect 585 23581 651 23598
rect 681 23836 747 23853
rect 681 23802 697 23836
rect 731 23802 747 23836
rect 681 23768 747 23802
rect 681 23734 697 23768
rect 731 23734 747 23768
rect 681 23700 747 23734
rect 681 23666 697 23700
rect 731 23666 747 23700
rect 681 23632 747 23666
rect 681 23598 697 23632
rect 731 23598 747 23632
rect 681 23581 747 23598
rect 777 23836 843 23853
rect 777 23802 793 23836
rect 827 23802 843 23836
rect 777 23768 843 23802
rect 777 23734 793 23768
rect 827 23734 843 23768
rect 777 23700 843 23734
rect 777 23666 793 23700
rect 827 23666 843 23700
rect 777 23632 843 23666
rect 777 23598 793 23632
rect 827 23598 843 23632
rect 777 23581 843 23598
rect 873 23836 939 23853
rect 873 23802 889 23836
rect 923 23802 939 23836
rect 873 23768 939 23802
rect 873 23734 889 23768
rect 923 23734 939 23768
rect 873 23700 939 23734
rect 873 23666 889 23700
rect 923 23666 939 23700
rect 873 23632 939 23666
rect 873 23598 889 23632
rect 923 23598 939 23632
rect 873 23581 939 23598
rect 969 23836 1035 23853
rect 969 23802 985 23836
rect 1019 23802 1035 23836
rect 969 23768 1035 23802
rect 969 23734 985 23768
rect 1019 23734 1035 23768
rect 969 23700 1035 23734
rect 969 23666 985 23700
rect 1019 23666 1035 23700
rect 969 23632 1035 23666
rect 969 23598 985 23632
rect 1019 23598 1035 23632
rect 969 23581 1035 23598
rect 1065 23836 1131 23853
rect 1065 23802 1081 23836
rect 1115 23802 1131 23836
rect 1065 23768 1131 23802
rect 1065 23734 1081 23768
rect 1115 23734 1131 23768
rect 1065 23700 1131 23734
rect 1065 23666 1081 23700
rect 1115 23666 1131 23700
rect 1065 23632 1131 23666
rect 1065 23598 1081 23632
rect 1115 23598 1131 23632
rect 1065 23581 1131 23598
rect 1161 23836 1227 23853
rect 1161 23802 1177 23836
rect 1211 23802 1227 23836
rect 1161 23768 1227 23802
rect 1161 23734 1177 23768
rect 1211 23734 1227 23768
rect 1161 23700 1227 23734
rect 1161 23666 1177 23700
rect 1211 23666 1227 23700
rect 1161 23632 1227 23666
rect 1161 23598 1177 23632
rect 1211 23598 1227 23632
rect 1161 23581 1227 23598
rect 1257 23836 1319 23853
rect 1257 23802 1273 23836
rect 1307 23802 1319 23836
rect 1257 23768 1319 23802
rect 1257 23734 1273 23768
rect 1307 23734 1319 23768
rect 1257 23700 1319 23734
rect 1257 23666 1273 23700
rect 1307 23666 1319 23700
rect 1257 23632 1319 23666
rect 1257 23598 1273 23632
rect 1307 23598 1319 23632
rect 1257 23581 1319 23598
rect 2454 23840 2516 23857
rect 2454 23806 2466 23840
rect 2500 23806 2516 23840
rect 2454 23772 2516 23806
rect 2454 23738 2466 23772
rect 2500 23738 2516 23772
rect 2454 23704 2516 23738
rect 2454 23670 2466 23704
rect 2500 23670 2516 23704
rect 2454 23636 2516 23670
rect 2454 23602 2466 23636
rect 2500 23602 2516 23636
rect 2454 23585 2516 23602
rect 2546 23840 2612 23857
rect 2546 23806 2562 23840
rect 2596 23806 2612 23840
rect 2546 23772 2612 23806
rect 2546 23738 2562 23772
rect 2596 23738 2612 23772
rect 2546 23704 2612 23738
rect 2546 23670 2562 23704
rect 2596 23670 2612 23704
rect 2546 23636 2612 23670
rect 2546 23602 2562 23636
rect 2596 23602 2612 23636
rect 2546 23585 2612 23602
rect 2642 23840 2708 23857
rect 2642 23806 2658 23840
rect 2692 23806 2708 23840
rect 2642 23772 2708 23806
rect 2642 23738 2658 23772
rect 2692 23738 2708 23772
rect 2642 23704 2708 23738
rect 2642 23670 2658 23704
rect 2692 23670 2708 23704
rect 2642 23636 2708 23670
rect 2642 23602 2658 23636
rect 2692 23602 2708 23636
rect 2642 23585 2708 23602
rect 2738 23840 2804 23857
rect 2738 23806 2754 23840
rect 2788 23806 2804 23840
rect 2738 23772 2804 23806
rect 2738 23738 2754 23772
rect 2788 23738 2804 23772
rect 2738 23704 2804 23738
rect 2738 23670 2754 23704
rect 2788 23670 2804 23704
rect 2738 23636 2804 23670
rect 2738 23602 2754 23636
rect 2788 23602 2804 23636
rect 2738 23585 2804 23602
rect 2834 23840 2900 23857
rect 2834 23806 2850 23840
rect 2884 23806 2900 23840
rect 2834 23772 2900 23806
rect 2834 23738 2850 23772
rect 2884 23738 2900 23772
rect 2834 23704 2900 23738
rect 2834 23670 2850 23704
rect 2884 23670 2900 23704
rect 2834 23636 2900 23670
rect 2834 23602 2850 23636
rect 2884 23602 2900 23636
rect 2834 23585 2900 23602
rect 2930 23840 2996 23857
rect 2930 23806 2946 23840
rect 2980 23806 2996 23840
rect 2930 23772 2996 23806
rect 2930 23738 2946 23772
rect 2980 23738 2996 23772
rect 2930 23704 2996 23738
rect 2930 23670 2946 23704
rect 2980 23670 2996 23704
rect 2930 23636 2996 23670
rect 2930 23602 2946 23636
rect 2980 23602 2996 23636
rect 2930 23585 2996 23602
rect 3026 23840 3092 23857
rect 3026 23806 3042 23840
rect 3076 23806 3092 23840
rect 3026 23772 3092 23806
rect 3026 23738 3042 23772
rect 3076 23738 3092 23772
rect 3026 23704 3092 23738
rect 3026 23670 3042 23704
rect 3076 23670 3092 23704
rect 3026 23636 3092 23670
rect 3026 23602 3042 23636
rect 3076 23602 3092 23636
rect 3026 23585 3092 23602
rect 3122 23840 3188 23857
rect 3122 23806 3138 23840
rect 3172 23806 3188 23840
rect 3122 23772 3188 23806
rect 3122 23738 3138 23772
rect 3172 23738 3188 23772
rect 3122 23704 3188 23738
rect 3122 23670 3138 23704
rect 3172 23670 3188 23704
rect 3122 23636 3188 23670
rect 3122 23602 3138 23636
rect 3172 23602 3188 23636
rect 3122 23585 3188 23602
rect 3218 23840 3284 23857
rect 3218 23806 3234 23840
rect 3268 23806 3284 23840
rect 3218 23772 3284 23806
rect 3218 23738 3234 23772
rect 3268 23738 3284 23772
rect 3218 23704 3284 23738
rect 3218 23670 3234 23704
rect 3268 23670 3284 23704
rect 3218 23636 3284 23670
rect 3218 23602 3234 23636
rect 3268 23602 3284 23636
rect 3218 23585 3284 23602
rect 3314 23840 3380 23857
rect 3314 23806 3330 23840
rect 3364 23806 3380 23840
rect 3314 23772 3380 23806
rect 3314 23738 3330 23772
rect 3364 23738 3380 23772
rect 3314 23704 3380 23738
rect 3314 23670 3330 23704
rect 3364 23670 3380 23704
rect 3314 23636 3380 23670
rect 3314 23602 3330 23636
rect 3364 23602 3380 23636
rect 3314 23585 3380 23602
rect 3410 23840 3472 23857
rect 3410 23806 3426 23840
rect 3460 23806 3472 23840
rect 3410 23772 3472 23806
rect 3410 23738 3426 23772
rect 3460 23738 3472 23772
rect 3410 23704 3472 23738
rect 3410 23670 3426 23704
rect 3460 23670 3472 23704
rect 3410 23636 3472 23670
rect 3410 23602 3426 23636
rect 3460 23602 3472 23636
rect 3410 23585 3472 23602
rect 3975 23840 4037 23857
rect 3975 23806 3987 23840
rect 4021 23806 4037 23840
rect 3975 23772 4037 23806
rect 3975 23738 3987 23772
rect 4021 23738 4037 23772
rect 3975 23704 4037 23738
rect 3975 23670 3987 23704
rect 4021 23670 4037 23704
rect 3975 23636 4037 23670
rect 3975 23602 3987 23636
rect 4021 23602 4037 23636
rect 3975 23585 4037 23602
rect 4067 23840 4133 23857
rect 4067 23806 4083 23840
rect 4117 23806 4133 23840
rect 4067 23772 4133 23806
rect 4067 23738 4083 23772
rect 4117 23738 4133 23772
rect 4067 23704 4133 23738
rect 4067 23670 4083 23704
rect 4117 23670 4133 23704
rect 4067 23636 4133 23670
rect 4067 23602 4083 23636
rect 4117 23602 4133 23636
rect 4067 23585 4133 23602
rect 4163 23840 4229 23857
rect 4163 23806 4179 23840
rect 4213 23806 4229 23840
rect 4163 23772 4229 23806
rect 4163 23738 4179 23772
rect 4213 23738 4229 23772
rect 4163 23704 4229 23738
rect 4163 23670 4179 23704
rect 4213 23670 4229 23704
rect 4163 23636 4229 23670
rect 4163 23602 4179 23636
rect 4213 23602 4229 23636
rect 4163 23585 4229 23602
rect 4259 23840 4325 23857
rect 4259 23806 4275 23840
rect 4309 23806 4325 23840
rect 4259 23772 4325 23806
rect 4259 23738 4275 23772
rect 4309 23738 4325 23772
rect 4259 23704 4325 23738
rect 4259 23670 4275 23704
rect 4309 23670 4325 23704
rect 4259 23636 4325 23670
rect 4259 23602 4275 23636
rect 4309 23602 4325 23636
rect 4259 23585 4325 23602
rect 4355 23840 4421 23857
rect 4355 23806 4371 23840
rect 4405 23806 4421 23840
rect 4355 23772 4421 23806
rect 4355 23738 4371 23772
rect 4405 23738 4421 23772
rect 4355 23704 4421 23738
rect 4355 23670 4371 23704
rect 4405 23670 4421 23704
rect 4355 23636 4421 23670
rect 4355 23602 4371 23636
rect 4405 23602 4421 23636
rect 4355 23585 4421 23602
rect 4451 23840 4517 23857
rect 4451 23806 4467 23840
rect 4501 23806 4517 23840
rect 4451 23772 4517 23806
rect 4451 23738 4467 23772
rect 4501 23738 4517 23772
rect 4451 23704 4517 23738
rect 4451 23670 4467 23704
rect 4501 23670 4517 23704
rect 4451 23636 4517 23670
rect 4451 23602 4467 23636
rect 4501 23602 4517 23636
rect 4451 23585 4517 23602
rect 4547 23840 4613 23857
rect 4547 23806 4563 23840
rect 4597 23806 4613 23840
rect 4547 23772 4613 23806
rect 4547 23738 4563 23772
rect 4597 23738 4613 23772
rect 4547 23704 4613 23738
rect 4547 23670 4563 23704
rect 4597 23670 4613 23704
rect 4547 23636 4613 23670
rect 4547 23602 4563 23636
rect 4597 23602 4613 23636
rect 4547 23585 4613 23602
rect 4643 23840 4709 23857
rect 4643 23806 4659 23840
rect 4693 23806 4709 23840
rect 4643 23772 4709 23806
rect 4643 23738 4659 23772
rect 4693 23738 4709 23772
rect 4643 23704 4709 23738
rect 4643 23670 4659 23704
rect 4693 23670 4709 23704
rect 4643 23636 4709 23670
rect 4643 23602 4659 23636
rect 4693 23602 4709 23636
rect 4643 23585 4709 23602
rect 4739 23840 4805 23857
rect 4739 23806 4755 23840
rect 4789 23806 4805 23840
rect 4739 23772 4805 23806
rect 4739 23738 4755 23772
rect 4789 23738 4805 23772
rect 4739 23704 4805 23738
rect 4739 23670 4755 23704
rect 4789 23670 4805 23704
rect 4739 23636 4805 23670
rect 4739 23602 4755 23636
rect 4789 23602 4805 23636
rect 4739 23585 4805 23602
rect 4835 23840 4901 23857
rect 4835 23806 4851 23840
rect 4885 23806 4901 23840
rect 4835 23772 4901 23806
rect 4835 23738 4851 23772
rect 4885 23738 4901 23772
rect 4835 23704 4901 23738
rect 4835 23670 4851 23704
rect 4885 23670 4901 23704
rect 4835 23636 4901 23670
rect 4835 23602 4851 23636
rect 4885 23602 4901 23636
rect 4835 23585 4901 23602
rect 4931 23840 4993 23857
rect 4931 23806 4947 23840
rect 4981 23806 4993 23840
rect 4931 23772 4993 23806
rect 4931 23738 4947 23772
rect 4981 23738 4993 23772
rect 4931 23704 4993 23738
rect 4931 23670 4947 23704
rect 4981 23670 4993 23704
rect 4931 23636 4993 23670
rect 4931 23602 4947 23636
rect 4981 23602 4993 23636
rect 4931 23585 4993 23602
rect 5348 23632 5400 23644
rect 5348 23598 5356 23632
rect 5390 23598 5400 23632
rect 5348 23564 5400 23598
rect 5348 23530 5356 23564
rect 5390 23530 5400 23564
rect 5348 23496 5400 23530
rect 5348 23462 5356 23496
rect 5390 23462 5400 23496
rect 5348 23444 5400 23462
rect 5430 23632 5482 23644
rect 5430 23598 5440 23632
rect 5474 23598 5482 23632
rect 5430 23564 5482 23598
rect 5430 23530 5440 23564
rect 5474 23530 5482 23564
rect 5430 23496 5482 23530
rect 5430 23462 5440 23496
rect 5474 23462 5482 23496
rect 5430 23444 5482 23462
rect 301 22549 363 22566
rect 301 22515 313 22549
rect 347 22515 363 22549
rect 301 22481 363 22515
rect 301 22447 313 22481
rect 347 22447 363 22481
rect 301 22413 363 22447
rect 301 22379 313 22413
rect 347 22379 363 22413
rect 301 22345 363 22379
rect 301 22311 313 22345
rect 347 22311 363 22345
rect 301 22294 363 22311
rect 393 22549 459 22566
rect 393 22515 409 22549
rect 443 22515 459 22549
rect 393 22481 459 22515
rect 393 22447 409 22481
rect 443 22447 459 22481
rect 393 22413 459 22447
rect 393 22379 409 22413
rect 443 22379 459 22413
rect 393 22345 459 22379
rect 393 22311 409 22345
rect 443 22311 459 22345
rect 393 22294 459 22311
rect 489 22549 555 22566
rect 489 22515 505 22549
rect 539 22515 555 22549
rect 489 22481 555 22515
rect 489 22447 505 22481
rect 539 22447 555 22481
rect 489 22413 555 22447
rect 489 22379 505 22413
rect 539 22379 555 22413
rect 489 22345 555 22379
rect 489 22311 505 22345
rect 539 22311 555 22345
rect 489 22294 555 22311
rect 585 22549 651 22566
rect 585 22515 601 22549
rect 635 22515 651 22549
rect 585 22481 651 22515
rect 585 22447 601 22481
rect 635 22447 651 22481
rect 585 22413 651 22447
rect 585 22379 601 22413
rect 635 22379 651 22413
rect 585 22345 651 22379
rect 585 22311 601 22345
rect 635 22311 651 22345
rect 585 22294 651 22311
rect 681 22549 747 22566
rect 681 22515 697 22549
rect 731 22515 747 22549
rect 681 22481 747 22515
rect 681 22447 697 22481
rect 731 22447 747 22481
rect 681 22413 747 22447
rect 681 22379 697 22413
rect 731 22379 747 22413
rect 681 22345 747 22379
rect 681 22311 697 22345
rect 731 22311 747 22345
rect 681 22294 747 22311
rect 777 22549 843 22566
rect 777 22515 793 22549
rect 827 22515 843 22549
rect 777 22481 843 22515
rect 777 22447 793 22481
rect 827 22447 843 22481
rect 777 22413 843 22447
rect 777 22379 793 22413
rect 827 22379 843 22413
rect 777 22345 843 22379
rect 777 22311 793 22345
rect 827 22311 843 22345
rect 777 22294 843 22311
rect 873 22549 939 22566
rect 873 22515 889 22549
rect 923 22515 939 22549
rect 873 22481 939 22515
rect 873 22447 889 22481
rect 923 22447 939 22481
rect 873 22413 939 22447
rect 873 22379 889 22413
rect 923 22379 939 22413
rect 873 22345 939 22379
rect 873 22311 889 22345
rect 923 22311 939 22345
rect 873 22294 939 22311
rect 969 22549 1035 22566
rect 969 22515 985 22549
rect 1019 22515 1035 22549
rect 969 22481 1035 22515
rect 969 22447 985 22481
rect 1019 22447 1035 22481
rect 969 22413 1035 22447
rect 969 22379 985 22413
rect 1019 22379 1035 22413
rect 969 22345 1035 22379
rect 969 22311 985 22345
rect 1019 22311 1035 22345
rect 969 22294 1035 22311
rect 1065 22549 1131 22566
rect 1065 22515 1081 22549
rect 1115 22515 1131 22549
rect 1065 22481 1131 22515
rect 1065 22447 1081 22481
rect 1115 22447 1131 22481
rect 1065 22413 1131 22447
rect 1065 22379 1081 22413
rect 1115 22379 1131 22413
rect 1065 22345 1131 22379
rect 1065 22311 1081 22345
rect 1115 22311 1131 22345
rect 1065 22294 1131 22311
rect 1161 22549 1227 22566
rect 1161 22515 1177 22549
rect 1211 22515 1227 22549
rect 1161 22481 1227 22515
rect 1161 22447 1177 22481
rect 1211 22447 1227 22481
rect 1161 22413 1227 22447
rect 1161 22379 1177 22413
rect 1211 22379 1227 22413
rect 1161 22345 1227 22379
rect 1161 22311 1177 22345
rect 1211 22311 1227 22345
rect 1161 22294 1227 22311
rect 1257 22549 1319 22566
rect 1257 22515 1273 22549
rect 1307 22515 1319 22549
rect 1257 22481 1319 22515
rect 1257 22447 1273 22481
rect 1307 22447 1319 22481
rect 1257 22413 1319 22447
rect 1257 22379 1273 22413
rect 1307 22379 1319 22413
rect 1257 22345 1319 22379
rect 1257 22311 1273 22345
rect 1307 22311 1319 22345
rect 1257 22294 1319 22311
rect 2454 22553 2516 22570
rect 2454 22519 2466 22553
rect 2500 22519 2516 22553
rect 2454 22485 2516 22519
rect 2454 22451 2466 22485
rect 2500 22451 2516 22485
rect 2454 22417 2516 22451
rect 2454 22383 2466 22417
rect 2500 22383 2516 22417
rect 2454 22349 2516 22383
rect 2454 22315 2466 22349
rect 2500 22315 2516 22349
rect 2454 22298 2516 22315
rect 2546 22553 2612 22570
rect 2546 22519 2562 22553
rect 2596 22519 2612 22553
rect 2546 22485 2612 22519
rect 2546 22451 2562 22485
rect 2596 22451 2612 22485
rect 2546 22417 2612 22451
rect 2546 22383 2562 22417
rect 2596 22383 2612 22417
rect 2546 22349 2612 22383
rect 2546 22315 2562 22349
rect 2596 22315 2612 22349
rect 2546 22298 2612 22315
rect 2642 22553 2708 22570
rect 2642 22519 2658 22553
rect 2692 22519 2708 22553
rect 2642 22485 2708 22519
rect 2642 22451 2658 22485
rect 2692 22451 2708 22485
rect 2642 22417 2708 22451
rect 2642 22383 2658 22417
rect 2692 22383 2708 22417
rect 2642 22349 2708 22383
rect 2642 22315 2658 22349
rect 2692 22315 2708 22349
rect 2642 22298 2708 22315
rect 2738 22553 2804 22570
rect 2738 22519 2754 22553
rect 2788 22519 2804 22553
rect 2738 22485 2804 22519
rect 2738 22451 2754 22485
rect 2788 22451 2804 22485
rect 2738 22417 2804 22451
rect 2738 22383 2754 22417
rect 2788 22383 2804 22417
rect 2738 22349 2804 22383
rect 2738 22315 2754 22349
rect 2788 22315 2804 22349
rect 2738 22298 2804 22315
rect 2834 22553 2900 22570
rect 2834 22519 2850 22553
rect 2884 22519 2900 22553
rect 2834 22485 2900 22519
rect 2834 22451 2850 22485
rect 2884 22451 2900 22485
rect 2834 22417 2900 22451
rect 2834 22383 2850 22417
rect 2884 22383 2900 22417
rect 2834 22349 2900 22383
rect 2834 22315 2850 22349
rect 2884 22315 2900 22349
rect 2834 22298 2900 22315
rect 2930 22553 2996 22570
rect 2930 22519 2946 22553
rect 2980 22519 2996 22553
rect 2930 22485 2996 22519
rect 2930 22451 2946 22485
rect 2980 22451 2996 22485
rect 2930 22417 2996 22451
rect 2930 22383 2946 22417
rect 2980 22383 2996 22417
rect 2930 22349 2996 22383
rect 2930 22315 2946 22349
rect 2980 22315 2996 22349
rect 2930 22298 2996 22315
rect 3026 22553 3092 22570
rect 3026 22519 3042 22553
rect 3076 22519 3092 22553
rect 3026 22485 3092 22519
rect 3026 22451 3042 22485
rect 3076 22451 3092 22485
rect 3026 22417 3092 22451
rect 3026 22383 3042 22417
rect 3076 22383 3092 22417
rect 3026 22349 3092 22383
rect 3026 22315 3042 22349
rect 3076 22315 3092 22349
rect 3026 22298 3092 22315
rect 3122 22553 3188 22570
rect 3122 22519 3138 22553
rect 3172 22519 3188 22553
rect 3122 22485 3188 22519
rect 3122 22451 3138 22485
rect 3172 22451 3188 22485
rect 3122 22417 3188 22451
rect 3122 22383 3138 22417
rect 3172 22383 3188 22417
rect 3122 22349 3188 22383
rect 3122 22315 3138 22349
rect 3172 22315 3188 22349
rect 3122 22298 3188 22315
rect 3218 22553 3284 22570
rect 3218 22519 3234 22553
rect 3268 22519 3284 22553
rect 3218 22485 3284 22519
rect 3218 22451 3234 22485
rect 3268 22451 3284 22485
rect 3218 22417 3284 22451
rect 3218 22383 3234 22417
rect 3268 22383 3284 22417
rect 3218 22349 3284 22383
rect 3218 22315 3234 22349
rect 3268 22315 3284 22349
rect 3218 22298 3284 22315
rect 3314 22553 3380 22570
rect 3314 22519 3330 22553
rect 3364 22519 3380 22553
rect 3314 22485 3380 22519
rect 3314 22451 3330 22485
rect 3364 22451 3380 22485
rect 3314 22417 3380 22451
rect 3314 22383 3330 22417
rect 3364 22383 3380 22417
rect 3314 22349 3380 22383
rect 3314 22315 3330 22349
rect 3364 22315 3380 22349
rect 3314 22298 3380 22315
rect 3410 22553 3472 22570
rect 3410 22519 3426 22553
rect 3460 22519 3472 22553
rect 3410 22485 3472 22519
rect 3410 22451 3426 22485
rect 3460 22451 3472 22485
rect 3410 22417 3472 22451
rect 3410 22383 3426 22417
rect 3460 22383 3472 22417
rect 3410 22349 3472 22383
rect 3410 22315 3426 22349
rect 3460 22315 3472 22349
rect 3410 22298 3472 22315
rect 3975 22553 4037 22570
rect 3975 22519 3987 22553
rect 4021 22519 4037 22553
rect 3975 22485 4037 22519
rect 3975 22451 3987 22485
rect 4021 22451 4037 22485
rect 3975 22417 4037 22451
rect 3975 22383 3987 22417
rect 4021 22383 4037 22417
rect 3975 22349 4037 22383
rect 3975 22315 3987 22349
rect 4021 22315 4037 22349
rect 3975 22298 4037 22315
rect 4067 22553 4133 22570
rect 4067 22519 4083 22553
rect 4117 22519 4133 22553
rect 4067 22485 4133 22519
rect 4067 22451 4083 22485
rect 4117 22451 4133 22485
rect 4067 22417 4133 22451
rect 4067 22383 4083 22417
rect 4117 22383 4133 22417
rect 4067 22349 4133 22383
rect 4067 22315 4083 22349
rect 4117 22315 4133 22349
rect 4067 22298 4133 22315
rect 4163 22553 4229 22570
rect 4163 22519 4179 22553
rect 4213 22519 4229 22553
rect 4163 22485 4229 22519
rect 4163 22451 4179 22485
rect 4213 22451 4229 22485
rect 4163 22417 4229 22451
rect 4163 22383 4179 22417
rect 4213 22383 4229 22417
rect 4163 22349 4229 22383
rect 4163 22315 4179 22349
rect 4213 22315 4229 22349
rect 4163 22298 4229 22315
rect 4259 22553 4325 22570
rect 4259 22519 4275 22553
rect 4309 22519 4325 22553
rect 4259 22485 4325 22519
rect 4259 22451 4275 22485
rect 4309 22451 4325 22485
rect 4259 22417 4325 22451
rect 4259 22383 4275 22417
rect 4309 22383 4325 22417
rect 4259 22349 4325 22383
rect 4259 22315 4275 22349
rect 4309 22315 4325 22349
rect 4259 22298 4325 22315
rect 4355 22553 4421 22570
rect 4355 22519 4371 22553
rect 4405 22519 4421 22553
rect 4355 22485 4421 22519
rect 4355 22451 4371 22485
rect 4405 22451 4421 22485
rect 4355 22417 4421 22451
rect 4355 22383 4371 22417
rect 4405 22383 4421 22417
rect 4355 22349 4421 22383
rect 4355 22315 4371 22349
rect 4405 22315 4421 22349
rect 4355 22298 4421 22315
rect 4451 22553 4517 22570
rect 4451 22519 4467 22553
rect 4501 22519 4517 22553
rect 4451 22485 4517 22519
rect 4451 22451 4467 22485
rect 4501 22451 4517 22485
rect 4451 22417 4517 22451
rect 4451 22383 4467 22417
rect 4501 22383 4517 22417
rect 4451 22349 4517 22383
rect 4451 22315 4467 22349
rect 4501 22315 4517 22349
rect 4451 22298 4517 22315
rect 4547 22553 4613 22570
rect 4547 22519 4563 22553
rect 4597 22519 4613 22553
rect 4547 22485 4613 22519
rect 4547 22451 4563 22485
rect 4597 22451 4613 22485
rect 4547 22417 4613 22451
rect 4547 22383 4563 22417
rect 4597 22383 4613 22417
rect 4547 22349 4613 22383
rect 4547 22315 4563 22349
rect 4597 22315 4613 22349
rect 4547 22298 4613 22315
rect 4643 22553 4709 22570
rect 4643 22519 4659 22553
rect 4693 22519 4709 22553
rect 4643 22485 4709 22519
rect 4643 22451 4659 22485
rect 4693 22451 4709 22485
rect 4643 22417 4709 22451
rect 4643 22383 4659 22417
rect 4693 22383 4709 22417
rect 4643 22349 4709 22383
rect 4643 22315 4659 22349
rect 4693 22315 4709 22349
rect 4643 22298 4709 22315
rect 4739 22553 4805 22570
rect 4739 22519 4755 22553
rect 4789 22519 4805 22553
rect 4739 22485 4805 22519
rect 4739 22451 4755 22485
rect 4789 22451 4805 22485
rect 4739 22417 4805 22451
rect 4739 22383 4755 22417
rect 4789 22383 4805 22417
rect 4739 22349 4805 22383
rect 4739 22315 4755 22349
rect 4789 22315 4805 22349
rect 4739 22298 4805 22315
rect 4835 22553 4901 22570
rect 4835 22519 4851 22553
rect 4885 22519 4901 22553
rect 4835 22485 4901 22519
rect 4835 22451 4851 22485
rect 4885 22451 4901 22485
rect 4835 22417 4901 22451
rect 4835 22383 4851 22417
rect 4885 22383 4901 22417
rect 4835 22349 4901 22383
rect 4835 22315 4851 22349
rect 4885 22315 4901 22349
rect 4835 22298 4901 22315
rect 4931 22553 4993 22570
rect 4931 22519 4947 22553
rect 4981 22519 4993 22553
rect 4931 22485 4993 22519
rect 4931 22451 4947 22485
rect 4981 22451 4993 22485
rect 4931 22417 4993 22451
rect 4931 22383 4947 22417
rect 4981 22383 4993 22417
rect 4931 22349 4993 22383
rect 4931 22315 4947 22349
rect 4981 22315 4993 22349
rect 4931 22298 4993 22315
rect 5348 22345 5400 22357
rect 5348 22311 5356 22345
rect 5390 22311 5400 22345
rect 5348 22277 5400 22311
rect 5348 22243 5356 22277
rect 5390 22243 5400 22277
rect 5348 22209 5400 22243
rect 5348 22175 5356 22209
rect 5390 22175 5400 22209
rect 5348 22157 5400 22175
rect 5430 22345 5482 22357
rect 5430 22311 5440 22345
rect 5474 22311 5482 22345
rect 5430 22277 5482 22311
rect 5430 22243 5440 22277
rect 5474 22243 5482 22277
rect 5430 22209 5482 22243
rect 5430 22175 5440 22209
rect 5474 22175 5482 22209
rect 5430 22157 5482 22175
rect 301 21262 363 21279
rect 301 21228 313 21262
rect 347 21228 363 21262
rect 301 21194 363 21228
rect 301 21160 313 21194
rect 347 21160 363 21194
rect 301 21126 363 21160
rect 301 21092 313 21126
rect 347 21092 363 21126
rect 301 21058 363 21092
rect 301 21024 313 21058
rect 347 21024 363 21058
rect 301 21007 363 21024
rect 393 21262 459 21279
rect 393 21228 409 21262
rect 443 21228 459 21262
rect 393 21194 459 21228
rect 393 21160 409 21194
rect 443 21160 459 21194
rect 393 21126 459 21160
rect 393 21092 409 21126
rect 443 21092 459 21126
rect 393 21058 459 21092
rect 393 21024 409 21058
rect 443 21024 459 21058
rect 393 21007 459 21024
rect 489 21262 555 21279
rect 489 21228 505 21262
rect 539 21228 555 21262
rect 489 21194 555 21228
rect 489 21160 505 21194
rect 539 21160 555 21194
rect 489 21126 555 21160
rect 489 21092 505 21126
rect 539 21092 555 21126
rect 489 21058 555 21092
rect 489 21024 505 21058
rect 539 21024 555 21058
rect 489 21007 555 21024
rect 585 21262 651 21279
rect 585 21228 601 21262
rect 635 21228 651 21262
rect 585 21194 651 21228
rect 585 21160 601 21194
rect 635 21160 651 21194
rect 585 21126 651 21160
rect 585 21092 601 21126
rect 635 21092 651 21126
rect 585 21058 651 21092
rect 585 21024 601 21058
rect 635 21024 651 21058
rect 585 21007 651 21024
rect 681 21262 747 21279
rect 681 21228 697 21262
rect 731 21228 747 21262
rect 681 21194 747 21228
rect 681 21160 697 21194
rect 731 21160 747 21194
rect 681 21126 747 21160
rect 681 21092 697 21126
rect 731 21092 747 21126
rect 681 21058 747 21092
rect 681 21024 697 21058
rect 731 21024 747 21058
rect 681 21007 747 21024
rect 777 21262 843 21279
rect 777 21228 793 21262
rect 827 21228 843 21262
rect 777 21194 843 21228
rect 777 21160 793 21194
rect 827 21160 843 21194
rect 777 21126 843 21160
rect 777 21092 793 21126
rect 827 21092 843 21126
rect 777 21058 843 21092
rect 777 21024 793 21058
rect 827 21024 843 21058
rect 777 21007 843 21024
rect 873 21262 939 21279
rect 873 21228 889 21262
rect 923 21228 939 21262
rect 873 21194 939 21228
rect 873 21160 889 21194
rect 923 21160 939 21194
rect 873 21126 939 21160
rect 873 21092 889 21126
rect 923 21092 939 21126
rect 873 21058 939 21092
rect 873 21024 889 21058
rect 923 21024 939 21058
rect 873 21007 939 21024
rect 969 21262 1035 21279
rect 969 21228 985 21262
rect 1019 21228 1035 21262
rect 969 21194 1035 21228
rect 969 21160 985 21194
rect 1019 21160 1035 21194
rect 969 21126 1035 21160
rect 969 21092 985 21126
rect 1019 21092 1035 21126
rect 969 21058 1035 21092
rect 969 21024 985 21058
rect 1019 21024 1035 21058
rect 969 21007 1035 21024
rect 1065 21262 1131 21279
rect 1065 21228 1081 21262
rect 1115 21228 1131 21262
rect 1065 21194 1131 21228
rect 1065 21160 1081 21194
rect 1115 21160 1131 21194
rect 1065 21126 1131 21160
rect 1065 21092 1081 21126
rect 1115 21092 1131 21126
rect 1065 21058 1131 21092
rect 1065 21024 1081 21058
rect 1115 21024 1131 21058
rect 1065 21007 1131 21024
rect 1161 21262 1227 21279
rect 1161 21228 1177 21262
rect 1211 21228 1227 21262
rect 1161 21194 1227 21228
rect 1161 21160 1177 21194
rect 1211 21160 1227 21194
rect 1161 21126 1227 21160
rect 1161 21092 1177 21126
rect 1211 21092 1227 21126
rect 1161 21058 1227 21092
rect 1161 21024 1177 21058
rect 1211 21024 1227 21058
rect 1161 21007 1227 21024
rect 1257 21262 1319 21279
rect 1257 21228 1273 21262
rect 1307 21228 1319 21262
rect 1257 21194 1319 21228
rect 1257 21160 1273 21194
rect 1307 21160 1319 21194
rect 1257 21126 1319 21160
rect 1257 21092 1273 21126
rect 1307 21092 1319 21126
rect 1257 21058 1319 21092
rect 1257 21024 1273 21058
rect 1307 21024 1319 21058
rect 1257 21007 1319 21024
rect 2454 21266 2516 21283
rect 2454 21232 2466 21266
rect 2500 21232 2516 21266
rect 2454 21198 2516 21232
rect 2454 21164 2466 21198
rect 2500 21164 2516 21198
rect 2454 21130 2516 21164
rect 2454 21096 2466 21130
rect 2500 21096 2516 21130
rect 2454 21062 2516 21096
rect 2454 21028 2466 21062
rect 2500 21028 2516 21062
rect 2454 21011 2516 21028
rect 2546 21266 2612 21283
rect 2546 21232 2562 21266
rect 2596 21232 2612 21266
rect 2546 21198 2612 21232
rect 2546 21164 2562 21198
rect 2596 21164 2612 21198
rect 2546 21130 2612 21164
rect 2546 21096 2562 21130
rect 2596 21096 2612 21130
rect 2546 21062 2612 21096
rect 2546 21028 2562 21062
rect 2596 21028 2612 21062
rect 2546 21011 2612 21028
rect 2642 21266 2708 21283
rect 2642 21232 2658 21266
rect 2692 21232 2708 21266
rect 2642 21198 2708 21232
rect 2642 21164 2658 21198
rect 2692 21164 2708 21198
rect 2642 21130 2708 21164
rect 2642 21096 2658 21130
rect 2692 21096 2708 21130
rect 2642 21062 2708 21096
rect 2642 21028 2658 21062
rect 2692 21028 2708 21062
rect 2642 21011 2708 21028
rect 2738 21266 2804 21283
rect 2738 21232 2754 21266
rect 2788 21232 2804 21266
rect 2738 21198 2804 21232
rect 2738 21164 2754 21198
rect 2788 21164 2804 21198
rect 2738 21130 2804 21164
rect 2738 21096 2754 21130
rect 2788 21096 2804 21130
rect 2738 21062 2804 21096
rect 2738 21028 2754 21062
rect 2788 21028 2804 21062
rect 2738 21011 2804 21028
rect 2834 21266 2900 21283
rect 2834 21232 2850 21266
rect 2884 21232 2900 21266
rect 2834 21198 2900 21232
rect 2834 21164 2850 21198
rect 2884 21164 2900 21198
rect 2834 21130 2900 21164
rect 2834 21096 2850 21130
rect 2884 21096 2900 21130
rect 2834 21062 2900 21096
rect 2834 21028 2850 21062
rect 2884 21028 2900 21062
rect 2834 21011 2900 21028
rect 2930 21266 2996 21283
rect 2930 21232 2946 21266
rect 2980 21232 2996 21266
rect 2930 21198 2996 21232
rect 2930 21164 2946 21198
rect 2980 21164 2996 21198
rect 2930 21130 2996 21164
rect 2930 21096 2946 21130
rect 2980 21096 2996 21130
rect 2930 21062 2996 21096
rect 2930 21028 2946 21062
rect 2980 21028 2996 21062
rect 2930 21011 2996 21028
rect 3026 21266 3092 21283
rect 3026 21232 3042 21266
rect 3076 21232 3092 21266
rect 3026 21198 3092 21232
rect 3026 21164 3042 21198
rect 3076 21164 3092 21198
rect 3026 21130 3092 21164
rect 3026 21096 3042 21130
rect 3076 21096 3092 21130
rect 3026 21062 3092 21096
rect 3026 21028 3042 21062
rect 3076 21028 3092 21062
rect 3026 21011 3092 21028
rect 3122 21266 3188 21283
rect 3122 21232 3138 21266
rect 3172 21232 3188 21266
rect 3122 21198 3188 21232
rect 3122 21164 3138 21198
rect 3172 21164 3188 21198
rect 3122 21130 3188 21164
rect 3122 21096 3138 21130
rect 3172 21096 3188 21130
rect 3122 21062 3188 21096
rect 3122 21028 3138 21062
rect 3172 21028 3188 21062
rect 3122 21011 3188 21028
rect 3218 21266 3284 21283
rect 3218 21232 3234 21266
rect 3268 21232 3284 21266
rect 3218 21198 3284 21232
rect 3218 21164 3234 21198
rect 3268 21164 3284 21198
rect 3218 21130 3284 21164
rect 3218 21096 3234 21130
rect 3268 21096 3284 21130
rect 3218 21062 3284 21096
rect 3218 21028 3234 21062
rect 3268 21028 3284 21062
rect 3218 21011 3284 21028
rect 3314 21266 3380 21283
rect 3314 21232 3330 21266
rect 3364 21232 3380 21266
rect 3314 21198 3380 21232
rect 3314 21164 3330 21198
rect 3364 21164 3380 21198
rect 3314 21130 3380 21164
rect 3314 21096 3330 21130
rect 3364 21096 3380 21130
rect 3314 21062 3380 21096
rect 3314 21028 3330 21062
rect 3364 21028 3380 21062
rect 3314 21011 3380 21028
rect 3410 21266 3472 21283
rect 3410 21232 3426 21266
rect 3460 21232 3472 21266
rect 3410 21198 3472 21232
rect 3410 21164 3426 21198
rect 3460 21164 3472 21198
rect 3410 21130 3472 21164
rect 3410 21096 3426 21130
rect 3460 21096 3472 21130
rect 3410 21062 3472 21096
rect 3410 21028 3426 21062
rect 3460 21028 3472 21062
rect 3410 21011 3472 21028
rect 3975 21266 4037 21283
rect 3975 21232 3987 21266
rect 4021 21232 4037 21266
rect 3975 21198 4037 21232
rect 3975 21164 3987 21198
rect 4021 21164 4037 21198
rect 3975 21130 4037 21164
rect 3975 21096 3987 21130
rect 4021 21096 4037 21130
rect 3975 21062 4037 21096
rect 3975 21028 3987 21062
rect 4021 21028 4037 21062
rect 3975 21011 4037 21028
rect 4067 21266 4133 21283
rect 4067 21232 4083 21266
rect 4117 21232 4133 21266
rect 4067 21198 4133 21232
rect 4067 21164 4083 21198
rect 4117 21164 4133 21198
rect 4067 21130 4133 21164
rect 4067 21096 4083 21130
rect 4117 21096 4133 21130
rect 4067 21062 4133 21096
rect 4067 21028 4083 21062
rect 4117 21028 4133 21062
rect 4067 21011 4133 21028
rect 4163 21266 4229 21283
rect 4163 21232 4179 21266
rect 4213 21232 4229 21266
rect 4163 21198 4229 21232
rect 4163 21164 4179 21198
rect 4213 21164 4229 21198
rect 4163 21130 4229 21164
rect 4163 21096 4179 21130
rect 4213 21096 4229 21130
rect 4163 21062 4229 21096
rect 4163 21028 4179 21062
rect 4213 21028 4229 21062
rect 4163 21011 4229 21028
rect 4259 21266 4325 21283
rect 4259 21232 4275 21266
rect 4309 21232 4325 21266
rect 4259 21198 4325 21232
rect 4259 21164 4275 21198
rect 4309 21164 4325 21198
rect 4259 21130 4325 21164
rect 4259 21096 4275 21130
rect 4309 21096 4325 21130
rect 4259 21062 4325 21096
rect 4259 21028 4275 21062
rect 4309 21028 4325 21062
rect 4259 21011 4325 21028
rect 4355 21266 4421 21283
rect 4355 21232 4371 21266
rect 4405 21232 4421 21266
rect 4355 21198 4421 21232
rect 4355 21164 4371 21198
rect 4405 21164 4421 21198
rect 4355 21130 4421 21164
rect 4355 21096 4371 21130
rect 4405 21096 4421 21130
rect 4355 21062 4421 21096
rect 4355 21028 4371 21062
rect 4405 21028 4421 21062
rect 4355 21011 4421 21028
rect 4451 21266 4517 21283
rect 4451 21232 4467 21266
rect 4501 21232 4517 21266
rect 4451 21198 4517 21232
rect 4451 21164 4467 21198
rect 4501 21164 4517 21198
rect 4451 21130 4517 21164
rect 4451 21096 4467 21130
rect 4501 21096 4517 21130
rect 4451 21062 4517 21096
rect 4451 21028 4467 21062
rect 4501 21028 4517 21062
rect 4451 21011 4517 21028
rect 4547 21266 4613 21283
rect 4547 21232 4563 21266
rect 4597 21232 4613 21266
rect 4547 21198 4613 21232
rect 4547 21164 4563 21198
rect 4597 21164 4613 21198
rect 4547 21130 4613 21164
rect 4547 21096 4563 21130
rect 4597 21096 4613 21130
rect 4547 21062 4613 21096
rect 4547 21028 4563 21062
rect 4597 21028 4613 21062
rect 4547 21011 4613 21028
rect 4643 21266 4709 21283
rect 4643 21232 4659 21266
rect 4693 21232 4709 21266
rect 4643 21198 4709 21232
rect 4643 21164 4659 21198
rect 4693 21164 4709 21198
rect 4643 21130 4709 21164
rect 4643 21096 4659 21130
rect 4693 21096 4709 21130
rect 4643 21062 4709 21096
rect 4643 21028 4659 21062
rect 4693 21028 4709 21062
rect 4643 21011 4709 21028
rect 4739 21266 4805 21283
rect 4739 21232 4755 21266
rect 4789 21232 4805 21266
rect 4739 21198 4805 21232
rect 4739 21164 4755 21198
rect 4789 21164 4805 21198
rect 4739 21130 4805 21164
rect 4739 21096 4755 21130
rect 4789 21096 4805 21130
rect 4739 21062 4805 21096
rect 4739 21028 4755 21062
rect 4789 21028 4805 21062
rect 4739 21011 4805 21028
rect 4835 21266 4901 21283
rect 4835 21232 4851 21266
rect 4885 21232 4901 21266
rect 4835 21198 4901 21232
rect 4835 21164 4851 21198
rect 4885 21164 4901 21198
rect 4835 21130 4901 21164
rect 4835 21096 4851 21130
rect 4885 21096 4901 21130
rect 4835 21062 4901 21096
rect 4835 21028 4851 21062
rect 4885 21028 4901 21062
rect 4835 21011 4901 21028
rect 4931 21266 4993 21283
rect 4931 21232 4947 21266
rect 4981 21232 4993 21266
rect 4931 21198 4993 21232
rect 4931 21164 4947 21198
rect 4981 21164 4993 21198
rect 4931 21130 4993 21164
rect 4931 21096 4947 21130
rect 4981 21096 4993 21130
rect 4931 21062 4993 21096
rect 4931 21028 4947 21062
rect 4981 21028 4993 21062
rect 4931 21011 4993 21028
rect 5348 21058 5400 21070
rect 5348 21024 5356 21058
rect 5390 21024 5400 21058
rect 5348 20990 5400 21024
rect 5348 20956 5356 20990
rect 5390 20956 5400 20990
rect 5348 20922 5400 20956
rect 5348 20888 5356 20922
rect 5390 20888 5400 20922
rect 5348 20870 5400 20888
rect 5430 21058 5482 21070
rect 5430 21024 5440 21058
rect 5474 21024 5482 21058
rect 5430 20990 5482 21024
rect 5430 20956 5440 20990
rect 5474 20956 5482 20990
rect 5430 20922 5482 20956
rect 5430 20888 5440 20922
rect 5474 20888 5482 20922
rect 5430 20870 5482 20888
rect 301 19975 363 19992
rect 301 19941 313 19975
rect 347 19941 363 19975
rect 301 19907 363 19941
rect 301 19873 313 19907
rect 347 19873 363 19907
rect 301 19839 363 19873
rect 301 19805 313 19839
rect 347 19805 363 19839
rect 301 19771 363 19805
rect 301 19737 313 19771
rect 347 19737 363 19771
rect 301 19720 363 19737
rect 393 19975 459 19992
rect 393 19941 409 19975
rect 443 19941 459 19975
rect 393 19907 459 19941
rect 393 19873 409 19907
rect 443 19873 459 19907
rect 393 19839 459 19873
rect 393 19805 409 19839
rect 443 19805 459 19839
rect 393 19771 459 19805
rect 393 19737 409 19771
rect 443 19737 459 19771
rect 393 19720 459 19737
rect 489 19975 555 19992
rect 489 19941 505 19975
rect 539 19941 555 19975
rect 489 19907 555 19941
rect 489 19873 505 19907
rect 539 19873 555 19907
rect 489 19839 555 19873
rect 489 19805 505 19839
rect 539 19805 555 19839
rect 489 19771 555 19805
rect 489 19737 505 19771
rect 539 19737 555 19771
rect 489 19720 555 19737
rect 585 19975 651 19992
rect 585 19941 601 19975
rect 635 19941 651 19975
rect 585 19907 651 19941
rect 585 19873 601 19907
rect 635 19873 651 19907
rect 585 19839 651 19873
rect 585 19805 601 19839
rect 635 19805 651 19839
rect 585 19771 651 19805
rect 585 19737 601 19771
rect 635 19737 651 19771
rect 585 19720 651 19737
rect 681 19975 747 19992
rect 681 19941 697 19975
rect 731 19941 747 19975
rect 681 19907 747 19941
rect 681 19873 697 19907
rect 731 19873 747 19907
rect 681 19839 747 19873
rect 681 19805 697 19839
rect 731 19805 747 19839
rect 681 19771 747 19805
rect 681 19737 697 19771
rect 731 19737 747 19771
rect 681 19720 747 19737
rect 777 19975 843 19992
rect 777 19941 793 19975
rect 827 19941 843 19975
rect 777 19907 843 19941
rect 777 19873 793 19907
rect 827 19873 843 19907
rect 777 19839 843 19873
rect 777 19805 793 19839
rect 827 19805 843 19839
rect 777 19771 843 19805
rect 777 19737 793 19771
rect 827 19737 843 19771
rect 777 19720 843 19737
rect 873 19975 939 19992
rect 873 19941 889 19975
rect 923 19941 939 19975
rect 873 19907 939 19941
rect 873 19873 889 19907
rect 923 19873 939 19907
rect 873 19839 939 19873
rect 873 19805 889 19839
rect 923 19805 939 19839
rect 873 19771 939 19805
rect 873 19737 889 19771
rect 923 19737 939 19771
rect 873 19720 939 19737
rect 969 19975 1035 19992
rect 969 19941 985 19975
rect 1019 19941 1035 19975
rect 969 19907 1035 19941
rect 969 19873 985 19907
rect 1019 19873 1035 19907
rect 969 19839 1035 19873
rect 969 19805 985 19839
rect 1019 19805 1035 19839
rect 969 19771 1035 19805
rect 969 19737 985 19771
rect 1019 19737 1035 19771
rect 969 19720 1035 19737
rect 1065 19975 1131 19992
rect 1065 19941 1081 19975
rect 1115 19941 1131 19975
rect 1065 19907 1131 19941
rect 1065 19873 1081 19907
rect 1115 19873 1131 19907
rect 1065 19839 1131 19873
rect 1065 19805 1081 19839
rect 1115 19805 1131 19839
rect 1065 19771 1131 19805
rect 1065 19737 1081 19771
rect 1115 19737 1131 19771
rect 1065 19720 1131 19737
rect 1161 19975 1227 19992
rect 1161 19941 1177 19975
rect 1211 19941 1227 19975
rect 1161 19907 1227 19941
rect 1161 19873 1177 19907
rect 1211 19873 1227 19907
rect 1161 19839 1227 19873
rect 1161 19805 1177 19839
rect 1211 19805 1227 19839
rect 1161 19771 1227 19805
rect 1161 19737 1177 19771
rect 1211 19737 1227 19771
rect 1161 19720 1227 19737
rect 1257 19975 1319 19992
rect 1257 19941 1273 19975
rect 1307 19941 1319 19975
rect 1257 19907 1319 19941
rect 1257 19873 1273 19907
rect 1307 19873 1319 19907
rect 1257 19839 1319 19873
rect 1257 19805 1273 19839
rect 1307 19805 1319 19839
rect 1257 19771 1319 19805
rect 1257 19737 1273 19771
rect 1307 19737 1319 19771
rect 1257 19720 1319 19737
rect 2454 19979 2516 19996
rect 2454 19945 2466 19979
rect 2500 19945 2516 19979
rect 2454 19911 2516 19945
rect 2454 19877 2466 19911
rect 2500 19877 2516 19911
rect 2454 19843 2516 19877
rect 2454 19809 2466 19843
rect 2500 19809 2516 19843
rect 2454 19775 2516 19809
rect 2454 19741 2466 19775
rect 2500 19741 2516 19775
rect 2454 19724 2516 19741
rect 2546 19979 2612 19996
rect 2546 19945 2562 19979
rect 2596 19945 2612 19979
rect 2546 19911 2612 19945
rect 2546 19877 2562 19911
rect 2596 19877 2612 19911
rect 2546 19843 2612 19877
rect 2546 19809 2562 19843
rect 2596 19809 2612 19843
rect 2546 19775 2612 19809
rect 2546 19741 2562 19775
rect 2596 19741 2612 19775
rect 2546 19724 2612 19741
rect 2642 19979 2708 19996
rect 2642 19945 2658 19979
rect 2692 19945 2708 19979
rect 2642 19911 2708 19945
rect 2642 19877 2658 19911
rect 2692 19877 2708 19911
rect 2642 19843 2708 19877
rect 2642 19809 2658 19843
rect 2692 19809 2708 19843
rect 2642 19775 2708 19809
rect 2642 19741 2658 19775
rect 2692 19741 2708 19775
rect 2642 19724 2708 19741
rect 2738 19979 2804 19996
rect 2738 19945 2754 19979
rect 2788 19945 2804 19979
rect 2738 19911 2804 19945
rect 2738 19877 2754 19911
rect 2788 19877 2804 19911
rect 2738 19843 2804 19877
rect 2738 19809 2754 19843
rect 2788 19809 2804 19843
rect 2738 19775 2804 19809
rect 2738 19741 2754 19775
rect 2788 19741 2804 19775
rect 2738 19724 2804 19741
rect 2834 19979 2900 19996
rect 2834 19945 2850 19979
rect 2884 19945 2900 19979
rect 2834 19911 2900 19945
rect 2834 19877 2850 19911
rect 2884 19877 2900 19911
rect 2834 19843 2900 19877
rect 2834 19809 2850 19843
rect 2884 19809 2900 19843
rect 2834 19775 2900 19809
rect 2834 19741 2850 19775
rect 2884 19741 2900 19775
rect 2834 19724 2900 19741
rect 2930 19979 2996 19996
rect 2930 19945 2946 19979
rect 2980 19945 2996 19979
rect 2930 19911 2996 19945
rect 2930 19877 2946 19911
rect 2980 19877 2996 19911
rect 2930 19843 2996 19877
rect 2930 19809 2946 19843
rect 2980 19809 2996 19843
rect 2930 19775 2996 19809
rect 2930 19741 2946 19775
rect 2980 19741 2996 19775
rect 2930 19724 2996 19741
rect 3026 19979 3092 19996
rect 3026 19945 3042 19979
rect 3076 19945 3092 19979
rect 3026 19911 3092 19945
rect 3026 19877 3042 19911
rect 3076 19877 3092 19911
rect 3026 19843 3092 19877
rect 3026 19809 3042 19843
rect 3076 19809 3092 19843
rect 3026 19775 3092 19809
rect 3026 19741 3042 19775
rect 3076 19741 3092 19775
rect 3026 19724 3092 19741
rect 3122 19979 3188 19996
rect 3122 19945 3138 19979
rect 3172 19945 3188 19979
rect 3122 19911 3188 19945
rect 3122 19877 3138 19911
rect 3172 19877 3188 19911
rect 3122 19843 3188 19877
rect 3122 19809 3138 19843
rect 3172 19809 3188 19843
rect 3122 19775 3188 19809
rect 3122 19741 3138 19775
rect 3172 19741 3188 19775
rect 3122 19724 3188 19741
rect 3218 19979 3284 19996
rect 3218 19945 3234 19979
rect 3268 19945 3284 19979
rect 3218 19911 3284 19945
rect 3218 19877 3234 19911
rect 3268 19877 3284 19911
rect 3218 19843 3284 19877
rect 3218 19809 3234 19843
rect 3268 19809 3284 19843
rect 3218 19775 3284 19809
rect 3218 19741 3234 19775
rect 3268 19741 3284 19775
rect 3218 19724 3284 19741
rect 3314 19979 3380 19996
rect 3314 19945 3330 19979
rect 3364 19945 3380 19979
rect 3314 19911 3380 19945
rect 3314 19877 3330 19911
rect 3364 19877 3380 19911
rect 3314 19843 3380 19877
rect 3314 19809 3330 19843
rect 3364 19809 3380 19843
rect 3314 19775 3380 19809
rect 3314 19741 3330 19775
rect 3364 19741 3380 19775
rect 3314 19724 3380 19741
rect 3410 19979 3472 19996
rect 3410 19945 3426 19979
rect 3460 19945 3472 19979
rect 3410 19911 3472 19945
rect 3410 19877 3426 19911
rect 3460 19877 3472 19911
rect 3410 19843 3472 19877
rect 3410 19809 3426 19843
rect 3460 19809 3472 19843
rect 3410 19775 3472 19809
rect 3410 19741 3426 19775
rect 3460 19741 3472 19775
rect 3410 19724 3472 19741
rect 3975 19979 4037 19996
rect 3975 19945 3987 19979
rect 4021 19945 4037 19979
rect 3975 19911 4037 19945
rect 3975 19877 3987 19911
rect 4021 19877 4037 19911
rect 3975 19843 4037 19877
rect 3975 19809 3987 19843
rect 4021 19809 4037 19843
rect 3975 19775 4037 19809
rect 3975 19741 3987 19775
rect 4021 19741 4037 19775
rect 3975 19724 4037 19741
rect 4067 19979 4133 19996
rect 4067 19945 4083 19979
rect 4117 19945 4133 19979
rect 4067 19911 4133 19945
rect 4067 19877 4083 19911
rect 4117 19877 4133 19911
rect 4067 19843 4133 19877
rect 4067 19809 4083 19843
rect 4117 19809 4133 19843
rect 4067 19775 4133 19809
rect 4067 19741 4083 19775
rect 4117 19741 4133 19775
rect 4067 19724 4133 19741
rect 4163 19979 4229 19996
rect 4163 19945 4179 19979
rect 4213 19945 4229 19979
rect 4163 19911 4229 19945
rect 4163 19877 4179 19911
rect 4213 19877 4229 19911
rect 4163 19843 4229 19877
rect 4163 19809 4179 19843
rect 4213 19809 4229 19843
rect 4163 19775 4229 19809
rect 4163 19741 4179 19775
rect 4213 19741 4229 19775
rect 4163 19724 4229 19741
rect 4259 19979 4325 19996
rect 4259 19945 4275 19979
rect 4309 19945 4325 19979
rect 4259 19911 4325 19945
rect 4259 19877 4275 19911
rect 4309 19877 4325 19911
rect 4259 19843 4325 19877
rect 4259 19809 4275 19843
rect 4309 19809 4325 19843
rect 4259 19775 4325 19809
rect 4259 19741 4275 19775
rect 4309 19741 4325 19775
rect 4259 19724 4325 19741
rect 4355 19979 4421 19996
rect 4355 19945 4371 19979
rect 4405 19945 4421 19979
rect 4355 19911 4421 19945
rect 4355 19877 4371 19911
rect 4405 19877 4421 19911
rect 4355 19843 4421 19877
rect 4355 19809 4371 19843
rect 4405 19809 4421 19843
rect 4355 19775 4421 19809
rect 4355 19741 4371 19775
rect 4405 19741 4421 19775
rect 4355 19724 4421 19741
rect 4451 19979 4517 19996
rect 4451 19945 4467 19979
rect 4501 19945 4517 19979
rect 4451 19911 4517 19945
rect 4451 19877 4467 19911
rect 4501 19877 4517 19911
rect 4451 19843 4517 19877
rect 4451 19809 4467 19843
rect 4501 19809 4517 19843
rect 4451 19775 4517 19809
rect 4451 19741 4467 19775
rect 4501 19741 4517 19775
rect 4451 19724 4517 19741
rect 4547 19979 4613 19996
rect 4547 19945 4563 19979
rect 4597 19945 4613 19979
rect 4547 19911 4613 19945
rect 4547 19877 4563 19911
rect 4597 19877 4613 19911
rect 4547 19843 4613 19877
rect 4547 19809 4563 19843
rect 4597 19809 4613 19843
rect 4547 19775 4613 19809
rect 4547 19741 4563 19775
rect 4597 19741 4613 19775
rect 4547 19724 4613 19741
rect 4643 19979 4709 19996
rect 4643 19945 4659 19979
rect 4693 19945 4709 19979
rect 4643 19911 4709 19945
rect 4643 19877 4659 19911
rect 4693 19877 4709 19911
rect 4643 19843 4709 19877
rect 4643 19809 4659 19843
rect 4693 19809 4709 19843
rect 4643 19775 4709 19809
rect 4643 19741 4659 19775
rect 4693 19741 4709 19775
rect 4643 19724 4709 19741
rect 4739 19979 4805 19996
rect 4739 19945 4755 19979
rect 4789 19945 4805 19979
rect 4739 19911 4805 19945
rect 4739 19877 4755 19911
rect 4789 19877 4805 19911
rect 4739 19843 4805 19877
rect 4739 19809 4755 19843
rect 4789 19809 4805 19843
rect 4739 19775 4805 19809
rect 4739 19741 4755 19775
rect 4789 19741 4805 19775
rect 4739 19724 4805 19741
rect 4835 19979 4901 19996
rect 4835 19945 4851 19979
rect 4885 19945 4901 19979
rect 4835 19911 4901 19945
rect 4835 19877 4851 19911
rect 4885 19877 4901 19911
rect 4835 19843 4901 19877
rect 4835 19809 4851 19843
rect 4885 19809 4901 19843
rect 4835 19775 4901 19809
rect 4835 19741 4851 19775
rect 4885 19741 4901 19775
rect 4835 19724 4901 19741
rect 4931 19979 4993 19996
rect 4931 19945 4947 19979
rect 4981 19945 4993 19979
rect 4931 19911 4993 19945
rect 4931 19877 4947 19911
rect 4981 19877 4993 19911
rect 4931 19843 4993 19877
rect 4931 19809 4947 19843
rect 4981 19809 4993 19843
rect 4931 19775 4993 19809
rect 4931 19741 4947 19775
rect 4981 19741 4993 19775
rect 4931 19724 4993 19741
rect 5348 19771 5400 19783
rect 5348 19737 5356 19771
rect 5390 19737 5400 19771
rect 5348 19703 5400 19737
rect 5348 19669 5356 19703
rect 5390 19669 5400 19703
rect 5348 19635 5400 19669
rect 5348 19601 5356 19635
rect 5390 19601 5400 19635
rect 5348 19583 5400 19601
rect 5430 19771 5482 19783
rect 5430 19737 5440 19771
rect 5474 19737 5482 19771
rect 5430 19703 5482 19737
rect 5430 19669 5440 19703
rect 5474 19669 5482 19703
rect 5430 19635 5482 19669
rect 5430 19601 5440 19635
rect 5474 19601 5482 19635
rect 5430 19583 5482 19601
rect 301 18688 363 18705
rect 301 18654 313 18688
rect 347 18654 363 18688
rect 301 18620 363 18654
rect 301 18586 313 18620
rect 347 18586 363 18620
rect 301 18552 363 18586
rect 301 18518 313 18552
rect 347 18518 363 18552
rect 301 18484 363 18518
rect 301 18450 313 18484
rect 347 18450 363 18484
rect 301 18433 363 18450
rect 393 18688 459 18705
rect 393 18654 409 18688
rect 443 18654 459 18688
rect 393 18620 459 18654
rect 393 18586 409 18620
rect 443 18586 459 18620
rect 393 18552 459 18586
rect 393 18518 409 18552
rect 443 18518 459 18552
rect 393 18484 459 18518
rect 393 18450 409 18484
rect 443 18450 459 18484
rect 393 18433 459 18450
rect 489 18688 555 18705
rect 489 18654 505 18688
rect 539 18654 555 18688
rect 489 18620 555 18654
rect 489 18586 505 18620
rect 539 18586 555 18620
rect 489 18552 555 18586
rect 489 18518 505 18552
rect 539 18518 555 18552
rect 489 18484 555 18518
rect 489 18450 505 18484
rect 539 18450 555 18484
rect 489 18433 555 18450
rect 585 18688 651 18705
rect 585 18654 601 18688
rect 635 18654 651 18688
rect 585 18620 651 18654
rect 585 18586 601 18620
rect 635 18586 651 18620
rect 585 18552 651 18586
rect 585 18518 601 18552
rect 635 18518 651 18552
rect 585 18484 651 18518
rect 585 18450 601 18484
rect 635 18450 651 18484
rect 585 18433 651 18450
rect 681 18688 747 18705
rect 681 18654 697 18688
rect 731 18654 747 18688
rect 681 18620 747 18654
rect 681 18586 697 18620
rect 731 18586 747 18620
rect 681 18552 747 18586
rect 681 18518 697 18552
rect 731 18518 747 18552
rect 681 18484 747 18518
rect 681 18450 697 18484
rect 731 18450 747 18484
rect 681 18433 747 18450
rect 777 18688 843 18705
rect 777 18654 793 18688
rect 827 18654 843 18688
rect 777 18620 843 18654
rect 777 18586 793 18620
rect 827 18586 843 18620
rect 777 18552 843 18586
rect 777 18518 793 18552
rect 827 18518 843 18552
rect 777 18484 843 18518
rect 777 18450 793 18484
rect 827 18450 843 18484
rect 777 18433 843 18450
rect 873 18688 939 18705
rect 873 18654 889 18688
rect 923 18654 939 18688
rect 873 18620 939 18654
rect 873 18586 889 18620
rect 923 18586 939 18620
rect 873 18552 939 18586
rect 873 18518 889 18552
rect 923 18518 939 18552
rect 873 18484 939 18518
rect 873 18450 889 18484
rect 923 18450 939 18484
rect 873 18433 939 18450
rect 969 18688 1035 18705
rect 969 18654 985 18688
rect 1019 18654 1035 18688
rect 969 18620 1035 18654
rect 969 18586 985 18620
rect 1019 18586 1035 18620
rect 969 18552 1035 18586
rect 969 18518 985 18552
rect 1019 18518 1035 18552
rect 969 18484 1035 18518
rect 969 18450 985 18484
rect 1019 18450 1035 18484
rect 969 18433 1035 18450
rect 1065 18688 1131 18705
rect 1065 18654 1081 18688
rect 1115 18654 1131 18688
rect 1065 18620 1131 18654
rect 1065 18586 1081 18620
rect 1115 18586 1131 18620
rect 1065 18552 1131 18586
rect 1065 18518 1081 18552
rect 1115 18518 1131 18552
rect 1065 18484 1131 18518
rect 1065 18450 1081 18484
rect 1115 18450 1131 18484
rect 1065 18433 1131 18450
rect 1161 18688 1227 18705
rect 1161 18654 1177 18688
rect 1211 18654 1227 18688
rect 1161 18620 1227 18654
rect 1161 18586 1177 18620
rect 1211 18586 1227 18620
rect 1161 18552 1227 18586
rect 1161 18518 1177 18552
rect 1211 18518 1227 18552
rect 1161 18484 1227 18518
rect 1161 18450 1177 18484
rect 1211 18450 1227 18484
rect 1161 18433 1227 18450
rect 1257 18688 1319 18705
rect 1257 18654 1273 18688
rect 1307 18654 1319 18688
rect 1257 18620 1319 18654
rect 1257 18586 1273 18620
rect 1307 18586 1319 18620
rect 1257 18552 1319 18586
rect 1257 18518 1273 18552
rect 1307 18518 1319 18552
rect 1257 18484 1319 18518
rect 1257 18450 1273 18484
rect 1307 18450 1319 18484
rect 1257 18433 1319 18450
rect 2454 18692 2516 18709
rect 2454 18658 2466 18692
rect 2500 18658 2516 18692
rect 2454 18624 2516 18658
rect 2454 18590 2466 18624
rect 2500 18590 2516 18624
rect 2454 18556 2516 18590
rect 2454 18522 2466 18556
rect 2500 18522 2516 18556
rect 2454 18488 2516 18522
rect 2454 18454 2466 18488
rect 2500 18454 2516 18488
rect 2454 18437 2516 18454
rect 2546 18692 2612 18709
rect 2546 18658 2562 18692
rect 2596 18658 2612 18692
rect 2546 18624 2612 18658
rect 2546 18590 2562 18624
rect 2596 18590 2612 18624
rect 2546 18556 2612 18590
rect 2546 18522 2562 18556
rect 2596 18522 2612 18556
rect 2546 18488 2612 18522
rect 2546 18454 2562 18488
rect 2596 18454 2612 18488
rect 2546 18437 2612 18454
rect 2642 18692 2708 18709
rect 2642 18658 2658 18692
rect 2692 18658 2708 18692
rect 2642 18624 2708 18658
rect 2642 18590 2658 18624
rect 2692 18590 2708 18624
rect 2642 18556 2708 18590
rect 2642 18522 2658 18556
rect 2692 18522 2708 18556
rect 2642 18488 2708 18522
rect 2642 18454 2658 18488
rect 2692 18454 2708 18488
rect 2642 18437 2708 18454
rect 2738 18692 2804 18709
rect 2738 18658 2754 18692
rect 2788 18658 2804 18692
rect 2738 18624 2804 18658
rect 2738 18590 2754 18624
rect 2788 18590 2804 18624
rect 2738 18556 2804 18590
rect 2738 18522 2754 18556
rect 2788 18522 2804 18556
rect 2738 18488 2804 18522
rect 2738 18454 2754 18488
rect 2788 18454 2804 18488
rect 2738 18437 2804 18454
rect 2834 18692 2900 18709
rect 2834 18658 2850 18692
rect 2884 18658 2900 18692
rect 2834 18624 2900 18658
rect 2834 18590 2850 18624
rect 2884 18590 2900 18624
rect 2834 18556 2900 18590
rect 2834 18522 2850 18556
rect 2884 18522 2900 18556
rect 2834 18488 2900 18522
rect 2834 18454 2850 18488
rect 2884 18454 2900 18488
rect 2834 18437 2900 18454
rect 2930 18692 2996 18709
rect 2930 18658 2946 18692
rect 2980 18658 2996 18692
rect 2930 18624 2996 18658
rect 2930 18590 2946 18624
rect 2980 18590 2996 18624
rect 2930 18556 2996 18590
rect 2930 18522 2946 18556
rect 2980 18522 2996 18556
rect 2930 18488 2996 18522
rect 2930 18454 2946 18488
rect 2980 18454 2996 18488
rect 2930 18437 2996 18454
rect 3026 18692 3092 18709
rect 3026 18658 3042 18692
rect 3076 18658 3092 18692
rect 3026 18624 3092 18658
rect 3026 18590 3042 18624
rect 3076 18590 3092 18624
rect 3026 18556 3092 18590
rect 3026 18522 3042 18556
rect 3076 18522 3092 18556
rect 3026 18488 3092 18522
rect 3026 18454 3042 18488
rect 3076 18454 3092 18488
rect 3026 18437 3092 18454
rect 3122 18692 3188 18709
rect 3122 18658 3138 18692
rect 3172 18658 3188 18692
rect 3122 18624 3188 18658
rect 3122 18590 3138 18624
rect 3172 18590 3188 18624
rect 3122 18556 3188 18590
rect 3122 18522 3138 18556
rect 3172 18522 3188 18556
rect 3122 18488 3188 18522
rect 3122 18454 3138 18488
rect 3172 18454 3188 18488
rect 3122 18437 3188 18454
rect 3218 18692 3284 18709
rect 3218 18658 3234 18692
rect 3268 18658 3284 18692
rect 3218 18624 3284 18658
rect 3218 18590 3234 18624
rect 3268 18590 3284 18624
rect 3218 18556 3284 18590
rect 3218 18522 3234 18556
rect 3268 18522 3284 18556
rect 3218 18488 3284 18522
rect 3218 18454 3234 18488
rect 3268 18454 3284 18488
rect 3218 18437 3284 18454
rect 3314 18692 3380 18709
rect 3314 18658 3330 18692
rect 3364 18658 3380 18692
rect 3314 18624 3380 18658
rect 3314 18590 3330 18624
rect 3364 18590 3380 18624
rect 3314 18556 3380 18590
rect 3314 18522 3330 18556
rect 3364 18522 3380 18556
rect 3314 18488 3380 18522
rect 3314 18454 3330 18488
rect 3364 18454 3380 18488
rect 3314 18437 3380 18454
rect 3410 18692 3472 18709
rect 3410 18658 3426 18692
rect 3460 18658 3472 18692
rect 3410 18624 3472 18658
rect 3410 18590 3426 18624
rect 3460 18590 3472 18624
rect 3410 18556 3472 18590
rect 3410 18522 3426 18556
rect 3460 18522 3472 18556
rect 3410 18488 3472 18522
rect 3410 18454 3426 18488
rect 3460 18454 3472 18488
rect 3410 18437 3472 18454
rect 3975 18692 4037 18709
rect 3975 18658 3987 18692
rect 4021 18658 4037 18692
rect 3975 18624 4037 18658
rect 3975 18590 3987 18624
rect 4021 18590 4037 18624
rect 3975 18556 4037 18590
rect 3975 18522 3987 18556
rect 4021 18522 4037 18556
rect 3975 18488 4037 18522
rect 3975 18454 3987 18488
rect 4021 18454 4037 18488
rect 3975 18437 4037 18454
rect 4067 18692 4133 18709
rect 4067 18658 4083 18692
rect 4117 18658 4133 18692
rect 4067 18624 4133 18658
rect 4067 18590 4083 18624
rect 4117 18590 4133 18624
rect 4067 18556 4133 18590
rect 4067 18522 4083 18556
rect 4117 18522 4133 18556
rect 4067 18488 4133 18522
rect 4067 18454 4083 18488
rect 4117 18454 4133 18488
rect 4067 18437 4133 18454
rect 4163 18692 4229 18709
rect 4163 18658 4179 18692
rect 4213 18658 4229 18692
rect 4163 18624 4229 18658
rect 4163 18590 4179 18624
rect 4213 18590 4229 18624
rect 4163 18556 4229 18590
rect 4163 18522 4179 18556
rect 4213 18522 4229 18556
rect 4163 18488 4229 18522
rect 4163 18454 4179 18488
rect 4213 18454 4229 18488
rect 4163 18437 4229 18454
rect 4259 18692 4325 18709
rect 4259 18658 4275 18692
rect 4309 18658 4325 18692
rect 4259 18624 4325 18658
rect 4259 18590 4275 18624
rect 4309 18590 4325 18624
rect 4259 18556 4325 18590
rect 4259 18522 4275 18556
rect 4309 18522 4325 18556
rect 4259 18488 4325 18522
rect 4259 18454 4275 18488
rect 4309 18454 4325 18488
rect 4259 18437 4325 18454
rect 4355 18692 4421 18709
rect 4355 18658 4371 18692
rect 4405 18658 4421 18692
rect 4355 18624 4421 18658
rect 4355 18590 4371 18624
rect 4405 18590 4421 18624
rect 4355 18556 4421 18590
rect 4355 18522 4371 18556
rect 4405 18522 4421 18556
rect 4355 18488 4421 18522
rect 4355 18454 4371 18488
rect 4405 18454 4421 18488
rect 4355 18437 4421 18454
rect 4451 18692 4517 18709
rect 4451 18658 4467 18692
rect 4501 18658 4517 18692
rect 4451 18624 4517 18658
rect 4451 18590 4467 18624
rect 4501 18590 4517 18624
rect 4451 18556 4517 18590
rect 4451 18522 4467 18556
rect 4501 18522 4517 18556
rect 4451 18488 4517 18522
rect 4451 18454 4467 18488
rect 4501 18454 4517 18488
rect 4451 18437 4517 18454
rect 4547 18692 4613 18709
rect 4547 18658 4563 18692
rect 4597 18658 4613 18692
rect 4547 18624 4613 18658
rect 4547 18590 4563 18624
rect 4597 18590 4613 18624
rect 4547 18556 4613 18590
rect 4547 18522 4563 18556
rect 4597 18522 4613 18556
rect 4547 18488 4613 18522
rect 4547 18454 4563 18488
rect 4597 18454 4613 18488
rect 4547 18437 4613 18454
rect 4643 18692 4709 18709
rect 4643 18658 4659 18692
rect 4693 18658 4709 18692
rect 4643 18624 4709 18658
rect 4643 18590 4659 18624
rect 4693 18590 4709 18624
rect 4643 18556 4709 18590
rect 4643 18522 4659 18556
rect 4693 18522 4709 18556
rect 4643 18488 4709 18522
rect 4643 18454 4659 18488
rect 4693 18454 4709 18488
rect 4643 18437 4709 18454
rect 4739 18692 4805 18709
rect 4739 18658 4755 18692
rect 4789 18658 4805 18692
rect 4739 18624 4805 18658
rect 4739 18590 4755 18624
rect 4789 18590 4805 18624
rect 4739 18556 4805 18590
rect 4739 18522 4755 18556
rect 4789 18522 4805 18556
rect 4739 18488 4805 18522
rect 4739 18454 4755 18488
rect 4789 18454 4805 18488
rect 4739 18437 4805 18454
rect 4835 18692 4901 18709
rect 4835 18658 4851 18692
rect 4885 18658 4901 18692
rect 4835 18624 4901 18658
rect 4835 18590 4851 18624
rect 4885 18590 4901 18624
rect 4835 18556 4901 18590
rect 4835 18522 4851 18556
rect 4885 18522 4901 18556
rect 4835 18488 4901 18522
rect 4835 18454 4851 18488
rect 4885 18454 4901 18488
rect 4835 18437 4901 18454
rect 4931 18692 4993 18709
rect 4931 18658 4947 18692
rect 4981 18658 4993 18692
rect 4931 18624 4993 18658
rect 4931 18590 4947 18624
rect 4981 18590 4993 18624
rect 4931 18556 4993 18590
rect 4931 18522 4947 18556
rect 4981 18522 4993 18556
rect 4931 18488 4993 18522
rect 4931 18454 4947 18488
rect 4981 18454 4993 18488
rect 4931 18437 4993 18454
rect 5348 18484 5400 18496
rect 5348 18450 5356 18484
rect 5390 18450 5400 18484
rect 5348 18416 5400 18450
rect 5348 18382 5356 18416
rect 5390 18382 5400 18416
rect 5348 18348 5400 18382
rect 5348 18314 5356 18348
rect 5390 18314 5400 18348
rect 5348 18296 5400 18314
rect 5430 18484 5482 18496
rect 5430 18450 5440 18484
rect 5474 18450 5482 18484
rect 5430 18416 5482 18450
rect 5430 18382 5440 18416
rect 5474 18382 5482 18416
rect 5430 18348 5482 18382
rect 5430 18314 5440 18348
rect 5474 18314 5482 18348
rect 5430 18296 5482 18314
rect 301 17401 363 17418
rect 301 17367 313 17401
rect 347 17367 363 17401
rect 301 17333 363 17367
rect 301 17299 313 17333
rect 347 17299 363 17333
rect 301 17265 363 17299
rect 301 17231 313 17265
rect 347 17231 363 17265
rect 301 17197 363 17231
rect 301 17163 313 17197
rect 347 17163 363 17197
rect 301 17146 363 17163
rect 393 17401 459 17418
rect 393 17367 409 17401
rect 443 17367 459 17401
rect 393 17333 459 17367
rect 393 17299 409 17333
rect 443 17299 459 17333
rect 393 17265 459 17299
rect 393 17231 409 17265
rect 443 17231 459 17265
rect 393 17197 459 17231
rect 393 17163 409 17197
rect 443 17163 459 17197
rect 393 17146 459 17163
rect 489 17401 555 17418
rect 489 17367 505 17401
rect 539 17367 555 17401
rect 489 17333 555 17367
rect 489 17299 505 17333
rect 539 17299 555 17333
rect 489 17265 555 17299
rect 489 17231 505 17265
rect 539 17231 555 17265
rect 489 17197 555 17231
rect 489 17163 505 17197
rect 539 17163 555 17197
rect 489 17146 555 17163
rect 585 17401 651 17418
rect 585 17367 601 17401
rect 635 17367 651 17401
rect 585 17333 651 17367
rect 585 17299 601 17333
rect 635 17299 651 17333
rect 585 17265 651 17299
rect 585 17231 601 17265
rect 635 17231 651 17265
rect 585 17197 651 17231
rect 585 17163 601 17197
rect 635 17163 651 17197
rect 585 17146 651 17163
rect 681 17401 747 17418
rect 681 17367 697 17401
rect 731 17367 747 17401
rect 681 17333 747 17367
rect 681 17299 697 17333
rect 731 17299 747 17333
rect 681 17265 747 17299
rect 681 17231 697 17265
rect 731 17231 747 17265
rect 681 17197 747 17231
rect 681 17163 697 17197
rect 731 17163 747 17197
rect 681 17146 747 17163
rect 777 17401 843 17418
rect 777 17367 793 17401
rect 827 17367 843 17401
rect 777 17333 843 17367
rect 777 17299 793 17333
rect 827 17299 843 17333
rect 777 17265 843 17299
rect 777 17231 793 17265
rect 827 17231 843 17265
rect 777 17197 843 17231
rect 777 17163 793 17197
rect 827 17163 843 17197
rect 777 17146 843 17163
rect 873 17401 939 17418
rect 873 17367 889 17401
rect 923 17367 939 17401
rect 873 17333 939 17367
rect 873 17299 889 17333
rect 923 17299 939 17333
rect 873 17265 939 17299
rect 873 17231 889 17265
rect 923 17231 939 17265
rect 873 17197 939 17231
rect 873 17163 889 17197
rect 923 17163 939 17197
rect 873 17146 939 17163
rect 969 17401 1035 17418
rect 969 17367 985 17401
rect 1019 17367 1035 17401
rect 969 17333 1035 17367
rect 969 17299 985 17333
rect 1019 17299 1035 17333
rect 969 17265 1035 17299
rect 969 17231 985 17265
rect 1019 17231 1035 17265
rect 969 17197 1035 17231
rect 969 17163 985 17197
rect 1019 17163 1035 17197
rect 969 17146 1035 17163
rect 1065 17401 1131 17418
rect 1065 17367 1081 17401
rect 1115 17367 1131 17401
rect 1065 17333 1131 17367
rect 1065 17299 1081 17333
rect 1115 17299 1131 17333
rect 1065 17265 1131 17299
rect 1065 17231 1081 17265
rect 1115 17231 1131 17265
rect 1065 17197 1131 17231
rect 1065 17163 1081 17197
rect 1115 17163 1131 17197
rect 1065 17146 1131 17163
rect 1161 17401 1227 17418
rect 1161 17367 1177 17401
rect 1211 17367 1227 17401
rect 1161 17333 1227 17367
rect 1161 17299 1177 17333
rect 1211 17299 1227 17333
rect 1161 17265 1227 17299
rect 1161 17231 1177 17265
rect 1211 17231 1227 17265
rect 1161 17197 1227 17231
rect 1161 17163 1177 17197
rect 1211 17163 1227 17197
rect 1161 17146 1227 17163
rect 1257 17401 1319 17418
rect 1257 17367 1273 17401
rect 1307 17367 1319 17401
rect 1257 17333 1319 17367
rect 1257 17299 1273 17333
rect 1307 17299 1319 17333
rect 1257 17265 1319 17299
rect 1257 17231 1273 17265
rect 1307 17231 1319 17265
rect 1257 17197 1319 17231
rect 1257 17163 1273 17197
rect 1307 17163 1319 17197
rect 1257 17146 1319 17163
rect 2454 17405 2516 17422
rect 2454 17371 2466 17405
rect 2500 17371 2516 17405
rect 2454 17337 2516 17371
rect 2454 17303 2466 17337
rect 2500 17303 2516 17337
rect 2454 17269 2516 17303
rect 2454 17235 2466 17269
rect 2500 17235 2516 17269
rect 2454 17201 2516 17235
rect 2454 17167 2466 17201
rect 2500 17167 2516 17201
rect 2454 17150 2516 17167
rect 2546 17405 2612 17422
rect 2546 17371 2562 17405
rect 2596 17371 2612 17405
rect 2546 17337 2612 17371
rect 2546 17303 2562 17337
rect 2596 17303 2612 17337
rect 2546 17269 2612 17303
rect 2546 17235 2562 17269
rect 2596 17235 2612 17269
rect 2546 17201 2612 17235
rect 2546 17167 2562 17201
rect 2596 17167 2612 17201
rect 2546 17150 2612 17167
rect 2642 17405 2708 17422
rect 2642 17371 2658 17405
rect 2692 17371 2708 17405
rect 2642 17337 2708 17371
rect 2642 17303 2658 17337
rect 2692 17303 2708 17337
rect 2642 17269 2708 17303
rect 2642 17235 2658 17269
rect 2692 17235 2708 17269
rect 2642 17201 2708 17235
rect 2642 17167 2658 17201
rect 2692 17167 2708 17201
rect 2642 17150 2708 17167
rect 2738 17405 2804 17422
rect 2738 17371 2754 17405
rect 2788 17371 2804 17405
rect 2738 17337 2804 17371
rect 2738 17303 2754 17337
rect 2788 17303 2804 17337
rect 2738 17269 2804 17303
rect 2738 17235 2754 17269
rect 2788 17235 2804 17269
rect 2738 17201 2804 17235
rect 2738 17167 2754 17201
rect 2788 17167 2804 17201
rect 2738 17150 2804 17167
rect 2834 17405 2900 17422
rect 2834 17371 2850 17405
rect 2884 17371 2900 17405
rect 2834 17337 2900 17371
rect 2834 17303 2850 17337
rect 2884 17303 2900 17337
rect 2834 17269 2900 17303
rect 2834 17235 2850 17269
rect 2884 17235 2900 17269
rect 2834 17201 2900 17235
rect 2834 17167 2850 17201
rect 2884 17167 2900 17201
rect 2834 17150 2900 17167
rect 2930 17405 2996 17422
rect 2930 17371 2946 17405
rect 2980 17371 2996 17405
rect 2930 17337 2996 17371
rect 2930 17303 2946 17337
rect 2980 17303 2996 17337
rect 2930 17269 2996 17303
rect 2930 17235 2946 17269
rect 2980 17235 2996 17269
rect 2930 17201 2996 17235
rect 2930 17167 2946 17201
rect 2980 17167 2996 17201
rect 2930 17150 2996 17167
rect 3026 17405 3092 17422
rect 3026 17371 3042 17405
rect 3076 17371 3092 17405
rect 3026 17337 3092 17371
rect 3026 17303 3042 17337
rect 3076 17303 3092 17337
rect 3026 17269 3092 17303
rect 3026 17235 3042 17269
rect 3076 17235 3092 17269
rect 3026 17201 3092 17235
rect 3026 17167 3042 17201
rect 3076 17167 3092 17201
rect 3026 17150 3092 17167
rect 3122 17405 3188 17422
rect 3122 17371 3138 17405
rect 3172 17371 3188 17405
rect 3122 17337 3188 17371
rect 3122 17303 3138 17337
rect 3172 17303 3188 17337
rect 3122 17269 3188 17303
rect 3122 17235 3138 17269
rect 3172 17235 3188 17269
rect 3122 17201 3188 17235
rect 3122 17167 3138 17201
rect 3172 17167 3188 17201
rect 3122 17150 3188 17167
rect 3218 17405 3284 17422
rect 3218 17371 3234 17405
rect 3268 17371 3284 17405
rect 3218 17337 3284 17371
rect 3218 17303 3234 17337
rect 3268 17303 3284 17337
rect 3218 17269 3284 17303
rect 3218 17235 3234 17269
rect 3268 17235 3284 17269
rect 3218 17201 3284 17235
rect 3218 17167 3234 17201
rect 3268 17167 3284 17201
rect 3218 17150 3284 17167
rect 3314 17405 3380 17422
rect 3314 17371 3330 17405
rect 3364 17371 3380 17405
rect 3314 17337 3380 17371
rect 3314 17303 3330 17337
rect 3364 17303 3380 17337
rect 3314 17269 3380 17303
rect 3314 17235 3330 17269
rect 3364 17235 3380 17269
rect 3314 17201 3380 17235
rect 3314 17167 3330 17201
rect 3364 17167 3380 17201
rect 3314 17150 3380 17167
rect 3410 17405 3472 17422
rect 3410 17371 3426 17405
rect 3460 17371 3472 17405
rect 3410 17337 3472 17371
rect 3410 17303 3426 17337
rect 3460 17303 3472 17337
rect 3410 17269 3472 17303
rect 3410 17235 3426 17269
rect 3460 17235 3472 17269
rect 3410 17201 3472 17235
rect 3410 17167 3426 17201
rect 3460 17167 3472 17201
rect 3410 17150 3472 17167
rect 3975 17405 4037 17422
rect 3975 17371 3987 17405
rect 4021 17371 4037 17405
rect 3975 17337 4037 17371
rect 3975 17303 3987 17337
rect 4021 17303 4037 17337
rect 3975 17269 4037 17303
rect 3975 17235 3987 17269
rect 4021 17235 4037 17269
rect 3975 17201 4037 17235
rect 3975 17167 3987 17201
rect 4021 17167 4037 17201
rect 3975 17150 4037 17167
rect 4067 17405 4133 17422
rect 4067 17371 4083 17405
rect 4117 17371 4133 17405
rect 4067 17337 4133 17371
rect 4067 17303 4083 17337
rect 4117 17303 4133 17337
rect 4067 17269 4133 17303
rect 4067 17235 4083 17269
rect 4117 17235 4133 17269
rect 4067 17201 4133 17235
rect 4067 17167 4083 17201
rect 4117 17167 4133 17201
rect 4067 17150 4133 17167
rect 4163 17405 4229 17422
rect 4163 17371 4179 17405
rect 4213 17371 4229 17405
rect 4163 17337 4229 17371
rect 4163 17303 4179 17337
rect 4213 17303 4229 17337
rect 4163 17269 4229 17303
rect 4163 17235 4179 17269
rect 4213 17235 4229 17269
rect 4163 17201 4229 17235
rect 4163 17167 4179 17201
rect 4213 17167 4229 17201
rect 4163 17150 4229 17167
rect 4259 17405 4325 17422
rect 4259 17371 4275 17405
rect 4309 17371 4325 17405
rect 4259 17337 4325 17371
rect 4259 17303 4275 17337
rect 4309 17303 4325 17337
rect 4259 17269 4325 17303
rect 4259 17235 4275 17269
rect 4309 17235 4325 17269
rect 4259 17201 4325 17235
rect 4259 17167 4275 17201
rect 4309 17167 4325 17201
rect 4259 17150 4325 17167
rect 4355 17405 4421 17422
rect 4355 17371 4371 17405
rect 4405 17371 4421 17405
rect 4355 17337 4421 17371
rect 4355 17303 4371 17337
rect 4405 17303 4421 17337
rect 4355 17269 4421 17303
rect 4355 17235 4371 17269
rect 4405 17235 4421 17269
rect 4355 17201 4421 17235
rect 4355 17167 4371 17201
rect 4405 17167 4421 17201
rect 4355 17150 4421 17167
rect 4451 17405 4517 17422
rect 4451 17371 4467 17405
rect 4501 17371 4517 17405
rect 4451 17337 4517 17371
rect 4451 17303 4467 17337
rect 4501 17303 4517 17337
rect 4451 17269 4517 17303
rect 4451 17235 4467 17269
rect 4501 17235 4517 17269
rect 4451 17201 4517 17235
rect 4451 17167 4467 17201
rect 4501 17167 4517 17201
rect 4451 17150 4517 17167
rect 4547 17405 4613 17422
rect 4547 17371 4563 17405
rect 4597 17371 4613 17405
rect 4547 17337 4613 17371
rect 4547 17303 4563 17337
rect 4597 17303 4613 17337
rect 4547 17269 4613 17303
rect 4547 17235 4563 17269
rect 4597 17235 4613 17269
rect 4547 17201 4613 17235
rect 4547 17167 4563 17201
rect 4597 17167 4613 17201
rect 4547 17150 4613 17167
rect 4643 17405 4709 17422
rect 4643 17371 4659 17405
rect 4693 17371 4709 17405
rect 4643 17337 4709 17371
rect 4643 17303 4659 17337
rect 4693 17303 4709 17337
rect 4643 17269 4709 17303
rect 4643 17235 4659 17269
rect 4693 17235 4709 17269
rect 4643 17201 4709 17235
rect 4643 17167 4659 17201
rect 4693 17167 4709 17201
rect 4643 17150 4709 17167
rect 4739 17405 4805 17422
rect 4739 17371 4755 17405
rect 4789 17371 4805 17405
rect 4739 17337 4805 17371
rect 4739 17303 4755 17337
rect 4789 17303 4805 17337
rect 4739 17269 4805 17303
rect 4739 17235 4755 17269
rect 4789 17235 4805 17269
rect 4739 17201 4805 17235
rect 4739 17167 4755 17201
rect 4789 17167 4805 17201
rect 4739 17150 4805 17167
rect 4835 17405 4901 17422
rect 4835 17371 4851 17405
rect 4885 17371 4901 17405
rect 4835 17337 4901 17371
rect 4835 17303 4851 17337
rect 4885 17303 4901 17337
rect 4835 17269 4901 17303
rect 4835 17235 4851 17269
rect 4885 17235 4901 17269
rect 4835 17201 4901 17235
rect 4835 17167 4851 17201
rect 4885 17167 4901 17201
rect 4835 17150 4901 17167
rect 4931 17405 4993 17422
rect 4931 17371 4947 17405
rect 4981 17371 4993 17405
rect 4931 17337 4993 17371
rect 4931 17303 4947 17337
rect 4981 17303 4993 17337
rect 4931 17269 4993 17303
rect 4931 17235 4947 17269
rect 4981 17235 4993 17269
rect 4931 17201 4993 17235
rect 4931 17167 4947 17201
rect 4981 17167 4993 17201
rect 4931 17150 4993 17167
rect 5348 17197 5400 17209
rect 5348 17163 5356 17197
rect 5390 17163 5400 17197
rect 5348 17129 5400 17163
rect 5348 17095 5356 17129
rect 5390 17095 5400 17129
rect 5348 17061 5400 17095
rect 5348 17027 5356 17061
rect 5390 17027 5400 17061
rect 5348 17009 5400 17027
rect 5430 17197 5482 17209
rect 5430 17163 5440 17197
rect 5474 17163 5482 17197
rect 5430 17129 5482 17163
rect 5430 17095 5440 17129
rect 5474 17095 5482 17129
rect 5430 17061 5482 17095
rect 5430 17027 5440 17061
rect 5474 17027 5482 17061
rect 5430 17009 5482 17027
rect 301 16114 363 16131
rect 301 16080 313 16114
rect 347 16080 363 16114
rect 301 16046 363 16080
rect 301 16012 313 16046
rect 347 16012 363 16046
rect 301 15978 363 16012
rect 301 15944 313 15978
rect 347 15944 363 15978
rect 301 15910 363 15944
rect 301 15876 313 15910
rect 347 15876 363 15910
rect 301 15859 363 15876
rect 393 16114 459 16131
rect 393 16080 409 16114
rect 443 16080 459 16114
rect 393 16046 459 16080
rect 393 16012 409 16046
rect 443 16012 459 16046
rect 393 15978 459 16012
rect 393 15944 409 15978
rect 443 15944 459 15978
rect 393 15910 459 15944
rect 393 15876 409 15910
rect 443 15876 459 15910
rect 393 15859 459 15876
rect 489 16114 555 16131
rect 489 16080 505 16114
rect 539 16080 555 16114
rect 489 16046 555 16080
rect 489 16012 505 16046
rect 539 16012 555 16046
rect 489 15978 555 16012
rect 489 15944 505 15978
rect 539 15944 555 15978
rect 489 15910 555 15944
rect 489 15876 505 15910
rect 539 15876 555 15910
rect 489 15859 555 15876
rect 585 16114 651 16131
rect 585 16080 601 16114
rect 635 16080 651 16114
rect 585 16046 651 16080
rect 585 16012 601 16046
rect 635 16012 651 16046
rect 585 15978 651 16012
rect 585 15944 601 15978
rect 635 15944 651 15978
rect 585 15910 651 15944
rect 585 15876 601 15910
rect 635 15876 651 15910
rect 585 15859 651 15876
rect 681 16114 747 16131
rect 681 16080 697 16114
rect 731 16080 747 16114
rect 681 16046 747 16080
rect 681 16012 697 16046
rect 731 16012 747 16046
rect 681 15978 747 16012
rect 681 15944 697 15978
rect 731 15944 747 15978
rect 681 15910 747 15944
rect 681 15876 697 15910
rect 731 15876 747 15910
rect 681 15859 747 15876
rect 777 16114 843 16131
rect 777 16080 793 16114
rect 827 16080 843 16114
rect 777 16046 843 16080
rect 777 16012 793 16046
rect 827 16012 843 16046
rect 777 15978 843 16012
rect 777 15944 793 15978
rect 827 15944 843 15978
rect 777 15910 843 15944
rect 777 15876 793 15910
rect 827 15876 843 15910
rect 777 15859 843 15876
rect 873 16114 939 16131
rect 873 16080 889 16114
rect 923 16080 939 16114
rect 873 16046 939 16080
rect 873 16012 889 16046
rect 923 16012 939 16046
rect 873 15978 939 16012
rect 873 15944 889 15978
rect 923 15944 939 15978
rect 873 15910 939 15944
rect 873 15876 889 15910
rect 923 15876 939 15910
rect 873 15859 939 15876
rect 969 16114 1035 16131
rect 969 16080 985 16114
rect 1019 16080 1035 16114
rect 969 16046 1035 16080
rect 969 16012 985 16046
rect 1019 16012 1035 16046
rect 969 15978 1035 16012
rect 969 15944 985 15978
rect 1019 15944 1035 15978
rect 969 15910 1035 15944
rect 969 15876 985 15910
rect 1019 15876 1035 15910
rect 969 15859 1035 15876
rect 1065 16114 1131 16131
rect 1065 16080 1081 16114
rect 1115 16080 1131 16114
rect 1065 16046 1131 16080
rect 1065 16012 1081 16046
rect 1115 16012 1131 16046
rect 1065 15978 1131 16012
rect 1065 15944 1081 15978
rect 1115 15944 1131 15978
rect 1065 15910 1131 15944
rect 1065 15876 1081 15910
rect 1115 15876 1131 15910
rect 1065 15859 1131 15876
rect 1161 16114 1227 16131
rect 1161 16080 1177 16114
rect 1211 16080 1227 16114
rect 1161 16046 1227 16080
rect 1161 16012 1177 16046
rect 1211 16012 1227 16046
rect 1161 15978 1227 16012
rect 1161 15944 1177 15978
rect 1211 15944 1227 15978
rect 1161 15910 1227 15944
rect 1161 15876 1177 15910
rect 1211 15876 1227 15910
rect 1161 15859 1227 15876
rect 1257 16114 1319 16131
rect 1257 16080 1273 16114
rect 1307 16080 1319 16114
rect 1257 16046 1319 16080
rect 1257 16012 1273 16046
rect 1307 16012 1319 16046
rect 1257 15978 1319 16012
rect 1257 15944 1273 15978
rect 1307 15944 1319 15978
rect 1257 15910 1319 15944
rect 1257 15876 1273 15910
rect 1307 15876 1319 15910
rect 1257 15859 1319 15876
rect 2454 16118 2516 16135
rect 2454 16084 2466 16118
rect 2500 16084 2516 16118
rect 2454 16050 2516 16084
rect 2454 16016 2466 16050
rect 2500 16016 2516 16050
rect 2454 15982 2516 16016
rect 2454 15948 2466 15982
rect 2500 15948 2516 15982
rect 2454 15914 2516 15948
rect 2454 15880 2466 15914
rect 2500 15880 2516 15914
rect 2454 15863 2516 15880
rect 2546 16118 2612 16135
rect 2546 16084 2562 16118
rect 2596 16084 2612 16118
rect 2546 16050 2612 16084
rect 2546 16016 2562 16050
rect 2596 16016 2612 16050
rect 2546 15982 2612 16016
rect 2546 15948 2562 15982
rect 2596 15948 2612 15982
rect 2546 15914 2612 15948
rect 2546 15880 2562 15914
rect 2596 15880 2612 15914
rect 2546 15863 2612 15880
rect 2642 16118 2708 16135
rect 2642 16084 2658 16118
rect 2692 16084 2708 16118
rect 2642 16050 2708 16084
rect 2642 16016 2658 16050
rect 2692 16016 2708 16050
rect 2642 15982 2708 16016
rect 2642 15948 2658 15982
rect 2692 15948 2708 15982
rect 2642 15914 2708 15948
rect 2642 15880 2658 15914
rect 2692 15880 2708 15914
rect 2642 15863 2708 15880
rect 2738 16118 2804 16135
rect 2738 16084 2754 16118
rect 2788 16084 2804 16118
rect 2738 16050 2804 16084
rect 2738 16016 2754 16050
rect 2788 16016 2804 16050
rect 2738 15982 2804 16016
rect 2738 15948 2754 15982
rect 2788 15948 2804 15982
rect 2738 15914 2804 15948
rect 2738 15880 2754 15914
rect 2788 15880 2804 15914
rect 2738 15863 2804 15880
rect 2834 16118 2900 16135
rect 2834 16084 2850 16118
rect 2884 16084 2900 16118
rect 2834 16050 2900 16084
rect 2834 16016 2850 16050
rect 2884 16016 2900 16050
rect 2834 15982 2900 16016
rect 2834 15948 2850 15982
rect 2884 15948 2900 15982
rect 2834 15914 2900 15948
rect 2834 15880 2850 15914
rect 2884 15880 2900 15914
rect 2834 15863 2900 15880
rect 2930 16118 2996 16135
rect 2930 16084 2946 16118
rect 2980 16084 2996 16118
rect 2930 16050 2996 16084
rect 2930 16016 2946 16050
rect 2980 16016 2996 16050
rect 2930 15982 2996 16016
rect 2930 15948 2946 15982
rect 2980 15948 2996 15982
rect 2930 15914 2996 15948
rect 2930 15880 2946 15914
rect 2980 15880 2996 15914
rect 2930 15863 2996 15880
rect 3026 16118 3092 16135
rect 3026 16084 3042 16118
rect 3076 16084 3092 16118
rect 3026 16050 3092 16084
rect 3026 16016 3042 16050
rect 3076 16016 3092 16050
rect 3026 15982 3092 16016
rect 3026 15948 3042 15982
rect 3076 15948 3092 15982
rect 3026 15914 3092 15948
rect 3026 15880 3042 15914
rect 3076 15880 3092 15914
rect 3026 15863 3092 15880
rect 3122 16118 3188 16135
rect 3122 16084 3138 16118
rect 3172 16084 3188 16118
rect 3122 16050 3188 16084
rect 3122 16016 3138 16050
rect 3172 16016 3188 16050
rect 3122 15982 3188 16016
rect 3122 15948 3138 15982
rect 3172 15948 3188 15982
rect 3122 15914 3188 15948
rect 3122 15880 3138 15914
rect 3172 15880 3188 15914
rect 3122 15863 3188 15880
rect 3218 16118 3284 16135
rect 3218 16084 3234 16118
rect 3268 16084 3284 16118
rect 3218 16050 3284 16084
rect 3218 16016 3234 16050
rect 3268 16016 3284 16050
rect 3218 15982 3284 16016
rect 3218 15948 3234 15982
rect 3268 15948 3284 15982
rect 3218 15914 3284 15948
rect 3218 15880 3234 15914
rect 3268 15880 3284 15914
rect 3218 15863 3284 15880
rect 3314 16118 3380 16135
rect 3314 16084 3330 16118
rect 3364 16084 3380 16118
rect 3314 16050 3380 16084
rect 3314 16016 3330 16050
rect 3364 16016 3380 16050
rect 3314 15982 3380 16016
rect 3314 15948 3330 15982
rect 3364 15948 3380 15982
rect 3314 15914 3380 15948
rect 3314 15880 3330 15914
rect 3364 15880 3380 15914
rect 3314 15863 3380 15880
rect 3410 16118 3472 16135
rect 3410 16084 3426 16118
rect 3460 16084 3472 16118
rect 3410 16050 3472 16084
rect 3410 16016 3426 16050
rect 3460 16016 3472 16050
rect 3410 15982 3472 16016
rect 3410 15948 3426 15982
rect 3460 15948 3472 15982
rect 3410 15914 3472 15948
rect 3410 15880 3426 15914
rect 3460 15880 3472 15914
rect 3410 15863 3472 15880
rect 3975 16118 4037 16135
rect 3975 16084 3987 16118
rect 4021 16084 4037 16118
rect 3975 16050 4037 16084
rect 3975 16016 3987 16050
rect 4021 16016 4037 16050
rect 3975 15982 4037 16016
rect 3975 15948 3987 15982
rect 4021 15948 4037 15982
rect 3975 15914 4037 15948
rect 3975 15880 3987 15914
rect 4021 15880 4037 15914
rect 3975 15863 4037 15880
rect 4067 16118 4133 16135
rect 4067 16084 4083 16118
rect 4117 16084 4133 16118
rect 4067 16050 4133 16084
rect 4067 16016 4083 16050
rect 4117 16016 4133 16050
rect 4067 15982 4133 16016
rect 4067 15948 4083 15982
rect 4117 15948 4133 15982
rect 4067 15914 4133 15948
rect 4067 15880 4083 15914
rect 4117 15880 4133 15914
rect 4067 15863 4133 15880
rect 4163 16118 4229 16135
rect 4163 16084 4179 16118
rect 4213 16084 4229 16118
rect 4163 16050 4229 16084
rect 4163 16016 4179 16050
rect 4213 16016 4229 16050
rect 4163 15982 4229 16016
rect 4163 15948 4179 15982
rect 4213 15948 4229 15982
rect 4163 15914 4229 15948
rect 4163 15880 4179 15914
rect 4213 15880 4229 15914
rect 4163 15863 4229 15880
rect 4259 16118 4325 16135
rect 4259 16084 4275 16118
rect 4309 16084 4325 16118
rect 4259 16050 4325 16084
rect 4259 16016 4275 16050
rect 4309 16016 4325 16050
rect 4259 15982 4325 16016
rect 4259 15948 4275 15982
rect 4309 15948 4325 15982
rect 4259 15914 4325 15948
rect 4259 15880 4275 15914
rect 4309 15880 4325 15914
rect 4259 15863 4325 15880
rect 4355 16118 4421 16135
rect 4355 16084 4371 16118
rect 4405 16084 4421 16118
rect 4355 16050 4421 16084
rect 4355 16016 4371 16050
rect 4405 16016 4421 16050
rect 4355 15982 4421 16016
rect 4355 15948 4371 15982
rect 4405 15948 4421 15982
rect 4355 15914 4421 15948
rect 4355 15880 4371 15914
rect 4405 15880 4421 15914
rect 4355 15863 4421 15880
rect 4451 16118 4517 16135
rect 4451 16084 4467 16118
rect 4501 16084 4517 16118
rect 4451 16050 4517 16084
rect 4451 16016 4467 16050
rect 4501 16016 4517 16050
rect 4451 15982 4517 16016
rect 4451 15948 4467 15982
rect 4501 15948 4517 15982
rect 4451 15914 4517 15948
rect 4451 15880 4467 15914
rect 4501 15880 4517 15914
rect 4451 15863 4517 15880
rect 4547 16118 4613 16135
rect 4547 16084 4563 16118
rect 4597 16084 4613 16118
rect 4547 16050 4613 16084
rect 4547 16016 4563 16050
rect 4597 16016 4613 16050
rect 4547 15982 4613 16016
rect 4547 15948 4563 15982
rect 4597 15948 4613 15982
rect 4547 15914 4613 15948
rect 4547 15880 4563 15914
rect 4597 15880 4613 15914
rect 4547 15863 4613 15880
rect 4643 16118 4709 16135
rect 4643 16084 4659 16118
rect 4693 16084 4709 16118
rect 4643 16050 4709 16084
rect 4643 16016 4659 16050
rect 4693 16016 4709 16050
rect 4643 15982 4709 16016
rect 4643 15948 4659 15982
rect 4693 15948 4709 15982
rect 4643 15914 4709 15948
rect 4643 15880 4659 15914
rect 4693 15880 4709 15914
rect 4643 15863 4709 15880
rect 4739 16118 4805 16135
rect 4739 16084 4755 16118
rect 4789 16084 4805 16118
rect 4739 16050 4805 16084
rect 4739 16016 4755 16050
rect 4789 16016 4805 16050
rect 4739 15982 4805 16016
rect 4739 15948 4755 15982
rect 4789 15948 4805 15982
rect 4739 15914 4805 15948
rect 4739 15880 4755 15914
rect 4789 15880 4805 15914
rect 4739 15863 4805 15880
rect 4835 16118 4901 16135
rect 4835 16084 4851 16118
rect 4885 16084 4901 16118
rect 4835 16050 4901 16084
rect 4835 16016 4851 16050
rect 4885 16016 4901 16050
rect 4835 15982 4901 16016
rect 4835 15948 4851 15982
rect 4885 15948 4901 15982
rect 4835 15914 4901 15948
rect 4835 15880 4851 15914
rect 4885 15880 4901 15914
rect 4835 15863 4901 15880
rect 4931 16118 4993 16135
rect 4931 16084 4947 16118
rect 4981 16084 4993 16118
rect 4931 16050 4993 16084
rect 4931 16016 4947 16050
rect 4981 16016 4993 16050
rect 4931 15982 4993 16016
rect 4931 15948 4947 15982
rect 4981 15948 4993 15982
rect 4931 15914 4993 15948
rect 4931 15880 4947 15914
rect 4981 15880 4993 15914
rect 4931 15863 4993 15880
rect 5348 15910 5400 15922
rect 5348 15876 5356 15910
rect 5390 15876 5400 15910
rect 5348 15842 5400 15876
rect 5348 15808 5356 15842
rect 5390 15808 5400 15842
rect 5348 15774 5400 15808
rect 5348 15740 5356 15774
rect 5390 15740 5400 15774
rect 5348 15722 5400 15740
rect 5430 15910 5482 15922
rect 5430 15876 5440 15910
rect 5474 15876 5482 15910
rect 5430 15842 5482 15876
rect 5430 15808 5440 15842
rect 5474 15808 5482 15842
rect 5430 15774 5482 15808
rect 5430 15740 5440 15774
rect 5474 15740 5482 15774
rect 5430 15722 5482 15740
rect 301 14827 363 14844
rect 301 14793 313 14827
rect 347 14793 363 14827
rect 301 14759 363 14793
rect 301 14725 313 14759
rect 347 14725 363 14759
rect 301 14691 363 14725
rect 301 14657 313 14691
rect 347 14657 363 14691
rect 301 14623 363 14657
rect 301 14589 313 14623
rect 347 14589 363 14623
rect 301 14572 363 14589
rect 393 14827 459 14844
rect 393 14793 409 14827
rect 443 14793 459 14827
rect 393 14759 459 14793
rect 393 14725 409 14759
rect 443 14725 459 14759
rect 393 14691 459 14725
rect 393 14657 409 14691
rect 443 14657 459 14691
rect 393 14623 459 14657
rect 393 14589 409 14623
rect 443 14589 459 14623
rect 393 14572 459 14589
rect 489 14827 555 14844
rect 489 14793 505 14827
rect 539 14793 555 14827
rect 489 14759 555 14793
rect 489 14725 505 14759
rect 539 14725 555 14759
rect 489 14691 555 14725
rect 489 14657 505 14691
rect 539 14657 555 14691
rect 489 14623 555 14657
rect 489 14589 505 14623
rect 539 14589 555 14623
rect 489 14572 555 14589
rect 585 14827 651 14844
rect 585 14793 601 14827
rect 635 14793 651 14827
rect 585 14759 651 14793
rect 585 14725 601 14759
rect 635 14725 651 14759
rect 585 14691 651 14725
rect 585 14657 601 14691
rect 635 14657 651 14691
rect 585 14623 651 14657
rect 585 14589 601 14623
rect 635 14589 651 14623
rect 585 14572 651 14589
rect 681 14827 747 14844
rect 681 14793 697 14827
rect 731 14793 747 14827
rect 681 14759 747 14793
rect 681 14725 697 14759
rect 731 14725 747 14759
rect 681 14691 747 14725
rect 681 14657 697 14691
rect 731 14657 747 14691
rect 681 14623 747 14657
rect 681 14589 697 14623
rect 731 14589 747 14623
rect 681 14572 747 14589
rect 777 14827 843 14844
rect 777 14793 793 14827
rect 827 14793 843 14827
rect 777 14759 843 14793
rect 777 14725 793 14759
rect 827 14725 843 14759
rect 777 14691 843 14725
rect 777 14657 793 14691
rect 827 14657 843 14691
rect 777 14623 843 14657
rect 777 14589 793 14623
rect 827 14589 843 14623
rect 777 14572 843 14589
rect 873 14827 939 14844
rect 873 14793 889 14827
rect 923 14793 939 14827
rect 873 14759 939 14793
rect 873 14725 889 14759
rect 923 14725 939 14759
rect 873 14691 939 14725
rect 873 14657 889 14691
rect 923 14657 939 14691
rect 873 14623 939 14657
rect 873 14589 889 14623
rect 923 14589 939 14623
rect 873 14572 939 14589
rect 969 14827 1035 14844
rect 969 14793 985 14827
rect 1019 14793 1035 14827
rect 969 14759 1035 14793
rect 969 14725 985 14759
rect 1019 14725 1035 14759
rect 969 14691 1035 14725
rect 969 14657 985 14691
rect 1019 14657 1035 14691
rect 969 14623 1035 14657
rect 969 14589 985 14623
rect 1019 14589 1035 14623
rect 969 14572 1035 14589
rect 1065 14827 1131 14844
rect 1065 14793 1081 14827
rect 1115 14793 1131 14827
rect 1065 14759 1131 14793
rect 1065 14725 1081 14759
rect 1115 14725 1131 14759
rect 1065 14691 1131 14725
rect 1065 14657 1081 14691
rect 1115 14657 1131 14691
rect 1065 14623 1131 14657
rect 1065 14589 1081 14623
rect 1115 14589 1131 14623
rect 1065 14572 1131 14589
rect 1161 14827 1227 14844
rect 1161 14793 1177 14827
rect 1211 14793 1227 14827
rect 1161 14759 1227 14793
rect 1161 14725 1177 14759
rect 1211 14725 1227 14759
rect 1161 14691 1227 14725
rect 1161 14657 1177 14691
rect 1211 14657 1227 14691
rect 1161 14623 1227 14657
rect 1161 14589 1177 14623
rect 1211 14589 1227 14623
rect 1161 14572 1227 14589
rect 1257 14827 1319 14844
rect 1257 14793 1273 14827
rect 1307 14793 1319 14827
rect 1257 14759 1319 14793
rect 1257 14725 1273 14759
rect 1307 14725 1319 14759
rect 1257 14691 1319 14725
rect 1257 14657 1273 14691
rect 1307 14657 1319 14691
rect 1257 14623 1319 14657
rect 1257 14589 1273 14623
rect 1307 14589 1319 14623
rect 1257 14572 1319 14589
rect 2454 14831 2516 14848
rect 2454 14797 2466 14831
rect 2500 14797 2516 14831
rect 2454 14763 2516 14797
rect 2454 14729 2466 14763
rect 2500 14729 2516 14763
rect 2454 14695 2516 14729
rect 2454 14661 2466 14695
rect 2500 14661 2516 14695
rect 2454 14627 2516 14661
rect 2454 14593 2466 14627
rect 2500 14593 2516 14627
rect 2454 14576 2516 14593
rect 2546 14831 2612 14848
rect 2546 14797 2562 14831
rect 2596 14797 2612 14831
rect 2546 14763 2612 14797
rect 2546 14729 2562 14763
rect 2596 14729 2612 14763
rect 2546 14695 2612 14729
rect 2546 14661 2562 14695
rect 2596 14661 2612 14695
rect 2546 14627 2612 14661
rect 2546 14593 2562 14627
rect 2596 14593 2612 14627
rect 2546 14576 2612 14593
rect 2642 14831 2708 14848
rect 2642 14797 2658 14831
rect 2692 14797 2708 14831
rect 2642 14763 2708 14797
rect 2642 14729 2658 14763
rect 2692 14729 2708 14763
rect 2642 14695 2708 14729
rect 2642 14661 2658 14695
rect 2692 14661 2708 14695
rect 2642 14627 2708 14661
rect 2642 14593 2658 14627
rect 2692 14593 2708 14627
rect 2642 14576 2708 14593
rect 2738 14831 2804 14848
rect 2738 14797 2754 14831
rect 2788 14797 2804 14831
rect 2738 14763 2804 14797
rect 2738 14729 2754 14763
rect 2788 14729 2804 14763
rect 2738 14695 2804 14729
rect 2738 14661 2754 14695
rect 2788 14661 2804 14695
rect 2738 14627 2804 14661
rect 2738 14593 2754 14627
rect 2788 14593 2804 14627
rect 2738 14576 2804 14593
rect 2834 14831 2900 14848
rect 2834 14797 2850 14831
rect 2884 14797 2900 14831
rect 2834 14763 2900 14797
rect 2834 14729 2850 14763
rect 2884 14729 2900 14763
rect 2834 14695 2900 14729
rect 2834 14661 2850 14695
rect 2884 14661 2900 14695
rect 2834 14627 2900 14661
rect 2834 14593 2850 14627
rect 2884 14593 2900 14627
rect 2834 14576 2900 14593
rect 2930 14831 2996 14848
rect 2930 14797 2946 14831
rect 2980 14797 2996 14831
rect 2930 14763 2996 14797
rect 2930 14729 2946 14763
rect 2980 14729 2996 14763
rect 2930 14695 2996 14729
rect 2930 14661 2946 14695
rect 2980 14661 2996 14695
rect 2930 14627 2996 14661
rect 2930 14593 2946 14627
rect 2980 14593 2996 14627
rect 2930 14576 2996 14593
rect 3026 14831 3092 14848
rect 3026 14797 3042 14831
rect 3076 14797 3092 14831
rect 3026 14763 3092 14797
rect 3026 14729 3042 14763
rect 3076 14729 3092 14763
rect 3026 14695 3092 14729
rect 3026 14661 3042 14695
rect 3076 14661 3092 14695
rect 3026 14627 3092 14661
rect 3026 14593 3042 14627
rect 3076 14593 3092 14627
rect 3026 14576 3092 14593
rect 3122 14831 3188 14848
rect 3122 14797 3138 14831
rect 3172 14797 3188 14831
rect 3122 14763 3188 14797
rect 3122 14729 3138 14763
rect 3172 14729 3188 14763
rect 3122 14695 3188 14729
rect 3122 14661 3138 14695
rect 3172 14661 3188 14695
rect 3122 14627 3188 14661
rect 3122 14593 3138 14627
rect 3172 14593 3188 14627
rect 3122 14576 3188 14593
rect 3218 14831 3284 14848
rect 3218 14797 3234 14831
rect 3268 14797 3284 14831
rect 3218 14763 3284 14797
rect 3218 14729 3234 14763
rect 3268 14729 3284 14763
rect 3218 14695 3284 14729
rect 3218 14661 3234 14695
rect 3268 14661 3284 14695
rect 3218 14627 3284 14661
rect 3218 14593 3234 14627
rect 3268 14593 3284 14627
rect 3218 14576 3284 14593
rect 3314 14831 3380 14848
rect 3314 14797 3330 14831
rect 3364 14797 3380 14831
rect 3314 14763 3380 14797
rect 3314 14729 3330 14763
rect 3364 14729 3380 14763
rect 3314 14695 3380 14729
rect 3314 14661 3330 14695
rect 3364 14661 3380 14695
rect 3314 14627 3380 14661
rect 3314 14593 3330 14627
rect 3364 14593 3380 14627
rect 3314 14576 3380 14593
rect 3410 14831 3472 14848
rect 3410 14797 3426 14831
rect 3460 14797 3472 14831
rect 3410 14763 3472 14797
rect 3410 14729 3426 14763
rect 3460 14729 3472 14763
rect 3410 14695 3472 14729
rect 3410 14661 3426 14695
rect 3460 14661 3472 14695
rect 3410 14627 3472 14661
rect 3410 14593 3426 14627
rect 3460 14593 3472 14627
rect 3410 14576 3472 14593
rect 3975 14831 4037 14848
rect 3975 14797 3987 14831
rect 4021 14797 4037 14831
rect 3975 14763 4037 14797
rect 3975 14729 3987 14763
rect 4021 14729 4037 14763
rect 3975 14695 4037 14729
rect 3975 14661 3987 14695
rect 4021 14661 4037 14695
rect 3975 14627 4037 14661
rect 3975 14593 3987 14627
rect 4021 14593 4037 14627
rect 3975 14576 4037 14593
rect 4067 14831 4133 14848
rect 4067 14797 4083 14831
rect 4117 14797 4133 14831
rect 4067 14763 4133 14797
rect 4067 14729 4083 14763
rect 4117 14729 4133 14763
rect 4067 14695 4133 14729
rect 4067 14661 4083 14695
rect 4117 14661 4133 14695
rect 4067 14627 4133 14661
rect 4067 14593 4083 14627
rect 4117 14593 4133 14627
rect 4067 14576 4133 14593
rect 4163 14831 4229 14848
rect 4163 14797 4179 14831
rect 4213 14797 4229 14831
rect 4163 14763 4229 14797
rect 4163 14729 4179 14763
rect 4213 14729 4229 14763
rect 4163 14695 4229 14729
rect 4163 14661 4179 14695
rect 4213 14661 4229 14695
rect 4163 14627 4229 14661
rect 4163 14593 4179 14627
rect 4213 14593 4229 14627
rect 4163 14576 4229 14593
rect 4259 14831 4325 14848
rect 4259 14797 4275 14831
rect 4309 14797 4325 14831
rect 4259 14763 4325 14797
rect 4259 14729 4275 14763
rect 4309 14729 4325 14763
rect 4259 14695 4325 14729
rect 4259 14661 4275 14695
rect 4309 14661 4325 14695
rect 4259 14627 4325 14661
rect 4259 14593 4275 14627
rect 4309 14593 4325 14627
rect 4259 14576 4325 14593
rect 4355 14831 4421 14848
rect 4355 14797 4371 14831
rect 4405 14797 4421 14831
rect 4355 14763 4421 14797
rect 4355 14729 4371 14763
rect 4405 14729 4421 14763
rect 4355 14695 4421 14729
rect 4355 14661 4371 14695
rect 4405 14661 4421 14695
rect 4355 14627 4421 14661
rect 4355 14593 4371 14627
rect 4405 14593 4421 14627
rect 4355 14576 4421 14593
rect 4451 14831 4517 14848
rect 4451 14797 4467 14831
rect 4501 14797 4517 14831
rect 4451 14763 4517 14797
rect 4451 14729 4467 14763
rect 4501 14729 4517 14763
rect 4451 14695 4517 14729
rect 4451 14661 4467 14695
rect 4501 14661 4517 14695
rect 4451 14627 4517 14661
rect 4451 14593 4467 14627
rect 4501 14593 4517 14627
rect 4451 14576 4517 14593
rect 4547 14831 4613 14848
rect 4547 14797 4563 14831
rect 4597 14797 4613 14831
rect 4547 14763 4613 14797
rect 4547 14729 4563 14763
rect 4597 14729 4613 14763
rect 4547 14695 4613 14729
rect 4547 14661 4563 14695
rect 4597 14661 4613 14695
rect 4547 14627 4613 14661
rect 4547 14593 4563 14627
rect 4597 14593 4613 14627
rect 4547 14576 4613 14593
rect 4643 14831 4709 14848
rect 4643 14797 4659 14831
rect 4693 14797 4709 14831
rect 4643 14763 4709 14797
rect 4643 14729 4659 14763
rect 4693 14729 4709 14763
rect 4643 14695 4709 14729
rect 4643 14661 4659 14695
rect 4693 14661 4709 14695
rect 4643 14627 4709 14661
rect 4643 14593 4659 14627
rect 4693 14593 4709 14627
rect 4643 14576 4709 14593
rect 4739 14831 4805 14848
rect 4739 14797 4755 14831
rect 4789 14797 4805 14831
rect 4739 14763 4805 14797
rect 4739 14729 4755 14763
rect 4789 14729 4805 14763
rect 4739 14695 4805 14729
rect 4739 14661 4755 14695
rect 4789 14661 4805 14695
rect 4739 14627 4805 14661
rect 4739 14593 4755 14627
rect 4789 14593 4805 14627
rect 4739 14576 4805 14593
rect 4835 14831 4901 14848
rect 4835 14797 4851 14831
rect 4885 14797 4901 14831
rect 4835 14763 4901 14797
rect 4835 14729 4851 14763
rect 4885 14729 4901 14763
rect 4835 14695 4901 14729
rect 4835 14661 4851 14695
rect 4885 14661 4901 14695
rect 4835 14627 4901 14661
rect 4835 14593 4851 14627
rect 4885 14593 4901 14627
rect 4835 14576 4901 14593
rect 4931 14831 4993 14848
rect 4931 14797 4947 14831
rect 4981 14797 4993 14831
rect 4931 14763 4993 14797
rect 4931 14729 4947 14763
rect 4981 14729 4993 14763
rect 4931 14695 4993 14729
rect 4931 14661 4947 14695
rect 4981 14661 4993 14695
rect 4931 14627 4993 14661
rect 4931 14593 4947 14627
rect 4981 14593 4993 14627
rect 4931 14576 4993 14593
rect 5348 14623 5400 14635
rect 5348 14589 5356 14623
rect 5390 14589 5400 14623
rect 5348 14555 5400 14589
rect 5348 14521 5356 14555
rect 5390 14521 5400 14555
rect 5348 14487 5400 14521
rect 5348 14453 5356 14487
rect 5390 14453 5400 14487
rect 5348 14435 5400 14453
rect 5430 14623 5482 14635
rect 5430 14589 5440 14623
rect 5474 14589 5482 14623
rect 5430 14555 5482 14589
rect 5430 14521 5440 14555
rect 5474 14521 5482 14555
rect 5430 14487 5482 14521
rect 5430 14453 5440 14487
rect 5474 14453 5482 14487
rect 5430 14435 5482 14453
rect 301 13540 363 13557
rect 301 13506 313 13540
rect 347 13506 363 13540
rect 301 13472 363 13506
rect 301 13438 313 13472
rect 347 13438 363 13472
rect 301 13404 363 13438
rect 301 13370 313 13404
rect 347 13370 363 13404
rect 301 13336 363 13370
rect 301 13302 313 13336
rect 347 13302 363 13336
rect 301 13285 363 13302
rect 393 13540 459 13557
rect 393 13506 409 13540
rect 443 13506 459 13540
rect 393 13472 459 13506
rect 393 13438 409 13472
rect 443 13438 459 13472
rect 393 13404 459 13438
rect 393 13370 409 13404
rect 443 13370 459 13404
rect 393 13336 459 13370
rect 393 13302 409 13336
rect 443 13302 459 13336
rect 393 13285 459 13302
rect 489 13540 555 13557
rect 489 13506 505 13540
rect 539 13506 555 13540
rect 489 13472 555 13506
rect 489 13438 505 13472
rect 539 13438 555 13472
rect 489 13404 555 13438
rect 489 13370 505 13404
rect 539 13370 555 13404
rect 489 13336 555 13370
rect 489 13302 505 13336
rect 539 13302 555 13336
rect 489 13285 555 13302
rect 585 13540 651 13557
rect 585 13506 601 13540
rect 635 13506 651 13540
rect 585 13472 651 13506
rect 585 13438 601 13472
rect 635 13438 651 13472
rect 585 13404 651 13438
rect 585 13370 601 13404
rect 635 13370 651 13404
rect 585 13336 651 13370
rect 585 13302 601 13336
rect 635 13302 651 13336
rect 585 13285 651 13302
rect 681 13540 747 13557
rect 681 13506 697 13540
rect 731 13506 747 13540
rect 681 13472 747 13506
rect 681 13438 697 13472
rect 731 13438 747 13472
rect 681 13404 747 13438
rect 681 13370 697 13404
rect 731 13370 747 13404
rect 681 13336 747 13370
rect 681 13302 697 13336
rect 731 13302 747 13336
rect 681 13285 747 13302
rect 777 13540 843 13557
rect 777 13506 793 13540
rect 827 13506 843 13540
rect 777 13472 843 13506
rect 777 13438 793 13472
rect 827 13438 843 13472
rect 777 13404 843 13438
rect 777 13370 793 13404
rect 827 13370 843 13404
rect 777 13336 843 13370
rect 777 13302 793 13336
rect 827 13302 843 13336
rect 777 13285 843 13302
rect 873 13540 939 13557
rect 873 13506 889 13540
rect 923 13506 939 13540
rect 873 13472 939 13506
rect 873 13438 889 13472
rect 923 13438 939 13472
rect 873 13404 939 13438
rect 873 13370 889 13404
rect 923 13370 939 13404
rect 873 13336 939 13370
rect 873 13302 889 13336
rect 923 13302 939 13336
rect 873 13285 939 13302
rect 969 13540 1035 13557
rect 969 13506 985 13540
rect 1019 13506 1035 13540
rect 969 13472 1035 13506
rect 969 13438 985 13472
rect 1019 13438 1035 13472
rect 969 13404 1035 13438
rect 969 13370 985 13404
rect 1019 13370 1035 13404
rect 969 13336 1035 13370
rect 969 13302 985 13336
rect 1019 13302 1035 13336
rect 969 13285 1035 13302
rect 1065 13540 1131 13557
rect 1065 13506 1081 13540
rect 1115 13506 1131 13540
rect 1065 13472 1131 13506
rect 1065 13438 1081 13472
rect 1115 13438 1131 13472
rect 1065 13404 1131 13438
rect 1065 13370 1081 13404
rect 1115 13370 1131 13404
rect 1065 13336 1131 13370
rect 1065 13302 1081 13336
rect 1115 13302 1131 13336
rect 1065 13285 1131 13302
rect 1161 13540 1227 13557
rect 1161 13506 1177 13540
rect 1211 13506 1227 13540
rect 1161 13472 1227 13506
rect 1161 13438 1177 13472
rect 1211 13438 1227 13472
rect 1161 13404 1227 13438
rect 1161 13370 1177 13404
rect 1211 13370 1227 13404
rect 1161 13336 1227 13370
rect 1161 13302 1177 13336
rect 1211 13302 1227 13336
rect 1161 13285 1227 13302
rect 1257 13540 1319 13557
rect 1257 13506 1273 13540
rect 1307 13506 1319 13540
rect 1257 13472 1319 13506
rect 1257 13438 1273 13472
rect 1307 13438 1319 13472
rect 1257 13404 1319 13438
rect 1257 13370 1273 13404
rect 1307 13370 1319 13404
rect 1257 13336 1319 13370
rect 1257 13302 1273 13336
rect 1307 13302 1319 13336
rect 1257 13285 1319 13302
rect 2454 13544 2516 13561
rect 2454 13510 2466 13544
rect 2500 13510 2516 13544
rect 2454 13476 2516 13510
rect 2454 13442 2466 13476
rect 2500 13442 2516 13476
rect 2454 13408 2516 13442
rect 2454 13374 2466 13408
rect 2500 13374 2516 13408
rect 2454 13340 2516 13374
rect 2454 13306 2466 13340
rect 2500 13306 2516 13340
rect 2454 13289 2516 13306
rect 2546 13544 2612 13561
rect 2546 13510 2562 13544
rect 2596 13510 2612 13544
rect 2546 13476 2612 13510
rect 2546 13442 2562 13476
rect 2596 13442 2612 13476
rect 2546 13408 2612 13442
rect 2546 13374 2562 13408
rect 2596 13374 2612 13408
rect 2546 13340 2612 13374
rect 2546 13306 2562 13340
rect 2596 13306 2612 13340
rect 2546 13289 2612 13306
rect 2642 13544 2708 13561
rect 2642 13510 2658 13544
rect 2692 13510 2708 13544
rect 2642 13476 2708 13510
rect 2642 13442 2658 13476
rect 2692 13442 2708 13476
rect 2642 13408 2708 13442
rect 2642 13374 2658 13408
rect 2692 13374 2708 13408
rect 2642 13340 2708 13374
rect 2642 13306 2658 13340
rect 2692 13306 2708 13340
rect 2642 13289 2708 13306
rect 2738 13544 2804 13561
rect 2738 13510 2754 13544
rect 2788 13510 2804 13544
rect 2738 13476 2804 13510
rect 2738 13442 2754 13476
rect 2788 13442 2804 13476
rect 2738 13408 2804 13442
rect 2738 13374 2754 13408
rect 2788 13374 2804 13408
rect 2738 13340 2804 13374
rect 2738 13306 2754 13340
rect 2788 13306 2804 13340
rect 2738 13289 2804 13306
rect 2834 13544 2900 13561
rect 2834 13510 2850 13544
rect 2884 13510 2900 13544
rect 2834 13476 2900 13510
rect 2834 13442 2850 13476
rect 2884 13442 2900 13476
rect 2834 13408 2900 13442
rect 2834 13374 2850 13408
rect 2884 13374 2900 13408
rect 2834 13340 2900 13374
rect 2834 13306 2850 13340
rect 2884 13306 2900 13340
rect 2834 13289 2900 13306
rect 2930 13544 2996 13561
rect 2930 13510 2946 13544
rect 2980 13510 2996 13544
rect 2930 13476 2996 13510
rect 2930 13442 2946 13476
rect 2980 13442 2996 13476
rect 2930 13408 2996 13442
rect 2930 13374 2946 13408
rect 2980 13374 2996 13408
rect 2930 13340 2996 13374
rect 2930 13306 2946 13340
rect 2980 13306 2996 13340
rect 2930 13289 2996 13306
rect 3026 13544 3092 13561
rect 3026 13510 3042 13544
rect 3076 13510 3092 13544
rect 3026 13476 3092 13510
rect 3026 13442 3042 13476
rect 3076 13442 3092 13476
rect 3026 13408 3092 13442
rect 3026 13374 3042 13408
rect 3076 13374 3092 13408
rect 3026 13340 3092 13374
rect 3026 13306 3042 13340
rect 3076 13306 3092 13340
rect 3026 13289 3092 13306
rect 3122 13544 3188 13561
rect 3122 13510 3138 13544
rect 3172 13510 3188 13544
rect 3122 13476 3188 13510
rect 3122 13442 3138 13476
rect 3172 13442 3188 13476
rect 3122 13408 3188 13442
rect 3122 13374 3138 13408
rect 3172 13374 3188 13408
rect 3122 13340 3188 13374
rect 3122 13306 3138 13340
rect 3172 13306 3188 13340
rect 3122 13289 3188 13306
rect 3218 13544 3284 13561
rect 3218 13510 3234 13544
rect 3268 13510 3284 13544
rect 3218 13476 3284 13510
rect 3218 13442 3234 13476
rect 3268 13442 3284 13476
rect 3218 13408 3284 13442
rect 3218 13374 3234 13408
rect 3268 13374 3284 13408
rect 3218 13340 3284 13374
rect 3218 13306 3234 13340
rect 3268 13306 3284 13340
rect 3218 13289 3284 13306
rect 3314 13544 3380 13561
rect 3314 13510 3330 13544
rect 3364 13510 3380 13544
rect 3314 13476 3380 13510
rect 3314 13442 3330 13476
rect 3364 13442 3380 13476
rect 3314 13408 3380 13442
rect 3314 13374 3330 13408
rect 3364 13374 3380 13408
rect 3314 13340 3380 13374
rect 3314 13306 3330 13340
rect 3364 13306 3380 13340
rect 3314 13289 3380 13306
rect 3410 13544 3472 13561
rect 3410 13510 3426 13544
rect 3460 13510 3472 13544
rect 3410 13476 3472 13510
rect 3410 13442 3426 13476
rect 3460 13442 3472 13476
rect 3410 13408 3472 13442
rect 3410 13374 3426 13408
rect 3460 13374 3472 13408
rect 3410 13340 3472 13374
rect 3410 13306 3426 13340
rect 3460 13306 3472 13340
rect 3410 13289 3472 13306
rect 3975 13544 4037 13561
rect 3975 13510 3987 13544
rect 4021 13510 4037 13544
rect 3975 13476 4037 13510
rect 3975 13442 3987 13476
rect 4021 13442 4037 13476
rect 3975 13408 4037 13442
rect 3975 13374 3987 13408
rect 4021 13374 4037 13408
rect 3975 13340 4037 13374
rect 3975 13306 3987 13340
rect 4021 13306 4037 13340
rect 3975 13289 4037 13306
rect 4067 13544 4133 13561
rect 4067 13510 4083 13544
rect 4117 13510 4133 13544
rect 4067 13476 4133 13510
rect 4067 13442 4083 13476
rect 4117 13442 4133 13476
rect 4067 13408 4133 13442
rect 4067 13374 4083 13408
rect 4117 13374 4133 13408
rect 4067 13340 4133 13374
rect 4067 13306 4083 13340
rect 4117 13306 4133 13340
rect 4067 13289 4133 13306
rect 4163 13544 4229 13561
rect 4163 13510 4179 13544
rect 4213 13510 4229 13544
rect 4163 13476 4229 13510
rect 4163 13442 4179 13476
rect 4213 13442 4229 13476
rect 4163 13408 4229 13442
rect 4163 13374 4179 13408
rect 4213 13374 4229 13408
rect 4163 13340 4229 13374
rect 4163 13306 4179 13340
rect 4213 13306 4229 13340
rect 4163 13289 4229 13306
rect 4259 13544 4325 13561
rect 4259 13510 4275 13544
rect 4309 13510 4325 13544
rect 4259 13476 4325 13510
rect 4259 13442 4275 13476
rect 4309 13442 4325 13476
rect 4259 13408 4325 13442
rect 4259 13374 4275 13408
rect 4309 13374 4325 13408
rect 4259 13340 4325 13374
rect 4259 13306 4275 13340
rect 4309 13306 4325 13340
rect 4259 13289 4325 13306
rect 4355 13544 4421 13561
rect 4355 13510 4371 13544
rect 4405 13510 4421 13544
rect 4355 13476 4421 13510
rect 4355 13442 4371 13476
rect 4405 13442 4421 13476
rect 4355 13408 4421 13442
rect 4355 13374 4371 13408
rect 4405 13374 4421 13408
rect 4355 13340 4421 13374
rect 4355 13306 4371 13340
rect 4405 13306 4421 13340
rect 4355 13289 4421 13306
rect 4451 13544 4517 13561
rect 4451 13510 4467 13544
rect 4501 13510 4517 13544
rect 4451 13476 4517 13510
rect 4451 13442 4467 13476
rect 4501 13442 4517 13476
rect 4451 13408 4517 13442
rect 4451 13374 4467 13408
rect 4501 13374 4517 13408
rect 4451 13340 4517 13374
rect 4451 13306 4467 13340
rect 4501 13306 4517 13340
rect 4451 13289 4517 13306
rect 4547 13544 4613 13561
rect 4547 13510 4563 13544
rect 4597 13510 4613 13544
rect 4547 13476 4613 13510
rect 4547 13442 4563 13476
rect 4597 13442 4613 13476
rect 4547 13408 4613 13442
rect 4547 13374 4563 13408
rect 4597 13374 4613 13408
rect 4547 13340 4613 13374
rect 4547 13306 4563 13340
rect 4597 13306 4613 13340
rect 4547 13289 4613 13306
rect 4643 13544 4709 13561
rect 4643 13510 4659 13544
rect 4693 13510 4709 13544
rect 4643 13476 4709 13510
rect 4643 13442 4659 13476
rect 4693 13442 4709 13476
rect 4643 13408 4709 13442
rect 4643 13374 4659 13408
rect 4693 13374 4709 13408
rect 4643 13340 4709 13374
rect 4643 13306 4659 13340
rect 4693 13306 4709 13340
rect 4643 13289 4709 13306
rect 4739 13544 4805 13561
rect 4739 13510 4755 13544
rect 4789 13510 4805 13544
rect 4739 13476 4805 13510
rect 4739 13442 4755 13476
rect 4789 13442 4805 13476
rect 4739 13408 4805 13442
rect 4739 13374 4755 13408
rect 4789 13374 4805 13408
rect 4739 13340 4805 13374
rect 4739 13306 4755 13340
rect 4789 13306 4805 13340
rect 4739 13289 4805 13306
rect 4835 13544 4901 13561
rect 4835 13510 4851 13544
rect 4885 13510 4901 13544
rect 4835 13476 4901 13510
rect 4835 13442 4851 13476
rect 4885 13442 4901 13476
rect 4835 13408 4901 13442
rect 4835 13374 4851 13408
rect 4885 13374 4901 13408
rect 4835 13340 4901 13374
rect 4835 13306 4851 13340
rect 4885 13306 4901 13340
rect 4835 13289 4901 13306
rect 4931 13544 4993 13561
rect 4931 13510 4947 13544
rect 4981 13510 4993 13544
rect 4931 13476 4993 13510
rect 4931 13442 4947 13476
rect 4981 13442 4993 13476
rect 4931 13408 4993 13442
rect 4931 13374 4947 13408
rect 4981 13374 4993 13408
rect 4931 13340 4993 13374
rect 4931 13306 4947 13340
rect 4981 13306 4993 13340
rect 4931 13289 4993 13306
rect 5348 13336 5400 13348
rect 5348 13302 5356 13336
rect 5390 13302 5400 13336
rect 5348 13268 5400 13302
rect 5348 13234 5356 13268
rect 5390 13234 5400 13268
rect 5348 13200 5400 13234
rect 5348 13166 5356 13200
rect 5390 13166 5400 13200
rect 5348 13148 5400 13166
rect 5430 13336 5482 13348
rect 5430 13302 5440 13336
rect 5474 13302 5482 13336
rect 5430 13268 5482 13302
rect 5430 13234 5440 13268
rect 5474 13234 5482 13268
rect 5430 13200 5482 13234
rect 5430 13166 5440 13200
rect 5474 13166 5482 13200
rect 5430 13148 5482 13166
rect 301 12253 363 12270
rect 301 12219 313 12253
rect 347 12219 363 12253
rect 301 12185 363 12219
rect 301 12151 313 12185
rect 347 12151 363 12185
rect 301 12117 363 12151
rect 301 12083 313 12117
rect 347 12083 363 12117
rect 301 12049 363 12083
rect 301 12015 313 12049
rect 347 12015 363 12049
rect 301 11998 363 12015
rect 393 12253 459 12270
rect 393 12219 409 12253
rect 443 12219 459 12253
rect 393 12185 459 12219
rect 393 12151 409 12185
rect 443 12151 459 12185
rect 393 12117 459 12151
rect 393 12083 409 12117
rect 443 12083 459 12117
rect 393 12049 459 12083
rect 393 12015 409 12049
rect 443 12015 459 12049
rect 393 11998 459 12015
rect 489 12253 555 12270
rect 489 12219 505 12253
rect 539 12219 555 12253
rect 489 12185 555 12219
rect 489 12151 505 12185
rect 539 12151 555 12185
rect 489 12117 555 12151
rect 489 12083 505 12117
rect 539 12083 555 12117
rect 489 12049 555 12083
rect 489 12015 505 12049
rect 539 12015 555 12049
rect 489 11998 555 12015
rect 585 12253 651 12270
rect 585 12219 601 12253
rect 635 12219 651 12253
rect 585 12185 651 12219
rect 585 12151 601 12185
rect 635 12151 651 12185
rect 585 12117 651 12151
rect 585 12083 601 12117
rect 635 12083 651 12117
rect 585 12049 651 12083
rect 585 12015 601 12049
rect 635 12015 651 12049
rect 585 11998 651 12015
rect 681 12253 747 12270
rect 681 12219 697 12253
rect 731 12219 747 12253
rect 681 12185 747 12219
rect 681 12151 697 12185
rect 731 12151 747 12185
rect 681 12117 747 12151
rect 681 12083 697 12117
rect 731 12083 747 12117
rect 681 12049 747 12083
rect 681 12015 697 12049
rect 731 12015 747 12049
rect 681 11998 747 12015
rect 777 12253 843 12270
rect 777 12219 793 12253
rect 827 12219 843 12253
rect 777 12185 843 12219
rect 777 12151 793 12185
rect 827 12151 843 12185
rect 777 12117 843 12151
rect 777 12083 793 12117
rect 827 12083 843 12117
rect 777 12049 843 12083
rect 777 12015 793 12049
rect 827 12015 843 12049
rect 777 11998 843 12015
rect 873 12253 939 12270
rect 873 12219 889 12253
rect 923 12219 939 12253
rect 873 12185 939 12219
rect 873 12151 889 12185
rect 923 12151 939 12185
rect 873 12117 939 12151
rect 873 12083 889 12117
rect 923 12083 939 12117
rect 873 12049 939 12083
rect 873 12015 889 12049
rect 923 12015 939 12049
rect 873 11998 939 12015
rect 969 12253 1035 12270
rect 969 12219 985 12253
rect 1019 12219 1035 12253
rect 969 12185 1035 12219
rect 969 12151 985 12185
rect 1019 12151 1035 12185
rect 969 12117 1035 12151
rect 969 12083 985 12117
rect 1019 12083 1035 12117
rect 969 12049 1035 12083
rect 969 12015 985 12049
rect 1019 12015 1035 12049
rect 969 11998 1035 12015
rect 1065 12253 1131 12270
rect 1065 12219 1081 12253
rect 1115 12219 1131 12253
rect 1065 12185 1131 12219
rect 1065 12151 1081 12185
rect 1115 12151 1131 12185
rect 1065 12117 1131 12151
rect 1065 12083 1081 12117
rect 1115 12083 1131 12117
rect 1065 12049 1131 12083
rect 1065 12015 1081 12049
rect 1115 12015 1131 12049
rect 1065 11998 1131 12015
rect 1161 12253 1227 12270
rect 1161 12219 1177 12253
rect 1211 12219 1227 12253
rect 1161 12185 1227 12219
rect 1161 12151 1177 12185
rect 1211 12151 1227 12185
rect 1161 12117 1227 12151
rect 1161 12083 1177 12117
rect 1211 12083 1227 12117
rect 1161 12049 1227 12083
rect 1161 12015 1177 12049
rect 1211 12015 1227 12049
rect 1161 11998 1227 12015
rect 1257 12253 1319 12270
rect 1257 12219 1273 12253
rect 1307 12219 1319 12253
rect 1257 12185 1319 12219
rect 1257 12151 1273 12185
rect 1307 12151 1319 12185
rect 1257 12117 1319 12151
rect 1257 12083 1273 12117
rect 1307 12083 1319 12117
rect 1257 12049 1319 12083
rect 1257 12015 1273 12049
rect 1307 12015 1319 12049
rect 1257 11998 1319 12015
rect 2454 12257 2516 12274
rect 2454 12223 2466 12257
rect 2500 12223 2516 12257
rect 2454 12189 2516 12223
rect 2454 12155 2466 12189
rect 2500 12155 2516 12189
rect 2454 12121 2516 12155
rect 2454 12087 2466 12121
rect 2500 12087 2516 12121
rect 2454 12053 2516 12087
rect 2454 12019 2466 12053
rect 2500 12019 2516 12053
rect 2454 12002 2516 12019
rect 2546 12257 2612 12274
rect 2546 12223 2562 12257
rect 2596 12223 2612 12257
rect 2546 12189 2612 12223
rect 2546 12155 2562 12189
rect 2596 12155 2612 12189
rect 2546 12121 2612 12155
rect 2546 12087 2562 12121
rect 2596 12087 2612 12121
rect 2546 12053 2612 12087
rect 2546 12019 2562 12053
rect 2596 12019 2612 12053
rect 2546 12002 2612 12019
rect 2642 12257 2708 12274
rect 2642 12223 2658 12257
rect 2692 12223 2708 12257
rect 2642 12189 2708 12223
rect 2642 12155 2658 12189
rect 2692 12155 2708 12189
rect 2642 12121 2708 12155
rect 2642 12087 2658 12121
rect 2692 12087 2708 12121
rect 2642 12053 2708 12087
rect 2642 12019 2658 12053
rect 2692 12019 2708 12053
rect 2642 12002 2708 12019
rect 2738 12257 2804 12274
rect 2738 12223 2754 12257
rect 2788 12223 2804 12257
rect 2738 12189 2804 12223
rect 2738 12155 2754 12189
rect 2788 12155 2804 12189
rect 2738 12121 2804 12155
rect 2738 12087 2754 12121
rect 2788 12087 2804 12121
rect 2738 12053 2804 12087
rect 2738 12019 2754 12053
rect 2788 12019 2804 12053
rect 2738 12002 2804 12019
rect 2834 12257 2900 12274
rect 2834 12223 2850 12257
rect 2884 12223 2900 12257
rect 2834 12189 2900 12223
rect 2834 12155 2850 12189
rect 2884 12155 2900 12189
rect 2834 12121 2900 12155
rect 2834 12087 2850 12121
rect 2884 12087 2900 12121
rect 2834 12053 2900 12087
rect 2834 12019 2850 12053
rect 2884 12019 2900 12053
rect 2834 12002 2900 12019
rect 2930 12257 2996 12274
rect 2930 12223 2946 12257
rect 2980 12223 2996 12257
rect 2930 12189 2996 12223
rect 2930 12155 2946 12189
rect 2980 12155 2996 12189
rect 2930 12121 2996 12155
rect 2930 12087 2946 12121
rect 2980 12087 2996 12121
rect 2930 12053 2996 12087
rect 2930 12019 2946 12053
rect 2980 12019 2996 12053
rect 2930 12002 2996 12019
rect 3026 12257 3092 12274
rect 3026 12223 3042 12257
rect 3076 12223 3092 12257
rect 3026 12189 3092 12223
rect 3026 12155 3042 12189
rect 3076 12155 3092 12189
rect 3026 12121 3092 12155
rect 3026 12087 3042 12121
rect 3076 12087 3092 12121
rect 3026 12053 3092 12087
rect 3026 12019 3042 12053
rect 3076 12019 3092 12053
rect 3026 12002 3092 12019
rect 3122 12257 3188 12274
rect 3122 12223 3138 12257
rect 3172 12223 3188 12257
rect 3122 12189 3188 12223
rect 3122 12155 3138 12189
rect 3172 12155 3188 12189
rect 3122 12121 3188 12155
rect 3122 12087 3138 12121
rect 3172 12087 3188 12121
rect 3122 12053 3188 12087
rect 3122 12019 3138 12053
rect 3172 12019 3188 12053
rect 3122 12002 3188 12019
rect 3218 12257 3284 12274
rect 3218 12223 3234 12257
rect 3268 12223 3284 12257
rect 3218 12189 3284 12223
rect 3218 12155 3234 12189
rect 3268 12155 3284 12189
rect 3218 12121 3284 12155
rect 3218 12087 3234 12121
rect 3268 12087 3284 12121
rect 3218 12053 3284 12087
rect 3218 12019 3234 12053
rect 3268 12019 3284 12053
rect 3218 12002 3284 12019
rect 3314 12257 3380 12274
rect 3314 12223 3330 12257
rect 3364 12223 3380 12257
rect 3314 12189 3380 12223
rect 3314 12155 3330 12189
rect 3364 12155 3380 12189
rect 3314 12121 3380 12155
rect 3314 12087 3330 12121
rect 3364 12087 3380 12121
rect 3314 12053 3380 12087
rect 3314 12019 3330 12053
rect 3364 12019 3380 12053
rect 3314 12002 3380 12019
rect 3410 12257 3472 12274
rect 3410 12223 3426 12257
rect 3460 12223 3472 12257
rect 3410 12189 3472 12223
rect 3410 12155 3426 12189
rect 3460 12155 3472 12189
rect 3410 12121 3472 12155
rect 3410 12087 3426 12121
rect 3460 12087 3472 12121
rect 3410 12053 3472 12087
rect 3410 12019 3426 12053
rect 3460 12019 3472 12053
rect 3410 12002 3472 12019
rect 3975 12257 4037 12274
rect 3975 12223 3987 12257
rect 4021 12223 4037 12257
rect 3975 12189 4037 12223
rect 3975 12155 3987 12189
rect 4021 12155 4037 12189
rect 3975 12121 4037 12155
rect 3975 12087 3987 12121
rect 4021 12087 4037 12121
rect 3975 12053 4037 12087
rect 3975 12019 3987 12053
rect 4021 12019 4037 12053
rect 3975 12002 4037 12019
rect 4067 12257 4133 12274
rect 4067 12223 4083 12257
rect 4117 12223 4133 12257
rect 4067 12189 4133 12223
rect 4067 12155 4083 12189
rect 4117 12155 4133 12189
rect 4067 12121 4133 12155
rect 4067 12087 4083 12121
rect 4117 12087 4133 12121
rect 4067 12053 4133 12087
rect 4067 12019 4083 12053
rect 4117 12019 4133 12053
rect 4067 12002 4133 12019
rect 4163 12257 4229 12274
rect 4163 12223 4179 12257
rect 4213 12223 4229 12257
rect 4163 12189 4229 12223
rect 4163 12155 4179 12189
rect 4213 12155 4229 12189
rect 4163 12121 4229 12155
rect 4163 12087 4179 12121
rect 4213 12087 4229 12121
rect 4163 12053 4229 12087
rect 4163 12019 4179 12053
rect 4213 12019 4229 12053
rect 4163 12002 4229 12019
rect 4259 12257 4325 12274
rect 4259 12223 4275 12257
rect 4309 12223 4325 12257
rect 4259 12189 4325 12223
rect 4259 12155 4275 12189
rect 4309 12155 4325 12189
rect 4259 12121 4325 12155
rect 4259 12087 4275 12121
rect 4309 12087 4325 12121
rect 4259 12053 4325 12087
rect 4259 12019 4275 12053
rect 4309 12019 4325 12053
rect 4259 12002 4325 12019
rect 4355 12257 4421 12274
rect 4355 12223 4371 12257
rect 4405 12223 4421 12257
rect 4355 12189 4421 12223
rect 4355 12155 4371 12189
rect 4405 12155 4421 12189
rect 4355 12121 4421 12155
rect 4355 12087 4371 12121
rect 4405 12087 4421 12121
rect 4355 12053 4421 12087
rect 4355 12019 4371 12053
rect 4405 12019 4421 12053
rect 4355 12002 4421 12019
rect 4451 12257 4517 12274
rect 4451 12223 4467 12257
rect 4501 12223 4517 12257
rect 4451 12189 4517 12223
rect 4451 12155 4467 12189
rect 4501 12155 4517 12189
rect 4451 12121 4517 12155
rect 4451 12087 4467 12121
rect 4501 12087 4517 12121
rect 4451 12053 4517 12087
rect 4451 12019 4467 12053
rect 4501 12019 4517 12053
rect 4451 12002 4517 12019
rect 4547 12257 4613 12274
rect 4547 12223 4563 12257
rect 4597 12223 4613 12257
rect 4547 12189 4613 12223
rect 4547 12155 4563 12189
rect 4597 12155 4613 12189
rect 4547 12121 4613 12155
rect 4547 12087 4563 12121
rect 4597 12087 4613 12121
rect 4547 12053 4613 12087
rect 4547 12019 4563 12053
rect 4597 12019 4613 12053
rect 4547 12002 4613 12019
rect 4643 12257 4709 12274
rect 4643 12223 4659 12257
rect 4693 12223 4709 12257
rect 4643 12189 4709 12223
rect 4643 12155 4659 12189
rect 4693 12155 4709 12189
rect 4643 12121 4709 12155
rect 4643 12087 4659 12121
rect 4693 12087 4709 12121
rect 4643 12053 4709 12087
rect 4643 12019 4659 12053
rect 4693 12019 4709 12053
rect 4643 12002 4709 12019
rect 4739 12257 4805 12274
rect 4739 12223 4755 12257
rect 4789 12223 4805 12257
rect 4739 12189 4805 12223
rect 4739 12155 4755 12189
rect 4789 12155 4805 12189
rect 4739 12121 4805 12155
rect 4739 12087 4755 12121
rect 4789 12087 4805 12121
rect 4739 12053 4805 12087
rect 4739 12019 4755 12053
rect 4789 12019 4805 12053
rect 4739 12002 4805 12019
rect 4835 12257 4901 12274
rect 4835 12223 4851 12257
rect 4885 12223 4901 12257
rect 4835 12189 4901 12223
rect 4835 12155 4851 12189
rect 4885 12155 4901 12189
rect 4835 12121 4901 12155
rect 4835 12087 4851 12121
rect 4885 12087 4901 12121
rect 4835 12053 4901 12087
rect 4835 12019 4851 12053
rect 4885 12019 4901 12053
rect 4835 12002 4901 12019
rect 4931 12257 4993 12274
rect 4931 12223 4947 12257
rect 4981 12223 4993 12257
rect 4931 12189 4993 12223
rect 4931 12155 4947 12189
rect 4981 12155 4993 12189
rect 4931 12121 4993 12155
rect 4931 12087 4947 12121
rect 4981 12087 4993 12121
rect 4931 12053 4993 12087
rect 4931 12019 4947 12053
rect 4981 12019 4993 12053
rect 4931 12002 4993 12019
rect 5348 12049 5400 12061
rect 5348 12015 5356 12049
rect 5390 12015 5400 12049
rect 5348 11981 5400 12015
rect 5348 11947 5356 11981
rect 5390 11947 5400 11981
rect 5348 11913 5400 11947
rect 5348 11879 5356 11913
rect 5390 11879 5400 11913
rect 5348 11861 5400 11879
rect 5430 12049 5482 12061
rect 5430 12015 5440 12049
rect 5474 12015 5482 12049
rect 5430 11981 5482 12015
rect 5430 11947 5440 11981
rect 5474 11947 5482 11981
rect 5430 11913 5482 11947
rect 5430 11879 5440 11913
rect 5474 11879 5482 11913
rect 5430 11861 5482 11879
rect 301 10966 363 10983
rect 301 10932 313 10966
rect 347 10932 363 10966
rect 301 10898 363 10932
rect 301 10864 313 10898
rect 347 10864 363 10898
rect 301 10830 363 10864
rect 301 10796 313 10830
rect 347 10796 363 10830
rect 301 10762 363 10796
rect 301 10728 313 10762
rect 347 10728 363 10762
rect 301 10711 363 10728
rect 393 10966 459 10983
rect 393 10932 409 10966
rect 443 10932 459 10966
rect 393 10898 459 10932
rect 393 10864 409 10898
rect 443 10864 459 10898
rect 393 10830 459 10864
rect 393 10796 409 10830
rect 443 10796 459 10830
rect 393 10762 459 10796
rect 393 10728 409 10762
rect 443 10728 459 10762
rect 393 10711 459 10728
rect 489 10966 555 10983
rect 489 10932 505 10966
rect 539 10932 555 10966
rect 489 10898 555 10932
rect 489 10864 505 10898
rect 539 10864 555 10898
rect 489 10830 555 10864
rect 489 10796 505 10830
rect 539 10796 555 10830
rect 489 10762 555 10796
rect 489 10728 505 10762
rect 539 10728 555 10762
rect 489 10711 555 10728
rect 585 10966 651 10983
rect 585 10932 601 10966
rect 635 10932 651 10966
rect 585 10898 651 10932
rect 585 10864 601 10898
rect 635 10864 651 10898
rect 585 10830 651 10864
rect 585 10796 601 10830
rect 635 10796 651 10830
rect 585 10762 651 10796
rect 585 10728 601 10762
rect 635 10728 651 10762
rect 585 10711 651 10728
rect 681 10966 747 10983
rect 681 10932 697 10966
rect 731 10932 747 10966
rect 681 10898 747 10932
rect 681 10864 697 10898
rect 731 10864 747 10898
rect 681 10830 747 10864
rect 681 10796 697 10830
rect 731 10796 747 10830
rect 681 10762 747 10796
rect 681 10728 697 10762
rect 731 10728 747 10762
rect 681 10711 747 10728
rect 777 10966 843 10983
rect 777 10932 793 10966
rect 827 10932 843 10966
rect 777 10898 843 10932
rect 777 10864 793 10898
rect 827 10864 843 10898
rect 777 10830 843 10864
rect 777 10796 793 10830
rect 827 10796 843 10830
rect 777 10762 843 10796
rect 777 10728 793 10762
rect 827 10728 843 10762
rect 777 10711 843 10728
rect 873 10966 939 10983
rect 873 10932 889 10966
rect 923 10932 939 10966
rect 873 10898 939 10932
rect 873 10864 889 10898
rect 923 10864 939 10898
rect 873 10830 939 10864
rect 873 10796 889 10830
rect 923 10796 939 10830
rect 873 10762 939 10796
rect 873 10728 889 10762
rect 923 10728 939 10762
rect 873 10711 939 10728
rect 969 10966 1035 10983
rect 969 10932 985 10966
rect 1019 10932 1035 10966
rect 969 10898 1035 10932
rect 969 10864 985 10898
rect 1019 10864 1035 10898
rect 969 10830 1035 10864
rect 969 10796 985 10830
rect 1019 10796 1035 10830
rect 969 10762 1035 10796
rect 969 10728 985 10762
rect 1019 10728 1035 10762
rect 969 10711 1035 10728
rect 1065 10966 1131 10983
rect 1065 10932 1081 10966
rect 1115 10932 1131 10966
rect 1065 10898 1131 10932
rect 1065 10864 1081 10898
rect 1115 10864 1131 10898
rect 1065 10830 1131 10864
rect 1065 10796 1081 10830
rect 1115 10796 1131 10830
rect 1065 10762 1131 10796
rect 1065 10728 1081 10762
rect 1115 10728 1131 10762
rect 1065 10711 1131 10728
rect 1161 10966 1227 10983
rect 1161 10932 1177 10966
rect 1211 10932 1227 10966
rect 1161 10898 1227 10932
rect 1161 10864 1177 10898
rect 1211 10864 1227 10898
rect 1161 10830 1227 10864
rect 1161 10796 1177 10830
rect 1211 10796 1227 10830
rect 1161 10762 1227 10796
rect 1161 10728 1177 10762
rect 1211 10728 1227 10762
rect 1161 10711 1227 10728
rect 1257 10966 1319 10983
rect 1257 10932 1273 10966
rect 1307 10932 1319 10966
rect 1257 10898 1319 10932
rect 1257 10864 1273 10898
rect 1307 10864 1319 10898
rect 1257 10830 1319 10864
rect 1257 10796 1273 10830
rect 1307 10796 1319 10830
rect 1257 10762 1319 10796
rect 1257 10728 1273 10762
rect 1307 10728 1319 10762
rect 1257 10711 1319 10728
rect 2454 10970 2516 10987
rect 2454 10936 2466 10970
rect 2500 10936 2516 10970
rect 2454 10902 2516 10936
rect 2454 10868 2466 10902
rect 2500 10868 2516 10902
rect 2454 10834 2516 10868
rect 2454 10800 2466 10834
rect 2500 10800 2516 10834
rect 2454 10766 2516 10800
rect 2454 10732 2466 10766
rect 2500 10732 2516 10766
rect 2454 10715 2516 10732
rect 2546 10970 2612 10987
rect 2546 10936 2562 10970
rect 2596 10936 2612 10970
rect 2546 10902 2612 10936
rect 2546 10868 2562 10902
rect 2596 10868 2612 10902
rect 2546 10834 2612 10868
rect 2546 10800 2562 10834
rect 2596 10800 2612 10834
rect 2546 10766 2612 10800
rect 2546 10732 2562 10766
rect 2596 10732 2612 10766
rect 2546 10715 2612 10732
rect 2642 10970 2708 10987
rect 2642 10936 2658 10970
rect 2692 10936 2708 10970
rect 2642 10902 2708 10936
rect 2642 10868 2658 10902
rect 2692 10868 2708 10902
rect 2642 10834 2708 10868
rect 2642 10800 2658 10834
rect 2692 10800 2708 10834
rect 2642 10766 2708 10800
rect 2642 10732 2658 10766
rect 2692 10732 2708 10766
rect 2642 10715 2708 10732
rect 2738 10970 2804 10987
rect 2738 10936 2754 10970
rect 2788 10936 2804 10970
rect 2738 10902 2804 10936
rect 2738 10868 2754 10902
rect 2788 10868 2804 10902
rect 2738 10834 2804 10868
rect 2738 10800 2754 10834
rect 2788 10800 2804 10834
rect 2738 10766 2804 10800
rect 2738 10732 2754 10766
rect 2788 10732 2804 10766
rect 2738 10715 2804 10732
rect 2834 10970 2900 10987
rect 2834 10936 2850 10970
rect 2884 10936 2900 10970
rect 2834 10902 2900 10936
rect 2834 10868 2850 10902
rect 2884 10868 2900 10902
rect 2834 10834 2900 10868
rect 2834 10800 2850 10834
rect 2884 10800 2900 10834
rect 2834 10766 2900 10800
rect 2834 10732 2850 10766
rect 2884 10732 2900 10766
rect 2834 10715 2900 10732
rect 2930 10970 2996 10987
rect 2930 10936 2946 10970
rect 2980 10936 2996 10970
rect 2930 10902 2996 10936
rect 2930 10868 2946 10902
rect 2980 10868 2996 10902
rect 2930 10834 2996 10868
rect 2930 10800 2946 10834
rect 2980 10800 2996 10834
rect 2930 10766 2996 10800
rect 2930 10732 2946 10766
rect 2980 10732 2996 10766
rect 2930 10715 2996 10732
rect 3026 10970 3092 10987
rect 3026 10936 3042 10970
rect 3076 10936 3092 10970
rect 3026 10902 3092 10936
rect 3026 10868 3042 10902
rect 3076 10868 3092 10902
rect 3026 10834 3092 10868
rect 3026 10800 3042 10834
rect 3076 10800 3092 10834
rect 3026 10766 3092 10800
rect 3026 10732 3042 10766
rect 3076 10732 3092 10766
rect 3026 10715 3092 10732
rect 3122 10970 3188 10987
rect 3122 10936 3138 10970
rect 3172 10936 3188 10970
rect 3122 10902 3188 10936
rect 3122 10868 3138 10902
rect 3172 10868 3188 10902
rect 3122 10834 3188 10868
rect 3122 10800 3138 10834
rect 3172 10800 3188 10834
rect 3122 10766 3188 10800
rect 3122 10732 3138 10766
rect 3172 10732 3188 10766
rect 3122 10715 3188 10732
rect 3218 10970 3284 10987
rect 3218 10936 3234 10970
rect 3268 10936 3284 10970
rect 3218 10902 3284 10936
rect 3218 10868 3234 10902
rect 3268 10868 3284 10902
rect 3218 10834 3284 10868
rect 3218 10800 3234 10834
rect 3268 10800 3284 10834
rect 3218 10766 3284 10800
rect 3218 10732 3234 10766
rect 3268 10732 3284 10766
rect 3218 10715 3284 10732
rect 3314 10970 3380 10987
rect 3314 10936 3330 10970
rect 3364 10936 3380 10970
rect 3314 10902 3380 10936
rect 3314 10868 3330 10902
rect 3364 10868 3380 10902
rect 3314 10834 3380 10868
rect 3314 10800 3330 10834
rect 3364 10800 3380 10834
rect 3314 10766 3380 10800
rect 3314 10732 3330 10766
rect 3364 10732 3380 10766
rect 3314 10715 3380 10732
rect 3410 10970 3472 10987
rect 3410 10936 3426 10970
rect 3460 10936 3472 10970
rect 3410 10902 3472 10936
rect 3410 10868 3426 10902
rect 3460 10868 3472 10902
rect 3410 10834 3472 10868
rect 3410 10800 3426 10834
rect 3460 10800 3472 10834
rect 3410 10766 3472 10800
rect 3410 10732 3426 10766
rect 3460 10732 3472 10766
rect 3410 10715 3472 10732
rect 3975 10970 4037 10987
rect 3975 10936 3987 10970
rect 4021 10936 4037 10970
rect 3975 10902 4037 10936
rect 3975 10868 3987 10902
rect 4021 10868 4037 10902
rect 3975 10834 4037 10868
rect 3975 10800 3987 10834
rect 4021 10800 4037 10834
rect 3975 10766 4037 10800
rect 3975 10732 3987 10766
rect 4021 10732 4037 10766
rect 3975 10715 4037 10732
rect 4067 10970 4133 10987
rect 4067 10936 4083 10970
rect 4117 10936 4133 10970
rect 4067 10902 4133 10936
rect 4067 10868 4083 10902
rect 4117 10868 4133 10902
rect 4067 10834 4133 10868
rect 4067 10800 4083 10834
rect 4117 10800 4133 10834
rect 4067 10766 4133 10800
rect 4067 10732 4083 10766
rect 4117 10732 4133 10766
rect 4067 10715 4133 10732
rect 4163 10970 4229 10987
rect 4163 10936 4179 10970
rect 4213 10936 4229 10970
rect 4163 10902 4229 10936
rect 4163 10868 4179 10902
rect 4213 10868 4229 10902
rect 4163 10834 4229 10868
rect 4163 10800 4179 10834
rect 4213 10800 4229 10834
rect 4163 10766 4229 10800
rect 4163 10732 4179 10766
rect 4213 10732 4229 10766
rect 4163 10715 4229 10732
rect 4259 10970 4325 10987
rect 4259 10936 4275 10970
rect 4309 10936 4325 10970
rect 4259 10902 4325 10936
rect 4259 10868 4275 10902
rect 4309 10868 4325 10902
rect 4259 10834 4325 10868
rect 4259 10800 4275 10834
rect 4309 10800 4325 10834
rect 4259 10766 4325 10800
rect 4259 10732 4275 10766
rect 4309 10732 4325 10766
rect 4259 10715 4325 10732
rect 4355 10970 4421 10987
rect 4355 10936 4371 10970
rect 4405 10936 4421 10970
rect 4355 10902 4421 10936
rect 4355 10868 4371 10902
rect 4405 10868 4421 10902
rect 4355 10834 4421 10868
rect 4355 10800 4371 10834
rect 4405 10800 4421 10834
rect 4355 10766 4421 10800
rect 4355 10732 4371 10766
rect 4405 10732 4421 10766
rect 4355 10715 4421 10732
rect 4451 10970 4517 10987
rect 4451 10936 4467 10970
rect 4501 10936 4517 10970
rect 4451 10902 4517 10936
rect 4451 10868 4467 10902
rect 4501 10868 4517 10902
rect 4451 10834 4517 10868
rect 4451 10800 4467 10834
rect 4501 10800 4517 10834
rect 4451 10766 4517 10800
rect 4451 10732 4467 10766
rect 4501 10732 4517 10766
rect 4451 10715 4517 10732
rect 4547 10970 4613 10987
rect 4547 10936 4563 10970
rect 4597 10936 4613 10970
rect 4547 10902 4613 10936
rect 4547 10868 4563 10902
rect 4597 10868 4613 10902
rect 4547 10834 4613 10868
rect 4547 10800 4563 10834
rect 4597 10800 4613 10834
rect 4547 10766 4613 10800
rect 4547 10732 4563 10766
rect 4597 10732 4613 10766
rect 4547 10715 4613 10732
rect 4643 10970 4709 10987
rect 4643 10936 4659 10970
rect 4693 10936 4709 10970
rect 4643 10902 4709 10936
rect 4643 10868 4659 10902
rect 4693 10868 4709 10902
rect 4643 10834 4709 10868
rect 4643 10800 4659 10834
rect 4693 10800 4709 10834
rect 4643 10766 4709 10800
rect 4643 10732 4659 10766
rect 4693 10732 4709 10766
rect 4643 10715 4709 10732
rect 4739 10970 4805 10987
rect 4739 10936 4755 10970
rect 4789 10936 4805 10970
rect 4739 10902 4805 10936
rect 4739 10868 4755 10902
rect 4789 10868 4805 10902
rect 4739 10834 4805 10868
rect 4739 10800 4755 10834
rect 4789 10800 4805 10834
rect 4739 10766 4805 10800
rect 4739 10732 4755 10766
rect 4789 10732 4805 10766
rect 4739 10715 4805 10732
rect 4835 10970 4901 10987
rect 4835 10936 4851 10970
rect 4885 10936 4901 10970
rect 4835 10902 4901 10936
rect 4835 10868 4851 10902
rect 4885 10868 4901 10902
rect 4835 10834 4901 10868
rect 4835 10800 4851 10834
rect 4885 10800 4901 10834
rect 4835 10766 4901 10800
rect 4835 10732 4851 10766
rect 4885 10732 4901 10766
rect 4835 10715 4901 10732
rect 4931 10970 4993 10987
rect 4931 10936 4947 10970
rect 4981 10936 4993 10970
rect 4931 10902 4993 10936
rect 4931 10868 4947 10902
rect 4981 10868 4993 10902
rect 4931 10834 4993 10868
rect 4931 10800 4947 10834
rect 4981 10800 4993 10834
rect 4931 10766 4993 10800
rect 4931 10732 4947 10766
rect 4981 10732 4993 10766
rect 4931 10715 4993 10732
rect 5348 10762 5400 10774
rect 5348 10728 5356 10762
rect 5390 10728 5400 10762
rect 5348 10694 5400 10728
rect 5348 10660 5356 10694
rect 5390 10660 5400 10694
rect 5348 10626 5400 10660
rect 5348 10592 5356 10626
rect 5390 10592 5400 10626
rect 5348 10574 5400 10592
rect 5430 10762 5482 10774
rect 5430 10728 5440 10762
rect 5474 10728 5482 10762
rect 5430 10694 5482 10728
rect 5430 10660 5440 10694
rect 5474 10660 5482 10694
rect 5430 10626 5482 10660
rect 5430 10592 5440 10626
rect 5474 10592 5482 10626
rect 5430 10574 5482 10592
rect 301 9679 363 9696
rect 301 9645 313 9679
rect 347 9645 363 9679
rect 301 9611 363 9645
rect 301 9577 313 9611
rect 347 9577 363 9611
rect 301 9543 363 9577
rect 301 9509 313 9543
rect 347 9509 363 9543
rect 301 9475 363 9509
rect 301 9441 313 9475
rect 347 9441 363 9475
rect 301 9424 363 9441
rect 393 9679 459 9696
rect 393 9645 409 9679
rect 443 9645 459 9679
rect 393 9611 459 9645
rect 393 9577 409 9611
rect 443 9577 459 9611
rect 393 9543 459 9577
rect 393 9509 409 9543
rect 443 9509 459 9543
rect 393 9475 459 9509
rect 393 9441 409 9475
rect 443 9441 459 9475
rect 393 9424 459 9441
rect 489 9679 555 9696
rect 489 9645 505 9679
rect 539 9645 555 9679
rect 489 9611 555 9645
rect 489 9577 505 9611
rect 539 9577 555 9611
rect 489 9543 555 9577
rect 489 9509 505 9543
rect 539 9509 555 9543
rect 489 9475 555 9509
rect 489 9441 505 9475
rect 539 9441 555 9475
rect 489 9424 555 9441
rect 585 9679 651 9696
rect 585 9645 601 9679
rect 635 9645 651 9679
rect 585 9611 651 9645
rect 585 9577 601 9611
rect 635 9577 651 9611
rect 585 9543 651 9577
rect 585 9509 601 9543
rect 635 9509 651 9543
rect 585 9475 651 9509
rect 585 9441 601 9475
rect 635 9441 651 9475
rect 585 9424 651 9441
rect 681 9679 747 9696
rect 681 9645 697 9679
rect 731 9645 747 9679
rect 681 9611 747 9645
rect 681 9577 697 9611
rect 731 9577 747 9611
rect 681 9543 747 9577
rect 681 9509 697 9543
rect 731 9509 747 9543
rect 681 9475 747 9509
rect 681 9441 697 9475
rect 731 9441 747 9475
rect 681 9424 747 9441
rect 777 9679 843 9696
rect 777 9645 793 9679
rect 827 9645 843 9679
rect 777 9611 843 9645
rect 777 9577 793 9611
rect 827 9577 843 9611
rect 777 9543 843 9577
rect 777 9509 793 9543
rect 827 9509 843 9543
rect 777 9475 843 9509
rect 777 9441 793 9475
rect 827 9441 843 9475
rect 777 9424 843 9441
rect 873 9679 939 9696
rect 873 9645 889 9679
rect 923 9645 939 9679
rect 873 9611 939 9645
rect 873 9577 889 9611
rect 923 9577 939 9611
rect 873 9543 939 9577
rect 873 9509 889 9543
rect 923 9509 939 9543
rect 873 9475 939 9509
rect 873 9441 889 9475
rect 923 9441 939 9475
rect 873 9424 939 9441
rect 969 9679 1035 9696
rect 969 9645 985 9679
rect 1019 9645 1035 9679
rect 969 9611 1035 9645
rect 969 9577 985 9611
rect 1019 9577 1035 9611
rect 969 9543 1035 9577
rect 969 9509 985 9543
rect 1019 9509 1035 9543
rect 969 9475 1035 9509
rect 969 9441 985 9475
rect 1019 9441 1035 9475
rect 969 9424 1035 9441
rect 1065 9679 1131 9696
rect 1065 9645 1081 9679
rect 1115 9645 1131 9679
rect 1065 9611 1131 9645
rect 1065 9577 1081 9611
rect 1115 9577 1131 9611
rect 1065 9543 1131 9577
rect 1065 9509 1081 9543
rect 1115 9509 1131 9543
rect 1065 9475 1131 9509
rect 1065 9441 1081 9475
rect 1115 9441 1131 9475
rect 1065 9424 1131 9441
rect 1161 9679 1227 9696
rect 1161 9645 1177 9679
rect 1211 9645 1227 9679
rect 1161 9611 1227 9645
rect 1161 9577 1177 9611
rect 1211 9577 1227 9611
rect 1161 9543 1227 9577
rect 1161 9509 1177 9543
rect 1211 9509 1227 9543
rect 1161 9475 1227 9509
rect 1161 9441 1177 9475
rect 1211 9441 1227 9475
rect 1161 9424 1227 9441
rect 1257 9679 1319 9696
rect 1257 9645 1273 9679
rect 1307 9645 1319 9679
rect 1257 9611 1319 9645
rect 1257 9577 1273 9611
rect 1307 9577 1319 9611
rect 1257 9543 1319 9577
rect 1257 9509 1273 9543
rect 1307 9509 1319 9543
rect 1257 9475 1319 9509
rect 1257 9441 1273 9475
rect 1307 9441 1319 9475
rect 1257 9424 1319 9441
rect 2454 9683 2516 9700
rect 2454 9649 2466 9683
rect 2500 9649 2516 9683
rect 2454 9615 2516 9649
rect 2454 9581 2466 9615
rect 2500 9581 2516 9615
rect 2454 9547 2516 9581
rect 2454 9513 2466 9547
rect 2500 9513 2516 9547
rect 2454 9479 2516 9513
rect 2454 9445 2466 9479
rect 2500 9445 2516 9479
rect 2454 9428 2516 9445
rect 2546 9683 2612 9700
rect 2546 9649 2562 9683
rect 2596 9649 2612 9683
rect 2546 9615 2612 9649
rect 2546 9581 2562 9615
rect 2596 9581 2612 9615
rect 2546 9547 2612 9581
rect 2546 9513 2562 9547
rect 2596 9513 2612 9547
rect 2546 9479 2612 9513
rect 2546 9445 2562 9479
rect 2596 9445 2612 9479
rect 2546 9428 2612 9445
rect 2642 9683 2708 9700
rect 2642 9649 2658 9683
rect 2692 9649 2708 9683
rect 2642 9615 2708 9649
rect 2642 9581 2658 9615
rect 2692 9581 2708 9615
rect 2642 9547 2708 9581
rect 2642 9513 2658 9547
rect 2692 9513 2708 9547
rect 2642 9479 2708 9513
rect 2642 9445 2658 9479
rect 2692 9445 2708 9479
rect 2642 9428 2708 9445
rect 2738 9683 2804 9700
rect 2738 9649 2754 9683
rect 2788 9649 2804 9683
rect 2738 9615 2804 9649
rect 2738 9581 2754 9615
rect 2788 9581 2804 9615
rect 2738 9547 2804 9581
rect 2738 9513 2754 9547
rect 2788 9513 2804 9547
rect 2738 9479 2804 9513
rect 2738 9445 2754 9479
rect 2788 9445 2804 9479
rect 2738 9428 2804 9445
rect 2834 9683 2900 9700
rect 2834 9649 2850 9683
rect 2884 9649 2900 9683
rect 2834 9615 2900 9649
rect 2834 9581 2850 9615
rect 2884 9581 2900 9615
rect 2834 9547 2900 9581
rect 2834 9513 2850 9547
rect 2884 9513 2900 9547
rect 2834 9479 2900 9513
rect 2834 9445 2850 9479
rect 2884 9445 2900 9479
rect 2834 9428 2900 9445
rect 2930 9683 2996 9700
rect 2930 9649 2946 9683
rect 2980 9649 2996 9683
rect 2930 9615 2996 9649
rect 2930 9581 2946 9615
rect 2980 9581 2996 9615
rect 2930 9547 2996 9581
rect 2930 9513 2946 9547
rect 2980 9513 2996 9547
rect 2930 9479 2996 9513
rect 2930 9445 2946 9479
rect 2980 9445 2996 9479
rect 2930 9428 2996 9445
rect 3026 9683 3092 9700
rect 3026 9649 3042 9683
rect 3076 9649 3092 9683
rect 3026 9615 3092 9649
rect 3026 9581 3042 9615
rect 3076 9581 3092 9615
rect 3026 9547 3092 9581
rect 3026 9513 3042 9547
rect 3076 9513 3092 9547
rect 3026 9479 3092 9513
rect 3026 9445 3042 9479
rect 3076 9445 3092 9479
rect 3026 9428 3092 9445
rect 3122 9683 3188 9700
rect 3122 9649 3138 9683
rect 3172 9649 3188 9683
rect 3122 9615 3188 9649
rect 3122 9581 3138 9615
rect 3172 9581 3188 9615
rect 3122 9547 3188 9581
rect 3122 9513 3138 9547
rect 3172 9513 3188 9547
rect 3122 9479 3188 9513
rect 3122 9445 3138 9479
rect 3172 9445 3188 9479
rect 3122 9428 3188 9445
rect 3218 9683 3284 9700
rect 3218 9649 3234 9683
rect 3268 9649 3284 9683
rect 3218 9615 3284 9649
rect 3218 9581 3234 9615
rect 3268 9581 3284 9615
rect 3218 9547 3284 9581
rect 3218 9513 3234 9547
rect 3268 9513 3284 9547
rect 3218 9479 3284 9513
rect 3218 9445 3234 9479
rect 3268 9445 3284 9479
rect 3218 9428 3284 9445
rect 3314 9683 3380 9700
rect 3314 9649 3330 9683
rect 3364 9649 3380 9683
rect 3314 9615 3380 9649
rect 3314 9581 3330 9615
rect 3364 9581 3380 9615
rect 3314 9547 3380 9581
rect 3314 9513 3330 9547
rect 3364 9513 3380 9547
rect 3314 9479 3380 9513
rect 3314 9445 3330 9479
rect 3364 9445 3380 9479
rect 3314 9428 3380 9445
rect 3410 9683 3472 9700
rect 3410 9649 3426 9683
rect 3460 9649 3472 9683
rect 3410 9615 3472 9649
rect 3410 9581 3426 9615
rect 3460 9581 3472 9615
rect 3410 9547 3472 9581
rect 3410 9513 3426 9547
rect 3460 9513 3472 9547
rect 3410 9479 3472 9513
rect 3410 9445 3426 9479
rect 3460 9445 3472 9479
rect 3410 9428 3472 9445
rect 3975 9683 4037 9700
rect 3975 9649 3987 9683
rect 4021 9649 4037 9683
rect 3975 9615 4037 9649
rect 3975 9581 3987 9615
rect 4021 9581 4037 9615
rect 3975 9547 4037 9581
rect 3975 9513 3987 9547
rect 4021 9513 4037 9547
rect 3975 9479 4037 9513
rect 3975 9445 3987 9479
rect 4021 9445 4037 9479
rect 3975 9428 4037 9445
rect 4067 9683 4133 9700
rect 4067 9649 4083 9683
rect 4117 9649 4133 9683
rect 4067 9615 4133 9649
rect 4067 9581 4083 9615
rect 4117 9581 4133 9615
rect 4067 9547 4133 9581
rect 4067 9513 4083 9547
rect 4117 9513 4133 9547
rect 4067 9479 4133 9513
rect 4067 9445 4083 9479
rect 4117 9445 4133 9479
rect 4067 9428 4133 9445
rect 4163 9683 4229 9700
rect 4163 9649 4179 9683
rect 4213 9649 4229 9683
rect 4163 9615 4229 9649
rect 4163 9581 4179 9615
rect 4213 9581 4229 9615
rect 4163 9547 4229 9581
rect 4163 9513 4179 9547
rect 4213 9513 4229 9547
rect 4163 9479 4229 9513
rect 4163 9445 4179 9479
rect 4213 9445 4229 9479
rect 4163 9428 4229 9445
rect 4259 9683 4325 9700
rect 4259 9649 4275 9683
rect 4309 9649 4325 9683
rect 4259 9615 4325 9649
rect 4259 9581 4275 9615
rect 4309 9581 4325 9615
rect 4259 9547 4325 9581
rect 4259 9513 4275 9547
rect 4309 9513 4325 9547
rect 4259 9479 4325 9513
rect 4259 9445 4275 9479
rect 4309 9445 4325 9479
rect 4259 9428 4325 9445
rect 4355 9683 4421 9700
rect 4355 9649 4371 9683
rect 4405 9649 4421 9683
rect 4355 9615 4421 9649
rect 4355 9581 4371 9615
rect 4405 9581 4421 9615
rect 4355 9547 4421 9581
rect 4355 9513 4371 9547
rect 4405 9513 4421 9547
rect 4355 9479 4421 9513
rect 4355 9445 4371 9479
rect 4405 9445 4421 9479
rect 4355 9428 4421 9445
rect 4451 9683 4517 9700
rect 4451 9649 4467 9683
rect 4501 9649 4517 9683
rect 4451 9615 4517 9649
rect 4451 9581 4467 9615
rect 4501 9581 4517 9615
rect 4451 9547 4517 9581
rect 4451 9513 4467 9547
rect 4501 9513 4517 9547
rect 4451 9479 4517 9513
rect 4451 9445 4467 9479
rect 4501 9445 4517 9479
rect 4451 9428 4517 9445
rect 4547 9683 4613 9700
rect 4547 9649 4563 9683
rect 4597 9649 4613 9683
rect 4547 9615 4613 9649
rect 4547 9581 4563 9615
rect 4597 9581 4613 9615
rect 4547 9547 4613 9581
rect 4547 9513 4563 9547
rect 4597 9513 4613 9547
rect 4547 9479 4613 9513
rect 4547 9445 4563 9479
rect 4597 9445 4613 9479
rect 4547 9428 4613 9445
rect 4643 9683 4709 9700
rect 4643 9649 4659 9683
rect 4693 9649 4709 9683
rect 4643 9615 4709 9649
rect 4643 9581 4659 9615
rect 4693 9581 4709 9615
rect 4643 9547 4709 9581
rect 4643 9513 4659 9547
rect 4693 9513 4709 9547
rect 4643 9479 4709 9513
rect 4643 9445 4659 9479
rect 4693 9445 4709 9479
rect 4643 9428 4709 9445
rect 4739 9683 4805 9700
rect 4739 9649 4755 9683
rect 4789 9649 4805 9683
rect 4739 9615 4805 9649
rect 4739 9581 4755 9615
rect 4789 9581 4805 9615
rect 4739 9547 4805 9581
rect 4739 9513 4755 9547
rect 4789 9513 4805 9547
rect 4739 9479 4805 9513
rect 4739 9445 4755 9479
rect 4789 9445 4805 9479
rect 4739 9428 4805 9445
rect 4835 9683 4901 9700
rect 4835 9649 4851 9683
rect 4885 9649 4901 9683
rect 4835 9615 4901 9649
rect 4835 9581 4851 9615
rect 4885 9581 4901 9615
rect 4835 9547 4901 9581
rect 4835 9513 4851 9547
rect 4885 9513 4901 9547
rect 4835 9479 4901 9513
rect 4835 9445 4851 9479
rect 4885 9445 4901 9479
rect 4835 9428 4901 9445
rect 4931 9683 4993 9700
rect 4931 9649 4947 9683
rect 4981 9649 4993 9683
rect 4931 9615 4993 9649
rect 4931 9581 4947 9615
rect 4981 9581 4993 9615
rect 4931 9547 4993 9581
rect 4931 9513 4947 9547
rect 4981 9513 4993 9547
rect 4931 9479 4993 9513
rect 4931 9445 4947 9479
rect 4981 9445 4993 9479
rect 4931 9428 4993 9445
rect 5348 9475 5400 9487
rect 5348 9441 5356 9475
rect 5390 9441 5400 9475
rect 5348 9407 5400 9441
rect 5348 9373 5356 9407
rect 5390 9373 5400 9407
rect 5348 9339 5400 9373
rect 5348 9305 5356 9339
rect 5390 9305 5400 9339
rect 5348 9287 5400 9305
rect 5430 9475 5482 9487
rect 5430 9441 5440 9475
rect 5474 9441 5482 9475
rect 5430 9407 5482 9441
rect 5430 9373 5440 9407
rect 5474 9373 5482 9407
rect 5430 9339 5482 9373
rect 5430 9305 5440 9339
rect 5474 9305 5482 9339
rect 5430 9287 5482 9305
rect 301 8392 363 8409
rect 301 8358 313 8392
rect 347 8358 363 8392
rect 301 8324 363 8358
rect 301 8290 313 8324
rect 347 8290 363 8324
rect 301 8256 363 8290
rect 301 8222 313 8256
rect 347 8222 363 8256
rect 301 8188 363 8222
rect 301 8154 313 8188
rect 347 8154 363 8188
rect 301 8137 363 8154
rect 393 8392 459 8409
rect 393 8358 409 8392
rect 443 8358 459 8392
rect 393 8324 459 8358
rect 393 8290 409 8324
rect 443 8290 459 8324
rect 393 8256 459 8290
rect 393 8222 409 8256
rect 443 8222 459 8256
rect 393 8188 459 8222
rect 393 8154 409 8188
rect 443 8154 459 8188
rect 393 8137 459 8154
rect 489 8392 555 8409
rect 489 8358 505 8392
rect 539 8358 555 8392
rect 489 8324 555 8358
rect 489 8290 505 8324
rect 539 8290 555 8324
rect 489 8256 555 8290
rect 489 8222 505 8256
rect 539 8222 555 8256
rect 489 8188 555 8222
rect 489 8154 505 8188
rect 539 8154 555 8188
rect 489 8137 555 8154
rect 585 8392 651 8409
rect 585 8358 601 8392
rect 635 8358 651 8392
rect 585 8324 651 8358
rect 585 8290 601 8324
rect 635 8290 651 8324
rect 585 8256 651 8290
rect 585 8222 601 8256
rect 635 8222 651 8256
rect 585 8188 651 8222
rect 585 8154 601 8188
rect 635 8154 651 8188
rect 585 8137 651 8154
rect 681 8392 747 8409
rect 681 8358 697 8392
rect 731 8358 747 8392
rect 681 8324 747 8358
rect 681 8290 697 8324
rect 731 8290 747 8324
rect 681 8256 747 8290
rect 681 8222 697 8256
rect 731 8222 747 8256
rect 681 8188 747 8222
rect 681 8154 697 8188
rect 731 8154 747 8188
rect 681 8137 747 8154
rect 777 8392 843 8409
rect 777 8358 793 8392
rect 827 8358 843 8392
rect 777 8324 843 8358
rect 777 8290 793 8324
rect 827 8290 843 8324
rect 777 8256 843 8290
rect 777 8222 793 8256
rect 827 8222 843 8256
rect 777 8188 843 8222
rect 777 8154 793 8188
rect 827 8154 843 8188
rect 777 8137 843 8154
rect 873 8392 939 8409
rect 873 8358 889 8392
rect 923 8358 939 8392
rect 873 8324 939 8358
rect 873 8290 889 8324
rect 923 8290 939 8324
rect 873 8256 939 8290
rect 873 8222 889 8256
rect 923 8222 939 8256
rect 873 8188 939 8222
rect 873 8154 889 8188
rect 923 8154 939 8188
rect 873 8137 939 8154
rect 969 8392 1035 8409
rect 969 8358 985 8392
rect 1019 8358 1035 8392
rect 969 8324 1035 8358
rect 969 8290 985 8324
rect 1019 8290 1035 8324
rect 969 8256 1035 8290
rect 969 8222 985 8256
rect 1019 8222 1035 8256
rect 969 8188 1035 8222
rect 969 8154 985 8188
rect 1019 8154 1035 8188
rect 969 8137 1035 8154
rect 1065 8392 1131 8409
rect 1065 8358 1081 8392
rect 1115 8358 1131 8392
rect 1065 8324 1131 8358
rect 1065 8290 1081 8324
rect 1115 8290 1131 8324
rect 1065 8256 1131 8290
rect 1065 8222 1081 8256
rect 1115 8222 1131 8256
rect 1065 8188 1131 8222
rect 1065 8154 1081 8188
rect 1115 8154 1131 8188
rect 1065 8137 1131 8154
rect 1161 8392 1227 8409
rect 1161 8358 1177 8392
rect 1211 8358 1227 8392
rect 1161 8324 1227 8358
rect 1161 8290 1177 8324
rect 1211 8290 1227 8324
rect 1161 8256 1227 8290
rect 1161 8222 1177 8256
rect 1211 8222 1227 8256
rect 1161 8188 1227 8222
rect 1161 8154 1177 8188
rect 1211 8154 1227 8188
rect 1161 8137 1227 8154
rect 1257 8392 1319 8409
rect 1257 8358 1273 8392
rect 1307 8358 1319 8392
rect 1257 8324 1319 8358
rect 1257 8290 1273 8324
rect 1307 8290 1319 8324
rect 1257 8256 1319 8290
rect 1257 8222 1273 8256
rect 1307 8222 1319 8256
rect 1257 8188 1319 8222
rect 1257 8154 1273 8188
rect 1307 8154 1319 8188
rect 1257 8137 1319 8154
rect 2454 8396 2516 8413
rect 2454 8362 2466 8396
rect 2500 8362 2516 8396
rect 2454 8328 2516 8362
rect 2454 8294 2466 8328
rect 2500 8294 2516 8328
rect 2454 8260 2516 8294
rect 2454 8226 2466 8260
rect 2500 8226 2516 8260
rect 2454 8192 2516 8226
rect 2454 8158 2466 8192
rect 2500 8158 2516 8192
rect 2454 8141 2516 8158
rect 2546 8396 2612 8413
rect 2546 8362 2562 8396
rect 2596 8362 2612 8396
rect 2546 8328 2612 8362
rect 2546 8294 2562 8328
rect 2596 8294 2612 8328
rect 2546 8260 2612 8294
rect 2546 8226 2562 8260
rect 2596 8226 2612 8260
rect 2546 8192 2612 8226
rect 2546 8158 2562 8192
rect 2596 8158 2612 8192
rect 2546 8141 2612 8158
rect 2642 8396 2708 8413
rect 2642 8362 2658 8396
rect 2692 8362 2708 8396
rect 2642 8328 2708 8362
rect 2642 8294 2658 8328
rect 2692 8294 2708 8328
rect 2642 8260 2708 8294
rect 2642 8226 2658 8260
rect 2692 8226 2708 8260
rect 2642 8192 2708 8226
rect 2642 8158 2658 8192
rect 2692 8158 2708 8192
rect 2642 8141 2708 8158
rect 2738 8396 2804 8413
rect 2738 8362 2754 8396
rect 2788 8362 2804 8396
rect 2738 8328 2804 8362
rect 2738 8294 2754 8328
rect 2788 8294 2804 8328
rect 2738 8260 2804 8294
rect 2738 8226 2754 8260
rect 2788 8226 2804 8260
rect 2738 8192 2804 8226
rect 2738 8158 2754 8192
rect 2788 8158 2804 8192
rect 2738 8141 2804 8158
rect 2834 8396 2900 8413
rect 2834 8362 2850 8396
rect 2884 8362 2900 8396
rect 2834 8328 2900 8362
rect 2834 8294 2850 8328
rect 2884 8294 2900 8328
rect 2834 8260 2900 8294
rect 2834 8226 2850 8260
rect 2884 8226 2900 8260
rect 2834 8192 2900 8226
rect 2834 8158 2850 8192
rect 2884 8158 2900 8192
rect 2834 8141 2900 8158
rect 2930 8396 2996 8413
rect 2930 8362 2946 8396
rect 2980 8362 2996 8396
rect 2930 8328 2996 8362
rect 2930 8294 2946 8328
rect 2980 8294 2996 8328
rect 2930 8260 2996 8294
rect 2930 8226 2946 8260
rect 2980 8226 2996 8260
rect 2930 8192 2996 8226
rect 2930 8158 2946 8192
rect 2980 8158 2996 8192
rect 2930 8141 2996 8158
rect 3026 8396 3092 8413
rect 3026 8362 3042 8396
rect 3076 8362 3092 8396
rect 3026 8328 3092 8362
rect 3026 8294 3042 8328
rect 3076 8294 3092 8328
rect 3026 8260 3092 8294
rect 3026 8226 3042 8260
rect 3076 8226 3092 8260
rect 3026 8192 3092 8226
rect 3026 8158 3042 8192
rect 3076 8158 3092 8192
rect 3026 8141 3092 8158
rect 3122 8396 3188 8413
rect 3122 8362 3138 8396
rect 3172 8362 3188 8396
rect 3122 8328 3188 8362
rect 3122 8294 3138 8328
rect 3172 8294 3188 8328
rect 3122 8260 3188 8294
rect 3122 8226 3138 8260
rect 3172 8226 3188 8260
rect 3122 8192 3188 8226
rect 3122 8158 3138 8192
rect 3172 8158 3188 8192
rect 3122 8141 3188 8158
rect 3218 8396 3284 8413
rect 3218 8362 3234 8396
rect 3268 8362 3284 8396
rect 3218 8328 3284 8362
rect 3218 8294 3234 8328
rect 3268 8294 3284 8328
rect 3218 8260 3284 8294
rect 3218 8226 3234 8260
rect 3268 8226 3284 8260
rect 3218 8192 3284 8226
rect 3218 8158 3234 8192
rect 3268 8158 3284 8192
rect 3218 8141 3284 8158
rect 3314 8396 3380 8413
rect 3314 8362 3330 8396
rect 3364 8362 3380 8396
rect 3314 8328 3380 8362
rect 3314 8294 3330 8328
rect 3364 8294 3380 8328
rect 3314 8260 3380 8294
rect 3314 8226 3330 8260
rect 3364 8226 3380 8260
rect 3314 8192 3380 8226
rect 3314 8158 3330 8192
rect 3364 8158 3380 8192
rect 3314 8141 3380 8158
rect 3410 8396 3472 8413
rect 3410 8362 3426 8396
rect 3460 8362 3472 8396
rect 3410 8328 3472 8362
rect 3410 8294 3426 8328
rect 3460 8294 3472 8328
rect 3410 8260 3472 8294
rect 3410 8226 3426 8260
rect 3460 8226 3472 8260
rect 3410 8192 3472 8226
rect 3410 8158 3426 8192
rect 3460 8158 3472 8192
rect 3410 8141 3472 8158
rect 3975 8396 4037 8413
rect 3975 8362 3987 8396
rect 4021 8362 4037 8396
rect 3975 8328 4037 8362
rect 3975 8294 3987 8328
rect 4021 8294 4037 8328
rect 3975 8260 4037 8294
rect 3975 8226 3987 8260
rect 4021 8226 4037 8260
rect 3975 8192 4037 8226
rect 3975 8158 3987 8192
rect 4021 8158 4037 8192
rect 3975 8141 4037 8158
rect 4067 8396 4133 8413
rect 4067 8362 4083 8396
rect 4117 8362 4133 8396
rect 4067 8328 4133 8362
rect 4067 8294 4083 8328
rect 4117 8294 4133 8328
rect 4067 8260 4133 8294
rect 4067 8226 4083 8260
rect 4117 8226 4133 8260
rect 4067 8192 4133 8226
rect 4067 8158 4083 8192
rect 4117 8158 4133 8192
rect 4067 8141 4133 8158
rect 4163 8396 4229 8413
rect 4163 8362 4179 8396
rect 4213 8362 4229 8396
rect 4163 8328 4229 8362
rect 4163 8294 4179 8328
rect 4213 8294 4229 8328
rect 4163 8260 4229 8294
rect 4163 8226 4179 8260
rect 4213 8226 4229 8260
rect 4163 8192 4229 8226
rect 4163 8158 4179 8192
rect 4213 8158 4229 8192
rect 4163 8141 4229 8158
rect 4259 8396 4325 8413
rect 4259 8362 4275 8396
rect 4309 8362 4325 8396
rect 4259 8328 4325 8362
rect 4259 8294 4275 8328
rect 4309 8294 4325 8328
rect 4259 8260 4325 8294
rect 4259 8226 4275 8260
rect 4309 8226 4325 8260
rect 4259 8192 4325 8226
rect 4259 8158 4275 8192
rect 4309 8158 4325 8192
rect 4259 8141 4325 8158
rect 4355 8396 4421 8413
rect 4355 8362 4371 8396
rect 4405 8362 4421 8396
rect 4355 8328 4421 8362
rect 4355 8294 4371 8328
rect 4405 8294 4421 8328
rect 4355 8260 4421 8294
rect 4355 8226 4371 8260
rect 4405 8226 4421 8260
rect 4355 8192 4421 8226
rect 4355 8158 4371 8192
rect 4405 8158 4421 8192
rect 4355 8141 4421 8158
rect 4451 8396 4517 8413
rect 4451 8362 4467 8396
rect 4501 8362 4517 8396
rect 4451 8328 4517 8362
rect 4451 8294 4467 8328
rect 4501 8294 4517 8328
rect 4451 8260 4517 8294
rect 4451 8226 4467 8260
rect 4501 8226 4517 8260
rect 4451 8192 4517 8226
rect 4451 8158 4467 8192
rect 4501 8158 4517 8192
rect 4451 8141 4517 8158
rect 4547 8396 4613 8413
rect 4547 8362 4563 8396
rect 4597 8362 4613 8396
rect 4547 8328 4613 8362
rect 4547 8294 4563 8328
rect 4597 8294 4613 8328
rect 4547 8260 4613 8294
rect 4547 8226 4563 8260
rect 4597 8226 4613 8260
rect 4547 8192 4613 8226
rect 4547 8158 4563 8192
rect 4597 8158 4613 8192
rect 4547 8141 4613 8158
rect 4643 8396 4709 8413
rect 4643 8362 4659 8396
rect 4693 8362 4709 8396
rect 4643 8328 4709 8362
rect 4643 8294 4659 8328
rect 4693 8294 4709 8328
rect 4643 8260 4709 8294
rect 4643 8226 4659 8260
rect 4693 8226 4709 8260
rect 4643 8192 4709 8226
rect 4643 8158 4659 8192
rect 4693 8158 4709 8192
rect 4643 8141 4709 8158
rect 4739 8396 4805 8413
rect 4739 8362 4755 8396
rect 4789 8362 4805 8396
rect 4739 8328 4805 8362
rect 4739 8294 4755 8328
rect 4789 8294 4805 8328
rect 4739 8260 4805 8294
rect 4739 8226 4755 8260
rect 4789 8226 4805 8260
rect 4739 8192 4805 8226
rect 4739 8158 4755 8192
rect 4789 8158 4805 8192
rect 4739 8141 4805 8158
rect 4835 8396 4901 8413
rect 4835 8362 4851 8396
rect 4885 8362 4901 8396
rect 4835 8328 4901 8362
rect 4835 8294 4851 8328
rect 4885 8294 4901 8328
rect 4835 8260 4901 8294
rect 4835 8226 4851 8260
rect 4885 8226 4901 8260
rect 4835 8192 4901 8226
rect 4835 8158 4851 8192
rect 4885 8158 4901 8192
rect 4835 8141 4901 8158
rect 4931 8396 4993 8413
rect 4931 8362 4947 8396
rect 4981 8362 4993 8396
rect 4931 8328 4993 8362
rect 4931 8294 4947 8328
rect 4981 8294 4993 8328
rect 4931 8260 4993 8294
rect 4931 8226 4947 8260
rect 4981 8226 4993 8260
rect 4931 8192 4993 8226
rect 4931 8158 4947 8192
rect 4981 8158 4993 8192
rect 4931 8141 4993 8158
rect 5348 8188 5400 8200
rect 5348 8154 5356 8188
rect 5390 8154 5400 8188
rect 5348 8120 5400 8154
rect 5348 8086 5356 8120
rect 5390 8086 5400 8120
rect 5348 8052 5400 8086
rect 5348 8018 5356 8052
rect 5390 8018 5400 8052
rect 5348 8000 5400 8018
rect 5430 8188 5482 8200
rect 5430 8154 5440 8188
rect 5474 8154 5482 8188
rect 5430 8120 5482 8154
rect 5430 8086 5440 8120
rect 5474 8086 5482 8120
rect 5430 8052 5482 8086
rect 5430 8018 5440 8052
rect 5474 8018 5482 8052
rect 5430 8000 5482 8018
rect 301 7105 363 7122
rect 301 7071 313 7105
rect 347 7071 363 7105
rect 301 7037 363 7071
rect 301 7003 313 7037
rect 347 7003 363 7037
rect 301 6969 363 7003
rect 301 6935 313 6969
rect 347 6935 363 6969
rect 301 6901 363 6935
rect 301 6867 313 6901
rect 347 6867 363 6901
rect 301 6850 363 6867
rect 393 7105 459 7122
rect 393 7071 409 7105
rect 443 7071 459 7105
rect 393 7037 459 7071
rect 393 7003 409 7037
rect 443 7003 459 7037
rect 393 6969 459 7003
rect 393 6935 409 6969
rect 443 6935 459 6969
rect 393 6901 459 6935
rect 393 6867 409 6901
rect 443 6867 459 6901
rect 393 6850 459 6867
rect 489 7105 555 7122
rect 489 7071 505 7105
rect 539 7071 555 7105
rect 489 7037 555 7071
rect 489 7003 505 7037
rect 539 7003 555 7037
rect 489 6969 555 7003
rect 489 6935 505 6969
rect 539 6935 555 6969
rect 489 6901 555 6935
rect 489 6867 505 6901
rect 539 6867 555 6901
rect 489 6850 555 6867
rect 585 7105 651 7122
rect 585 7071 601 7105
rect 635 7071 651 7105
rect 585 7037 651 7071
rect 585 7003 601 7037
rect 635 7003 651 7037
rect 585 6969 651 7003
rect 585 6935 601 6969
rect 635 6935 651 6969
rect 585 6901 651 6935
rect 585 6867 601 6901
rect 635 6867 651 6901
rect 585 6850 651 6867
rect 681 7105 747 7122
rect 681 7071 697 7105
rect 731 7071 747 7105
rect 681 7037 747 7071
rect 681 7003 697 7037
rect 731 7003 747 7037
rect 681 6969 747 7003
rect 681 6935 697 6969
rect 731 6935 747 6969
rect 681 6901 747 6935
rect 681 6867 697 6901
rect 731 6867 747 6901
rect 681 6850 747 6867
rect 777 7105 843 7122
rect 777 7071 793 7105
rect 827 7071 843 7105
rect 777 7037 843 7071
rect 777 7003 793 7037
rect 827 7003 843 7037
rect 777 6969 843 7003
rect 777 6935 793 6969
rect 827 6935 843 6969
rect 777 6901 843 6935
rect 777 6867 793 6901
rect 827 6867 843 6901
rect 777 6850 843 6867
rect 873 7105 939 7122
rect 873 7071 889 7105
rect 923 7071 939 7105
rect 873 7037 939 7071
rect 873 7003 889 7037
rect 923 7003 939 7037
rect 873 6969 939 7003
rect 873 6935 889 6969
rect 923 6935 939 6969
rect 873 6901 939 6935
rect 873 6867 889 6901
rect 923 6867 939 6901
rect 873 6850 939 6867
rect 969 7105 1035 7122
rect 969 7071 985 7105
rect 1019 7071 1035 7105
rect 969 7037 1035 7071
rect 969 7003 985 7037
rect 1019 7003 1035 7037
rect 969 6969 1035 7003
rect 969 6935 985 6969
rect 1019 6935 1035 6969
rect 969 6901 1035 6935
rect 969 6867 985 6901
rect 1019 6867 1035 6901
rect 969 6850 1035 6867
rect 1065 7105 1131 7122
rect 1065 7071 1081 7105
rect 1115 7071 1131 7105
rect 1065 7037 1131 7071
rect 1065 7003 1081 7037
rect 1115 7003 1131 7037
rect 1065 6969 1131 7003
rect 1065 6935 1081 6969
rect 1115 6935 1131 6969
rect 1065 6901 1131 6935
rect 1065 6867 1081 6901
rect 1115 6867 1131 6901
rect 1065 6850 1131 6867
rect 1161 7105 1227 7122
rect 1161 7071 1177 7105
rect 1211 7071 1227 7105
rect 1161 7037 1227 7071
rect 1161 7003 1177 7037
rect 1211 7003 1227 7037
rect 1161 6969 1227 7003
rect 1161 6935 1177 6969
rect 1211 6935 1227 6969
rect 1161 6901 1227 6935
rect 1161 6867 1177 6901
rect 1211 6867 1227 6901
rect 1161 6850 1227 6867
rect 1257 7105 1319 7122
rect 1257 7071 1273 7105
rect 1307 7071 1319 7105
rect 1257 7037 1319 7071
rect 1257 7003 1273 7037
rect 1307 7003 1319 7037
rect 1257 6969 1319 7003
rect 1257 6935 1273 6969
rect 1307 6935 1319 6969
rect 1257 6901 1319 6935
rect 1257 6867 1273 6901
rect 1307 6867 1319 6901
rect 1257 6850 1319 6867
rect 2454 7109 2516 7126
rect 2454 7075 2466 7109
rect 2500 7075 2516 7109
rect 2454 7041 2516 7075
rect 2454 7007 2466 7041
rect 2500 7007 2516 7041
rect 2454 6973 2516 7007
rect 2454 6939 2466 6973
rect 2500 6939 2516 6973
rect 2454 6905 2516 6939
rect 2454 6871 2466 6905
rect 2500 6871 2516 6905
rect 2454 6854 2516 6871
rect 2546 7109 2612 7126
rect 2546 7075 2562 7109
rect 2596 7075 2612 7109
rect 2546 7041 2612 7075
rect 2546 7007 2562 7041
rect 2596 7007 2612 7041
rect 2546 6973 2612 7007
rect 2546 6939 2562 6973
rect 2596 6939 2612 6973
rect 2546 6905 2612 6939
rect 2546 6871 2562 6905
rect 2596 6871 2612 6905
rect 2546 6854 2612 6871
rect 2642 7109 2708 7126
rect 2642 7075 2658 7109
rect 2692 7075 2708 7109
rect 2642 7041 2708 7075
rect 2642 7007 2658 7041
rect 2692 7007 2708 7041
rect 2642 6973 2708 7007
rect 2642 6939 2658 6973
rect 2692 6939 2708 6973
rect 2642 6905 2708 6939
rect 2642 6871 2658 6905
rect 2692 6871 2708 6905
rect 2642 6854 2708 6871
rect 2738 7109 2804 7126
rect 2738 7075 2754 7109
rect 2788 7075 2804 7109
rect 2738 7041 2804 7075
rect 2738 7007 2754 7041
rect 2788 7007 2804 7041
rect 2738 6973 2804 7007
rect 2738 6939 2754 6973
rect 2788 6939 2804 6973
rect 2738 6905 2804 6939
rect 2738 6871 2754 6905
rect 2788 6871 2804 6905
rect 2738 6854 2804 6871
rect 2834 7109 2900 7126
rect 2834 7075 2850 7109
rect 2884 7075 2900 7109
rect 2834 7041 2900 7075
rect 2834 7007 2850 7041
rect 2884 7007 2900 7041
rect 2834 6973 2900 7007
rect 2834 6939 2850 6973
rect 2884 6939 2900 6973
rect 2834 6905 2900 6939
rect 2834 6871 2850 6905
rect 2884 6871 2900 6905
rect 2834 6854 2900 6871
rect 2930 7109 2996 7126
rect 2930 7075 2946 7109
rect 2980 7075 2996 7109
rect 2930 7041 2996 7075
rect 2930 7007 2946 7041
rect 2980 7007 2996 7041
rect 2930 6973 2996 7007
rect 2930 6939 2946 6973
rect 2980 6939 2996 6973
rect 2930 6905 2996 6939
rect 2930 6871 2946 6905
rect 2980 6871 2996 6905
rect 2930 6854 2996 6871
rect 3026 7109 3092 7126
rect 3026 7075 3042 7109
rect 3076 7075 3092 7109
rect 3026 7041 3092 7075
rect 3026 7007 3042 7041
rect 3076 7007 3092 7041
rect 3026 6973 3092 7007
rect 3026 6939 3042 6973
rect 3076 6939 3092 6973
rect 3026 6905 3092 6939
rect 3026 6871 3042 6905
rect 3076 6871 3092 6905
rect 3026 6854 3092 6871
rect 3122 7109 3188 7126
rect 3122 7075 3138 7109
rect 3172 7075 3188 7109
rect 3122 7041 3188 7075
rect 3122 7007 3138 7041
rect 3172 7007 3188 7041
rect 3122 6973 3188 7007
rect 3122 6939 3138 6973
rect 3172 6939 3188 6973
rect 3122 6905 3188 6939
rect 3122 6871 3138 6905
rect 3172 6871 3188 6905
rect 3122 6854 3188 6871
rect 3218 7109 3284 7126
rect 3218 7075 3234 7109
rect 3268 7075 3284 7109
rect 3218 7041 3284 7075
rect 3218 7007 3234 7041
rect 3268 7007 3284 7041
rect 3218 6973 3284 7007
rect 3218 6939 3234 6973
rect 3268 6939 3284 6973
rect 3218 6905 3284 6939
rect 3218 6871 3234 6905
rect 3268 6871 3284 6905
rect 3218 6854 3284 6871
rect 3314 7109 3380 7126
rect 3314 7075 3330 7109
rect 3364 7075 3380 7109
rect 3314 7041 3380 7075
rect 3314 7007 3330 7041
rect 3364 7007 3380 7041
rect 3314 6973 3380 7007
rect 3314 6939 3330 6973
rect 3364 6939 3380 6973
rect 3314 6905 3380 6939
rect 3314 6871 3330 6905
rect 3364 6871 3380 6905
rect 3314 6854 3380 6871
rect 3410 7109 3472 7126
rect 3410 7075 3426 7109
rect 3460 7075 3472 7109
rect 3410 7041 3472 7075
rect 3410 7007 3426 7041
rect 3460 7007 3472 7041
rect 3410 6973 3472 7007
rect 3410 6939 3426 6973
rect 3460 6939 3472 6973
rect 3410 6905 3472 6939
rect 3410 6871 3426 6905
rect 3460 6871 3472 6905
rect 3410 6854 3472 6871
rect 3975 7109 4037 7126
rect 3975 7075 3987 7109
rect 4021 7075 4037 7109
rect 3975 7041 4037 7075
rect 3975 7007 3987 7041
rect 4021 7007 4037 7041
rect 3975 6973 4037 7007
rect 3975 6939 3987 6973
rect 4021 6939 4037 6973
rect 3975 6905 4037 6939
rect 3975 6871 3987 6905
rect 4021 6871 4037 6905
rect 3975 6854 4037 6871
rect 4067 7109 4133 7126
rect 4067 7075 4083 7109
rect 4117 7075 4133 7109
rect 4067 7041 4133 7075
rect 4067 7007 4083 7041
rect 4117 7007 4133 7041
rect 4067 6973 4133 7007
rect 4067 6939 4083 6973
rect 4117 6939 4133 6973
rect 4067 6905 4133 6939
rect 4067 6871 4083 6905
rect 4117 6871 4133 6905
rect 4067 6854 4133 6871
rect 4163 7109 4229 7126
rect 4163 7075 4179 7109
rect 4213 7075 4229 7109
rect 4163 7041 4229 7075
rect 4163 7007 4179 7041
rect 4213 7007 4229 7041
rect 4163 6973 4229 7007
rect 4163 6939 4179 6973
rect 4213 6939 4229 6973
rect 4163 6905 4229 6939
rect 4163 6871 4179 6905
rect 4213 6871 4229 6905
rect 4163 6854 4229 6871
rect 4259 7109 4325 7126
rect 4259 7075 4275 7109
rect 4309 7075 4325 7109
rect 4259 7041 4325 7075
rect 4259 7007 4275 7041
rect 4309 7007 4325 7041
rect 4259 6973 4325 7007
rect 4259 6939 4275 6973
rect 4309 6939 4325 6973
rect 4259 6905 4325 6939
rect 4259 6871 4275 6905
rect 4309 6871 4325 6905
rect 4259 6854 4325 6871
rect 4355 7109 4421 7126
rect 4355 7075 4371 7109
rect 4405 7075 4421 7109
rect 4355 7041 4421 7075
rect 4355 7007 4371 7041
rect 4405 7007 4421 7041
rect 4355 6973 4421 7007
rect 4355 6939 4371 6973
rect 4405 6939 4421 6973
rect 4355 6905 4421 6939
rect 4355 6871 4371 6905
rect 4405 6871 4421 6905
rect 4355 6854 4421 6871
rect 4451 7109 4517 7126
rect 4451 7075 4467 7109
rect 4501 7075 4517 7109
rect 4451 7041 4517 7075
rect 4451 7007 4467 7041
rect 4501 7007 4517 7041
rect 4451 6973 4517 7007
rect 4451 6939 4467 6973
rect 4501 6939 4517 6973
rect 4451 6905 4517 6939
rect 4451 6871 4467 6905
rect 4501 6871 4517 6905
rect 4451 6854 4517 6871
rect 4547 7109 4613 7126
rect 4547 7075 4563 7109
rect 4597 7075 4613 7109
rect 4547 7041 4613 7075
rect 4547 7007 4563 7041
rect 4597 7007 4613 7041
rect 4547 6973 4613 7007
rect 4547 6939 4563 6973
rect 4597 6939 4613 6973
rect 4547 6905 4613 6939
rect 4547 6871 4563 6905
rect 4597 6871 4613 6905
rect 4547 6854 4613 6871
rect 4643 7109 4709 7126
rect 4643 7075 4659 7109
rect 4693 7075 4709 7109
rect 4643 7041 4709 7075
rect 4643 7007 4659 7041
rect 4693 7007 4709 7041
rect 4643 6973 4709 7007
rect 4643 6939 4659 6973
rect 4693 6939 4709 6973
rect 4643 6905 4709 6939
rect 4643 6871 4659 6905
rect 4693 6871 4709 6905
rect 4643 6854 4709 6871
rect 4739 7109 4805 7126
rect 4739 7075 4755 7109
rect 4789 7075 4805 7109
rect 4739 7041 4805 7075
rect 4739 7007 4755 7041
rect 4789 7007 4805 7041
rect 4739 6973 4805 7007
rect 4739 6939 4755 6973
rect 4789 6939 4805 6973
rect 4739 6905 4805 6939
rect 4739 6871 4755 6905
rect 4789 6871 4805 6905
rect 4739 6854 4805 6871
rect 4835 7109 4901 7126
rect 4835 7075 4851 7109
rect 4885 7075 4901 7109
rect 4835 7041 4901 7075
rect 4835 7007 4851 7041
rect 4885 7007 4901 7041
rect 4835 6973 4901 7007
rect 4835 6939 4851 6973
rect 4885 6939 4901 6973
rect 4835 6905 4901 6939
rect 4835 6871 4851 6905
rect 4885 6871 4901 6905
rect 4835 6854 4901 6871
rect 4931 7109 4993 7126
rect 4931 7075 4947 7109
rect 4981 7075 4993 7109
rect 4931 7041 4993 7075
rect 4931 7007 4947 7041
rect 4981 7007 4993 7041
rect 4931 6973 4993 7007
rect 4931 6939 4947 6973
rect 4981 6939 4993 6973
rect 4931 6905 4993 6939
rect 4931 6871 4947 6905
rect 4981 6871 4993 6905
rect 4931 6854 4993 6871
rect 5348 6901 5400 6913
rect 5348 6867 5356 6901
rect 5390 6867 5400 6901
rect 5348 6833 5400 6867
rect 5348 6799 5356 6833
rect 5390 6799 5400 6833
rect 5348 6765 5400 6799
rect 5348 6731 5356 6765
rect 5390 6731 5400 6765
rect 5348 6713 5400 6731
rect 5430 6901 5482 6913
rect 5430 6867 5440 6901
rect 5474 6867 5482 6901
rect 5430 6833 5482 6867
rect 5430 6799 5440 6833
rect 5474 6799 5482 6833
rect 5430 6765 5482 6799
rect 5430 6731 5440 6765
rect 5474 6731 5482 6765
rect 5430 6713 5482 6731
rect 301 5818 363 5835
rect 301 5784 313 5818
rect 347 5784 363 5818
rect 301 5750 363 5784
rect 301 5716 313 5750
rect 347 5716 363 5750
rect 301 5682 363 5716
rect 301 5648 313 5682
rect 347 5648 363 5682
rect 301 5614 363 5648
rect 301 5580 313 5614
rect 347 5580 363 5614
rect 301 5563 363 5580
rect 393 5818 459 5835
rect 393 5784 409 5818
rect 443 5784 459 5818
rect 393 5750 459 5784
rect 393 5716 409 5750
rect 443 5716 459 5750
rect 393 5682 459 5716
rect 393 5648 409 5682
rect 443 5648 459 5682
rect 393 5614 459 5648
rect 393 5580 409 5614
rect 443 5580 459 5614
rect 393 5563 459 5580
rect 489 5818 555 5835
rect 489 5784 505 5818
rect 539 5784 555 5818
rect 489 5750 555 5784
rect 489 5716 505 5750
rect 539 5716 555 5750
rect 489 5682 555 5716
rect 489 5648 505 5682
rect 539 5648 555 5682
rect 489 5614 555 5648
rect 489 5580 505 5614
rect 539 5580 555 5614
rect 489 5563 555 5580
rect 585 5818 651 5835
rect 585 5784 601 5818
rect 635 5784 651 5818
rect 585 5750 651 5784
rect 585 5716 601 5750
rect 635 5716 651 5750
rect 585 5682 651 5716
rect 585 5648 601 5682
rect 635 5648 651 5682
rect 585 5614 651 5648
rect 585 5580 601 5614
rect 635 5580 651 5614
rect 585 5563 651 5580
rect 681 5818 747 5835
rect 681 5784 697 5818
rect 731 5784 747 5818
rect 681 5750 747 5784
rect 681 5716 697 5750
rect 731 5716 747 5750
rect 681 5682 747 5716
rect 681 5648 697 5682
rect 731 5648 747 5682
rect 681 5614 747 5648
rect 681 5580 697 5614
rect 731 5580 747 5614
rect 681 5563 747 5580
rect 777 5818 843 5835
rect 777 5784 793 5818
rect 827 5784 843 5818
rect 777 5750 843 5784
rect 777 5716 793 5750
rect 827 5716 843 5750
rect 777 5682 843 5716
rect 777 5648 793 5682
rect 827 5648 843 5682
rect 777 5614 843 5648
rect 777 5580 793 5614
rect 827 5580 843 5614
rect 777 5563 843 5580
rect 873 5818 939 5835
rect 873 5784 889 5818
rect 923 5784 939 5818
rect 873 5750 939 5784
rect 873 5716 889 5750
rect 923 5716 939 5750
rect 873 5682 939 5716
rect 873 5648 889 5682
rect 923 5648 939 5682
rect 873 5614 939 5648
rect 873 5580 889 5614
rect 923 5580 939 5614
rect 873 5563 939 5580
rect 969 5818 1035 5835
rect 969 5784 985 5818
rect 1019 5784 1035 5818
rect 969 5750 1035 5784
rect 969 5716 985 5750
rect 1019 5716 1035 5750
rect 969 5682 1035 5716
rect 969 5648 985 5682
rect 1019 5648 1035 5682
rect 969 5614 1035 5648
rect 969 5580 985 5614
rect 1019 5580 1035 5614
rect 969 5563 1035 5580
rect 1065 5818 1131 5835
rect 1065 5784 1081 5818
rect 1115 5784 1131 5818
rect 1065 5750 1131 5784
rect 1065 5716 1081 5750
rect 1115 5716 1131 5750
rect 1065 5682 1131 5716
rect 1065 5648 1081 5682
rect 1115 5648 1131 5682
rect 1065 5614 1131 5648
rect 1065 5580 1081 5614
rect 1115 5580 1131 5614
rect 1065 5563 1131 5580
rect 1161 5818 1227 5835
rect 1161 5784 1177 5818
rect 1211 5784 1227 5818
rect 1161 5750 1227 5784
rect 1161 5716 1177 5750
rect 1211 5716 1227 5750
rect 1161 5682 1227 5716
rect 1161 5648 1177 5682
rect 1211 5648 1227 5682
rect 1161 5614 1227 5648
rect 1161 5580 1177 5614
rect 1211 5580 1227 5614
rect 1161 5563 1227 5580
rect 1257 5818 1319 5835
rect 1257 5784 1273 5818
rect 1307 5784 1319 5818
rect 1257 5750 1319 5784
rect 1257 5716 1273 5750
rect 1307 5716 1319 5750
rect 1257 5682 1319 5716
rect 1257 5648 1273 5682
rect 1307 5648 1319 5682
rect 1257 5614 1319 5648
rect 1257 5580 1273 5614
rect 1307 5580 1319 5614
rect 1257 5563 1319 5580
rect 2454 5822 2516 5839
rect 2454 5788 2466 5822
rect 2500 5788 2516 5822
rect 2454 5754 2516 5788
rect 2454 5720 2466 5754
rect 2500 5720 2516 5754
rect 2454 5686 2516 5720
rect 2454 5652 2466 5686
rect 2500 5652 2516 5686
rect 2454 5618 2516 5652
rect 2454 5584 2466 5618
rect 2500 5584 2516 5618
rect 2454 5567 2516 5584
rect 2546 5822 2612 5839
rect 2546 5788 2562 5822
rect 2596 5788 2612 5822
rect 2546 5754 2612 5788
rect 2546 5720 2562 5754
rect 2596 5720 2612 5754
rect 2546 5686 2612 5720
rect 2546 5652 2562 5686
rect 2596 5652 2612 5686
rect 2546 5618 2612 5652
rect 2546 5584 2562 5618
rect 2596 5584 2612 5618
rect 2546 5567 2612 5584
rect 2642 5822 2708 5839
rect 2642 5788 2658 5822
rect 2692 5788 2708 5822
rect 2642 5754 2708 5788
rect 2642 5720 2658 5754
rect 2692 5720 2708 5754
rect 2642 5686 2708 5720
rect 2642 5652 2658 5686
rect 2692 5652 2708 5686
rect 2642 5618 2708 5652
rect 2642 5584 2658 5618
rect 2692 5584 2708 5618
rect 2642 5567 2708 5584
rect 2738 5822 2804 5839
rect 2738 5788 2754 5822
rect 2788 5788 2804 5822
rect 2738 5754 2804 5788
rect 2738 5720 2754 5754
rect 2788 5720 2804 5754
rect 2738 5686 2804 5720
rect 2738 5652 2754 5686
rect 2788 5652 2804 5686
rect 2738 5618 2804 5652
rect 2738 5584 2754 5618
rect 2788 5584 2804 5618
rect 2738 5567 2804 5584
rect 2834 5822 2900 5839
rect 2834 5788 2850 5822
rect 2884 5788 2900 5822
rect 2834 5754 2900 5788
rect 2834 5720 2850 5754
rect 2884 5720 2900 5754
rect 2834 5686 2900 5720
rect 2834 5652 2850 5686
rect 2884 5652 2900 5686
rect 2834 5618 2900 5652
rect 2834 5584 2850 5618
rect 2884 5584 2900 5618
rect 2834 5567 2900 5584
rect 2930 5822 2996 5839
rect 2930 5788 2946 5822
rect 2980 5788 2996 5822
rect 2930 5754 2996 5788
rect 2930 5720 2946 5754
rect 2980 5720 2996 5754
rect 2930 5686 2996 5720
rect 2930 5652 2946 5686
rect 2980 5652 2996 5686
rect 2930 5618 2996 5652
rect 2930 5584 2946 5618
rect 2980 5584 2996 5618
rect 2930 5567 2996 5584
rect 3026 5822 3092 5839
rect 3026 5788 3042 5822
rect 3076 5788 3092 5822
rect 3026 5754 3092 5788
rect 3026 5720 3042 5754
rect 3076 5720 3092 5754
rect 3026 5686 3092 5720
rect 3026 5652 3042 5686
rect 3076 5652 3092 5686
rect 3026 5618 3092 5652
rect 3026 5584 3042 5618
rect 3076 5584 3092 5618
rect 3026 5567 3092 5584
rect 3122 5822 3188 5839
rect 3122 5788 3138 5822
rect 3172 5788 3188 5822
rect 3122 5754 3188 5788
rect 3122 5720 3138 5754
rect 3172 5720 3188 5754
rect 3122 5686 3188 5720
rect 3122 5652 3138 5686
rect 3172 5652 3188 5686
rect 3122 5618 3188 5652
rect 3122 5584 3138 5618
rect 3172 5584 3188 5618
rect 3122 5567 3188 5584
rect 3218 5822 3284 5839
rect 3218 5788 3234 5822
rect 3268 5788 3284 5822
rect 3218 5754 3284 5788
rect 3218 5720 3234 5754
rect 3268 5720 3284 5754
rect 3218 5686 3284 5720
rect 3218 5652 3234 5686
rect 3268 5652 3284 5686
rect 3218 5618 3284 5652
rect 3218 5584 3234 5618
rect 3268 5584 3284 5618
rect 3218 5567 3284 5584
rect 3314 5822 3380 5839
rect 3314 5788 3330 5822
rect 3364 5788 3380 5822
rect 3314 5754 3380 5788
rect 3314 5720 3330 5754
rect 3364 5720 3380 5754
rect 3314 5686 3380 5720
rect 3314 5652 3330 5686
rect 3364 5652 3380 5686
rect 3314 5618 3380 5652
rect 3314 5584 3330 5618
rect 3364 5584 3380 5618
rect 3314 5567 3380 5584
rect 3410 5822 3472 5839
rect 3410 5788 3426 5822
rect 3460 5788 3472 5822
rect 3410 5754 3472 5788
rect 3410 5720 3426 5754
rect 3460 5720 3472 5754
rect 3410 5686 3472 5720
rect 3410 5652 3426 5686
rect 3460 5652 3472 5686
rect 3410 5618 3472 5652
rect 3410 5584 3426 5618
rect 3460 5584 3472 5618
rect 3410 5567 3472 5584
rect 3975 5822 4037 5839
rect 3975 5788 3987 5822
rect 4021 5788 4037 5822
rect 3975 5754 4037 5788
rect 3975 5720 3987 5754
rect 4021 5720 4037 5754
rect 3975 5686 4037 5720
rect 3975 5652 3987 5686
rect 4021 5652 4037 5686
rect 3975 5618 4037 5652
rect 3975 5584 3987 5618
rect 4021 5584 4037 5618
rect 3975 5567 4037 5584
rect 4067 5822 4133 5839
rect 4067 5788 4083 5822
rect 4117 5788 4133 5822
rect 4067 5754 4133 5788
rect 4067 5720 4083 5754
rect 4117 5720 4133 5754
rect 4067 5686 4133 5720
rect 4067 5652 4083 5686
rect 4117 5652 4133 5686
rect 4067 5618 4133 5652
rect 4067 5584 4083 5618
rect 4117 5584 4133 5618
rect 4067 5567 4133 5584
rect 4163 5822 4229 5839
rect 4163 5788 4179 5822
rect 4213 5788 4229 5822
rect 4163 5754 4229 5788
rect 4163 5720 4179 5754
rect 4213 5720 4229 5754
rect 4163 5686 4229 5720
rect 4163 5652 4179 5686
rect 4213 5652 4229 5686
rect 4163 5618 4229 5652
rect 4163 5584 4179 5618
rect 4213 5584 4229 5618
rect 4163 5567 4229 5584
rect 4259 5822 4325 5839
rect 4259 5788 4275 5822
rect 4309 5788 4325 5822
rect 4259 5754 4325 5788
rect 4259 5720 4275 5754
rect 4309 5720 4325 5754
rect 4259 5686 4325 5720
rect 4259 5652 4275 5686
rect 4309 5652 4325 5686
rect 4259 5618 4325 5652
rect 4259 5584 4275 5618
rect 4309 5584 4325 5618
rect 4259 5567 4325 5584
rect 4355 5822 4421 5839
rect 4355 5788 4371 5822
rect 4405 5788 4421 5822
rect 4355 5754 4421 5788
rect 4355 5720 4371 5754
rect 4405 5720 4421 5754
rect 4355 5686 4421 5720
rect 4355 5652 4371 5686
rect 4405 5652 4421 5686
rect 4355 5618 4421 5652
rect 4355 5584 4371 5618
rect 4405 5584 4421 5618
rect 4355 5567 4421 5584
rect 4451 5822 4517 5839
rect 4451 5788 4467 5822
rect 4501 5788 4517 5822
rect 4451 5754 4517 5788
rect 4451 5720 4467 5754
rect 4501 5720 4517 5754
rect 4451 5686 4517 5720
rect 4451 5652 4467 5686
rect 4501 5652 4517 5686
rect 4451 5618 4517 5652
rect 4451 5584 4467 5618
rect 4501 5584 4517 5618
rect 4451 5567 4517 5584
rect 4547 5822 4613 5839
rect 4547 5788 4563 5822
rect 4597 5788 4613 5822
rect 4547 5754 4613 5788
rect 4547 5720 4563 5754
rect 4597 5720 4613 5754
rect 4547 5686 4613 5720
rect 4547 5652 4563 5686
rect 4597 5652 4613 5686
rect 4547 5618 4613 5652
rect 4547 5584 4563 5618
rect 4597 5584 4613 5618
rect 4547 5567 4613 5584
rect 4643 5822 4709 5839
rect 4643 5788 4659 5822
rect 4693 5788 4709 5822
rect 4643 5754 4709 5788
rect 4643 5720 4659 5754
rect 4693 5720 4709 5754
rect 4643 5686 4709 5720
rect 4643 5652 4659 5686
rect 4693 5652 4709 5686
rect 4643 5618 4709 5652
rect 4643 5584 4659 5618
rect 4693 5584 4709 5618
rect 4643 5567 4709 5584
rect 4739 5822 4805 5839
rect 4739 5788 4755 5822
rect 4789 5788 4805 5822
rect 4739 5754 4805 5788
rect 4739 5720 4755 5754
rect 4789 5720 4805 5754
rect 4739 5686 4805 5720
rect 4739 5652 4755 5686
rect 4789 5652 4805 5686
rect 4739 5618 4805 5652
rect 4739 5584 4755 5618
rect 4789 5584 4805 5618
rect 4739 5567 4805 5584
rect 4835 5822 4901 5839
rect 4835 5788 4851 5822
rect 4885 5788 4901 5822
rect 4835 5754 4901 5788
rect 4835 5720 4851 5754
rect 4885 5720 4901 5754
rect 4835 5686 4901 5720
rect 4835 5652 4851 5686
rect 4885 5652 4901 5686
rect 4835 5618 4901 5652
rect 4835 5584 4851 5618
rect 4885 5584 4901 5618
rect 4835 5567 4901 5584
rect 4931 5822 4993 5839
rect 4931 5788 4947 5822
rect 4981 5788 4993 5822
rect 4931 5754 4993 5788
rect 4931 5720 4947 5754
rect 4981 5720 4993 5754
rect 4931 5686 4993 5720
rect 4931 5652 4947 5686
rect 4981 5652 4993 5686
rect 4931 5618 4993 5652
rect 4931 5584 4947 5618
rect 4981 5584 4993 5618
rect 4931 5567 4993 5584
rect 5348 5614 5400 5626
rect 5348 5580 5356 5614
rect 5390 5580 5400 5614
rect 5348 5546 5400 5580
rect 5348 5512 5356 5546
rect 5390 5512 5400 5546
rect 5348 5478 5400 5512
rect 5348 5444 5356 5478
rect 5390 5444 5400 5478
rect 5348 5426 5400 5444
rect 5430 5614 5482 5626
rect 5430 5580 5440 5614
rect 5474 5580 5482 5614
rect 5430 5546 5482 5580
rect 5430 5512 5440 5546
rect 5474 5512 5482 5546
rect 5430 5478 5482 5512
rect 5430 5444 5440 5478
rect 5474 5444 5482 5478
rect 5430 5426 5482 5444
rect 301 4531 363 4548
rect 301 4497 313 4531
rect 347 4497 363 4531
rect 301 4463 363 4497
rect 301 4429 313 4463
rect 347 4429 363 4463
rect 301 4395 363 4429
rect 301 4361 313 4395
rect 347 4361 363 4395
rect 301 4327 363 4361
rect 301 4293 313 4327
rect 347 4293 363 4327
rect 301 4276 363 4293
rect 393 4531 459 4548
rect 393 4497 409 4531
rect 443 4497 459 4531
rect 393 4463 459 4497
rect 393 4429 409 4463
rect 443 4429 459 4463
rect 393 4395 459 4429
rect 393 4361 409 4395
rect 443 4361 459 4395
rect 393 4327 459 4361
rect 393 4293 409 4327
rect 443 4293 459 4327
rect 393 4276 459 4293
rect 489 4531 555 4548
rect 489 4497 505 4531
rect 539 4497 555 4531
rect 489 4463 555 4497
rect 489 4429 505 4463
rect 539 4429 555 4463
rect 489 4395 555 4429
rect 489 4361 505 4395
rect 539 4361 555 4395
rect 489 4327 555 4361
rect 489 4293 505 4327
rect 539 4293 555 4327
rect 489 4276 555 4293
rect 585 4531 651 4548
rect 585 4497 601 4531
rect 635 4497 651 4531
rect 585 4463 651 4497
rect 585 4429 601 4463
rect 635 4429 651 4463
rect 585 4395 651 4429
rect 585 4361 601 4395
rect 635 4361 651 4395
rect 585 4327 651 4361
rect 585 4293 601 4327
rect 635 4293 651 4327
rect 585 4276 651 4293
rect 681 4531 747 4548
rect 681 4497 697 4531
rect 731 4497 747 4531
rect 681 4463 747 4497
rect 681 4429 697 4463
rect 731 4429 747 4463
rect 681 4395 747 4429
rect 681 4361 697 4395
rect 731 4361 747 4395
rect 681 4327 747 4361
rect 681 4293 697 4327
rect 731 4293 747 4327
rect 681 4276 747 4293
rect 777 4531 843 4548
rect 777 4497 793 4531
rect 827 4497 843 4531
rect 777 4463 843 4497
rect 777 4429 793 4463
rect 827 4429 843 4463
rect 777 4395 843 4429
rect 777 4361 793 4395
rect 827 4361 843 4395
rect 777 4327 843 4361
rect 777 4293 793 4327
rect 827 4293 843 4327
rect 777 4276 843 4293
rect 873 4531 939 4548
rect 873 4497 889 4531
rect 923 4497 939 4531
rect 873 4463 939 4497
rect 873 4429 889 4463
rect 923 4429 939 4463
rect 873 4395 939 4429
rect 873 4361 889 4395
rect 923 4361 939 4395
rect 873 4327 939 4361
rect 873 4293 889 4327
rect 923 4293 939 4327
rect 873 4276 939 4293
rect 969 4531 1035 4548
rect 969 4497 985 4531
rect 1019 4497 1035 4531
rect 969 4463 1035 4497
rect 969 4429 985 4463
rect 1019 4429 1035 4463
rect 969 4395 1035 4429
rect 969 4361 985 4395
rect 1019 4361 1035 4395
rect 969 4327 1035 4361
rect 969 4293 985 4327
rect 1019 4293 1035 4327
rect 969 4276 1035 4293
rect 1065 4531 1131 4548
rect 1065 4497 1081 4531
rect 1115 4497 1131 4531
rect 1065 4463 1131 4497
rect 1065 4429 1081 4463
rect 1115 4429 1131 4463
rect 1065 4395 1131 4429
rect 1065 4361 1081 4395
rect 1115 4361 1131 4395
rect 1065 4327 1131 4361
rect 1065 4293 1081 4327
rect 1115 4293 1131 4327
rect 1065 4276 1131 4293
rect 1161 4531 1227 4548
rect 1161 4497 1177 4531
rect 1211 4497 1227 4531
rect 1161 4463 1227 4497
rect 1161 4429 1177 4463
rect 1211 4429 1227 4463
rect 1161 4395 1227 4429
rect 1161 4361 1177 4395
rect 1211 4361 1227 4395
rect 1161 4327 1227 4361
rect 1161 4293 1177 4327
rect 1211 4293 1227 4327
rect 1161 4276 1227 4293
rect 1257 4531 1319 4548
rect 1257 4497 1273 4531
rect 1307 4497 1319 4531
rect 1257 4463 1319 4497
rect 1257 4429 1273 4463
rect 1307 4429 1319 4463
rect 1257 4395 1319 4429
rect 1257 4361 1273 4395
rect 1307 4361 1319 4395
rect 1257 4327 1319 4361
rect 1257 4293 1273 4327
rect 1307 4293 1319 4327
rect 1257 4276 1319 4293
rect 2454 4535 2516 4552
rect 2454 4501 2466 4535
rect 2500 4501 2516 4535
rect 2454 4467 2516 4501
rect 2454 4433 2466 4467
rect 2500 4433 2516 4467
rect 2454 4399 2516 4433
rect 2454 4365 2466 4399
rect 2500 4365 2516 4399
rect 2454 4331 2516 4365
rect 2454 4297 2466 4331
rect 2500 4297 2516 4331
rect 2454 4280 2516 4297
rect 2546 4535 2612 4552
rect 2546 4501 2562 4535
rect 2596 4501 2612 4535
rect 2546 4467 2612 4501
rect 2546 4433 2562 4467
rect 2596 4433 2612 4467
rect 2546 4399 2612 4433
rect 2546 4365 2562 4399
rect 2596 4365 2612 4399
rect 2546 4331 2612 4365
rect 2546 4297 2562 4331
rect 2596 4297 2612 4331
rect 2546 4280 2612 4297
rect 2642 4535 2708 4552
rect 2642 4501 2658 4535
rect 2692 4501 2708 4535
rect 2642 4467 2708 4501
rect 2642 4433 2658 4467
rect 2692 4433 2708 4467
rect 2642 4399 2708 4433
rect 2642 4365 2658 4399
rect 2692 4365 2708 4399
rect 2642 4331 2708 4365
rect 2642 4297 2658 4331
rect 2692 4297 2708 4331
rect 2642 4280 2708 4297
rect 2738 4535 2804 4552
rect 2738 4501 2754 4535
rect 2788 4501 2804 4535
rect 2738 4467 2804 4501
rect 2738 4433 2754 4467
rect 2788 4433 2804 4467
rect 2738 4399 2804 4433
rect 2738 4365 2754 4399
rect 2788 4365 2804 4399
rect 2738 4331 2804 4365
rect 2738 4297 2754 4331
rect 2788 4297 2804 4331
rect 2738 4280 2804 4297
rect 2834 4535 2900 4552
rect 2834 4501 2850 4535
rect 2884 4501 2900 4535
rect 2834 4467 2900 4501
rect 2834 4433 2850 4467
rect 2884 4433 2900 4467
rect 2834 4399 2900 4433
rect 2834 4365 2850 4399
rect 2884 4365 2900 4399
rect 2834 4331 2900 4365
rect 2834 4297 2850 4331
rect 2884 4297 2900 4331
rect 2834 4280 2900 4297
rect 2930 4535 2996 4552
rect 2930 4501 2946 4535
rect 2980 4501 2996 4535
rect 2930 4467 2996 4501
rect 2930 4433 2946 4467
rect 2980 4433 2996 4467
rect 2930 4399 2996 4433
rect 2930 4365 2946 4399
rect 2980 4365 2996 4399
rect 2930 4331 2996 4365
rect 2930 4297 2946 4331
rect 2980 4297 2996 4331
rect 2930 4280 2996 4297
rect 3026 4535 3092 4552
rect 3026 4501 3042 4535
rect 3076 4501 3092 4535
rect 3026 4467 3092 4501
rect 3026 4433 3042 4467
rect 3076 4433 3092 4467
rect 3026 4399 3092 4433
rect 3026 4365 3042 4399
rect 3076 4365 3092 4399
rect 3026 4331 3092 4365
rect 3026 4297 3042 4331
rect 3076 4297 3092 4331
rect 3026 4280 3092 4297
rect 3122 4535 3188 4552
rect 3122 4501 3138 4535
rect 3172 4501 3188 4535
rect 3122 4467 3188 4501
rect 3122 4433 3138 4467
rect 3172 4433 3188 4467
rect 3122 4399 3188 4433
rect 3122 4365 3138 4399
rect 3172 4365 3188 4399
rect 3122 4331 3188 4365
rect 3122 4297 3138 4331
rect 3172 4297 3188 4331
rect 3122 4280 3188 4297
rect 3218 4535 3284 4552
rect 3218 4501 3234 4535
rect 3268 4501 3284 4535
rect 3218 4467 3284 4501
rect 3218 4433 3234 4467
rect 3268 4433 3284 4467
rect 3218 4399 3284 4433
rect 3218 4365 3234 4399
rect 3268 4365 3284 4399
rect 3218 4331 3284 4365
rect 3218 4297 3234 4331
rect 3268 4297 3284 4331
rect 3218 4280 3284 4297
rect 3314 4535 3380 4552
rect 3314 4501 3330 4535
rect 3364 4501 3380 4535
rect 3314 4467 3380 4501
rect 3314 4433 3330 4467
rect 3364 4433 3380 4467
rect 3314 4399 3380 4433
rect 3314 4365 3330 4399
rect 3364 4365 3380 4399
rect 3314 4331 3380 4365
rect 3314 4297 3330 4331
rect 3364 4297 3380 4331
rect 3314 4280 3380 4297
rect 3410 4535 3472 4552
rect 3410 4501 3426 4535
rect 3460 4501 3472 4535
rect 3410 4467 3472 4501
rect 3410 4433 3426 4467
rect 3460 4433 3472 4467
rect 3410 4399 3472 4433
rect 3410 4365 3426 4399
rect 3460 4365 3472 4399
rect 3410 4331 3472 4365
rect 3410 4297 3426 4331
rect 3460 4297 3472 4331
rect 3410 4280 3472 4297
rect 3975 4535 4037 4552
rect 3975 4501 3987 4535
rect 4021 4501 4037 4535
rect 3975 4467 4037 4501
rect 3975 4433 3987 4467
rect 4021 4433 4037 4467
rect 3975 4399 4037 4433
rect 3975 4365 3987 4399
rect 4021 4365 4037 4399
rect 3975 4331 4037 4365
rect 3975 4297 3987 4331
rect 4021 4297 4037 4331
rect 3975 4280 4037 4297
rect 4067 4535 4133 4552
rect 4067 4501 4083 4535
rect 4117 4501 4133 4535
rect 4067 4467 4133 4501
rect 4067 4433 4083 4467
rect 4117 4433 4133 4467
rect 4067 4399 4133 4433
rect 4067 4365 4083 4399
rect 4117 4365 4133 4399
rect 4067 4331 4133 4365
rect 4067 4297 4083 4331
rect 4117 4297 4133 4331
rect 4067 4280 4133 4297
rect 4163 4535 4229 4552
rect 4163 4501 4179 4535
rect 4213 4501 4229 4535
rect 4163 4467 4229 4501
rect 4163 4433 4179 4467
rect 4213 4433 4229 4467
rect 4163 4399 4229 4433
rect 4163 4365 4179 4399
rect 4213 4365 4229 4399
rect 4163 4331 4229 4365
rect 4163 4297 4179 4331
rect 4213 4297 4229 4331
rect 4163 4280 4229 4297
rect 4259 4535 4325 4552
rect 4259 4501 4275 4535
rect 4309 4501 4325 4535
rect 4259 4467 4325 4501
rect 4259 4433 4275 4467
rect 4309 4433 4325 4467
rect 4259 4399 4325 4433
rect 4259 4365 4275 4399
rect 4309 4365 4325 4399
rect 4259 4331 4325 4365
rect 4259 4297 4275 4331
rect 4309 4297 4325 4331
rect 4259 4280 4325 4297
rect 4355 4535 4421 4552
rect 4355 4501 4371 4535
rect 4405 4501 4421 4535
rect 4355 4467 4421 4501
rect 4355 4433 4371 4467
rect 4405 4433 4421 4467
rect 4355 4399 4421 4433
rect 4355 4365 4371 4399
rect 4405 4365 4421 4399
rect 4355 4331 4421 4365
rect 4355 4297 4371 4331
rect 4405 4297 4421 4331
rect 4355 4280 4421 4297
rect 4451 4535 4517 4552
rect 4451 4501 4467 4535
rect 4501 4501 4517 4535
rect 4451 4467 4517 4501
rect 4451 4433 4467 4467
rect 4501 4433 4517 4467
rect 4451 4399 4517 4433
rect 4451 4365 4467 4399
rect 4501 4365 4517 4399
rect 4451 4331 4517 4365
rect 4451 4297 4467 4331
rect 4501 4297 4517 4331
rect 4451 4280 4517 4297
rect 4547 4535 4613 4552
rect 4547 4501 4563 4535
rect 4597 4501 4613 4535
rect 4547 4467 4613 4501
rect 4547 4433 4563 4467
rect 4597 4433 4613 4467
rect 4547 4399 4613 4433
rect 4547 4365 4563 4399
rect 4597 4365 4613 4399
rect 4547 4331 4613 4365
rect 4547 4297 4563 4331
rect 4597 4297 4613 4331
rect 4547 4280 4613 4297
rect 4643 4535 4709 4552
rect 4643 4501 4659 4535
rect 4693 4501 4709 4535
rect 4643 4467 4709 4501
rect 4643 4433 4659 4467
rect 4693 4433 4709 4467
rect 4643 4399 4709 4433
rect 4643 4365 4659 4399
rect 4693 4365 4709 4399
rect 4643 4331 4709 4365
rect 4643 4297 4659 4331
rect 4693 4297 4709 4331
rect 4643 4280 4709 4297
rect 4739 4535 4805 4552
rect 4739 4501 4755 4535
rect 4789 4501 4805 4535
rect 4739 4467 4805 4501
rect 4739 4433 4755 4467
rect 4789 4433 4805 4467
rect 4739 4399 4805 4433
rect 4739 4365 4755 4399
rect 4789 4365 4805 4399
rect 4739 4331 4805 4365
rect 4739 4297 4755 4331
rect 4789 4297 4805 4331
rect 4739 4280 4805 4297
rect 4835 4535 4901 4552
rect 4835 4501 4851 4535
rect 4885 4501 4901 4535
rect 4835 4467 4901 4501
rect 4835 4433 4851 4467
rect 4885 4433 4901 4467
rect 4835 4399 4901 4433
rect 4835 4365 4851 4399
rect 4885 4365 4901 4399
rect 4835 4331 4901 4365
rect 4835 4297 4851 4331
rect 4885 4297 4901 4331
rect 4835 4280 4901 4297
rect 4931 4535 4993 4552
rect 4931 4501 4947 4535
rect 4981 4501 4993 4535
rect 4931 4467 4993 4501
rect 4931 4433 4947 4467
rect 4981 4433 4993 4467
rect 4931 4399 4993 4433
rect 4931 4365 4947 4399
rect 4981 4365 4993 4399
rect 4931 4331 4993 4365
rect 4931 4297 4947 4331
rect 4981 4297 4993 4331
rect 4931 4280 4993 4297
rect 5348 4327 5400 4339
rect 5348 4293 5356 4327
rect 5390 4293 5400 4327
rect 5348 4259 5400 4293
rect 5348 4225 5356 4259
rect 5390 4225 5400 4259
rect 5348 4191 5400 4225
rect 5348 4157 5356 4191
rect 5390 4157 5400 4191
rect 5348 4139 5400 4157
rect 5430 4327 5482 4339
rect 5430 4293 5440 4327
rect 5474 4293 5482 4327
rect 5430 4259 5482 4293
rect 5430 4225 5440 4259
rect 5474 4225 5482 4259
rect 5430 4191 5482 4225
rect 5430 4157 5440 4191
rect 5474 4157 5482 4191
rect 5430 4139 5482 4157
rect 301 3244 363 3261
rect 301 3210 313 3244
rect 347 3210 363 3244
rect 301 3176 363 3210
rect 301 3142 313 3176
rect 347 3142 363 3176
rect 301 3108 363 3142
rect 301 3074 313 3108
rect 347 3074 363 3108
rect 301 3040 363 3074
rect 301 3006 313 3040
rect 347 3006 363 3040
rect 301 2989 363 3006
rect 393 3244 459 3261
rect 393 3210 409 3244
rect 443 3210 459 3244
rect 393 3176 459 3210
rect 393 3142 409 3176
rect 443 3142 459 3176
rect 393 3108 459 3142
rect 393 3074 409 3108
rect 443 3074 459 3108
rect 393 3040 459 3074
rect 393 3006 409 3040
rect 443 3006 459 3040
rect 393 2989 459 3006
rect 489 3244 555 3261
rect 489 3210 505 3244
rect 539 3210 555 3244
rect 489 3176 555 3210
rect 489 3142 505 3176
rect 539 3142 555 3176
rect 489 3108 555 3142
rect 489 3074 505 3108
rect 539 3074 555 3108
rect 489 3040 555 3074
rect 489 3006 505 3040
rect 539 3006 555 3040
rect 489 2989 555 3006
rect 585 3244 651 3261
rect 585 3210 601 3244
rect 635 3210 651 3244
rect 585 3176 651 3210
rect 585 3142 601 3176
rect 635 3142 651 3176
rect 585 3108 651 3142
rect 585 3074 601 3108
rect 635 3074 651 3108
rect 585 3040 651 3074
rect 585 3006 601 3040
rect 635 3006 651 3040
rect 585 2989 651 3006
rect 681 3244 747 3261
rect 681 3210 697 3244
rect 731 3210 747 3244
rect 681 3176 747 3210
rect 681 3142 697 3176
rect 731 3142 747 3176
rect 681 3108 747 3142
rect 681 3074 697 3108
rect 731 3074 747 3108
rect 681 3040 747 3074
rect 681 3006 697 3040
rect 731 3006 747 3040
rect 681 2989 747 3006
rect 777 3244 843 3261
rect 777 3210 793 3244
rect 827 3210 843 3244
rect 777 3176 843 3210
rect 777 3142 793 3176
rect 827 3142 843 3176
rect 777 3108 843 3142
rect 777 3074 793 3108
rect 827 3074 843 3108
rect 777 3040 843 3074
rect 777 3006 793 3040
rect 827 3006 843 3040
rect 777 2989 843 3006
rect 873 3244 939 3261
rect 873 3210 889 3244
rect 923 3210 939 3244
rect 873 3176 939 3210
rect 873 3142 889 3176
rect 923 3142 939 3176
rect 873 3108 939 3142
rect 873 3074 889 3108
rect 923 3074 939 3108
rect 873 3040 939 3074
rect 873 3006 889 3040
rect 923 3006 939 3040
rect 873 2989 939 3006
rect 969 3244 1035 3261
rect 969 3210 985 3244
rect 1019 3210 1035 3244
rect 969 3176 1035 3210
rect 969 3142 985 3176
rect 1019 3142 1035 3176
rect 969 3108 1035 3142
rect 969 3074 985 3108
rect 1019 3074 1035 3108
rect 969 3040 1035 3074
rect 969 3006 985 3040
rect 1019 3006 1035 3040
rect 969 2989 1035 3006
rect 1065 3244 1131 3261
rect 1065 3210 1081 3244
rect 1115 3210 1131 3244
rect 1065 3176 1131 3210
rect 1065 3142 1081 3176
rect 1115 3142 1131 3176
rect 1065 3108 1131 3142
rect 1065 3074 1081 3108
rect 1115 3074 1131 3108
rect 1065 3040 1131 3074
rect 1065 3006 1081 3040
rect 1115 3006 1131 3040
rect 1065 2989 1131 3006
rect 1161 3244 1227 3261
rect 1161 3210 1177 3244
rect 1211 3210 1227 3244
rect 1161 3176 1227 3210
rect 1161 3142 1177 3176
rect 1211 3142 1227 3176
rect 1161 3108 1227 3142
rect 1161 3074 1177 3108
rect 1211 3074 1227 3108
rect 1161 3040 1227 3074
rect 1161 3006 1177 3040
rect 1211 3006 1227 3040
rect 1161 2989 1227 3006
rect 1257 3244 1319 3261
rect 1257 3210 1273 3244
rect 1307 3210 1319 3244
rect 1257 3176 1319 3210
rect 1257 3142 1273 3176
rect 1307 3142 1319 3176
rect 1257 3108 1319 3142
rect 1257 3074 1273 3108
rect 1307 3074 1319 3108
rect 1257 3040 1319 3074
rect 1257 3006 1273 3040
rect 1307 3006 1319 3040
rect 1257 2989 1319 3006
rect 2454 3248 2516 3265
rect 2454 3214 2466 3248
rect 2500 3214 2516 3248
rect 2454 3180 2516 3214
rect 2454 3146 2466 3180
rect 2500 3146 2516 3180
rect 2454 3112 2516 3146
rect 2454 3078 2466 3112
rect 2500 3078 2516 3112
rect 2454 3044 2516 3078
rect 2454 3010 2466 3044
rect 2500 3010 2516 3044
rect 2454 2993 2516 3010
rect 2546 3248 2612 3265
rect 2546 3214 2562 3248
rect 2596 3214 2612 3248
rect 2546 3180 2612 3214
rect 2546 3146 2562 3180
rect 2596 3146 2612 3180
rect 2546 3112 2612 3146
rect 2546 3078 2562 3112
rect 2596 3078 2612 3112
rect 2546 3044 2612 3078
rect 2546 3010 2562 3044
rect 2596 3010 2612 3044
rect 2546 2993 2612 3010
rect 2642 3248 2708 3265
rect 2642 3214 2658 3248
rect 2692 3214 2708 3248
rect 2642 3180 2708 3214
rect 2642 3146 2658 3180
rect 2692 3146 2708 3180
rect 2642 3112 2708 3146
rect 2642 3078 2658 3112
rect 2692 3078 2708 3112
rect 2642 3044 2708 3078
rect 2642 3010 2658 3044
rect 2692 3010 2708 3044
rect 2642 2993 2708 3010
rect 2738 3248 2804 3265
rect 2738 3214 2754 3248
rect 2788 3214 2804 3248
rect 2738 3180 2804 3214
rect 2738 3146 2754 3180
rect 2788 3146 2804 3180
rect 2738 3112 2804 3146
rect 2738 3078 2754 3112
rect 2788 3078 2804 3112
rect 2738 3044 2804 3078
rect 2738 3010 2754 3044
rect 2788 3010 2804 3044
rect 2738 2993 2804 3010
rect 2834 3248 2900 3265
rect 2834 3214 2850 3248
rect 2884 3214 2900 3248
rect 2834 3180 2900 3214
rect 2834 3146 2850 3180
rect 2884 3146 2900 3180
rect 2834 3112 2900 3146
rect 2834 3078 2850 3112
rect 2884 3078 2900 3112
rect 2834 3044 2900 3078
rect 2834 3010 2850 3044
rect 2884 3010 2900 3044
rect 2834 2993 2900 3010
rect 2930 3248 2996 3265
rect 2930 3214 2946 3248
rect 2980 3214 2996 3248
rect 2930 3180 2996 3214
rect 2930 3146 2946 3180
rect 2980 3146 2996 3180
rect 2930 3112 2996 3146
rect 2930 3078 2946 3112
rect 2980 3078 2996 3112
rect 2930 3044 2996 3078
rect 2930 3010 2946 3044
rect 2980 3010 2996 3044
rect 2930 2993 2996 3010
rect 3026 3248 3092 3265
rect 3026 3214 3042 3248
rect 3076 3214 3092 3248
rect 3026 3180 3092 3214
rect 3026 3146 3042 3180
rect 3076 3146 3092 3180
rect 3026 3112 3092 3146
rect 3026 3078 3042 3112
rect 3076 3078 3092 3112
rect 3026 3044 3092 3078
rect 3026 3010 3042 3044
rect 3076 3010 3092 3044
rect 3026 2993 3092 3010
rect 3122 3248 3188 3265
rect 3122 3214 3138 3248
rect 3172 3214 3188 3248
rect 3122 3180 3188 3214
rect 3122 3146 3138 3180
rect 3172 3146 3188 3180
rect 3122 3112 3188 3146
rect 3122 3078 3138 3112
rect 3172 3078 3188 3112
rect 3122 3044 3188 3078
rect 3122 3010 3138 3044
rect 3172 3010 3188 3044
rect 3122 2993 3188 3010
rect 3218 3248 3284 3265
rect 3218 3214 3234 3248
rect 3268 3214 3284 3248
rect 3218 3180 3284 3214
rect 3218 3146 3234 3180
rect 3268 3146 3284 3180
rect 3218 3112 3284 3146
rect 3218 3078 3234 3112
rect 3268 3078 3284 3112
rect 3218 3044 3284 3078
rect 3218 3010 3234 3044
rect 3268 3010 3284 3044
rect 3218 2993 3284 3010
rect 3314 3248 3380 3265
rect 3314 3214 3330 3248
rect 3364 3214 3380 3248
rect 3314 3180 3380 3214
rect 3314 3146 3330 3180
rect 3364 3146 3380 3180
rect 3314 3112 3380 3146
rect 3314 3078 3330 3112
rect 3364 3078 3380 3112
rect 3314 3044 3380 3078
rect 3314 3010 3330 3044
rect 3364 3010 3380 3044
rect 3314 2993 3380 3010
rect 3410 3248 3472 3265
rect 3410 3214 3426 3248
rect 3460 3214 3472 3248
rect 3410 3180 3472 3214
rect 3410 3146 3426 3180
rect 3460 3146 3472 3180
rect 3410 3112 3472 3146
rect 3410 3078 3426 3112
rect 3460 3078 3472 3112
rect 3410 3044 3472 3078
rect 3410 3010 3426 3044
rect 3460 3010 3472 3044
rect 3410 2993 3472 3010
rect 3975 3248 4037 3265
rect 3975 3214 3987 3248
rect 4021 3214 4037 3248
rect 3975 3180 4037 3214
rect 3975 3146 3987 3180
rect 4021 3146 4037 3180
rect 3975 3112 4037 3146
rect 3975 3078 3987 3112
rect 4021 3078 4037 3112
rect 3975 3044 4037 3078
rect 3975 3010 3987 3044
rect 4021 3010 4037 3044
rect 3975 2993 4037 3010
rect 4067 3248 4133 3265
rect 4067 3214 4083 3248
rect 4117 3214 4133 3248
rect 4067 3180 4133 3214
rect 4067 3146 4083 3180
rect 4117 3146 4133 3180
rect 4067 3112 4133 3146
rect 4067 3078 4083 3112
rect 4117 3078 4133 3112
rect 4067 3044 4133 3078
rect 4067 3010 4083 3044
rect 4117 3010 4133 3044
rect 4067 2993 4133 3010
rect 4163 3248 4229 3265
rect 4163 3214 4179 3248
rect 4213 3214 4229 3248
rect 4163 3180 4229 3214
rect 4163 3146 4179 3180
rect 4213 3146 4229 3180
rect 4163 3112 4229 3146
rect 4163 3078 4179 3112
rect 4213 3078 4229 3112
rect 4163 3044 4229 3078
rect 4163 3010 4179 3044
rect 4213 3010 4229 3044
rect 4163 2993 4229 3010
rect 4259 3248 4325 3265
rect 4259 3214 4275 3248
rect 4309 3214 4325 3248
rect 4259 3180 4325 3214
rect 4259 3146 4275 3180
rect 4309 3146 4325 3180
rect 4259 3112 4325 3146
rect 4259 3078 4275 3112
rect 4309 3078 4325 3112
rect 4259 3044 4325 3078
rect 4259 3010 4275 3044
rect 4309 3010 4325 3044
rect 4259 2993 4325 3010
rect 4355 3248 4421 3265
rect 4355 3214 4371 3248
rect 4405 3214 4421 3248
rect 4355 3180 4421 3214
rect 4355 3146 4371 3180
rect 4405 3146 4421 3180
rect 4355 3112 4421 3146
rect 4355 3078 4371 3112
rect 4405 3078 4421 3112
rect 4355 3044 4421 3078
rect 4355 3010 4371 3044
rect 4405 3010 4421 3044
rect 4355 2993 4421 3010
rect 4451 3248 4517 3265
rect 4451 3214 4467 3248
rect 4501 3214 4517 3248
rect 4451 3180 4517 3214
rect 4451 3146 4467 3180
rect 4501 3146 4517 3180
rect 4451 3112 4517 3146
rect 4451 3078 4467 3112
rect 4501 3078 4517 3112
rect 4451 3044 4517 3078
rect 4451 3010 4467 3044
rect 4501 3010 4517 3044
rect 4451 2993 4517 3010
rect 4547 3248 4613 3265
rect 4547 3214 4563 3248
rect 4597 3214 4613 3248
rect 4547 3180 4613 3214
rect 4547 3146 4563 3180
rect 4597 3146 4613 3180
rect 4547 3112 4613 3146
rect 4547 3078 4563 3112
rect 4597 3078 4613 3112
rect 4547 3044 4613 3078
rect 4547 3010 4563 3044
rect 4597 3010 4613 3044
rect 4547 2993 4613 3010
rect 4643 3248 4709 3265
rect 4643 3214 4659 3248
rect 4693 3214 4709 3248
rect 4643 3180 4709 3214
rect 4643 3146 4659 3180
rect 4693 3146 4709 3180
rect 4643 3112 4709 3146
rect 4643 3078 4659 3112
rect 4693 3078 4709 3112
rect 4643 3044 4709 3078
rect 4643 3010 4659 3044
rect 4693 3010 4709 3044
rect 4643 2993 4709 3010
rect 4739 3248 4805 3265
rect 4739 3214 4755 3248
rect 4789 3214 4805 3248
rect 4739 3180 4805 3214
rect 4739 3146 4755 3180
rect 4789 3146 4805 3180
rect 4739 3112 4805 3146
rect 4739 3078 4755 3112
rect 4789 3078 4805 3112
rect 4739 3044 4805 3078
rect 4739 3010 4755 3044
rect 4789 3010 4805 3044
rect 4739 2993 4805 3010
rect 4835 3248 4901 3265
rect 4835 3214 4851 3248
rect 4885 3214 4901 3248
rect 4835 3180 4901 3214
rect 4835 3146 4851 3180
rect 4885 3146 4901 3180
rect 4835 3112 4901 3146
rect 4835 3078 4851 3112
rect 4885 3078 4901 3112
rect 4835 3044 4901 3078
rect 4835 3010 4851 3044
rect 4885 3010 4901 3044
rect 4835 2993 4901 3010
rect 4931 3248 4993 3265
rect 4931 3214 4947 3248
rect 4981 3214 4993 3248
rect 4931 3180 4993 3214
rect 4931 3146 4947 3180
rect 4981 3146 4993 3180
rect 4931 3112 4993 3146
rect 4931 3078 4947 3112
rect 4981 3078 4993 3112
rect 4931 3044 4993 3078
rect 4931 3010 4947 3044
rect 4981 3010 4993 3044
rect 4931 2993 4993 3010
rect 5348 3040 5400 3052
rect 5348 3006 5356 3040
rect 5390 3006 5400 3040
rect 5348 2972 5400 3006
rect 5348 2938 5356 2972
rect 5390 2938 5400 2972
rect 5348 2904 5400 2938
rect 5348 2870 5356 2904
rect 5390 2870 5400 2904
rect 5348 2852 5400 2870
rect 5430 3040 5482 3052
rect 5430 3006 5440 3040
rect 5474 3006 5482 3040
rect 5430 2972 5482 3006
rect 5430 2938 5440 2972
rect 5474 2938 5482 2972
rect 5430 2904 5482 2938
rect 5430 2870 5440 2904
rect 5474 2870 5482 2904
rect 5430 2852 5482 2870
rect 301 1957 363 1974
rect 301 1923 313 1957
rect 347 1923 363 1957
rect 301 1889 363 1923
rect 301 1855 313 1889
rect 347 1855 363 1889
rect 301 1821 363 1855
rect 301 1787 313 1821
rect 347 1787 363 1821
rect 301 1753 363 1787
rect 301 1719 313 1753
rect 347 1719 363 1753
rect 301 1702 363 1719
rect 393 1957 459 1974
rect 393 1923 409 1957
rect 443 1923 459 1957
rect 393 1889 459 1923
rect 393 1855 409 1889
rect 443 1855 459 1889
rect 393 1821 459 1855
rect 393 1787 409 1821
rect 443 1787 459 1821
rect 393 1753 459 1787
rect 393 1719 409 1753
rect 443 1719 459 1753
rect 393 1702 459 1719
rect 489 1957 555 1974
rect 489 1923 505 1957
rect 539 1923 555 1957
rect 489 1889 555 1923
rect 489 1855 505 1889
rect 539 1855 555 1889
rect 489 1821 555 1855
rect 489 1787 505 1821
rect 539 1787 555 1821
rect 489 1753 555 1787
rect 489 1719 505 1753
rect 539 1719 555 1753
rect 489 1702 555 1719
rect 585 1957 651 1974
rect 585 1923 601 1957
rect 635 1923 651 1957
rect 585 1889 651 1923
rect 585 1855 601 1889
rect 635 1855 651 1889
rect 585 1821 651 1855
rect 585 1787 601 1821
rect 635 1787 651 1821
rect 585 1753 651 1787
rect 585 1719 601 1753
rect 635 1719 651 1753
rect 585 1702 651 1719
rect 681 1957 747 1974
rect 681 1923 697 1957
rect 731 1923 747 1957
rect 681 1889 747 1923
rect 681 1855 697 1889
rect 731 1855 747 1889
rect 681 1821 747 1855
rect 681 1787 697 1821
rect 731 1787 747 1821
rect 681 1753 747 1787
rect 681 1719 697 1753
rect 731 1719 747 1753
rect 681 1702 747 1719
rect 777 1957 843 1974
rect 777 1923 793 1957
rect 827 1923 843 1957
rect 777 1889 843 1923
rect 777 1855 793 1889
rect 827 1855 843 1889
rect 777 1821 843 1855
rect 777 1787 793 1821
rect 827 1787 843 1821
rect 777 1753 843 1787
rect 777 1719 793 1753
rect 827 1719 843 1753
rect 777 1702 843 1719
rect 873 1957 939 1974
rect 873 1923 889 1957
rect 923 1923 939 1957
rect 873 1889 939 1923
rect 873 1855 889 1889
rect 923 1855 939 1889
rect 873 1821 939 1855
rect 873 1787 889 1821
rect 923 1787 939 1821
rect 873 1753 939 1787
rect 873 1719 889 1753
rect 923 1719 939 1753
rect 873 1702 939 1719
rect 969 1957 1035 1974
rect 969 1923 985 1957
rect 1019 1923 1035 1957
rect 969 1889 1035 1923
rect 969 1855 985 1889
rect 1019 1855 1035 1889
rect 969 1821 1035 1855
rect 969 1787 985 1821
rect 1019 1787 1035 1821
rect 969 1753 1035 1787
rect 969 1719 985 1753
rect 1019 1719 1035 1753
rect 969 1702 1035 1719
rect 1065 1957 1131 1974
rect 1065 1923 1081 1957
rect 1115 1923 1131 1957
rect 1065 1889 1131 1923
rect 1065 1855 1081 1889
rect 1115 1855 1131 1889
rect 1065 1821 1131 1855
rect 1065 1787 1081 1821
rect 1115 1787 1131 1821
rect 1065 1753 1131 1787
rect 1065 1719 1081 1753
rect 1115 1719 1131 1753
rect 1065 1702 1131 1719
rect 1161 1957 1227 1974
rect 1161 1923 1177 1957
rect 1211 1923 1227 1957
rect 1161 1889 1227 1923
rect 1161 1855 1177 1889
rect 1211 1855 1227 1889
rect 1161 1821 1227 1855
rect 1161 1787 1177 1821
rect 1211 1787 1227 1821
rect 1161 1753 1227 1787
rect 1161 1719 1177 1753
rect 1211 1719 1227 1753
rect 1161 1702 1227 1719
rect 1257 1957 1319 1974
rect 1257 1923 1273 1957
rect 1307 1923 1319 1957
rect 1257 1889 1319 1923
rect 1257 1855 1273 1889
rect 1307 1855 1319 1889
rect 1257 1821 1319 1855
rect 1257 1787 1273 1821
rect 1307 1787 1319 1821
rect 1257 1753 1319 1787
rect 1257 1719 1273 1753
rect 1307 1719 1319 1753
rect 1257 1702 1319 1719
rect 2454 1961 2516 1978
rect 2454 1927 2466 1961
rect 2500 1927 2516 1961
rect 2454 1893 2516 1927
rect 2454 1859 2466 1893
rect 2500 1859 2516 1893
rect 2454 1825 2516 1859
rect 2454 1791 2466 1825
rect 2500 1791 2516 1825
rect 2454 1757 2516 1791
rect 2454 1723 2466 1757
rect 2500 1723 2516 1757
rect 2454 1706 2516 1723
rect 2546 1961 2612 1978
rect 2546 1927 2562 1961
rect 2596 1927 2612 1961
rect 2546 1893 2612 1927
rect 2546 1859 2562 1893
rect 2596 1859 2612 1893
rect 2546 1825 2612 1859
rect 2546 1791 2562 1825
rect 2596 1791 2612 1825
rect 2546 1757 2612 1791
rect 2546 1723 2562 1757
rect 2596 1723 2612 1757
rect 2546 1706 2612 1723
rect 2642 1961 2708 1978
rect 2642 1927 2658 1961
rect 2692 1927 2708 1961
rect 2642 1893 2708 1927
rect 2642 1859 2658 1893
rect 2692 1859 2708 1893
rect 2642 1825 2708 1859
rect 2642 1791 2658 1825
rect 2692 1791 2708 1825
rect 2642 1757 2708 1791
rect 2642 1723 2658 1757
rect 2692 1723 2708 1757
rect 2642 1706 2708 1723
rect 2738 1961 2804 1978
rect 2738 1927 2754 1961
rect 2788 1927 2804 1961
rect 2738 1893 2804 1927
rect 2738 1859 2754 1893
rect 2788 1859 2804 1893
rect 2738 1825 2804 1859
rect 2738 1791 2754 1825
rect 2788 1791 2804 1825
rect 2738 1757 2804 1791
rect 2738 1723 2754 1757
rect 2788 1723 2804 1757
rect 2738 1706 2804 1723
rect 2834 1961 2900 1978
rect 2834 1927 2850 1961
rect 2884 1927 2900 1961
rect 2834 1893 2900 1927
rect 2834 1859 2850 1893
rect 2884 1859 2900 1893
rect 2834 1825 2900 1859
rect 2834 1791 2850 1825
rect 2884 1791 2900 1825
rect 2834 1757 2900 1791
rect 2834 1723 2850 1757
rect 2884 1723 2900 1757
rect 2834 1706 2900 1723
rect 2930 1961 2996 1978
rect 2930 1927 2946 1961
rect 2980 1927 2996 1961
rect 2930 1893 2996 1927
rect 2930 1859 2946 1893
rect 2980 1859 2996 1893
rect 2930 1825 2996 1859
rect 2930 1791 2946 1825
rect 2980 1791 2996 1825
rect 2930 1757 2996 1791
rect 2930 1723 2946 1757
rect 2980 1723 2996 1757
rect 2930 1706 2996 1723
rect 3026 1961 3092 1978
rect 3026 1927 3042 1961
rect 3076 1927 3092 1961
rect 3026 1893 3092 1927
rect 3026 1859 3042 1893
rect 3076 1859 3092 1893
rect 3026 1825 3092 1859
rect 3026 1791 3042 1825
rect 3076 1791 3092 1825
rect 3026 1757 3092 1791
rect 3026 1723 3042 1757
rect 3076 1723 3092 1757
rect 3026 1706 3092 1723
rect 3122 1961 3188 1978
rect 3122 1927 3138 1961
rect 3172 1927 3188 1961
rect 3122 1893 3188 1927
rect 3122 1859 3138 1893
rect 3172 1859 3188 1893
rect 3122 1825 3188 1859
rect 3122 1791 3138 1825
rect 3172 1791 3188 1825
rect 3122 1757 3188 1791
rect 3122 1723 3138 1757
rect 3172 1723 3188 1757
rect 3122 1706 3188 1723
rect 3218 1961 3284 1978
rect 3218 1927 3234 1961
rect 3268 1927 3284 1961
rect 3218 1893 3284 1927
rect 3218 1859 3234 1893
rect 3268 1859 3284 1893
rect 3218 1825 3284 1859
rect 3218 1791 3234 1825
rect 3268 1791 3284 1825
rect 3218 1757 3284 1791
rect 3218 1723 3234 1757
rect 3268 1723 3284 1757
rect 3218 1706 3284 1723
rect 3314 1961 3380 1978
rect 3314 1927 3330 1961
rect 3364 1927 3380 1961
rect 3314 1893 3380 1927
rect 3314 1859 3330 1893
rect 3364 1859 3380 1893
rect 3314 1825 3380 1859
rect 3314 1791 3330 1825
rect 3364 1791 3380 1825
rect 3314 1757 3380 1791
rect 3314 1723 3330 1757
rect 3364 1723 3380 1757
rect 3314 1706 3380 1723
rect 3410 1961 3472 1978
rect 3410 1927 3426 1961
rect 3460 1927 3472 1961
rect 3410 1893 3472 1927
rect 3410 1859 3426 1893
rect 3460 1859 3472 1893
rect 3410 1825 3472 1859
rect 3410 1791 3426 1825
rect 3460 1791 3472 1825
rect 3410 1757 3472 1791
rect 3410 1723 3426 1757
rect 3460 1723 3472 1757
rect 3410 1706 3472 1723
rect 3975 1961 4037 1978
rect 3975 1927 3987 1961
rect 4021 1927 4037 1961
rect 3975 1893 4037 1927
rect 3975 1859 3987 1893
rect 4021 1859 4037 1893
rect 3975 1825 4037 1859
rect 3975 1791 3987 1825
rect 4021 1791 4037 1825
rect 3975 1757 4037 1791
rect 3975 1723 3987 1757
rect 4021 1723 4037 1757
rect 3975 1706 4037 1723
rect 4067 1961 4133 1978
rect 4067 1927 4083 1961
rect 4117 1927 4133 1961
rect 4067 1893 4133 1927
rect 4067 1859 4083 1893
rect 4117 1859 4133 1893
rect 4067 1825 4133 1859
rect 4067 1791 4083 1825
rect 4117 1791 4133 1825
rect 4067 1757 4133 1791
rect 4067 1723 4083 1757
rect 4117 1723 4133 1757
rect 4067 1706 4133 1723
rect 4163 1961 4229 1978
rect 4163 1927 4179 1961
rect 4213 1927 4229 1961
rect 4163 1893 4229 1927
rect 4163 1859 4179 1893
rect 4213 1859 4229 1893
rect 4163 1825 4229 1859
rect 4163 1791 4179 1825
rect 4213 1791 4229 1825
rect 4163 1757 4229 1791
rect 4163 1723 4179 1757
rect 4213 1723 4229 1757
rect 4163 1706 4229 1723
rect 4259 1961 4325 1978
rect 4259 1927 4275 1961
rect 4309 1927 4325 1961
rect 4259 1893 4325 1927
rect 4259 1859 4275 1893
rect 4309 1859 4325 1893
rect 4259 1825 4325 1859
rect 4259 1791 4275 1825
rect 4309 1791 4325 1825
rect 4259 1757 4325 1791
rect 4259 1723 4275 1757
rect 4309 1723 4325 1757
rect 4259 1706 4325 1723
rect 4355 1961 4421 1978
rect 4355 1927 4371 1961
rect 4405 1927 4421 1961
rect 4355 1893 4421 1927
rect 4355 1859 4371 1893
rect 4405 1859 4421 1893
rect 4355 1825 4421 1859
rect 4355 1791 4371 1825
rect 4405 1791 4421 1825
rect 4355 1757 4421 1791
rect 4355 1723 4371 1757
rect 4405 1723 4421 1757
rect 4355 1706 4421 1723
rect 4451 1961 4517 1978
rect 4451 1927 4467 1961
rect 4501 1927 4517 1961
rect 4451 1893 4517 1927
rect 4451 1859 4467 1893
rect 4501 1859 4517 1893
rect 4451 1825 4517 1859
rect 4451 1791 4467 1825
rect 4501 1791 4517 1825
rect 4451 1757 4517 1791
rect 4451 1723 4467 1757
rect 4501 1723 4517 1757
rect 4451 1706 4517 1723
rect 4547 1961 4613 1978
rect 4547 1927 4563 1961
rect 4597 1927 4613 1961
rect 4547 1893 4613 1927
rect 4547 1859 4563 1893
rect 4597 1859 4613 1893
rect 4547 1825 4613 1859
rect 4547 1791 4563 1825
rect 4597 1791 4613 1825
rect 4547 1757 4613 1791
rect 4547 1723 4563 1757
rect 4597 1723 4613 1757
rect 4547 1706 4613 1723
rect 4643 1961 4709 1978
rect 4643 1927 4659 1961
rect 4693 1927 4709 1961
rect 4643 1893 4709 1927
rect 4643 1859 4659 1893
rect 4693 1859 4709 1893
rect 4643 1825 4709 1859
rect 4643 1791 4659 1825
rect 4693 1791 4709 1825
rect 4643 1757 4709 1791
rect 4643 1723 4659 1757
rect 4693 1723 4709 1757
rect 4643 1706 4709 1723
rect 4739 1961 4805 1978
rect 4739 1927 4755 1961
rect 4789 1927 4805 1961
rect 4739 1893 4805 1927
rect 4739 1859 4755 1893
rect 4789 1859 4805 1893
rect 4739 1825 4805 1859
rect 4739 1791 4755 1825
rect 4789 1791 4805 1825
rect 4739 1757 4805 1791
rect 4739 1723 4755 1757
rect 4789 1723 4805 1757
rect 4739 1706 4805 1723
rect 4835 1961 4901 1978
rect 4835 1927 4851 1961
rect 4885 1927 4901 1961
rect 4835 1893 4901 1927
rect 4835 1859 4851 1893
rect 4885 1859 4901 1893
rect 4835 1825 4901 1859
rect 4835 1791 4851 1825
rect 4885 1791 4901 1825
rect 4835 1757 4901 1791
rect 4835 1723 4851 1757
rect 4885 1723 4901 1757
rect 4835 1706 4901 1723
rect 4931 1961 4993 1978
rect 4931 1927 4947 1961
rect 4981 1927 4993 1961
rect 4931 1893 4993 1927
rect 4931 1859 4947 1893
rect 4981 1859 4993 1893
rect 4931 1825 4993 1859
rect 4931 1791 4947 1825
rect 4981 1791 4993 1825
rect 4931 1757 4993 1791
rect 4931 1723 4947 1757
rect 4981 1723 4993 1757
rect 4931 1706 4993 1723
rect 5348 1753 5400 1765
rect 5348 1719 5356 1753
rect 5390 1719 5400 1753
rect 5348 1685 5400 1719
rect 5348 1651 5356 1685
rect 5390 1651 5400 1685
rect 5348 1617 5400 1651
rect 5348 1583 5356 1617
rect 5390 1583 5400 1617
rect 5348 1565 5400 1583
rect 5430 1753 5482 1765
rect 5430 1719 5440 1753
rect 5474 1719 5482 1753
rect 5430 1685 5482 1719
rect 5430 1651 5440 1685
rect 5474 1651 5482 1685
rect 5430 1617 5482 1651
rect 5430 1583 5440 1617
rect 5474 1583 5482 1617
rect 5430 1565 5482 1583
<< ndiffc >>
rect 313 41222 347 41256
rect 409 41222 443 41256
rect 505 41222 539 41256
rect 601 41222 635 41256
rect 697 41222 731 41256
rect 793 41222 827 41256
rect 889 41222 923 41256
rect 985 41222 1019 41256
rect 1081 41222 1115 41256
rect 1177 41222 1211 41256
rect 1273 41222 1307 41256
rect 2466 41226 2500 41260
rect 2562 41226 2596 41260
rect 2658 41226 2692 41260
rect 2754 41226 2788 41260
rect 2850 41226 2884 41260
rect 2946 41226 2980 41260
rect 3042 41226 3076 41260
rect 3138 41226 3172 41260
rect 3234 41226 3268 41260
rect 3330 41226 3364 41260
rect 3426 41226 3460 41260
rect 3647 41211 3681 41287
rect 3735 41211 3769 41287
rect 3987 41226 4021 41260
rect 4083 41226 4117 41260
rect 4179 41226 4213 41260
rect 4275 41226 4309 41260
rect 4371 41226 4405 41260
rect 4467 41226 4501 41260
rect 4563 41226 4597 41260
rect 4659 41226 4693 41260
rect 4755 41226 4789 41260
rect 4851 41226 4885 41260
rect 4947 41226 4981 41260
rect 5356 41296 5390 41330
rect 5356 41228 5390 41262
rect 5440 41296 5474 41330
rect 5440 41228 5474 41262
rect 313 39935 347 39969
rect 409 39935 443 39969
rect 505 39935 539 39969
rect 601 39935 635 39969
rect 697 39935 731 39969
rect 793 39935 827 39969
rect 889 39935 923 39969
rect 985 39935 1019 39969
rect 1081 39935 1115 39969
rect 1177 39935 1211 39969
rect 1273 39935 1307 39969
rect 2466 39939 2500 39973
rect 2562 39939 2596 39973
rect 2658 39939 2692 39973
rect 2754 39939 2788 39973
rect 2850 39939 2884 39973
rect 2946 39939 2980 39973
rect 3042 39939 3076 39973
rect 3138 39939 3172 39973
rect 3234 39939 3268 39973
rect 3330 39939 3364 39973
rect 3426 39939 3460 39973
rect 3647 39924 3681 40000
rect 3735 39924 3769 40000
rect 3987 39939 4021 39973
rect 4083 39939 4117 39973
rect 4179 39939 4213 39973
rect 4275 39939 4309 39973
rect 4371 39939 4405 39973
rect 4467 39939 4501 39973
rect 4563 39939 4597 39973
rect 4659 39939 4693 39973
rect 4755 39939 4789 39973
rect 4851 39939 4885 39973
rect 4947 39939 4981 39973
rect 5356 40009 5390 40043
rect 5356 39941 5390 39975
rect 5440 40009 5474 40043
rect 5440 39941 5474 39975
rect 313 38648 347 38682
rect 409 38648 443 38682
rect 505 38648 539 38682
rect 601 38648 635 38682
rect 697 38648 731 38682
rect 793 38648 827 38682
rect 889 38648 923 38682
rect 985 38648 1019 38682
rect 1081 38648 1115 38682
rect 1177 38648 1211 38682
rect 1273 38648 1307 38682
rect 2466 38652 2500 38686
rect 2562 38652 2596 38686
rect 2658 38652 2692 38686
rect 2754 38652 2788 38686
rect 2850 38652 2884 38686
rect 2946 38652 2980 38686
rect 3042 38652 3076 38686
rect 3138 38652 3172 38686
rect 3234 38652 3268 38686
rect 3330 38652 3364 38686
rect 3426 38652 3460 38686
rect 3647 38637 3681 38713
rect 3735 38637 3769 38713
rect 3987 38652 4021 38686
rect 4083 38652 4117 38686
rect 4179 38652 4213 38686
rect 4275 38652 4309 38686
rect 4371 38652 4405 38686
rect 4467 38652 4501 38686
rect 4563 38652 4597 38686
rect 4659 38652 4693 38686
rect 4755 38652 4789 38686
rect 4851 38652 4885 38686
rect 4947 38652 4981 38686
rect 5356 38722 5390 38756
rect 5356 38654 5390 38688
rect 5440 38722 5474 38756
rect 5440 38654 5474 38688
rect 313 37361 347 37395
rect 409 37361 443 37395
rect 505 37361 539 37395
rect 601 37361 635 37395
rect 697 37361 731 37395
rect 793 37361 827 37395
rect 889 37361 923 37395
rect 985 37361 1019 37395
rect 1081 37361 1115 37395
rect 1177 37361 1211 37395
rect 1273 37361 1307 37395
rect 2466 37365 2500 37399
rect 2562 37365 2596 37399
rect 2658 37365 2692 37399
rect 2754 37365 2788 37399
rect 2850 37365 2884 37399
rect 2946 37365 2980 37399
rect 3042 37365 3076 37399
rect 3138 37365 3172 37399
rect 3234 37365 3268 37399
rect 3330 37365 3364 37399
rect 3426 37365 3460 37399
rect 3647 37350 3681 37426
rect 3735 37350 3769 37426
rect 3987 37365 4021 37399
rect 4083 37365 4117 37399
rect 4179 37365 4213 37399
rect 4275 37365 4309 37399
rect 4371 37365 4405 37399
rect 4467 37365 4501 37399
rect 4563 37365 4597 37399
rect 4659 37365 4693 37399
rect 4755 37365 4789 37399
rect 4851 37365 4885 37399
rect 4947 37365 4981 37399
rect 5356 37435 5390 37469
rect 5356 37367 5390 37401
rect 5440 37435 5474 37469
rect 5440 37367 5474 37401
rect 313 36074 347 36108
rect 409 36074 443 36108
rect 505 36074 539 36108
rect 601 36074 635 36108
rect 697 36074 731 36108
rect 793 36074 827 36108
rect 889 36074 923 36108
rect 985 36074 1019 36108
rect 1081 36074 1115 36108
rect 1177 36074 1211 36108
rect 1273 36074 1307 36108
rect 2466 36078 2500 36112
rect 2562 36078 2596 36112
rect 2658 36078 2692 36112
rect 2754 36078 2788 36112
rect 2850 36078 2884 36112
rect 2946 36078 2980 36112
rect 3042 36078 3076 36112
rect 3138 36078 3172 36112
rect 3234 36078 3268 36112
rect 3330 36078 3364 36112
rect 3426 36078 3460 36112
rect 3647 36063 3681 36139
rect 3735 36063 3769 36139
rect 3987 36078 4021 36112
rect 4083 36078 4117 36112
rect 4179 36078 4213 36112
rect 4275 36078 4309 36112
rect 4371 36078 4405 36112
rect 4467 36078 4501 36112
rect 4563 36078 4597 36112
rect 4659 36078 4693 36112
rect 4755 36078 4789 36112
rect 4851 36078 4885 36112
rect 4947 36078 4981 36112
rect 5356 36148 5390 36182
rect 5356 36080 5390 36114
rect 5440 36148 5474 36182
rect 5440 36080 5474 36114
rect 313 34787 347 34821
rect 409 34787 443 34821
rect 505 34787 539 34821
rect 601 34787 635 34821
rect 697 34787 731 34821
rect 793 34787 827 34821
rect 889 34787 923 34821
rect 985 34787 1019 34821
rect 1081 34787 1115 34821
rect 1177 34787 1211 34821
rect 1273 34787 1307 34821
rect 2466 34791 2500 34825
rect 2562 34791 2596 34825
rect 2658 34791 2692 34825
rect 2754 34791 2788 34825
rect 2850 34791 2884 34825
rect 2946 34791 2980 34825
rect 3042 34791 3076 34825
rect 3138 34791 3172 34825
rect 3234 34791 3268 34825
rect 3330 34791 3364 34825
rect 3426 34791 3460 34825
rect 3647 34776 3681 34852
rect 3735 34776 3769 34852
rect 3987 34791 4021 34825
rect 4083 34791 4117 34825
rect 4179 34791 4213 34825
rect 4275 34791 4309 34825
rect 4371 34791 4405 34825
rect 4467 34791 4501 34825
rect 4563 34791 4597 34825
rect 4659 34791 4693 34825
rect 4755 34791 4789 34825
rect 4851 34791 4885 34825
rect 4947 34791 4981 34825
rect 5356 34861 5390 34895
rect 5356 34793 5390 34827
rect 5440 34861 5474 34895
rect 5440 34793 5474 34827
rect 313 33500 347 33534
rect 409 33500 443 33534
rect 505 33500 539 33534
rect 601 33500 635 33534
rect 697 33500 731 33534
rect 793 33500 827 33534
rect 889 33500 923 33534
rect 985 33500 1019 33534
rect 1081 33500 1115 33534
rect 1177 33500 1211 33534
rect 1273 33500 1307 33534
rect 2466 33504 2500 33538
rect 2562 33504 2596 33538
rect 2658 33504 2692 33538
rect 2754 33504 2788 33538
rect 2850 33504 2884 33538
rect 2946 33504 2980 33538
rect 3042 33504 3076 33538
rect 3138 33504 3172 33538
rect 3234 33504 3268 33538
rect 3330 33504 3364 33538
rect 3426 33504 3460 33538
rect 3647 33489 3681 33565
rect 3735 33489 3769 33565
rect 3987 33504 4021 33538
rect 4083 33504 4117 33538
rect 4179 33504 4213 33538
rect 4275 33504 4309 33538
rect 4371 33504 4405 33538
rect 4467 33504 4501 33538
rect 4563 33504 4597 33538
rect 4659 33504 4693 33538
rect 4755 33504 4789 33538
rect 4851 33504 4885 33538
rect 4947 33504 4981 33538
rect 5356 33574 5390 33608
rect 5356 33506 5390 33540
rect 5440 33574 5474 33608
rect 5440 33506 5474 33540
rect 313 32213 347 32247
rect 409 32213 443 32247
rect 505 32213 539 32247
rect 601 32213 635 32247
rect 697 32213 731 32247
rect 793 32213 827 32247
rect 889 32213 923 32247
rect 985 32213 1019 32247
rect 1081 32213 1115 32247
rect 1177 32213 1211 32247
rect 1273 32213 1307 32247
rect 2466 32217 2500 32251
rect 2562 32217 2596 32251
rect 2658 32217 2692 32251
rect 2754 32217 2788 32251
rect 2850 32217 2884 32251
rect 2946 32217 2980 32251
rect 3042 32217 3076 32251
rect 3138 32217 3172 32251
rect 3234 32217 3268 32251
rect 3330 32217 3364 32251
rect 3426 32217 3460 32251
rect 3647 32202 3681 32278
rect 3735 32202 3769 32278
rect 3987 32217 4021 32251
rect 4083 32217 4117 32251
rect 4179 32217 4213 32251
rect 4275 32217 4309 32251
rect 4371 32217 4405 32251
rect 4467 32217 4501 32251
rect 4563 32217 4597 32251
rect 4659 32217 4693 32251
rect 4755 32217 4789 32251
rect 4851 32217 4885 32251
rect 4947 32217 4981 32251
rect 5356 32287 5390 32321
rect 5356 32219 5390 32253
rect 5440 32287 5474 32321
rect 5440 32219 5474 32253
rect 313 30926 347 30960
rect 409 30926 443 30960
rect 505 30926 539 30960
rect 601 30926 635 30960
rect 697 30926 731 30960
rect 793 30926 827 30960
rect 889 30926 923 30960
rect 985 30926 1019 30960
rect 1081 30926 1115 30960
rect 1177 30926 1211 30960
rect 1273 30926 1307 30960
rect 2466 30930 2500 30964
rect 2562 30930 2596 30964
rect 2658 30930 2692 30964
rect 2754 30930 2788 30964
rect 2850 30930 2884 30964
rect 2946 30930 2980 30964
rect 3042 30930 3076 30964
rect 3138 30930 3172 30964
rect 3234 30930 3268 30964
rect 3330 30930 3364 30964
rect 3426 30930 3460 30964
rect 3647 30915 3681 30991
rect 3735 30915 3769 30991
rect 3987 30930 4021 30964
rect 4083 30930 4117 30964
rect 4179 30930 4213 30964
rect 4275 30930 4309 30964
rect 4371 30930 4405 30964
rect 4467 30930 4501 30964
rect 4563 30930 4597 30964
rect 4659 30930 4693 30964
rect 4755 30930 4789 30964
rect 4851 30930 4885 30964
rect 4947 30930 4981 30964
rect 5356 31000 5390 31034
rect 5356 30932 5390 30966
rect 5440 31000 5474 31034
rect 5440 30932 5474 30966
rect 313 29639 347 29673
rect 409 29639 443 29673
rect 505 29639 539 29673
rect 601 29639 635 29673
rect 697 29639 731 29673
rect 793 29639 827 29673
rect 889 29639 923 29673
rect 985 29639 1019 29673
rect 1081 29639 1115 29673
rect 1177 29639 1211 29673
rect 1273 29639 1307 29673
rect 2466 29643 2500 29677
rect 2562 29643 2596 29677
rect 2658 29643 2692 29677
rect 2754 29643 2788 29677
rect 2850 29643 2884 29677
rect 2946 29643 2980 29677
rect 3042 29643 3076 29677
rect 3138 29643 3172 29677
rect 3234 29643 3268 29677
rect 3330 29643 3364 29677
rect 3426 29643 3460 29677
rect 3647 29628 3681 29704
rect 3735 29628 3769 29704
rect 3987 29643 4021 29677
rect 4083 29643 4117 29677
rect 4179 29643 4213 29677
rect 4275 29643 4309 29677
rect 4371 29643 4405 29677
rect 4467 29643 4501 29677
rect 4563 29643 4597 29677
rect 4659 29643 4693 29677
rect 4755 29643 4789 29677
rect 4851 29643 4885 29677
rect 4947 29643 4981 29677
rect 5356 29713 5390 29747
rect 5356 29645 5390 29679
rect 5440 29713 5474 29747
rect 5440 29645 5474 29679
rect 313 28352 347 28386
rect 409 28352 443 28386
rect 505 28352 539 28386
rect 601 28352 635 28386
rect 697 28352 731 28386
rect 793 28352 827 28386
rect 889 28352 923 28386
rect 985 28352 1019 28386
rect 1081 28352 1115 28386
rect 1177 28352 1211 28386
rect 1273 28352 1307 28386
rect 2466 28356 2500 28390
rect 2562 28356 2596 28390
rect 2658 28356 2692 28390
rect 2754 28356 2788 28390
rect 2850 28356 2884 28390
rect 2946 28356 2980 28390
rect 3042 28356 3076 28390
rect 3138 28356 3172 28390
rect 3234 28356 3268 28390
rect 3330 28356 3364 28390
rect 3426 28356 3460 28390
rect 3647 28341 3681 28417
rect 3735 28341 3769 28417
rect 3987 28356 4021 28390
rect 4083 28356 4117 28390
rect 4179 28356 4213 28390
rect 4275 28356 4309 28390
rect 4371 28356 4405 28390
rect 4467 28356 4501 28390
rect 4563 28356 4597 28390
rect 4659 28356 4693 28390
rect 4755 28356 4789 28390
rect 4851 28356 4885 28390
rect 4947 28356 4981 28390
rect 5356 28426 5390 28460
rect 5356 28358 5390 28392
rect 5440 28426 5474 28460
rect 5440 28358 5474 28392
rect 313 27065 347 27099
rect 409 27065 443 27099
rect 505 27065 539 27099
rect 601 27065 635 27099
rect 697 27065 731 27099
rect 793 27065 827 27099
rect 889 27065 923 27099
rect 985 27065 1019 27099
rect 1081 27065 1115 27099
rect 1177 27065 1211 27099
rect 1273 27065 1307 27099
rect 2466 27069 2500 27103
rect 2562 27069 2596 27103
rect 2658 27069 2692 27103
rect 2754 27069 2788 27103
rect 2850 27069 2884 27103
rect 2946 27069 2980 27103
rect 3042 27069 3076 27103
rect 3138 27069 3172 27103
rect 3234 27069 3268 27103
rect 3330 27069 3364 27103
rect 3426 27069 3460 27103
rect 3647 27054 3681 27130
rect 3735 27054 3769 27130
rect 3987 27069 4021 27103
rect 4083 27069 4117 27103
rect 4179 27069 4213 27103
rect 4275 27069 4309 27103
rect 4371 27069 4405 27103
rect 4467 27069 4501 27103
rect 4563 27069 4597 27103
rect 4659 27069 4693 27103
rect 4755 27069 4789 27103
rect 4851 27069 4885 27103
rect 4947 27069 4981 27103
rect 5356 27139 5390 27173
rect 5356 27071 5390 27105
rect 5440 27139 5474 27173
rect 5440 27071 5474 27105
rect 313 25778 347 25812
rect 409 25778 443 25812
rect 505 25778 539 25812
rect 601 25778 635 25812
rect 697 25778 731 25812
rect 793 25778 827 25812
rect 889 25778 923 25812
rect 985 25778 1019 25812
rect 1081 25778 1115 25812
rect 1177 25778 1211 25812
rect 1273 25778 1307 25812
rect 2466 25782 2500 25816
rect 2562 25782 2596 25816
rect 2658 25782 2692 25816
rect 2754 25782 2788 25816
rect 2850 25782 2884 25816
rect 2946 25782 2980 25816
rect 3042 25782 3076 25816
rect 3138 25782 3172 25816
rect 3234 25782 3268 25816
rect 3330 25782 3364 25816
rect 3426 25782 3460 25816
rect 3647 25767 3681 25843
rect 3735 25767 3769 25843
rect 3987 25782 4021 25816
rect 4083 25782 4117 25816
rect 4179 25782 4213 25816
rect 4275 25782 4309 25816
rect 4371 25782 4405 25816
rect 4467 25782 4501 25816
rect 4563 25782 4597 25816
rect 4659 25782 4693 25816
rect 4755 25782 4789 25816
rect 4851 25782 4885 25816
rect 4947 25782 4981 25816
rect 5356 25852 5390 25886
rect 5356 25784 5390 25818
rect 5440 25852 5474 25886
rect 5440 25784 5474 25818
rect 313 24491 347 24525
rect 409 24491 443 24525
rect 505 24491 539 24525
rect 601 24491 635 24525
rect 697 24491 731 24525
rect 793 24491 827 24525
rect 889 24491 923 24525
rect 985 24491 1019 24525
rect 1081 24491 1115 24525
rect 1177 24491 1211 24525
rect 1273 24491 1307 24525
rect 2466 24495 2500 24529
rect 2562 24495 2596 24529
rect 2658 24495 2692 24529
rect 2754 24495 2788 24529
rect 2850 24495 2884 24529
rect 2946 24495 2980 24529
rect 3042 24495 3076 24529
rect 3138 24495 3172 24529
rect 3234 24495 3268 24529
rect 3330 24495 3364 24529
rect 3426 24495 3460 24529
rect 3647 24480 3681 24556
rect 3735 24480 3769 24556
rect 3987 24495 4021 24529
rect 4083 24495 4117 24529
rect 4179 24495 4213 24529
rect 4275 24495 4309 24529
rect 4371 24495 4405 24529
rect 4467 24495 4501 24529
rect 4563 24495 4597 24529
rect 4659 24495 4693 24529
rect 4755 24495 4789 24529
rect 4851 24495 4885 24529
rect 4947 24495 4981 24529
rect 5356 24565 5390 24599
rect 5356 24497 5390 24531
rect 5440 24565 5474 24599
rect 5440 24497 5474 24531
rect 313 23204 347 23238
rect 409 23204 443 23238
rect 505 23204 539 23238
rect 601 23204 635 23238
rect 697 23204 731 23238
rect 793 23204 827 23238
rect 889 23204 923 23238
rect 985 23204 1019 23238
rect 1081 23204 1115 23238
rect 1177 23204 1211 23238
rect 1273 23204 1307 23238
rect 2466 23208 2500 23242
rect 2562 23208 2596 23242
rect 2658 23208 2692 23242
rect 2754 23208 2788 23242
rect 2850 23208 2884 23242
rect 2946 23208 2980 23242
rect 3042 23208 3076 23242
rect 3138 23208 3172 23242
rect 3234 23208 3268 23242
rect 3330 23208 3364 23242
rect 3426 23208 3460 23242
rect 3647 23193 3681 23269
rect 3735 23193 3769 23269
rect 3987 23208 4021 23242
rect 4083 23208 4117 23242
rect 4179 23208 4213 23242
rect 4275 23208 4309 23242
rect 4371 23208 4405 23242
rect 4467 23208 4501 23242
rect 4563 23208 4597 23242
rect 4659 23208 4693 23242
rect 4755 23208 4789 23242
rect 4851 23208 4885 23242
rect 4947 23208 4981 23242
rect 5356 23278 5390 23312
rect 5356 23210 5390 23244
rect 5440 23278 5474 23312
rect 5440 23210 5474 23244
rect 313 21917 347 21951
rect 409 21917 443 21951
rect 505 21917 539 21951
rect 601 21917 635 21951
rect 697 21917 731 21951
rect 793 21917 827 21951
rect 889 21917 923 21951
rect 985 21917 1019 21951
rect 1081 21917 1115 21951
rect 1177 21917 1211 21951
rect 1273 21917 1307 21951
rect 2466 21921 2500 21955
rect 2562 21921 2596 21955
rect 2658 21921 2692 21955
rect 2754 21921 2788 21955
rect 2850 21921 2884 21955
rect 2946 21921 2980 21955
rect 3042 21921 3076 21955
rect 3138 21921 3172 21955
rect 3234 21921 3268 21955
rect 3330 21921 3364 21955
rect 3426 21921 3460 21955
rect 3647 21906 3681 21982
rect 3735 21906 3769 21982
rect 3987 21921 4021 21955
rect 4083 21921 4117 21955
rect 4179 21921 4213 21955
rect 4275 21921 4309 21955
rect 4371 21921 4405 21955
rect 4467 21921 4501 21955
rect 4563 21921 4597 21955
rect 4659 21921 4693 21955
rect 4755 21921 4789 21955
rect 4851 21921 4885 21955
rect 4947 21921 4981 21955
rect 5356 21991 5390 22025
rect 5356 21923 5390 21957
rect 5440 21991 5474 22025
rect 5440 21923 5474 21957
rect 313 20630 347 20664
rect 409 20630 443 20664
rect 505 20630 539 20664
rect 601 20630 635 20664
rect 697 20630 731 20664
rect 793 20630 827 20664
rect 889 20630 923 20664
rect 985 20630 1019 20664
rect 1081 20630 1115 20664
rect 1177 20630 1211 20664
rect 1273 20630 1307 20664
rect 2466 20634 2500 20668
rect 2562 20634 2596 20668
rect 2658 20634 2692 20668
rect 2754 20634 2788 20668
rect 2850 20634 2884 20668
rect 2946 20634 2980 20668
rect 3042 20634 3076 20668
rect 3138 20634 3172 20668
rect 3234 20634 3268 20668
rect 3330 20634 3364 20668
rect 3426 20634 3460 20668
rect 3647 20619 3681 20695
rect 3735 20619 3769 20695
rect 3987 20634 4021 20668
rect 4083 20634 4117 20668
rect 4179 20634 4213 20668
rect 4275 20634 4309 20668
rect 4371 20634 4405 20668
rect 4467 20634 4501 20668
rect 4563 20634 4597 20668
rect 4659 20634 4693 20668
rect 4755 20634 4789 20668
rect 4851 20634 4885 20668
rect 4947 20634 4981 20668
rect 5356 20704 5390 20738
rect 5356 20636 5390 20670
rect 5440 20704 5474 20738
rect 5440 20636 5474 20670
rect 313 19343 347 19377
rect 409 19343 443 19377
rect 505 19343 539 19377
rect 601 19343 635 19377
rect 697 19343 731 19377
rect 793 19343 827 19377
rect 889 19343 923 19377
rect 985 19343 1019 19377
rect 1081 19343 1115 19377
rect 1177 19343 1211 19377
rect 1273 19343 1307 19377
rect 2466 19347 2500 19381
rect 2562 19347 2596 19381
rect 2658 19347 2692 19381
rect 2754 19347 2788 19381
rect 2850 19347 2884 19381
rect 2946 19347 2980 19381
rect 3042 19347 3076 19381
rect 3138 19347 3172 19381
rect 3234 19347 3268 19381
rect 3330 19347 3364 19381
rect 3426 19347 3460 19381
rect 3647 19332 3681 19408
rect 3735 19332 3769 19408
rect 3987 19347 4021 19381
rect 4083 19347 4117 19381
rect 4179 19347 4213 19381
rect 4275 19347 4309 19381
rect 4371 19347 4405 19381
rect 4467 19347 4501 19381
rect 4563 19347 4597 19381
rect 4659 19347 4693 19381
rect 4755 19347 4789 19381
rect 4851 19347 4885 19381
rect 4947 19347 4981 19381
rect 5356 19417 5390 19451
rect 5356 19349 5390 19383
rect 5440 19417 5474 19451
rect 5440 19349 5474 19383
rect 313 18056 347 18090
rect 409 18056 443 18090
rect 505 18056 539 18090
rect 601 18056 635 18090
rect 697 18056 731 18090
rect 793 18056 827 18090
rect 889 18056 923 18090
rect 985 18056 1019 18090
rect 1081 18056 1115 18090
rect 1177 18056 1211 18090
rect 1273 18056 1307 18090
rect 2466 18060 2500 18094
rect 2562 18060 2596 18094
rect 2658 18060 2692 18094
rect 2754 18060 2788 18094
rect 2850 18060 2884 18094
rect 2946 18060 2980 18094
rect 3042 18060 3076 18094
rect 3138 18060 3172 18094
rect 3234 18060 3268 18094
rect 3330 18060 3364 18094
rect 3426 18060 3460 18094
rect 3647 18045 3681 18121
rect 3735 18045 3769 18121
rect 3987 18060 4021 18094
rect 4083 18060 4117 18094
rect 4179 18060 4213 18094
rect 4275 18060 4309 18094
rect 4371 18060 4405 18094
rect 4467 18060 4501 18094
rect 4563 18060 4597 18094
rect 4659 18060 4693 18094
rect 4755 18060 4789 18094
rect 4851 18060 4885 18094
rect 4947 18060 4981 18094
rect 5356 18130 5390 18164
rect 5356 18062 5390 18096
rect 5440 18130 5474 18164
rect 5440 18062 5474 18096
rect 313 16769 347 16803
rect 409 16769 443 16803
rect 505 16769 539 16803
rect 601 16769 635 16803
rect 697 16769 731 16803
rect 793 16769 827 16803
rect 889 16769 923 16803
rect 985 16769 1019 16803
rect 1081 16769 1115 16803
rect 1177 16769 1211 16803
rect 1273 16769 1307 16803
rect 2466 16773 2500 16807
rect 2562 16773 2596 16807
rect 2658 16773 2692 16807
rect 2754 16773 2788 16807
rect 2850 16773 2884 16807
rect 2946 16773 2980 16807
rect 3042 16773 3076 16807
rect 3138 16773 3172 16807
rect 3234 16773 3268 16807
rect 3330 16773 3364 16807
rect 3426 16773 3460 16807
rect 3647 16758 3681 16834
rect 3735 16758 3769 16834
rect 3987 16773 4021 16807
rect 4083 16773 4117 16807
rect 4179 16773 4213 16807
rect 4275 16773 4309 16807
rect 4371 16773 4405 16807
rect 4467 16773 4501 16807
rect 4563 16773 4597 16807
rect 4659 16773 4693 16807
rect 4755 16773 4789 16807
rect 4851 16773 4885 16807
rect 4947 16773 4981 16807
rect 5356 16843 5390 16877
rect 5356 16775 5390 16809
rect 5440 16843 5474 16877
rect 5440 16775 5474 16809
rect 313 15482 347 15516
rect 409 15482 443 15516
rect 505 15482 539 15516
rect 601 15482 635 15516
rect 697 15482 731 15516
rect 793 15482 827 15516
rect 889 15482 923 15516
rect 985 15482 1019 15516
rect 1081 15482 1115 15516
rect 1177 15482 1211 15516
rect 1273 15482 1307 15516
rect 2466 15486 2500 15520
rect 2562 15486 2596 15520
rect 2658 15486 2692 15520
rect 2754 15486 2788 15520
rect 2850 15486 2884 15520
rect 2946 15486 2980 15520
rect 3042 15486 3076 15520
rect 3138 15486 3172 15520
rect 3234 15486 3268 15520
rect 3330 15486 3364 15520
rect 3426 15486 3460 15520
rect 3647 15471 3681 15547
rect 3735 15471 3769 15547
rect 3987 15486 4021 15520
rect 4083 15486 4117 15520
rect 4179 15486 4213 15520
rect 4275 15486 4309 15520
rect 4371 15486 4405 15520
rect 4467 15486 4501 15520
rect 4563 15486 4597 15520
rect 4659 15486 4693 15520
rect 4755 15486 4789 15520
rect 4851 15486 4885 15520
rect 4947 15486 4981 15520
rect 5356 15556 5390 15590
rect 5356 15488 5390 15522
rect 5440 15556 5474 15590
rect 5440 15488 5474 15522
rect 313 14195 347 14229
rect 409 14195 443 14229
rect 505 14195 539 14229
rect 601 14195 635 14229
rect 697 14195 731 14229
rect 793 14195 827 14229
rect 889 14195 923 14229
rect 985 14195 1019 14229
rect 1081 14195 1115 14229
rect 1177 14195 1211 14229
rect 1273 14195 1307 14229
rect 2466 14199 2500 14233
rect 2562 14199 2596 14233
rect 2658 14199 2692 14233
rect 2754 14199 2788 14233
rect 2850 14199 2884 14233
rect 2946 14199 2980 14233
rect 3042 14199 3076 14233
rect 3138 14199 3172 14233
rect 3234 14199 3268 14233
rect 3330 14199 3364 14233
rect 3426 14199 3460 14233
rect 3647 14184 3681 14260
rect 3735 14184 3769 14260
rect 3987 14199 4021 14233
rect 4083 14199 4117 14233
rect 4179 14199 4213 14233
rect 4275 14199 4309 14233
rect 4371 14199 4405 14233
rect 4467 14199 4501 14233
rect 4563 14199 4597 14233
rect 4659 14199 4693 14233
rect 4755 14199 4789 14233
rect 4851 14199 4885 14233
rect 4947 14199 4981 14233
rect 5356 14269 5390 14303
rect 5356 14201 5390 14235
rect 5440 14269 5474 14303
rect 5440 14201 5474 14235
rect 313 12908 347 12942
rect 409 12908 443 12942
rect 505 12908 539 12942
rect 601 12908 635 12942
rect 697 12908 731 12942
rect 793 12908 827 12942
rect 889 12908 923 12942
rect 985 12908 1019 12942
rect 1081 12908 1115 12942
rect 1177 12908 1211 12942
rect 1273 12908 1307 12942
rect 2466 12912 2500 12946
rect 2562 12912 2596 12946
rect 2658 12912 2692 12946
rect 2754 12912 2788 12946
rect 2850 12912 2884 12946
rect 2946 12912 2980 12946
rect 3042 12912 3076 12946
rect 3138 12912 3172 12946
rect 3234 12912 3268 12946
rect 3330 12912 3364 12946
rect 3426 12912 3460 12946
rect 3647 12897 3681 12973
rect 3735 12897 3769 12973
rect 3987 12912 4021 12946
rect 4083 12912 4117 12946
rect 4179 12912 4213 12946
rect 4275 12912 4309 12946
rect 4371 12912 4405 12946
rect 4467 12912 4501 12946
rect 4563 12912 4597 12946
rect 4659 12912 4693 12946
rect 4755 12912 4789 12946
rect 4851 12912 4885 12946
rect 4947 12912 4981 12946
rect 5356 12982 5390 13016
rect 5356 12914 5390 12948
rect 5440 12982 5474 13016
rect 5440 12914 5474 12948
rect 313 11621 347 11655
rect 409 11621 443 11655
rect 505 11621 539 11655
rect 601 11621 635 11655
rect 697 11621 731 11655
rect 793 11621 827 11655
rect 889 11621 923 11655
rect 985 11621 1019 11655
rect 1081 11621 1115 11655
rect 1177 11621 1211 11655
rect 1273 11621 1307 11655
rect 2466 11625 2500 11659
rect 2562 11625 2596 11659
rect 2658 11625 2692 11659
rect 2754 11625 2788 11659
rect 2850 11625 2884 11659
rect 2946 11625 2980 11659
rect 3042 11625 3076 11659
rect 3138 11625 3172 11659
rect 3234 11625 3268 11659
rect 3330 11625 3364 11659
rect 3426 11625 3460 11659
rect 3647 11610 3681 11686
rect 3735 11610 3769 11686
rect 3987 11625 4021 11659
rect 4083 11625 4117 11659
rect 4179 11625 4213 11659
rect 4275 11625 4309 11659
rect 4371 11625 4405 11659
rect 4467 11625 4501 11659
rect 4563 11625 4597 11659
rect 4659 11625 4693 11659
rect 4755 11625 4789 11659
rect 4851 11625 4885 11659
rect 4947 11625 4981 11659
rect 5356 11695 5390 11729
rect 5356 11627 5390 11661
rect 5440 11695 5474 11729
rect 5440 11627 5474 11661
rect 313 10334 347 10368
rect 409 10334 443 10368
rect 505 10334 539 10368
rect 601 10334 635 10368
rect 697 10334 731 10368
rect 793 10334 827 10368
rect 889 10334 923 10368
rect 985 10334 1019 10368
rect 1081 10334 1115 10368
rect 1177 10334 1211 10368
rect 1273 10334 1307 10368
rect 2466 10338 2500 10372
rect 2562 10338 2596 10372
rect 2658 10338 2692 10372
rect 2754 10338 2788 10372
rect 2850 10338 2884 10372
rect 2946 10338 2980 10372
rect 3042 10338 3076 10372
rect 3138 10338 3172 10372
rect 3234 10338 3268 10372
rect 3330 10338 3364 10372
rect 3426 10338 3460 10372
rect 3647 10323 3681 10399
rect 3735 10323 3769 10399
rect 3987 10338 4021 10372
rect 4083 10338 4117 10372
rect 4179 10338 4213 10372
rect 4275 10338 4309 10372
rect 4371 10338 4405 10372
rect 4467 10338 4501 10372
rect 4563 10338 4597 10372
rect 4659 10338 4693 10372
rect 4755 10338 4789 10372
rect 4851 10338 4885 10372
rect 4947 10338 4981 10372
rect 5356 10408 5390 10442
rect 5356 10340 5390 10374
rect 5440 10408 5474 10442
rect 5440 10340 5474 10374
rect 313 9047 347 9081
rect 409 9047 443 9081
rect 505 9047 539 9081
rect 601 9047 635 9081
rect 697 9047 731 9081
rect 793 9047 827 9081
rect 889 9047 923 9081
rect 985 9047 1019 9081
rect 1081 9047 1115 9081
rect 1177 9047 1211 9081
rect 1273 9047 1307 9081
rect 2466 9051 2500 9085
rect 2562 9051 2596 9085
rect 2658 9051 2692 9085
rect 2754 9051 2788 9085
rect 2850 9051 2884 9085
rect 2946 9051 2980 9085
rect 3042 9051 3076 9085
rect 3138 9051 3172 9085
rect 3234 9051 3268 9085
rect 3330 9051 3364 9085
rect 3426 9051 3460 9085
rect 3647 9036 3681 9112
rect 3735 9036 3769 9112
rect 3987 9051 4021 9085
rect 4083 9051 4117 9085
rect 4179 9051 4213 9085
rect 4275 9051 4309 9085
rect 4371 9051 4405 9085
rect 4467 9051 4501 9085
rect 4563 9051 4597 9085
rect 4659 9051 4693 9085
rect 4755 9051 4789 9085
rect 4851 9051 4885 9085
rect 4947 9051 4981 9085
rect 5356 9121 5390 9155
rect 5356 9053 5390 9087
rect 5440 9121 5474 9155
rect 5440 9053 5474 9087
rect 313 7760 347 7794
rect 409 7760 443 7794
rect 505 7760 539 7794
rect 601 7760 635 7794
rect 697 7760 731 7794
rect 793 7760 827 7794
rect 889 7760 923 7794
rect 985 7760 1019 7794
rect 1081 7760 1115 7794
rect 1177 7760 1211 7794
rect 1273 7760 1307 7794
rect 2466 7764 2500 7798
rect 2562 7764 2596 7798
rect 2658 7764 2692 7798
rect 2754 7764 2788 7798
rect 2850 7764 2884 7798
rect 2946 7764 2980 7798
rect 3042 7764 3076 7798
rect 3138 7764 3172 7798
rect 3234 7764 3268 7798
rect 3330 7764 3364 7798
rect 3426 7764 3460 7798
rect 3647 7749 3681 7825
rect 3735 7749 3769 7825
rect 3987 7764 4021 7798
rect 4083 7764 4117 7798
rect 4179 7764 4213 7798
rect 4275 7764 4309 7798
rect 4371 7764 4405 7798
rect 4467 7764 4501 7798
rect 4563 7764 4597 7798
rect 4659 7764 4693 7798
rect 4755 7764 4789 7798
rect 4851 7764 4885 7798
rect 4947 7764 4981 7798
rect 5356 7834 5390 7868
rect 5356 7766 5390 7800
rect 5440 7834 5474 7868
rect 5440 7766 5474 7800
rect 313 6473 347 6507
rect 409 6473 443 6507
rect 505 6473 539 6507
rect 601 6473 635 6507
rect 697 6473 731 6507
rect 793 6473 827 6507
rect 889 6473 923 6507
rect 985 6473 1019 6507
rect 1081 6473 1115 6507
rect 1177 6473 1211 6507
rect 1273 6473 1307 6507
rect 2466 6477 2500 6511
rect 2562 6477 2596 6511
rect 2658 6477 2692 6511
rect 2754 6477 2788 6511
rect 2850 6477 2884 6511
rect 2946 6477 2980 6511
rect 3042 6477 3076 6511
rect 3138 6477 3172 6511
rect 3234 6477 3268 6511
rect 3330 6477 3364 6511
rect 3426 6477 3460 6511
rect 3647 6462 3681 6538
rect 3735 6462 3769 6538
rect 3987 6477 4021 6511
rect 4083 6477 4117 6511
rect 4179 6477 4213 6511
rect 4275 6477 4309 6511
rect 4371 6477 4405 6511
rect 4467 6477 4501 6511
rect 4563 6477 4597 6511
rect 4659 6477 4693 6511
rect 4755 6477 4789 6511
rect 4851 6477 4885 6511
rect 4947 6477 4981 6511
rect 5356 6547 5390 6581
rect 5356 6479 5390 6513
rect 5440 6547 5474 6581
rect 5440 6479 5474 6513
rect 313 5186 347 5220
rect 409 5186 443 5220
rect 505 5186 539 5220
rect 601 5186 635 5220
rect 697 5186 731 5220
rect 793 5186 827 5220
rect 889 5186 923 5220
rect 985 5186 1019 5220
rect 1081 5186 1115 5220
rect 1177 5186 1211 5220
rect 1273 5186 1307 5220
rect 2466 5190 2500 5224
rect 2562 5190 2596 5224
rect 2658 5190 2692 5224
rect 2754 5190 2788 5224
rect 2850 5190 2884 5224
rect 2946 5190 2980 5224
rect 3042 5190 3076 5224
rect 3138 5190 3172 5224
rect 3234 5190 3268 5224
rect 3330 5190 3364 5224
rect 3426 5190 3460 5224
rect 3647 5175 3681 5251
rect 3735 5175 3769 5251
rect 3987 5190 4021 5224
rect 4083 5190 4117 5224
rect 4179 5190 4213 5224
rect 4275 5190 4309 5224
rect 4371 5190 4405 5224
rect 4467 5190 4501 5224
rect 4563 5190 4597 5224
rect 4659 5190 4693 5224
rect 4755 5190 4789 5224
rect 4851 5190 4885 5224
rect 4947 5190 4981 5224
rect 5356 5260 5390 5294
rect 5356 5192 5390 5226
rect 5440 5260 5474 5294
rect 5440 5192 5474 5226
rect 313 3899 347 3933
rect 409 3899 443 3933
rect 505 3899 539 3933
rect 601 3899 635 3933
rect 697 3899 731 3933
rect 793 3899 827 3933
rect 889 3899 923 3933
rect 985 3899 1019 3933
rect 1081 3899 1115 3933
rect 1177 3899 1211 3933
rect 1273 3899 1307 3933
rect 2466 3903 2500 3937
rect 2562 3903 2596 3937
rect 2658 3903 2692 3937
rect 2754 3903 2788 3937
rect 2850 3903 2884 3937
rect 2946 3903 2980 3937
rect 3042 3903 3076 3937
rect 3138 3903 3172 3937
rect 3234 3903 3268 3937
rect 3330 3903 3364 3937
rect 3426 3903 3460 3937
rect 3647 3888 3681 3964
rect 3735 3888 3769 3964
rect 3987 3903 4021 3937
rect 4083 3903 4117 3937
rect 4179 3903 4213 3937
rect 4275 3903 4309 3937
rect 4371 3903 4405 3937
rect 4467 3903 4501 3937
rect 4563 3903 4597 3937
rect 4659 3903 4693 3937
rect 4755 3903 4789 3937
rect 4851 3903 4885 3937
rect 4947 3903 4981 3937
rect 5356 3973 5390 4007
rect 5356 3905 5390 3939
rect 5440 3973 5474 4007
rect 5440 3905 5474 3939
rect 313 2612 347 2646
rect 409 2612 443 2646
rect 505 2612 539 2646
rect 601 2612 635 2646
rect 697 2612 731 2646
rect 793 2612 827 2646
rect 889 2612 923 2646
rect 985 2612 1019 2646
rect 1081 2612 1115 2646
rect 1177 2612 1211 2646
rect 1273 2612 1307 2646
rect 2466 2616 2500 2650
rect 2562 2616 2596 2650
rect 2658 2616 2692 2650
rect 2754 2616 2788 2650
rect 2850 2616 2884 2650
rect 2946 2616 2980 2650
rect 3042 2616 3076 2650
rect 3138 2616 3172 2650
rect 3234 2616 3268 2650
rect 3330 2616 3364 2650
rect 3426 2616 3460 2650
rect 3647 2601 3681 2677
rect 3735 2601 3769 2677
rect 3987 2616 4021 2650
rect 4083 2616 4117 2650
rect 4179 2616 4213 2650
rect 4275 2616 4309 2650
rect 4371 2616 4405 2650
rect 4467 2616 4501 2650
rect 4563 2616 4597 2650
rect 4659 2616 4693 2650
rect 4755 2616 4789 2650
rect 4851 2616 4885 2650
rect 4947 2616 4981 2650
rect 5356 2686 5390 2720
rect 5356 2618 5390 2652
rect 5440 2686 5474 2720
rect 5440 2618 5474 2652
rect 313 1325 347 1359
rect 409 1325 443 1359
rect 505 1325 539 1359
rect 601 1325 635 1359
rect 697 1325 731 1359
rect 793 1325 827 1359
rect 889 1325 923 1359
rect 985 1325 1019 1359
rect 1081 1325 1115 1359
rect 1177 1325 1211 1359
rect 1273 1325 1307 1359
rect 2466 1329 2500 1363
rect 2562 1329 2596 1363
rect 2658 1329 2692 1363
rect 2754 1329 2788 1363
rect 2850 1329 2884 1363
rect 2946 1329 2980 1363
rect 3042 1329 3076 1363
rect 3138 1329 3172 1363
rect 3234 1329 3268 1363
rect 3330 1329 3364 1363
rect 3426 1329 3460 1363
rect 3647 1314 3681 1390
rect 3735 1314 3769 1390
rect 3987 1329 4021 1363
rect 4083 1329 4117 1363
rect 4179 1329 4213 1363
rect 4275 1329 4309 1363
rect 4371 1329 4405 1363
rect 4467 1329 4501 1363
rect 4563 1329 4597 1363
rect 4659 1329 4693 1363
rect 4755 1329 4789 1363
rect 4851 1329 4885 1363
rect 4947 1329 4981 1363
rect 5356 1399 5390 1433
rect 5356 1331 5390 1365
rect 5440 1399 5474 1433
rect 5440 1331 5474 1365
<< pdiffc >>
rect 313 41820 347 41854
rect 313 41752 347 41786
rect 313 41684 347 41718
rect 313 41616 347 41650
rect 409 41820 443 41854
rect 409 41752 443 41786
rect 409 41684 443 41718
rect 409 41616 443 41650
rect 505 41820 539 41854
rect 505 41752 539 41786
rect 505 41684 539 41718
rect 505 41616 539 41650
rect 601 41820 635 41854
rect 601 41752 635 41786
rect 601 41684 635 41718
rect 601 41616 635 41650
rect 697 41820 731 41854
rect 697 41752 731 41786
rect 697 41684 731 41718
rect 697 41616 731 41650
rect 793 41820 827 41854
rect 793 41752 827 41786
rect 793 41684 827 41718
rect 793 41616 827 41650
rect 889 41820 923 41854
rect 889 41752 923 41786
rect 889 41684 923 41718
rect 889 41616 923 41650
rect 985 41820 1019 41854
rect 985 41752 1019 41786
rect 985 41684 1019 41718
rect 985 41616 1019 41650
rect 1081 41820 1115 41854
rect 1081 41752 1115 41786
rect 1081 41684 1115 41718
rect 1081 41616 1115 41650
rect 1177 41820 1211 41854
rect 1177 41752 1211 41786
rect 1177 41684 1211 41718
rect 1177 41616 1211 41650
rect 1273 41820 1307 41854
rect 1273 41752 1307 41786
rect 1273 41684 1307 41718
rect 1273 41616 1307 41650
rect 2466 41824 2500 41858
rect 2466 41756 2500 41790
rect 2466 41688 2500 41722
rect 2466 41620 2500 41654
rect 2562 41824 2596 41858
rect 2562 41756 2596 41790
rect 2562 41688 2596 41722
rect 2562 41620 2596 41654
rect 2658 41824 2692 41858
rect 2658 41756 2692 41790
rect 2658 41688 2692 41722
rect 2658 41620 2692 41654
rect 2754 41824 2788 41858
rect 2754 41756 2788 41790
rect 2754 41688 2788 41722
rect 2754 41620 2788 41654
rect 2850 41824 2884 41858
rect 2850 41756 2884 41790
rect 2850 41688 2884 41722
rect 2850 41620 2884 41654
rect 2946 41824 2980 41858
rect 2946 41756 2980 41790
rect 2946 41688 2980 41722
rect 2946 41620 2980 41654
rect 3042 41824 3076 41858
rect 3042 41756 3076 41790
rect 3042 41688 3076 41722
rect 3042 41620 3076 41654
rect 3138 41824 3172 41858
rect 3138 41756 3172 41790
rect 3138 41688 3172 41722
rect 3138 41620 3172 41654
rect 3234 41824 3268 41858
rect 3234 41756 3268 41790
rect 3234 41688 3268 41722
rect 3234 41620 3268 41654
rect 3330 41824 3364 41858
rect 3330 41756 3364 41790
rect 3330 41688 3364 41722
rect 3330 41620 3364 41654
rect 3426 41824 3460 41858
rect 3426 41756 3460 41790
rect 3426 41688 3460 41722
rect 3426 41620 3460 41654
rect 3987 41824 4021 41858
rect 3987 41756 4021 41790
rect 3987 41688 4021 41722
rect 3987 41620 4021 41654
rect 4083 41824 4117 41858
rect 4083 41756 4117 41790
rect 4083 41688 4117 41722
rect 4083 41620 4117 41654
rect 4179 41824 4213 41858
rect 4179 41756 4213 41790
rect 4179 41688 4213 41722
rect 4179 41620 4213 41654
rect 4275 41824 4309 41858
rect 4275 41756 4309 41790
rect 4275 41688 4309 41722
rect 4275 41620 4309 41654
rect 4371 41824 4405 41858
rect 4371 41756 4405 41790
rect 4371 41688 4405 41722
rect 4371 41620 4405 41654
rect 4467 41824 4501 41858
rect 4467 41756 4501 41790
rect 4467 41688 4501 41722
rect 4467 41620 4501 41654
rect 4563 41824 4597 41858
rect 4563 41756 4597 41790
rect 4563 41688 4597 41722
rect 4563 41620 4597 41654
rect 4659 41824 4693 41858
rect 4659 41756 4693 41790
rect 4659 41688 4693 41722
rect 4659 41620 4693 41654
rect 4755 41824 4789 41858
rect 4755 41756 4789 41790
rect 4755 41688 4789 41722
rect 4755 41620 4789 41654
rect 4851 41824 4885 41858
rect 4851 41756 4885 41790
rect 4851 41688 4885 41722
rect 4851 41620 4885 41654
rect 4947 41824 4981 41858
rect 4947 41756 4981 41790
rect 4947 41688 4981 41722
rect 4947 41620 4981 41654
rect 5356 41616 5390 41650
rect 5356 41548 5390 41582
rect 5356 41480 5390 41514
rect 5440 41616 5474 41650
rect 5440 41548 5474 41582
rect 5440 41480 5474 41514
rect 313 40533 347 40567
rect 313 40465 347 40499
rect 313 40397 347 40431
rect 313 40329 347 40363
rect 409 40533 443 40567
rect 409 40465 443 40499
rect 409 40397 443 40431
rect 409 40329 443 40363
rect 505 40533 539 40567
rect 505 40465 539 40499
rect 505 40397 539 40431
rect 505 40329 539 40363
rect 601 40533 635 40567
rect 601 40465 635 40499
rect 601 40397 635 40431
rect 601 40329 635 40363
rect 697 40533 731 40567
rect 697 40465 731 40499
rect 697 40397 731 40431
rect 697 40329 731 40363
rect 793 40533 827 40567
rect 793 40465 827 40499
rect 793 40397 827 40431
rect 793 40329 827 40363
rect 889 40533 923 40567
rect 889 40465 923 40499
rect 889 40397 923 40431
rect 889 40329 923 40363
rect 985 40533 1019 40567
rect 985 40465 1019 40499
rect 985 40397 1019 40431
rect 985 40329 1019 40363
rect 1081 40533 1115 40567
rect 1081 40465 1115 40499
rect 1081 40397 1115 40431
rect 1081 40329 1115 40363
rect 1177 40533 1211 40567
rect 1177 40465 1211 40499
rect 1177 40397 1211 40431
rect 1177 40329 1211 40363
rect 1273 40533 1307 40567
rect 1273 40465 1307 40499
rect 1273 40397 1307 40431
rect 1273 40329 1307 40363
rect 2466 40537 2500 40571
rect 2466 40469 2500 40503
rect 2466 40401 2500 40435
rect 2466 40333 2500 40367
rect 2562 40537 2596 40571
rect 2562 40469 2596 40503
rect 2562 40401 2596 40435
rect 2562 40333 2596 40367
rect 2658 40537 2692 40571
rect 2658 40469 2692 40503
rect 2658 40401 2692 40435
rect 2658 40333 2692 40367
rect 2754 40537 2788 40571
rect 2754 40469 2788 40503
rect 2754 40401 2788 40435
rect 2754 40333 2788 40367
rect 2850 40537 2884 40571
rect 2850 40469 2884 40503
rect 2850 40401 2884 40435
rect 2850 40333 2884 40367
rect 2946 40537 2980 40571
rect 2946 40469 2980 40503
rect 2946 40401 2980 40435
rect 2946 40333 2980 40367
rect 3042 40537 3076 40571
rect 3042 40469 3076 40503
rect 3042 40401 3076 40435
rect 3042 40333 3076 40367
rect 3138 40537 3172 40571
rect 3138 40469 3172 40503
rect 3138 40401 3172 40435
rect 3138 40333 3172 40367
rect 3234 40537 3268 40571
rect 3234 40469 3268 40503
rect 3234 40401 3268 40435
rect 3234 40333 3268 40367
rect 3330 40537 3364 40571
rect 3330 40469 3364 40503
rect 3330 40401 3364 40435
rect 3330 40333 3364 40367
rect 3426 40537 3460 40571
rect 3426 40469 3460 40503
rect 3426 40401 3460 40435
rect 3426 40333 3460 40367
rect 3987 40537 4021 40571
rect 3987 40469 4021 40503
rect 3987 40401 4021 40435
rect 3987 40333 4021 40367
rect 4083 40537 4117 40571
rect 4083 40469 4117 40503
rect 4083 40401 4117 40435
rect 4083 40333 4117 40367
rect 4179 40537 4213 40571
rect 4179 40469 4213 40503
rect 4179 40401 4213 40435
rect 4179 40333 4213 40367
rect 4275 40537 4309 40571
rect 4275 40469 4309 40503
rect 4275 40401 4309 40435
rect 4275 40333 4309 40367
rect 4371 40537 4405 40571
rect 4371 40469 4405 40503
rect 4371 40401 4405 40435
rect 4371 40333 4405 40367
rect 4467 40537 4501 40571
rect 4467 40469 4501 40503
rect 4467 40401 4501 40435
rect 4467 40333 4501 40367
rect 4563 40537 4597 40571
rect 4563 40469 4597 40503
rect 4563 40401 4597 40435
rect 4563 40333 4597 40367
rect 4659 40537 4693 40571
rect 4659 40469 4693 40503
rect 4659 40401 4693 40435
rect 4659 40333 4693 40367
rect 4755 40537 4789 40571
rect 4755 40469 4789 40503
rect 4755 40401 4789 40435
rect 4755 40333 4789 40367
rect 4851 40537 4885 40571
rect 4851 40469 4885 40503
rect 4851 40401 4885 40435
rect 4851 40333 4885 40367
rect 4947 40537 4981 40571
rect 4947 40469 4981 40503
rect 4947 40401 4981 40435
rect 4947 40333 4981 40367
rect 5356 40329 5390 40363
rect 5356 40261 5390 40295
rect 5356 40193 5390 40227
rect 5440 40329 5474 40363
rect 5440 40261 5474 40295
rect 5440 40193 5474 40227
rect 313 39246 347 39280
rect 313 39178 347 39212
rect 313 39110 347 39144
rect 313 39042 347 39076
rect 409 39246 443 39280
rect 409 39178 443 39212
rect 409 39110 443 39144
rect 409 39042 443 39076
rect 505 39246 539 39280
rect 505 39178 539 39212
rect 505 39110 539 39144
rect 505 39042 539 39076
rect 601 39246 635 39280
rect 601 39178 635 39212
rect 601 39110 635 39144
rect 601 39042 635 39076
rect 697 39246 731 39280
rect 697 39178 731 39212
rect 697 39110 731 39144
rect 697 39042 731 39076
rect 793 39246 827 39280
rect 793 39178 827 39212
rect 793 39110 827 39144
rect 793 39042 827 39076
rect 889 39246 923 39280
rect 889 39178 923 39212
rect 889 39110 923 39144
rect 889 39042 923 39076
rect 985 39246 1019 39280
rect 985 39178 1019 39212
rect 985 39110 1019 39144
rect 985 39042 1019 39076
rect 1081 39246 1115 39280
rect 1081 39178 1115 39212
rect 1081 39110 1115 39144
rect 1081 39042 1115 39076
rect 1177 39246 1211 39280
rect 1177 39178 1211 39212
rect 1177 39110 1211 39144
rect 1177 39042 1211 39076
rect 1273 39246 1307 39280
rect 1273 39178 1307 39212
rect 1273 39110 1307 39144
rect 1273 39042 1307 39076
rect 2466 39250 2500 39284
rect 2466 39182 2500 39216
rect 2466 39114 2500 39148
rect 2466 39046 2500 39080
rect 2562 39250 2596 39284
rect 2562 39182 2596 39216
rect 2562 39114 2596 39148
rect 2562 39046 2596 39080
rect 2658 39250 2692 39284
rect 2658 39182 2692 39216
rect 2658 39114 2692 39148
rect 2658 39046 2692 39080
rect 2754 39250 2788 39284
rect 2754 39182 2788 39216
rect 2754 39114 2788 39148
rect 2754 39046 2788 39080
rect 2850 39250 2884 39284
rect 2850 39182 2884 39216
rect 2850 39114 2884 39148
rect 2850 39046 2884 39080
rect 2946 39250 2980 39284
rect 2946 39182 2980 39216
rect 2946 39114 2980 39148
rect 2946 39046 2980 39080
rect 3042 39250 3076 39284
rect 3042 39182 3076 39216
rect 3042 39114 3076 39148
rect 3042 39046 3076 39080
rect 3138 39250 3172 39284
rect 3138 39182 3172 39216
rect 3138 39114 3172 39148
rect 3138 39046 3172 39080
rect 3234 39250 3268 39284
rect 3234 39182 3268 39216
rect 3234 39114 3268 39148
rect 3234 39046 3268 39080
rect 3330 39250 3364 39284
rect 3330 39182 3364 39216
rect 3330 39114 3364 39148
rect 3330 39046 3364 39080
rect 3426 39250 3460 39284
rect 3426 39182 3460 39216
rect 3426 39114 3460 39148
rect 3426 39046 3460 39080
rect 3987 39250 4021 39284
rect 3987 39182 4021 39216
rect 3987 39114 4021 39148
rect 3987 39046 4021 39080
rect 4083 39250 4117 39284
rect 4083 39182 4117 39216
rect 4083 39114 4117 39148
rect 4083 39046 4117 39080
rect 4179 39250 4213 39284
rect 4179 39182 4213 39216
rect 4179 39114 4213 39148
rect 4179 39046 4213 39080
rect 4275 39250 4309 39284
rect 4275 39182 4309 39216
rect 4275 39114 4309 39148
rect 4275 39046 4309 39080
rect 4371 39250 4405 39284
rect 4371 39182 4405 39216
rect 4371 39114 4405 39148
rect 4371 39046 4405 39080
rect 4467 39250 4501 39284
rect 4467 39182 4501 39216
rect 4467 39114 4501 39148
rect 4467 39046 4501 39080
rect 4563 39250 4597 39284
rect 4563 39182 4597 39216
rect 4563 39114 4597 39148
rect 4563 39046 4597 39080
rect 4659 39250 4693 39284
rect 4659 39182 4693 39216
rect 4659 39114 4693 39148
rect 4659 39046 4693 39080
rect 4755 39250 4789 39284
rect 4755 39182 4789 39216
rect 4755 39114 4789 39148
rect 4755 39046 4789 39080
rect 4851 39250 4885 39284
rect 4851 39182 4885 39216
rect 4851 39114 4885 39148
rect 4851 39046 4885 39080
rect 4947 39250 4981 39284
rect 4947 39182 4981 39216
rect 4947 39114 4981 39148
rect 4947 39046 4981 39080
rect 5356 39042 5390 39076
rect 5356 38974 5390 39008
rect 5356 38906 5390 38940
rect 5440 39042 5474 39076
rect 5440 38974 5474 39008
rect 5440 38906 5474 38940
rect 313 37959 347 37993
rect 313 37891 347 37925
rect 313 37823 347 37857
rect 313 37755 347 37789
rect 409 37959 443 37993
rect 409 37891 443 37925
rect 409 37823 443 37857
rect 409 37755 443 37789
rect 505 37959 539 37993
rect 505 37891 539 37925
rect 505 37823 539 37857
rect 505 37755 539 37789
rect 601 37959 635 37993
rect 601 37891 635 37925
rect 601 37823 635 37857
rect 601 37755 635 37789
rect 697 37959 731 37993
rect 697 37891 731 37925
rect 697 37823 731 37857
rect 697 37755 731 37789
rect 793 37959 827 37993
rect 793 37891 827 37925
rect 793 37823 827 37857
rect 793 37755 827 37789
rect 889 37959 923 37993
rect 889 37891 923 37925
rect 889 37823 923 37857
rect 889 37755 923 37789
rect 985 37959 1019 37993
rect 985 37891 1019 37925
rect 985 37823 1019 37857
rect 985 37755 1019 37789
rect 1081 37959 1115 37993
rect 1081 37891 1115 37925
rect 1081 37823 1115 37857
rect 1081 37755 1115 37789
rect 1177 37959 1211 37993
rect 1177 37891 1211 37925
rect 1177 37823 1211 37857
rect 1177 37755 1211 37789
rect 1273 37959 1307 37993
rect 1273 37891 1307 37925
rect 1273 37823 1307 37857
rect 1273 37755 1307 37789
rect 2466 37963 2500 37997
rect 2466 37895 2500 37929
rect 2466 37827 2500 37861
rect 2466 37759 2500 37793
rect 2562 37963 2596 37997
rect 2562 37895 2596 37929
rect 2562 37827 2596 37861
rect 2562 37759 2596 37793
rect 2658 37963 2692 37997
rect 2658 37895 2692 37929
rect 2658 37827 2692 37861
rect 2658 37759 2692 37793
rect 2754 37963 2788 37997
rect 2754 37895 2788 37929
rect 2754 37827 2788 37861
rect 2754 37759 2788 37793
rect 2850 37963 2884 37997
rect 2850 37895 2884 37929
rect 2850 37827 2884 37861
rect 2850 37759 2884 37793
rect 2946 37963 2980 37997
rect 2946 37895 2980 37929
rect 2946 37827 2980 37861
rect 2946 37759 2980 37793
rect 3042 37963 3076 37997
rect 3042 37895 3076 37929
rect 3042 37827 3076 37861
rect 3042 37759 3076 37793
rect 3138 37963 3172 37997
rect 3138 37895 3172 37929
rect 3138 37827 3172 37861
rect 3138 37759 3172 37793
rect 3234 37963 3268 37997
rect 3234 37895 3268 37929
rect 3234 37827 3268 37861
rect 3234 37759 3268 37793
rect 3330 37963 3364 37997
rect 3330 37895 3364 37929
rect 3330 37827 3364 37861
rect 3330 37759 3364 37793
rect 3426 37963 3460 37997
rect 3426 37895 3460 37929
rect 3426 37827 3460 37861
rect 3426 37759 3460 37793
rect 3987 37963 4021 37997
rect 3987 37895 4021 37929
rect 3987 37827 4021 37861
rect 3987 37759 4021 37793
rect 4083 37963 4117 37997
rect 4083 37895 4117 37929
rect 4083 37827 4117 37861
rect 4083 37759 4117 37793
rect 4179 37963 4213 37997
rect 4179 37895 4213 37929
rect 4179 37827 4213 37861
rect 4179 37759 4213 37793
rect 4275 37963 4309 37997
rect 4275 37895 4309 37929
rect 4275 37827 4309 37861
rect 4275 37759 4309 37793
rect 4371 37963 4405 37997
rect 4371 37895 4405 37929
rect 4371 37827 4405 37861
rect 4371 37759 4405 37793
rect 4467 37963 4501 37997
rect 4467 37895 4501 37929
rect 4467 37827 4501 37861
rect 4467 37759 4501 37793
rect 4563 37963 4597 37997
rect 4563 37895 4597 37929
rect 4563 37827 4597 37861
rect 4563 37759 4597 37793
rect 4659 37963 4693 37997
rect 4659 37895 4693 37929
rect 4659 37827 4693 37861
rect 4659 37759 4693 37793
rect 4755 37963 4789 37997
rect 4755 37895 4789 37929
rect 4755 37827 4789 37861
rect 4755 37759 4789 37793
rect 4851 37963 4885 37997
rect 4851 37895 4885 37929
rect 4851 37827 4885 37861
rect 4851 37759 4885 37793
rect 4947 37963 4981 37997
rect 4947 37895 4981 37929
rect 4947 37827 4981 37861
rect 4947 37759 4981 37793
rect 5356 37755 5390 37789
rect 5356 37687 5390 37721
rect 5356 37619 5390 37653
rect 5440 37755 5474 37789
rect 5440 37687 5474 37721
rect 5440 37619 5474 37653
rect 313 36672 347 36706
rect 313 36604 347 36638
rect 313 36536 347 36570
rect 313 36468 347 36502
rect 409 36672 443 36706
rect 409 36604 443 36638
rect 409 36536 443 36570
rect 409 36468 443 36502
rect 505 36672 539 36706
rect 505 36604 539 36638
rect 505 36536 539 36570
rect 505 36468 539 36502
rect 601 36672 635 36706
rect 601 36604 635 36638
rect 601 36536 635 36570
rect 601 36468 635 36502
rect 697 36672 731 36706
rect 697 36604 731 36638
rect 697 36536 731 36570
rect 697 36468 731 36502
rect 793 36672 827 36706
rect 793 36604 827 36638
rect 793 36536 827 36570
rect 793 36468 827 36502
rect 889 36672 923 36706
rect 889 36604 923 36638
rect 889 36536 923 36570
rect 889 36468 923 36502
rect 985 36672 1019 36706
rect 985 36604 1019 36638
rect 985 36536 1019 36570
rect 985 36468 1019 36502
rect 1081 36672 1115 36706
rect 1081 36604 1115 36638
rect 1081 36536 1115 36570
rect 1081 36468 1115 36502
rect 1177 36672 1211 36706
rect 1177 36604 1211 36638
rect 1177 36536 1211 36570
rect 1177 36468 1211 36502
rect 1273 36672 1307 36706
rect 1273 36604 1307 36638
rect 1273 36536 1307 36570
rect 1273 36468 1307 36502
rect 2466 36676 2500 36710
rect 2466 36608 2500 36642
rect 2466 36540 2500 36574
rect 2466 36472 2500 36506
rect 2562 36676 2596 36710
rect 2562 36608 2596 36642
rect 2562 36540 2596 36574
rect 2562 36472 2596 36506
rect 2658 36676 2692 36710
rect 2658 36608 2692 36642
rect 2658 36540 2692 36574
rect 2658 36472 2692 36506
rect 2754 36676 2788 36710
rect 2754 36608 2788 36642
rect 2754 36540 2788 36574
rect 2754 36472 2788 36506
rect 2850 36676 2884 36710
rect 2850 36608 2884 36642
rect 2850 36540 2884 36574
rect 2850 36472 2884 36506
rect 2946 36676 2980 36710
rect 2946 36608 2980 36642
rect 2946 36540 2980 36574
rect 2946 36472 2980 36506
rect 3042 36676 3076 36710
rect 3042 36608 3076 36642
rect 3042 36540 3076 36574
rect 3042 36472 3076 36506
rect 3138 36676 3172 36710
rect 3138 36608 3172 36642
rect 3138 36540 3172 36574
rect 3138 36472 3172 36506
rect 3234 36676 3268 36710
rect 3234 36608 3268 36642
rect 3234 36540 3268 36574
rect 3234 36472 3268 36506
rect 3330 36676 3364 36710
rect 3330 36608 3364 36642
rect 3330 36540 3364 36574
rect 3330 36472 3364 36506
rect 3426 36676 3460 36710
rect 3426 36608 3460 36642
rect 3426 36540 3460 36574
rect 3426 36472 3460 36506
rect 3987 36676 4021 36710
rect 3987 36608 4021 36642
rect 3987 36540 4021 36574
rect 3987 36472 4021 36506
rect 4083 36676 4117 36710
rect 4083 36608 4117 36642
rect 4083 36540 4117 36574
rect 4083 36472 4117 36506
rect 4179 36676 4213 36710
rect 4179 36608 4213 36642
rect 4179 36540 4213 36574
rect 4179 36472 4213 36506
rect 4275 36676 4309 36710
rect 4275 36608 4309 36642
rect 4275 36540 4309 36574
rect 4275 36472 4309 36506
rect 4371 36676 4405 36710
rect 4371 36608 4405 36642
rect 4371 36540 4405 36574
rect 4371 36472 4405 36506
rect 4467 36676 4501 36710
rect 4467 36608 4501 36642
rect 4467 36540 4501 36574
rect 4467 36472 4501 36506
rect 4563 36676 4597 36710
rect 4563 36608 4597 36642
rect 4563 36540 4597 36574
rect 4563 36472 4597 36506
rect 4659 36676 4693 36710
rect 4659 36608 4693 36642
rect 4659 36540 4693 36574
rect 4659 36472 4693 36506
rect 4755 36676 4789 36710
rect 4755 36608 4789 36642
rect 4755 36540 4789 36574
rect 4755 36472 4789 36506
rect 4851 36676 4885 36710
rect 4851 36608 4885 36642
rect 4851 36540 4885 36574
rect 4851 36472 4885 36506
rect 4947 36676 4981 36710
rect 4947 36608 4981 36642
rect 4947 36540 4981 36574
rect 4947 36472 4981 36506
rect 5356 36468 5390 36502
rect 5356 36400 5390 36434
rect 5356 36332 5390 36366
rect 5440 36468 5474 36502
rect 5440 36400 5474 36434
rect 5440 36332 5474 36366
rect 313 35385 347 35419
rect 313 35317 347 35351
rect 313 35249 347 35283
rect 313 35181 347 35215
rect 409 35385 443 35419
rect 409 35317 443 35351
rect 409 35249 443 35283
rect 409 35181 443 35215
rect 505 35385 539 35419
rect 505 35317 539 35351
rect 505 35249 539 35283
rect 505 35181 539 35215
rect 601 35385 635 35419
rect 601 35317 635 35351
rect 601 35249 635 35283
rect 601 35181 635 35215
rect 697 35385 731 35419
rect 697 35317 731 35351
rect 697 35249 731 35283
rect 697 35181 731 35215
rect 793 35385 827 35419
rect 793 35317 827 35351
rect 793 35249 827 35283
rect 793 35181 827 35215
rect 889 35385 923 35419
rect 889 35317 923 35351
rect 889 35249 923 35283
rect 889 35181 923 35215
rect 985 35385 1019 35419
rect 985 35317 1019 35351
rect 985 35249 1019 35283
rect 985 35181 1019 35215
rect 1081 35385 1115 35419
rect 1081 35317 1115 35351
rect 1081 35249 1115 35283
rect 1081 35181 1115 35215
rect 1177 35385 1211 35419
rect 1177 35317 1211 35351
rect 1177 35249 1211 35283
rect 1177 35181 1211 35215
rect 1273 35385 1307 35419
rect 1273 35317 1307 35351
rect 1273 35249 1307 35283
rect 1273 35181 1307 35215
rect 2466 35389 2500 35423
rect 2466 35321 2500 35355
rect 2466 35253 2500 35287
rect 2466 35185 2500 35219
rect 2562 35389 2596 35423
rect 2562 35321 2596 35355
rect 2562 35253 2596 35287
rect 2562 35185 2596 35219
rect 2658 35389 2692 35423
rect 2658 35321 2692 35355
rect 2658 35253 2692 35287
rect 2658 35185 2692 35219
rect 2754 35389 2788 35423
rect 2754 35321 2788 35355
rect 2754 35253 2788 35287
rect 2754 35185 2788 35219
rect 2850 35389 2884 35423
rect 2850 35321 2884 35355
rect 2850 35253 2884 35287
rect 2850 35185 2884 35219
rect 2946 35389 2980 35423
rect 2946 35321 2980 35355
rect 2946 35253 2980 35287
rect 2946 35185 2980 35219
rect 3042 35389 3076 35423
rect 3042 35321 3076 35355
rect 3042 35253 3076 35287
rect 3042 35185 3076 35219
rect 3138 35389 3172 35423
rect 3138 35321 3172 35355
rect 3138 35253 3172 35287
rect 3138 35185 3172 35219
rect 3234 35389 3268 35423
rect 3234 35321 3268 35355
rect 3234 35253 3268 35287
rect 3234 35185 3268 35219
rect 3330 35389 3364 35423
rect 3330 35321 3364 35355
rect 3330 35253 3364 35287
rect 3330 35185 3364 35219
rect 3426 35389 3460 35423
rect 3426 35321 3460 35355
rect 3426 35253 3460 35287
rect 3426 35185 3460 35219
rect 3987 35389 4021 35423
rect 3987 35321 4021 35355
rect 3987 35253 4021 35287
rect 3987 35185 4021 35219
rect 4083 35389 4117 35423
rect 4083 35321 4117 35355
rect 4083 35253 4117 35287
rect 4083 35185 4117 35219
rect 4179 35389 4213 35423
rect 4179 35321 4213 35355
rect 4179 35253 4213 35287
rect 4179 35185 4213 35219
rect 4275 35389 4309 35423
rect 4275 35321 4309 35355
rect 4275 35253 4309 35287
rect 4275 35185 4309 35219
rect 4371 35389 4405 35423
rect 4371 35321 4405 35355
rect 4371 35253 4405 35287
rect 4371 35185 4405 35219
rect 4467 35389 4501 35423
rect 4467 35321 4501 35355
rect 4467 35253 4501 35287
rect 4467 35185 4501 35219
rect 4563 35389 4597 35423
rect 4563 35321 4597 35355
rect 4563 35253 4597 35287
rect 4563 35185 4597 35219
rect 4659 35389 4693 35423
rect 4659 35321 4693 35355
rect 4659 35253 4693 35287
rect 4659 35185 4693 35219
rect 4755 35389 4789 35423
rect 4755 35321 4789 35355
rect 4755 35253 4789 35287
rect 4755 35185 4789 35219
rect 4851 35389 4885 35423
rect 4851 35321 4885 35355
rect 4851 35253 4885 35287
rect 4851 35185 4885 35219
rect 4947 35389 4981 35423
rect 4947 35321 4981 35355
rect 4947 35253 4981 35287
rect 4947 35185 4981 35219
rect 5356 35181 5390 35215
rect 5356 35113 5390 35147
rect 5356 35045 5390 35079
rect 5440 35181 5474 35215
rect 5440 35113 5474 35147
rect 5440 35045 5474 35079
rect 313 34098 347 34132
rect 313 34030 347 34064
rect 313 33962 347 33996
rect 313 33894 347 33928
rect 409 34098 443 34132
rect 409 34030 443 34064
rect 409 33962 443 33996
rect 409 33894 443 33928
rect 505 34098 539 34132
rect 505 34030 539 34064
rect 505 33962 539 33996
rect 505 33894 539 33928
rect 601 34098 635 34132
rect 601 34030 635 34064
rect 601 33962 635 33996
rect 601 33894 635 33928
rect 697 34098 731 34132
rect 697 34030 731 34064
rect 697 33962 731 33996
rect 697 33894 731 33928
rect 793 34098 827 34132
rect 793 34030 827 34064
rect 793 33962 827 33996
rect 793 33894 827 33928
rect 889 34098 923 34132
rect 889 34030 923 34064
rect 889 33962 923 33996
rect 889 33894 923 33928
rect 985 34098 1019 34132
rect 985 34030 1019 34064
rect 985 33962 1019 33996
rect 985 33894 1019 33928
rect 1081 34098 1115 34132
rect 1081 34030 1115 34064
rect 1081 33962 1115 33996
rect 1081 33894 1115 33928
rect 1177 34098 1211 34132
rect 1177 34030 1211 34064
rect 1177 33962 1211 33996
rect 1177 33894 1211 33928
rect 1273 34098 1307 34132
rect 1273 34030 1307 34064
rect 1273 33962 1307 33996
rect 1273 33894 1307 33928
rect 2466 34102 2500 34136
rect 2466 34034 2500 34068
rect 2466 33966 2500 34000
rect 2466 33898 2500 33932
rect 2562 34102 2596 34136
rect 2562 34034 2596 34068
rect 2562 33966 2596 34000
rect 2562 33898 2596 33932
rect 2658 34102 2692 34136
rect 2658 34034 2692 34068
rect 2658 33966 2692 34000
rect 2658 33898 2692 33932
rect 2754 34102 2788 34136
rect 2754 34034 2788 34068
rect 2754 33966 2788 34000
rect 2754 33898 2788 33932
rect 2850 34102 2884 34136
rect 2850 34034 2884 34068
rect 2850 33966 2884 34000
rect 2850 33898 2884 33932
rect 2946 34102 2980 34136
rect 2946 34034 2980 34068
rect 2946 33966 2980 34000
rect 2946 33898 2980 33932
rect 3042 34102 3076 34136
rect 3042 34034 3076 34068
rect 3042 33966 3076 34000
rect 3042 33898 3076 33932
rect 3138 34102 3172 34136
rect 3138 34034 3172 34068
rect 3138 33966 3172 34000
rect 3138 33898 3172 33932
rect 3234 34102 3268 34136
rect 3234 34034 3268 34068
rect 3234 33966 3268 34000
rect 3234 33898 3268 33932
rect 3330 34102 3364 34136
rect 3330 34034 3364 34068
rect 3330 33966 3364 34000
rect 3330 33898 3364 33932
rect 3426 34102 3460 34136
rect 3426 34034 3460 34068
rect 3426 33966 3460 34000
rect 3426 33898 3460 33932
rect 3987 34102 4021 34136
rect 3987 34034 4021 34068
rect 3987 33966 4021 34000
rect 3987 33898 4021 33932
rect 4083 34102 4117 34136
rect 4083 34034 4117 34068
rect 4083 33966 4117 34000
rect 4083 33898 4117 33932
rect 4179 34102 4213 34136
rect 4179 34034 4213 34068
rect 4179 33966 4213 34000
rect 4179 33898 4213 33932
rect 4275 34102 4309 34136
rect 4275 34034 4309 34068
rect 4275 33966 4309 34000
rect 4275 33898 4309 33932
rect 4371 34102 4405 34136
rect 4371 34034 4405 34068
rect 4371 33966 4405 34000
rect 4371 33898 4405 33932
rect 4467 34102 4501 34136
rect 4467 34034 4501 34068
rect 4467 33966 4501 34000
rect 4467 33898 4501 33932
rect 4563 34102 4597 34136
rect 4563 34034 4597 34068
rect 4563 33966 4597 34000
rect 4563 33898 4597 33932
rect 4659 34102 4693 34136
rect 4659 34034 4693 34068
rect 4659 33966 4693 34000
rect 4659 33898 4693 33932
rect 4755 34102 4789 34136
rect 4755 34034 4789 34068
rect 4755 33966 4789 34000
rect 4755 33898 4789 33932
rect 4851 34102 4885 34136
rect 4851 34034 4885 34068
rect 4851 33966 4885 34000
rect 4851 33898 4885 33932
rect 4947 34102 4981 34136
rect 4947 34034 4981 34068
rect 4947 33966 4981 34000
rect 4947 33898 4981 33932
rect 5356 33894 5390 33928
rect 5356 33826 5390 33860
rect 5356 33758 5390 33792
rect 5440 33894 5474 33928
rect 5440 33826 5474 33860
rect 5440 33758 5474 33792
rect 313 32811 347 32845
rect 313 32743 347 32777
rect 313 32675 347 32709
rect 313 32607 347 32641
rect 409 32811 443 32845
rect 409 32743 443 32777
rect 409 32675 443 32709
rect 409 32607 443 32641
rect 505 32811 539 32845
rect 505 32743 539 32777
rect 505 32675 539 32709
rect 505 32607 539 32641
rect 601 32811 635 32845
rect 601 32743 635 32777
rect 601 32675 635 32709
rect 601 32607 635 32641
rect 697 32811 731 32845
rect 697 32743 731 32777
rect 697 32675 731 32709
rect 697 32607 731 32641
rect 793 32811 827 32845
rect 793 32743 827 32777
rect 793 32675 827 32709
rect 793 32607 827 32641
rect 889 32811 923 32845
rect 889 32743 923 32777
rect 889 32675 923 32709
rect 889 32607 923 32641
rect 985 32811 1019 32845
rect 985 32743 1019 32777
rect 985 32675 1019 32709
rect 985 32607 1019 32641
rect 1081 32811 1115 32845
rect 1081 32743 1115 32777
rect 1081 32675 1115 32709
rect 1081 32607 1115 32641
rect 1177 32811 1211 32845
rect 1177 32743 1211 32777
rect 1177 32675 1211 32709
rect 1177 32607 1211 32641
rect 1273 32811 1307 32845
rect 1273 32743 1307 32777
rect 1273 32675 1307 32709
rect 1273 32607 1307 32641
rect 2466 32815 2500 32849
rect 2466 32747 2500 32781
rect 2466 32679 2500 32713
rect 2466 32611 2500 32645
rect 2562 32815 2596 32849
rect 2562 32747 2596 32781
rect 2562 32679 2596 32713
rect 2562 32611 2596 32645
rect 2658 32815 2692 32849
rect 2658 32747 2692 32781
rect 2658 32679 2692 32713
rect 2658 32611 2692 32645
rect 2754 32815 2788 32849
rect 2754 32747 2788 32781
rect 2754 32679 2788 32713
rect 2754 32611 2788 32645
rect 2850 32815 2884 32849
rect 2850 32747 2884 32781
rect 2850 32679 2884 32713
rect 2850 32611 2884 32645
rect 2946 32815 2980 32849
rect 2946 32747 2980 32781
rect 2946 32679 2980 32713
rect 2946 32611 2980 32645
rect 3042 32815 3076 32849
rect 3042 32747 3076 32781
rect 3042 32679 3076 32713
rect 3042 32611 3076 32645
rect 3138 32815 3172 32849
rect 3138 32747 3172 32781
rect 3138 32679 3172 32713
rect 3138 32611 3172 32645
rect 3234 32815 3268 32849
rect 3234 32747 3268 32781
rect 3234 32679 3268 32713
rect 3234 32611 3268 32645
rect 3330 32815 3364 32849
rect 3330 32747 3364 32781
rect 3330 32679 3364 32713
rect 3330 32611 3364 32645
rect 3426 32815 3460 32849
rect 3426 32747 3460 32781
rect 3426 32679 3460 32713
rect 3426 32611 3460 32645
rect 3987 32815 4021 32849
rect 3987 32747 4021 32781
rect 3987 32679 4021 32713
rect 3987 32611 4021 32645
rect 4083 32815 4117 32849
rect 4083 32747 4117 32781
rect 4083 32679 4117 32713
rect 4083 32611 4117 32645
rect 4179 32815 4213 32849
rect 4179 32747 4213 32781
rect 4179 32679 4213 32713
rect 4179 32611 4213 32645
rect 4275 32815 4309 32849
rect 4275 32747 4309 32781
rect 4275 32679 4309 32713
rect 4275 32611 4309 32645
rect 4371 32815 4405 32849
rect 4371 32747 4405 32781
rect 4371 32679 4405 32713
rect 4371 32611 4405 32645
rect 4467 32815 4501 32849
rect 4467 32747 4501 32781
rect 4467 32679 4501 32713
rect 4467 32611 4501 32645
rect 4563 32815 4597 32849
rect 4563 32747 4597 32781
rect 4563 32679 4597 32713
rect 4563 32611 4597 32645
rect 4659 32815 4693 32849
rect 4659 32747 4693 32781
rect 4659 32679 4693 32713
rect 4659 32611 4693 32645
rect 4755 32815 4789 32849
rect 4755 32747 4789 32781
rect 4755 32679 4789 32713
rect 4755 32611 4789 32645
rect 4851 32815 4885 32849
rect 4851 32747 4885 32781
rect 4851 32679 4885 32713
rect 4851 32611 4885 32645
rect 4947 32815 4981 32849
rect 4947 32747 4981 32781
rect 4947 32679 4981 32713
rect 4947 32611 4981 32645
rect 5356 32607 5390 32641
rect 5356 32539 5390 32573
rect 5356 32471 5390 32505
rect 5440 32607 5474 32641
rect 5440 32539 5474 32573
rect 5440 32471 5474 32505
rect 313 31524 347 31558
rect 313 31456 347 31490
rect 313 31388 347 31422
rect 313 31320 347 31354
rect 409 31524 443 31558
rect 409 31456 443 31490
rect 409 31388 443 31422
rect 409 31320 443 31354
rect 505 31524 539 31558
rect 505 31456 539 31490
rect 505 31388 539 31422
rect 505 31320 539 31354
rect 601 31524 635 31558
rect 601 31456 635 31490
rect 601 31388 635 31422
rect 601 31320 635 31354
rect 697 31524 731 31558
rect 697 31456 731 31490
rect 697 31388 731 31422
rect 697 31320 731 31354
rect 793 31524 827 31558
rect 793 31456 827 31490
rect 793 31388 827 31422
rect 793 31320 827 31354
rect 889 31524 923 31558
rect 889 31456 923 31490
rect 889 31388 923 31422
rect 889 31320 923 31354
rect 985 31524 1019 31558
rect 985 31456 1019 31490
rect 985 31388 1019 31422
rect 985 31320 1019 31354
rect 1081 31524 1115 31558
rect 1081 31456 1115 31490
rect 1081 31388 1115 31422
rect 1081 31320 1115 31354
rect 1177 31524 1211 31558
rect 1177 31456 1211 31490
rect 1177 31388 1211 31422
rect 1177 31320 1211 31354
rect 1273 31524 1307 31558
rect 1273 31456 1307 31490
rect 1273 31388 1307 31422
rect 1273 31320 1307 31354
rect 2466 31528 2500 31562
rect 2466 31460 2500 31494
rect 2466 31392 2500 31426
rect 2466 31324 2500 31358
rect 2562 31528 2596 31562
rect 2562 31460 2596 31494
rect 2562 31392 2596 31426
rect 2562 31324 2596 31358
rect 2658 31528 2692 31562
rect 2658 31460 2692 31494
rect 2658 31392 2692 31426
rect 2658 31324 2692 31358
rect 2754 31528 2788 31562
rect 2754 31460 2788 31494
rect 2754 31392 2788 31426
rect 2754 31324 2788 31358
rect 2850 31528 2884 31562
rect 2850 31460 2884 31494
rect 2850 31392 2884 31426
rect 2850 31324 2884 31358
rect 2946 31528 2980 31562
rect 2946 31460 2980 31494
rect 2946 31392 2980 31426
rect 2946 31324 2980 31358
rect 3042 31528 3076 31562
rect 3042 31460 3076 31494
rect 3042 31392 3076 31426
rect 3042 31324 3076 31358
rect 3138 31528 3172 31562
rect 3138 31460 3172 31494
rect 3138 31392 3172 31426
rect 3138 31324 3172 31358
rect 3234 31528 3268 31562
rect 3234 31460 3268 31494
rect 3234 31392 3268 31426
rect 3234 31324 3268 31358
rect 3330 31528 3364 31562
rect 3330 31460 3364 31494
rect 3330 31392 3364 31426
rect 3330 31324 3364 31358
rect 3426 31528 3460 31562
rect 3426 31460 3460 31494
rect 3426 31392 3460 31426
rect 3426 31324 3460 31358
rect 3987 31528 4021 31562
rect 3987 31460 4021 31494
rect 3987 31392 4021 31426
rect 3987 31324 4021 31358
rect 4083 31528 4117 31562
rect 4083 31460 4117 31494
rect 4083 31392 4117 31426
rect 4083 31324 4117 31358
rect 4179 31528 4213 31562
rect 4179 31460 4213 31494
rect 4179 31392 4213 31426
rect 4179 31324 4213 31358
rect 4275 31528 4309 31562
rect 4275 31460 4309 31494
rect 4275 31392 4309 31426
rect 4275 31324 4309 31358
rect 4371 31528 4405 31562
rect 4371 31460 4405 31494
rect 4371 31392 4405 31426
rect 4371 31324 4405 31358
rect 4467 31528 4501 31562
rect 4467 31460 4501 31494
rect 4467 31392 4501 31426
rect 4467 31324 4501 31358
rect 4563 31528 4597 31562
rect 4563 31460 4597 31494
rect 4563 31392 4597 31426
rect 4563 31324 4597 31358
rect 4659 31528 4693 31562
rect 4659 31460 4693 31494
rect 4659 31392 4693 31426
rect 4659 31324 4693 31358
rect 4755 31528 4789 31562
rect 4755 31460 4789 31494
rect 4755 31392 4789 31426
rect 4755 31324 4789 31358
rect 4851 31528 4885 31562
rect 4851 31460 4885 31494
rect 4851 31392 4885 31426
rect 4851 31324 4885 31358
rect 4947 31528 4981 31562
rect 4947 31460 4981 31494
rect 4947 31392 4981 31426
rect 4947 31324 4981 31358
rect 5356 31320 5390 31354
rect 5356 31252 5390 31286
rect 5356 31184 5390 31218
rect 5440 31320 5474 31354
rect 5440 31252 5474 31286
rect 5440 31184 5474 31218
rect 313 30237 347 30271
rect 313 30169 347 30203
rect 313 30101 347 30135
rect 313 30033 347 30067
rect 409 30237 443 30271
rect 409 30169 443 30203
rect 409 30101 443 30135
rect 409 30033 443 30067
rect 505 30237 539 30271
rect 505 30169 539 30203
rect 505 30101 539 30135
rect 505 30033 539 30067
rect 601 30237 635 30271
rect 601 30169 635 30203
rect 601 30101 635 30135
rect 601 30033 635 30067
rect 697 30237 731 30271
rect 697 30169 731 30203
rect 697 30101 731 30135
rect 697 30033 731 30067
rect 793 30237 827 30271
rect 793 30169 827 30203
rect 793 30101 827 30135
rect 793 30033 827 30067
rect 889 30237 923 30271
rect 889 30169 923 30203
rect 889 30101 923 30135
rect 889 30033 923 30067
rect 985 30237 1019 30271
rect 985 30169 1019 30203
rect 985 30101 1019 30135
rect 985 30033 1019 30067
rect 1081 30237 1115 30271
rect 1081 30169 1115 30203
rect 1081 30101 1115 30135
rect 1081 30033 1115 30067
rect 1177 30237 1211 30271
rect 1177 30169 1211 30203
rect 1177 30101 1211 30135
rect 1177 30033 1211 30067
rect 1273 30237 1307 30271
rect 1273 30169 1307 30203
rect 1273 30101 1307 30135
rect 1273 30033 1307 30067
rect 2466 30241 2500 30275
rect 2466 30173 2500 30207
rect 2466 30105 2500 30139
rect 2466 30037 2500 30071
rect 2562 30241 2596 30275
rect 2562 30173 2596 30207
rect 2562 30105 2596 30139
rect 2562 30037 2596 30071
rect 2658 30241 2692 30275
rect 2658 30173 2692 30207
rect 2658 30105 2692 30139
rect 2658 30037 2692 30071
rect 2754 30241 2788 30275
rect 2754 30173 2788 30207
rect 2754 30105 2788 30139
rect 2754 30037 2788 30071
rect 2850 30241 2884 30275
rect 2850 30173 2884 30207
rect 2850 30105 2884 30139
rect 2850 30037 2884 30071
rect 2946 30241 2980 30275
rect 2946 30173 2980 30207
rect 2946 30105 2980 30139
rect 2946 30037 2980 30071
rect 3042 30241 3076 30275
rect 3042 30173 3076 30207
rect 3042 30105 3076 30139
rect 3042 30037 3076 30071
rect 3138 30241 3172 30275
rect 3138 30173 3172 30207
rect 3138 30105 3172 30139
rect 3138 30037 3172 30071
rect 3234 30241 3268 30275
rect 3234 30173 3268 30207
rect 3234 30105 3268 30139
rect 3234 30037 3268 30071
rect 3330 30241 3364 30275
rect 3330 30173 3364 30207
rect 3330 30105 3364 30139
rect 3330 30037 3364 30071
rect 3426 30241 3460 30275
rect 3426 30173 3460 30207
rect 3426 30105 3460 30139
rect 3426 30037 3460 30071
rect 3987 30241 4021 30275
rect 3987 30173 4021 30207
rect 3987 30105 4021 30139
rect 3987 30037 4021 30071
rect 4083 30241 4117 30275
rect 4083 30173 4117 30207
rect 4083 30105 4117 30139
rect 4083 30037 4117 30071
rect 4179 30241 4213 30275
rect 4179 30173 4213 30207
rect 4179 30105 4213 30139
rect 4179 30037 4213 30071
rect 4275 30241 4309 30275
rect 4275 30173 4309 30207
rect 4275 30105 4309 30139
rect 4275 30037 4309 30071
rect 4371 30241 4405 30275
rect 4371 30173 4405 30207
rect 4371 30105 4405 30139
rect 4371 30037 4405 30071
rect 4467 30241 4501 30275
rect 4467 30173 4501 30207
rect 4467 30105 4501 30139
rect 4467 30037 4501 30071
rect 4563 30241 4597 30275
rect 4563 30173 4597 30207
rect 4563 30105 4597 30139
rect 4563 30037 4597 30071
rect 4659 30241 4693 30275
rect 4659 30173 4693 30207
rect 4659 30105 4693 30139
rect 4659 30037 4693 30071
rect 4755 30241 4789 30275
rect 4755 30173 4789 30207
rect 4755 30105 4789 30139
rect 4755 30037 4789 30071
rect 4851 30241 4885 30275
rect 4851 30173 4885 30207
rect 4851 30105 4885 30139
rect 4851 30037 4885 30071
rect 4947 30241 4981 30275
rect 4947 30173 4981 30207
rect 4947 30105 4981 30139
rect 4947 30037 4981 30071
rect 5356 30033 5390 30067
rect 5356 29965 5390 29999
rect 5356 29897 5390 29931
rect 5440 30033 5474 30067
rect 5440 29965 5474 29999
rect 5440 29897 5474 29931
rect 313 28950 347 28984
rect 313 28882 347 28916
rect 313 28814 347 28848
rect 313 28746 347 28780
rect 409 28950 443 28984
rect 409 28882 443 28916
rect 409 28814 443 28848
rect 409 28746 443 28780
rect 505 28950 539 28984
rect 505 28882 539 28916
rect 505 28814 539 28848
rect 505 28746 539 28780
rect 601 28950 635 28984
rect 601 28882 635 28916
rect 601 28814 635 28848
rect 601 28746 635 28780
rect 697 28950 731 28984
rect 697 28882 731 28916
rect 697 28814 731 28848
rect 697 28746 731 28780
rect 793 28950 827 28984
rect 793 28882 827 28916
rect 793 28814 827 28848
rect 793 28746 827 28780
rect 889 28950 923 28984
rect 889 28882 923 28916
rect 889 28814 923 28848
rect 889 28746 923 28780
rect 985 28950 1019 28984
rect 985 28882 1019 28916
rect 985 28814 1019 28848
rect 985 28746 1019 28780
rect 1081 28950 1115 28984
rect 1081 28882 1115 28916
rect 1081 28814 1115 28848
rect 1081 28746 1115 28780
rect 1177 28950 1211 28984
rect 1177 28882 1211 28916
rect 1177 28814 1211 28848
rect 1177 28746 1211 28780
rect 1273 28950 1307 28984
rect 1273 28882 1307 28916
rect 1273 28814 1307 28848
rect 1273 28746 1307 28780
rect 2466 28954 2500 28988
rect 2466 28886 2500 28920
rect 2466 28818 2500 28852
rect 2466 28750 2500 28784
rect 2562 28954 2596 28988
rect 2562 28886 2596 28920
rect 2562 28818 2596 28852
rect 2562 28750 2596 28784
rect 2658 28954 2692 28988
rect 2658 28886 2692 28920
rect 2658 28818 2692 28852
rect 2658 28750 2692 28784
rect 2754 28954 2788 28988
rect 2754 28886 2788 28920
rect 2754 28818 2788 28852
rect 2754 28750 2788 28784
rect 2850 28954 2884 28988
rect 2850 28886 2884 28920
rect 2850 28818 2884 28852
rect 2850 28750 2884 28784
rect 2946 28954 2980 28988
rect 2946 28886 2980 28920
rect 2946 28818 2980 28852
rect 2946 28750 2980 28784
rect 3042 28954 3076 28988
rect 3042 28886 3076 28920
rect 3042 28818 3076 28852
rect 3042 28750 3076 28784
rect 3138 28954 3172 28988
rect 3138 28886 3172 28920
rect 3138 28818 3172 28852
rect 3138 28750 3172 28784
rect 3234 28954 3268 28988
rect 3234 28886 3268 28920
rect 3234 28818 3268 28852
rect 3234 28750 3268 28784
rect 3330 28954 3364 28988
rect 3330 28886 3364 28920
rect 3330 28818 3364 28852
rect 3330 28750 3364 28784
rect 3426 28954 3460 28988
rect 3426 28886 3460 28920
rect 3426 28818 3460 28852
rect 3426 28750 3460 28784
rect 3987 28954 4021 28988
rect 3987 28886 4021 28920
rect 3987 28818 4021 28852
rect 3987 28750 4021 28784
rect 4083 28954 4117 28988
rect 4083 28886 4117 28920
rect 4083 28818 4117 28852
rect 4083 28750 4117 28784
rect 4179 28954 4213 28988
rect 4179 28886 4213 28920
rect 4179 28818 4213 28852
rect 4179 28750 4213 28784
rect 4275 28954 4309 28988
rect 4275 28886 4309 28920
rect 4275 28818 4309 28852
rect 4275 28750 4309 28784
rect 4371 28954 4405 28988
rect 4371 28886 4405 28920
rect 4371 28818 4405 28852
rect 4371 28750 4405 28784
rect 4467 28954 4501 28988
rect 4467 28886 4501 28920
rect 4467 28818 4501 28852
rect 4467 28750 4501 28784
rect 4563 28954 4597 28988
rect 4563 28886 4597 28920
rect 4563 28818 4597 28852
rect 4563 28750 4597 28784
rect 4659 28954 4693 28988
rect 4659 28886 4693 28920
rect 4659 28818 4693 28852
rect 4659 28750 4693 28784
rect 4755 28954 4789 28988
rect 4755 28886 4789 28920
rect 4755 28818 4789 28852
rect 4755 28750 4789 28784
rect 4851 28954 4885 28988
rect 4851 28886 4885 28920
rect 4851 28818 4885 28852
rect 4851 28750 4885 28784
rect 4947 28954 4981 28988
rect 4947 28886 4981 28920
rect 4947 28818 4981 28852
rect 4947 28750 4981 28784
rect 5356 28746 5390 28780
rect 5356 28678 5390 28712
rect 5356 28610 5390 28644
rect 5440 28746 5474 28780
rect 5440 28678 5474 28712
rect 5440 28610 5474 28644
rect 313 27663 347 27697
rect 313 27595 347 27629
rect 313 27527 347 27561
rect 313 27459 347 27493
rect 409 27663 443 27697
rect 409 27595 443 27629
rect 409 27527 443 27561
rect 409 27459 443 27493
rect 505 27663 539 27697
rect 505 27595 539 27629
rect 505 27527 539 27561
rect 505 27459 539 27493
rect 601 27663 635 27697
rect 601 27595 635 27629
rect 601 27527 635 27561
rect 601 27459 635 27493
rect 697 27663 731 27697
rect 697 27595 731 27629
rect 697 27527 731 27561
rect 697 27459 731 27493
rect 793 27663 827 27697
rect 793 27595 827 27629
rect 793 27527 827 27561
rect 793 27459 827 27493
rect 889 27663 923 27697
rect 889 27595 923 27629
rect 889 27527 923 27561
rect 889 27459 923 27493
rect 985 27663 1019 27697
rect 985 27595 1019 27629
rect 985 27527 1019 27561
rect 985 27459 1019 27493
rect 1081 27663 1115 27697
rect 1081 27595 1115 27629
rect 1081 27527 1115 27561
rect 1081 27459 1115 27493
rect 1177 27663 1211 27697
rect 1177 27595 1211 27629
rect 1177 27527 1211 27561
rect 1177 27459 1211 27493
rect 1273 27663 1307 27697
rect 1273 27595 1307 27629
rect 1273 27527 1307 27561
rect 1273 27459 1307 27493
rect 2466 27667 2500 27701
rect 2466 27599 2500 27633
rect 2466 27531 2500 27565
rect 2466 27463 2500 27497
rect 2562 27667 2596 27701
rect 2562 27599 2596 27633
rect 2562 27531 2596 27565
rect 2562 27463 2596 27497
rect 2658 27667 2692 27701
rect 2658 27599 2692 27633
rect 2658 27531 2692 27565
rect 2658 27463 2692 27497
rect 2754 27667 2788 27701
rect 2754 27599 2788 27633
rect 2754 27531 2788 27565
rect 2754 27463 2788 27497
rect 2850 27667 2884 27701
rect 2850 27599 2884 27633
rect 2850 27531 2884 27565
rect 2850 27463 2884 27497
rect 2946 27667 2980 27701
rect 2946 27599 2980 27633
rect 2946 27531 2980 27565
rect 2946 27463 2980 27497
rect 3042 27667 3076 27701
rect 3042 27599 3076 27633
rect 3042 27531 3076 27565
rect 3042 27463 3076 27497
rect 3138 27667 3172 27701
rect 3138 27599 3172 27633
rect 3138 27531 3172 27565
rect 3138 27463 3172 27497
rect 3234 27667 3268 27701
rect 3234 27599 3268 27633
rect 3234 27531 3268 27565
rect 3234 27463 3268 27497
rect 3330 27667 3364 27701
rect 3330 27599 3364 27633
rect 3330 27531 3364 27565
rect 3330 27463 3364 27497
rect 3426 27667 3460 27701
rect 3426 27599 3460 27633
rect 3426 27531 3460 27565
rect 3426 27463 3460 27497
rect 3987 27667 4021 27701
rect 3987 27599 4021 27633
rect 3987 27531 4021 27565
rect 3987 27463 4021 27497
rect 4083 27667 4117 27701
rect 4083 27599 4117 27633
rect 4083 27531 4117 27565
rect 4083 27463 4117 27497
rect 4179 27667 4213 27701
rect 4179 27599 4213 27633
rect 4179 27531 4213 27565
rect 4179 27463 4213 27497
rect 4275 27667 4309 27701
rect 4275 27599 4309 27633
rect 4275 27531 4309 27565
rect 4275 27463 4309 27497
rect 4371 27667 4405 27701
rect 4371 27599 4405 27633
rect 4371 27531 4405 27565
rect 4371 27463 4405 27497
rect 4467 27667 4501 27701
rect 4467 27599 4501 27633
rect 4467 27531 4501 27565
rect 4467 27463 4501 27497
rect 4563 27667 4597 27701
rect 4563 27599 4597 27633
rect 4563 27531 4597 27565
rect 4563 27463 4597 27497
rect 4659 27667 4693 27701
rect 4659 27599 4693 27633
rect 4659 27531 4693 27565
rect 4659 27463 4693 27497
rect 4755 27667 4789 27701
rect 4755 27599 4789 27633
rect 4755 27531 4789 27565
rect 4755 27463 4789 27497
rect 4851 27667 4885 27701
rect 4851 27599 4885 27633
rect 4851 27531 4885 27565
rect 4851 27463 4885 27497
rect 4947 27667 4981 27701
rect 4947 27599 4981 27633
rect 4947 27531 4981 27565
rect 4947 27463 4981 27497
rect 5356 27459 5390 27493
rect 5356 27391 5390 27425
rect 5356 27323 5390 27357
rect 5440 27459 5474 27493
rect 5440 27391 5474 27425
rect 5440 27323 5474 27357
rect 313 26376 347 26410
rect 313 26308 347 26342
rect 313 26240 347 26274
rect 313 26172 347 26206
rect 409 26376 443 26410
rect 409 26308 443 26342
rect 409 26240 443 26274
rect 409 26172 443 26206
rect 505 26376 539 26410
rect 505 26308 539 26342
rect 505 26240 539 26274
rect 505 26172 539 26206
rect 601 26376 635 26410
rect 601 26308 635 26342
rect 601 26240 635 26274
rect 601 26172 635 26206
rect 697 26376 731 26410
rect 697 26308 731 26342
rect 697 26240 731 26274
rect 697 26172 731 26206
rect 793 26376 827 26410
rect 793 26308 827 26342
rect 793 26240 827 26274
rect 793 26172 827 26206
rect 889 26376 923 26410
rect 889 26308 923 26342
rect 889 26240 923 26274
rect 889 26172 923 26206
rect 985 26376 1019 26410
rect 985 26308 1019 26342
rect 985 26240 1019 26274
rect 985 26172 1019 26206
rect 1081 26376 1115 26410
rect 1081 26308 1115 26342
rect 1081 26240 1115 26274
rect 1081 26172 1115 26206
rect 1177 26376 1211 26410
rect 1177 26308 1211 26342
rect 1177 26240 1211 26274
rect 1177 26172 1211 26206
rect 1273 26376 1307 26410
rect 1273 26308 1307 26342
rect 1273 26240 1307 26274
rect 1273 26172 1307 26206
rect 2466 26380 2500 26414
rect 2466 26312 2500 26346
rect 2466 26244 2500 26278
rect 2466 26176 2500 26210
rect 2562 26380 2596 26414
rect 2562 26312 2596 26346
rect 2562 26244 2596 26278
rect 2562 26176 2596 26210
rect 2658 26380 2692 26414
rect 2658 26312 2692 26346
rect 2658 26244 2692 26278
rect 2658 26176 2692 26210
rect 2754 26380 2788 26414
rect 2754 26312 2788 26346
rect 2754 26244 2788 26278
rect 2754 26176 2788 26210
rect 2850 26380 2884 26414
rect 2850 26312 2884 26346
rect 2850 26244 2884 26278
rect 2850 26176 2884 26210
rect 2946 26380 2980 26414
rect 2946 26312 2980 26346
rect 2946 26244 2980 26278
rect 2946 26176 2980 26210
rect 3042 26380 3076 26414
rect 3042 26312 3076 26346
rect 3042 26244 3076 26278
rect 3042 26176 3076 26210
rect 3138 26380 3172 26414
rect 3138 26312 3172 26346
rect 3138 26244 3172 26278
rect 3138 26176 3172 26210
rect 3234 26380 3268 26414
rect 3234 26312 3268 26346
rect 3234 26244 3268 26278
rect 3234 26176 3268 26210
rect 3330 26380 3364 26414
rect 3330 26312 3364 26346
rect 3330 26244 3364 26278
rect 3330 26176 3364 26210
rect 3426 26380 3460 26414
rect 3426 26312 3460 26346
rect 3426 26244 3460 26278
rect 3426 26176 3460 26210
rect 3987 26380 4021 26414
rect 3987 26312 4021 26346
rect 3987 26244 4021 26278
rect 3987 26176 4021 26210
rect 4083 26380 4117 26414
rect 4083 26312 4117 26346
rect 4083 26244 4117 26278
rect 4083 26176 4117 26210
rect 4179 26380 4213 26414
rect 4179 26312 4213 26346
rect 4179 26244 4213 26278
rect 4179 26176 4213 26210
rect 4275 26380 4309 26414
rect 4275 26312 4309 26346
rect 4275 26244 4309 26278
rect 4275 26176 4309 26210
rect 4371 26380 4405 26414
rect 4371 26312 4405 26346
rect 4371 26244 4405 26278
rect 4371 26176 4405 26210
rect 4467 26380 4501 26414
rect 4467 26312 4501 26346
rect 4467 26244 4501 26278
rect 4467 26176 4501 26210
rect 4563 26380 4597 26414
rect 4563 26312 4597 26346
rect 4563 26244 4597 26278
rect 4563 26176 4597 26210
rect 4659 26380 4693 26414
rect 4659 26312 4693 26346
rect 4659 26244 4693 26278
rect 4659 26176 4693 26210
rect 4755 26380 4789 26414
rect 4755 26312 4789 26346
rect 4755 26244 4789 26278
rect 4755 26176 4789 26210
rect 4851 26380 4885 26414
rect 4851 26312 4885 26346
rect 4851 26244 4885 26278
rect 4851 26176 4885 26210
rect 4947 26380 4981 26414
rect 4947 26312 4981 26346
rect 4947 26244 4981 26278
rect 4947 26176 4981 26210
rect 5356 26172 5390 26206
rect 5356 26104 5390 26138
rect 5356 26036 5390 26070
rect 5440 26172 5474 26206
rect 5440 26104 5474 26138
rect 5440 26036 5474 26070
rect 313 25089 347 25123
rect 313 25021 347 25055
rect 313 24953 347 24987
rect 313 24885 347 24919
rect 409 25089 443 25123
rect 409 25021 443 25055
rect 409 24953 443 24987
rect 409 24885 443 24919
rect 505 25089 539 25123
rect 505 25021 539 25055
rect 505 24953 539 24987
rect 505 24885 539 24919
rect 601 25089 635 25123
rect 601 25021 635 25055
rect 601 24953 635 24987
rect 601 24885 635 24919
rect 697 25089 731 25123
rect 697 25021 731 25055
rect 697 24953 731 24987
rect 697 24885 731 24919
rect 793 25089 827 25123
rect 793 25021 827 25055
rect 793 24953 827 24987
rect 793 24885 827 24919
rect 889 25089 923 25123
rect 889 25021 923 25055
rect 889 24953 923 24987
rect 889 24885 923 24919
rect 985 25089 1019 25123
rect 985 25021 1019 25055
rect 985 24953 1019 24987
rect 985 24885 1019 24919
rect 1081 25089 1115 25123
rect 1081 25021 1115 25055
rect 1081 24953 1115 24987
rect 1081 24885 1115 24919
rect 1177 25089 1211 25123
rect 1177 25021 1211 25055
rect 1177 24953 1211 24987
rect 1177 24885 1211 24919
rect 1273 25089 1307 25123
rect 1273 25021 1307 25055
rect 1273 24953 1307 24987
rect 1273 24885 1307 24919
rect 2466 25093 2500 25127
rect 2466 25025 2500 25059
rect 2466 24957 2500 24991
rect 2466 24889 2500 24923
rect 2562 25093 2596 25127
rect 2562 25025 2596 25059
rect 2562 24957 2596 24991
rect 2562 24889 2596 24923
rect 2658 25093 2692 25127
rect 2658 25025 2692 25059
rect 2658 24957 2692 24991
rect 2658 24889 2692 24923
rect 2754 25093 2788 25127
rect 2754 25025 2788 25059
rect 2754 24957 2788 24991
rect 2754 24889 2788 24923
rect 2850 25093 2884 25127
rect 2850 25025 2884 25059
rect 2850 24957 2884 24991
rect 2850 24889 2884 24923
rect 2946 25093 2980 25127
rect 2946 25025 2980 25059
rect 2946 24957 2980 24991
rect 2946 24889 2980 24923
rect 3042 25093 3076 25127
rect 3042 25025 3076 25059
rect 3042 24957 3076 24991
rect 3042 24889 3076 24923
rect 3138 25093 3172 25127
rect 3138 25025 3172 25059
rect 3138 24957 3172 24991
rect 3138 24889 3172 24923
rect 3234 25093 3268 25127
rect 3234 25025 3268 25059
rect 3234 24957 3268 24991
rect 3234 24889 3268 24923
rect 3330 25093 3364 25127
rect 3330 25025 3364 25059
rect 3330 24957 3364 24991
rect 3330 24889 3364 24923
rect 3426 25093 3460 25127
rect 3426 25025 3460 25059
rect 3426 24957 3460 24991
rect 3426 24889 3460 24923
rect 3987 25093 4021 25127
rect 3987 25025 4021 25059
rect 3987 24957 4021 24991
rect 3987 24889 4021 24923
rect 4083 25093 4117 25127
rect 4083 25025 4117 25059
rect 4083 24957 4117 24991
rect 4083 24889 4117 24923
rect 4179 25093 4213 25127
rect 4179 25025 4213 25059
rect 4179 24957 4213 24991
rect 4179 24889 4213 24923
rect 4275 25093 4309 25127
rect 4275 25025 4309 25059
rect 4275 24957 4309 24991
rect 4275 24889 4309 24923
rect 4371 25093 4405 25127
rect 4371 25025 4405 25059
rect 4371 24957 4405 24991
rect 4371 24889 4405 24923
rect 4467 25093 4501 25127
rect 4467 25025 4501 25059
rect 4467 24957 4501 24991
rect 4467 24889 4501 24923
rect 4563 25093 4597 25127
rect 4563 25025 4597 25059
rect 4563 24957 4597 24991
rect 4563 24889 4597 24923
rect 4659 25093 4693 25127
rect 4659 25025 4693 25059
rect 4659 24957 4693 24991
rect 4659 24889 4693 24923
rect 4755 25093 4789 25127
rect 4755 25025 4789 25059
rect 4755 24957 4789 24991
rect 4755 24889 4789 24923
rect 4851 25093 4885 25127
rect 4851 25025 4885 25059
rect 4851 24957 4885 24991
rect 4851 24889 4885 24923
rect 4947 25093 4981 25127
rect 4947 25025 4981 25059
rect 4947 24957 4981 24991
rect 4947 24889 4981 24923
rect 5356 24885 5390 24919
rect 5356 24817 5390 24851
rect 5356 24749 5390 24783
rect 5440 24885 5474 24919
rect 5440 24817 5474 24851
rect 5440 24749 5474 24783
rect 313 23802 347 23836
rect 313 23734 347 23768
rect 313 23666 347 23700
rect 313 23598 347 23632
rect 409 23802 443 23836
rect 409 23734 443 23768
rect 409 23666 443 23700
rect 409 23598 443 23632
rect 505 23802 539 23836
rect 505 23734 539 23768
rect 505 23666 539 23700
rect 505 23598 539 23632
rect 601 23802 635 23836
rect 601 23734 635 23768
rect 601 23666 635 23700
rect 601 23598 635 23632
rect 697 23802 731 23836
rect 697 23734 731 23768
rect 697 23666 731 23700
rect 697 23598 731 23632
rect 793 23802 827 23836
rect 793 23734 827 23768
rect 793 23666 827 23700
rect 793 23598 827 23632
rect 889 23802 923 23836
rect 889 23734 923 23768
rect 889 23666 923 23700
rect 889 23598 923 23632
rect 985 23802 1019 23836
rect 985 23734 1019 23768
rect 985 23666 1019 23700
rect 985 23598 1019 23632
rect 1081 23802 1115 23836
rect 1081 23734 1115 23768
rect 1081 23666 1115 23700
rect 1081 23598 1115 23632
rect 1177 23802 1211 23836
rect 1177 23734 1211 23768
rect 1177 23666 1211 23700
rect 1177 23598 1211 23632
rect 1273 23802 1307 23836
rect 1273 23734 1307 23768
rect 1273 23666 1307 23700
rect 1273 23598 1307 23632
rect 2466 23806 2500 23840
rect 2466 23738 2500 23772
rect 2466 23670 2500 23704
rect 2466 23602 2500 23636
rect 2562 23806 2596 23840
rect 2562 23738 2596 23772
rect 2562 23670 2596 23704
rect 2562 23602 2596 23636
rect 2658 23806 2692 23840
rect 2658 23738 2692 23772
rect 2658 23670 2692 23704
rect 2658 23602 2692 23636
rect 2754 23806 2788 23840
rect 2754 23738 2788 23772
rect 2754 23670 2788 23704
rect 2754 23602 2788 23636
rect 2850 23806 2884 23840
rect 2850 23738 2884 23772
rect 2850 23670 2884 23704
rect 2850 23602 2884 23636
rect 2946 23806 2980 23840
rect 2946 23738 2980 23772
rect 2946 23670 2980 23704
rect 2946 23602 2980 23636
rect 3042 23806 3076 23840
rect 3042 23738 3076 23772
rect 3042 23670 3076 23704
rect 3042 23602 3076 23636
rect 3138 23806 3172 23840
rect 3138 23738 3172 23772
rect 3138 23670 3172 23704
rect 3138 23602 3172 23636
rect 3234 23806 3268 23840
rect 3234 23738 3268 23772
rect 3234 23670 3268 23704
rect 3234 23602 3268 23636
rect 3330 23806 3364 23840
rect 3330 23738 3364 23772
rect 3330 23670 3364 23704
rect 3330 23602 3364 23636
rect 3426 23806 3460 23840
rect 3426 23738 3460 23772
rect 3426 23670 3460 23704
rect 3426 23602 3460 23636
rect 3987 23806 4021 23840
rect 3987 23738 4021 23772
rect 3987 23670 4021 23704
rect 3987 23602 4021 23636
rect 4083 23806 4117 23840
rect 4083 23738 4117 23772
rect 4083 23670 4117 23704
rect 4083 23602 4117 23636
rect 4179 23806 4213 23840
rect 4179 23738 4213 23772
rect 4179 23670 4213 23704
rect 4179 23602 4213 23636
rect 4275 23806 4309 23840
rect 4275 23738 4309 23772
rect 4275 23670 4309 23704
rect 4275 23602 4309 23636
rect 4371 23806 4405 23840
rect 4371 23738 4405 23772
rect 4371 23670 4405 23704
rect 4371 23602 4405 23636
rect 4467 23806 4501 23840
rect 4467 23738 4501 23772
rect 4467 23670 4501 23704
rect 4467 23602 4501 23636
rect 4563 23806 4597 23840
rect 4563 23738 4597 23772
rect 4563 23670 4597 23704
rect 4563 23602 4597 23636
rect 4659 23806 4693 23840
rect 4659 23738 4693 23772
rect 4659 23670 4693 23704
rect 4659 23602 4693 23636
rect 4755 23806 4789 23840
rect 4755 23738 4789 23772
rect 4755 23670 4789 23704
rect 4755 23602 4789 23636
rect 4851 23806 4885 23840
rect 4851 23738 4885 23772
rect 4851 23670 4885 23704
rect 4851 23602 4885 23636
rect 4947 23806 4981 23840
rect 4947 23738 4981 23772
rect 4947 23670 4981 23704
rect 4947 23602 4981 23636
rect 5356 23598 5390 23632
rect 5356 23530 5390 23564
rect 5356 23462 5390 23496
rect 5440 23598 5474 23632
rect 5440 23530 5474 23564
rect 5440 23462 5474 23496
rect 313 22515 347 22549
rect 313 22447 347 22481
rect 313 22379 347 22413
rect 313 22311 347 22345
rect 409 22515 443 22549
rect 409 22447 443 22481
rect 409 22379 443 22413
rect 409 22311 443 22345
rect 505 22515 539 22549
rect 505 22447 539 22481
rect 505 22379 539 22413
rect 505 22311 539 22345
rect 601 22515 635 22549
rect 601 22447 635 22481
rect 601 22379 635 22413
rect 601 22311 635 22345
rect 697 22515 731 22549
rect 697 22447 731 22481
rect 697 22379 731 22413
rect 697 22311 731 22345
rect 793 22515 827 22549
rect 793 22447 827 22481
rect 793 22379 827 22413
rect 793 22311 827 22345
rect 889 22515 923 22549
rect 889 22447 923 22481
rect 889 22379 923 22413
rect 889 22311 923 22345
rect 985 22515 1019 22549
rect 985 22447 1019 22481
rect 985 22379 1019 22413
rect 985 22311 1019 22345
rect 1081 22515 1115 22549
rect 1081 22447 1115 22481
rect 1081 22379 1115 22413
rect 1081 22311 1115 22345
rect 1177 22515 1211 22549
rect 1177 22447 1211 22481
rect 1177 22379 1211 22413
rect 1177 22311 1211 22345
rect 1273 22515 1307 22549
rect 1273 22447 1307 22481
rect 1273 22379 1307 22413
rect 1273 22311 1307 22345
rect 2466 22519 2500 22553
rect 2466 22451 2500 22485
rect 2466 22383 2500 22417
rect 2466 22315 2500 22349
rect 2562 22519 2596 22553
rect 2562 22451 2596 22485
rect 2562 22383 2596 22417
rect 2562 22315 2596 22349
rect 2658 22519 2692 22553
rect 2658 22451 2692 22485
rect 2658 22383 2692 22417
rect 2658 22315 2692 22349
rect 2754 22519 2788 22553
rect 2754 22451 2788 22485
rect 2754 22383 2788 22417
rect 2754 22315 2788 22349
rect 2850 22519 2884 22553
rect 2850 22451 2884 22485
rect 2850 22383 2884 22417
rect 2850 22315 2884 22349
rect 2946 22519 2980 22553
rect 2946 22451 2980 22485
rect 2946 22383 2980 22417
rect 2946 22315 2980 22349
rect 3042 22519 3076 22553
rect 3042 22451 3076 22485
rect 3042 22383 3076 22417
rect 3042 22315 3076 22349
rect 3138 22519 3172 22553
rect 3138 22451 3172 22485
rect 3138 22383 3172 22417
rect 3138 22315 3172 22349
rect 3234 22519 3268 22553
rect 3234 22451 3268 22485
rect 3234 22383 3268 22417
rect 3234 22315 3268 22349
rect 3330 22519 3364 22553
rect 3330 22451 3364 22485
rect 3330 22383 3364 22417
rect 3330 22315 3364 22349
rect 3426 22519 3460 22553
rect 3426 22451 3460 22485
rect 3426 22383 3460 22417
rect 3426 22315 3460 22349
rect 3987 22519 4021 22553
rect 3987 22451 4021 22485
rect 3987 22383 4021 22417
rect 3987 22315 4021 22349
rect 4083 22519 4117 22553
rect 4083 22451 4117 22485
rect 4083 22383 4117 22417
rect 4083 22315 4117 22349
rect 4179 22519 4213 22553
rect 4179 22451 4213 22485
rect 4179 22383 4213 22417
rect 4179 22315 4213 22349
rect 4275 22519 4309 22553
rect 4275 22451 4309 22485
rect 4275 22383 4309 22417
rect 4275 22315 4309 22349
rect 4371 22519 4405 22553
rect 4371 22451 4405 22485
rect 4371 22383 4405 22417
rect 4371 22315 4405 22349
rect 4467 22519 4501 22553
rect 4467 22451 4501 22485
rect 4467 22383 4501 22417
rect 4467 22315 4501 22349
rect 4563 22519 4597 22553
rect 4563 22451 4597 22485
rect 4563 22383 4597 22417
rect 4563 22315 4597 22349
rect 4659 22519 4693 22553
rect 4659 22451 4693 22485
rect 4659 22383 4693 22417
rect 4659 22315 4693 22349
rect 4755 22519 4789 22553
rect 4755 22451 4789 22485
rect 4755 22383 4789 22417
rect 4755 22315 4789 22349
rect 4851 22519 4885 22553
rect 4851 22451 4885 22485
rect 4851 22383 4885 22417
rect 4851 22315 4885 22349
rect 4947 22519 4981 22553
rect 4947 22451 4981 22485
rect 4947 22383 4981 22417
rect 4947 22315 4981 22349
rect 5356 22311 5390 22345
rect 5356 22243 5390 22277
rect 5356 22175 5390 22209
rect 5440 22311 5474 22345
rect 5440 22243 5474 22277
rect 5440 22175 5474 22209
rect 313 21228 347 21262
rect 313 21160 347 21194
rect 313 21092 347 21126
rect 313 21024 347 21058
rect 409 21228 443 21262
rect 409 21160 443 21194
rect 409 21092 443 21126
rect 409 21024 443 21058
rect 505 21228 539 21262
rect 505 21160 539 21194
rect 505 21092 539 21126
rect 505 21024 539 21058
rect 601 21228 635 21262
rect 601 21160 635 21194
rect 601 21092 635 21126
rect 601 21024 635 21058
rect 697 21228 731 21262
rect 697 21160 731 21194
rect 697 21092 731 21126
rect 697 21024 731 21058
rect 793 21228 827 21262
rect 793 21160 827 21194
rect 793 21092 827 21126
rect 793 21024 827 21058
rect 889 21228 923 21262
rect 889 21160 923 21194
rect 889 21092 923 21126
rect 889 21024 923 21058
rect 985 21228 1019 21262
rect 985 21160 1019 21194
rect 985 21092 1019 21126
rect 985 21024 1019 21058
rect 1081 21228 1115 21262
rect 1081 21160 1115 21194
rect 1081 21092 1115 21126
rect 1081 21024 1115 21058
rect 1177 21228 1211 21262
rect 1177 21160 1211 21194
rect 1177 21092 1211 21126
rect 1177 21024 1211 21058
rect 1273 21228 1307 21262
rect 1273 21160 1307 21194
rect 1273 21092 1307 21126
rect 1273 21024 1307 21058
rect 2466 21232 2500 21266
rect 2466 21164 2500 21198
rect 2466 21096 2500 21130
rect 2466 21028 2500 21062
rect 2562 21232 2596 21266
rect 2562 21164 2596 21198
rect 2562 21096 2596 21130
rect 2562 21028 2596 21062
rect 2658 21232 2692 21266
rect 2658 21164 2692 21198
rect 2658 21096 2692 21130
rect 2658 21028 2692 21062
rect 2754 21232 2788 21266
rect 2754 21164 2788 21198
rect 2754 21096 2788 21130
rect 2754 21028 2788 21062
rect 2850 21232 2884 21266
rect 2850 21164 2884 21198
rect 2850 21096 2884 21130
rect 2850 21028 2884 21062
rect 2946 21232 2980 21266
rect 2946 21164 2980 21198
rect 2946 21096 2980 21130
rect 2946 21028 2980 21062
rect 3042 21232 3076 21266
rect 3042 21164 3076 21198
rect 3042 21096 3076 21130
rect 3042 21028 3076 21062
rect 3138 21232 3172 21266
rect 3138 21164 3172 21198
rect 3138 21096 3172 21130
rect 3138 21028 3172 21062
rect 3234 21232 3268 21266
rect 3234 21164 3268 21198
rect 3234 21096 3268 21130
rect 3234 21028 3268 21062
rect 3330 21232 3364 21266
rect 3330 21164 3364 21198
rect 3330 21096 3364 21130
rect 3330 21028 3364 21062
rect 3426 21232 3460 21266
rect 3426 21164 3460 21198
rect 3426 21096 3460 21130
rect 3426 21028 3460 21062
rect 3987 21232 4021 21266
rect 3987 21164 4021 21198
rect 3987 21096 4021 21130
rect 3987 21028 4021 21062
rect 4083 21232 4117 21266
rect 4083 21164 4117 21198
rect 4083 21096 4117 21130
rect 4083 21028 4117 21062
rect 4179 21232 4213 21266
rect 4179 21164 4213 21198
rect 4179 21096 4213 21130
rect 4179 21028 4213 21062
rect 4275 21232 4309 21266
rect 4275 21164 4309 21198
rect 4275 21096 4309 21130
rect 4275 21028 4309 21062
rect 4371 21232 4405 21266
rect 4371 21164 4405 21198
rect 4371 21096 4405 21130
rect 4371 21028 4405 21062
rect 4467 21232 4501 21266
rect 4467 21164 4501 21198
rect 4467 21096 4501 21130
rect 4467 21028 4501 21062
rect 4563 21232 4597 21266
rect 4563 21164 4597 21198
rect 4563 21096 4597 21130
rect 4563 21028 4597 21062
rect 4659 21232 4693 21266
rect 4659 21164 4693 21198
rect 4659 21096 4693 21130
rect 4659 21028 4693 21062
rect 4755 21232 4789 21266
rect 4755 21164 4789 21198
rect 4755 21096 4789 21130
rect 4755 21028 4789 21062
rect 4851 21232 4885 21266
rect 4851 21164 4885 21198
rect 4851 21096 4885 21130
rect 4851 21028 4885 21062
rect 4947 21232 4981 21266
rect 4947 21164 4981 21198
rect 4947 21096 4981 21130
rect 4947 21028 4981 21062
rect 5356 21024 5390 21058
rect 5356 20956 5390 20990
rect 5356 20888 5390 20922
rect 5440 21024 5474 21058
rect 5440 20956 5474 20990
rect 5440 20888 5474 20922
rect 313 19941 347 19975
rect 313 19873 347 19907
rect 313 19805 347 19839
rect 313 19737 347 19771
rect 409 19941 443 19975
rect 409 19873 443 19907
rect 409 19805 443 19839
rect 409 19737 443 19771
rect 505 19941 539 19975
rect 505 19873 539 19907
rect 505 19805 539 19839
rect 505 19737 539 19771
rect 601 19941 635 19975
rect 601 19873 635 19907
rect 601 19805 635 19839
rect 601 19737 635 19771
rect 697 19941 731 19975
rect 697 19873 731 19907
rect 697 19805 731 19839
rect 697 19737 731 19771
rect 793 19941 827 19975
rect 793 19873 827 19907
rect 793 19805 827 19839
rect 793 19737 827 19771
rect 889 19941 923 19975
rect 889 19873 923 19907
rect 889 19805 923 19839
rect 889 19737 923 19771
rect 985 19941 1019 19975
rect 985 19873 1019 19907
rect 985 19805 1019 19839
rect 985 19737 1019 19771
rect 1081 19941 1115 19975
rect 1081 19873 1115 19907
rect 1081 19805 1115 19839
rect 1081 19737 1115 19771
rect 1177 19941 1211 19975
rect 1177 19873 1211 19907
rect 1177 19805 1211 19839
rect 1177 19737 1211 19771
rect 1273 19941 1307 19975
rect 1273 19873 1307 19907
rect 1273 19805 1307 19839
rect 1273 19737 1307 19771
rect 2466 19945 2500 19979
rect 2466 19877 2500 19911
rect 2466 19809 2500 19843
rect 2466 19741 2500 19775
rect 2562 19945 2596 19979
rect 2562 19877 2596 19911
rect 2562 19809 2596 19843
rect 2562 19741 2596 19775
rect 2658 19945 2692 19979
rect 2658 19877 2692 19911
rect 2658 19809 2692 19843
rect 2658 19741 2692 19775
rect 2754 19945 2788 19979
rect 2754 19877 2788 19911
rect 2754 19809 2788 19843
rect 2754 19741 2788 19775
rect 2850 19945 2884 19979
rect 2850 19877 2884 19911
rect 2850 19809 2884 19843
rect 2850 19741 2884 19775
rect 2946 19945 2980 19979
rect 2946 19877 2980 19911
rect 2946 19809 2980 19843
rect 2946 19741 2980 19775
rect 3042 19945 3076 19979
rect 3042 19877 3076 19911
rect 3042 19809 3076 19843
rect 3042 19741 3076 19775
rect 3138 19945 3172 19979
rect 3138 19877 3172 19911
rect 3138 19809 3172 19843
rect 3138 19741 3172 19775
rect 3234 19945 3268 19979
rect 3234 19877 3268 19911
rect 3234 19809 3268 19843
rect 3234 19741 3268 19775
rect 3330 19945 3364 19979
rect 3330 19877 3364 19911
rect 3330 19809 3364 19843
rect 3330 19741 3364 19775
rect 3426 19945 3460 19979
rect 3426 19877 3460 19911
rect 3426 19809 3460 19843
rect 3426 19741 3460 19775
rect 3987 19945 4021 19979
rect 3987 19877 4021 19911
rect 3987 19809 4021 19843
rect 3987 19741 4021 19775
rect 4083 19945 4117 19979
rect 4083 19877 4117 19911
rect 4083 19809 4117 19843
rect 4083 19741 4117 19775
rect 4179 19945 4213 19979
rect 4179 19877 4213 19911
rect 4179 19809 4213 19843
rect 4179 19741 4213 19775
rect 4275 19945 4309 19979
rect 4275 19877 4309 19911
rect 4275 19809 4309 19843
rect 4275 19741 4309 19775
rect 4371 19945 4405 19979
rect 4371 19877 4405 19911
rect 4371 19809 4405 19843
rect 4371 19741 4405 19775
rect 4467 19945 4501 19979
rect 4467 19877 4501 19911
rect 4467 19809 4501 19843
rect 4467 19741 4501 19775
rect 4563 19945 4597 19979
rect 4563 19877 4597 19911
rect 4563 19809 4597 19843
rect 4563 19741 4597 19775
rect 4659 19945 4693 19979
rect 4659 19877 4693 19911
rect 4659 19809 4693 19843
rect 4659 19741 4693 19775
rect 4755 19945 4789 19979
rect 4755 19877 4789 19911
rect 4755 19809 4789 19843
rect 4755 19741 4789 19775
rect 4851 19945 4885 19979
rect 4851 19877 4885 19911
rect 4851 19809 4885 19843
rect 4851 19741 4885 19775
rect 4947 19945 4981 19979
rect 4947 19877 4981 19911
rect 4947 19809 4981 19843
rect 4947 19741 4981 19775
rect 5356 19737 5390 19771
rect 5356 19669 5390 19703
rect 5356 19601 5390 19635
rect 5440 19737 5474 19771
rect 5440 19669 5474 19703
rect 5440 19601 5474 19635
rect 313 18654 347 18688
rect 313 18586 347 18620
rect 313 18518 347 18552
rect 313 18450 347 18484
rect 409 18654 443 18688
rect 409 18586 443 18620
rect 409 18518 443 18552
rect 409 18450 443 18484
rect 505 18654 539 18688
rect 505 18586 539 18620
rect 505 18518 539 18552
rect 505 18450 539 18484
rect 601 18654 635 18688
rect 601 18586 635 18620
rect 601 18518 635 18552
rect 601 18450 635 18484
rect 697 18654 731 18688
rect 697 18586 731 18620
rect 697 18518 731 18552
rect 697 18450 731 18484
rect 793 18654 827 18688
rect 793 18586 827 18620
rect 793 18518 827 18552
rect 793 18450 827 18484
rect 889 18654 923 18688
rect 889 18586 923 18620
rect 889 18518 923 18552
rect 889 18450 923 18484
rect 985 18654 1019 18688
rect 985 18586 1019 18620
rect 985 18518 1019 18552
rect 985 18450 1019 18484
rect 1081 18654 1115 18688
rect 1081 18586 1115 18620
rect 1081 18518 1115 18552
rect 1081 18450 1115 18484
rect 1177 18654 1211 18688
rect 1177 18586 1211 18620
rect 1177 18518 1211 18552
rect 1177 18450 1211 18484
rect 1273 18654 1307 18688
rect 1273 18586 1307 18620
rect 1273 18518 1307 18552
rect 1273 18450 1307 18484
rect 2466 18658 2500 18692
rect 2466 18590 2500 18624
rect 2466 18522 2500 18556
rect 2466 18454 2500 18488
rect 2562 18658 2596 18692
rect 2562 18590 2596 18624
rect 2562 18522 2596 18556
rect 2562 18454 2596 18488
rect 2658 18658 2692 18692
rect 2658 18590 2692 18624
rect 2658 18522 2692 18556
rect 2658 18454 2692 18488
rect 2754 18658 2788 18692
rect 2754 18590 2788 18624
rect 2754 18522 2788 18556
rect 2754 18454 2788 18488
rect 2850 18658 2884 18692
rect 2850 18590 2884 18624
rect 2850 18522 2884 18556
rect 2850 18454 2884 18488
rect 2946 18658 2980 18692
rect 2946 18590 2980 18624
rect 2946 18522 2980 18556
rect 2946 18454 2980 18488
rect 3042 18658 3076 18692
rect 3042 18590 3076 18624
rect 3042 18522 3076 18556
rect 3042 18454 3076 18488
rect 3138 18658 3172 18692
rect 3138 18590 3172 18624
rect 3138 18522 3172 18556
rect 3138 18454 3172 18488
rect 3234 18658 3268 18692
rect 3234 18590 3268 18624
rect 3234 18522 3268 18556
rect 3234 18454 3268 18488
rect 3330 18658 3364 18692
rect 3330 18590 3364 18624
rect 3330 18522 3364 18556
rect 3330 18454 3364 18488
rect 3426 18658 3460 18692
rect 3426 18590 3460 18624
rect 3426 18522 3460 18556
rect 3426 18454 3460 18488
rect 3987 18658 4021 18692
rect 3987 18590 4021 18624
rect 3987 18522 4021 18556
rect 3987 18454 4021 18488
rect 4083 18658 4117 18692
rect 4083 18590 4117 18624
rect 4083 18522 4117 18556
rect 4083 18454 4117 18488
rect 4179 18658 4213 18692
rect 4179 18590 4213 18624
rect 4179 18522 4213 18556
rect 4179 18454 4213 18488
rect 4275 18658 4309 18692
rect 4275 18590 4309 18624
rect 4275 18522 4309 18556
rect 4275 18454 4309 18488
rect 4371 18658 4405 18692
rect 4371 18590 4405 18624
rect 4371 18522 4405 18556
rect 4371 18454 4405 18488
rect 4467 18658 4501 18692
rect 4467 18590 4501 18624
rect 4467 18522 4501 18556
rect 4467 18454 4501 18488
rect 4563 18658 4597 18692
rect 4563 18590 4597 18624
rect 4563 18522 4597 18556
rect 4563 18454 4597 18488
rect 4659 18658 4693 18692
rect 4659 18590 4693 18624
rect 4659 18522 4693 18556
rect 4659 18454 4693 18488
rect 4755 18658 4789 18692
rect 4755 18590 4789 18624
rect 4755 18522 4789 18556
rect 4755 18454 4789 18488
rect 4851 18658 4885 18692
rect 4851 18590 4885 18624
rect 4851 18522 4885 18556
rect 4851 18454 4885 18488
rect 4947 18658 4981 18692
rect 4947 18590 4981 18624
rect 4947 18522 4981 18556
rect 4947 18454 4981 18488
rect 5356 18450 5390 18484
rect 5356 18382 5390 18416
rect 5356 18314 5390 18348
rect 5440 18450 5474 18484
rect 5440 18382 5474 18416
rect 5440 18314 5474 18348
rect 313 17367 347 17401
rect 313 17299 347 17333
rect 313 17231 347 17265
rect 313 17163 347 17197
rect 409 17367 443 17401
rect 409 17299 443 17333
rect 409 17231 443 17265
rect 409 17163 443 17197
rect 505 17367 539 17401
rect 505 17299 539 17333
rect 505 17231 539 17265
rect 505 17163 539 17197
rect 601 17367 635 17401
rect 601 17299 635 17333
rect 601 17231 635 17265
rect 601 17163 635 17197
rect 697 17367 731 17401
rect 697 17299 731 17333
rect 697 17231 731 17265
rect 697 17163 731 17197
rect 793 17367 827 17401
rect 793 17299 827 17333
rect 793 17231 827 17265
rect 793 17163 827 17197
rect 889 17367 923 17401
rect 889 17299 923 17333
rect 889 17231 923 17265
rect 889 17163 923 17197
rect 985 17367 1019 17401
rect 985 17299 1019 17333
rect 985 17231 1019 17265
rect 985 17163 1019 17197
rect 1081 17367 1115 17401
rect 1081 17299 1115 17333
rect 1081 17231 1115 17265
rect 1081 17163 1115 17197
rect 1177 17367 1211 17401
rect 1177 17299 1211 17333
rect 1177 17231 1211 17265
rect 1177 17163 1211 17197
rect 1273 17367 1307 17401
rect 1273 17299 1307 17333
rect 1273 17231 1307 17265
rect 1273 17163 1307 17197
rect 2466 17371 2500 17405
rect 2466 17303 2500 17337
rect 2466 17235 2500 17269
rect 2466 17167 2500 17201
rect 2562 17371 2596 17405
rect 2562 17303 2596 17337
rect 2562 17235 2596 17269
rect 2562 17167 2596 17201
rect 2658 17371 2692 17405
rect 2658 17303 2692 17337
rect 2658 17235 2692 17269
rect 2658 17167 2692 17201
rect 2754 17371 2788 17405
rect 2754 17303 2788 17337
rect 2754 17235 2788 17269
rect 2754 17167 2788 17201
rect 2850 17371 2884 17405
rect 2850 17303 2884 17337
rect 2850 17235 2884 17269
rect 2850 17167 2884 17201
rect 2946 17371 2980 17405
rect 2946 17303 2980 17337
rect 2946 17235 2980 17269
rect 2946 17167 2980 17201
rect 3042 17371 3076 17405
rect 3042 17303 3076 17337
rect 3042 17235 3076 17269
rect 3042 17167 3076 17201
rect 3138 17371 3172 17405
rect 3138 17303 3172 17337
rect 3138 17235 3172 17269
rect 3138 17167 3172 17201
rect 3234 17371 3268 17405
rect 3234 17303 3268 17337
rect 3234 17235 3268 17269
rect 3234 17167 3268 17201
rect 3330 17371 3364 17405
rect 3330 17303 3364 17337
rect 3330 17235 3364 17269
rect 3330 17167 3364 17201
rect 3426 17371 3460 17405
rect 3426 17303 3460 17337
rect 3426 17235 3460 17269
rect 3426 17167 3460 17201
rect 3987 17371 4021 17405
rect 3987 17303 4021 17337
rect 3987 17235 4021 17269
rect 3987 17167 4021 17201
rect 4083 17371 4117 17405
rect 4083 17303 4117 17337
rect 4083 17235 4117 17269
rect 4083 17167 4117 17201
rect 4179 17371 4213 17405
rect 4179 17303 4213 17337
rect 4179 17235 4213 17269
rect 4179 17167 4213 17201
rect 4275 17371 4309 17405
rect 4275 17303 4309 17337
rect 4275 17235 4309 17269
rect 4275 17167 4309 17201
rect 4371 17371 4405 17405
rect 4371 17303 4405 17337
rect 4371 17235 4405 17269
rect 4371 17167 4405 17201
rect 4467 17371 4501 17405
rect 4467 17303 4501 17337
rect 4467 17235 4501 17269
rect 4467 17167 4501 17201
rect 4563 17371 4597 17405
rect 4563 17303 4597 17337
rect 4563 17235 4597 17269
rect 4563 17167 4597 17201
rect 4659 17371 4693 17405
rect 4659 17303 4693 17337
rect 4659 17235 4693 17269
rect 4659 17167 4693 17201
rect 4755 17371 4789 17405
rect 4755 17303 4789 17337
rect 4755 17235 4789 17269
rect 4755 17167 4789 17201
rect 4851 17371 4885 17405
rect 4851 17303 4885 17337
rect 4851 17235 4885 17269
rect 4851 17167 4885 17201
rect 4947 17371 4981 17405
rect 4947 17303 4981 17337
rect 4947 17235 4981 17269
rect 4947 17167 4981 17201
rect 5356 17163 5390 17197
rect 5356 17095 5390 17129
rect 5356 17027 5390 17061
rect 5440 17163 5474 17197
rect 5440 17095 5474 17129
rect 5440 17027 5474 17061
rect 313 16080 347 16114
rect 313 16012 347 16046
rect 313 15944 347 15978
rect 313 15876 347 15910
rect 409 16080 443 16114
rect 409 16012 443 16046
rect 409 15944 443 15978
rect 409 15876 443 15910
rect 505 16080 539 16114
rect 505 16012 539 16046
rect 505 15944 539 15978
rect 505 15876 539 15910
rect 601 16080 635 16114
rect 601 16012 635 16046
rect 601 15944 635 15978
rect 601 15876 635 15910
rect 697 16080 731 16114
rect 697 16012 731 16046
rect 697 15944 731 15978
rect 697 15876 731 15910
rect 793 16080 827 16114
rect 793 16012 827 16046
rect 793 15944 827 15978
rect 793 15876 827 15910
rect 889 16080 923 16114
rect 889 16012 923 16046
rect 889 15944 923 15978
rect 889 15876 923 15910
rect 985 16080 1019 16114
rect 985 16012 1019 16046
rect 985 15944 1019 15978
rect 985 15876 1019 15910
rect 1081 16080 1115 16114
rect 1081 16012 1115 16046
rect 1081 15944 1115 15978
rect 1081 15876 1115 15910
rect 1177 16080 1211 16114
rect 1177 16012 1211 16046
rect 1177 15944 1211 15978
rect 1177 15876 1211 15910
rect 1273 16080 1307 16114
rect 1273 16012 1307 16046
rect 1273 15944 1307 15978
rect 1273 15876 1307 15910
rect 2466 16084 2500 16118
rect 2466 16016 2500 16050
rect 2466 15948 2500 15982
rect 2466 15880 2500 15914
rect 2562 16084 2596 16118
rect 2562 16016 2596 16050
rect 2562 15948 2596 15982
rect 2562 15880 2596 15914
rect 2658 16084 2692 16118
rect 2658 16016 2692 16050
rect 2658 15948 2692 15982
rect 2658 15880 2692 15914
rect 2754 16084 2788 16118
rect 2754 16016 2788 16050
rect 2754 15948 2788 15982
rect 2754 15880 2788 15914
rect 2850 16084 2884 16118
rect 2850 16016 2884 16050
rect 2850 15948 2884 15982
rect 2850 15880 2884 15914
rect 2946 16084 2980 16118
rect 2946 16016 2980 16050
rect 2946 15948 2980 15982
rect 2946 15880 2980 15914
rect 3042 16084 3076 16118
rect 3042 16016 3076 16050
rect 3042 15948 3076 15982
rect 3042 15880 3076 15914
rect 3138 16084 3172 16118
rect 3138 16016 3172 16050
rect 3138 15948 3172 15982
rect 3138 15880 3172 15914
rect 3234 16084 3268 16118
rect 3234 16016 3268 16050
rect 3234 15948 3268 15982
rect 3234 15880 3268 15914
rect 3330 16084 3364 16118
rect 3330 16016 3364 16050
rect 3330 15948 3364 15982
rect 3330 15880 3364 15914
rect 3426 16084 3460 16118
rect 3426 16016 3460 16050
rect 3426 15948 3460 15982
rect 3426 15880 3460 15914
rect 3987 16084 4021 16118
rect 3987 16016 4021 16050
rect 3987 15948 4021 15982
rect 3987 15880 4021 15914
rect 4083 16084 4117 16118
rect 4083 16016 4117 16050
rect 4083 15948 4117 15982
rect 4083 15880 4117 15914
rect 4179 16084 4213 16118
rect 4179 16016 4213 16050
rect 4179 15948 4213 15982
rect 4179 15880 4213 15914
rect 4275 16084 4309 16118
rect 4275 16016 4309 16050
rect 4275 15948 4309 15982
rect 4275 15880 4309 15914
rect 4371 16084 4405 16118
rect 4371 16016 4405 16050
rect 4371 15948 4405 15982
rect 4371 15880 4405 15914
rect 4467 16084 4501 16118
rect 4467 16016 4501 16050
rect 4467 15948 4501 15982
rect 4467 15880 4501 15914
rect 4563 16084 4597 16118
rect 4563 16016 4597 16050
rect 4563 15948 4597 15982
rect 4563 15880 4597 15914
rect 4659 16084 4693 16118
rect 4659 16016 4693 16050
rect 4659 15948 4693 15982
rect 4659 15880 4693 15914
rect 4755 16084 4789 16118
rect 4755 16016 4789 16050
rect 4755 15948 4789 15982
rect 4755 15880 4789 15914
rect 4851 16084 4885 16118
rect 4851 16016 4885 16050
rect 4851 15948 4885 15982
rect 4851 15880 4885 15914
rect 4947 16084 4981 16118
rect 4947 16016 4981 16050
rect 4947 15948 4981 15982
rect 4947 15880 4981 15914
rect 5356 15876 5390 15910
rect 5356 15808 5390 15842
rect 5356 15740 5390 15774
rect 5440 15876 5474 15910
rect 5440 15808 5474 15842
rect 5440 15740 5474 15774
rect 313 14793 347 14827
rect 313 14725 347 14759
rect 313 14657 347 14691
rect 313 14589 347 14623
rect 409 14793 443 14827
rect 409 14725 443 14759
rect 409 14657 443 14691
rect 409 14589 443 14623
rect 505 14793 539 14827
rect 505 14725 539 14759
rect 505 14657 539 14691
rect 505 14589 539 14623
rect 601 14793 635 14827
rect 601 14725 635 14759
rect 601 14657 635 14691
rect 601 14589 635 14623
rect 697 14793 731 14827
rect 697 14725 731 14759
rect 697 14657 731 14691
rect 697 14589 731 14623
rect 793 14793 827 14827
rect 793 14725 827 14759
rect 793 14657 827 14691
rect 793 14589 827 14623
rect 889 14793 923 14827
rect 889 14725 923 14759
rect 889 14657 923 14691
rect 889 14589 923 14623
rect 985 14793 1019 14827
rect 985 14725 1019 14759
rect 985 14657 1019 14691
rect 985 14589 1019 14623
rect 1081 14793 1115 14827
rect 1081 14725 1115 14759
rect 1081 14657 1115 14691
rect 1081 14589 1115 14623
rect 1177 14793 1211 14827
rect 1177 14725 1211 14759
rect 1177 14657 1211 14691
rect 1177 14589 1211 14623
rect 1273 14793 1307 14827
rect 1273 14725 1307 14759
rect 1273 14657 1307 14691
rect 1273 14589 1307 14623
rect 2466 14797 2500 14831
rect 2466 14729 2500 14763
rect 2466 14661 2500 14695
rect 2466 14593 2500 14627
rect 2562 14797 2596 14831
rect 2562 14729 2596 14763
rect 2562 14661 2596 14695
rect 2562 14593 2596 14627
rect 2658 14797 2692 14831
rect 2658 14729 2692 14763
rect 2658 14661 2692 14695
rect 2658 14593 2692 14627
rect 2754 14797 2788 14831
rect 2754 14729 2788 14763
rect 2754 14661 2788 14695
rect 2754 14593 2788 14627
rect 2850 14797 2884 14831
rect 2850 14729 2884 14763
rect 2850 14661 2884 14695
rect 2850 14593 2884 14627
rect 2946 14797 2980 14831
rect 2946 14729 2980 14763
rect 2946 14661 2980 14695
rect 2946 14593 2980 14627
rect 3042 14797 3076 14831
rect 3042 14729 3076 14763
rect 3042 14661 3076 14695
rect 3042 14593 3076 14627
rect 3138 14797 3172 14831
rect 3138 14729 3172 14763
rect 3138 14661 3172 14695
rect 3138 14593 3172 14627
rect 3234 14797 3268 14831
rect 3234 14729 3268 14763
rect 3234 14661 3268 14695
rect 3234 14593 3268 14627
rect 3330 14797 3364 14831
rect 3330 14729 3364 14763
rect 3330 14661 3364 14695
rect 3330 14593 3364 14627
rect 3426 14797 3460 14831
rect 3426 14729 3460 14763
rect 3426 14661 3460 14695
rect 3426 14593 3460 14627
rect 3987 14797 4021 14831
rect 3987 14729 4021 14763
rect 3987 14661 4021 14695
rect 3987 14593 4021 14627
rect 4083 14797 4117 14831
rect 4083 14729 4117 14763
rect 4083 14661 4117 14695
rect 4083 14593 4117 14627
rect 4179 14797 4213 14831
rect 4179 14729 4213 14763
rect 4179 14661 4213 14695
rect 4179 14593 4213 14627
rect 4275 14797 4309 14831
rect 4275 14729 4309 14763
rect 4275 14661 4309 14695
rect 4275 14593 4309 14627
rect 4371 14797 4405 14831
rect 4371 14729 4405 14763
rect 4371 14661 4405 14695
rect 4371 14593 4405 14627
rect 4467 14797 4501 14831
rect 4467 14729 4501 14763
rect 4467 14661 4501 14695
rect 4467 14593 4501 14627
rect 4563 14797 4597 14831
rect 4563 14729 4597 14763
rect 4563 14661 4597 14695
rect 4563 14593 4597 14627
rect 4659 14797 4693 14831
rect 4659 14729 4693 14763
rect 4659 14661 4693 14695
rect 4659 14593 4693 14627
rect 4755 14797 4789 14831
rect 4755 14729 4789 14763
rect 4755 14661 4789 14695
rect 4755 14593 4789 14627
rect 4851 14797 4885 14831
rect 4851 14729 4885 14763
rect 4851 14661 4885 14695
rect 4851 14593 4885 14627
rect 4947 14797 4981 14831
rect 4947 14729 4981 14763
rect 4947 14661 4981 14695
rect 4947 14593 4981 14627
rect 5356 14589 5390 14623
rect 5356 14521 5390 14555
rect 5356 14453 5390 14487
rect 5440 14589 5474 14623
rect 5440 14521 5474 14555
rect 5440 14453 5474 14487
rect 313 13506 347 13540
rect 313 13438 347 13472
rect 313 13370 347 13404
rect 313 13302 347 13336
rect 409 13506 443 13540
rect 409 13438 443 13472
rect 409 13370 443 13404
rect 409 13302 443 13336
rect 505 13506 539 13540
rect 505 13438 539 13472
rect 505 13370 539 13404
rect 505 13302 539 13336
rect 601 13506 635 13540
rect 601 13438 635 13472
rect 601 13370 635 13404
rect 601 13302 635 13336
rect 697 13506 731 13540
rect 697 13438 731 13472
rect 697 13370 731 13404
rect 697 13302 731 13336
rect 793 13506 827 13540
rect 793 13438 827 13472
rect 793 13370 827 13404
rect 793 13302 827 13336
rect 889 13506 923 13540
rect 889 13438 923 13472
rect 889 13370 923 13404
rect 889 13302 923 13336
rect 985 13506 1019 13540
rect 985 13438 1019 13472
rect 985 13370 1019 13404
rect 985 13302 1019 13336
rect 1081 13506 1115 13540
rect 1081 13438 1115 13472
rect 1081 13370 1115 13404
rect 1081 13302 1115 13336
rect 1177 13506 1211 13540
rect 1177 13438 1211 13472
rect 1177 13370 1211 13404
rect 1177 13302 1211 13336
rect 1273 13506 1307 13540
rect 1273 13438 1307 13472
rect 1273 13370 1307 13404
rect 1273 13302 1307 13336
rect 2466 13510 2500 13544
rect 2466 13442 2500 13476
rect 2466 13374 2500 13408
rect 2466 13306 2500 13340
rect 2562 13510 2596 13544
rect 2562 13442 2596 13476
rect 2562 13374 2596 13408
rect 2562 13306 2596 13340
rect 2658 13510 2692 13544
rect 2658 13442 2692 13476
rect 2658 13374 2692 13408
rect 2658 13306 2692 13340
rect 2754 13510 2788 13544
rect 2754 13442 2788 13476
rect 2754 13374 2788 13408
rect 2754 13306 2788 13340
rect 2850 13510 2884 13544
rect 2850 13442 2884 13476
rect 2850 13374 2884 13408
rect 2850 13306 2884 13340
rect 2946 13510 2980 13544
rect 2946 13442 2980 13476
rect 2946 13374 2980 13408
rect 2946 13306 2980 13340
rect 3042 13510 3076 13544
rect 3042 13442 3076 13476
rect 3042 13374 3076 13408
rect 3042 13306 3076 13340
rect 3138 13510 3172 13544
rect 3138 13442 3172 13476
rect 3138 13374 3172 13408
rect 3138 13306 3172 13340
rect 3234 13510 3268 13544
rect 3234 13442 3268 13476
rect 3234 13374 3268 13408
rect 3234 13306 3268 13340
rect 3330 13510 3364 13544
rect 3330 13442 3364 13476
rect 3330 13374 3364 13408
rect 3330 13306 3364 13340
rect 3426 13510 3460 13544
rect 3426 13442 3460 13476
rect 3426 13374 3460 13408
rect 3426 13306 3460 13340
rect 3987 13510 4021 13544
rect 3987 13442 4021 13476
rect 3987 13374 4021 13408
rect 3987 13306 4021 13340
rect 4083 13510 4117 13544
rect 4083 13442 4117 13476
rect 4083 13374 4117 13408
rect 4083 13306 4117 13340
rect 4179 13510 4213 13544
rect 4179 13442 4213 13476
rect 4179 13374 4213 13408
rect 4179 13306 4213 13340
rect 4275 13510 4309 13544
rect 4275 13442 4309 13476
rect 4275 13374 4309 13408
rect 4275 13306 4309 13340
rect 4371 13510 4405 13544
rect 4371 13442 4405 13476
rect 4371 13374 4405 13408
rect 4371 13306 4405 13340
rect 4467 13510 4501 13544
rect 4467 13442 4501 13476
rect 4467 13374 4501 13408
rect 4467 13306 4501 13340
rect 4563 13510 4597 13544
rect 4563 13442 4597 13476
rect 4563 13374 4597 13408
rect 4563 13306 4597 13340
rect 4659 13510 4693 13544
rect 4659 13442 4693 13476
rect 4659 13374 4693 13408
rect 4659 13306 4693 13340
rect 4755 13510 4789 13544
rect 4755 13442 4789 13476
rect 4755 13374 4789 13408
rect 4755 13306 4789 13340
rect 4851 13510 4885 13544
rect 4851 13442 4885 13476
rect 4851 13374 4885 13408
rect 4851 13306 4885 13340
rect 4947 13510 4981 13544
rect 4947 13442 4981 13476
rect 4947 13374 4981 13408
rect 4947 13306 4981 13340
rect 5356 13302 5390 13336
rect 5356 13234 5390 13268
rect 5356 13166 5390 13200
rect 5440 13302 5474 13336
rect 5440 13234 5474 13268
rect 5440 13166 5474 13200
rect 313 12219 347 12253
rect 313 12151 347 12185
rect 313 12083 347 12117
rect 313 12015 347 12049
rect 409 12219 443 12253
rect 409 12151 443 12185
rect 409 12083 443 12117
rect 409 12015 443 12049
rect 505 12219 539 12253
rect 505 12151 539 12185
rect 505 12083 539 12117
rect 505 12015 539 12049
rect 601 12219 635 12253
rect 601 12151 635 12185
rect 601 12083 635 12117
rect 601 12015 635 12049
rect 697 12219 731 12253
rect 697 12151 731 12185
rect 697 12083 731 12117
rect 697 12015 731 12049
rect 793 12219 827 12253
rect 793 12151 827 12185
rect 793 12083 827 12117
rect 793 12015 827 12049
rect 889 12219 923 12253
rect 889 12151 923 12185
rect 889 12083 923 12117
rect 889 12015 923 12049
rect 985 12219 1019 12253
rect 985 12151 1019 12185
rect 985 12083 1019 12117
rect 985 12015 1019 12049
rect 1081 12219 1115 12253
rect 1081 12151 1115 12185
rect 1081 12083 1115 12117
rect 1081 12015 1115 12049
rect 1177 12219 1211 12253
rect 1177 12151 1211 12185
rect 1177 12083 1211 12117
rect 1177 12015 1211 12049
rect 1273 12219 1307 12253
rect 1273 12151 1307 12185
rect 1273 12083 1307 12117
rect 1273 12015 1307 12049
rect 2466 12223 2500 12257
rect 2466 12155 2500 12189
rect 2466 12087 2500 12121
rect 2466 12019 2500 12053
rect 2562 12223 2596 12257
rect 2562 12155 2596 12189
rect 2562 12087 2596 12121
rect 2562 12019 2596 12053
rect 2658 12223 2692 12257
rect 2658 12155 2692 12189
rect 2658 12087 2692 12121
rect 2658 12019 2692 12053
rect 2754 12223 2788 12257
rect 2754 12155 2788 12189
rect 2754 12087 2788 12121
rect 2754 12019 2788 12053
rect 2850 12223 2884 12257
rect 2850 12155 2884 12189
rect 2850 12087 2884 12121
rect 2850 12019 2884 12053
rect 2946 12223 2980 12257
rect 2946 12155 2980 12189
rect 2946 12087 2980 12121
rect 2946 12019 2980 12053
rect 3042 12223 3076 12257
rect 3042 12155 3076 12189
rect 3042 12087 3076 12121
rect 3042 12019 3076 12053
rect 3138 12223 3172 12257
rect 3138 12155 3172 12189
rect 3138 12087 3172 12121
rect 3138 12019 3172 12053
rect 3234 12223 3268 12257
rect 3234 12155 3268 12189
rect 3234 12087 3268 12121
rect 3234 12019 3268 12053
rect 3330 12223 3364 12257
rect 3330 12155 3364 12189
rect 3330 12087 3364 12121
rect 3330 12019 3364 12053
rect 3426 12223 3460 12257
rect 3426 12155 3460 12189
rect 3426 12087 3460 12121
rect 3426 12019 3460 12053
rect 3987 12223 4021 12257
rect 3987 12155 4021 12189
rect 3987 12087 4021 12121
rect 3987 12019 4021 12053
rect 4083 12223 4117 12257
rect 4083 12155 4117 12189
rect 4083 12087 4117 12121
rect 4083 12019 4117 12053
rect 4179 12223 4213 12257
rect 4179 12155 4213 12189
rect 4179 12087 4213 12121
rect 4179 12019 4213 12053
rect 4275 12223 4309 12257
rect 4275 12155 4309 12189
rect 4275 12087 4309 12121
rect 4275 12019 4309 12053
rect 4371 12223 4405 12257
rect 4371 12155 4405 12189
rect 4371 12087 4405 12121
rect 4371 12019 4405 12053
rect 4467 12223 4501 12257
rect 4467 12155 4501 12189
rect 4467 12087 4501 12121
rect 4467 12019 4501 12053
rect 4563 12223 4597 12257
rect 4563 12155 4597 12189
rect 4563 12087 4597 12121
rect 4563 12019 4597 12053
rect 4659 12223 4693 12257
rect 4659 12155 4693 12189
rect 4659 12087 4693 12121
rect 4659 12019 4693 12053
rect 4755 12223 4789 12257
rect 4755 12155 4789 12189
rect 4755 12087 4789 12121
rect 4755 12019 4789 12053
rect 4851 12223 4885 12257
rect 4851 12155 4885 12189
rect 4851 12087 4885 12121
rect 4851 12019 4885 12053
rect 4947 12223 4981 12257
rect 4947 12155 4981 12189
rect 4947 12087 4981 12121
rect 4947 12019 4981 12053
rect 5356 12015 5390 12049
rect 5356 11947 5390 11981
rect 5356 11879 5390 11913
rect 5440 12015 5474 12049
rect 5440 11947 5474 11981
rect 5440 11879 5474 11913
rect 313 10932 347 10966
rect 313 10864 347 10898
rect 313 10796 347 10830
rect 313 10728 347 10762
rect 409 10932 443 10966
rect 409 10864 443 10898
rect 409 10796 443 10830
rect 409 10728 443 10762
rect 505 10932 539 10966
rect 505 10864 539 10898
rect 505 10796 539 10830
rect 505 10728 539 10762
rect 601 10932 635 10966
rect 601 10864 635 10898
rect 601 10796 635 10830
rect 601 10728 635 10762
rect 697 10932 731 10966
rect 697 10864 731 10898
rect 697 10796 731 10830
rect 697 10728 731 10762
rect 793 10932 827 10966
rect 793 10864 827 10898
rect 793 10796 827 10830
rect 793 10728 827 10762
rect 889 10932 923 10966
rect 889 10864 923 10898
rect 889 10796 923 10830
rect 889 10728 923 10762
rect 985 10932 1019 10966
rect 985 10864 1019 10898
rect 985 10796 1019 10830
rect 985 10728 1019 10762
rect 1081 10932 1115 10966
rect 1081 10864 1115 10898
rect 1081 10796 1115 10830
rect 1081 10728 1115 10762
rect 1177 10932 1211 10966
rect 1177 10864 1211 10898
rect 1177 10796 1211 10830
rect 1177 10728 1211 10762
rect 1273 10932 1307 10966
rect 1273 10864 1307 10898
rect 1273 10796 1307 10830
rect 1273 10728 1307 10762
rect 2466 10936 2500 10970
rect 2466 10868 2500 10902
rect 2466 10800 2500 10834
rect 2466 10732 2500 10766
rect 2562 10936 2596 10970
rect 2562 10868 2596 10902
rect 2562 10800 2596 10834
rect 2562 10732 2596 10766
rect 2658 10936 2692 10970
rect 2658 10868 2692 10902
rect 2658 10800 2692 10834
rect 2658 10732 2692 10766
rect 2754 10936 2788 10970
rect 2754 10868 2788 10902
rect 2754 10800 2788 10834
rect 2754 10732 2788 10766
rect 2850 10936 2884 10970
rect 2850 10868 2884 10902
rect 2850 10800 2884 10834
rect 2850 10732 2884 10766
rect 2946 10936 2980 10970
rect 2946 10868 2980 10902
rect 2946 10800 2980 10834
rect 2946 10732 2980 10766
rect 3042 10936 3076 10970
rect 3042 10868 3076 10902
rect 3042 10800 3076 10834
rect 3042 10732 3076 10766
rect 3138 10936 3172 10970
rect 3138 10868 3172 10902
rect 3138 10800 3172 10834
rect 3138 10732 3172 10766
rect 3234 10936 3268 10970
rect 3234 10868 3268 10902
rect 3234 10800 3268 10834
rect 3234 10732 3268 10766
rect 3330 10936 3364 10970
rect 3330 10868 3364 10902
rect 3330 10800 3364 10834
rect 3330 10732 3364 10766
rect 3426 10936 3460 10970
rect 3426 10868 3460 10902
rect 3426 10800 3460 10834
rect 3426 10732 3460 10766
rect 3987 10936 4021 10970
rect 3987 10868 4021 10902
rect 3987 10800 4021 10834
rect 3987 10732 4021 10766
rect 4083 10936 4117 10970
rect 4083 10868 4117 10902
rect 4083 10800 4117 10834
rect 4083 10732 4117 10766
rect 4179 10936 4213 10970
rect 4179 10868 4213 10902
rect 4179 10800 4213 10834
rect 4179 10732 4213 10766
rect 4275 10936 4309 10970
rect 4275 10868 4309 10902
rect 4275 10800 4309 10834
rect 4275 10732 4309 10766
rect 4371 10936 4405 10970
rect 4371 10868 4405 10902
rect 4371 10800 4405 10834
rect 4371 10732 4405 10766
rect 4467 10936 4501 10970
rect 4467 10868 4501 10902
rect 4467 10800 4501 10834
rect 4467 10732 4501 10766
rect 4563 10936 4597 10970
rect 4563 10868 4597 10902
rect 4563 10800 4597 10834
rect 4563 10732 4597 10766
rect 4659 10936 4693 10970
rect 4659 10868 4693 10902
rect 4659 10800 4693 10834
rect 4659 10732 4693 10766
rect 4755 10936 4789 10970
rect 4755 10868 4789 10902
rect 4755 10800 4789 10834
rect 4755 10732 4789 10766
rect 4851 10936 4885 10970
rect 4851 10868 4885 10902
rect 4851 10800 4885 10834
rect 4851 10732 4885 10766
rect 4947 10936 4981 10970
rect 4947 10868 4981 10902
rect 4947 10800 4981 10834
rect 4947 10732 4981 10766
rect 5356 10728 5390 10762
rect 5356 10660 5390 10694
rect 5356 10592 5390 10626
rect 5440 10728 5474 10762
rect 5440 10660 5474 10694
rect 5440 10592 5474 10626
rect 313 9645 347 9679
rect 313 9577 347 9611
rect 313 9509 347 9543
rect 313 9441 347 9475
rect 409 9645 443 9679
rect 409 9577 443 9611
rect 409 9509 443 9543
rect 409 9441 443 9475
rect 505 9645 539 9679
rect 505 9577 539 9611
rect 505 9509 539 9543
rect 505 9441 539 9475
rect 601 9645 635 9679
rect 601 9577 635 9611
rect 601 9509 635 9543
rect 601 9441 635 9475
rect 697 9645 731 9679
rect 697 9577 731 9611
rect 697 9509 731 9543
rect 697 9441 731 9475
rect 793 9645 827 9679
rect 793 9577 827 9611
rect 793 9509 827 9543
rect 793 9441 827 9475
rect 889 9645 923 9679
rect 889 9577 923 9611
rect 889 9509 923 9543
rect 889 9441 923 9475
rect 985 9645 1019 9679
rect 985 9577 1019 9611
rect 985 9509 1019 9543
rect 985 9441 1019 9475
rect 1081 9645 1115 9679
rect 1081 9577 1115 9611
rect 1081 9509 1115 9543
rect 1081 9441 1115 9475
rect 1177 9645 1211 9679
rect 1177 9577 1211 9611
rect 1177 9509 1211 9543
rect 1177 9441 1211 9475
rect 1273 9645 1307 9679
rect 1273 9577 1307 9611
rect 1273 9509 1307 9543
rect 1273 9441 1307 9475
rect 2466 9649 2500 9683
rect 2466 9581 2500 9615
rect 2466 9513 2500 9547
rect 2466 9445 2500 9479
rect 2562 9649 2596 9683
rect 2562 9581 2596 9615
rect 2562 9513 2596 9547
rect 2562 9445 2596 9479
rect 2658 9649 2692 9683
rect 2658 9581 2692 9615
rect 2658 9513 2692 9547
rect 2658 9445 2692 9479
rect 2754 9649 2788 9683
rect 2754 9581 2788 9615
rect 2754 9513 2788 9547
rect 2754 9445 2788 9479
rect 2850 9649 2884 9683
rect 2850 9581 2884 9615
rect 2850 9513 2884 9547
rect 2850 9445 2884 9479
rect 2946 9649 2980 9683
rect 2946 9581 2980 9615
rect 2946 9513 2980 9547
rect 2946 9445 2980 9479
rect 3042 9649 3076 9683
rect 3042 9581 3076 9615
rect 3042 9513 3076 9547
rect 3042 9445 3076 9479
rect 3138 9649 3172 9683
rect 3138 9581 3172 9615
rect 3138 9513 3172 9547
rect 3138 9445 3172 9479
rect 3234 9649 3268 9683
rect 3234 9581 3268 9615
rect 3234 9513 3268 9547
rect 3234 9445 3268 9479
rect 3330 9649 3364 9683
rect 3330 9581 3364 9615
rect 3330 9513 3364 9547
rect 3330 9445 3364 9479
rect 3426 9649 3460 9683
rect 3426 9581 3460 9615
rect 3426 9513 3460 9547
rect 3426 9445 3460 9479
rect 3987 9649 4021 9683
rect 3987 9581 4021 9615
rect 3987 9513 4021 9547
rect 3987 9445 4021 9479
rect 4083 9649 4117 9683
rect 4083 9581 4117 9615
rect 4083 9513 4117 9547
rect 4083 9445 4117 9479
rect 4179 9649 4213 9683
rect 4179 9581 4213 9615
rect 4179 9513 4213 9547
rect 4179 9445 4213 9479
rect 4275 9649 4309 9683
rect 4275 9581 4309 9615
rect 4275 9513 4309 9547
rect 4275 9445 4309 9479
rect 4371 9649 4405 9683
rect 4371 9581 4405 9615
rect 4371 9513 4405 9547
rect 4371 9445 4405 9479
rect 4467 9649 4501 9683
rect 4467 9581 4501 9615
rect 4467 9513 4501 9547
rect 4467 9445 4501 9479
rect 4563 9649 4597 9683
rect 4563 9581 4597 9615
rect 4563 9513 4597 9547
rect 4563 9445 4597 9479
rect 4659 9649 4693 9683
rect 4659 9581 4693 9615
rect 4659 9513 4693 9547
rect 4659 9445 4693 9479
rect 4755 9649 4789 9683
rect 4755 9581 4789 9615
rect 4755 9513 4789 9547
rect 4755 9445 4789 9479
rect 4851 9649 4885 9683
rect 4851 9581 4885 9615
rect 4851 9513 4885 9547
rect 4851 9445 4885 9479
rect 4947 9649 4981 9683
rect 4947 9581 4981 9615
rect 4947 9513 4981 9547
rect 4947 9445 4981 9479
rect 5356 9441 5390 9475
rect 5356 9373 5390 9407
rect 5356 9305 5390 9339
rect 5440 9441 5474 9475
rect 5440 9373 5474 9407
rect 5440 9305 5474 9339
rect 313 8358 347 8392
rect 313 8290 347 8324
rect 313 8222 347 8256
rect 313 8154 347 8188
rect 409 8358 443 8392
rect 409 8290 443 8324
rect 409 8222 443 8256
rect 409 8154 443 8188
rect 505 8358 539 8392
rect 505 8290 539 8324
rect 505 8222 539 8256
rect 505 8154 539 8188
rect 601 8358 635 8392
rect 601 8290 635 8324
rect 601 8222 635 8256
rect 601 8154 635 8188
rect 697 8358 731 8392
rect 697 8290 731 8324
rect 697 8222 731 8256
rect 697 8154 731 8188
rect 793 8358 827 8392
rect 793 8290 827 8324
rect 793 8222 827 8256
rect 793 8154 827 8188
rect 889 8358 923 8392
rect 889 8290 923 8324
rect 889 8222 923 8256
rect 889 8154 923 8188
rect 985 8358 1019 8392
rect 985 8290 1019 8324
rect 985 8222 1019 8256
rect 985 8154 1019 8188
rect 1081 8358 1115 8392
rect 1081 8290 1115 8324
rect 1081 8222 1115 8256
rect 1081 8154 1115 8188
rect 1177 8358 1211 8392
rect 1177 8290 1211 8324
rect 1177 8222 1211 8256
rect 1177 8154 1211 8188
rect 1273 8358 1307 8392
rect 1273 8290 1307 8324
rect 1273 8222 1307 8256
rect 1273 8154 1307 8188
rect 2466 8362 2500 8396
rect 2466 8294 2500 8328
rect 2466 8226 2500 8260
rect 2466 8158 2500 8192
rect 2562 8362 2596 8396
rect 2562 8294 2596 8328
rect 2562 8226 2596 8260
rect 2562 8158 2596 8192
rect 2658 8362 2692 8396
rect 2658 8294 2692 8328
rect 2658 8226 2692 8260
rect 2658 8158 2692 8192
rect 2754 8362 2788 8396
rect 2754 8294 2788 8328
rect 2754 8226 2788 8260
rect 2754 8158 2788 8192
rect 2850 8362 2884 8396
rect 2850 8294 2884 8328
rect 2850 8226 2884 8260
rect 2850 8158 2884 8192
rect 2946 8362 2980 8396
rect 2946 8294 2980 8328
rect 2946 8226 2980 8260
rect 2946 8158 2980 8192
rect 3042 8362 3076 8396
rect 3042 8294 3076 8328
rect 3042 8226 3076 8260
rect 3042 8158 3076 8192
rect 3138 8362 3172 8396
rect 3138 8294 3172 8328
rect 3138 8226 3172 8260
rect 3138 8158 3172 8192
rect 3234 8362 3268 8396
rect 3234 8294 3268 8328
rect 3234 8226 3268 8260
rect 3234 8158 3268 8192
rect 3330 8362 3364 8396
rect 3330 8294 3364 8328
rect 3330 8226 3364 8260
rect 3330 8158 3364 8192
rect 3426 8362 3460 8396
rect 3426 8294 3460 8328
rect 3426 8226 3460 8260
rect 3426 8158 3460 8192
rect 3987 8362 4021 8396
rect 3987 8294 4021 8328
rect 3987 8226 4021 8260
rect 3987 8158 4021 8192
rect 4083 8362 4117 8396
rect 4083 8294 4117 8328
rect 4083 8226 4117 8260
rect 4083 8158 4117 8192
rect 4179 8362 4213 8396
rect 4179 8294 4213 8328
rect 4179 8226 4213 8260
rect 4179 8158 4213 8192
rect 4275 8362 4309 8396
rect 4275 8294 4309 8328
rect 4275 8226 4309 8260
rect 4275 8158 4309 8192
rect 4371 8362 4405 8396
rect 4371 8294 4405 8328
rect 4371 8226 4405 8260
rect 4371 8158 4405 8192
rect 4467 8362 4501 8396
rect 4467 8294 4501 8328
rect 4467 8226 4501 8260
rect 4467 8158 4501 8192
rect 4563 8362 4597 8396
rect 4563 8294 4597 8328
rect 4563 8226 4597 8260
rect 4563 8158 4597 8192
rect 4659 8362 4693 8396
rect 4659 8294 4693 8328
rect 4659 8226 4693 8260
rect 4659 8158 4693 8192
rect 4755 8362 4789 8396
rect 4755 8294 4789 8328
rect 4755 8226 4789 8260
rect 4755 8158 4789 8192
rect 4851 8362 4885 8396
rect 4851 8294 4885 8328
rect 4851 8226 4885 8260
rect 4851 8158 4885 8192
rect 4947 8362 4981 8396
rect 4947 8294 4981 8328
rect 4947 8226 4981 8260
rect 4947 8158 4981 8192
rect 5356 8154 5390 8188
rect 5356 8086 5390 8120
rect 5356 8018 5390 8052
rect 5440 8154 5474 8188
rect 5440 8086 5474 8120
rect 5440 8018 5474 8052
rect 313 7071 347 7105
rect 313 7003 347 7037
rect 313 6935 347 6969
rect 313 6867 347 6901
rect 409 7071 443 7105
rect 409 7003 443 7037
rect 409 6935 443 6969
rect 409 6867 443 6901
rect 505 7071 539 7105
rect 505 7003 539 7037
rect 505 6935 539 6969
rect 505 6867 539 6901
rect 601 7071 635 7105
rect 601 7003 635 7037
rect 601 6935 635 6969
rect 601 6867 635 6901
rect 697 7071 731 7105
rect 697 7003 731 7037
rect 697 6935 731 6969
rect 697 6867 731 6901
rect 793 7071 827 7105
rect 793 7003 827 7037
rect 793 6935 827 6969
rect 793 6867 827 6901
rect 889 7071 923 7105
rect 889 7003 923 7037
rect 889 6935 923 6969
rect 889 6867 923 6901
rect 985 7071 1019 7105
rect 985 7003 1019 7037
rect 985 6935 1019 6969
rect 985 6867 1019 6901
rect 1081 7071 1115 7105
rect 1081 7003 1115 7037
rect 1081 6935 1115 6969
rect 1081 6867 1115 6901
rect 1177 7071 1211 7105
rect 1177 7003 1211 7037
rect 1177 6935 1211 6969
rect 1177 6867 1211 6901
rect 1273 7071 1307 7105
rect 1273 7003 1307 7037
rect 1273 6935 1307 6969
rect 1273 6867 1307 6901
rect 2466 7075 2500 7109
rect 2466 7007 2500 7041
rect 2466 6939 2500 6973
rect 2466 6871 2500 6905
rect 2562 7075 2596 7109
rect 2562 7007 2596 7041
rect 2562 6939 2596 6973
rect 2562 6871 2596 6905
rect 2658 7075 2692 7109
rect 2658 7007 2692 7041
rect 2658 6939 2692 6973
rect 2658 6871 2692 6905
rect 2754 7075 2788 7109
rect 2754 7007 2788 7041
rect 2754 6939 2788 6973
rect 2754 6871 2788 6905
rect 2850 7075 2884 7109
rect 2850 7007 2884 7041
rect 2850 6939 2884 6973
rect 2850 6871 2884 6905
rect 2946 7075 2980 7109
rect 2946 7007 2980 7041
rect 2946 6939 2980 6973
rect 2946 6871 2980 6905
rect 3042 7075 3076 7109
rect 3042 7007 3076 7041
rect 3042 6939 3076 6973
rect 3042 6871 3076 6905
rect 3138 7075 3172 7109
rect 3138 7007 3172 7041
rect 3138 6939 3172 6973
rect 3138 6871 3172 6905
rect 3234 7075 3268 7109
rect 3234 7007 3268 7041
rect 3234 6939 3268 6973
rect 3234 6871 3268 6905
rect 3330 7075 3364 7109
rect 3330 7007 3364 7041
rect 3330 6939 3364 6973
rect 3330 6871 3364 6905
rect 3426 7075 3460 7109
rect 3426 7007 3460 7041
rect 3426 6939 3460 6973
rect 3426 6871 3460 6905
rect 3987 7075 4021 7109
rect 3987 7007 4021 7041
rect 3987 6939 4021 6973
rect 3987 6871 4021 6905
rect 4083 7075 4117 7109
rect 4083 7007 4117 7041
rect 4083 6939 4117 6973
rect 4083 6871 4117 6905
rect 4179 7075 4213 7109
rect 4179 7007 4213 7041
rect 4179 6939 4213 6973
rect 4179 6871 4213 6905
rect 4275 7075 4309 7109
rect 4275 7007 4309 7041
rect 4275 6939 4309 6973
rect 4275 6871 4309 6905
rect 4371 7075 4405 7109
rect 4371 7007 4405 7041
rect 4371 6939 4405 6973
rect 4371 6871 4405 6905
rect 4467 7075 4501 7109
rect 4467 7007 4501 7041
rect 4467 6939 4501 6973
rect 4467 6871 4501 6905
rect 4563 7075 4597 7109
rect 4563 7007 4597 7041
rect 4563 6939 4597 6973
rect 4563 6871 4597 6905
rect 4659 7075 4693 7109
rect 4659 7007 4693 7041
rect 4659 6939 4693 6973
rect 4659 6871 4693 6905
rect 4755 7075 4789 7109
rect 4755 7007 4789 7041
rect 4755 6939 4789 6973
rect 4755 6871 4789 6905
rect 4851 7075 4885 7109
rect 4851 7007 4885 7041
rect 4851 6939 4885 6973
rect 4851 6871 4885 6905
rect 4947 7075 4981 7109
rect 4947 7007 4981 7041
rect 4947 6939 4981 6973
rect 4947 6871 4981 6905
rect 5356 6867 5390 6901
rect 5356 6799 5390 6833
rect 5356 6731 5390 6765
rect 5440 6867 5474 6901
rect 5440 6799 5474 6833
rect 5440 6731 5474 6765
rect 313 5784 347 5818
rect 313 5716 347 5750
rect 313 5648 347 5682
rect 313 5580 347 5614
rect 409 5784 443 5818
rect 409 5716 443 5750
rect 409 5648 443 5682
rect 409 5580 443 5614
rect 505 5784 539 5818
rect 505 5716 539 5750
rect 505 5648 539 5682
rect 505 5580 539 5614
rect 601 5784 635 5818
rect 601 5716 635 5750
rect 601 5648 635 5682
rect 601 5580 635 5614
rect 697 5784 731 5818
rect 697 5716 731 5750
rect 697 5648 731 5682
rect 697 5580 731 5614
rect 793 5784 827 5818
rect 793 5716 827 5750
rect 793 5648 827 5682
rect 793 5580 827 5614
rect 889 5784 923 5818
rect 889 5716 923 5750
rect 889 5648 923 5682
rect 889 5580 923 5614
rect 985 5784 1019 5818
rect 985 5716 1019 5750
rect 985 5648 1019 5682
rect 985 5580 1019 5614
rect 1081 5784 1115 5818
rect 1081 5716 1115 5750
rect 1081 5648 1115 5682
rect 1081 5580 1115 5614
rect 1177 5784 1211 5818
rect 1177 5716 1211 5750
rect 1177 5648 1211 5682
rect 1177 5580 1211 5614
rect 1273 5784 1307 5818
rect 1273 5716 1307 5750
rect 1273 5648 1307 5682
rect 1273 5580 1307 5614
rect 2466 5788 2500 5822
rect 2466 5720 2500 5754
rect 2466 5652 2500 5686
rect 2466 5584 2500 5618
rect 2562 5788 2596 5822
rect 2562 5720 2596 5754
rect 2562 5652 2596 5686
rect 2562 5584 2596 5618
rect 2658 5788 2692 5822
rect 2658 5720 2692 5754
rect 2658 5652 2692 5686
rect 2658 5584 2692 5618
rect 2754 5788 2788 5822
rect 2754 5720 2788 5754
rect 2754 5652 2788 5686
rect 2754 5584 2788 5618
rect 2850 5788 2884 5822
rect 2850 5720 2884 5754
rect 2850 5652 2884 5686
rect 2850 5584 2884 5618
rect 2946 5788 2980 5822
rect 2946 5720 2980 5754
rect 2946 5652 2980 5686
rect 2946 5584 2980 5618
rect 3042 5788 3076 5822
rect 3042 5720 3076 5754
rect 3042 5652 3076 5686
rect 3042 5584 3076 5618
rect 3138 5788 3172 5822
rect 3138 5720 3172 5754
rect 3138 5652 3172 5686
rect 3138 5584 3172 5618
rect 3234 5788 3268 5822
rect 3234 5720 3268 5754
rect 3234 5652 3268 5686
rect 3234 5584 3268 5618
rect 3330 5788 3364 5822
rect 3330 5720 3364 5754
rect 3330 5652 3364 5686
rect 3330 5584 3364 5618
rect 3426 5788 3460 5822
rect 3426 5720 3460 5754
rect 3426 5652 3460 5686
rect 3426 5584 3460 5618
rect 3987 5788 4021 5822
rect 3987 5720 4021 5754
rect 3987 5652 4021 5686
rect 3987 5584 4021 5618
rect 4083 5788 4117 5822
rect 4083 5720 4117 5754
rect 4083 5652 4117 5686
rect 4083 5584 4117 5618
rect 4179 5788 4213 5822
rect 4179 5720 4213 5754
rect 4179 5652 4213 5686
rect 4179 5584 4213 5618
rect 4275 5788 4309 5822
rect 4275 5720 4309 5754
rect 4275 5652 4309 5686
rect 4275 5584 4309 5618
rect 4371 5788 4405 5822
rect 4371 5720 4405 5754
rect 4371 5652 4405 5686
rect 4371 5584 4405 5618
rect 4467 5788 4501 5822
rect 4467 5720 4501 5754
rect 4467 5652 4501 5686
rect 4467 5584 4501 5618
rect 4563 5788 4597 5822
rect 4563 5720 4597 5754
rect 4563 5652 4597 5686
rect 4563 5584 4597 5618
rect 4659 5788 4693 5822
rect 4659 5720 4693 5754
rect 4659 5652 4693 5686
rect 4659 5584 4693 5618
rect 4755 5788 4789 5822
rect 4755 5720 4789 5754
rect 4755 5652 4789 5686
rect 4755 5584 4789 5618
rect 4851 5788 4885 5822
rect 4851 5720 4885 5754
rect 4851 5652 4885 5686
rect 4851 5584 4885 5618
rect 4947 5788 4981 5822
rect 4947 5720 4981 5754
rect 4947 5652 4981 5686
rect 4947 5584 4981 5618
rect 5356 5580 5390 5614
rect 5356 5512 5390 5546
rect 5356 5444 5390 5478
rect 5440 5580 5474 5614
rect 5440 5512 5474 5546
rect 5440 5444 5474 5478
rect 313 4497 347 4531
rect 313 4429 347 4463
rect 313 4361 347 4395
rect 313 4293 347 4327
rect 409 4497 443 4531
rect 409 4429 443 4463
rect 409 4361 443 4395
rect 409 4293 443 4327
rect 505 4497 539 4531
rect 505 4429 539 4463
rect 505 4361 539 4395
rect 505 4293 539 4327
rect 601 4497 635 4531
rect 601 4429 635 4463
rect 601 4361 635 4395
rect 601 4293 635 4327
rect 697 4497 731 4531
rect 697 4429 731 4463
rect 697 4361 731 4395
rect 697 4293 731 4327
rect 793 4497 827 4531
rect 793 4429 827 4463
rect 793 4361 827 4395
rect 793 4293 827 4327
rect 889 4497 923 4531
rect 889 4429 923 4463
rect 889 4361 923 4395
rect 889 4293 923 4327
rect 985 4497 1019 4531
rect 985 4429 1019 4463
rect 985 4361 1019 4395
rect 985 4293 1019 4327
rect 1081 4497 1115 4531
rect 1081 4429 1115 4463
rect 1081 4361 1115 4395
rect 1081 4293 1115 4327
rect 1177 4497 1211 4531
rect 1177 4429 1211 4463
rect 1177 4361 1211 4395
rect 1177 4293 1211 4327
rect 1273 4497 1307 4531
rect 1273 4429 1307 4463
rect 1273 4361 1307 4395
rect 1273 4293 1307 4327
rect 2466 4501 2500 4535
rect 2466 4433 2500 4467
rect 2466 4365 2500 4399
rect 2466 4297 2500 4331
rect 2562 4501 2596 4535
rect 2562 4433 2596 4467
rect 2562 4365 2596 4399
rect 2562 4297 2596 4331
rect 2658 4501 2692 4535
rect 2658 4433 2692 4467
rect 2658 4365 2692 4399
rect 2658 4297 2692 4331
rect 2754 4501 2788 4535
rect 2754 4433 2788 4467
rect 2754 4365 2788 4399
rect 2754 4297 2788 4331
rect 2850 4501 2884 4535
rect 2850 4433 2884 4467
rect 2850 4365 2884 4399
rect 2850 4297 2884 4331
rect 2946 4501 2980 4535
rect 2946 4433 2980 4467
rect 2946 4365 2980 4399
rect 2946 4297 2980 4331
rect 3042 4501 3076 4535
rect 3042 4433 3076 4467
rect 3042 4365 3076 4399
rect 3042 4297 3076 4331
rect 3138 4501 3172 4535
rect 3138 4433 3172 4467
rect 3138 4365 3172 4399
rect 3138 4297 3172 4331
rect 3234 4501 3268 4535
rect 3234 4433 3268 4467
rect 3234 4365 3268 4399
rect 3234 4297 3268 4331
rect 3330 4501 3364 4535
rect 3330 4433 3364 4467
rect 3330 4365 3364 4399
rect 3330 4297 3364 4331
rect 3426 4501 3460 4535
rect 3426 4433 3460 4467
rect 3426 4365 3460 4399
rect 3426 4297 3460 4331
rect 3987 4501 4021 4535
rect 3987 4433 4021 4467
rect 3987 4365 4021 4399
rect 3987 4297 4021 4331
rect 4083 4501 4117 4535
rect 4083 4433 4117 4467
rect 4083 4365 4117 4399
rect 4083 4297 4117 4331
rect 4179 4501 4213 4535
rect 4179 4433 4213 4467
rect 4179 4365 4213 4399
rect 4179 4297 4213 4331
rect 4275 4501 4309 4535
rect 4275 4433 4309 4467
rect 4275 4365 4309 4399
rect 4275 4297 4309 4331
rect 4371 4501 4405 4535
rect 4371 4433 4405 4467
rect 4371 4365 4405 4399
rect 4371 4297 4405 4331
rect 4467 4501 4501 4535
rect 4467 4433 4501 4467
rect 4467 4365 4501 4399
rect 4467 4297 4501 4331
rect 4563 4501 4597 4535
rect 4563 4433 4597 4467
rect 4563 4365 4597 4399
rect 4563 4297 4597 4331
rect 4659 4501 4693 4535
rect 4659 4433 4693 4467
rect 4659 4365 4693 4399
rect 4659 4297 4693 4331
rect 4755 4501 4789 4535
rect 4755 4433 4789 4467
rect 4755 4365 4789 4399
rect 4755 4297 4789 4331
rect 4851 4501 4885 4535
rect 4851 4433 4885 4467
rect 4851 4365 4885 4399
rect 4851 4297 4885 4331
rect 4947 4501 4981 4535
rect 4947 4433 4981 4467
rect 4947 4365 4981 4399
rect 4947 4297 4981 4331
rect 5356 4293 5390 4327
rect 5356 4225 5390 4259
rect 5356 4157 5390 4191
rect 5440 4293 5474 4327
rect 5440 4225 5474 4259
rect 5440 4157 5474 4191
rect 313 3210 347 3244
rect 313 3142 347 3176
rect 313 3074 347 3108
rect 313 3006 347 3040
rect 409 3210 443 3244
rect 409 3142 443 3176
rect 409 3074 443 3108
rect 409 3006 443 3040
rect 505 3210 539 3244
rect 505 3142 539 3176
rect 505 3074 539 3108
rect 505 3006 539 3040
rect 601 3210 635 3244
rect 601 3142 635 3176
rect 601 3074 635 3108
rect 601 3006 635 3040
rect 697 3210 731 3244
rect 697 3142 731 3176
rect 697 3074 731 3108
rect 697 3006 731 3040
rect 793 3210 827 3244
rect 793 3142 827 3176
rect 793 3074 827 3108
rect 793 3006 827 3040
rect 889 3210 923 3244
rect 889 3142 923 3176
rect 889 3074 923 3108
rect 889 3006 923 3040
rect 985 3210 1019 3244
rect 985 3142 1019 3176
rect 985 3074 1019 3108
rect 985 3006 1019 3040
rect 1081 3210 1115 3244
rect 1081 3142 1115 3176
rect 1081 3074 1115 3108
rect 1081 3006 1115 3040
rect 1177 3210 1211 3244
rect 1177 3142 1211 3176
rect 1177 3074 1211 3108
rect 1177 3006 1211 3040
rect 1273 3210 1307 3244
rect 1273 3142 1307 3176
rect 1273 3074 1307 3108
rect 1273 3006 1307 3040
rect 2466 3214 2500 3248
rect 2466 3146 2500 3180
rect 2466 3078 2500 3112
rect 2466 3010 2500 3044
rect 2562 3214 2596 3248
rect 2562 3146 2596 3180
rect 2562 3078 2596 3112
rect 2562 3010 2596 3044
rect 2658 3214 2692 3248
rect 2658 3146 2692 3180
rect 2658 3078 2692 3112
rect 2658 3010 2692 3044
rect 2754 3214 2788 3248
rect 2754 3146 2788 3180
rect 2754 3078 2788 3112
rect 2754 3010 2788 3044
rect 2850 3214 2884 3248
rect 2850 3146 2884 3180
rect 2850 3078 2884 3112
rect 2850 3010 2884 3044
rect 2946 3214 2980 3248
rect 2946 3146 2980 3180
rect 2946 3078 2980 3112
rect 2946 3010 2980 3044
rect 3042 3214 3076 3248
rect 3042 3146 3076 3180
rect 3042 3078 3076 3112
rect 3042 3010 3076 3044
rect 3138 3214 3172 3248
rect 3138 3146 3172 3180
rect 3138 3078 3172 3112
rect 3138 3010 3172 3044
rect 3234 3214 3268 3248
rect 3234 3146 3268 3180
rect 3234 3078 3268 3112
rect 3234 3010 3268 3044
rect 3330 3214 3364 3248
rect 3330 3146 3364 3180
rect 3330 3078 3364 3112
rect 3330 3010 3364 3044
rect 3426 3214 3460 3248
rect 3426 3146 3460 3180
rect 3426 3078 3460 3112
rect 3426 3010 3460 3044
rect 3987 3214 4021 3248
rect 3987 3146 4021 3180
rect 3987 3078 4021 3112
rect 3987 3010 4021 3044
rect 4083 3214 4117 3248
rect 4083 3146 4117 3180
rect 4083 3078 4117 3112
rect 4083 3010 4117 3044
rect 4179 3214 4213 3248
rect 4179 3146 4213 3180
rect 4179 3078 4213 3112
rect 4179 3010 4213 3044
rect 4275 3214 4309 3248
rect 4275 3146 4309 3180
rect 4275 3078 4309 3112
rect 4275 3010 4309 3044
rect 4371 3214 4405 3248
rect 4371 3146 4405 3180
rect 4371 3078 4405 3112
rect 4371 3010 4405 3044
rect 4467 3214 4501 3248
rect 4467 3146 4501 3180
rect 4467 3078 4501 3112
rect 4467 3010 4501 3044
rect 4563 3214 4597 3248
rect 4563 3146 4597 3180
rect 4563 3078 4597 3112
rect 4563 3010 4597 3044
rect 4659 3214 4693 3248
rect 4659 3146 4693 3180
rect 4659 3078 4693 3112
rect 4659 3010 4693 3044
rect 4755 3214 4789 3248
rect 4755 3146 4789 3180
rect 4755 3078 4789 3112
rect 4755 3010 4789 3044
rect 4851 3214 4885 3248
rect 4851 3146 4885 3180
rect 4851 3078 4885 3112
rect 4851 3010 4885 3044
rect 4947 3214 4981 3248
rect 4947 3146 4981 3180
rect 4947 3078 4981 3112
rect 4947 3010 4981 3044
rect 5356 3006 5390 3040
rect 5356 2938 5390 2972
rect 5356 2870 5390 2904
rect 5440 3006 5474 3040
rect 5440 2938 5474 2972
rect 5440 2870 5474 2904
rect 313 1923 347 1957
rect 313 1855 347 1889
rect 313 1787 347 1821
rect 313 1719 347 1753
rect 409 1923 443 1957
rect 409 1855 443 1889
rect 409 1787 443 1821
rect 409 1719 443 1753
rect 505 1923 539 1957
rect 505 1855 539 1889
rect 505 1787 539 1821
rect 505 1719 539 1753
rect 601 1923 635 1957
rect 601 1855 635 1889
rect 601 1787 635 1821
rect 601 1719 635 1753
rect 697 1923 731 1957
rect 697 1855 731 1889
rect 697 1787 731 1821
rect 697 1719 731 1753
rect 793 1923 827 1957
rect 793 1855 827 1889
rect 793 1787 827 1821
rect 793 1719 827 1753
rect 889 1923 923 1957
rect 889 1855 923 1889
rect 889 1787 923 1821
rect 889 1719 923 1753
rect 985 1923 1019 1957
rect 985 1855 1019 1889
rect 985 1787 1019 1821
rect 985 1719 1019 1753
rect 1081 1923 1115 1957
rect 1081 1855 1115 1889
rect 1081 1787 1115 1821
rect 1081 1719 1115 1753
rect 1177 1923 1211 1957
rect 1177 1855 1211 1889
rect 1177 1787 1211 1821
rect 1177 1719 1211 1753
rect 1273 1923 1307 1957
rect 1273 1855 1307 1889
rect 1273 1787 1307 1821
rect 1273 1719 1307 1753
rect 2466 1927 2500 1961
rect 2466 1859 2500 1893
rect 2466 1791 2500 1825
rect 2466 1723 2500 1757
rect 2562 1927 2596 1961
rect 2562 1859 2596 1893
rect 2562 1791 2596 1825
rect 2562 1723 2596 1757
rect 2658 1927 2692 1961
rect 2658 1859 2692 1893
rect 2658 1791 2692 1825
rect 2658 1723 2692 1757
rect 2754 1927 2788 1961
rect 2754 1859 2788 1893
rect 2754 1791 2788 1825
rect 2754 1723 2788 1757
rect 2850 1927 2884 1961
rect 2850 1859 2884 1893
rect 2850 1791 2884 1825
rect 2850 1723 2884 1757
rect 2946 1927 2980 1961
rect 2946 1859 2980 1893
rect 2946 1791 2980 1825
rect 2946 1723 2980 1757
rect 3042 1927 3076 1961
rect 3042 1859 3076 1893
rect 3042 1791 3076 1825
rect 3042 1723 3076 1757
rect 3138 1927 3172 1961
rect 3138 1859 3172 1893
rect 3138 1791 3172 1825
rect 3138 1723 3172 1757
rect 3234 1927 3268 1961
rect 3234 1859 3268 1893
rect 3234 1791 3268 1825
rect 3234 1723 3268 1757
rect 3330 1927 3364 1961
rect 3330 1859 3364 1893
rect 3330 1791 3364 1825
rect 3330 1723 3364 1757
rect 3426 1927 3460 1961
rect 3426 1859 3460 1893
rect 3426 1791 3460 1825
rect 3426 1723 3460 1757
rect 3987 1927 4021 1961
rect 3987 1859 4021 1893
rect 3987 1791 4021 1825
rect 3987 1723 4021 1757
rect 4083 1927 4117 1961
rect 4083 1859 4117 1893
rect 4083 1791 4117 1825
rect 4083 1723 4117 1757
rect 4179 1927 4213 1961
rect 4179 1859 4213 1893
rect 4179 1791 4213 1825
rect 4179 1723 4213 1757
rect 4275 1927 4309 1961
rect 4275 1859 4309 1893
rect 4275 1791 4309 1825
rect 4275 1723 4309 1757
rect 4371 1927 4405 1961
rect 4371 1859 4405 1893
rect 4371 1791 4405 1825
rect 4371 1723 4405 1757
rect 4467 1927 4501 1961
rect 4467 1859 4501 1893
rect 4467 1791 4501 1825
rect 4467 1723 4501 1757
rect 4563 1927 4597 1961
rect 4563 1859 4597 1893
rect 4563 1791 4597 1825
rect 4563 1723 4597 1757
rect 4659 1927 4693 1961
rect 4659 1859 4693 1893
rect 4659 1791 4693 1825
rect 4659 1723 4693 1757
rect 4755 1927 4789 1961
rect 4755 1859 4789 1893
rect 4755 1791 4789 1825
rect 4755 1723 4789 1757
rect 4851 1927 4885 1961
rect 4851 1859 4885 1893
rect 4851 1791 4885 1825
rect 4851 1723 4885 1757
rect 4947 1927 4981 1961
rect 4947 1859 4981 1893
rect 4947 1791 4981 1825
rect 4947 1723 4981 1757
rect 5356 1719 5390 1753
rect 5356 1651 5390 1685
rect 5356 1583 5390 1617
rect 5440 1719 5474 1753
rect 5440 1651 5474 1685
rect 5440 1583 5474 1617
<< psubdiff >>
rect 199 41369 317 41403
rect 351 41369 385 41403
rect 419 41369 453 41403
rect 487 41369 521 41403
rect 555 41369 589 41403
rect 623 41369 657 41403
rect 691 41369 725 41403
rect 759 41369 793 41403
rect 827 41369 861 41403
rect 895 41369 929 41403
rect 963 41369 997 41403
rect 1031 41369 1065 41403
rect 1099 41369 1133 41403
rect 1167 41369 1201 41403
rect 1235 41369 1269 41403
rect 1303 41369 1421 41403
rect 199 41293 233 41369
rect 1387 41293 1421 41369
rect 199 41225 233 41259
rect 199 41157 233 41191
rect 1387 41225 1421 41259
rect 199 41047 233 41123
rect 1387 41157 1421 41191
rect 1387 41047 1421 41123
rect 199 41013 317 41047
rect 351 41013 385 41047
rect 419 41013 453 41047
rect 487 41013 521 41047
rect 555 41013 589 41047
rect 623 41013 657 41047
rect 691 41013 725 41047
rect 759 41013 793 41047
rect 827 41013 861 41047
rect 895 41013 929 41047
rect 963 41013 997 41047
rect 1031 41013 1065 41047
rect 1099 41013 1133 41047
rect 1167 41013 1201 41047
rect 1235 41013 1269 41047
rect 1303 41013 1421 41047
rect 2352 41373 2470 41407
rect 2504 41373 2538 41407
rect 2572 41373 2606 41407
rect 2640 41373 2674 41407
rect 2708 41373 2742 41407
rect 2776 41373 2810 41407
rect 2844 41373 2878 41407
rect 2912 41373 2946 41407
rect 2980 41373 3014 41407
rect 3048 41373 3082 41407
rect 3116 41373 3150 41407
rect 3184 41373 3218 41407
rect 3252 41373 3286 41407
rect 3320 41373 3354 41407
rect 3388 41373 3422 41407
rect 3456 41373 3574 41407
rect 2352 41297 2386 41373
rect 3540 41297 3574 41373
rect 3873 41373 3991 41407
rect 4025 41373 4059 41407
rect 4093 41373 4127 41407
rect 4161 41373 4195 41407
rect 4229 41373 4263 41407
rect 4297 41373 4331 41407
rect 4365 41373 4399 41407
rect 4433 41373 4467 41407
rect 4501 41373 4535 41407
rect 4569 41373 4603 41407
rect 4637 41373 4671 41407
rect 4705 41373 4739 41407
rect 4773 41373 4807 41407
rect 4841 41373 4875 41407
rect 4909 41373 4943 41407
rect 4977 41373 5095 41407
rect 2352 41229 2386 41263
rect 2352 41161 2386 41195
rect 3540 41229 3574 41263
rect 3873 41297 3907 41373
rect 5061 41297 5095 41373
rect 3873 41229 3907 41263
rect 2352 41051 2386 41127
rect 3540 41161 3574 41195
rect 3540 41051 3574 41127
rect 2352 41017 2470 41051
rect 2504 41017 2538 41051
rect 2572 41017 2606 41051
rect 2640 41017 2674 41051
rect 2708 41017 2742 41051
rect 2776 41017 2810 41051
rect 2844 41017 2878 41051
rect 2912 41017 2946 41051
rect 2980 41017 3014 41051
rect 3048 41017 3082 41051
rect 3116 41017 3150 41051
rect 3184 41017 3218 41051
rect 3252 41017 3286 41051
rect 3320 41017 3354 41051
rect 3388 41017 3422 41051
rect 3456 41017 3574 41051
rect 3873 41161 3907 41195
rect 5061 41229 5095 41263
rect 3873 41051 3907 41127
rect 5061 41161 5095 41195
rect 5061 41051 5095 41127
rect 3873 41017 3991 41051
rect 4025 41017 4059 41051
rect 4093 41017 4127 41051
rect 4161 41017 4195 41051
rect 4229 41017 4263 41051
rect 4297 41017 4331 41051
rect 4365 41017 4399 41051
rect 4433 41017 4467 41051
rect 4501 41017 4535 41051
rect 4569 41017 4603 41051
rect 4637 41017 4671 41051
rect 4705 41017 4739 41051
rect 4773 41017 4807 41051
rect 4841 41017 4875 41051
rect 4909 41017 4943 41051
rect 4977 41017 5095 41051
rect 199 40082 317 40116
rect 351 40082 385 40116
rect 419 40082 453 40116
rect 487 40082 521 40116
rect 555 40082 589 40116
rect 623 40082 657 40116
rect 691 40082 725 40116
rect 759 40082 793 40116
rect 827 40082 861 40116
rect 895 40082 929 40116
rect 963 40082 997 40116
rect 1031 40082 1065 40116
rect 1099 40082 1133 40116
rect 1167 40082 1201 40116
rect 1235 40082 1269 40116
rect 1303 40082 1421 40116
rect 199 40006 233 40082
rect 1387 40006 1421 40082
rect 199 39938 233 39972
rect 199 39870 233 39904
rect 1387 39938 1421 39972
rect 199 39760 233 39836
rect 1387 39870 1421 39904
rect 1387 39760 1421 39836
rect 199 39726 317 39760
rect 351 39726 385 39760
rect 419 39726 453 39760
rect 487 39726 521 39760
rect 555 39726 589 39760
rect 623 39726 657 39760
rect 691 39726 725 39760
rect 759 39726 793 39760
rect 827 39726 861 39760
rect 895 39726 929 39760
rect 963 39726 997 39760
rect 1031 39726 1065 39760
rect 1099 39726 1133 39760
rect 1167 39726 1201 39760
rect 1235 39726 1269 39760
rect 1303 39726 1421 39760
rect 2352 40086 2470 40120
rect 2504 40086 2538 40120
rect 2572 40086 2606 40120
rect 2640 40086 2674 40120
rect 2708 40086 2742 40120
rect 2776 40086 2810 40120
rect 2844 40086 2878 40120
rect 2912 40086 2946 40120
rect 2980 40086 3014 40120
rect 3048 40086 3082 40120
rect 3116 40086 3150 40120
rect 3184 40086 3218 40120
rect 3252 40086 3286 40120
rect 3320 40086 3354 40120
rect 3388 40086 3422 40120
rect 3456 40086 3574 40120
rect 2352 40010 2386 40086
rect 3540 40010 3574 40086
rect 3873 40086 3991 40120
rect 4025 40086 4059 40120
rect 4093 40086 4127 40120
rect 4161 40086 4195 40120
rect 4229 40086 4263 40120
rect 4297 40086 4331 40120
rect 4365 40086 4399 40120
rect 4433 40086 4467 40120
rect 4501 40086 4535 40120
rect 4569 40086 4603 40120
rect 4637 40086 4671 40120
rect 4705 40086 4739 40120
rect 4773 40086 4807 40120
rect 4841 40086 4875 40120
rect 4909 40086 4943 40120
rect 4977 40086 5095 40120
rect 2352 39942 2386 39976
rect 2352 39874 2386 39908
rect 3540 39942 3574 39976
rect 3873 40010 3907 40086
rect 5061 40010 5095 40086
rect 3873 39942 3907 39976
rect 2352 39764 2386 39840
rect 3540 39874 3574 39908
rect 3540 39764 3574 39840
rect 2352 39730 2470 39764
rect 2504 39730 2538 39764
rect 2572 39730 2606 39764
rect 2640 39730 2674 39764
rect 2708 39730 2742 39764
rect 2776 39730 2810 39764
rect 2844 39730 2878 39764
rect 2912 39730 2946 39764
rect 2980 39730 3014 39764
rect 3048 39730 3082 39764
rect 3116 39730 3150 39764
rect 3184 39730 3218 39764
rect 3252 39730 3286 39764
rect 3320 39730 3354 39764
rect 3388 39730 3422 39764
rect 3456 39730 3574 39764
rect 3873 39874 3907 39908
rect 5061 39942 5095 39976
rect 3873 39764 3907 39840
rect 5061 39874 5095 39908
rect 5061 39764 5095 39840
rect 3873 39730 3991 39764
rect 4025 39730 4059 39764
rect 4093 39730 4127 39764
rect 4161 39730 4195 39764
rect 4229 39730 4263 39764
rect 4297 39730 4331 39764
rect 4365 39730 4399 39764
rect 4433 39730 4467 39764
rect 4501 39730 4535 39764
rect 4569 39730 4603 39764
rect 4637 39730 4671 39764
rect 4705 39730 4739 39764
rect 4773 39730 4807 39764
rect 4841 39730 4875 39764
rect 4909 39730 4943 39764
rect 4977 39730 5095 39764
rect 199 38795 317 38829
rect 351 38795 385 38829
rect 419 38795 453 38829
rect 487 38795 521 38829
rect 555 38795 589 38829
rect 623 38795 657 38829
rect 691 38795 725 38829
rect 759 38795 793 38829
rect 827 38795 861 38829
rect 895 38795 929 38829
rect 963 38795 997 38829
rect 1031 38795 1065 38829
rect 1099 38795 1133 38829
rect 1167 38795 1201 38829
rect 1235 38795 1269 38829
rect 1303 38795 1421 38829
rect 199 38719 233 38795
rect 1387 38719 1421 38795
rect 199 38651 233 38685
rect 199 38583 233 38617
rect 1387 38651 1421 38685
rect 199 38473 233 38549
rect 1387 38583 1421 38617
rect 1387 38473 1421 38549
rect 199 38439 317 38473
rect 351 38439 385 38473
rect 419 38439 453 38473
rect 487 38439 521 38473
rect 555 38439 589 38473
rect 623 38439 657 38473
rect 691 38439 725 38473
rect 759 38439 793 38473
rect 827 38439 861 38473
rect 895 38439 929 38473
rect 963 38439 997 38473
rect 1031 38439 1065 38473
rect 1099 38439 1133 38473
rect 1167 38439 1201 38473
rect 1235 38439 1269 38473
rect 1303 38439 1421 38473
rect 2352 38799 2470 38833
rect 2504 38799 2538 38833
rect 2572 38799 2606 38833
rect 2640 38799 2674 38833
rect 2708 38799 2742 38833
rect 2776 38799 2810 38833
rect 2844 38799 2878 38833
rect 2912 38799 2946 38833
rect 2980 38799 3014 38833
rect 3048 38799 3082 38833
rect 3116 38799 3150 38833
rect 3184 38799 3218 38833
rect 3252 38799 3286 38833
rect 3320 38799 3354 38833
rect 3388 38799 3422 38833
rect 3456 38799 3574 38833
rect 2352 38723 2386 38799
rect 3540 38723 3574 38799
rect 3873 38799 3991 38833
rect 4025 38799 4059 38833
rect 4093 38799 4127 38833
rect 4161 38799 4195 38833
rect 4229 38799 4263 38833
rect 4297 38799 4331 38833
rect 4365 38799 4399 38833
rect 4433 38799 4467 38833
rect 4501 38799 4535 38833
rect 4569 38799 4603 38833
rect 4637 38799 4671 38833
rect 4705 38799 4739 38833
rect 4773 38799 4807 38833
rect 4841 38799 4875 38833
rect 4909 38799 4943 38833
rect 4977 38799 5095 38833
rect 2352 38655 2386 38689
rect 2352 38587 2386 38621
rect 3540 38655 3574 38689
rect 3873 38723 3907 38799
rect 5061 38723 5095 38799
rect 3873 38655 3907 38689
rect 2352 38477 2386 38553
rect 3540 38587 3574 38621
rect 3540 38477 3574 38553
rect 2352 38443 2470 38477
rect 2504 38443 2538 38477
rect 2572 38443 2606 38477
rect 2640 38443 2674 38477
rect 2708 38443 2742 38477
rect 2776 38443 2810 38477
rect 2844 38443 2878 38477
rect 2912 38443 2946 38477
rect 2980 38443 3014 38477
rect 3048 38443 3082 38477
rect 3116 38443 3150 38477
rect 3184 38443 3218 38477
rect 3252 38443 3286 38477
rect 3320 38443 3354 38477
rect 3388 38443 3422 38477
rect 3456 38443 3574 38477
rect 3873 38587 3907 38621
rect 5061 38655 5095 38689
rect 3873 38477 3907 38553
rect 5061 38587 5095 38621
rect 5061 38477 5095 38553
rect 3873 38443 3991 38477
rect 4025 38443 4059 38477
rect 4093 38443 4127 38477
rect 4161 38443 4195 38477
rect 4229 38443 4263 38477
rect 4297 38443 4331 38477
rect 4365 38443 4399 38477
rect 4433 38443 4467 38477
rect 4501 38443 4535 38477
rect 4569 38443 4603 38477
rect 4637 38443 4671 38477
rect 4705 38443 4739 38477
rect 4773 38443 4807 38477
rect 4841 38443 4875 38477
rect 4909 38443 4943 38477
rect 4977 38443 5095 38477
rect 199 37508 317 37542
rect 351 37508 385 37542
rect 419 37508 453 37542
rect 487 37508 521 37542
rect 555 37508 589 37542
rect 623 37508 657 37542
rect 691 37508 725 37542
rect 759 37508 793 37542
rect 827 37508 861 37542
rect 895 37508 929 37542
rect 963 37508 997 37542
rect 1031 37508 1065 37542
rect 1099 37508 1133 37542
rect 1167 37508 1201 37542
rect 1235 37508 1269 37542
rect 1303 37508 1421 37542
rect 199 37432 233 37508
rect 1387 37432 1421 37508
rect 199 37364 233 37398
rect 199 37296 233 37330
rect 1387 37364 1421 37398
rect 199 37186 233 37262
rect 1387 37296 1421 37330
rect 1387 37186 1421 37262
rect 199 37152 317 37186
rect 351 37152 385 37186
rect 419 37152 453 37186
rect 487 37152 521 37186
rect 555 37152 589 37186
rect 623 37152 657 37186
rect 691 37152 725 37186
rect 759 37152 793 37186
rect 827 37152 861 37186
rect 895 37152 929 37186
rect 963 37152 997 37186
rect 1031 37152 1065 37186
rect 1099 37152 1133 37186
rect 1167 37152 1201 37186
rect 1235 37152 1269 37186
rect 1303 37152 1421 37186
rect 2352 37512 2470 37546
rect 2504 37512 2538 37546
rect 2572 37512 2606 37546
rect 2640 37512 2674 37546
rect 2708 37512 2742 37546
rect 2776 37512 2810 37546
rect 2844 37512 2878 37546
rect 2912 37512 2946 37546
rect 2980 37512 3014 37546
rect 3048 37512 3082 37546
rect 3116 37512 3150 37546
rect 3184 37512 3218 37546
rect 3252 37512 3286 37546
rect 3320 37512 3354 37546
rect 3388 37512 3422 37546
rect 3456 37512 3574 37546
rect 2352 37436 2386 37512
rect 3540 37436 3574 37512
rect 3873 37512 3991 37546
rect 4025 37512 4059 37546
rect 4093 37512 4127 37546
rect 4161 37512 4195 37546
rect 4229 37512 4263 37546
rect 4297 37512 4331 37546
rect 4365 37512 4399 37546
rect 4433 37512 4467 37546
rect 4501 37512 4535 37546
rect 4569 37512 4603 37546
rect 4637 37512 4671 37546
rect 4705 37512 4739 37546
rect 4773 37512 4807 37546
rect 4841 37512 4875 37546
rect 4909 37512 4943 37546
rect 4977 37512 5095 37546
rect 2352 37368 2386 37402
rect 2352 37300 2386 37334
rect 3540 37368 3574 37402
rect 3873 37436 3907 37512
rect 5061 37436 5095 37512
rect 3873 37368 3907 37402
rect 2352 37190 2386 37266
rect 3540 37300 3574 37334
rect 3540 37190 3574 37266
rect 2352 37156 2470 37190
rect 2504 37156 2538 37190
rect 2572 37156 2606 37190
rect 2640 37156 2674 37190
rect 2708 37156 2742 37190
rect 2776 37156 2810 37190
rect 2844 37156 2878 37190
rect 2912 37156 2946 37190
rect 2980 37156 3014 37190
rect 3048 37156 3082 37190
rect 3116 37156 3150 37190
rect 3184 37156 3218 37190
rect 3252 37156 3286 37190
rect 3320 37156 3354 37190
rect 3388 37156 3422 37190
rect 3456 37156 3574 37190
rect 3873 37300 3907 37334
rect 5061 37368 5095 37402
rect 3873 37190 3907 37266
rect 5061 37300 5095 37334
rect 5061 37190 5095 37266
rect 3873 37156 3991 37190
rect 4025 37156 4059 37190
rect 4093 37156 4127 37190
rect 4161 37156 4195 37190
rect 4229 37156 4263 37190
rect 4297 37156 4331 37190
rect 4365 37156 4399 37190
rect 4433 37156 4467 37190
rect 4501 37156 4535 37190
rect 4569 37156 4603 37190
rect 4637 37156 4671 37190
rect 4705 37156 4739 37190
rect 4773 37156 4807 37190
rect 4841 37156 4875 37190
rect 4909 37156 4943 37190
rect 4977 37156 5095 37190
rect 199 36221 317 36255
rect 351 36221 385 36255
rect 419 36221 453 36255
rect 487 36221 521 36255
rect 555 36221 589 36255
rect 623 36221 657 36255
rect 691 36221 725 36255
rect 759 36221 793 36255
rect 827 36221 861 36255
rect 895 36221 929 36255
rect 963 36221 997 36255
rect 1031 36221 1065 36255
rect 1099 36221 1133 36255
rect 1167 36221 1201 36255
rect 1235 36221 1269 36255
rect 1303 36221 1421 36255
rect 199 36145 233 36221
rect 1387 36145 1421 36221
rect 199 36077 233 36111
rect 199 36009 233 36043
rect 1387 36077 1421 36111
rect 199 35899 233 35975
rect 1387 36009 1421 36043
rect 1387 35899 1421 35975
rect 199 35865 317 35899
rect 351 35865 385 35899
rect 419 35865 453 35899
rect 487 35865 521 35899
rect 555 35865 589 35899
rect 623 35865 657 35899
rect 691 35865 725 35899
rect 759 35865 793 35899
rect 827 35865 861 35899
rect 895 35865 929 35899
rect 963 35865 997 35899
rect 1031 35865 1065 35899
rect 1099 35865 1133 35899
rect 1167 35865 1201 35899
rect 1235 35865 1269 35899
rect 1303 35865 1421 35899
rect 2352 36225 2470 36259
rect 2504 36225 2538 36259
rect 2572 36225 2606 36259
rect 2640 36225 2674 36259
rect 2708 36225 2742 36259
rect 2776 36225 2810 36259
rect 2844 36225 2878 36259
rect 2912 36225 2946 36259
rect 2980 36225 3014 36259
rect 3048 36225 3082 36259
rect 3116 36225 3150 36259
rect 3184 36225 3218 36259
rect 3252 36225 3286 36259
rect 3320 36225 3354 36259
rect 3388 36225 3422 36259
rect 3456 36225 3574 36259
rect 2352 36149 2386 36225
rect 3540 36149 3574 36225
rect 3873 36225 3991 36259
rect 4025 36225 4059 36259
rect 4093 36225 4127 36259
rect 4161 36225 4195 36259
rect 4229 36225 4263 36259
rect 4297 36225 4331 36259
rect 4365 36225 4399 36259
rect 4433 36225 4467 36259
rect 4501 36225 4535 36259
rect 4569 36225 4603 36259
rect 4637 36225 4671 36259
rect 4705 36225 4739 36259
rect 4773 36225 4807 36259
rect 4841 36225 4875 36259
rect 4909 36225 4943 36259
rect 4977 36225 5095 36259
rect 2352 36081 2386 36115
rect 2352 36013 2386 36047
rect 3540 36081 3574 36115
rect 3873 36149 3907 36225
rect 5061 36149 5095 36225
rect 3873 36081 3907 36115
rect 2352 35903 2386 35979
rect 3540 36013 3574 36047
rect 3540 35903 3574 35979
rect 2352 35869 2470 35903
rect 2504 35869 2538 35903
rect 2572 35869 2606 35903
rect 2640 35869 2674 35903
rect 2708 35869 2742 35903
rect 2776 35869 2810 35903
rect 2844 35869 2878 35903
rect 2912 35869 2946 35903
rect 2980 35869 3014 35903
rect 3048 35869 3082 35903
rect 3116 35869 3150 35903
rect 3184 35869 3218 35903
rect 3252 35869 3286 35903
rect 3320 35869 3354 35903
rect 3388 35869 3422 35903
rect 3456 35869 3574 35903
rect 3873 36013 3907 36047
rect 5061 36081 5095 36115
rect 3873 35903 3907 35979
rect 5061 36013 5095 36047
rect 5061 35903 5095 35979
rect 3873 35869 3991 35903
rect 4025 35869 4059 35903
rect 4093 35869 4127 35903
rect 4161 35869 4195 35903
rect 4229 35869 4263 35903
rect 4297 35869 4331 35903
rect 4365 35869 4399 35903
rect 4433 35869 4467 35903
rect 4501 35869 4535 35903
rect 4569 35869 4603 35903
rect 4637 35869 4671 35903
rect 4705 35869 4739 35903
rect 4773 35869 4807 35903
rect 4841 35869 4875 35903
rect 4909 35869 4943 35903
rect 4977 35869 5095 35903
rect 199 34934 317 34968
rect 351 34934 385 34968
rect 419 34934 453 34968
rect 487 34934 521 34968
rect 555 34934 589 34968
rect 623 34934 657 34968
rect 691 34934 725 34968
rect 759 34934 793 34968
rect 827 34934 861 34968
rect 895 34934 929 34968
rect 963 34934 997 34968
rect 1031 34934 1065 34968
rect 1099 34934 1133 34968
rect 1167 34934 1201 34968
rect 1235 34934 1269 34968
rect 1303 34934 1421 34968
rect 199 34858 233 34934
rect 1387 34858 1421 34934
rect 199 34790 233 34824
rect 199 34722 233 34756
rect 1387 34790 1421 34824
rect 199 34612 233 34688
rect 1387 34722 1421 34756
rect 1387 34612 1421 34688
rect 199 34578 317 34612
rect 351 34578 385 34612
rect 419 34578 453 34612
rect 487 34578 521 34612
rect 555 34578 589 34612
rect 623 34578 657 34612
rect 691 34578 725 34612
rect 759 34578 793 34612
rect 827 34578 861 34612
rect 895 34578 929 34612
rect 963 34578 997 34612
rect 1031 34578 1065 34612
rect 1099 34578 1133 34612
rect 1167 34578 1201 34612
rect 1235 34578 1269 34612
rect 1303 34578 1421 34612
rect 2352 34938 2470 34972
rect 2504 34938 2538 34972
rect 2572 34938 2606 34972
rect 2640 34938 2674 34972
rect 2708 34938 2742 34972
rect 2776 34938 2810 34972
rect 2844 34938 2878 34972
rect 2912 34938 2946 34972
rect 2980 34938 3014 34972
rect 3048 34938 3082 34972
rect 3116 34938 3150 34972
rect 3184 34938 3218 34972
rect 3252 34938 3286 34972
rect 3320 34938 3354 34972
rect 3388 34938 3422 34972
rect 3456 34938 3574 34972
rect 2352 34862 2386 34938
rect 3540 34862 3574 34938
rect 3873 34938 3991 34972
rect 4025 34938 4059 34972
rect 4093 34938 4127 34972
rect 4161 34938 4195 34972
rect 4229 34938 4263 34972
rect 4297 34938 4331 34972
rect 4365 34938 4399 34972
rect 4433 34938 4467 34972
rect 4501 34938 4535 34972
rect 4569 34938 4603 34972
rect 4637 34938 4671 34972
rect 4705 34938 4739 34972
rect 4773 34938 4807 34972
rect 4841 34938 4875 34972
rect 4909 34938 4943 34972
rect 4977 34938 5095 34972
rect 2352 34794 2386 34828
rect 2352 34726 2386 34760
rect 3540 34794 3574 34828
rect 3873 34862 3907 34938
rect 5061 34862 5095 34938
rect 3873 34794 3907 34828
rect 2352 34616 2386 34692
rect 3540 34726 3574 34760
rect 3540 34616 3574 34692
rect 2352 34582 2470 34616
rect 2504 34582 2538 34616
rect 2572 34582 2606 34616
rect 2640 34582 2674 34616
rect 2708 34582 2742 34616
rect 2776 34582 2810 34616
rect 2844 34582 2878 34616
rect 2912 34582 2946 34616
rect 2980 34582 3014 34616
rect 3048 34582 3082 34616
rect 3116 34582 3150 34616
rect 3184 34582 3218 34616
rect 3252 34582 3286 34616
rect 3320 34582 3354 34616
rect 3388 34582 3422 34616
rect 3456 34582 3574 34616
rect 3873 34726 3907 34760
rect 5061 34794 5095 34828
rect 3873 34616 3907 34692
rect 5061 34726 5095 34760
rect 5061 34616 5095 34692
rect 3873 34582 3991 34616
rect 4025 34582 4059 34616
rect 4093 34582 4127 34616
rect 4161 34582 4195 34616
rect 4229 34582 4263 34616
rect 4297 34582 4331 34616
rect 4365 34582 4399 34616
rect 4433 34582 4467 34616
rect 4501 34582 4535 34616
rect 4569 34582 4603 34616
rect 4637 34582 4671 34616
rect 4705 34582 4739 34616
rect 4773 34582 4807 34616
rect 4841 34582 4875 34616
rect 4909 34582 4943 34616
rect 4977 34582 5095 34616
rect 199 33647 317 33681
rect 351 33647 385 33681
rect 419 33647 453 33681
rect 487 33647 521 33681
rect 555 33647 589 33681
rect 623 33647 657 33681
rect 691 33647 725 33681
rect 759 33647 793 33681
rect 827 33647 861 33681
rect 895 33647 929 33681
rect 963 33647 997 33681
rect 1031 33647 1065 33681
rect 1099 33647 1133 33681
rect 1167 33647 1201 33681
rect 1235 33647 1269 33681
rect 1303 33647 1421 33681
rect 199 33571 233 33647
rect 1387 33571 1421 33647
rect 199 33503 233 33537
rect 199 33435 233 33469
rect 1387 33503 1421 33537
rect 199 33325 233 33401
rect 1387 33435 1421 33469
rect 1387 33325 1421 33401
rect 199 33291 317 33325
rect 351 33291 385 33325
rect 419 33291 453 33325
rect 487 33291 521 33325
rect 555 33291 589 33325
rect 623 33291 657 33325
rect 691 33291 725 33325
rect 759 33291 793 33325
rect 827 33291 861 33325
rect 895 33291 929 33325
rect 963 33291 997 33325
rect 1031 33291 1065 33325
rect 1099 33291 1133 33325
rect 1167 33291 1201 33325
rect 1235 33291 1269 33325
rect 1303 33291 1421 33325
rect 2352 33651 2470 33685
rect 2504 33651 2538 33685
rect 2572 33651 2606 33685
rect 2640 33651 2674 33685
rect 2708 33651 2742 33685
rect 2776 33651 2810 33685
rect 2844 33651 2878 33685
rect 2912 33651 2946 33685
rect 2980 33651 3014 33685
rect 3048 33651 3082 33685
rect 3116 33651 3150 33685
rect 3184 33651 3218 33685
rect 3252 33651 3286 33685
rect 3320 33651 3354 33685
rect 3388 33651 3422 33685
rect 3456 33651 3574 33685
rect 2352 33575 2386 33651
rect 3540 33575 3574 33651
rect 3873 33651 3991 33685
rect 4025 33651 4059 33685
rect 4093 33651 4127 33685
rect 4161 33651 4195 33685
rect 4229 33651 4263 33685
rect 4297 33651 4331 33685
rect 4365 33651 4399 33685
rect 4433 33651 4467 33685
rect 4501 33651 4535 33685
rect 4569 33651 4603 33685
rect 4637 33651 4671 33685
rect 4705 33651 4739 33685
rect 4773 33651 4807 33685
rect 4841 33651 4875 33685
rect 4909 33651 4943 33685
rect 4977 33651 5095 33685
rect 2352 33507 2386 33541
rect 2352 33439 2386 33473
rect 3540 33507 3574 33541
rect 3873 33575 3907 33651
rect 5061 33575 5095 33651
rect 3873 33507 3907 33541
rect 2352 33329 2386 33405
rect 3540 33439 3574 33473
rect 3540 33329 3574 33405
rect 2352 33295 2470 33329
rect 2504 33295 2538 33329
rect 2572 33295 2606 33329
rect 2640 33295 2674 33329
rect 2708 33295 2742 33329
rect 2776 33295 2810 33329
rect 2844 33295 2878 33329
rect 2912 33295 2946 33329
rect 2980 33295 3014 33329
rect 3048 33295 3082 33329
rect 3116 33295 3150 33329
rect 3184 33295 3218 33329
rect 3252 33295 3286 33329
rect 3320 33295 3354 33329
rect 3388 33295 3422 33329
rect 3456 33295 3574 33329
rect 3873 33439 3907 33473
rect 5061 33507 5095 33541
rect 3873 33329 3907 33405
rect 5061 33439 5095 33473
rect 5061 33329 5095 33405
rect 3873 33295 3991 33329
rect 4025 33295 4059 33329
rect 4093 33295 4127 33329
rect 4161 33295 4195 33329
rect 4229 33295 4263 33329
rect 4297 33295 4331 33329
rect 4365 33295 4399 33329
rect 4433 33295 4467 33329
rect 4501 33295 4535 33329
rect 4569 33295 4603 33329
rect 4637 33295 4671 33329
rect 4705 33295 4739 33329
rect 4773 33295 4807 33329
rect 4841 33295 4875 33329
rect 4909 33295 4943 33329
rect 4977 33295 5095 33329
rect 199 32360 317 32394
rect 351 32360 385 32394
rect 419 32360 453 32394
rect 487 32360 521 32394
rect 555 32360 589 32394
rect 623 32360 657 32394
rect 691 32360 725 32394
rect 759 32360 793 32394
rect 827 32360 861 32394
rect 895 32360 929 32394
rect 963 32360 997 32394
rect 1031 32360 1065 32394
rect 1099 32360 1133 32394
rect 1167 32360 1201 32394
rect 1235 32360 1269 32394
rect 1303 32360 1421 32394
rect 199 32284 233 32360
rect 1387 32284 1421 32360
rect 199 32216 233 32250
rect 199 32148 233 32182
rect 1387 32216 1421 32250
rect 199 32038 233 32114
rect 1387 32148 1421 32182
rect 1387 32038 1421 32114
rect 199 32004 317 32038
rect 351 32004 385 32038
rect 419 32004 453 32038
rect 487 32004 521 32038
rect 555 32004 589 32038
rect 623 32004 657 32038
rect 691 32004 725 32038
rect 759 32004 793 32038
rect 827 32004 861 32038
rect 895 32004 929 32038
rect 963 32004 997 32038
rect 1031 32004 1065 32038
rect 1099 32004 1133 32038
rect 1167 32004 1201 32038
rect 1235 32004 1269 32038
rect 1303 32004 1421 32038
rect 2352 32364 2470 32398
rect 2504 32364 2538 32398
rect 2572 32364 2606 32398
rect 2640 32364 2674 32398
rect 2708 32364 2742 32398
rect 2776 32364 2810 32398
rect 2844 32364 2878 32398
rect 2912 32364 2946 32398
rect 2980 32364 3014 32398
rect 3048 32364 3082 32398
rect 3116 32364 3150 32398
rect 3184 32364 3218 32398
rect 3252 32364 3286 32398
rect 3320 32364 3354 32398
rect 3388 32364 3422 32398
rect 3456 32364 3574 32398
rect 2352 32288 2386 32364
rect 3540 32288 3574 32364
rect 3873 32364 3991 32398
rect 4025 32364 4059 32398
rect 4093 32364 4127 32398
rect 4161 32364 4195 32398
rect 4229 32364 4263 32398
rect 4297 32364 4331 32398
rect 4365 32364 4399 32398
rect 4433 32364 4467 32398
rect 4501 32364 4535 32398
rect 4569 32364 4603 32398
rect 4637 32364 4671 32398
rect 4705 32364 4739 32398
rect 4773 32364 4807 32398
rect 4841 32364 4875 32398
rect 4909 32364 4943 32398
rect 4977 32364 5095 32398
rect 2352 32220 2386 32254
rect 2352 32152 2386 32186
rect 3540 32220 3574 32254
rect 3873 32288 3907 32364
rect 5061 32288 5095 32364
rect 3873 32220 3907 32254
rect 2352 32042 2386 32118
rect 3540 32152 3574 32186
rect 3540 32042 3574 32118
rect 2352 32008 2470 32042
rect 2504 32008 2538 32042
rect 2572 32008 2606 32042
rect 2640 32008 2674 32042
rect 2708 32008 2742 32042
rect 2776 32008 2810 32042
rect 2844 32008 2878 32042
rect 2912 32008 2946 32042
rect 2980 32008 3014 32042
rect 3048 32008 3082 32042
rect 3116 32008 3150 32042
rect 3184 32008 3218 32042
rect 3252 32008 3286 32042
rect 3320 32008 3354 32042
rect 3388 32008 3422 32042
rect 3456 32008 3574 32042
rect 3873 32152 3907 32186
rect 5061 32220 5095 32254
rect 3873 32042 3907 32118
rect 5061 32152 5095 32186
rect 5061 32042 5095 32118
rect 3873 32008 3991 32042
rect 4025 32008 4059 32042
rect 4093 32008 4127 32042
rect 4161 32008 4195 32042
rect 4229 32008 4263 32042
rect 4297 32008 4331 32042
rect 4365 32008 4399 32042
rect 4433 32008 4467 32042
rect 4501 32008 4535 32042
rect 4569 32008 4603 32042
rect 4637 32008 4671 32042
rect 4705 32008 4739 32042
rect 4773 32008 4807 32042
rect 4841 32008 4875 32042
rect 4909 32008 4943 32042
rect 4977 32008 5095 32042
rect 199 31073 317 31107
rect 351 31073 385 31107
rect 419 31073 453 31107
rect 487 31073 521 31107
rect 555 31073 589 31107
rect 623 31073 657 31107
rect 691 31073 725 31107
rect 759 31073 793 31107
rect 827 31073 861 31107
rect 895 31073 929 31107
rect 963 31073 997 31107
rect 1031 31073 1065 31107
rect 1099 31073 1133 31107
rect 1167 31073 1201 31107
rect 1235 31073 1269 31107
rect 1303 31073 1421 31107
rect 199 30997 233 31073
rect 1387 30997 1421 31073
rect 199 30929 233 30963
rect 199 30861 233 30895
rect 1387 30929 1421 30963
rect 199 30751 233 30827
rect 1387 30861 1421 30895
rect 1387 30751 1421 30827
rect 199 30717 317 30751
rect 351 30717 385 30751
rect 419 30717 453 30751
rect 487 30717 521 30751
rect 555 30717 589 30751
rect 623 30717 657 30751
rect 691 30717 725 30751
rect 759 30717 793 30751
rect 827 30717 861 30751
rect 895 30717 929 30751
rect 963 30717 997 30751
rect 1031 30717 1065 30751
rect 1099 30717 1133 30751
rect 1167 30717 1201 30751
rect 1235 30717 1269 30751
rect 1303 30717 1421 30751
rect 2352 31077 2470 31111
rect 2504 31077 2538 31111
rect 2572 31077 2606 31111
rect 2640 31077 2674 31111
rect 2708 31077 2742 31111
rect 2776 31077 2810 31111
rect 2844 31077 2878 31111
rect 2912 31077 2946 31111
rect 2980 31077 3014 31111
rect 3048 31077 3082 31111
rect 3116 31077 3150 31111
rect 3184 31077 3218 31111
rect 3252 31077 3286 31111
rect 3320 31077 3354 31111
rect 3388 31077 3422 31111
rect 3456 31077 3574 31111
rect 2352 31001 2386 31077
rect 3540 31001 3574 31077
rect 3873 31077 3991 31111
rect 4025 31077 4059 31111
rect 4093 31077 4127 31111
rect 4161 31077 4195 31111
rect 4229 31077 4263 31111
rect 4297 31077 4331 31111
rect 4365 31077 4399 31111
rect 4433 31077 4467 31111
rect 4501 31077 4535 31111
rect 4569 31077 4603 31111
rect 4637 31077 4671 31111
rect 4705 31077 4739 31111
rect 4773 31077 4807 31111
rect 4841 31077 4875 31111
rect 4909 31077 4943 31111
rect 4977 31077 5095 31111
rect 2352 30933 2386 30967
rect 2352 30865 2386 30899
rect 3540 30933 3574 30967
rect 3873 31001 3907 31077
rect 5061 31001 5095 31077
rect 3873 30933 3907 30967
rect 2352 30755 2386 30831
rect 3540 30865 3574 30899
rect 3540 30755 3574 30831
rect 2352 30721 2470 30755
rect 2504 30721 2538 30755
rect 2572 30721 2606 30755
rect 2640 30721 2674 30755
rect 2708 30721 2742 30755
rect 2776 30721 2810 30755
rect 2844 30721 2878 30755
rect 2912 30721 2946 30755
rect 2980 30721 3014 30755
rect 3048 30721 3082 30755
rect 3116 30721 3150 30755
rect 3184 30721 3218 30755
rect 3252 30721 3286 30755
rect 3320 30721 3354 30755
rect 3388 30721 3422 30755
rect 3456 30721 3574 30755
rect 3873 30865 3907 30899
rect 5061 30933 5095 30967
rect 3873 30755 3907 30831
rect 5061 30865 5095 30899
rect 5061 30755 5095 30831
rect 3873 30721 3991 30755
rect 4025 30721 4059 30755
rect 4093 30721 4127 30755
rect 4161 30721 4195 30755
rect 4229 30721 4263 30755
rect 4297 30721 4331 30755
rect 4365 30721 4399 30755
rect 4433 30721 4467 30755
rect 4501 30721 4535 30755
rect 4569 30721 4603 30755
rect 4637 30721 4671 30755
rect 4705 30721 4739 30755
rect 4773 30721 4807 30755
rect 4841 30721 4875 30755
rect 4909 30721 4943 30755
rect 4977 30721 5095 30755
rect 199 29786 317 29820
rect 351 29786 385 29820
rect 419 29786 453 29820
rect 487 29786 521 29820
rect 555 29786 589 29820
rect 623 29786 657 29820
rect 691 29786 725 29820
rect 759 29786 793 29820
rect 827 29786 861 29820
rect 895 29786 929 29820
rect 963 29786 997 29820
rect 1031 29786 1065 29820
rect 1099 29786 1133 29820
rect 1167 29786 1201 29820
rect 1235 29786 1269 29820
rect 1303 29786 1421 29820
rect 199 29710 233 29786
rect 1387 29710 1421 29786
rect 199 29642 233 29676
rect 199 29574 233 29608
rect 1387 29642 1421 29676
rect 199 29464 233 29540
rect 1387 29574 1421 29608
rect 1387 29464 1421 29540
rect 199 29430 317 29464
rect 351 29430 385 29464
rect 419 29430 453 29464
rect 487 29430 521 29464
rect 555 29430 589 29464
rect 623 29430 657 29464
rect 691 29430 725 29464
rect 759 29430 793 29464
rect 827 29430 861 29464
rect 895 29430 929 29464
rect 963 29430 997 29464
rect 1031 29430 1065 29464
rect 1099 29430 1133 29464
rect 1167 29430 1201 29464
rect 1235 29430 1269 29464
rect 1303 29430 1421 29464
rect 2352 29790 2470 29824
rect 2504 29790 2538 29824
rect 2572 29790 2606 29824
rect 2640 29790 2674 29824
rect 2708 29790 2742 29824
rect 2776 29790 2810 29824
rect 2844 29790 2878 29824
rect 2912 29790 2946 29824
rect 2980 29790 3014 29824
rect 3048 29790 3082 29824
rect 3116 29790 3150 29824
rect 3184 29790 3218 29824
rect 3252 29790 3286 29824
rect 3320 29790 3354 29824
rect 3388 29790 3422 29824
rect 3456 29790 3574 29824
rect 2352 29714 2386 29790
rect 3540 29714 3574 29790
rect 3873 29790 3991 29824
rect 4025 29790 4059 29824
rect 4093 29790 4127 29824
rect 4161 29790 4195 29824
rect 4229 29790 4263 29824
rect 4297 29790 4331 29824
rect 4365 29790 4399 29824
rect 4433 29790 4467 29824
rect 4501 29790 4535 29824
rect 4569 29790 4603 29824
rect 4637 29790 4671 29824
rect 4705 29790 4739 29824
rect 4773 29790 4807 29824
rect 4841 29790 4875 29824
rect 4909 29790 4943 29824
rect 4977 29790 5095 29824
rect 2352 29646 2386 29680
rect 2352 29578 2386 29612
rect 3540 29646 3574 29680
rect 3873 29714 3907 29790
rect 5061 29714 5095 29790
rect 3873 29646 3907 29680
rect 2352 29468 2386 29544
rect 3540 29578 3574 29612
rect 3540 29468 3574 29544
rect 2352 29434 2470 29468
rect 2504 29434 2538 29468
rect 2572 29434 2606 29468
rect 2640 29434 2674 29468
rect 2708 29434 2742 29468
rect 2776 29434 2810 29468
rect 2844 29434 2878 29468
rect 2912 29434 2946 29468
rect 2980 29434 3014 29468
rect 3048 29434 3082 29468
rect 3116 29434 3150 29468
rect 3184 29434 3218 29468
rect 3252 29434 3286 29468
rect 3320 29434 3354 29468
rect 3388 29434 3422 29468
rect 3456 29434 3574 29468
rect 3873 29578 3907 29612
rect 5061 29646 5095 29680
rect 3873 29468 3907 29544
rect 5061 29578 5095 29612
rect 5061 29468 5095 29544
rect 3873 29434 3991 29468
rect 4025 29434 4059 29468
rect 4093 29434 4127 29468
rect 4161 29434 4195 29468
rect 4229 29434 4263 29468
rect 4297 29434 4331 29468
rect 4365 29434 4399 29468
rect 4433 29434 4467 29468
rect 4501 29434 4535 29468
rect 4569 29434 4603 29468
rect 4637 29434 4671 29468
rect 4705 29434 4739 29468
rect 4773 29434 4807 29468
rect 4841 29434 4875 29468
rect 4909 29434 4943 29468
rect 4977 29434 5095 29468
rect 199 28499 317 28533
rect 351 28499 385 28533
rect 419 28499 453 28533
rect 487 28499 521 28533
rect 555 28499 589 28533
rect 623 28499 657 28533
rect 691 28499 725 28533
rect 759 28499 793 28533
rect 827 28499 861 28533
rect 895 28499 929 28533
rect 963 28499 997 28533
rect 1031 28499 1065 28533
rect 1099 28499 1133 28533
rect 1167 28499 1201 28533
rect 1235 28499 1269 28533
rect 1303 28499 1421 28533
rect 199 28423 233 28499
rect 1387 28423 1421 28499
rect 199 28355 233 28389
rect 199 28287 233 28321
rect 1387 28355 1421 28389
rect 199 28177 233 28253
rect 1387 28287 1421 28321
rect 1387 28177 1421 28253
rect 199 28143 317 28177
rect 351 28143 385 28177
rect 419 28143 453 28177
rect 487 28143 521 28177
rect 555 28143 589 28177
rect 623 28143 657 28177
rect 691 28143 725 28177
rect 759 28143 793 28177
rect 827 28143 861 28177
rect 895 28143 929 28177
rect 963 28143 997 28177
rect 1031 28143 1065 28177
rect 1099 28143 1133 28177
rect 1167 28143 1201 28177
rect 1235 28143 1269 28177
rect 1303 28143 1421 28177
rect 2352 28503 2470 28537
rect 2504 28503 2538 28537
rect 2572 28503 2606 28537
rect 2640 28503 2674 28537
rect 2708 28503 2742 28537
rect 2776 28503 2810 28537
rect 2844 28503 2878 28537
rect 2912 28503 2946 28537
rect 2980 28503 3014 28537
rect 3048 28503 3082 28537
rect 3116 28503 3150 28537
rect 3184 28503 3218 28537
rect 3252 28503 3286 28537
rect 3320 28503 3354 28537
rect 3388 28503 3422 28537
rect 3456 28503 3574 28537
rect 2352 28427 2386 28503
rect 3540 28427 3574 28503
rect 3873 28503 3991 28537
rect 4025 28503 4059 28537
rect 4093 28503 4127 28537
rect 4161 28503 4195 28537
rect 4229 28503 4263 28537
rect 4297 28503 4331 28537
rect 4365 28503 4399 28537
rect 4433 28503 4467 28537
rect 4501 28503 4535 28537
rect 4569 28503 4603 28537
rect 4637 28503 4671 28537
rect 4705 28503 4739 28537
rect 4773 28503 4807 28537
rect 4841 28503 4875 28537
rect 4909 28503 4943 28537
rect 4977 28503 5095 28537
rect 2352 28359 2386 28393
rect 2352 28291 2386 28325
rect 3540 28359 3574 28393
rect 3873 28427 3907 28503
rect 5061 28427 5095 28503
rect 3873 28359 3907 28393
rect 2352 28181 2386 28257
rect 3540 28291 3574 28325
rect 3540 28181 3574 28257
rect 2352 28147 2470 28181
rect 2504 28147 2538 28181
rect 2572 28147 2606 28181
rect 2640 28147 2674 28181
rect 2708 28147 2742 28181
rect 2776 28147 2810 28181
rect 2844 28147 2878 28181
rect 2912 28147 2946 28181
rect 2980 28147 3014 28181
rect 3048 28147 3082 28181
rect 3116 28147 3150 28181
rect 3184 28147 3218 28181
rect 3252 28147 3286 28181
rect 3320 28147 3354 28181
rect 3388 28147 3422 28181
rect 3456 28147 3574 28181
rect 3873 28291 3907 28325
rect 5061 28359 5095 28393
rect 3873 28181 3907 28257
rect 5061 28291 5095 28325
rect 5061 28181 5095 28257
rect 3873 28147 3991 28181
rect 4025 28147 4059 28181
rect 4093 28147 4127 28181
rect 4161 28147 4195 28181
rect 4229 28147 4263 28181
rect 4297 28147 4331 28181
rect 4365 28147 4399 28181
rect 4433 28147 4467 28181
rect 4501 28147 4535 28181
rect 4569 28147 4603 28181
rect 4637 28147 4671 28181
rect 4705 28147 4739 28181
rect 4773 28147 4807 28181
rect 4841 28147 4875 28181
rect 4909 28147 4943 28181
rect 4977 28147 5095 28181
rect 199 27212 317 27246
rect 351 27212 385 27246
rect 419 27212 453 27246
rect 487 27212 521 27246
rect 555 27212 589 27246
rect 623 27212 657 27246
rect 691 27212 725 27246
rect 759 27212 793 27246
rect 827 27212 861 27246
rect 895 27212 929 27246
rect 963 27212 997 27246
rect 1031 27212 1065 27246
rect 1099 27212 1133 27246
rect 1167 27212 1201 27246
rect 1235 27212 1269 27246
rect 1303 27212 1421 27246
rect 199 27136 233 27212
rect 1387 27136 1421 27212
rect 199 27068 233 27102
rect 199 27000 233 27034
rect 1387 27068 1421 27102
rect 199 26890 233 26966
rect 1387 27000 1421 27034
rect 1387 26890 1421 26966
rect 199 26856 317 26890
rect 351 26856 385 26890
rect 419 26856 453 26890
rect 487 26856 521 26890
rect 555 26856 589 26890
rect 623 26856 657 26890
rect 691 26856 725 26890
rect 759 26856 793 26890
rect 827 26856 861 26890
rect 895 26856 929 26890
rect 963 26856 997 26890
rect 1031 26856 1065 26890
rect 1099 26856 1133 26890
rect 1167 26856 1201 26890
rect 1235 26856 1269 26890
rect 1303 26856 1421 26890
rect 2352 27216 2470 27250
rect 2504 27216 2538 27250
rect 2572 27216 2606 27250
rect 2640 27216 2674 27250
rect 2708 27216 2742 27250
rect 2776 27216 2810 27250
rect 2844 27216 2878 27250
rect 2912 27216 2946 27250
rect 2980 27216 3014 27250
rect 3048 27216 3082 27250
rect 3116 27216 3150 27250
rect 3184 27216 3218 27250
rect 3252 27216 3286 27250
rect 3320 27216 3354 27250
rect 3388 27216 3422 27250
rect 3456 27216 3574 27250
rect 2352 27140 2386 27216
rect 3540 27140 3574 27216
rect 3873 27216 3991 27250
rect 4025 27216 4059 27250
rect 4093 27216 4127 27250
rect 4161 27216 4195 27250
rect 4229 27216 4263 27250
rect 4297 27216 4331 27250
rect 4365 27216 4399 27250
rect 4433 27216 4467 27250
rect 4501 27216 4535 27250
rect 4569 27216 4603 27250
rect 4637 27216 4671 27250
rect 4705 27216 4739 27250
rect 4773 27216 4807 27250
rect 4841 27216 4875 27250
rect 4909 27216 4943 27250
rect 4977 27216 5095 27250
rect 2352 27072 2386 27106
rect 2352 27004 2386 27038
rect 3540 27072 3574 27106
rect 3873 27140 3907 27216
rect 5061 27140 5095 27216
rect 3873 27072 3907 27106
rect 2352 26894 2386 26970
rect 3540 27004 3574 27038
rect 3540 26894 3574 26970
rect 2352 26860 2470 26894
rect 2504 26860 2538 26894
rect 2572 26860 2606 26894
rect 2640 26860 2674 26894
rect 2708 26860 2742 26894
rect 2776 26860 2810 26894
rect 2844 26860 2878 26894
rect 2912 26860 2946 26894
rect 2980 26860 3014 26894
rect 3048 26860 3082 26894
rect 3116 26860 3150 26894
rect 3184 26860 3218 26894
rect 3252 26860 3286 26894
rect 3320 26860 3354 26894
rect 3388 26860 3422 26894
rect 3456 26860 3574 26894
rect 3873 27004 3907 27038
rect 5061 27072 5095 27106
rect 3873 26894 3907 26970
rect 5061 27004 5095 27038
rect 5061 26894 5095 26970
rect 3873 26860 3991 26894
rect 4025 26860 4059 26894
rect 4093 26860 4127 26894
rect 4161 26860 4195 26894
rect 4229 26860 4263 26894
rect 4297 26860 4331 26894
rect 4365 26860 4399 26894
rect 4433 26860 4467 26894
rect 4501 26860 4535 26894
rect 4569 26860 4603 26894
rect 4637 26860 4671 26894
rect 4705 26860 4739 26894
rect 4773 26860 4807 26894
rect 4841 26860 4875 26894
rect 4909 26860 4943 26894
rect 4977 26860 5095 26894
rect 199 25925 317 25959
rect 351 25925 385 25959
rect 419 25925 453 25959
rect 487 25925 521 25959
rect 555 25925 589 25959
rect 623 25925 657 25959
rect 691 25925 725 25959
rect 759 25925 793 25959
rect 827 25925 861 25959
rect 895 25925 929 25959
rect 963 25925 997 25959
rect 1031 25925 1065 25959
rect 1099 25925 1133 25959
rect 1167 25925 1201 25959
rect 1235 25925 1269 25959
rect 1303 25925 1421 25959
rect 199 25849 233 25925
rect 1387 25849 1421 25925
rect 199 25781 233 25815
rect 199 25713 233 25747
rect 1387 25781 1421 25815
rect 199 25603 233 25679
rect 1387 25713 1421 25747
rect 1387 25603 1421 25679
rect 199 25569 317 25603
rect 351 25569 385 25603
rect 419 25569 453 25603
rect 487 25569 521 25603
rect 555 25569 589 25603
rect 623 25569 657 25603
rect 691 25569 725 25603
rect 759 25569 793 25603
rect 827 25569 861 25603
rect 895 25569 929 25603
rect 963 25569 997 25603
rect 1031 25569 1065 25603
rect 1099 25569 1133 25603
rect 1167 25569 1201 25603
rect 1235 25569 1269 25603
rect 1303 25569 1421 25603
rect 2352 25929 2470 25963
rect 2504 25929 2538 25963
rect 2572 25929 2606 25963
rect 2640 25929 2674 25963
rect 2708 25929 2742 25963
rect 2776 25929 2810 25963
rect 2844 25929 2878 25963
rect 2912 25929 2946 25963
rect 2980 25929 3014 25963
rect 3048 25929 3082 25963
rect 3116 25929 3150 25963
rect 3184 25929 3218 25963
rect 3252 25929 3286 25963
rect 3320 25929 3354 25963
rect 3388 25929 3422 25963
rect 3456 25929 3574 25963
rect 2352 25853 2386 25929
rect 3540 25853 3574 25929
rect 3873 25929 3991 25963
rect 4025 25929 4059 25963
rect 4093 25929 4127 25963
rect 4161 25929 4195 25963
rect 4229 25929 4263 25963
rect 4297 25929 4331 25963
rect 4365 25929 4399 25963
rect 4433 25929 4467 25963
rect 4501 25929 4535 25963
rect 4569 25929 4603 25963
rect 4637 25929 4671 25963
rect 4705 25929 4739 25963
rect 4773 25929 4807 25963
rect 4841 25929 4875 25963
rect 4909 25929 4943 25963
rect 4977 25929 5095 25963
rect 2352 25785 2386 25819
rect 2352 25717 2386 25751
rect 3540 25785 3574 25819
rect 3873 25853 3907 25929
rect 5061 25853 5095 25929
rect 3873 25785 3907 25819
rect 2352 25607 2386 25683
rect 3540 25717 3574 25751
rect 3540 25607 3574 25683
rect 2352 25573 2470 25607
rect 2504 25573 2538 25607
rect 2572 25573 2606 25607
rect 2640 25573 2674 25607
rect 2708 25573 2742 25607
rect 2776 25573 2810 25607
rect 2844 25573 2878 25607
rect 2912 25573 2946 25607
rect 2980 25573 3014 25607
rect 3048 25573 3082 25607
rect 3116 25573 3150 25607
rect 3184 25573 3218 25607
rect 3252 25573 3286 25607
rect 3320 25573 3354 25607
rect 3388 25573 3422 25607
rect 3456 25573 3574 25607
rect 3873 25717 3907 25751
rect 5061 25785 5095 25819
rect 3873 25607 3907 25683
rect 5061 25717 5095 25751
rect 5061 25607 5095 25683
rect 3873 25573 3991 25607
rect 4025 25573 4059 25607
rect 4093 25573 4127 25607
rect 4161 25573 4195 25607
rect 4229 25573 4263 25607
rect 4297 25573 4331 25607
rect 4365 25573 4399 25607
rect 4433 25573 4467 25607
rect 4501 25573 4535 25607
rect 4569 25573 4603 25607
rect 4637 25573 4671 25607
rect 4705 25573 4739 25607
rect 4773 25573 4807 25607
rect 4841 25573 4875 25607
rect 4909 25573 4943 25607
rect 4977 25573 5095 25607
rect 199 24638 317 24672
rect 351 24638 385 24672
rect 419 24638 453 24672
rect 487 24638 521 24672
rect 555 24638 589 24672
rect 623 24638 657 24672
rect 691 24638 725 24672
rect 759 24638 793 24672
rect 827 24638 861 24672
rect 895 24638 929 24672
rect 963 24638 997 24672
rect 1031 24638 1065 24672
rect 1099 24638 1133 24672
rect 1167 24638 1201 24672
rect 1235 24638 1269 24672
rect 1303 24638 1421 24672
rect 199 24562 233 24638
rect 1387 24562 1421 24638
rect 199 24494 233 24528
rect 199 24426 233 24460
rect 1387 24494 1421 24528
rect 199 24316 233 24392
rect 1387 24426 1421 24460
rect 1387 24316 1421 24392
rect 199 24282 317 24316
rect 351 24282 385 24316
rect 419 24282 453 24316
rect 487 24282 521 24316
rect 555 24282 589 24316
rect 623 24282 657 24316
rect 691 24282 725 24316
rect 759 24282 793 24316
rect 827 24282 861 24316
rect 895 24282 929 24316
rect 963 24282 997 24316
rect 1031 24282 1065 24316
rect 1099 24282 1133 24316
rect 1167 24282 1201 24316
rect 1235 24282 1269 24316
rect 1303 24282 1421 24316
rect 2352 24642 2470 24676
rect 2504 24642 2538 24676
rect 2572 24642 2606 24676
rect 2640 24642 2674 24676
rect 2708 24642 2742 24676
rect 2776 24642 2810 24676
rect 2844 24642 2878 24676
rect 2912 24642 2946 24676
rect 2980 24642 3014 24676
rect 3048 24642 3082 24676
rect 3116 24642 3150 24676
rect 3184 24642 3218 24676
rect 3252 24642 3286 24676
rect 3320 24642 3354 24676
rect 3388 24642 3422 24676
rect 3456 24642 3574 24676
rect 2352 24566 2386 24642
rect 3540 24566 3574 24642
rect 3873 24642 3991 24676
rect 4025 24642 4059 24676
rect 4093 24642 4127 24676
rect 4161 24642 4195 24676
rect 4229 24642 4263 24676
rect 4297 24642 4331 24676
rect 4365 24642 4399 24676
rect 4433 24642 4467 24676
rect 4501 24642 4535 24676
rect 4569 24642 4603 24676
rect 4637 24642 4671 24676
rect 4705 24642 4739 24676
rect 4773 24642 4807 24676
rect 4841 24642 4875 24676
rect 4909 24642 4943 24676
rect 4977 24642 5095 24676
rect 2352 24498 2386 24532
rect 2352 24430 2386 24464
rect 3540 24498 3574 24532
rect 3873 24566 3907 24642
rect 5061 24566 5095 24642
rect 3873 24498 3907 24532
rect 2352 24320 2386 24396
rect 3540 24430 3574 24464
rect 3540 24320 3574 24396
rect 2352 24286 2470 24320
rect 2504 24286 2538 24320
rect 2572 24286 2606 24320
rect 2640 24286 2674 24320
rect 2708 24286 2742 24320
rect 2776 24286 2810 24320
rect 2844 24286 2878 24320
rect 2912 24286 2946 24320
rect 2980 24286 3014 24320
rect 3048 24286 3082 24320
rect 3116 24286 3150 24320
rect 3184 24286 3218 24320
rect 3252 24286 3286 24320
rect 3320 24286 3354 24320
rect 3388 24286 3422 24320
rect 3456 24286 3574 24320
rect 3873 24430 3907 24464
rect 5061 24498 5095 24532
rect 3873 24320 3907 24396
rect 5061 24430 5095 24464
rect 5061 24320 5095 24396
rect 3873 24286 3991 24320
rect 4025 24286 4059 24320
rect 4093 24286 4127 24320
rect 4161 24286 4195 24320
rect 4229 24286 4263 24320
rect 4297 24286 4331 24320
rect 4365 24286 4399 24320
rect 4433 24286 4467 24320
rect 4501 24286 4535 24320
rect 4569 24286 4603 24320
rect 4637 24286 4671 24320
rect 4705 24286 4739 24320
rect 4773 24286 4807 24320
rect 4841 24286 4875 24320
rect 4909 24286 4943 24320
rect 4977 24286 5095 24320
rect 199 23351 317 23385
rect 351 23351 385 23385
rect 419 23351 453 23385
rect 487 23351 521 23385
rect 555 23351 589 23385
rect 623 23351 657 23385
rect 691 23351 725 23385
rect 759 23351 793 23385
rect 827 23351 861 23385
rect 895 23351 929 23385
rect 963 23351 997 23385
rect 1031 23351 1065 23385
rect 1099 23351 1133 23385
rect 1167 23351 1201 23385
rect 1235 23351 1269 23385
rect 1303 23351 1421 23385
rect 199 23275 233 23351
rect 1387 23275 1421 23351
rect 199 23207 233 23241
rect 199 23139 233 23173
rect 1387 23207 1421 23241
rect 199 23029 233 23105
rect 1387 23139 1421 23173
rect 1387 23029 1421 23105
rect 199 22995 317 23029
rect 351 22995 385 23029
rect 419 22995 453 23029
rect 487 22995 521 23029
rect 555 22995 589 23029
rect 623 22995 657 23029
rect 691 22995 725 23029
rect 759 22995 793 23029
rect 827 22995 861 23029
rect 895 22995 929 23029
rect 963 22995 997 23029
rect 1031 22995 1065 23029
rect 1099 22995 1133 23029
rect 1167 22995 1201 23029
rect 1235 22995 1269 23029
rect 1303 22995 1421 23029
rect 2352 23355 2470 23389
rect 2504 23355 2538 23389
rect 2572 23355 2606 23389
rect 2640 23355 2674 23389
rect 2708 23355 2742 23389
rect 2776 23355 2810 23389
rect 2844 23355 2878 23389
rect 2912 23355 2946 23389
rect 2980 23355 3014 23389
rect 3048 23355 3082 23389
rect 3116 23355 3150 23389
rect 3184 23355 3218 23389
rect 3252 23355 3286 23389
rect 3320 23355 3354 23389
rect 3388 23355 3422 23389
rect 3456 23355 3574 23389
rect 2352 23279 2386 23355
rect 3540 23279 3574 23355
rect 3873 23355 3991 23389
rect 4025 23355 4059 23389
rect 4093 23355 4127 23389
rect 4161 23355 4195 23389
rect 4229 23355 4263 23389
rect 4297 23355 4331 23389
rect 4365 23355 4399 23389
rect 4433 23355 4467 23389
rect 4501 23355 4535 23389
rect 4569 23355 4603 23389
rect 4637 23355 4671 23389
rect 4705 23355 4739 23389
rect 4773 23355 4807 23389
rect 4841 23355 4875 23389
rect 4909 23355 4943 23389
rect 4977 23355 5095 23389
rect 2352 23211 2386 23245
rect 2352 23143 2386 23177
rect 3540 23211 3574 23245
rect 3873 23279 3907 23355
rect 5061 23279 5095 23355
rect 3873 23211 3907 23245
rect 2352 23033 2386 23109
rect 3540 23143 3574 23177
rect 3540 23033 3574 23109
rect 2352 22999 2470 23033
rect 2504 22999 2538 23033
rect 2572 22999 2606 23033
rect 2640 22999 2674 23033
rect 2708 22999 2742 23033
rect 2776 22999 2810 23033
rect 2844 22999 2878 23033
rect 2912 22999 2946 23033
rect 2980 22999 3014 23033
rect 3048 22999 3082 23033
rect 3116 22999 3150 23033
rect 3184 22999 3218 23033
rect 3252 22999 3286 23033
rect 3320 22999 3354 23033
rect 3388 22999 3422 23033
rect 3456 22999 3574 23033
rect 3873 23143 3907 23177
rect 5061 23211 5095 23245
rect 3873 23033 3907 23109
rect 5061 23143 5095 23177
rect 5061 23033 5095 23109
rect 3873 22999 3991 23033
rect 4025 22999 4059 23033
rect 4093 22999 4127 23033
rect 4161 22999 4195 23033
rect 4229 22999 4263 23033
rect 4297 22999 4331 23033
rect 4365 22999 4399 23033
rect 4433 22999 4467 23033
rect 4501 22999 4535 23033
rect 4569 22999 4603 23033
rect 4637 22999 4671 23033
rect 4705 22999 4739 23033
rect 4773 22999 4807 23033
rect 4841 22999 4875 23033
rect 4909 22999 4943 23033
rect 4977 22999 5095 23033
rect 199 22064 317 22098
rect 351 22064 385 22098
rect 419 22064 453 22098
rect 487 22064 521 22098
rect 555 22064 589 22098
rect 623 22064 657 22098
rect 691 22064 725 22098
rect 759 22064 793 22098
rect 827 22064 861 22098
rect 895 22064 929 22098
rect 963 22064 997 22098
rect 1031 22064 1065 22098
rect 1099 22064 1133 22098
rect 1167 22064 1201 22098
rect 1235 22064 1269 22098
rect 1303 22064 1421 22098
rect 199 21988 233 22064
rect 1387 21988 1421 22064
rect 199 21920 233 21954
rect 199 21852 233 21886
rect 1387 21920 1421 21954
rect 199 21742 233 21818
rect 1387 21852 1421 21886
rect 1387 21742 1421 21818
rect 199 21708 317 21742
rect 351 21708 385 21742
rect 419 21708 453 21742
rect 487 21708 521 21742
rect 555 21708 589 21742
rect 623 21708 657 21742
rect 691 21708 725 21742
rect 759 21708 793 21742
rect 827 21708 861 21742
rect 895 21708 929 21742
rect 963 21708 997 21742
rect 1031 21708 1065 21742
rect 1099 21708 1133 21742
rect 1167 21708 1201 21742
rect 1235 21708 1269 21742
rect 1303 21708 1421 21742
rect 2352 22068 2470 22102
rect 2504 22068 2538 22102
rect 2572 22068 2606 22102
rect 2640 22068 2674 22102
rect 2708 22068 2742 22102
rect 2776 22068 2810 22102
rect 2844 22068 2878 22102
rect 2912 22068 2946 22102
rect 2980 22068 3014 22102
rect 3048 22068 3082 22102
rect 3116 22068 3150 22102
rect 3184 22068 3218 22102
rect 3252 22068 3286 22102
rect 3320 22068 3354 22102
rect 3388 22068 3422 22102
rect 3456 22068 3574 22102
rect 2352 21992 2386 22068
rect 3540 21992 3574 22068
rect 3873 22068 3991 22102
rect 4025 22068 4059 22102
rect 4093 22068 4127 22102
rect 4161 22068 4195 22102
rect 4229 22068 4263 22102
rect 4297 22068 4331 22102
rect 4365 22068 4399 22102
rect 4433 22068 4467 22102
rect 4501 22068 4535 22102
rect 4569 22068 4603 22102
rect 4637 22068 4671 22102
rect 4705 22068 4739 22102
rect 4773 22068 4807 22102
rect 4841 22068 4875 22102
rect 4909 22068 4943 22102
rect 4977 22068 5095 22102
rect 2352 21924 2386 21958
rect 2352 21856 2386 21890
rect 3540 21924 3574 21958
rect 3873 21992 3907 22068
rect 5061 21992 5095 22068
rect 3873 21924 3907 21958
rect 2352 21746 2386 21822
rect 3540 21856 3574 21890
rect 3540 21746 3574 21822
rect 2352 21712 2470 21746
rect 2504 21712 2538 21746
rect 2572 21712 2606 21746
rect 2640 21712 2674 21746
rect 2708 21712 2742 21746
rect 2776 21712 2810 21746
rect 2844 21712 2878 21746
rect 2912 21712 2946 21746
rect 2980 21712 3014 21746
rect 3048 21712 3082 21746
rect 3116 21712 3150 21746
rect 3184 21712 3218 21746
rect 3252 21712 3286 21746
rect 3320 21712 3354 21746
rect 3388 21712 3422 21746
rect 3456 21712 3574 21746
rect 3873 21856 3907 21890
rect 5061 21924 5095 21958
rect 3873 21746 3907 21822
rect 5061 21856 5095 21890
rect 5061 21746 5095 21822
rect 3873 21712 3991 21746
rect 4025 21712 4059 21746
rect 4093 21712 4127 21746
rect 4161 21712 4195 21746
rect 4229 21712 4263 21746
rect 4297 21712 4331 21746
rect 4365 21712 4399 21746
rect 4433 21712 4467 21746
rect 4501 21712 4535 21746
rect 4569 21712 4603 21746
rect 4637 21712 4671 21746
rect 4705 21712 4739 21746
rect 4773 21712 4807 21746
rect 4841 21712 4875 21746
rect 4909 21712 4943 21746
rect 4977 21712 5095 21746
rect 199 20777 317 20811
rect 351 20777 385 20811
rect 419 20777 453 20811
rect 487 20777 521 20811
rect 555 20777 589 20811
rect 623 20777 657 20811
rect 691 20777 725 20811
rect 759 20777 793 20811
rect 827 20777 861 20811
rect 895 20777 929 20811
rect 963 20777 997 20811
rect 1031 20777 1065 20811
rect 1099 20777 1133 20811
rect 1167 20777 1201 20811
rect 1235 20777 1269 20811
rect 1303 20777 1421 20811
rect 199 20701 233 20777
rect 1387 20701 1421 20777
rect 199 20633 233 20667
rect 199 20565 233 20599
rect 1387 20633 1421 20667
rect 199 20455 233 20531
rect 1387 20565 1421 20599
rect 1387 20455 1421 20531
rect 199 20421 317 20455
rect 351 20421 385 20455
rect 419 20421 453 20455
rect 487 20421 521 20455
rect 555 20421 589 20455
rect 623 20421 657 20455
rect 691 20421 725 20455
rect 759 20421 793 20455
rect 827 20421 861 20455
rect 895 20421 929 20455
rect 963 20421 997 20455
rect 1031 20421 1065 20455
rect 1099 20421 1133 20455
rect 1167 20421 1201 20455
rect 1235 20421 1269 20455
rect 1303 20421 1421 20455
rect 2352 20781 2470 20815
rect 2504 20781 2538 20815
rect 2572 20781 2606 20815
rect 2640 20781 2674 20815
rect 2708 20781 2742 20815
rect 2776 20781 2810 20815
rect 2844 20781 2878 20815
rect 2912 20781 2946 20815
rect 2980 20781 3014 20815
rect 3048 20781 3082 20815
rect 3116 20781 3150 20815
rect 3184 20781 3218 20815
rect 3252 20781 3286 20815
rect 3320 20781 3354 20815
rect 3388 20781 3422 20815
rect 3456 20781 3574 20815
rect 2352 20705 2386 20781
rect 3540 20705 3574 20781
rect 3873 20781 3991 20815
rect 4025 20781 4059 20815
rect 4093 20781 4127 20815
rect 4161 20781 4195 20815
rect 4229 20781 4263 20815
rect 4297 20781 4331 20815
rect 4365 20781 4399 20815
rect 4433 20781 4467 20815
rect 4501 20781 4535 20815
rect 4569 20781 4603 20815
rect 4637 20781 4671 20815
rect 4705 20781 4739 20815
rect 4773 20781 4807 20815
rect 4841 20781 4875 20815
rect 4909 20781 4943 20815
rect 4977 20781 5095 20815
rect 2352 20637 2386 20671
rect 2352 20569 2386 20603
rect 3540 20637 3574 20671
rect 3873 20705 3907 20781
rect 5061 20705 5095 20781
rect 3873 20637 3907 20671
rect 2352 20459 2386 20535
rect 3540 20569 3574 20603
rect 3540 20459 3574 20535
rect 2352 20425 2470 20459
rect 2504 20425 2538 20459
rect 2572 20425 2606 20459
rect 2640 20425 2674 20459
rect 2708 20425 2742 20459
rect 2776 20425 2810 20459
rect 2844 20425 2878 20459
rect 2912 20425 2946 20459
rect 2980 20425 3014 20459
rect 3048 20425 3082 20459
rect 3116 20425 3150 20459
rect 3184 20425 3218 20459
rect 3252 20425 3286 20459
rect 3320 20425 3354 20459
rect 3388 20425 3422 20459
rect 3456 20425 3574 20459
rect 3873 20569 3907 20603
rect 5061 20637 5095 20671
rect 3873 20459 3907 20535
rect 5061 20569 5095 20603
rect 5061 20459 5095 20535
rect 3873 20425 3991 20459
rect 4025 20425 4059 20459
rect 4093 20425 4127 20459
rect 4161 20425 4195 20459
rect 4229 20425 4263 20459
rect 4297 20425 4331 20459
rect 4365 20425 4399 20459
rect 4433 20425 4467 20459
rect 4501 20425 4535 20459
rect 4569 20425 4603 20459
rect 4637 20425 4671 20459
rect 4705 20425 4739 20459
rect 4773 20425 4807 20459
rect 4841 20425 4875 20459
rect 4909 20425 4943 20459
rect 4977 20425 5095 20459
rect 199 19490 317 19524
rect 351 19490 385 19524
rect 419 19490 453 19524
rect 487 19490 521 19524
rect 555 19490 589 19524
rect 623 19490 657 19524
rect 691 19490 725 19524
rect 759 19490 793 19524
rect 827 19490 861 19524
rect 895 19490 929 19524
rect 963 19490 997 19524
rect 1031 19490 1065 19524
rect 1099 19490 1133 19524
rect 1167 19490 1201 19524
rect 1235 19490 1269 19524
rect 1303 19490 1421 19524
rect 199 19414 233 19490
rect 1387 19414 1421 19490
rect 199 19346 233 19380
rect 199 19278 233 19312
rect 1387 19346 1421 19380
rect 199 19168 233 19244
rect 1387 19278 1421 19312
rect 1387 19168 1421 19244
rect 199 19134 317 19168
rect 351 19134 385 19168
rect 419 19134 453 19168
rect 487 19134 521 19168
rect 555 19134 589 19168
rect 623 19134 657 19168
rect 691 19134 725 19168
rect 759 19134 793 19168
rect 827 19134 861 19168
rect 895 19134 929 19168
rect 963 19134 997 19168
rect 1031 19134 1065 19168
rect 1099 19134 1133 19168
rect 1167 19134 1201 19168
rect 1235 19134 1269 19168
rect 1303 19134 1421 19168
rect 2352 19494 2470 19528
rect 2504 19494 2538 19528
rect 2572 19494 2606 19528
rect 2640 19494 2674 19528
rect 2708 19494 2742 19528
rect 2776 19494 2810 19528
rect 2844 19494 2878 19528
rect 2912 19494 2946 19528
rect 2980 19494 3014 19528
rect 3048 19494 3082 19528
rect 3116 19494 3150 19528
rect 3184 19494 3218 19528
rect 3252 19494 3286 19528
rect 3320 19494 3354 19528
rect 3388 19494 3422 19528
rect 3456 19494 3574 19528
rect 2352 19418 2386 19494
rect 3540 19418 3574 19494
rect 3873 19494 3991 19528
rect 4025 19494 4059 19528
rect 4093 19494 4127 19528
rect 4161 19494 4195 19528
rect 4229 19494 4263 19528
rect 4297 19494 4331 19528
rect 4365 19494 4399 19528
rect 4433 19494 4467 19528
rect 4501 19494 4535 19528
rect 4569 19494 4603 19528
rect 4637 19494 4671 19528
rect 4705 19494 4739 19528
rect 4773 19494 4807 19528
rect 4841 19494 4875 19528
rect 4909 19494 4943 19528
rect 4977 19494 5095 19528
rect 2352 19350 2386 19384
rect 2352 19282 2386 19316
rect 3540 19350 3574 19384
rect 3873 19418 3907 19494
rect 5061 19418 5095 19494
rect 3873 19350 3907 19384
rect 2352 19172 2386 19248
rect 3540 19282 3574 19316
rect 3540 19172 3574 19248
rect 2352 19138 2470 19172
rect 2504 19138 2538 19172
rect 2572 19138 2606 19172
rect 2640 19138 2674 19172
rect 2708 19138 2742 19172
rect 2776 19138 2810 19172
rect 2844 19138 2878 19172
rect 2912 19138 2946 19172
rect 2980 19138 3014 19172
rect 3048 19138 3082 19172
rect 3116 19138 3150 19172
rect 3184 19138 3218 19172
rect 3252 19138 3286 19172
rect 3320 19138 3354 19172
rect 3388 19138 3422 19172
rect 3456 19138 3574 19172
rect 3873 19282 3907 19316
rect 5061 19350 5095 19384
rect 3873 19172 3907 19248
rect 5061 19282 5095 19316
rect 5061 19172 5095 19248
rect 3873 19138 3991 19172
rect 4025 19138 4059 19172
rect 4093 19138 4127 19172
rect 4161 19138 4195 19172
rect 4229 19138 4263 19172
rect 4297 19138 4331 19172
rect 4365 19138 4399 19172
rect 4433 19138 4467 19172
rect 4501 19138 4535 19172
rect 4569 19138 4603 19172
rect 4637 19138 4671 19172
rect 4705 19138 4739 19172
rect 4773 19138 4807 19172
rect 4841 19138 4875 19172
rect 4909 19138 4943 19172
rect 4977 19138 5095 19172
rect 199 18203 317 18237
rect 351 18203 385 18237
rect 419 18203 453 18237
rect 487 18203 521 18237
rect 555 18203 589 18237
rect 623 18203 657 18237
rect 691 18203 725 18237
rect 759 18203 793 18237
rect 827 18203 861 18237
rect 895 18203 929 18237
rect 963 18203 997 18237
rect 1031 18203 1065 18237
rect 1099 18203 1133 18237
rect 1167 18203 1201 18237
rect 1235 18203 1269 18237
rect 1303 18203 1421 18237
rect 199 18127 233 18203
rect 1387 18127 1421 18203
rect 199 18059 233 18093
rect 199 17991 233 18025
rect 1387 18059 1421 18093
rect 199 17881 233 17957
rect 1387 17991 1421 18025
rect 1387 17881 1421 17957
rect 199 17847 317 17881
rect 351 17847 385 17881
rect 419 17847 453 17881
rect 487 17847 521 17881
rect 555 17847 589 17881
rect 623 17847 657 17881
rect 691 17847 725 17881
rect 759 17847 793 17881
rect 827 17847 861 17881
rect 895 17847 929 17881
rect 963 17847 997 17881
rect 1031 17847 1065 17881
rect 1099 17847 1133 17881
rect 1167 17847 1201 17881
rect 1235 17847 1269 17881
rect 1303 17847 1421 17881
rect 2352 18207 2470 18241
rect 2504 18207 2538 18241
rect 2572 18207 2606 18241
rect 2640 18207 2674 18241
rect 2708 18207 2742 18241
rect 2776 18207 2810 18241
rect 2844 18207 2878 18241
rect 2912 18207 2946 18241
rect 2980 18207 3014 18241
rect 3048 18207 3082 18241
rect 3116 18207 3150 18241
rect 3184 18207 3218 18241
rect 3252 18207 3286 18241
rect 3320 18207 3354 18241
rect 3388 18207 3422 18241
rect 3456 18207 3574 18241
rect 2352 18131 2386 18207
rect 3540 18131 3574 18207
rect 3873 18207 3991 18241
rect 4025 18207 4059 18241
rect 4093 18207 4127 18241
rect 4161 18207 4195 18241
rect 4229 18207 4263 18241
rect 4297 18207 4331 18241
rect 4365 18207 4399 18241
rect 4433 18207 4467 18241
rect 4501 18207 4535 18241
rect 4569 18207 4603 18241
rect 4637 18207 4671 18241
rect 4705 18207 4739 18241
rect 4773 18207 4807 18241
rect 4841 18207 4875 18241
rect 4909 18207 4943 18241
rect 4977 18207 5095 18241
rect 2352 18063 2386 18097
rect 2352 17995 2386 18029
rect 3540 18063 3574 18097
rect 3873 18131 3907 18207
rect 5061 18131 5095 18207
rect 3873 18063 3907 18097
rect 2352 17885 2386 17961
rect 3540 17995 3574 18029
rect 3540 17885 3574 17961
rect 2352 17851 2470 17885
rect 2504 17851 2538 17885
rect 2572 17851 2606 17885
rect 2640 17851 2674 17885
rect 2708 17851 2742 17885
rect 2776 17851 2810 17885
rect 2844 17851 2878 17885
rect 2912 17851 2946 17885
rect 2980 17851 3014 17885
rect 3048 17851 3082 17885
rect 3116 17851 3150 17885
rect 3184 17851 3218 17885
rect 3252 17851 3286 17885
rect 3320 17851 3354 17885
rect 3388 17851 3422 17885
rect 3456 17851 3574 17885
rect 3873 17995 3907 18029
rect 5061 18063 5095 18097
rect 3873 17885 3907 17961
rect 5061 17995 5095 18029
rect 5061 17885 5095 17961
rect 3873 17851 3991 17885
rect 4025 17851 4059 17885
rect 4093 17851 4127 17885
rect 4161 17851 4195 17885
rect 4229 17851 4263 17885
rect 4297 17851 4331 17885
rect 4365 17851 4399 17885
rect 4433 17851 4467 17885
rect 4501 17851 4535 17885
rect 4569 17851 4603 17885
rect 4637 17851 4671 17885
rect 4705 17851 4739 17885
rect 4773 17851 4807 17885
rect 4841 17851 4875 17885
rect 4909 17851 4943 17885
rect 4977 17851 5095 17885
rect 199 16916 317 16950
rect 351 16916 385 16950
rect 419 16916 453 16950
rect 487 16916 521 16950
rect 555 16916 589 16950
rect 623 16916 657 16950
rect 691 16916 725 16950
rect 759 16916 793 16950
rect 827 16916 861 16950
rect 895 16916 929 16950
rect 963 16916 997 16950
rect 1031 16916 1065 16950
rect 1099 16916 1133 16950
rect 1167 16916 1201 16950
rect 1235 16916 1269 16950
rect 1303 16916 1421 16950
rect 199 16840 233 16916
rect 1387 16840 1421 16916
rect 199 16772 233 16806
rect 199 16704 233 16738
rect 1387 16772 1421 16806
rect 199 16594 233 16670
rect 1387 16704 1421 16738
rect 1387 16594 1421 16670
rect 199 16560 317 16594
rect 351 16560 385 16594
rect 419 16560 453 16594
rect 487 16560 521 16594
rect 555 16560 589 16594
rect 623 16560 657 16594
rect 691 16560 725 16594
rect 759 16560 793 16594
rect 827 16560 861 16594
rect 895 16560 929 16594
rect 963 16560 997 16594
rect 1031 16560 1065 16594
rect 1099 16560 1133 16594
rect 1167 16560 1201 16594
rect 1235 16560 1269 16594
rect 1303 16560 1421 16594
rect 2352 16920 2470 16954
rect 2504 16920 2538 16954
rect 2572 16920 2606 16954
rect 2640 16920 2674 16954
rect 2708 16920 2742 16954
rect 2776 16920 2810 16954
rect 2844 16920 2878 16954
rect 2912 16920 2946 16954
rect 2980 16920 3014 16954
rect 3048 16920 3082 16954
rect 3116 16920 3150 16954
rect 3184 16920 3218 16954
rect 3252 16920 3286 16954
rect 3320 16920 3354 16954
rect 3388 16920 3422 16954
rect 3456 16920 3574 16954
rect 2352 16844 2386 16920
rect 3540 16844 3574 16920
rect 3873 16920 3991 16954
rect 4025 16920 4059 16954
rect 4093 16920 4127 16954
rect 4161 16920 4195 16954
rect 4229 16920 4263 16954
rect 4297 16920 4331 16954
rect 4365 16920 4399 16954
rect 4433 16920 4467 16954
rect 4501 16920 4535 16954
rect 4569 16920 4603 16954
rect 4637 16920 4671 16954
rect 4705 16920 4739 16954
rect 4773 16920 4807 16954
rect 4841 16920 4875 16954
rect 4909 16920 4943 16954
rect 4977 16920 5095 16954
rect 2352 16776 2386 16810
rect 2352 16708 2386 16742
rect 3540 16776 3574 16810
rect 3873 16844 3907 16920
rect 5061 16844 5095 16920
rect 3873 16776 3907 16810
rect 2352 16598 2386 16674
rect 3540 16708 3574 16742
rect 3540 16598 3574 16674
rect 2352 16564 2470 16598
rect 2504 16564 2538 16598
rect 2572 16564 2606 16598
rect 2640 16564 2674 16598
rect 2708 16564 2742 16598
rect 2776 16564 2810 16598
rect 2844 16564 2878 16598
rect 2912 16564 2946 16598
rect 2980 16564 3014 16598
rect 3048 16564 3082 16598
rect 3116 16564 3150 16598
rect 3184 16564 3218 16598
rect 3252 16564 3286 16598
rect 3320 16564 3354 16598
rect 3388 16564 3422 16598
rect 3456 16564 3574 16598
rect 3873 16708 3907 16742
rect 5061 16776 5095 16810
rect 3873 16598 3907 16674
rect 5061 16708 5095 16742
rect 5061 16598 5095 16674
rect 3873 16564 3991 16598
rect 4025 16564 4059 16598
rect 4093 16564 4127 16598
rect 4161 16564 4195 16598
rect 4229 16564 4263 16598
rect 4297 16564 4331 16598
rect 4365 16564 4399 16598
rect 4433 16564 4467 16598
rect 4501 16564 4535 16598
rect 4569 16564 4603 16598
rect 4637 16564 4671 16598
rect 4705 16564 4739 16598
rect 4773 16564 4807 16598
rect 4841 16564 4875 16598
rect 4909 16564 4943 16598
rect 4977 16564 5095 16598
rect 199 15629 317 15663
rect 351 15629 385 15663
rect 419 15629 453 15663
rect 487 15629 521 15663
rect 555 15629 589 15663
rect 623 15629 657 15663
rect 691 15629 725 15663
rect 759 15629 793 15663
rect 827 15629 861 15663
rect 895 15629 929 15663
rect 963 15629 997 15663
rect 1031 15629 1065 15663
rect 1099 15629 1133 15663
rect 1167 15629 1201 15663
rect 1235 15629 1269 15663
rect 1303 15629 1421 15663
rect 199 15553 233 15629
rect 1387 15553 1421 15629
rect 199 15485 233 15519
rect 199 15417 233 15451
rect 1387 15485 1421 15519
rect 199 15307 233 15383
rect 1387 15417 1421 15451
rect 1387 15307 1421 15383
rect 199 15273 317 15307
rect 351 15273 385 15307
rect 419 15273 453 15307
rect 487 15273 521 15307
rect 555 15273 589 15307
rect 623 15273 657 15307
rect 691 15273 725 15307
rect 759 15273 793 15307
rect 827 15273 861 15307
rect 895 15273 929 15307
rect 963 15273 997 15307
rect 1031 15273 1065 15307
rect 1099 15273 1133 15307
rect 1167 15273 1201 15307
rect 1235 15273 1269 15307
rect 1303 15273 1421 15307
rect 2352 15633 2470 15667
rect 2504 15633 2538 15667
rect 2572 15633 2606 15667
rect 2640 15633 2674 15667
rect 2708 15633 2742 15667
rect 2776 15633 2810 15667
rect 2844 15633 2878 15667
rect 2912 15633 2946 15667
rect 2980 15633 3014 15667
rect 3048 15633 3082 15667
rect 3116 15633 3150 15667
rect 3184 15633 3218 15667
rect 3252 15633 3286 15667
rect 3320 15633 3354 15667
rect 3388 15633 3422 15667
rect 3456 15633 3574 15667
rect 2352 15557 2386 15633
rect 3540 15557 3574 15633
rect 3873 15633 3991 15667
rect 4025 15633 4059 15667
rect 4093 15633 4127 15667
rect 4161 15633 4195 15667
rect 4229 15633 4263 15667
rect 4297 15633 4331 15667
rect 4365 15633 4399 15667
rect 4433 15633 4467 15667
rect 4501 15633 4535 15667
rect 4569 15633 4603 15667
rect 4637 15633 4671 15667
rect 4705 15633 4739 15667
rect 4773 15633 4807 15667
rect 4841 15633 4875 15667
rect 4909 15633 4943 15667
rect 4977 15633 5095 15667
rect 2352 15489 2386 15523
rect 2352 15421 2386 15455
rect 3540 15489 3574 15523
rect 3873 15557 3907 15633
rect 5061 15557 5095 15633
rect 3873 15489 3907 15523
rect 2352 15311 2386 15387
rect 3540 15421 3574 15455
rect 3540 15311 3574 15387
rect 2352 15277 2470 15311
rect 2504 15277 2538 15311
rect 2572 15277 2606 15311
rect 2640 15277 2674 15311
rect 2708 15277 2742 15311
rect 2776 15277 2810 15311
rect 2844 15277 2878 15311
rect 2912 15277 2946 15311
rect 2980 15277 3014 15311
rect 3048 15277 3082 15311
rect 3116 15277 3150 15311
rect 3184 15277 3218 15311
rect 3252 15277 3286 15311
rect 3320 15277 3354 15311
rect 3388 15277 3422 15311
rect 3456 15277 3574 15311
rect 3873 15421 3907 15455
rect 5061 15489 5095 15523
rect 3873 15311 3907 15387
rect 5061 15421 5095 15455
rect 5061 15311 5095 15387
rect 3873 15277 3991 15311
rect 4025 15277 4059 15311
rect 4093 15277 4127 15311
rect 4161 15277 4195 15311
rect 4229 15277 4263 15311
rect 4297 15277 4331 15311
rect 4365 15277 4399 15311
rect 4433 15277 4467 15311
rect 4501 15277 4535 15311
rect 4569 15277 4603 15311
rect 4637 15277 4671 15311
rect 4705 15277 4739 15311
rect 4773 15277 4807 15311
rect 4841 15277 4875 15311
rect 4909 15277 4943 15311
rect 4977 15277 5095 15311
rect 199 14342 317 14376
rect 351 14342 385 14376
rect 419 14342 453 14376
rect 487 14342 521 14376
rect 555 14342 589 14376
rect 623 14342 657 14376
rect 691 14342 725 14376
rect 759 14342 793 14376
rect 827 14342 861 14376
rect 895 14342 929 14376
rect 963 14342 997 14376
rect 1031 14342 1065 14376
rect 1099 14342 1133 14376
rect 1167 14342 1201 14376
rect 1235 14342 1269 14376
rect 1303 14342 1421 14376
rect 199 14266 233 14342
rect 1387 14266 1421 14342
rect 199 14198 233 14232
rect 199 14130 233 14164
rect 1387 14198 1421 14232
rect 199 14020 233 14096
rect 1387 14130 1421 14164
rect 1387 14020 1421 14096
rect 199 13986 317 14020
rect 351 13986 385 14020
rect 419 13986 453 14020
rect 487 13986 521 14020
rect 555 13986 589 14020
rect 623 13986 657 14020
rect 691 13986 725 14020
rect 759 13986 793 14020
rect 827 13986 861 14020
rect 895 13986 929 14020
rect 963 13986 997 14020
rect 1031 13986 1065 14020
rect 1099 13986 1133 14020
rect 1167 13986 1201 14020
rect 1235 13986 1269 14020
rect 1303 13986 1421 14020
rect 2352 14346 2470 14380
rect 2504 14346 2538 14380
rect 2572 14346 2606 14380
rect 2640 14346 2674 14380
rect 2708 14346 2742 14380
rect 2776 14346 2810 14380
rect 2844 14346 2878 14380
rect 2912 14346 2946 14380
rect 2980 14346 3014 14380
rect 3048 14346 3082 14380
rect 3116 14346 3150 14380
rect 3184 14346 3218 14380
rect 3252 14346 3286 14380
rect 3320 14346 3354 14380
rect 3388 14346 3422 14380
rect 3456 14346 3574 14380
rect 2352 14270 2386 14346
rect 3540 14270 3574 14346
rect 3873 14346 3991 14380
rect 4025 14346 4059 14380
rect 4093 14346 4127 14380
rect 4161 14346 4195 14380
rect 4229 14346 4263 14380
rect 4297 14346 4331 14380
rect 4365 14346 4399 14380
rect 4433 14346 4467 14380
rect 4501 14346 4535 14380
rect 4569 14346 4603 14380
rect 4637 14346 4671 14380
rect 4705 14346 4739 14380
rect 4773 14346 4807 14380
rect 4841 14346 4875 14380
rect 4909 14346 4943 14380
rect 4977 14346 5095 14380
rect 2352 14202 2386 14236
rect 2352 14134 2386 14168
rect 3540 14202 3574 14236
rect 3873 14270 3907 14346
rect 5061 14270 5095 14346
rect 3873 14202 3907 14236
rect 2352 14024 2386 14100
rect 3540 14134 3574 14168
rect 3540 14024 3574 14100
rect 2352 13990 2470 14024
rect 2504 13990 2538 14024
rect 2572 13990 2606 14024
rect 2640 13990 2674 14024
rect 2708 13990 2742 14024
rect 2776 13990 2810 14024
rect 2844 13990 2878 14024
rect 2912 13990 2946 14024
rect 2980 13990 3014 14024
rect 3048 13990 3082 14024
rect 3116 13990 3150 14024
rect 3184 13990 3218 14024
rect 3252 13990 3286 14024
rect 3320 13990 3354 14024
rect 3388 13990 3422 14024
rect 3456 13990 3574 14024
rect 3873 14134 3907 14168
rect 5061 14202 5095 14236
rect 3873 14024 3907 14100
rect 5061 14134 5095 14168
rect 5061 14024 5095 14100
rect 3873 13990 3991 14024
rect 4025 13990 4059 14024
rect 4093 13990 4127 14024
rect 4161 13990 4195 14024
rect 4229 13990 4263 14024
rect 4297 13990 4331 14024
rect 4365 13990 4399 14024
rect 4433 13990 4467 14024
rect 4501 13990 4535 14024
rect 4569 13990 4603 14024
rect 4637 13990 4671 14024
rect 4705 13990 4739 14024
rect 4773 13990 4807 14024
rect 4841 13990 4875 14024
rect 4909 13990 4943 14024
rect 4977 13990 5095 14024
rect 199 13055 317 13089
rect 351 13055 385 13089
rect 419 13055 453 13089
rect 487 13055 521 13089
rect 555 13055 589 13089
rect 623 13055 657 13089
rect 691 13055 725 13089
rect 759 13055 793 13089
rect 827 13055 861 13089
rect 895 13055 929 13089
rect 963 13055 997 13089
rect 1031 13055 1065 13089
rect 1099 13055 1133 13089
rect 1167 13055 1201 13089
rect 1235 13055 1269 13089
rect 1303 13055 1421 13089
rect 199 12979 233 13055
rect 1387 12979 1421 13055
rect 199 12911 233 12945
rect 199 12843 233 12877
rect 1387 12911 1421 12945
rect 199 12733 233 12809
rect 1387 12843 1421 12877
rect 1387 12733 1421 12809
rect 199 12699 317 12733
rect 351 12699 385 12733
rect 419 12699 453 12733
rect 487 12699 521 12733
rect 555 12699 589 12733
rect 623 12699 657 12733
rect 691 12699 725 12733
rect 759 12699 793 12733
rect 827 12699 861 12733
rect 895 12699 929 12733
rect 963 12699 997 12733
rect 1031 12699 1065 12733
rect 1099 12699 1133 12733
rect 1167 12699 1201 12733
rect 1235 12699 1269 12733
rect 1303 12699 1421 12733
rect 2352 13059 2470 13093
rect 2504 13059 2538 13093
rect 2572 13059 2606 13093
rect 2640 13059 2674 13093
rect 2708 13059 2742 13093
rect 2776 13059 2810 13093
rect 2844 13059 2878 13093
rect 2912 13059 2946 13093
rect 2980 13059 3014 13093
rect 3048 13059 3082 13093
rect 3116 13059 3150 13093
rect 3184 13059 3218 13093
rect 3252 13059 3286 13093
rect 3320 13059 3354 13093
rect 3388 13059 3422 13093
rect 3456 13059 3574 13093
rect 2352 12983 2386 13059
rect 3540 12983 3574 13059
rect 3873 13059 3991 13093
rect 4025 13059 4059 13093
rect 4093 13059 4127 13093
rect 4161 13059 4195 13093
rect 4229 13059 4263 13093
rect 4297 13059 4331 13093
rect 4365 13059 4399 13093
rect 4433 13059 4467 13093
rect 4501 13059 4535 13093
rect 4569 13059 4603 13093
rect 4637 13059 4671 13093
rect 4705 13059 4739 13093
rect 4773 13059 4807 13093
rect 4841 13059 4875 13093
rect 4909 13059 4943 13093
rect 4977 13059 5095 13093
rect 2352 12915 2386 12949
rect 2352 12847 2386 12881
rect 3540 12915 3574 12949
rect 3873 12983 3907 13059
rect 5061 12983 5095 13059
rect 3873 12915 3907 12949
rect 2352 12737 2386 12813
rect 3540 12847 3574 12881
rect 3540 12737 3574 12813
rect 2352 12703 2470 12737
rect 2504 12703 2538 12737
rect 2572 12703 2606 12737
rect 2640 12703 2674 12737
rect 2708 12703 2742 12737
rect 2776 12703 2810 12737
rect 2844 12703 2878 12737
rect 2912 12703 2946 12737
rect 2980 12703 3014 12737
rect 3048 12703 3082 12737
rect 3116 12703 3150 12737
rect 3184 12703 3218 12737
rect 3252 12703 3286 12737
rect 3320 12703 3354 12737
rect 3388 12703 3422 12737
rect 3456 12703 3574 12737
rect 3873 12847 3907 12881
rect 5061 12915 5095 12949
rect 3873 12737 3907 12813
rect 5061 12847 5095 12881
rect 5061 12737 5095 12813
rect 3873 12703 3991 12737
rect 4025 12703 4059 12737
rect 4093 12703 4127 12737
rect 4161 12703 4195 12737
rect 4229 12703 4263 12737
rect 4297 12703 4331 12737
rect 4365 12703 4399 12737
rect 4433 12703 4467 12737
rect 4501 12703 4535 12737
rect 4569 12703 4603 12737
rect 4637 12703 4671 12737
rect 4705 12703 4739 12737
rect 4773 12703 4807 12737
rect 4841 12703 4875 12737
rect 4909 12703 4943 12737
rect 4977 12703 5095 12737
rect 199 11768 317 11802
rect 351 11768 385 11802
rect 419 11768 453 11802
rect 487 11768 521 11802
rect 555 11768 589 11802
rect 623 11768 657 11802
rect 691 11768 725 11802
rect 759 11768 793 11802
rect 827 11768 861 11802
rect 895 11768 929 11802
rect 963 11768 997 11802
rect 1031 11768 1065 11802
rect 1099 11768 1133 11802
rect 1167 11768 1201 11802
rect 1235 11768 1269 11802
rect 1303 11768 1421 11802
rect 199 11692 233 11768
rect 1387 11692 1421 11768
rect 199 11624 233 11658
rect 199 11556 233 11590
rect 1387 11624 1421 11658
rect 199 11446 233 11522
rect 1387 11556 1421 11590
rect 1387 11446 1421 11522
rect 199 11412 317 11446
rect 351 11412 385 11446
rect 419 11412 453 11446
rect 487 11412 521 11446
rect 555 11412 589 11446
rect 623 11412 657 11446
rect 691 11412 725 11446
rect 759 11412 793 11446
rect 827 11412 861 11446
rect 895 11412 929 11446
rect 963 11412 997 11446
rect 1031 11412 1065 11446
rect 1099 11412 1133 11446
rect 1167 11412 1201 11446
rect 1235 11412 1269 11446
rect 1303 11412 1421 11446
rect 2352 11772 2470 11806
rect 2504 11772 2538 11806
rect 2572 11772 2606 11806
rect 2640 11772 2674 11806
rect 2708 11772 2742 11806
rect 2776 11772 2810 11806
rect 2844 11772 2878 11806
rect 2912 11772 2946 11806
rect 2980 11772 3014 11806
rect 3048 11772 3082 11806
rect 3116 11772 3150 11806
rect 3184 11772 3218 11806
rect 3252 11772 3286 11806
rect 3320 11772 3354 11806
rect 3388 11772 3422 11806
rect 3456 11772 3574 11806
rect 2352 11696 2386 11772
rect 3540 11696 3574 11772
rect 3873 11772 3991 11806
rect 4025 11772 4059 11806
rect 4093 11772 4127 11806
rect 4161 11772 4195 11806
rect 4229 11772 4263 11806
rect 4297 11772 4331 11806
rect 4365 11772 4399 11806
rect 4433 11772 4467 11806
rect 4501 11772 4535 11806
rect 4569 11772 4603 11806
rect 4637 11772 4671 11806
rect 4705 11772 4739 11806
rect 4773 11772 4807 11806
rect 4841 11772 4875 11806
rect 4909 11772 4943 11806
rect 4977 11772 5095 11806
rect 2352 11628 2386 11662
rect 2352 11560 2386 11594
rect 3540 11628 3574 11662
rect 3873 11696 3907 11772
rect 5061 11696 5095 11772
rect 3873 11628 3907 11662
rect 2352 11450 2386 11526
rect 3540 11560 3574 11594
rect 3540 11450 3574 11526
rect 2352 11416 2470 11450
rect 2504 11416 2538 11450
rect 2572 11416 2606 11450
rect 2640 11416 2674 11450
rect 2708 11416 2742 11450
rect 2776 11416 2810 11450
rect 2844 11416 2878 11450
rect 2912 11416 2946 11450
rect 2980 11416 3014 11450
rect 3048 11416 3082 11450
rect 3116 11416 3150 11450
rect 3184 11416 3218 11450
rect 3252 11416 3286 11450
rect 3320 11416 3354 11450
rect 3388 11416 3422 11450
rect 3456 11416 3574 11450
rect 3873 11560 3907 11594
rect 5061 11628 5095 11662
rect 3873 11450 3907 11526
rect 5061 11560 5095 11594
rect 5061 11450 5095 11526
rect 3873 11416 3991 11450
rect 4025 11416 4059 11450
rect 4093 11416 4127 11450
rect 4161 11416 4195 11450
rect 4229 11416 4263 11450
rect 4297 11416 4331 11450
rect 4365 11416 4399 11450
rect 4433 11416 4467 11450
rect 4501 11416 4535 11450
rect 4569 11416 4603 11450
rect 4637 11416 4671 11450
rect 4705 11416 4739 11450
rect 4773 11416 4807 11450
rect 4841 11416 4875 11450
rect 4909 11416 4943 11450
rect 4977 11416 5095 11450
rect 199 10481 317 10515
rect 351 10481 385 10515
rect 419 10481 453 10515
rect 487 10481 521 10515
rect 555 10481 589 10515
rect 623 10481 657 10515
rect 691 10481 725 10515
rect 759 10481 793 10515
rect 827 10481 861 10515
rect 895 10481 929 10515
rect 963 10481 997 10515
rect 1031 10481 1065 10515
rect 1099 10481 1133 10515
rect 1167 10481 1201 10515
rect 1235 10481 1269 10515
rect 1303 10481 1421 10515
rect 199 10405 233 10481
rect 1387 10405 1421 10481
rect 199 10337 233 10371
rect 199 10269 233 10303
rect 1387 10337 1421 10371
rect 199 10159 233 10235
rect 1387 10269 1421 10303
rect 1387 10159 1421 10235
rect 199 10125 317 10159
rect 351 10125 385 10159
rect 419 10125 453 10159
rect 487 10125 521 10159
rect 555 10125 589 10159
rect 623 10125 657 10159
rect 691 10125 725 10159
rect 759 10125 793 10159
rect 827 10125 861 10159
rect 895 10125 929 10159
rect 963 10125 997 10159
rect 1031 10125 1065 10159
rect 1099 10125 1133 10159
rect 1167 10125 1201 10159
rect 1235 10125 1269 10159
rect 1303 10125 1421 10159
rect 2352 10485 2470 10519
rect 2504 10485 2538 10519
rect 2572 10485 2606 10519
rect 2640 10485 2674 10519
rect 2708 10485 2742 10519
rect 2776 10485 2810 10519
rect 2844 10485 2878 10519
rect 2912 10485 2946 10519
rect 2980 10485 3014 10519
rect 3048 10485 3082 10519
rect 3116 10485 3150 10519
rect 3184 10485 3218 10519
rect 3252 10485 3286 10519
rect 3320 10485 3354 10519
rect 3388 10485 3422 10519
rect 3456 10485 3574 10519
rect 2352 10409 2386 10485
rect 3540 10409 3574 10485
rect 3873 10485 3991 10519
rect 4025 10485 4059 10519
rect 4093 10485 4127 10519
rect 4161 10485 4195 10519
rect 4229 10485 4263 10519
rect 4297 10485 4331 10519
rect 4365 10485 4399 10519
rect 4433 10485 4467 10519
rect 4501 10485 4535 10519
rect 4569 10485 4603 10519
rect 4637 10485 4671 10519
rect 4705 10485 4739 10519
rect 4773 10485 4807 10519
rect 4841 10485 4875 10519
rect 4909 10485 4943 10519
rect 4977 10485 5095 10519
rect 2352 10341 2386 10375
rect 2352 10273 2386 10307
rect 3540 10341 3574 10375
rect 3873 10409 3907 10485
rect 5061 10409 5095 10485
rect 3873 10341 3907 10375
rect 2352 10163 2386 10239
rect 3540 10273 3574 10307
rect 3540 10163 3574 10239
rect 2352 10129 2470 10163
rect 2504 10129 2538 10163
rect 2572 10129 2606 10163
rect 2640 10129 2674 10163
rect 2708 10129 2742 10163
rect 2776 10129 2810 10163
rect 2844 10129 2878 10163
rect 2912 10129 2946 10163
rect 2980 10129 3014 10163
rect 3048 10129 3082 10163
rect 3116 10129 3150 10163
rect 3184 10129 3218 10163
rect 3252 10129 3286 10163
rect 3320 10129 3354 10163
rect 3388 10129 3422 10163
rect 3456 10129 3574 10163
rect 3873 10273 3907 10307
rect 5061 10341 5095 10375
rect 3873 10163 3907 10239
rect 5061 10273 5095 10307
rect 5061 10163 5095 10239
rect 3873 10129 3991 10163
rect 4025 10129 4059 10163
rect 4093 10129 4127 10163
rect 4161 10129 4195 10163
rect 4229 10129 4263 10163
rect 4297 10129 4331 10163
rect 4365 10129 4399 10163
rect 4433 10129 4467 10163
rect 4501 10129 4535 10163
rect 4569 10129 4603 10163
rect 4637 10129 4671 10163
rect 4705 10129 4739 10163
rect 4773 10129 4807 10163
rect 4841 10129 4875 10163
rect 4909 10129 4943 10163
rect 4977 10129 5095 10163
rect 199 9194 317 9228
rect 351 9194 385 9228
rect 419 9194 453 9228
rect 487 9194 521 9228
rect 555 9194 589 9228
rect 623 9194 657 9228
rect 691 9194 725 9228
rect 759 9194 793 9228
rect 827 9194 861 9228
rect 895 9194 929 9228
rect 963 9194 997 9228
rect 1031 9194 1065 9228
rect 1099 9194 1133 9228
rect 1167 9194 1201 9228
rect 1235 9194 1269 9228
rect 1303 9194 1421 9228
rect 199 9118 233 9194
rect 1387 9118 1421 9194
rect 199 9050 233 9084
rect 199 8982 233 9016
rect 1387 9050 1421 9084
rect 199 8872 233 8948
rect 1387 8982 1421 9016
rect 1387 8872 1421 8948
rect 199 8838 317 8872
rect 351 8838 385 8872
rect 419 8838 453 8872
rect 487 8838 521 8872
rect 555 8838 589 8872
rect 623 8838 657 8872
rect 691 8838 725 8872
rect 759 8838 793 8872
rect 827 8838 861 8872
rect 895 8838 929 8872
rect 963 8838 997 8872
rect 1031 8838 1065 8872
rect 1099 8838 1133 8872
rect 1167 8838 1201 8872
rect 1235 8838 1269 8872
rect 1303 8838 1421 8872
rect 2352 9198 2470 9232
rect 2504 9198 2538 9232
rect 2572 9198 2606 9232
rect 2640 9198 2674 9232
rect 2708 9198 2742 9232
rect 2776 9198 2810 9232
rect 2844 9198 2878 9232
rect 2912 9198 2946 9232
rect 2980 9198 3014 9232
rect 3048 9198 3082 9232
rect 3116 9198 3150 9232
rect 3184 9198 3218 9232
rect 3252 9198 3286 9232
rect 3320 9198 3354 9232
rect 3388 9198 3422 9232
rect 3456 9198 3574 9232
rect 2352 9122 2386 9198
rect 3540 9122 3574 9198
rect 3873 9198 3991 9232
rect 4025 9198 4059 9232
rect 4093 9198 4127 9232
rect 4161 9198 4195 9232
rect 4229 9198 4263 9232
rect 4297 9198 4331 9232
rect 4365 9198 4399 9232
rect 4433 9198 4467 9232
rect 4501 9198 4535 9232
rect 4569 9198 4603 9232
rect 4637 9198 4671 9232
rect 4705 9198 4739 9232
rect 4773 9198 4807 9232
rect 4841 9198 4875 9232
rect 4909 9198 4943 9232
rect 4977 9198 5095 9232
rect 2352 9054 2386 9088
rect 2352 8986 2386 9020
rect 3540 9054 3574 9088
rect 3873 9122 3907 9198
rect 5061 9122 5095 9198
rect 3873 9054 3907 9088
rect 2352 8876 2386 8952
rect 3540 8986 3574 9020
rect 3540 8876 3574 8952
rect 2352 8842 2470 8876
rect 2504 8842 2538 8876
rect 2572 8842 2606 8876
rect 2640 8842 2674 8876
rect 2708 8842 2742 8876
rect 2776 8842 2810 8876
rect 2844 8842 2878 8876
rect 2912 8842 2946 8876
rect 2980 8842 3014 8876
rect 3048 8842 3082 8876
rect 3116 8842 3150 8876
rect 3184 8842 3218 8876
rect 3252 8842 3286 8876
rect 3320 8842 3354 8876
rect 3388 8842 3422 8876
rect 3456 8842 3574 8876
rect 3873 8986 3907 9020
rect 5061 9054 5095 9088
rect 3873 8876 3907 8952
rect 5061 8986 5095 9020
rect 5061 8876 5095 8952
rect 3873 8842 3991 8876
rect 4025 8842 4059 8876
rect 4093 8842 4127 8876
rect 4161 8842 4195 8876
rect 4229 8842 4263 8876
rect 4297 8842 4331 8876
rect 4365 8842 4399 8876
rect 4433 8842 4467 8876
rect 4501 8842 4535 8876
rect 4569 8842 4603 8876
rect 4637 8842 4671 8876
rect 4705 8842 4739 8876
rect 4773 8842 4807 8876
rect 4841 8842 4875 8876
rect 4909 8842 4943 8876
rect 4977 8842 5095 8876
rect 199 7907 317 7941
rect 351 7907 385 7941
rect 419 7907 453 7941
rect 487 7907 521 7941
rect 555 7907 589 7941
rect 623 7907 657 7941
rect 691 7907 725 7941
rect 759 7907 793 7941
rect 827 7907 861 7941
rect 895 7907 929 7941
rect 963 7907 997 7941
rect 1031 7907 1065 7941
rect 1099 7907 1133 7941
rect 1167 7907 1201 7941
rect 1235 7907 1269 7941
rect 1303 7907 1421 7941
rect 199 7831 233 7907
rect 1387 7831 1421 7907
rect 199 7763 233 7797
rect 199 7695 233 7729
rect 1387 7763 1421 7797
rect 199 7585 233 7661
rect 1387 7695 1421 7729
rect 1387 7585 1421 7661
rect 199 7551 317 7585
rect 351 7551 385 7585
rect 419 7551 453 7585
rect 487 7551 521 7585
rect 555 7551 589 7585
rect 623 7551 657 7585
rect 691 7551 725 7585
rect 759 7551 793 7585
rect 827 7551 861 7585
rect 895 7551 929 7585
rect 963 7551 997 7585
rect 1031 7551 1065 7585
rect 1099 7551 1133 7585
rect 1167 7551 1201 7585
rect 1235 7551 1269 7585
rect 1303 7551 1421 7585
rect 2352 7911 2470 7945
rect 2504 7911 2538 7945
rect 2572 7911 2606 7945
rect 2640 7911 2674 7945
rect 2708 7911 2742 7945
rect 2776 7911 2810 7945
rect 2844 7911 2878 7945
rect 2912 7911 2946 7945
rect 2980 7911 3014 7945
rect 3048 7911 3082 7945
rect 3116 7911 3150 7945
rect 3184 7911 3218 7945
rect 3252 7911 3286 7945
rect 3320 7911 3354 7945
rect 3388 7911 3422 7945
rect 3456 7911 3574 7945
rect 2352 7835 2386 7911
rect 3540 7835 3574 7911
rect 3873 7911 3991 7945
rect 4025 7911 4059 7945
rect 4093 7911 4127 7945
rect 4161 7911 4195 7945
rect 4229 7911 4263 7945
rect 4297 7911 4331 7945
rect 4365 7911 4399 7945
rect 4433 7911 4467 7945
rect 4501 7911 4535 7945
rect 4569 7911 4603 7945
rect 4637 7911 4671 7945
rect 4705 7911 4739 7945
rect 4773 7911 4807 7945
rect 4841 7911 4875 7945
rect 4909 7911 4943 7945
rect 4977 7911 5095 7945
rect 2352 7767 2386 7801
rect 2352 7699 2386 7733
rect 3540 7767 3574 7801
rect 3873 7835 3907 7911
rect 5061 7835 5095 7911
rect 3873 7767 3907 7801
rect 2352 7589 2386 7665
rect 3540 7699 3574 7733
rect 3540 7589 3574 7665
rect 2352 7555 2470 7589
rect 2504 7555 2538 7589
rect 2572 7555 2606 7589
rect 2640 7555 2674 7589
rect 2708 7555 2742 7589
rect 2776 7555 2810 7589
rect 2844 7555 2878 7589
rect 2912 7555 2946 7589
rect 2980 7555 3014 7589
rect 3048 7555 3082 7589
rect 3116 7555 3150 7589
rect 3184 7555 3218 7589
rect 3252 7555 3286 7589
rect 3320 7555 3354 7589
rect 3388 7555 3422 7589
rect 3456 7555 3574 7589
rect 3873 7699 3907 7733
rect 5061 7767 5095 7801
rect 3873 7589 3907 7665
rect 5061 7699 5095 7733
rect 5061 7589 5095 7665
rect 3873 7555 3991 7589
rect 4025 7555 4059 7589
rect 4093 7555 4127 7589
rect 4161 7555 4195 7589
rect 4229 7555 4263 7589
rect 4297 7555 4331 7589
rect 4365 7555 4399 7589
rect 4433 7555 4467 7589
rect 4501 7555 4535 7589
rect 4569 7555 4603 7589
rect 4637 7555 4671 7589
rect 4705 7555 4739 7589
rect 4773 7555 4807 7589
rect 4841 7555 4875 7589
rect 4909 7555 4943 7589
rect 4977 7555 5095 7589
rect 199 6620 317 6654
rect 351 6620 385 6654
rect 419 6620 453 6654
rect 487 6620 521 6654
rect 555 6620 589 6654
rect 623 6620 657 6654
rect 691 6620 725 6654
rect 759 6620 793 6654
rect 827 6620 861 6654
rect 895 6620 929 6654
rect 963 6620 997 6654
rect 1031 6620 1065 6654
rect 1099 6620 1133 6654
rect 1167 6620 1201 6654
rect 1235 6620 1269 6654
rect 1303 6620 1421 6654
rect 199 6544 233 6620
rect 1387 6544 1421 6620
rect 199 6476 233 6510
rect 199 6408 233 6442
rect 1387 6476 1421 6510
rect 199 6298 233 6374
rect 1387 6408 1421 6442
rect 1387 6298 1421 6374
rect 199 6264 317 6298
rect 351 6264 385 6298
rect 419 6264 453 6298
rect 487 6264 521 6298
rect 555 6264 589 6298
rect 623 6264 657 6298
rect 691 6264 725 6298
rect 759 6264 793 6298
rect 827 6264 861 6298
rect 895 6264 929 6298
rect 963 6264 997 6298
rect 1031 6264 1065 6298
rect 1099 6264 1133 6298
rect 1167 6264 1201 6298
rect 1235 6264 1269 6298
rect 1303 6264 1421 6298
rect 2352 6624 2470 6658
rect 2504 6624 2538 6658
rect 2572 6624 2606 6658
rect 2640 6624 2674 6658
rect 2708 6624 2742 6658
rect 2776 6624 2810 6658
rect 2844 6624 2878 6658
rect 2912 6624 2946 6658
rect 2980 6624 3014 6658
rect 3048 6624 3082 6658
rect 3116 6624 3150 6658
rect 3184 6624 3218 6658
rect 3252 6624 3286 6658
rect 3320 6624 3354 6658
rect 3388 6624 3422 6658
rect 3456 6624 3574 6658
rect 2352 6548 2386 6624
rect 3540 6548 3574 6624
rect 3873 6624 3991 6658
rect 4025 6624 4059 6658
rect 4093 6624 4127 6658
rect 4161 6624 4195 6658
rect 4229 6624 4263 6658
rect 4297 6624 4331 6658
rect 4365 6624 4399 6658
rect 4433 6624 4467 6658
rect 4501 6624 4535 6658
rect 4569 6624 4603 6658
rect 4637 6624 4671 6658
rect 4705 6624 4739 6658
rect 4773 6624 4807 6658
rect 4841 6624 4875 6658
rect 4909 6624 4943 6658
rect 4977 6624 5095 6658
rect 2352 6480 2386 6514
rect 2352 6412 2386 6446
rect 3540 6480 3574 6514
rect 3873 6548 3907 6624
rect 5061 6548 5095 6624
rect 3873 6480 3907 6514
rect 2352 6302 2386 6378
rect 3540 6412 3574 6446
rect 3540 6302 3574 6378
rect 2352 6268 2470 6302
rect 2504 6268 2538 6302
rect 2572 6268 2606 6302
rect 2640 6268 2674 6302
rect 2708 6268 2742 6302
rect 2776 6268 2810 6302
rect 2844 6268 2878 6302
rect 2912 6268 2946 6302
rect 2980 6268 3014 6302
rect 3048 6268 3082 6302
rect 3116 6268 3150 6302
rect 3184 6268 3218 6302
rect 3252 6268 3286 6302
rect 3320 6268 3354 6302
rect 3388 6268 3422 6302
rect 3456 6268 3574 6302
rect 3873 6412 3907 6446
rect 5061 6480 5095 6514
rect 3873 6302 3907 6378
rect 5061 6412 5095 6446
rect 5061 6302 5095 6378
rect 3873 6268 3991 6302
rect 4025 6268 4059 6302
rect 4093 6268 4127 6302
rect 4161 6268 4195 6302
rect 4229 6268 4263 6302
rect 4297 6268 4331 6302
rect 4365 6268 4399 6302
rect 4433 6268 4467 6302
rect 4501 6268 4535 6302
rect 4569 6268 4603 6302
rect 4637 6268 4671 6302
rect 4705 6268 4739 6302
rect 4773 6268 4807 6302
rect 4841 6268 4875 6302
rect 4909 6268 4943 6302
rect 4977 6268 5095 6302
rect 199 5333 317 5367
rect 351 5333 385 5367
rect 419 5333 453 5367
rect 487 5333 521 5367
rect 555 5333 589 5367
rect 623 5333 657 5367
rect 691 5333 725 5367
rect 759 5333 793 5367
rect 827 5333 861 5367
rect 895 5333 929 5367
rect 963 5333 997 5367
rect 1031 5333 1065 5367
rect 1099 5333 1133 5367
rect 1167 5333 1201 5367
rect 1235 5333 1269 5367
rect 1303 5333 1421 5367
rect 199 5257 233 5333
rect 1387 5257 1421 5333
rect 199 5189 233 5223
rect 199 5121 233 5155
rect 1387 5189 1421 5223
rect 199 5011 233 5087
rect 1387 5121 1421 5155
rect 1387 5011 1421 5087
rect 199 4977 317 5011
rect 351 4977 385 5011
rect 419 4977 453 5011
rect 487 4977 521 5011
rect 555 4977 589 5011
rect 623 4977 657 5011
rect 691 4977 725 5011
rect 759 4977 793 5011
rect 827 4977 861 5011
rect 895 4977 929 5011
rect 963 4977 997 5011
rect 1031 4977 1065 5011
rect 1099 4977 1133 5011
rect 1167 4977 1201 5011
rect 1235 4977 1269 5011
rect 1303 4977 1421 5011
rect 2352 5337 2470 5371
rect 2504 5337 2538 5371
rect 2572 5337 2606 5371
rect 2640 5337 2674 5371
rect 2708 5337 2742 5371
rect 2776 5337 2810 5371
rect 2844 5337 2878 5371
rect 2912 5337 2946 5371
rect 2980 5337 3014 5371
rect 3048 5337 3082 5371
rect 3116 5337 3150 5371
rect 3184 5337 3218 5371
rect 3252 5337 3286 5371
rect 3320 5337 3354 5371
rect 3388 5337 3422 5371
rect 3456 5337 3574 5371
rect 2352 5261 2386 5337
rect 3540 5261 3574 5337
rect 3873 5337 3991 5371
rect 4025 5337 4059 5371
rect 4093 5337 4127 5371
rect 4161 5337 4195 5371
rect 4229 5337 4263 5371
rect 4297 5337 4331 5371
rect 4365 5337 4399 5371
rect 4433 5337 4467 5371
rect 4501 5337 4535 5371
rect 4569 5337 4603 5371
rect 4637 5337 4671 5371
rect 4705 5337 4739 5371
rect 4773 5337 4807 5371
rect 4841 5337 4875 5371
rect 4909 5337 4943 5371
rect 4977 5337 5095 5371
rect 2352 5193 2386 5227
rect 2352 5125 2386 5159
rect 3540 5193 3574 5227
rect 3873 5261 3907 5337
rect 5061 5261 5095 5337
rect 3873 5193 3907 5227
rect 2352 5015 2386 5091
rect 3540 5125 3574 5159
rect 3540 5015 3574 5091
rect 2352 4981 2470 5015
rect 2504 4981 2538 5015
rect 2572 4981 2606 5015
rect 2640 4981 2674 5015
rect 2708 4981 2742 5015
rect 2776 4981 2810 5015
rect 2844 4981 2878 5015
rect 2912 4981 2946 5015
rect 2980 4981 3014 5015
rect 3048 4981 3082 5015
rect 3116 4981 3150 5015
rect 3184 4981 3218 5015
rect 3252 4981 3286 5015
rect 3320 4981 3354 5015
rect 3388 4981 3422 5015
rect 3456 4981 3574 5015
rect 3873 5125 3907 5159
rect 5061 5193 5095 5227
rect 3873 5015 3907 5091
rect 5061 5125 5095 5159
rect 5061 5015 5095 5091
rect 3873 4981 3991 5015
rect 4025 4981 4059 5015
rect 4093 4981 4127 5015
rect 4161 4981 4195 5015
rect 4229 4981 4263 5015
rect 4297 4981 4331 5015
rect 4365 4981 4399 5015
rect 4433 4981 4467 5015
rect 4501 4981 4535 5015
rect 4569 4981 4603 5015
rect 4637 4981 4671 5015
rect 4705 4981 4739 5015
rect 4773 4981 4807 5015
rect 4841 4981 4875 5015
rect 4909 4981 4943 5015
rect 4977 4981 5095 5015
rect 199 4046 317 4080
rect 351 4046 385 4080
rect 419 4046 453 4080
rect 487 4046 521 4080
rect 555 4046 589 4080
rect 623 4046 657 4080
rect 691 4046 725 4080
rect 759 4046 793 4080
rect 827 4046 861 4080
rect 895 4046 929 4080
rect 963 4046 997 4080
rect 1031 4046 1065 4080
rect 1099 4046 1133 4080
rect 1167 4046 1201 4080
rect 1235 4046 1269 4080
rect 1303 4046 1421 4080
rect 199 3970 233 4046
rect 1387 3970 1421 4046
rect 199 3902 233 3936
rect 199 3834 233 3868
rect 1387 3902 1421 3936
rect 199 3724 233 3800
rect 1387 3834 1421 3868
rect 1387 3724 1421 3800
rect 199 3690 317 3724
rect 351 3690 385 3724
rect 419 3690 453 3724
rect 487 3690 521 3724
rect 555 3690 589 3724
rect 623 3690 657 3724
rect 691 3690 725 3724
rect 759 3690 793 3724
rect 827 3690 861 3724
rect 895 3690 929 3724
rect 963 3690 997 3724
rect 1031 3690 1065 3724
rect 1099 3690 1133 3724
rect 1167 3690 1201 3724
rect 1235 3690 1269 3724
rect 1303 3690 1421 3724
rect 2352 4050 2470 4084
rect 2504 4050 2538 4084
rect 2572 4050 2606 4084
rect 2640 4050 2674 4084
rect 2708 4050 2742 4084
rect 2776 4050 2810 4084
rect 2844 4050 2878 4084
rect 2912 4050 2946 4084
rect 2980 4050 3014 4084
rect 3048 4050 3082 4084
rect 3116 4050 3150 4084
rect 3184 4050 3218 4084
rect 3252 4050 3286 4084
rect 3320 4050 3354 4084
rect 3388 4050 3422 4084
rect 3456 4050 3574 4084
rect 2352 3974 2386 4050
rect 3540 3974 3574 4050
rect 3873 4050 3991 4084
rect 4025 4050 4059 4084
rect 4093 4050 4127 4084
rect 4161 4050 4195 4084
rect 4229 4050 4263 4084
rect 4297 4050 4331 4084
rect 4365 4050 4399 4084
rect 4433 4050 4467 4084
rect 4501 4050 4535 4084
rect 4569 4050 4603 4084
rect 4637 4050 4671 4084
rect 4705 4050 4739 4084
rect 4773 4050 4807 4084
rect 4841 4050 4875 4084
rect 4909 4050 4943 4084
rect 4977 4050 5095 4084
rect 2352 3906 2386 3940
rect 2352 3838 2386 3872
rect 3540 3906 3574 3940
rect 3873 3974 3907 4050
rect 5061 3974 5095 4050
rect 3873 3906 3907 3940
rect 2352 3728 2386 3804
rect 3540 3838 3574 3872
rect 3540 3728 3574 3804
rect 2352 3694 2470 3728
rect 2504 3694 2538 3728
rect 2572 3694 2606 3728
rect 2640 3694 2674 3728
rect 2708 3694 2742 3728
rect 2776 3694 2810 3728
rect 2844 3694 2878 3728
rect 2912 3694 2946 3728
rect 2980 3694 3014 3728
rect 3048 3694 3082 3728
rect 3116 3694 3150 3728
rect 3184 3694 3218 3728
rect 3252 3694 3286 3728
rect 3320 3694 3354 3728
rect 3388 3694 3422 3728
rect 3456 3694 3574 3728
rect 3873 3838 3907 3872
rect 5061 3906 5095 3940
rect 3873 3728 3907 3804
rect 5061 3838 5095 3872
rect 5061 3728 5095 3804
rect 3873 3694 3991 3728
rect 4025 3694 4059 3728
rect 4093 3694 4127 3728
rect 4161 3694 4195 3728
rect 4229 3694 4263 3728
rect 4297 3694 4331 3728
rect 4365 3694 4399 3728
rect 4433 3694 4467 3728
rect 4501 3694 4535 3728
rect 4569 3694 4603 3728
rect 4637 3694 4671 3728
rect 4705 3694 4739 3728
rect 4773 3694 4807 3728
rect 4841 3694 4875 3728
rect 4909 3694 4943 3728
rect 4977 3694 5095 3728
rect 199 2759 317 2793
rect 351 2759 385 2793
rect 419 2759 453 2793
rect 487 2759 521 2793
rect 555 2759 589 2793
rect 623 2759 657 2793
rect 691 2759 725 2793
rect 759 2759 793 2793
rect 827 2759 861 2793
rect 895 2759 929 2793
rect 963 2759 997 2793
rect 1031 2759 1065 2793
rect 1099 2759 1133 2793
rect 1167 2759 1201 2793
rect 1235 2759 1269 2793
rect 1303 2759 1421 2793
rect 199 2683 233 2759
rect 1387 2683 1421 2759
rect 199 2615 233 2649
rect 199 2547 233 2581
rect 1387 2615 1421 2649
rect 199 2437 233 2513
rect 1387 2547 1421 2581
rect 1387 2437 1421 2513
rect 199 2403 317 2437
rect 351 2403 385 2437
rect 419 2403 453 2437
rect 487 2403 521 2437
rect 555 2403 589 2437
rect 623 2403 657 2437
rect 691 2403 725 2437
rect 759 2403 793 2437
rect 827 2403 861 2437
rect 895 2403 929 2437
rect 963 2403 997 2437
rect 1031 2403 1065 2437
rect 1099 2403 1133 2437
rect 1167 2403 1201 2437
rect 1235 2403 1269 2437
rect 1303 2403 1421 2437
rect 2352 2763 2470 2797
rect 2504 2763 2538 2797
rect 2572 2763 2606 2797
rect 2640 2763 2674 2797
rect 2708 2763 2742 2797
rect 2776 2763 2810 2797
rect 2844 2763 2878 2797
rect 2912 2763 2946 2797
rect 2980 2763 3014 2797
rect 3048 2763 3082 2797
rect 3116 2763 3150 2797
rect 3184 2763 3218 2797
rect 3252 2763 3286 2797
rect 3320 2763 3354 2797
rect 3388 2763 3422 2797
rect 3456 2763 3574 2797
rect 2352 2687 2386 2763
rect 3540 2687 3574 2763
rect 3873 2763 3991 2797
rect 4025 2763 4059 2797
rect 4093 2763 4127 2797
rect 4161 2763 4195 2797
rect 4229 2763 4263 2797
rect 4297 2763 4331 2797
rect 4365 2763 4399 2797
rect 4433 2763 4467 2797
rect 4501 2763 4535 2797
rect 4569 2763 4603 2797
rect 4637 2763 4671 2797
rect 4705 2763 4739 2797
rect 4773 2763 4807 2797
rect 4841 2763 4875 2797
rect 4909 2763 4943 2797
rect 4977 2763 5095 2797
rect 2352 2619 2386 2653
rect 2352 2551 2386 2585
rect 3540 2619 3574 2653
rect 3873 2687 3907 2763
rect 5061 2687 5095 2763
rect 3873 2619 3907 2653
rect 2352 2441 2386 2517
rect 3540 2551 3574 2585
rect 3540 2441 3574 2517
rect 2352 2407 2470 2441
rect 2504 2407 2538 2441
rect 2572 2407 2606 2441
rect 2640 2407 2674 2441
rect 2708 2407 2742 2441
rect 2776 2407 2810 2441
rect 2844 2407 2878 2441
rect 2912 2407 2946 2441
rect 2980 2407 3014 2441
rect 3048 2407 3082 2441
rect 3116 2407 3150 2441
rect 3184 2407 3218 2441
rect 3252 2407 3286 2441
rect 3320 2407 3354 2441
rect 3388 2407 3422 2441
rect 3456 2407 3574 2441
rect 3873 2551 3907 2585
rect 5061 2619 5095 2653
rect 3873 2441 3907 2517
rect 5061 2551 5095 2585
rect 5061 2441 5095 2517
rect 3873 2407 3991 2441
rect 4025 2407 4059 2441
rect 4093 2407 4127 2441
rect 4161 2407 4195 2441
rect 4229 2407 4263 2441
rect 4297 2407 4331 2441
rect 4365 2407 4399 2441
rect 4433 2407 4467 2441
rect 4501 2407 4535 2441
rect 4569 2407 4603 2441
rect 4637 2407 4671 2441
rect 4705 2407 4739 2441
rect 4773 2407 4807 2441
rect 4841 2407 4875 2441
rect 4909 2407 4943 2441
rect 4977 2407 5095 2441
rect 199 1472 317 1506
rect 351 1472 385 1506
rect 419 1472 453 1506
rect 487 1472 521 1506
rect 555 1472 589 1506
rect 623 1472 657 1506
rect 691 1472 725 1506
rect 759 1472 793 1506
rect 827 1472 861 1506
rect 895 1472 929 1506
rect 963 1472 997 1506
rect 1031 1472 1065 1506
rect 1099 1472 1133 1506
rect 1167 1472 1201 1506
rect 1235 1472 1269 1506
rect 1303 1472 1421 1506
rect 199 1396 233 1472
rect 1387 1396 1421 1472
rect 199 1328 233 1362
rect 199 1260 233 1294
rect 1387 1328 1421 1362
rect 199 1150 233 1226
rect 1387 1260 1421 1294
rect 1387 1150 1421 1226
rect 199 1116 317 1150
rect 351 1116 385 1150
rect 419 1116 453 1150
rect 487 1116 521 1150
rect 555 1116 589 1150
rect 623 1116 657 1150
rect 691 1116 725 1150
rect 759 1116 793 1150
rect 827 1116 861 1150
rect 895 1116 929 1150
rect 963 1116 997 1150
rect 1031 1116 1065 1150
rect 1099 1116 1133 1150
rect 1167 1116 1201 1150
rect 1235 1116 1269 1150
rect 1303 1116 1421 1150
rect 2352 1476 2470 1510
rect 2504 1476 2538 1510
rect 2572 1476 2606 1510
rect 2640 1476 2674 1510
rect 2708 1476 2742 1510
rect 2776 1476 2810 1510
rect 2844 1476 2878 1510
rect 2912 1476 2946 1510
rect 2980 1476 3014 1510
rect 3048 1476 3082 1510
rect 3116 1476 3150 1510
rect 3184 1476 3218 1510
rect 3252 1476 3286 1510
rect 3320 1476 3354 1510
rect 3388 1476 3422 1510
rect 3456 1476 3574 1510
rect 2352 1400 2386 1476
rect 3540 1400 3574 1476
rect 3873 1476 3991 1510
rect 4025 1476 4059 1510
rect 4093 1476 4127 1510
rect 4161 1476 4195 1510
rect 4229 1476 4263 1510
rect 4297 1476 4331 1510
rect 4365 1476 4399 1510
rect 4433 1476 4467 1510
rect 4501 1476 4535 1510
rect 4569 1476 4603 1510
rect 4637 1476 4671 1510
rect 4705 1476 4739 1510
rect 4773 1476 4807 1510
rect 4841 1476 4875 1510
rect 4909 1476 4943 1510
rect 4977 1476 5095 1510
rect 2352 1332 2386 1366
rect 2352 1264 2386 1298
rect 3540 1332 3574 1366
rect 3873 1400 3907 1476
rect 5061 1400 5095 1476
rect 3873 1332 3907 1366
rect 2352 1154 2386 1230
rect 3540 1264 3574 1298
rect 3540 1154 3574 1230
rect 2352 1120 2470 1154
rect 2504 1120 2538 1154
rect 2572 1120 2606 1154
rect 2640 1120 2674 1154
rect 2708 1120 2742 1154
rect 2776 1120 2810 1154
rect 2844 1120 2878 1154
rect 2912 1120 2946 1154
rect 2980 1120 3014 1154
rect 3048 1120 3082 1154
rect 3116 1120 3150 1154
rect 3184 1120 3218 1154
rect 3252 1120 3286 1154
rect 3320 1120 3354 1154
rect 3388 1120 3422 1154
rect 3456 1120 3574 1154
rect 3873 1264 3907 1298
rect 5061 1332 5095 1366
rect 3873 1154 3907 1230
rect 5061 1264 5095 1298
rect 5061 1154 5095 1230
rect 3873 1120 3991 1154
rect 4025 1120 4059 1154
rect 4093 1120 4127 1154
rect 4161 1120 4195 1154
rect 4229 1120 4263 1154
rect 4297 1120 4331 1154
rect 4365 1120 4399 1154
rect 4433 1120 4467 1154
rect 4501 1120 4535 1154
rect 4569 1120 4603 1154
rect 4637 1120 4671 1154
rect 4705 1120 4739 1154
rect 4773 1120 4807 1154
rect 4841 1120 4875 1154
rect 4909 1120 4943 1154
rect 4977 1120 5095 1154
<< nsubdiff >>
rect 199 42021 317 42055
rect 351 42021 385 42055
rect 419 42021 453 42055
rect 487 42021 521 42055
rect 555 42021 589 42055
rect 623 42021 657 42055
rect 691 42021 725 42055
rect 759 42021 793 42055
rect 827 42021 861 42055
rect 895 42021 929 42055
rect 963 42021 997 42055
rect 1031 42021 1065 42055
rect 1099 42021 1133 42055
rect 1167 42021 1201 42055
rect 1235 42021 1269 42055
rect 1303 42021 1421 42055
rect 199 41953 233 42021
rect 199 41885 233 41919
rect 1387 41953 1421 42021
rect 1387 41885 1421 41919
rect 199 41817 233 41851
rect 199 41749 233 41783
rect 199 41681 233 41715
rect 199 41613 233 41647
rect 1387 41817 1421 41851
rect 1387 41749 1421 41783
rect 1387 41681 1421 41715
rect 1387 41613 1421 41647
rect 199 41511 233 41579
rect 1387 41511 1421 41579
rect 199 41477 317 41511
rect 351 41477 385 41511
rect 419 41477 453 41511
rect 487 41477 521 41511
rect 555 41477 589 41511
rect 623 41477 657 41511
rect 691 41477 725 41511
rect 759 41477 793 41511
rect 827 41477 861 41511
rect 895 41477 929 41511
rect 963 41477 997 41511
rect 1031 41477 1065 41511
rect 1099 41477 1133 41511
rect 1167 41477 1201 41511
rect 1235 41477 1269 41511
rect 1303 41477 1421 41511
rect 2352 42025 2470 42059
rect 2504 42025 2538 42059
rect 2572 42025 2606 42059
rect 2640 42025 2674 42059
rect 2708 42025 2742 42059
rect 2776 42025 2810 42059
rect 2844 42025 2878 42059
rect 2912 42025 2946 42059
rect 2980 42025 3014 42059
rect 3048 42025 3082 42059
rect 3116 42025 3150 42059
rect 3184 42025 3218 42059
rect 3252 42025 3286 42059
rect 3320 42025 3354 42059
rect 3388 42025 3422 42059
rect 3456 42025 3574 42059
rect 2352 41957 2386 42025
rect 2352 41889 2386 41923
rect 3540 41957 3574 42025
rect 3540 41889 3574 41923
rect 2352 41821 2386 41855
rect 2352 41753 2386 41787
rect 2352 41685 2386 41719
rect 2352 41617 2386 41651
rect 3540 41821 3574 41855
rect 3540 41753 3574 41787
rect 3540 41685 3574 41719
rect 3540 41617 3574 41651
rect 2352 41515 2386 41583
rect 3540 41515 3574 41583
rect 2352 41481 2470 41515
rect 2504 41481 2538 41515
rect 2572 41481 2606 41515
rect 2640 41481 2674 41515
rect 2708 41481 2742 41515
rect 2776 41481 2810 41515
rect 2844 41481 2878 41515
rect 2912 41481 2946 41515
rect 2980 41481 3014 41515
rect 3048 41481 3082 41515
rect 3116 41481 3150 41515
rect 3184 41481 3218 41515
rect 3252 41481 3286 41515
rect 3320 41481 3354 41515
rect 3388 41481 3422 41515
rect 3456 41481 3574 41515
rect 3873 42025 3991 42059
rect 4025 42025 4059 42059
rect 4093 42025 4127 42059
rect 4161 42025 4195 42059
rect 4229 42025 4263 42059
rect 4297 42025 4331 42059
rect 4365 42025 4399 42059
rect 4433 42025 4467 42059
rect 4501 42025 4535 42059
rect 4569 42025 4603 42059
rect 4637 42025 4671 42059
rect 4705 42025 4739 42059
rect 4773 42025 4807 42059
rect 4841 42025 4875 42059
rect 4909 42025 4943 42059
rect 4977 42025 5095 42059
rect 3873 41957 3907 42025
rect 3873 41889 3907 41923
rect 5061 41957 5095 42025
rect 5061 41889 5095 41923
rect 3873 41821 3907 41855
rect 3873 41753 3907 41787
rect 3873 41685 3907 41719
rect 3873 41617 3907 41651
rect 5061 41821 5095 41855
rect 5061 41753 5095 41787
rect 5061 41685 5095 41719
rect 5061 41617 5095 41651
rect 3873 41515 3907 41583
rect 5061 41515 5095 41583
rect 3873 41481 3991 41515
rect 4025 41481 4059 41515
rect 4093 41481 4127 41515
rect 4161 41481 4195 41515
rect 4229 41481 4263 41515
rect 4297 41481 4331 41515
rect 4365 41481 4399 41515
rect 4433 41481 4467 41515
rect 4501 41481 4535 41515
rect 4569 41481 4603 41515
rect 4637 41481 4671 41515
rect 4705 41481 4739 41515
rect 4773 41481 4807 41515
rect 4841 41481 4875 41515
rect 4909 41481 4943 41515
rect 4977 41481 5095 41515
rect 199 40734 317 40768
rect 351 40734 385 40768
rect 419 40734 453 40768
rect 487 40734 521 40768
rect 555 40734 589 40768
rect 623 40734 657 40768
rect 691 40734 725 40768
rect 759 40734 793 40768
rect 827 40734 861 40768
rect 895 40734 929 40768
rect 963 40734 997 40768
rect 1031 40734 1065 40768
rect 1099 40734 1133 40768
rect 1167 40734 1201 40768
rect 1235 40734 1269 40768
rect 1303 40734 1421 40768
rect 199 40666 233 40734
rect 199 40598 233 40632
rect 1387 40666 1421 40734
rect 1387 40598 1421 40632
rect 199 40530 233 40564
rect 199 40462 233 40496
rect 199 40394 233 40428
rect 199 40326 233 40360
rect 1387 40530 1421 40564
rect 1387 40462 1421 40496
rect 1387 40394 1421 40428
rect 1387 40326 1421 40360
rect 199 40224 233 40292
rect 1387 40224 1421 40292
rect 199 40190 317 40224
rect 351 40190 385 40224
rect 419 40190 453 40224
rect 487 40190 521 40224
rect 555 40190 589 40224
rect 623 40190 657 40224
rect 691 40190 725 40224
rect 759 40190 793 40224
rect 827 40190 861 40224
rect 895 40190 929 40224
rect 963 40190 997 40224
rect 1031 40190 1065 40224
rect 1099 40190 1133 40224
rect 1167 40190 1201 40224
rect 1235 40190 1269 40224
rect 1303 40190 1421 40224
rect 2352 40738 2470 40772
rect 2504 40738 2538 40772
rect 2572 40738 2606 40772
rect 2640 40738 2674 40772
rect 2708 40738 2742 40772
rect 2776 40738 2810 40772
rect 2844 40738 2878 40772
rect 2912 40738 2946 40772
rect 2980 40738 3014 40772
rect 3048 40738 3082 40772
rect 3116 40738 3150 40772
rect 3184 40738 3218 40772
rect 3252 40738 3286 40772
rect 3320 40738 3354 40772
rect 3388 40738 3422 40772
rect 3456 40738 3574 40772
rect 2352 40670 2386 40738
rect 2352 40602 2386 40636
rect 3540 40670 3574 40738
rect 3540 40602 3574 40636
rect 2352 40534 2386 40568
rect 2352 40466 2386 40500
rect 2352 40398 2386 40432
rect 2352 40330 2386 40364
rect 3540 40534 3574 40568
rect 3540 40466 3574 40500
rect 3540 40398 3574 40432
rect 3540 40330 3574 40364
rect 2352 40228 2386 40296
rect 3540 40228 3574 40296
rect 2352 40194 2470 40228
rect 2504 40194 2538 40228
rect 2572 40194 2606 40228
rect 2640 40194 2674 40228
rect 2708 40194 2742 40228
rect 2776 40194 2810 40228
rect 2844 40194 2878 40228
rect 2912 40194 2946 40228
rect 2980 40194 3014 40228
rect 3048 40194 3082 40228
rect 3116 40194 3150 40228
rect 3184 40194 3218 40228
rect 3252 40194 3286 40228
rect 3320 40194 3354 40228
rect 3388 40194 3422 40228
rect 3456 40194 3574 40228
rect 3873 40738 3991 40772
rect 4025 40738 4059 40772
rect 4093 40738 4127 40772
rect 4161 40738 4195 40772
rect 4229 40738 4263 40772
rect 4297 40738 4331 40772
rect 4365 40738 4399 40772
rect 4433 40738 4467 40772
rect 4501 40738 4535 40772
rect 4569 40738 4603 40772
rect 4637 40738 4671 40772
rect 4705 40738 4739 40772
rect 4773 40738 4807 40772
rect 4841 40738 4875 40772
rect 4909 40738 4943 40772
rect 4977 40738 5095 40772
rect 3873 40670 3907 40738
rect 3873 40602 3907 40636
rect 5061 40670 5095 40738
rect 5061 40602 5095 40636
rect 3873 40534 3907 40568
rect 3873 40466 3907 40500
rect 3873 40398 3907 40432
rect 3873 40330 3907 40364
rect 5061 40534 5095 40568
rect 5061 40466 5095 40500
rect 5061 40398 5095 40432
rect 5061 40330 5095 40364
rect 3873 40228 3907 40296
rect 5061 40228 5095 40296
rect 3873 40194 3991 40228
rect 4025 40194 4059 40228
rect 4093 40194 4127 40228
rect 4161 40194 4195 40228
rect 4229 40194 4263 40228
rect 4297 40194 4331 40228
rect 4365 40194 4399 40228
rect 4433 40194 4467 40228
rect 4501 40194 4535 40228
rect 4569 40194 4603 40228
rect 4637 40194 4671 40228
rect 4705 40194 4739 40228
rect 4773 40194 4807 40228
rect 4841 40194 4875 40228
rect 4909 40194 4943 40228
rect 4977 40194 5095 40228
rect 199 39447 317 39481
rect 351 39447 385 39481
rect 419 39447 453 39481
rect 487 39447 521 39481
rect 555 39447 589 39481
rect 623 39447 657 39481
rect 691 39447 725 39481
rect 759 39447 793 39481
rect 827 39447 861 39481
rect 895 39447 929 39481
rect 963 39447 997 39481
rect 1031 39447 1065 39481
rect 1099 39447 1133 39481
rect 1167 39447 1201 39481
rect 1235 39447 1269 39481
rect 1303 39447 1421 39481
rect 199 39379 233 39447
rect 199 39311 233 39345
rect 1387 39379 1421 39447
rect 1387 39311 1421 39345
rect 199 39243 233 39277
rect 199 39175 233 39209
rect 199 39107 233 39141
rect 199 39039 233 39073
rect 1387 39243 1421 39277
rect 1387 39175 1421 39209
rect 1387 39107 1421 39141
rect 1387 39039 1421 39073
rect 199 38937 233 39005
rect 1387 38937 1421 39005
rect 199 38903 317 38937
rect 351 38903 385 38937
rect 419 38903 453 38937
rect 487 38903 521 38937
rect 555 38903 589 38937
rect 623 38903 657 38937
rect 691 38903 725 38937
rect 759 38903 793 38937
rect 827 38903 861 38937
rect 895 38903 929 38937
rect 963 38903 997 38937
rect 1031 38903 1065 38937
rect 1099 38903 1133 38937
rect 1167 38903 1201 38937
rect 1235 38903 1269 38937
rect 1303 38903 1421 38937
rect 2352 39451 2470 39485
rect 2504 39451 2538 39485
rect 2572 39451 2606 39485
rect 2640 39451 2674 39485
rect 2708 39451 2742 39485
rect 2776 39451 2810 39485
rect 2844 39451 2878 39485
rect 2912 39451 2946 39485
rect 2980 39451 3014 39485
rect 3048 39451 3082 39485
rect 3116 39451 3150 39485
rect 3184 39451 3218 39485
rect 3252 39451 3286 39485
rect 3320 39451 3354 39485
rect 3388 39451 3422 39485
rect 3456 39451 3574 39485
rect 2352 39383 2386 39451
rect 2352 39315 2386 39349
rect 3540 39383 3574 39451
rect 3540 39315 3574 39349
rect 2352 39247 2386 39281
rect 2352 39179 2386 39213
rect 2352 39111 2386 39145
rect 2352 39043 2386 39077
rect 3540 39247 3574 39281
rect 3540 39179 3574 39213
rect 3540 39111 3574 39145
rect 3540 39043 3574 39077
rect 2352 38941 2386 39009
rect 3540 38941 3574 39009
rect 2352 38907 2470 38941
rect 2504 38907 2538 38941
rect 2572 38907 2606 38941
rect 2640 38907 2674 38941
rect 2708 38907 2742 38941
rect 2776 38907 2810 38941
rect 2844 38907 2878 38941
rect 2912 38907 2946 38941
rect 2980 38907 3014 38941
rect 3048 38907 3082 38941
rect 3116 38907 3150 38941
rect 3184 38907 3218 38941
rect 3252 38907 3286 38941
rect 3320 38907 3354 38941
rect 3388 38907 3422 38941
rect 3456 38907 3574 38941
rect 3873 39451 3991 39485
rect 4025 39451 4059 39485
rect 4093 39451 4127 39485
rect 4161 39451 4195 39485
rect 4229 39451 4263 39485
rect 4297 39451 4331 39485
rect 4365 39451 4399 39485
rect 4433 39451 4467 39485
rect 4501 39451 4535 39485
rect 4569 39451 4603 39485
rect 4637 39451 4671 39485
rect 4705 39451 4739 39485
rect 4773 39451 4807 39485
rect 4841 39451 4875 39485
rect 4909 39451 4943 39485
rect 4977 39451 5095 39485
rect 3873 39383 3907 39451
rect 3873 39315 3907 39349
rect 5061 39383 5095 39451
rect 5061 39315 5095 39349
rect 3873 39247 3907 39281
rect 3873 39179 3907 39213
rect 3873 39111 3907 39145
rect 3873 39043 3907 39077
rect 5061 39247 5095 39281
rect 5061 39179 5095 39213
rect 5061 39111 5095 39145
rect 5061 39043 5095 39077
rect 3873 38941 3907 39009
rect 5061 38941 5095 39009
rect 3873 38907 3991 38941
rect 4025 38907 4059 38941
rect 4093 38907 4127 38941
rect 4161 38907 4195 38941
rect 4229 38907 4263 38941
rect 4297 38907 4331 38941
rect 4365 38907 4399 38941
rect 4433 38907 4467 38941
rect 4501 38907 4535 38941
rect 4569 38907 4603 38941
rect 4637 38907 4671 38941
rect 4705 38907 4739 38941
rect 4773 38907 4807 38941
rect 4841 38907 4875 38941
rect 4909 38907 4943 38941
rect 4977 38907 5095 38941
rect 199 38160 317 38194
rect 351 38160 385 38194
rect 419 38160 453 38194
rect 487 38160 521 38194
rect 555 38160 589 38194
rect 623 38160 657 38194
rect 691 38160 725 38194
rect 759 38160 793 38194
rect 827 38160 861 38194
rect 895 38160 929 38194
rect 963 38160 997 38194
rect 1031 38160 1065 38194
rect 1099 38160 1133 38194
rect 1167 38160 1201 38194
rect 1235 38160 1269 38194
rect 1303 38160 1421 38194
rect 199 38092 233 38160
rect 199 38024 233 38058
rect 1387 38092 1421 38160
rect 1387 38024 1421 38058
rect 199 37956 233 37990
rect 199 37888 233 37922
rect 199 37820 233 37854
rect 199 37752 233 37786
rect 1387 37956 1421 37990
rect 1387 37888 1421 37922
rect 1387 37820 1421 37854
rect 1387 37752 1421 37786
rect 199 37650 233 37718
rect 1387 37650 1421 37718
rect 199 37616 317 37650
rect 351 37616 385 37650
rect 419 37616 453 37650
rect 487 37616 521 37650
rect 555 37616 589 37650
rect 623 37616 657 37650
rect 691 37616 725 37650
rect 759 37616 793 37650
rect 827 37616 861 37650
rect 895 37616 929 37650
rect 963 37616 997 37650
rect 1031 37616 1065 37650
rect 1099 37616 1133 37650
rect 1167 37616 1201 37650
rect 1235 37616 1269 37650
rect 1303 37616 1421 37650
rect 2352 38164 2470 38198
rect 2504 38164 2538 38198
rect 2572 38164 2606 38198
rect 2640 38164 2674 38198
rect 2708 38164 2742 38198
rect 2776 38164 2810 38198
rect 2844 38164 2878 38198
rect 2912 38164 2946 38198
rect 2980 38164 3014 38198
rect 3048 38164 3082 38198
rect 3116 38164 3150 38198
rect 3184 38164 3218 38198
rect 3252 38164 3286 38198
rect 3320 38164 3354 38198
rect 3388 38164 3422 38198
rect 3456 38164 3574 38198
rect 2352 38096 2386 38164
rect 2352 38028 2386 38062
rect 3540 38096 3574 38164
rect 3540 38028 3574 38062
rect 2352 37960 2386 37994
rect 2352 37892 2386 37926
rect 2352 37824 2386 37858
rect 2352 37756 2386 37790
rect 3540 37960 3574 37994
rect 3540 37892 3574 37926
rect 3540 37824 3574 37858
rect 3540 37756 3574 37790
rect 2352 37654 2386 37722
rect 3540 37654 3574 37722
rect 2352 37620 2470 37654
rect 2504 37620 2538 37654
rect 2572 37620 2606 37654
rect 2640 37620 2674 37654
rect 2708 37620 2742 37654
rect 2776 37620 2810 37654
rect 2844 37620 2878 37654
rect 2912 37620 2946 37654
rect 2980 37620 3014 37654
rect 3048 37620 3082 37654
rect 3116 37620 3150 37654
rect 3184 37620 3218 37654
rect 3252 37620 3286 37654
rect 3320 37620 3354 37654
rect 3388 37620 3422 37654
rect 3456 37620 3574 37654
rect 3873 38164 3991 38198
rect 4025 38164 4059 38198
rect 4093 38164 4127 38198
rect 4161 38164 4195 38198
rect 4229 38164 4263 38198
rect 4297 38164 4331 38198
rect 4365 38164 4399 38198
rect 4433 38164 4467 38198
rect 4501 38164 4535 38198
rect 4569 38164 4603 38198
rect 4637 38164 4671 38198
rect 4705 38164 4739 38198
rect 4773 38164 4807 38198
rect 4841 38164 4875 38198
rect 4909 38164 4943 38198
rect 4977 38164 5095 38198
rect 3873 38096 3907 38164
rect 3873 38028 3907 38062
rect 5061 38096 5095 38164
rect 5061 38028 5095 38062
rect 3873 37960 3907 37994
rect 3873 37892 3907 37926
rect 3873 37824 3907 37858
rect 3873 37756 3907 37790
rect 5061 37960 5095 37994
rect 5061 37892 5095 37926
rect 5061 37824 5095 37858
rect 5061 37756 5095 37790
rect 3873 37654 3907 37722
rect 5061 37654 5095 37722
rect 3873 37620 3991 37654
rect 4025 37620 4059 37654
rect 4093 37620 4127 37654
rect 4161 37620 4195 37654
rect 4229 37620 4263 37654
rect 4297 37620 4331 37654
rect 4365 37620 4399 37654
rect 4433 37620 4467 37654
rect 4501 37620 4535 37654
rect 4569 37620 4603 37654
rect 4637 37620 4671 37654
rect 4705 37620 4739 37654
rect 4773 37620 4807 37654
rect 4841 37620 4875 37654
rect 4909 37620 4943 37654
rect 4977 37620 5095 37654
rect 199 36873 317 36907
rect 351 36873 385 36907
rect 419 36873 453 36907
rect 487 36873 521 36907
rect 555 36873 589 36907
rect 623 36873 657 36907
rect 691 36873 725 36907
rect 759 36873 793 36907
rect 827 36873 861 36907
rect 895 36873 929 36907
rect 963 36873 997 36907
rect 1031 36873 1065 36907
rect 1099 36873 1133 36907
rect 1167 36873 1201 36907
rect 1235 36873 1269 36907
rect 1303 36873 1421 36907
rect 199 36805 233 36873
rect 199 36737 233 36771
rect 1387 36805 1421 36873
rect 1387 36737 1421 36771
rect 199 36669 233 36703
rect 199 36601 233 36635
rect 199 36533 233 36567
rect 199 36465 233 36499
rect 1387 36669 1421 36703
rect 1387 36601 1421 36635
rect 1387 36533 1421 36567
rect 1387 36465 1421 36499
rect 199 36363 233 36431
rect 1387 36363 1421 36431
rect 199 36329 317 36363
rect 351 36329 385 36363
rect 419 36329 453 36363
rect 487 36329 521 36363
rect 555 36329 589 36363
rect 623 36329 657 36363
rect 691 36329 725 36363
rect 759 36329 793 36363
rect 827 36329 861 36363
rect 895 36329 929 36363
rect 963 36329 997 36363
rect 1031 36329 1065 36363
rect 1099 36329 1133 36363
rect 1167 36329 1201 36363
rect 1235 36329 1269 36363
rect 1303 36329 1421 36363
rect 2352 36877 2470 36911
rect 2504 36877 2538 36911
rect 2572 36877 2606 36911
rect 2640 36877 2674 36911
rect 2708 36877 2742 36911
rect 2776 36877 2810 36911
rect 2844 36877 2878 36911
rect 2912 36877 2946 36911
rect 2980 36877 3014 36911
rect 3048 36877 3082 36911
rect 3116 36877 3150 36911
rect 3184 36877 3218 36911
rect 3252 36877 3286 36911
rect 3320 36877 3354 36911
rect 3388 36877 3422 36911
rect 3456 36877 3574 36911
rect 2352 36809 2386 36877
rect 2352 36741 2386 36775
rect 3540 36809 3574 36877
rect 3540 36741 3574 36775
rect 2352 36673 2386 36707
rect 2352 36605 2386 36639
rect 2352 36537 2386 36571
rect 2352 36469 2386 36503
rect 3540 36673 3574 36707
rect 3540 36605 3574 36639
rect 3540 36537 3574 36571
rect 3540 36469 3574 36503
rect 2352 36367 2386 36435
rect 3540 36367 3574 36435
rect 2352 36333 2470 36367
rect 2504 36333 2538 36367
rect 2572 36333 2606 36367
rect 2640 36333 2674 36367
rect 2708 36333 2742 36367
rect 2776 36333 2810 36367
rect 2844 36333 2878 36367
rect 2912 36333 2946 36367
rect 2980 36333 3014 36367
rect 3048 36333 3082 36367
rect 3116 36333 3150 36367
rect 3184 36333 3218 36367
rect 3252 36333 3286 36367
rect 3320 36333 3354 36367
rect 3388 36333 3422 36367
rect 3456 36333 3574 36367
rect 3873 36877 3991 36911
rect 4025 36877 4059 36911
rect 4093 36877 4127 36911
rect 4161 36877 4195 36911
rect 4229 36877 4263 36911
rect 4297 36877 4331 36911
rect 4365 36877 4399 36911
rect 4433 36877 4467 36911
rect 4501 36877 4535 36911
rect 4569 36877 4603 36911
rect 4637 36877 4671 36911
rect 4705 36877 4739 36911
rect 4773 36877 4807 36911
rect 4841 36877 4875 36911
rect 4909 36877 4943 36911
rect 4977 36877 5095 36911
rect 3873 36809 3907 36877
rect 3873 36741 3907 36775
rect 5061 36809 5095 36877
rect 5061 36741 5095 36775
rect 3873 36673 3907 36707
rect 3873 36605 3907 36639
rect 3873 36537 3907 36571
rect 3873 36469 3907 36503
rect 5061 36673 5095 36707
rect 5061 36605 5095 36639
rect 5061 36537 5095 36571
rect 5061 36469 5095 36503
rect 3873 36367 3907 36435
rect 5061 36367 5095 36435
rect 3873 36333 3991 36367
rect 4025 36333 4059 36367
rect 4093 36333 4127 36367
rect 4161 36333 4195 36367
rect 4229 36333 4263 36367
rect 4297 36333 4331 36367
rect 4365 36333 4399 36367
rect 4433 36333 4467 36367
rect 4501 36333 4535 36367
rect 4569 36333 4603 36367
rect 4637 36333 4671 36367
rect 4705 36333 4739 36367
rect 4773 36333 4807 36367
rect 4841 36333 4875 36367
rect 4909 36333 4943 36367
rect 4977 36333 5095 36367
rect 199 35586 317 35620
rect 351 35586 385 35620
rect 419 35586 453 35620
rect 487 35586 521 35620
rect 555 35586 589 35620
rect 623 35586 657 35620
rect 691 35586 725 35620
rect 759 35586 793 35620
rect 827 35586 861 35620
rect 895 35586 929 35620
rect 963 35586 997 35620
rect 1031 35586 1065 35620
rect 1099 35586 1133 35620
rect 1167 35586 1201 35620
rect 1235 35586 1269 35620
rect 1303 35586 1421 35620
rect 199 35518 233 35586
rect 199 35450 233 35484
rect 1387 35518 1421 35586
rect 1387 35450 1421 35484
rect 199 35382 233 35416
rect 199 35314 233 35348
rect 199 35246 233 35280
rect 199 35178 233 35212
rect 1387 35382 1421 35416
rect 1387 35314 1421 35348
rect 1387 35246 1421 35280
rect 1387 35178 1421 35212
rect 199 35076 233 35144
rect 1387 35076 1421 35144
rect 199 35042 317 35076
rect 351 35042 385 35076
rect 419 35042 453 35076
rect 487 35042 521 35076
rect 555 35042 589 35076
rect 623 35042 657 35076
rect 691 35042 725 35076
rect 759 35042 793 35076
rect 827 35042 861 35076
rect 895 35042 929 35076
rect 963 35042 997 35076
rect 1031 35042 1065 35076
rect 1099 35042 1133 35076
rect 1167 35042 1201 35076
rect 1235 35042 1269 35076
rect 1303 35042 1421 35076
rect 2352 35590 2470 35624
rect 2504 35590 2538 35624
rect 2572 35590 2606 35624
rect 2640 35590 2674 35624
rect 2708 35590 2742 35624
rect 2776 35590 2810 35624
rect 2844 35590 2878 35624
rect 2912 35590 2946 35624
rect 2980 35590 3014 35624
rect 3048 35590 3082 35624
rect 3116 35590 3150 35624
rect 3184 35590 3218 35624
rect 3252 35590 3286 35624
rect 3320 35590 3354 35624
rect 3388 35590 3422 35624
rect 3456 35590 3574 35624
rect 2352 35522 2386 35590
rect 2352 35454 2386 35488
rect 3540 35522 3574 35590
rect 3540 35454 3574 35488
rect 2352 35386 2386 35420
rect 2352 35318 2386 35352
rect 2352 35250 2386 35284
rect 2352 35182 2386 35216
rect 3540 35386 3574 35420
rect 3540 35318 3574 35352
rect 3540 35250 3574 35284
rect 3540 35182 3574 35216
rect 2352 35080 2386 35148
rect 3540 35080 3574 35148
rect 2352 35046 2470 35080
rect 2504 35046 2538 35080
rect 2572 35046 2606 35080
rect 2640 35046 2674 35080
rect 2708 35046 2742 35080
rect 2776 35046 2810 35080
rect 2844 35046 2878 35080
rect 2912 35046 2946 35080
rect 2980 35046 3014 35080
rect 3048 35046 3082 35080
rect 3116 35046 3150 35080
rect 3184 35046 3218 35080
rect 3252 35046 3286 35080
rect 3320 35046 3354 35080
rect 3388 35046 3422 35080
rect 3456 35046 3574 35080
rect 3873 35590 3991 35624
rect 4025 35590 4059 35624
rect 4093 35590 4127 35624
rect 4161 35590 4195 35624
rect 4229 35590 4263 35624
rect 4297 35590 4331 35624
rect 4365 35590 4399 35624
rect 4433 35590 4467 35624
rect 4501 35590 4535 35624
rect 4569 35590 4603 35624
rect 4637 35590 4671 35624
rect 4705 35590 4739 35624
rect 4773 35590 4807 35624
rect 4841 35590 4875 35624
rect 4909 35590 4943 35624
rect 4977 35590 5095 35624
rect 3873 35522 3907 35590
rect 3873 35454 3907 35488
rect 5061 35522 5095 35590
rect 5061 35454 5095 35488
rect 3873 35386 3907 35420
rect 3873 35318 3907 35352
rect 3873 35250 3907 35284
rect 3873 35182 3907 35216
rect 5061 35386 5095 35420
rect 5061 35318 5095 35352
rect 5061 35250 5095 35284
rect 5061 35182 5095 35216
rect 3873 35080 3907 35148
rect 5061 35080 5095 35148
rect 3873 35046 3991 35080
rect 4025 35046 4059 35080
rect 4093 35046 4127 35080
rect 4161 35046 4195 35080
rect 4229 35046 4263 35080
rect 4297 35046 4331 35080
rect 4365 35046 4399 35080
rect 4433 35046 4467 35080
rect 4501 35046 4535 35080
rect 4569 35046 4603 35080
rect 4637 35046 4671 35080
rect 4705 35046 4739 35080
rect 4773 35046 4807 35080
rect 4841 35046 4875 35080
rect 4909 35046 4943 35080
rect 4977 35046 5095 35080
rect 199 34299 317 34333
rect 351 34299 385 34333
rect 419 34299 453 34333
rect 487 34299 521 34333
rect 555 34299 589 34333
rect 623 34299 657 34333
rect 691 34299 725 34333
rect 759 34299 793 34333
rect 827 34299 861 34333
rect 895 34299 929 34333
rect 963 34299 997 34333
rect 1031 34299 1065 34333
rect 1099 34299 1133 34333
rect 1167 34299 1201 34333
rect 1235 34299 1269 34333
rect 1303 34299 1421 34333
rect 199 34231 233 34299
rect 199 34163 233 34197
rect 1387 34231 1421 34299
rect 1387 34163 1421 34197
rect 199 34095 233 34129
rect 199 34027 233 34061
rect 199 33959 233 33993
rect 199 33891 233 33925
rect 1387 34095 1421 34129
rect 1387 34027 1421 34061
rect 1387 33959 1421 33993
rect 1387 33891 1421 33925
rect 199 33789 233 33857
rect 1387 33789 1421 33857
rect 199 33755 317 33789
rect 351 33755 385 33789
rect 419 33755 453 33789
rect 487 33755 521 33789
rect 555 33755 589 33789
rect 623 33755 657 33789
rect 691 33755 725 33789
rect 759 33755 793 33789
rect 827 33755 861 33789
rect 895 33755 929 33789
rect 963 33755 997 33789
rect 1031 33755 1065 33789
rect 1099 33755 1133 33789
rect 1167 33755 1201 33789
rect 1235 33755 1269 33789
rect 1303 33755 1421 33789
rect 2352 34303 2470 34337
rect 2504 34303 2538 34337
rect 2572 34303 2606 34337
rect 2640 34303 2674 34337
rect 2708 34303 2742 34337
rect 2776 34303 2810 34337
rect 2844 34303 2878 34337
rect 2912 34303 2946 34337
rect 2980 34303 3014 34337
rect 3048 34303 3082 34337
rect 3116 34303 3150 34337
rect 3184 34303 3218 34337
rect 3252 34303 3286 34337
rect 3320 34303 3354 34337
rect 3388 34303 3422 34337
rect 3456 34303 3574 34337
rect 2352 34235 2386 34303
rect 2352 34167 2386 34201
rect 3540 34235 3574 34303
rect 3540 34167 3574 34201
rect 2352 34099 2386 34133
rect 2352 34031 2386 34065
rect 2352 33963 2386 33997
rect 2352 33895 2386 33929
rect 3540 34099 3574 34133
rect 3540 34031 3574 34065
rect 3540 33963 3574 33997
rect 3540 33895 3574 33929
rect 2352 33793 2386 33861
rect 3540 33793 3574 33861
rect 2352 33759 2470 33793
rect 2504 33759 2538 33793
rect 2572 33759 2606 33793
rect 2640 33759 2674 33793
rect 2708 33759 2742 33793
rect 2776 33759 2810 33793
rect 2844 33759 2878 33793
rect 2912 33759 2946 33793
rect 2980 33759 3014 33793
rect 3048 33759 3082 33793
rect 3116 33759 3150 33793
rect 3184 33759 3218 33793
rect 3252 33759 3286 33793
rect 3320 33759 3354 33793
rect 3388 33759 3422 33793
rect 3456 33759 3574 33793
rect 3873 34303 3991 34337
rect 4025 34303 4059 34337
rect 4093 34303 4127 34337
rect 4161 34303 4195 34337
rect 4229 34303 4263 34337
rect 4297 34303 4331 34337
rect 4365 34303 4399 34337
rect 4433 34303 4467 34337
rect 4501 34303 4535 34337
rect 4569 34303 4603 34337
rect 4637 34303 4671 34337
rect 4705 34303 4739 34337
rect 4773 34303 4807 34337
rect 4841 34303 4875 34337
rect 4909 34303 4943 34337
rect 4977 34303 5095 34337
rect 3873 34235 3907 34303
rect 3873 34167 3907 34201
rect 5061 34235 5095 34303
rect 5061 34167 5095 34201
rect 3873 34099 3907 34133
rect 3873 34031 3907 34065
rect 3873 33963 3907 33997
rect 3873 33895 3907 33929
rect 5061 34099 5095 34133
rect 5061 34031 5095 34065
rect 5061 33963 5095 33997
rect 5061 33895 5095 33929
rect 3873 33793 3907 33861
rect 5061 33793 5095 33861
rect 3873 33759 3991 33793
rect 4025 33759 4059 33793
rect 4093 33759 4127 33793
rect 4161 33759 4195 33793
rect 4229 33759 4263 33793
rect 4297 33759 4331 33793
rect 4365 33759 4399 33793
rect 4433 33759 4467 33793
rect 4501 33759 4535 33793
rect 4569 33759 4603 33793
rect 4637 33759 4671 33793
rect 4705 33759 4739 33793
rect 4773 33759 4807 33793
rect 4841 33759 4875 33793
rect 4909 33759 4943 33793
rect 4977 33759 5095 33793
rect 199 33012 317 33046
rect 351 33012 385 33046
rect 419 33012 453 33046
rect 487 33012 521 33046
rect 555 33012 589 33046
rect 623 33012 657 33046
rect 691 33012 725 33046
rect 759 33012 793 33046
rect 827 33012 861 33046
rect 895 33012 929 33046
rect 963 33012 997 33046
rect 1031 33012 1065 33046
rect 1099 33012 1133 33046
rect 1167 33012 1201 33046
rect 1235 33012 1269 33046
rect 1303 33012 1421 33046
rect 199 32944 233 33012
rect 199 32876 233 32910
rect 1387 32944 1421 33012
rect 1387 32876 1421 32910
rect 199 32808 233 32842
rect 199 32740 233 32774
rect 199 32672 233 32706
rect 199 32604 233 32638
rect 1387 32808 1421 32842
rect 1387 32740 1421 32774
rect 1387 32672 1421 32706
rect 1387 32604 1421 32638
rect 199 32502 233 32570
rect 1387 32502 1421 32570
rect 199 32468 317 32502
rect 351 32468 385 32502
rect 419 32468 453 32502
rect 487 32468 521 32502
rect 555 32468 589 32502
rect 623 32468 657 32502
rect 691 32468 725 32502
rect 759 32468 793 32502
rect 827 32468 861 32502
rect 895 32468 929 32502
rect 963 32468 997 32502
rect 1031 32468 1065 32502
rect 1099 32468 1133 32502
rect 1167 32468 1201 32502
rect 1235 32468 1269 32502
rect 1303 32468 1421 32502
rect 2352 33016 2470 33050
rect 2504 33016 2538 33050
rect 2572 33016 2606 33050
rect 2640 33016 2674 33050
rect 2708 33016 2742 33050
rect 2776 33016 2810 33050
rect 2844 33016 2878 33050
rect 2912 33016 2946 33050
rect 2980 33016 3014 33050
rect 3048 33016 3082 33050
rect 3116 33016 3150 33050
rect 3184 33016 3218 33050
rect 3252 33016 3286 33050
rect 3320 33016 3354 33050
rect 3388 33016 3422 33050
rect 3456 33016 3574 33050
rect 2352 32948 2386 33016
rect 2352 32880 2386 32914
rect 3540 32948 3574 33016
rect 3540 32880 3574 32914
rect 2352 32812 2386 32846
rect 2352 32744 2386 32778
rect 2352 32676 2386 32710
rect 2352 32608 2386 32642
rect 3540 32812 3574 32846
rect 3540 32744 3574 32778
rect 3540 32676 3574 32710
rect 3540 32608 3574 32642
rect 2352 32506 2386 32574
rect 3540 32506 3574 32574
rect 2352 32472 2470 32506
rect 2504 32472 2538 32506
rect 2572 32472 2606 32506
rect 2640 32472 2674 32506
rect 2708 32472 2742 32506
rect 2776 32472 2810 32506
rect 2844 32472 2878 32506
rect 2912 32472 2946 32506
rect 2980 32472 3014 32506
rect 3048 32472 3082 32506
rect 3116 32472 3150 32506
rect 3184 32472 3218 32506
rect 3252 32472 3286 32506
rect 3320 32472 3354 32506
rect 3388 32472 3422 32506
rect 3456 32472 3574 32506
rect 3873 33016 3991 33050
rect 4025 33016 4059 33050
rect 4093 33016 4127 33050
rect 4161 33016 4195 33050
rect 4229 33016 4263 33050
rect 4297 33016 4331 33050
rect 4365 33016 4399 33050
rect 4433 33016 4467 33050
rect 4501 33016 4535 33050
rect 4569 33016 4603 33050
rect 4637 33016 4671 33050
rect 4705 33016 4739 33050
rect 4773 33016 4807 33050
rect 4841 33016 4875 33050
rect 4909 33016 4943 33050
rect 4977 33016 5095 33050
rect 3873 32948 3907 33016
rect 3873 32880 3907 32914
rect 5061 32948 5095 33016
rect 5061 32880 5095 32914
rect 3873 32812 3907 32846
rect 3873 32744 3907 32778
rect 3873 32676 3907 32710
rect 3873 32608 3907 32642
rect 5061 32812 5095 32846
rect 5061 32744 5095 32778
rect 5061 32676 5095 32710
rect 5061 32608 5095 32642
rect 3873 32506 3907 32574
rect 5061 32506 5095 32574
rect 3873 32472 3991 32506
rect 4025 32472 4059 32506
rect 4093 32472 4127 32506
rect 4161 32472 4195 32506
rect 4229 32472 4263 32506
rect 4297 32472 4331 32506
rect 4365 32472 4399 32506
rect 4433 32472 4467 32506
rect 4501 32472 4535 32506
rect 4569 32472 4603 32506
rect 4637 32472 4671 32506
rect 4705 32472 4739 32506
rect 4773 32472 4807 32506
rect 4841 32472 4875 32506
rect 4909 32472 4943 32506
rect 4977 32472 5095 32506
rect 199 31725 317 31759
rect 351 31725 385 31759
rect 419 31725 453 31759
rect 487 31725 521 31759
rect 555 31725 589 31759
rect 623 31725 657 31759
rect 691 31725 725 31759
rect 759 31725 793 31759
rect 827 31725 861 31759
rect 895 31725 929 31759
rect 963 31725 997 31759
rect 1031 31725 1065 31759
rect 1099 31725 1133 31759
rect 1167 31725 1201 31759
rect 1235 31725 1269 31759
rect 1303 31725 1421 31759
rect 199 31657 233 31725
rect 199 31589 233 31623
rect 1387 31657 1421 31725
rect 1387 31589 1421 31623
rect 199 31521 233 31555
rect 199 31453 233 31487
rect 199 31385 233 31419
rect 199 31317 233 31351
rect 1387 31521 1421 31555
rect 1387 31453 1421 31487
rect 1387 31385 1421 31419
rect 1387 31317 1421 31351
rect 199 31215 233 31283
rect 1387 31215 1421 31283
rect 199 31181 317 31215
rect 351 31181 385 31215
rect 419 31181 453 31215
rect 487 31181 521 31215
rect 555 31181 589 31215
rect 623 31181 657 31215
rect 691 31181 725 31215
rect 759 31181 793 31215
rect 827 31181 861 31215
rect 895 31181 929 31215
rect 963 31181 997 31215
rect 1031 31181 1065 31215
rect 1099 31181 1133 31215
rect 1167 31181 1201 31215
rect 1235 31181 1269 31215
rect 1303 31181 1421 31215
rect 2352 31729 2470 31763
rect 2504 31729 2538 31763
rect 2572 31729 2606 31763
rect 2640 31729 2674 31763
rect 2708 31729 2742 31763
rect 2776 31729 2810 31763
rect 2844 31729 2878 31763
rect 2912 31729 2946 31763
rect 2980 31729 3014 31763
rect 3048 31729 3082 31763
rect 3116 31729 3150 31763
rect 3184 31729 3218 31763
rect 3252 31729 3286 31763
rect 3320 31729 3354 31763
rect 3388 31729 3422 31763
rect 3456 31729 3574 31763
rect 2352 31661 2386 31729
rect 2352 31593 2386 31627
rect 3540 31661 3574 31729
rect 3540 31593 3574 31627
rect 2352 31525 2386 31559
rect 2352 31457 2386 31491
rect 2352 31389 2386 31423
rect 2352 31321 2386 31355
rect 3540 31525 3574 31559
rect 3540 31457 3574 31491
rect 3540 31389 3574 31423
rect 3540 31321 3574 31355
rect 2352 31219 2386 31287
rect 3540 31219 3574 31287
rect 2352 31185 2470 31219
rect 2504 31185 2538 31219
rect 2572 31185 2606 31219
rect 2640 31185 2674 31219
rect 2708 31185 2742 31219
rect 2776 31185 2810 31219
rect 2844 31185 2878 31219
rect 2912 31185 2946 31219
rect 2980 31185 3014 31219
rect 3048 31185 3082 31219
rect 3116 31185 3150 31219
rect 3184 31185 3218 31219
rect 3252 31185 3286 31219
rect 3320 31185 3354 31219
rect 3388 31185 3422 31219
rect 3456 31185 3574 31219
rect 3873 31729 3991 31763
rect 4025 31729 4059 31763
rect 4093 31729 4127 31763
rect 4161 31729 4195 31763
rect 4229 31729 4263 31763
rect 4297 31729 4331 31763
rect 4365 31729 4399 31763
rect 4433 31729 4467 31763
rect 4501 31729 4535 31763
rect 4569 31729 4603 31763
rect 4637 31729 4671 31763
rect 4705 31729 4739 31763
rect 4773 31729 4807 31763
rect 4841 31729 4875 31763
rect 4909 31729 4943 31763
rect 4977 31729 5095 31763
rect 3873 31661 3907 31729
rect 3873 31593 3907 31627
rect 5061 31661 5095 31729
rect 5061 31593 5095 31627
rect 3873 31525 3907 31559
rect 3873 31457 3907 31491
rect 3873 31389 3907 31423
rect 3873 31321 3907 31355
rect 5061 31525 5095 31559
rect 5061 31457 5095 31491
rect 5061 31389 5095 31423
rect 5061 31321 5095 31355
rect 3873 31219 3907 31287
rect 5061 31219 5095 31287
rect 3873 31185 3991 31219
rect 4025 31185 4059 31219
rect 4093 31185 4127 31219
rect 4161 31185 4195 31219
rect 4229 31185 4263 31219
rect 4297 31185 4331 31219
rect 4365 31185 4399 31219
rect 4433 31185 4467 31219
rect 4501 31185 4535 31219
rect 4569 31185 4603 31219
rect 4637 31185 4671 31219
rect 4705 31185 4739 31219
rect 4773 31185 4807 31219
rect 4841 31185 4875 31219
rect 4909 31185 4943 31219
rect 4977 31185 5095 31219
rect 199 30438 317 30472
rect 351 30438 385 30472
rect 419 30438 453 30472
rect 487 30438 521 30472
rect 555 30438 589 30472
rect 623 30438 657 30472
rect 691 30438 725 30472
rect 759 30438 793 30472
rect 827 30438 861 30472
rect 895 30438 929 30472
rect 963 30438 997 30472
rect 1031 30438 1065 30472
rect 1099 30438 1133 30472
rect 1167 30438 1201 30472
rect 1235 30438 1269 30472
rect 1303 30438 1421 30472
rect 199 30370 233 30438
rect 199 30302 233 30336
rect 1387 30370 1421 30438
rect 1387 30302 1421 30336
rect 199 30234 233 30268
rect 199 30166 233 30200
rect 199 30098 233 30132
rect 199 30030 233 30064
rect 1387 30234 1421 30268
rect 1387 30166 1421 30200
rect 1387 30098 1421 30132
rect 1387 30030 1421 30064
rect 199 29928 233 29996
rect 1387 29928 1421 29996
rect 199 29894 317 29928
rect 351 29894 385 29928
rect 419 29894 453 29928
rect 487 29894 521 29928
rect 555 29894 589 29928
rect 623 29894 657 29928
rect 691 29894 725 29928
rect 759 29894 793 29928
rect 827 29894 861 29928
rect 895 29894 929 29928
rect 963 29894 997 29928
rect 1031 29894 1065 29928
rect 1099 29894 1133 29928
rect 1167 29894 1201 29928
rect 1235 29894 1269 29928
rect 1303 29894 1421 29928
rect 2352 30442 2470 30476
rect 2504 30442 2538 30476
rect 2572 30442 2606 30476
rect 2640 30442 2674 30476
rect 2708 30442 2742 30476
rect 2776 30442 2810 30476
rect 2844 30442 2878 30476
rect 2912 30442 2946 30476
rect 2980 30442 3014 30476
rect 3048 30442 3082 30476
rect 3116 30442 3150 30476
rect 3184 30442 3218 30476
rect 3252 30442 3286 30476
rect 3320 30442 3354 30476
rect 3388 30442 3422 30476
rect 3456 30442 3574 30476
rect 2352 30374 2386 30442
rect 2352 30306 2386 30340
rect 3540 30374 3574 30442
rect 3540 30306 3574 30340
rect 2352 30238 2386 30272
rect 2352 30170 2386 30204
rect 2352 30102 2386 30136
rect 2352 30034 2386 30068
rect 3540 30238 3574 30272
rect 3540 30170 3574 30204
rect 3540 30102 3574 30136
rect 3540 30034 3574 30068
rect 2352 29932 2386 30000
rect 3540 29932 3574 30000
rect 2352 29898 2470 29932
rect 2504 29898 2538 29932
rect 2572 29898 2606 29932
rect 2640 29898 2674 29932
rect 2708 29898 2742 29932
rect 2776 29898 2810 29932
rect 2844 29898 2878 29932
rect 2912 29898 2946 29932
rect 2980 29898 3014 29932
rect 3048 29898 3082 29932
rect 3116 29898 3150 29932
rect 3184 29898 3218 29932
rect 3252 29898 3286 29932
rect 3320 29898 3354 29932
rect 3388 29898 3422 29932
rect 3456 29898 3574 29932
rect 3873 30442 3991 30476
rect 4025 30442 4059 30476
rect 4093 30442 4127 30476
rect 4161 30442 4195 30476
rect 4229 30442 4263 30476
rect 4297 30442 4331 30476
rect 4365 30442 4399 30476
rect 4433 30442 4467 30476
rect 4501 30442 4535 30476
rect 4569 30442 4603 30476
rect 4637 30442 4671 30476
rect 4705 30442 4739 30476
rect 4773 30442 4807 30476
rect 4841 30442 4875 30476
rect 4909 30442 4943 30476
rect 4977 30442 5095 30476
rect 3873 30374 3907 30442
rect 3873 30306 3907 30340
rect 5061 30374 5095 30442
rect 5061 30306 5095 30340
rect 3873 30238 3907 30272
rect 3873 30170 3907 30204
rect 3873 30102 3907 30136
rect 3873 30034 3907 30068
rect 5061 30238 5095 30272
rect 5061 30170 5095 30204
rect 5061 30102 5095 30136
rect 5061 30034 5095 30068
rect 3873 29932 3907 30000
rect 5061 29932 5095 30000
rect 3873 29898 3991 29932
rect 4025 29898 4059 29932
rect 4093 29898 4127 29932
rect 4161 29898 4195 29932
rect 4229 29898 4263 29932
rect 4297 29898 4331 29932
rect 4365 29898 4399 29932
rect 4433 29898 4467 29932
rect 4501 29898 4535 29932
rect 4569 29898 4603 29932
rect 4637 29898 4671 29932
rect 4705 29898 4739 29932
rect 4773 29898 4807 29932
rect 4841 29898 4875 29932
rect 4909 29898 4943 29932
rect 4977 29898 5095 29932
rect 199 29151 317 29185
rect 351 29151 385 29185
rect 419 29151 453 29185
rect 487 29151 521 29185
rect 555 29151 589 29185
rect 623 29151 657 29185
rect 691 29151 725 29185
rect 759 29151 793 29185
rect 827 29151 861 29185
rect 895 29151 929 29185
rect 963 29151 997 29185
rect 1031 29151 1065 29185
rect 1099 29151 1133 29185
rect 1167 29151 1201 29185
rect 1235 29151 1269 29185
rect 1303 29151 1421 29185
rect 199 29083 233 29151
rect 199 29015 233 29049
rect 1387 29083 1421 29151
rect 1387 29015 1421 29049
rect 199 28947 233 28981
rect 199 28879 233 28913
rect 199 28811 233 28845
rect 199 28743 233 28777
rect 1387 28947 1421 28981
rect 1387 28879 1421 28913
rect 1387 28811 1421 28845
rect 1387 28743 1421 28777
rect 199 28641 233 28709
rect 1387 28641 1421 28709
rect 199 28607 317 28641
rect 351 28607 385 28641
rect 419 28607 453 28641
rect 487 28607 521 28641
rect 555 28607 589 28641
rect 623 28607 657 28641
rect 691 28607 725 28641
rect 759 28607 793 28641
rect 827 28607 861 28641
rect 895 28607 929 28641
rect 963 28607 997 28641
rect 1031 28607 1065 28641
rect 1099 28607 1133 28641
rect 1167 28607 1201 28641
rect 1235 28607 1269 28641
rect 1303 28607 1421 28641
rect 2352 29155 2470 29189
rect 2504 29155 2538 29189
rect 2572 29155 2606 29189
rect 2640 29155 2674 29189
rect 2708 29155 2742 29189
rect 2776 29155 2810 29189
rect 2844 29155 2878 29189
rect 2912 29155 2946 29189
rect 2980 29155 3014 29189
rect 3048 29155 3082 29189
rect 3116 29155 3150 29189
rect 3184 29155 3218 29189
rect 3252 29155 3286 29189
rect 3320 29155 3354 29189
rect 3388 29155 3422 29189
rect 3456 29155 3574 29189
rect 2352 29087 2386 29155
rect 2352 29019 2386 29053
rect 3540 29087 3574 29155
rect 3540 29019 3574 29053
rect 2352 28951 2386 28985
rect 2352 28883 2386 28917
rect 2352 28815 2386 28849
rect 2352 28747 2386 28781
rect 3540 28951 3574 28985
rect 3540 28883 3574 28917
rect 3540 28815 3574 28849
rect 3540 28747 3574 28781
rect 2352 28645 2386 28713
rect 3540 28645 3574 28713
rect 2352 28611 2470 28645
rect 2504 28611 2538 28645
rect 2572 28611 2606 28645
rect 2640 28611 2674 28645
rect 2708 28611 2742 28645
rect 2776 28611 2810 28645
rect 2844 28611 2878 28645
rect 2912 28611 2946 28645
rect 2980 28611 3014 28645
rect 3048 28611 3082 28645
rect 3116 28611 3150 28645
rect 3184 28611 3218 28645
rect 3252 28611 3286 28645
rect 3320 28611 3354 28645
rect 3388 28611 3422 28645
rect 3456 28611 3574 28645
rect 3873 29155 3991 29189
rect 4025 29155 4059 29189
rect 4093 29155 4127 29189
rect 4161 29155 4195 29189
rect 4229 29155 4263 29189
rect 4297 29155 4331 29189
rect 4365 29155 4399 29189
rect 4433 29155 4467 29189
rect 4501 29155 4535 29189
rect 4569 29155 4603 29189
rect 4637 29155 4671 29189
rect 4705 29155 4739 29189
rect 4773 29155 4807 29189
rect 4841 29155 4875 29189
rect 4909 29155 4943 29189
rect 4977 29155 5095 29189
rect 3873 29087 3907 29155
rect 3873 29019 3907 29053
rect 5061 29087 5095 29155
rect 5061 29019 5095 29053
rect 3873 28951 3907 28985
rect 3873 28883 3907 28917
rect 3873 28815 3907 28849
rect 3873 28747 3907 28781
rect 5061 28951 5095 28985
rect 5061 28883 5095 28917
rect 5061 28815 5095 28849
rect 5061 28747 5095 28781
rect 3873 28645 3907 28713
rect 5061 28645 5095 28713
rect 3873 28611 3991 28645
rect 4025 28611 4059 28645
rect 4093 28611 4127 28645
rect 4161 28611 4195 28645
rect 4229 28611 4263 28645
rect 4297 28611 4331 28645
rect 4365 28611 4399 28645
rect 4433 28611 4467 28645
rect 4501 28611 4535 28645
rect 4569 28611 4603 28645
rect 4637 28611 4671 28645
rect 4705 28611 4739 28645
rect 4773 28611 4807 28645
rect 4841 28611 4875 28645
rect 4909 28611 4943 28645
rect 4977 28611 5095 28645
rect 199 27864 317 27898
rect 351 27864 385 27898
rect 419 27864 453 27898
rect 487 27864 521 27898
rect 555 27864 589 27898
rect 623 27864 657 27898
rect 691 27864 725 27898
rect 759 27864 793 27898
rect 827 27864 861 27898
rect 895 27864 929 27898
rect 963 27864 997 27898
rect 1031 27864 1065 27898
rect 1099 27864 1133 27898
rect 1167 27864 1201 27898
rect 1235 27864 1269 27898
rect 1303 27864 1421 27898
rect 199 27796 233 27864
rect 199 27728 233 27762
rect 1387 27796 1421 27864
rect 1387 27728 1421 27762
rect 199 27660 233 27694
rect 199 27592 233 27626
rect 199 27524 233 27558
rect 199 27456 233 27490
rect 1387 27660 1421 27694
rect 1387 27592 1421 27626
rect 1387 27524 1421 27558
rect 1387 27456 1421 27490
rect 199 27354 233 27422
rect 1387 27354 1421 27422
rect 199 27320 317 27354
rect 351 27320 385 27354
rect 419 27320 453 27354
rect 487 27320 521 27354
rect 555 27320 589 27354
rect 623 27320 657 27354
rect 691 27320 725 27354
rect 759 27320 793 27354
rect 827 27320 861 27354
rect 895 27320 929 27354
rect 963 27320 997 27354
rect 1031 27320 1065 27354
rect 1099 27320 1133 27354
rect 1167 27320 1201 27354
rect 1235 27320 1269 27354
rect 1303 27320 1421 27354
rect 2352 27868 2470 27902
rect 2504 27868 2538 27902
rect 2572 27868 2606 27902
rect 2640 27868 2674 27902
rect 2708 27868 2742 27902
rect 2776 27868 2810 27902
rect 2844 27868 2878 27902
rect 2912 27868 2946 27902
rect 2980 27868 3014 27902
rect 3048 27868 3082 27902
rect 3116 27868 3150 27902
rect 3184 27868 3218 27902
rect 3252 27868 3286 27902
rect 3320 27868 3354 27902
rect 3388 27868 3422 27902
rect 3456 27868 3574 27902
rect 2352 27800 2386 27868
rect 2352 27732 2386 27766
rect 3540 27800 3574 27868
rect 3540 27732 3574 27766
rect 2352 27664 2386 27698
rect 2352 27596 2386 27630
rect 2352 27528 2386 27562
rect 2352 27460 2386 27494
rect 3540 27664 3574 27698
rect 3540 27596 3574 27630
rect 3540 27528 3574 27562
rect 3540 27460 3574 27494
rect 2352 27358 2386 27426
rect 3540 27358 3574 27426
rect 2352 27324 2470 27358
rect 2504 27324 2538 27358
rect 2572 27324 2606 27358
rect 2640 27324 2674 27358
rect 2708 27324 2742 27358
rect 2776 27324 2810 27358
rect 2844 27324 2878 27358
rect 2912 27324 2946 27358
rect 2980 27324 3014 27358
rect 3048 27324 3082 27358
rect 3116 27324 3150 27358
rect 3184 27324 3218 27358
rect 3252 27324 3286 27358
rect 3320 27324 3354 27358
rect 3388 27324 3422 27358
rect 3456 27324 3574 27358
rect 3873 27868 3991 27902
rect 4025 27868 4059 27902
rect 4093 27868 4127 27902
rect 4161 27868 4195 27902
rect 4229 27868 4263 27902
rect 4297 27868 4331 27902
rect 4365 27868 4399 27902
rect 4433 27868 4467 27902
rect 4501 27868 4535 27902
rect 4569 27868 4603 27902
rect 4637 27868 4671 27902
rect 4705 27868 4739 27902
rect 4773 27868 4807 27902
rect 4841 27868 4875 27902
rect 4909 27868 4943 27902
rect 4977 27868 5095 27902
rect 3873 27800 3907 27868
rect 3873 27732 3907 27766
rect 5061 27800 5095 27868
rect 5061 27732 5095 27766
rect 3873 27664 3907 27698
rect 3873 27596 3907 27630
rect 3873 27528 3907 27562
rect 3873 27460 3907 27494
rect 5061 27664 5095 27698
rect 5061 27596 5095 27630
rect 5061 27528 5095 27562
rect 5061 27460 5095 27494
rect 3873 27358 3907 27426
rect 5061 27358 5095 27426
rect 3873 27324 3991 27358
rect 4025 27324 4059 27358
rect 4093 27324 4127 27358
rect 4161 27324 4195 27358
rect 4229 27324 4263 27358
rect 4297 27324 4331 27358
rect 4365 27324 4399 27358
rect 4433 27324 4467 27358
rect 4501 27324 4535 27358
rect 4569 27324 4603 27358
rect 4637 27324 4671 27358
rect 4705 27324 4739 27358
rect 4773 27324 4807 27358
rect 4841 27324 4875 27358
rect 4909 27324 4943 27358
rect 4977 27324 5095 27358
rect 199 26577 317 26611
rect 351 26577 385 26611
rect 419 26577 453 26611
rect 487 26577 521 26611
rect 555 26577 589 26611
rect 623 26577 657 26611
rect 691 26577 725 26611
rect 759 26577 793 26611
rect 827 26577 861 26611
rect 895 26577 929 26611
rect 963 26577 997 26611
rect 1031 26577 1065 26611
rect 1099 26577 1133 26611
rect 1167 26577 1201 26611
rect 1235 26577 1269 26611
rect 1303 26577 1421 26611
rect 199 26509 233 26577
rect 199 26441 233 26475
rect 1387 26509 1421 26577
rect 1387 26441 1421 26475
rect 199 26373 233 26407
rect 199 26305 233 26339
rect 199 26237 233 26271
rect 199 26169 233 26203
rect 1387 26373 1421 26407
rect 1387 26305 1421 26339
rect 1387 26237 1421 26271
rect 1387 26169 1421 26203
rect 199 26067 233 26135
rect 1387 26067 1421 26135
rect 199 26033 317 26067
rect 351 26033 385 26067
rect 419 26033 453 26067
rect 487 26033 521 26067
rect 555 26033 589 26067
rect 623 26033 657 26067
rect 691 26033 725 26067
rect 759 26033 793 26067
rect 827 26033 861 26067
rect 895 26033 929 26067
rect 963 26033 997 26067
rect 1031 26033 1065 26067
rect 1099 26033 1133 26067
rect 1167 26033 1201 26067
rect 1235 26033 1269 26067
rect 1303 26033 1421 26067
rect 2352 26581 2470 26615
rect 2504 26581 2538 26615
rect 2572 26581 2606 26615
rect 2640 26581 2674 26615
rect 2708 26581 2742 26615
rect 2776 26581 2810 26615
rect 2844 26581 2878 26615
rect 2912 26581 2946 26615
rect 2980 26581 3014 26615
rect 3048 26581 3082 26615
rect 3116 26581 3150 26615
rect 3184 26581 3218 26615
rect 3252 26581 3286 26615
rect 3320 26581 3354 26615
rect 3388 26581 3422 26615
rect 3456 26581 3574 26615
rect 2352 26513 2386 26581
rect 2352 26445 2386 26479
rect 3540 26513 3574 26581
rect 3540 26445 3574 26479
rect 2352 26377 2386 26411
rect 2352 26309 2386 26343
rect 2352 26241 2386 26275
rect 2352 26173 2386 26207
rect 3540 26377 3574 26411
rect 3540 26309 3574 26343
rect 3540 26241 3574 26275
rect 3540 26173 3574 26207
rect 2352 26071 2386 26139
rect 3540 26071 3574 26139
rect 2352 26037 2470 26071
rect 2504 26037 2538 26071
rect 2572 26037 2606 26071
rect 2640 26037 2674 26071
rect 2708 26037 2742 26071
rect 2776 26037 2810 26071
rect 2844 26037 2878 26071
rect 2912 26037 2946 26071
rect 2980 26037 3014 26071
rect 3048 26037 3082 26071
rect 3116 26037 3150 26071
rect 3184 26037 3218 26071
rect 3252 26037 3286 26071
rect 3320 26037 3354 26071
rect 3388 26037 3422 26071
rect 3456 26037 3574 26071
rect 3873 26581 3991 26615
rect 4025 26581 4059 26615
rect 4093 26581 4127 26615
rect 4161 26581 4195 26615
rect 4229 26581 4263 26615
rect 4297 26581 4331 26615
rect 4365 26581 4399 26615
rect 4433 26581 4467 26615
rect 4501 26581 4535 26615
rect 4569 26581 4603 26615
rect 4637 26581 4671 26615
rect 4705 26581 4739 26615
rect 4773 26581 4807 26615
rect 4841 26581 4875 26615
rect 4909 26581 4943 26615
rect 4977 26581 5095 26615
rect 3873 26513 3907 26581
rect 3873 26445 3907 26479
rect 5061 26513 5095 26581
rect 5061 26445 5095 26479
rect 3873 26377 3907 26411
rect 3873 26309 3907 26343
rect 3873 26241 3907 26275
rect 3873 26173 3907 26207
rect 5061 26377 5095 26411
rect 5061 26309 5095 26343
rect 5061 26241 5095 26275
rect 5061 26173 5095 26207
rect 3873 26071 3907 26139
rect 5061 26071 5095 26139
rect 3873 26037 3991 26071
rect 4025 26037 4059 26071
rect 4093 26037 4127 26071
rect 4161 26037 4195 26071
rect 4229 26037 4263 26071
rect 4297 26037 4331 26071
rect 4365 26037 4399 26071
rect 4433 26037 4467 26071
rect 4501 26037 4535 26071
rect 4569 26037 4603 26071
rect 4637 26037 4671 26071
rect 4705 26037 4739 26071
rect 4773 26037 4807 26071
rect 4841 26037 4875 26071
rect 4909 26037 4943 26071
rect 4977 26037 5095 26071
rect 199 25290 317 25324
rect 351 25290 385 25324
rect 419 25290 453 25324
rect 487 25290 521 25324
rect 555 25290 589 25324
rect 623 25290 657 25324
rect 691 25290 725 25324
rect 759 25290 793 25324
rect 827 25290 861 25324
rect 895 25290 929 25324
rect 963 25290 997 25324
rect 1031 25290 1065 25324
rect 1099 25290 1133 25324
rect 1167 25290 1201 25324
rect 1235 25290 1269 25324
rect 1303 25290 1421 25324
rect 199 25222 233 25290
rect 199 25154 233 25188
rect 1387 25222 1421 25290
rect 1387 25154 1421 25188
rect 199 25086 233 25120
rect 199 25018 233 25052
rect 199 24950 233 24984
rect 199 24882 233 24916
rect 1387 25086 1421 25120
rect 1387 25018 1421 25052
rect 1387 24950 1421 24984
rect 1387 24882 1421 24916
rect 199 24780 233 24848
rect 1387 24780 1421 24848
rect 199 24746 317 24780
rect 351 24746 385 24780
rect 419 24746 453 24780
rect 487 24746 521 24780
rect 555 24746 589 24780
rect 623 24746 657 24780
rect 691 24746 725 24780
rect 759 24746 793 24780
rect 827 24746 861 24780
rect 895 24746 929 24780
rect 963 24746 997 24780
rect 1031 24746 1065 24780
rect 1099 24746 1133 24780
rect 1167 24746 1201 24780
rect 1235 24746 1269 24780
rect 1303 24746 1421 24780
rect 2352 25294 2470 25328
rect 2504 25294 2538 25328
rect 2572 25294 2606 25328
rect 2640 25294 2674 25328
rect 2708 25294 2742 25328
rect 2776 25294 2810 25328
rect 2844 25294 2878 25328
rect 2912 25294 2946 25328
rect 2980 25294 3014 25328
rect 3048 25294 3082 25328
rect 3116 25294 3150 25328
rect 3184 25294 3218 25328
rect 3252 25294 3286 25328
rect 3320 25294 3354 25328
rect 3388 25294 3422 25328
rect 3456 25294 3574 25328
rect 2352 25226 2386 25294
rect 2352 25158 2386 25192
rect 3540 25226 3574 25294
rect 3540 25158 3574 25192
rect 2352 25090 2386 25124
rect 2352 25022 2386 25056
rect 2352 24954 2386 24988
rect 2352 24886 2386 24920
rect 3540 25090 3574 25124
rect 3540 25022 3574 25056
rect 3540 24954 3574 24988
rect 3540 24886 3574 24920
rect 2352 24784 2386 24852
rect 3540 24784 3574 24852
rect 2352 24750 2470 24784
rect 2504 24750 2538 24784
rect 2572 24750 2606 24784
rect 2640 24750 2674 24784
rect 2708 24750 2742 24784
rect 2776 24750 2810 24784
rect 2844 24750 2878 24784
rect 2912 24750 2946 24784
rect 2980 24750 3014 24784
rect 3048 24750 3082 24784
rect 3116 24750 3150 24784
rect 3184 24750 3218 24784
rect 3252 24750 3286 24784
rect 3320 24750 3354 24784
rect 3388 24750 3422 24784
rect 3456 24750 3574 24784
rect 3873 25294 3991 25328
rect 4025 25294 4059 25328
rect 4093 25294 4127 25328
rect 4161 25294 4195 25328
rect 4229 25294 4263 25328
rect 4297 25294 4331 25328
rect 4365 25294 4399 25328
rect 4433 25294 4467 25328
rect 4501 25294 4535 25328
rect 4569 25294 4603 25328
rect 4637 25294 4671 25328
rect 4705 25294 4739 25328
rect 4773 25294 4807 25328
rect 4841 25294 4875 25328
rect 4909 25294 4943 25328
rect 4977 25294 5095 25328
rect 3873 25226 3907 25294
rect 3873 25158 3907 25192
rect 5061 25226 5095 25294
rect 5061 25158 5095 25192
rect 3873 25090 3907 25124
rect 3873 25022 3907 25056
rect 3873 24954 3907 24988
rect 3873 24886 3907 24920
rect 5061 25090 5095 25124
rect 5061 25022 5095 25056
rect 5061 24954 5095 24988
rect 5061 24886 5095 24920
rect 3873 24784 3907 24852
rect 5061 24784 5095 24852
rect 3873 24750 3991 24784
rect 4025 24750 4059 24784
rect 4093 24750 4127 24784
rect 4161 24750 4195 24784
rect 4229 24750 4263 24784
rect 4297 24750 4331 24784
rect 4365 24750 4399 24784
rect 4433 24750 4467 24784
rect 4501 24750 4535 24784
rect 4569 24750 4603 24784
rect 4637 24750 4671 24784
rect 4705 24750 4739 24784
rect 4773 24750 4807 24784
rect 4841 24750 4875 24784
rect 4909 24750 4943 24784
rect 4977 24750 5095 24784
rect 199 24003 317 24037
rect 351 24003 385 24037
rect 419 24003 453 24037
rect 487 24003 521 24037
rect 555 24003 589 24037
rect 623 24003 657 24037
rect 691 24003 725 24037
rect 759 24003 793 24037
rect 827 24003 861 24037
rect 895 24003 929 24037
rect 963 24003 997 24037
rect 1031 24003 1065 24037
rect 1099 24003 1133 24037
rect 1167 24003 1201 24037
rect 1235 24003 1269 24037
rect 1303 24003 1421 24037
rect 199 23935 233 24003
rect 199 23867 233 23901
rect 1387 23935 1421 24003
rect 1387 23867 1421 23901
rect 199 23799 233 23833
rect 199 23731 233 23765
rect 199 23663 233 23697
rect 199 23595 233 23629
rect 1387 23799 1421 23833
rect 1387 23731 1421 23765
rect 1387 23663 1421 23697
rect 1387 23595 1421 23629
rect 199 23493 233 23561
rect 1387 23493 1421 23561
rect 199 23459 317 23493
rect 351 23459 385 23493
rect 419 23459 453 23493
rect 487 23459 521 23493
rect 555 23459 589 23493
rect 623 23459 657 23493
rect 691 23459 725 23493
rect 759 23459 793 23493
rect 827 23459 861 23493
rect 895 23459 929 23493
rect 963 23459 997 23493
rect 1031 23459 1065 23493
rect 1099 23459 1133 23493
rect 1167 23459 1201 23493
rect 1235 23459 1269 23493
rect 1303 23459 1421 23493
rect 2352 24007 2470 24041
rect 2504 24007 2538 24041
rect 2572 24007 2606 24041
rect 2640 24007 2674 24041
rect 2708 24007 2742 24041
rect 2776 24007 2810 24041
rect 2844 24007 2878 24041
rect 2912 24007 2946 24041
rect 2980 24007 3014 24041
rect 3048 24007 3082 24041
rect 3116 24007 3150 24041
rect 3184 24007 3218 24041
rect 3252 24007 3286 24041
rect 3320 24007 3354 24041
rect 3388 24007 3422 24041
rect 3456 24007 3574 24041
rect 2352 23939 2386 24007
rect 2352 23871 2386 23905
rect 3540 23939 3574 24007
rect 3540 23871 3574 23905
rect 2352 23803 2386 23837
rect 2352 23735 2386 23769
rect 2352 23667 2386 23701
rect 2352 23599 2386 23633
rect 3540 23803 3574 23837
rect 3540 23735 3574 23769
rect 3540 23667 3574 23701
rect 3540 23599 3574 23633
rect 2352 23497 2386 23565
rect 3540 23497 3574 23565
rect 2352 23463 2470 23497
rect 2504 23463 2538 23497
rect 2572 23463 2606 23497
rect 2640 23463 2674 23497
rect 2708 23463 2742 23497
rect 2776 23463 2810 23497
rect 2844 23463 2878 23497
rect 2912 23463 2946 23497
rect 2980 23463 3014 23497
rect 3048 23463 3082 23497
rect 3116 23463 3150 23497
rect 3184 23463 3218 23497
rect 3252 23463 3286 23497
rect 3320 23463 3354 23497
rect 3388 23463 3422 23497
rect 3456 23463 3574 23497
rect 3873 24007 3991 24041
rect 4025 24007 4059 24041
rect 4093 24007 4127 24041
rect 4161 24007 4195 24041
rect 4229 24007 4263 24041
rect 4297 24007 4331 24041
rect 4365 24007 4399 24041
rect 4433 24007 4467 24041
rect 4501 24007 4535 24041
rect 4569 24007 4603 24041
rect 4637 24007 4671 24041
rect 4705 24007 4739 24041
rect 4773 24007 4807 24041
rect 4841 24007 4875 24041
rect 4909 24007 4943 24041
rect 4977 24007 5095 24041
rect 3873 23939 3907 24007
rect 3873 23871 3907 23905
rect 5061 23939 5095 24007
rect 5061 23871 5095 23905
rect 3873 23803 3907 23837
rect 3873 23735 3907 23769
rect 3873 23667 3907 23701
rect 3873 23599 3907 23633
rect 5061 23803 5095 23837
rect 5061 23735 5095 23769
rect 5061 23667 5095 23701
rect 5061 23599 5095 23633
rect 3873 23497 3907 23565
rect 5061 23497 5095 23565
rect 3873 23463 3991 23497
rect 4025 23463 4059 23497
rect 4093 23463 4127 23497
rect 4161 23463 4195 23497
rect 4229 23463 4263 23497
rect 4297 23463 4331 23497
rect 4365 23463 4399 23497
rect 4433 23463 4467 23497
rect 4501 23463 4535 23497
rect 4569 23463 4603 23497
rect 4637 23463 4671 23497
rect 4705 23463 4739 23497
rect 4773 23463 4807 23497
rect 4841 23463 4875 23497
rect 4909 23463 4943 23497
rect 4977 23463 5095 23497
rect 199 22716 317 22750
rect 351 22716 385 22750
rect 419 22716 453 22750
rect 487 22716 521 22750
rect 555 22716 589 22750
rect 623 22716 657 22750
rect 691 22716 725 22750
rect 759 22716 793 22750
rect 827 22716 861 22750
rect 895 22716 929 22750
rect 963 22716 997 22750
rect 1031 22716 1065 22750
rect 1099 22716 1133 22750
rect 1167 22716 1201 22750
rect 1235 22716 1269 22750
rect 1303 22716 1421 22750
rect 199 22648 233 22716
rect 199 22580 233 22614
rect 1387 22648 1421 22716
rect 1387 22580 1421 22614
rect 199 22512 233 22546
rect 199 22444 233 22478
rect 199 22376 233 22410
rect 199 22308 233 22342
rect 1387 22512 1421 22546
rect 1387 22444 1421 22478
rect 1387 22376 1421 22410
rect 1387 22308 1421 22342
rect 199 22206 233 22274
rect 1387 22206 1421 22274
rect 199 22172 317 22206
rect 351 22172 385 22206
rect 419 22172 453 22206
rect 487 22172 521 22206
rect 555 22172 589 22206
rect 623 22172 657 22206
rect 691 22172 725 22206
rect 759 22172 793 22206
rect 827 22172 861 22206
rect 895 22172 929 22206
rect 963 22172 997 22206
rect 1031 22172 1065 22206
rect 1099 22172 1133 22206
rect 1167 22172 1201 22206
rect 1235 22172 1269 22206
rect 1303 22172 1421 22206
rect 2352 22720 2470 22754
rect 2504 22720 2538 22754
rect 2572 22720 2606 22754
rect 2640 22720 2674 22754
rect 2708 22720 2742 22754
rect 2776 22720 2810 22754
rect 2844 22720 2878 22754
rect 2912 22720 2946 22754
rect 2980 22720 3014 22754
rect 3048 22720 3082 22754
rect 3116 22720 3150 22754
rect 3184 22720 3218 22754
rect 3252 22720 3286 22754
rect 3320 22720 3354 22754
rect 3388 22720 3422 22754
rect 3456 22720 3574 22754
rect 2352 22652 2386 22720
rect 2352 22584 2386 22618
rect 3540 22652 3574 22720
rect 3540 22584 3574 22618
rect 2352 22516 2386 22550
rect 2352 22448 2386 22482
rect 2352 22380 2386 22414
rect 2352 22312 2386 22346
rect 3540 22516 3574 22550
rect 3540 22448 3574 22482
rect 3540 22380 3574 22414
rect 3540 22312 3574 22346
rect 2352 22210 2386 22278
rect 3540 22210 3574 22278
rect 2352 22176 2470 22210
rect 2504 22176 2538 22210
rect 2572 22176 2606 22210
rect 2640 22176 2674 22210
rect 2708 22176 2742 22210
rect 2776 22176 2810 22210
rect 2844 22176 2878 22210
rect 2912 22176 2946 22210
rect 2980 22176 3014 22210
rect 3048 22176 3082 22210
rect 3116 22176 3150 22210
rect 3184 22176 3218 22210
rect 3252 22176 3286 22210
rect 3320 22176 3354 22210
rect 3388 22176 3422 22210
rect 3456 22176 3574 22210
rect 3873 22720 3991 22754
rect 4025 22720 4059 22754
rect 4093 22720 4127 22754
rect 4161 22720 4195 22754
rect 4229 22720 4263 22754
rect 4297 22720 4331 22754
rect 4365 22720 4399 22754
rect 4433 22720 4467 22754
rect 4501 22720 4535 22754
rect 4569 22720 4603 22754
rect 4637 22720 4671 22754
rect 4705 22720 4739 22754
rect 4773 22720 4807 22754
rect 4841 22720 4875 22754
rect 4909 22720 4943 22754
rect 4977 22720 5095 22754
rect 3873 22652 3907 22720
rect 3873 22584 3907 22618
rect 5061 22652 5095 22720
rect 5061 22584 5095 22618
rect 3873 22516 3907 22550
rect 3873 22448 3907 22482
rect 3873 22380 3907 22414
rect 3873 22312 3907 22346
rect 5061 22516 5095 22550
rect 5061 22448 5095 22482
rect 5061 22380 5095 22414
rect 5061 22312 5095 22346
rect 3873 22210 3907 22278
rect 5061 22210 5095 22278
rect 3873 22176 3991 22210
rect 4025 22176 4059 22210
rect 4093 22176 4127 22210
rect 4161 22176 4195 22210
rect 4229 22176 4263 22210
rect 4297 22176 4331 22210
rect 4365 22176 4399 22210
rect 4433 22176 4467 22210
rect 4501 22176 4535 22210
rect 4569 22176 4603 22210
rect 4637 22176 4671 22210
rect 4705 22176 4739 22210
rect 4773 22176 4807 22210
rect 4841 22176 4875 22210
rect 4909 22176 4943 22210
rect 4977 22176 5095 22210
rect 199 21429 317 21463
rect 351 21429 385 21463
rect 419 21429 453 21463
rect 487 21429 521 21463
rect 555 21429 589 21463
rect 623 21429 657 21463
rect 691 21429 725 21463
rect 759 21429 793 21463
rect 827 21429 861 21463
rect 895 21429 929 21463
rect 963 21429 997 21463
rect 1031 21429 1065 21463
rect 1099 21429 1133 21463
rect 1167 21429 1201 21463
rect 1235 21429 1269 21463
rect 1303 21429 1421 21463
rect 199 21361 233 21429
rect 199 21293 233 21327
rect 1387 21361 1421 21429
rect 1387 21293 1421 21327
rect 199 21225 233 21259
rect 199 21157 233 21191
rect 199 21089 233 21123
rect 199 21021 233 21055
rect 1387 21225 1421 21259
rect 1387 21157 1421 21191
rect 1387 21089 1421 21123
rect 1387 21021 1421 21055
rect 199 20919 233 20987
rect 1387 20919 1421 20987
rect 199 20885 317 20919
rect 351 20885 385 20919
rect 419 20885 453 20919
rect 487 20885 521 20919
rect 555 20885 589 20919
rect 623 20885 657 20919
rect 691 20885 725 20919
rect 759 20885 793 20919
rect 827 20885 861 20919
rect 895 20885 929 20919
rect 963 20885 997 20919
rect 1031 20885 1065 20919
rect 1099 20885 1133 20919
rect 1167 20885 1201 20919
rect 1235 20885 1269 20919
rect 1303 20885 1421 20919
rect 2352 21433 2470 21467
rect 2504 21433 2538 21467
rect 2572 21433 2606 21467
rect 2640 21433 2674 21467
rect 2708 21433 2742 21467
rect 2776 21433 2810 21467
rect 2844 21433 2878 21467
rect 2912 21433 2946 21467
rect 2980 21433 3014 21467
rect 3048 21433 3082 21467
rect 3116 21433 3150 21467
rect 3184 21433 3218 21467
rect 3252 21433 3286 21467
rect 3320 21433 3354 21467
rect 3388 21433 3422 21467
rect 3456 21433 3574 21467
rect 2352 21365 2386 21433
rect 2352 21297 2386 21331
rect 3540 21365 3574 21433
rect 3540 21297 3574 21331
rect 2352 21229 2386 21263
rect 2352 21161 2386 21195
rect 2352 21093 2386 21127
rect 2352 21025 2386 21059
rect 3540 21229 3574 21263
rect 3540 21161 3574 21195
rect 3540 21093 3574 21127
rect 3540 21025 3574 21059
rect 2352 20923 2386 20991
rect 3540 20923 3574 20991
rect 2352 20889 2470 20923
rect 2504 20889 2538 20923
rect 2572 20889 2606 20923
rect 2640 20889 2674 20923
rect 2708 20889 2742 20923
rect 2776 20889 2810 20923
rect 2844 20889 2878 20923
rect 2912 20889 2946 20923
rect 2980 20889 3014 20923
rect 3048 20889 3082 20923
rect 3116 20889 3150 20923
rect 3184 20889 3218 20923
rect 3252 20889 3286 20923
rect 3320 20889 3354 20923
rect 3388 20889 3422 20923
rect 3456 20889 3574 20923
rect 3873 21433 3991 21467
rect 4025 21433 4059 21467
rect 4093 21433 4127 21467
rect 4161 21433 4195 21467
rect 4229 21433 4263 21467
rect 4297 21433 4331 21467
rect 4365 21433 4399 21467
rect 4433 21433 4467 21467
rect 4501 21433 4535 21467
rect 4569 21433 4603 21467
rect 4637 21433 4671 21467
rect 4705 21433 4739 21467
rect 4773 21433 4807 21467
rect 4841 21433 4875 21467
rect 4909 21433 4943 21467
rect 4977 21433 5095 21467
rect 3873 21365 3907 21433
rect 3873 21297 3907 21331
rect 5061 21365 5095 21433
rect 5061 21297 5095 21331
rect 3873 21229 3907 21263
rect 3873 21161 3907 21195
rect 3873 21093 3907 21127
rect 3873 21025 3907 21059
rect 5061 21229 5095 21263
rect 5061 21161 5095 21195
rect 5061 21093 5095 21127
rect 5061 21025 5095 21059
rect 3873 20923 3907 20991
rect 5061 20923 5095 20991
rect 3873 20889 3991 20923
rect 4025 20889 4059 20923
rect 4093 20889 4127 20923
rect 4161 20889 4195 20923
rect 4229 20889 4263 20923
rect 4297 20889 4331 20923
rect 4365 20889 4399 20923
rect 4433 20889 4467 20923
rect 4501 20889 4535 20923
rect 4569 20889 4603 20923
rect 4637 20889 4671 20923
rect 4705 20889 4739 20923
rect 4773 20889 4807 20923
rect 4841 20889 4875 20923
rect 4909 20889 4943 20923
rect 4977 20889 5095 20923
rect 199 20142 317 20176
rect 351 20142 385 20176
rect 419 20142 453 20176
rect 487 20142 521 20176
rect 555 20142 589 20176
rect 623 20142 657 20176
rect 691 20142 725 20176
rect 759 20142 793 20176
rect 827 20142 861 20176
rect 895 20142 929 20176
rect 963 20142 997 20176
rect 1031 20142 1065 20176
rect 1099 20142 1133 20176
rect 1167 20142 1201 20176
rect 1235 20142 1269 20176
rect 1303 20142 1421 20176
rect 199 20074 233 20142
rect 199 20006 233 20040
rect 1387 20074 1421 20142
rect 1387 20006 1421 20040
rect 199 19938 233 19972
rect 199 19870 233 19904
rect 199 19802 233 19836
rect 199 19734 233 19768
rect 1387 19938 1421 19972
rect 1387 19870 1421 19904
rect 1387 19802 1421 19836
rect 1387 19734 1421 19768
rect 199 19632 233 19700
rect 1387 19632 1421 19700
rect 199 19598 317 19632
rect 351 19598 385 19632
rect 419 19598 453 19632
rect 487 19598 521 19632
rect 555 19598 589 19632
rect 623 19598 657 19632
rect 691 19598 725 19632
rect 759 19598 793 19632
rect 827 19598 861 19632
rect 895 19598 929 19632
rect 963 19598 997 19632
rect 1031 19598 1065 19632
rect 1099 19598 1133 19632
rect 1167 19598 1201 19632
rect 1235 19598 1269 19632
rect 1303 19598 1421 19632
rect 2352 20146 2470 20180
rect 2504 20146 2538 20180
rect 2572 20146 2606 20180
rect 2640 20146 2674 20180
rect 2708 20146 2742 20180
rect 2776 20146 2810 20180
rect 2844 20146 2878 20180
rect 2912 20146 2946 20180
rect 2980 20146 3014 20180
rect 3048 20146 3082 20180
rect 3116 20146 3150 20180
rect 3184 20146 3218 20180
rect 3252 20146 3286 20180
rect 3320 20146 3354 20180
rect 3388 20146 3422 20180
rect 3456 20146 3574 20180
rect 2352 20078 2386 20146
rect 2352 20010 2386 20044
rect 3540 20078 3574 20146
rect 3540 20010 3574 20044
rect 2352 19942 2386 19976
rect 2352 19874 2386 19908
rect 2352 19806 2386 19840
rect 2352 19738 2386 19772
rect 3540 19942 3574 19976
rect 3540 19874 3574 19908
rect 3540 19806 3574 19840
rect 3540 19738 3574 19772
rect 2352 19636 2386 19704
rect 3540 19636 3574 19704
rect 2352 19602 2470 19636
rect 2504 19602 2538 19636
rect 2572 19602 2606 19636
rect 2640 19602 2674 19636
rect 2708 19602 2742 19636
rect 2776 19602 2810 19636
rect 2844 19602 2878 19636
rect 2912 19602 2946 19636
rect 2980 19602 3014 19636
rect 3048 19602 3082 19636
rect 3116 19602 3150 19636
rect 3184 19602 3218 19636
rect 3252 19602 3286 19636
rect 3320 19602 3354 19636
rect 3388 19602 3422 19636
rect 3456 19602 3574 19636
rect 3873 20146 3991 20180
rect 4025 20146 4059 20180
rect 4093 20146 4127 20180
rect 4161 20146 4195 20180
rect 4229 20146 4263 20180
rect 4297 20146 4331 20180
rect 4365 20146 4399 20180
rect 4433 20146 4467 20180
rect 4501 20146 4535 20180
rect 4569 20146 4603 20180
rect 4637 20146 4671 20180
rect 4705 20146 4739 20180
rect 4773 20146 4807 20180
rect 4841 20146 4875 20180
rect 4909 20146 4943 20180
rect 4977 20146 5095 20180
rect 3873 20078 3907 20146
rect 3873 20010 3907 20044
rect 5061 20078 5095 20146
rect 5061 20010 5095 20044
rect 3873 19942 3907 19976
rect 3873 19874 3907 19908
rect 3873 19806 3907 19840
rect 3873 19738 3907 19772
rect 5061 19942 5095 19976
rect 5061 19874 5095 19908
rect 5061 19806 5095 19840
rect 5061 19738 5095 19772
rect 3873 19636 3907 19704
rect 5061 19636 5095 19704
rect 3873 19602 3991 19636
rect 4025 19602 4059 19636
rect 4093 19602 4127 19636
rect 4161 19602 4195 19636
rect 4229 19602 4263 19636
rect 4297 19602 4331 19636
rect 4365 19602 4399 19636
rect 4433 19602 4467 19636
rect 4501 19602 4535 19636
rect 4569 19602 4603 19636
rect 4637 19602 4671 19636
rect 4705 19602 4739 19636
rect 4773 19602 4807 19636
rect 4841 19602 4875 19636
rect 4909 19602 4943 19636
rect 4977 19602 5095 19636
rect 199 18855 317 18889
rect 351 18855 385 18889
rect 419 18855 453 18889
rect 487 18855 521 18889
rect 555 18855 589 18889
rect 623 18855 657 18889
rect 691 18855 725 18889
rect 759 18855 793 18889
rect 827 18855 861 18889
rect 895 18855 929 18889
rect 963 18855 997 18889
rect 1031 18855 1065 18889
rect 1099 18855 1133 18889
rect 1167 18855 1201 18889
rect 1235 18855 1269 18889
rect 1303 18855 1421 18889
rect 199 18787 233 18855
rect 199 18719 233 18753
rect 1387 18787 1421 18855
rect 1387 18719 1421 18753
rect 199 18651 233 18685
rect 199 18583 233 18617
rect 199 18515 233 18549
rect 199 18447 233 18481
rect 1387 18651 1421 18685
rect 1387 18583 1421 18617
rect 1387 18515 1421 18549
rect 1387 18447 1421 18481
rect 199 18345 233 18413
rect 1387 18345 1421 18413
rect 199 18311 317 18345
rect 351 18311 385 18345
rect 419 18311 453 18345
rect 487 18311 521 18345
rect 555 18311 589 18345
rect 623 18311 657 18345
rect 691 18311 725 18345
rect 759 18311 793 18345
rect 827 18311 861 18345
rect 895 18311 929 18345
rect 963 18311 997 18345
rect 1031 18311 1065 18345
rect 1099 18311 1133 18345
rect 1167 18311 1201 18345
rect 1235 18311 1269 18345
rect 1303 18311 1421 18345
rect 2352 18859 2470 18893
rect 2504 18859 2538 18893
rect 2572 18859 2606 18893
rect 2640 18859 2674 18893
rect 2708 18859 2742 18893
rect 2776 18859 2810 18893
rect 2844 18859 2878 18893
rect 2912 18859 2946 18893
rect 2980 18859 3014 18893
rect 3048 18859 3082 18893
rect 3116 18859 3150 18893
rect 3184 18859 3218 18893
rect 3252 18859 3286 18893
rect 3320 18859 3354 18893
rect 3388 18859 3422 18893
rect 3456 18859 3574 18893
rect 2352 18791 2386 18859
rect 2352 18723 2386 18757
rect 3540 18791 3574 18859
rect 3540 18723 3574 18757
rect 2352 18655 2386 18689
rect 2352 18587 2386 18621
rect 2352 18519 2386 18553
rect 2352 18451 2386 18485
rect 3540 18655 3574 18689
rect 3540 18587 3574 18621
rect 3540 18519 3574 18553
rect 3540 18451 3574 18485
rect 2352 18349 2386 18417
rect 3540 18349 3574 18417
rect 2352 18315 2470 18349
rect 2504 18315 2538 18349
rect 2572 18315 2606 18349
rect 2640 18315 2674 18349
rect 2708 18315 2742 18349
rect 2776 18315 2810 18349
rect 2844 18315 2878 18349
rect 2912 18315 2946 18349
rect 2980 18315 3014 18349
rect 3048 18315 3082 18349
rect 3116 18315 3150 18349
rect 3184 18315 3218 18349
rect 3252 18315 3286 18349
rect 3320 18315 3354 18349
rect 3388 18315 3422 18349
rect 3456 18315 3574 18349
rect 3873 18859 3991 18893
rect 4025 18859 4059 18893
rect 4093 18859 4127 18893
rect 4161 18859 4195 18893
rect 4229 18859 4263 18893
rect 4297 18859 4331 18893
rect 4365 18859 4399 18893
rect 4433 18859 4467 18893
rect 4501 18859 4535 18893
rect 4569 18859 4603 18893
rect 4637 18859 4671 18893
rect 4705 18859 4739 18893
rect 4773 18859 4807 18893
rect 4841 18859 4875 18893
rect 4909 18859 4943 18893
rect 4977 18859 5095 18893
rect 3873 18791 3907 18859
rect 3873 18723 3907 18757
rect 5061 18791 5095 18859
rect 5061 18723 5095 18757
rect 3873 18655 3907 18689
rect 3873 18587 3907 18621
rect 3873 18519 3907 18553
rect 3873 18451 3907 18485
rect 5061 18655 5095 18689
rect 5061 18587 5095 18621
rect 5061 18519 5095 18553
rect 5061 18451 5095 18485
rect 3873 18349 3907 18417
rect 5061 18349 5095 18417
rect 3873 18315 3991 18349
rect 4025 18315 4059 18349
rect 4093 18315 4127 18349
rect 4161 18315 4195 18349
rect 4229 18315 4263 18349
rect 4297 18315 4331 18349
rect 4365 18315 4399 18349
rect 4433 18315 4467 18349
rect 4501 18315 4535 18349
rect 4569 18315 4603 18349
rect 4637 18315 4671 18349
rect 4705 18315 4739 18349
rect 4773 18315 4807 18349
rect 4841 18315 4875 18349
rect 4909 18315 4943 18349
rect 4977 18315 5095 18349
rect 199 17568 317 17602
rect 351 17568 385 17602
rect 419 17568 453 17602
rect 487 17568 521 17602
rect 555 17568 589 17602
rect 623 17568 657 17602
rect 691 17568 725 17602
rect 759 17568 793 17602
rect 827 17568 861 17602
rect 895 17568 929 17602
rect 963 17568 997 17602
rect 1031 17568 1065 17602
rect 1099 17568 1133 17602
rect 1167 17568 1201 17602
rect 1235 17568 1269 17602
rect 1303 17568 1421 17602
rect 199 17500 233 17568
rect 199 17432 233 17466
rect 1387 17500 1421 17568
rect 1387 17432 1421 17466
rect 199 17364 233 17398
rect 199 17296 233 17330
rect 199 17228 233 17262
rect 199 17160 233 17194
rect 1387 17364 1421 17398
rect 1387 17296 1421 17330
rect 1387 17228 1421 17262
rect 1387 17160 1421 17194
rect 199 17058 233 17126
rect 1387 17058 1421 17126
rect 199 17024 317 17058
rect 351 17024 385 17058
rect 419 17024 453 17058
rect 487 17024 521 17058
rect 555 17024 589 17058
rect 623 17024 657 17058
rect 691 17024 725 17058
rect 759 17024 793 17058
rect 827 17024 861 17058
rect 895 17024 929 17058
rect 963 17024 997 17058
rect 1031 17024 1065 17058
rect 1099 17024 1133 17058
rect 1167 17024 1201 17058
rect 1235 17024 1269 17058
rect 1303 17024 1421 17058
rect 2352 17572 2470 17606
rect 2504 17572 2538 17606
rect 2572 17572 2606 17606
rect 2640 17572 2674 17606
rect 2708 17572 2742 17606
rect 2776 17572 2810 17606
rect 2844 17572 2878 17606
rect 2912 17572 2946 17606
rect 2980 17572 3014 17606
rect 3048 17572 3082 17606
rect 3116 17572 3150 17606
rect 3184 17572 3218 17606
rect 3252 17572 3286 17606
rect 3320 17572 3354 17606
rect 3388 17572 3422 17606
rect 3456 17572 3574 17606
rect 2352 17504 2386 17572
rect 2352 17436 2386 17470
rect 3540 17504 3574 17572
rect 3540 17436 3574 17470
rect 2352 17368 2386 17402
rect 2352 17300 2386 17334
rect 2352 17232 2386 17266
rect 2352 17164 2386 17198
rect 3540 17368 3574 17402
rect 3540 17300 3574 17334
rect 3540 17232 3574 17266
rect 3540 17164 3574 17198
rect 2352 17062 2386 17130
rect 3540 17062 3574 17130
rect 2352 17028 2470 17062
rect 2504 17028 2538 17062
rect 2572 17028 2606 17062
rect 2640 17028 2674 17062
rect 2708 17028 2742 17062
rect 2776 17028 2810 17062
rect 2844 17028 2878 17062
rect 2912 17028 2946 17062
rect 2980 17028 3014 17062
rect 3048 17028 3082 17062
rect 3116 17028 3150 17062
rect 3184 17028 3218 17062
rect 3252 17028 3286 17062
rect 3320 17028 3354 17062
rect 3388 17028 3422 17062
rect 3456 17028 3574 17062
rect 3873 17572 3991 17606
rect 4025 17572 4059 17606
rect 4093 17572 4127 17606
rect 4161 17572 4195 17606
rect 4229 17572 4263 17606
rect 4297 17572 4331 17606
rect 4365 17572 4399 17606
rect 4433 17572 4467 17606
rect 4501 17572 4535 17606
rect 4569 17572 4603 17606
rect 4637 17572 4671 17606
rect 4705 17572 4739 17606
rect 4773 17572 4807 17606
rect 4841 17572 4875 17606
rect 4909 17572 4943 17606
rect 4977 17572 5095 17606
rect 3873 17504 3907 17572
rect 3873 17436 3907 17470
rect 5061 17504 5095 17572
rect 5061 17436 5095 17470
rect 3873 17368 3907 17402
rect 3873 17300 3907 17334
rect 3873 17232 3907 17266
rect 3873 17164 3907 17198
rect 5061 17368 5095 17402
rect 5061 17300 5095 17334
rect 5061 17232 5095 17266
rect 5061 17164 5095 17198
rect 3873 17062 3907 17130
rect 5061 17062 5095 17130
rect 3873 17028 3991 17062
rect 4025 17028 4059 17062
rect 4093 17028 4127 17062
rect 4161 17028 4195 17062
rect 4229 17028 4263 17062
rect 4297 17028 4331 17062
rect 4365 17028 4399 17062
rect 4433 17028 4467 17062
rect 4501 17028 4535 17062
rect 4569 17028 4603 17062
rect 4637 17028 4671 17062
rect 4705 17028 4739 17062
rect 4773 17028 4807 17062
rect 4841 17028 4875 17062
rect 4909 17028 4943 17062
rect 4977 17028 5095 17062
rect 199 16281 317 16315
rect 351 16281 385 16315
rect 419 16281 453 16315
rect 487 16281 521 16315
rect 555 16281 589 16315
rect 623 16281 657 16315
rect 691 16281 725 16315
rect 759 16281 793 16315
rect 827 16281 861 16315
rect 895 16281 929 16315
rect 963 16281 997 16315
rect 1031 16281 1065 16315
rect 1099 16281 1133 16315
rect 1167 16281 1201 16315
rect 1235 16281 1269 16315
rect 1303 16281 1421 16315
rect 199 16213 233 16281
rect 199 16145 233 16179
rect 1387 16213 1421 16281
rect 1387 16145 1421 16179
rect 199 16077 233 16111
rect 199 16009 233 16043
rect 199 15941 233 15975
rect 199 15873 233 15907
rect 1387 16077 1421 16111
rect 1387 16009 1421 16043
rect 1387 15941 1421 15975
rect 1387 15873 1421 15907
rect 199 15771 233 15839
rect 1387 15771 1421 15839
rect 199 15737 317 15771
rect 351 15737 385 15771
rect 419 15737 453 15771
rect 487 15737 521 15771
rect 555 15737 589 15771
rect 623 15737 657 15771
rect 691 15737 725 15771
rect 759 15737 793 15771
rect 827 15737 861 15771
rect 895 15737 929 15771
rect 963 15737 997 15771
rect 1031 15737 1065 15771
rect 1099 15737 1133 15771
rect 1167 15737 1201 15771
rect 1235 15737 1269 15771
rect 1303 15737 1421 15771
rect 2352 16285 2470 16319
rect 2504 16285 2538 16319
rect 2572 16285 2606 16319
rect 2640 16285 2674 16319
rect 2708 16285 2742 16319
rect 2776 16285 2810 16319
rect 2844 16285 2878 16319
rect 2912 16285 2946 16319
rect 2980 16285 3014 16319
rect 3048 16285 3082 16319
rect 3116 16285 3150 16319
rect 3184 16285 3218 16319
rect 3252 16285 3286 16319
rect 3320 16285 3354 16319
rect 3388 16285 3422 16319
rect 3456 16285 3574 16319
rect 2352 16217 2386 16285
rect 2352 16149 2386 16183
rect 3540 16217 3574 16285
rect 3540 16149 3574 16183
rect 2352 16081 2386 16115
rect 2352 16013 2386 16047
rect 2352 15945 2386 15979
rect 2352 15877 2386 15911
rect 3540 16081 3574 16115
rect 3540 16013 3574 16047
rect 3540 15945 3574 15979
rect 3540 15877 3574 15911
rect 2352 15775 2386 15843
rect 3540 15775 3574 15843
rect 2352 15741 2470 15775
rect 2504 15741 2538 15775
rect 2572 15741 2606 15775
rect 2640 15741 2674 15775
rect 2708 15741 2742 15775
rect 2776 15741 2810 15775
rect 2844 15741 2878 15775
rect 2912 15741 2946 15775
rect 2980 15741 3014 15775
rect 3048 15741 3082 15775
rect 3116 15741 3150 15775
rect 3184 15741 3218 15775
rect 3252 15741 3286 15775
rect 3320 15741 3354 15775
rect 3388 15741 3422 15775
rect 3456 15741 3574 15775
rect 3873 16285 3991 16319
rect 4025 16285 4059 16319
rect 4093 16285 4127 16319
rect 4161 16285 4195 16319
rect 4229 16285 4263 16319
rect 4297 16285 4331 16319
rect 4365 16285 4399 16319
rect 4433 16285 4467 16319
rect 4501 16285 4535 16319
rect 4569 16285 4603 16319
rect 4637 16285 4671 16319
rect 4705 16285 4739 16319
rect 4773 16285 4807 16319
rect 4841 16285 4875 16319
rect 4909 16285 4943 16319
rect 4977 16285 5095 16319
rect 3873 16217 3907 16285
rect 3873 16149 3907 16183
rect 5061 16217 5095 16285
rect 5061 16149 5095 16183
rect 3873 16081 3907 16115
rect 3873 16013 3907 16047
rect 3873 15945 3907 15979
rect 3873 15877 3907 15911
rect 5061 16081 5095 16115
rect 5061 16013 5095 16047
rect 5061 15945 5095 15979
rect 5061 15877 5095 15911
rect 3873 15775 3907 15843
rect 5061 15775 5095 15843
rect 3873 15741 3991 15775
rect 4025 15741 4059 15775
rect 4093 15741 4127 15775
rect 4161 15741 4195 15775
rect 4229 15741 4263 15775
rect 4297 15741 4331 15775
rect 4365 15741 4399 15775
rect 4433 15741 4467 15775
rect 4501 15741 4535 15775
rect 4569 15741 4603 15775
rect 4637 15741 4671 15775
rect 4705 15741 4739 15775
rect 4773 15741 4807 15775
rect 4841 15741 4875 15775
rect 4909 15741 4943 15775
rect 4977 15741 5095 15775
rect 199 14994 317 15028
rect 351 14994 385 15028
rect 419 14994 453 15028
rect 487 14994 521 15028
rect 555 14994 589 15028
rect 623 14994 657 15028
rect 691 14994 725 15028
rect 759 14994 793 15028
rect 827 14994 861 15028
rect 895 14994 929 15028
rect 963 14994 997 15028
rect 1031 14994 1065 15028
rect 1099 14994 1133 15028
rect 1167 14994 1201 15028
rect 1235 14994 1269 15028
rect 1303 14994 1421 15028
rect 199 14926 233 14994
rect 199 14858 233 14892
rect 1387 14926 1421 14994
rect 1387 14858 1421 14892
rect 199 14790 233 14824
rect 199 14722 233 14756
rect 199 14654 233 14688
rect 199 14586 233 14620
rect 1387 14790 1421 14824
rect 1387 14722 1421 14756
rect 1387 14654 1421 14688
rect 1387 14586 1421 14620
rect 199 14484 233 14552
rect 1387 14484 1421 14552
rect 199 14450 317 14484
rect 351 14450 385 14484
rect 419 14450 453 14484
rect 487 14450 521 14484
rect 555 14450 589 14484
rect 623 14450 657 14484
rect 691 14450 725 14484
rect 759 14450 793 14484
rect 827 14450 861 14484
rect 895 14450 929 14484
rect 963 14450 997 14484
rect 1031 14450 1065 14484
rect 1099 14450 1133 14484
rect 1167 14450 1201 14484
rect 1235 14450 1269 14484
rect 1303 14450 1421 14484
rect 2352 14998 2470 15032
rect 2504 14998 2538 15032
rect 2572 14998 2606 15032
rect 2640 14998 2674 15032
rect 2708 14998 2742 15032
rect 2776 14998 2810 15032
rect 2844 14998 2878 15032
rect 2912 14998 2946 15032
rect 2980 14998 3014 15032
rect 3048 14998 3082 15032
rect 3116 14998 3150 15032
rect 3184 14998 3218 15032
rect 3252 14998 3286 15032
rect 3320 14998 3354 15032
rect 3388 14998 3422 15032
rect 3456 14998 3574 15032
rect 2352 14930 2386 14998
rect 2352 14862 2386 14896
rect 3540 14930 3574 14998
rect 3540 14862 3574 14896
rect 2352 14794 2386 14828
rect 2352 14726 2386 14760
rect 2352 14658 2386 14692
rect 2352 14590 2386 14624
rect 3540 14794 3574 14828
rect 3540 14726 3574 14760
rect 3540 14658 3574 14692
rect 3540 14590 3574 14624
rect 2352 14488 2386 14556
rect 3540 14488 3574 14556
rect 2352 14454 2470 14488
rect 2504 14454 2538 14488
rect 2572 14454 2606 14488
rect 2640 14454 2674 14488
rect 2708 14454 2742 14488
rect 2776 14454 2810 14488
rect 2844 14454 2878 14488
rect 2912 14454 2946 14488
rect 2980 14454 3014 14488
rect 3048 14454 3082 14488
rect 3116 14454 3150 14488
rect 3184 14454 3218 14488
rect 3252 14454 3286 14488
rect 3320 14454 3354 14488
rect 3388 14454 3422 14488
rect 3456 14454 3574 14488
rect 3873 14998 3991 15032
rect 4025 14998 4059 15032
rect 4093 14998 4127 15032
rect 4161 14998 4195 15032
rect 4229 14998 4263 15032
rect 4297 14998 4331 15032
rect 4365 14998 4399 15032
rect 4433 14998 4467 15032
rect 4501 14998 4535 15032
rect 4569 14998 4603 15032
rect 4637 14998 4671 15032
rect 4705 14998 4739 15032
rect 4773 14998 4807 15032
rect 4841 14998 4875 15032
rect 4909 14998 4943 15032
rect 4977 14998 5095 15032
rect 3873 14930 3907 14998
rect 3873 14862 3907 14896
rect 5061 14930 5095 14998
rect 5061 14862 5095 14896
rect 3873 14794 3907 14828
rect 3873 14726 3907 14760
rect 3873 14658 3907 14692
rect 3873 14590 3907 14624
rect 5061 14794 5095 14828
rect 5061 14726 5095 14760
rect 5061 14658 5095 14692
rect 5061 14590 5095 14624
rect 3873 14488 3907 14556
rect 5061 14488 5095 14556
rect 3873 14454 3991 14488
rect 4025 14454 4059 14488
rect 4093 14454 4127 14488
rect 4161 14454 4195 14488
rect 4229 14454 4263 14488
rect 4297 14454 4331 14488
rect 4365 14454 4399 14488
rect 4433 14454 4467 14488
rect 4501 14454 4535 14488
rect 4569 14454 4603 14488
rect 4637 14454 4671 14488
rect 4705 14454 4739 14488
rect 4773 14454 4807 14488
rect 4841 14454 4875 14488
rect 4909 14454 4943 14488
rect 4977 14454 5095 14488
rect 199 13707 317 13741
rect 351 13707 385 13741
rect 419 13707 453 13741
rect 487 13707 521 13741
rect 555 13707 589 13741
rect 623 13707 657 13741
rect 691 13707 725 13741
rect 759 13707 793 13741
rect 827 13707 861 13741
rect 895 13707 929 13741
rect 963 13707 997 13741
rect 1031 13707 1065 13741
rect 1099 13707 1133 13741
rect 1167 13707 1201 13741
rect 1235 13707 1269 13741
rect 1303 13707 1421 13741
rect 199 13639 233 13707
rect 199 13571 233 13605
rect 1387 13639 1421 13707
rect 1387 13571 1421 13605
rect 199 13503 233 13537
rect 199 13435 233 13469
rect 199 13367 233 13401
rect 199 13299 233 13333
rect 1387 13503 1421 13537
rect 1387 13435 1421 13469
rect 1387 13367 1421 13401
rect 1387 13299 1421 13333
rect 199 13197 233 13265
rect 1387 13197 1421 13265
rect 199 13163 317 13197
rect 351 13163 385 13197
rect 419 13163 453 13197
rect 487 13163 521 13197
rect 555 13163 589 13197
rect 623 13163 657 13197
rect 691 13163 725 13197
rect 759 13163 793 13197
rect 827 13163 861 13197
rect 895 13163 929 13197
rect 963 13163 997 13197
rect 1031 13163 1065 13197
rect 1099 13163 1133 13197
rect 1167 13163 1201 13197
rect 1235 13163 1269 13197
rect 1303 13163 1421 13197
rect 2352 13711 2470 13745
rect 2504 13711 2538 13745
rect 2572 13711 2606 13745
rect 2640 13711 2674 13745
rect 2708 13711 2742 13745
rect 2776 13711 2810 13745
rect 2844 13711 2878 13745
rect 2912 13711 2946 13745
rect 2980 13711 3014 13745
rect 3048 13711 3082 13745
rect 3116 13711 3150 13745
rect 3184 13711 3218 13745
rect 3252 13711 3286 13745
rect 3320 13711 3354 13745
rect 3388 13711 3422 13745
rect 3456 13711 3574 13745
rect 2352 13643 2386 13711
rect 2352 13575 2386 13609
rect 3540 13643 3574 13711
rect 3540 13575 3574 13609
rect 2352 13507 2386 13541
rect 2352 13439 2386 13473
rect 2352 13371 2386 13405
rect 2352 13303 2386 13337
rect 3540 13507 3574 13541
rect 3540 13439 3574 13473
rect 3540 13371 3574 13405
rect 3540 13303 3574 13337
rect 2352 13201 2386 13269
rect 3540 13201 3574 13269
rect 2352 13167 2470 13201
rect 2504 13167 2538 13201
rect 2572 13167 2606 13201
rect 2640 13167 2674 13201
rect 2708 13167 2742 13201
rect 2776 13167 2810 13201
rect 2844 13167 2878 13201
rect 2912 13167 2946 13201
rect 2980 13167 3014 13201
rect 3048 13167 3082 13201
rect 3116 13167 3150 13201
rect 3184 13167 3218 13201
rect 3252 13167 3286 13201
rect 3320 13167 3354 13201
rect 3388 13167 3422 13201
rect 3456 13167 3574 13201
rect 3873 13711 3991 13745
rect 4025 13711 4059 13745
rect 4093 13711 4127 13745
rect 4161 13711 4195 13745
rect 4229 13711 4263 13745
rect 4297 13711 4331 13745
rect 4365 13711 4399 13745
rect 4433 13711 4467 13745
rect 4501 13711 4535 13745
rect 4569 13711 4603 13745
rect 4637 13711 4671 13745
rect 4705 13711 4739 13745
rect 4773 13711 4807 13745
rect 4841 13711 4875 13745
rect 4909 13711 4943 13745
rect 4977 13711 5095 13745
rect 3873 13643 3907 13711
rect 3873 13575 3907 13609
rect 5061 13643 5095 13711
rect 5061 13575 5095 13609
rect 3873 13507 3907 13541
rect 3873 13439 3907 13473
rect 3873 13371 3907 13405
rect 3873 13303 3907 13337
rect 5061 13507 5095 13541
rect 5061 13439 5095 13473
rect 5061 13371 5095 13405
rect 5061 13303 5095 13337
rect 3873 13201 3907 13269
rect 5061 13201 5095 13269
rect 3873 13167 3991 13201
rect 4025 13167 4059 13201
rect 4093 13167 4127 13201
rect 4161 13167 4195 13201
rect 4229 13167 4263 13201
rect 4297 13167 4331 13201
rect 4365 13167 4399 13201
rect 4433 13167 4467 13201
rect 4501 13167 4535 13201
rect 4569 13167 4603 13201
rect 4637 13167 4671 13201
rect 4705 13167 4739 13201
rect 4773 13167 4807 13201
rect 4841 13167 4875 13201
rect 4909 13167 4943 13201
rect 4977 13167 5095 13201
rect 199 12420 317 12454
rect 351 12420 385 12454
rect 419 12420 453 12454
rect 487 12420 521 12454
rect 555 12420 589 12454
rect 623 12420 657 12454
rect 691 12420 725 12454
rect 759 12420 793 12454
rect 827 12420 861 12454
rect 895 12420 929 12454
rect 963 12420 997 12454
rect 1031 12420 1065 12454
rect 1099 12420 1133 12454
rect 1167 12420 1201 12454
rect 1235 12420 1269 12454
rect 1303 12420 1421 12454
rect 199 12352 233 12420
rect 199 12284 233 12318
rect 1387 12352 1421 12420
rect 1387 12284 1421 12318
rect 199 12216 233 12250
rect 199 12148 233 12182
rect 199 12080 233 12114
rect 199 12012 233 12046
rect 1387 12216 1421 12250
rect 1387 12148 1421 12182
rect 1387 12080 1421 12114
rect 1387 12012 1421 12046
rect 199 11910 233 11978
rect 1387 11910 1421 11978
rect 199 11876 317 11910
rect 351 11876 385 11910
rect 419 11876 453 11910
rect 487 11876 521 11910
rect 555 11876 589 11910
rect 623 11876 657 11910
rect 691 11876 725 11910
rect 759 11876 793 11910
rect 827 11876 861 11910
rect 895 11876 929 11910
rect 963 11876 997 11910
rect 1031 11876 1065 11910
rect 1099 11876 1133 11910
rect 1167 11876 1201 11910
rect 1235 11876 1269 11910
rect 1303 11876 1421 11910
rect 2352 12424 2470 12458
rect 2504 12424 2538 12458
rect 2572 12424 2606 12458
rect 2640 12424 2674 12458
rect 2708 12424 2742 12458
rect 2776 12424 2810 12458
rect 2844 12424 2878 12458
rect 2912 12424 2946 12458
rect 2980 12424 3014 12458
rect 3048 12424 3082 12458
rect 3116 12424 3150 12458
rect 3184 12424 3218 12458
rect 3252 12424 3286 12458
rect 3320 12424 3354 12458
rect 3388 12424 3422 12458
rect 3456 12424 3574 12458
rect 2352 12356 2386 12424
rect 2352 12288 2386 12322
rect 3540 12356 3574 12424
rect 3540 12288 3574 12322
rect 2352 12220 2386 12254
rect 2352 12152 2386 12186
rect 2352 12084 2386 12118
rect 2352 12016 2386 12050
rect 3540 12220 3574 12254
rect 3540 12152 3574 12186
rect 3540 12084 3574 12118
rect 3540 12016 3574 12050
rect 2352 11914 2386 11982
rect 3540 11914 3574 11982
rect 2352 11880 2470 11914
rect 2504 11880 2538 11914
rect 2572 11880 2606 11914
rect 2640 11880 2674 11914
rect 2708 11880 2742 11914
rect 2776 11880 2810 11914
rect 2844 11880 2878 11914
rect 2912 11880 2946 11914
rect 2980 11880 3014 11914
rect 3048 11880 3082 11914
rect 3116 11880 3150 11914
rect 3184 11880 3218 11914
rect 3252 11880 3286 11914
rect 3320 11880 3354 11914
rect 3388 11880 3422 11914
rect 3456 11880 3574 11914
rect 3873 12424 3991 12458
rect 4025 12424 4059 12458
rect 4093 12424 4127 12458
rect 4161 12424 4195 12458
rect 4229 12424 4263 12458
rect 4297 12424 4331 12458
rect 4365 12424 4399 12458
rect 4433 12424 4467 12458
rect 4501 12424 4535 12458
rect 4569 12424 4603 12458
rect 4637 12424 4671 12458
rect 4705 12424 4739 12458
rect 4773 12424 4807 12458
rect 4841 12424 4875 12458
rect 4909 12424 4943 12458
rect 4977 12424 5095 12458
rect 3873 12356 3907 12424
rect 3873 12288 3907 12322
rect 5061 12356 5095 12424
rect 5061 12288 5095 12322
rect 3873 12220 3907 12254
rect 3873 12152 3907 12186
rect 3873 12084 3907 12118
rect 3873 12016 3907 12050
rect 5061 12220 5095 12254
rect 5061 12152 5095 12186
rect 5061 12084 5095 12118
rect 5061 12016 5095 12050
rect 3873 11914 3907 11982
rect 5061 11914 5095 11982
rect 3873 11880 3991 11914
rect 4025 11880 4059 11914
rect 4093 11880 4127 11914
rect 4161 11880 4195 11914
rect 4229 11880 4263 11914
rect 4297 11880 4331 11914
rect 4365 11880 4399 11914
rect 4433 11880 4467 11914
rect 4501 11880 4535 11914
rect 4569 11880 4603 11914
rect 4637 11880 4671 11914
rect 4705 11880 4739 11914
rect 4773 11880 4807 11914
rect 4841 11880 4875 11914
rect 4909 11880 4943 11914
rect 4977 11880 5095 11914
rect 199 11133 317 11167
rect 351 11133 385 11167
rect 419 11133 453 11167
rect 487 11133 521 11167
rect 555 11133 589 11167
rect 623 11133 657 11167
rect 691 11133 725 11167
rect 759 11133 793 11167
rect 827 11133 861 11167
rect 895 11133 929 11167
rect 963 11133 997 11167
rect 1031 11133 1065 11167
rect 1099 11133 1133 11167
rect 1167 11133 1201 11167
rect 1235 11133 1269 11167
rect 1303 11133 1421 11167
rect 199 11065 233 11133
rect 199 10997 233 11031
rect 1387 11065 1421 11133
rect 1387 10997 1421 11031
rect 199 10929 233 10963
rect 199 10861 233 10895
rect 199 10793 233 10827
rect 199 10725 233 10759
rect 1387 10929 1421 10963
rect 1387 10861 1421 10895
rect 1387 10793 1421 10827
rect 1387 10725 1421 10759
rect 199 10623 233 10691
rect 1387 10623 1421 10691
rect 199 10589 317 10623
rect 351 10589 385 10623
rect 419 10589 453 10623
rect 487 10589 521 10623
rect 555 10589 589 10623
rect 623 10589 657 10623
rect 691 10589 725 10623
rect 759 10589 793 10623
rect 827 10589 861 10623
rect 895 10589 929 10623
rect 963 10589 997 10623
rect 1031 10589 1065 10623
rect 1099 10589 1133 10623
rect 1167 10589 1201 10623
rect 1235 10589 1269 10623
rect 1303 10589 1421 10623
rect 2352 11137 2470 11171
rect 2504 11137 2538 11171
rect 2572 11137 2606 11171
rect 2640 11137 2674 11171
rect 2708 11137 2742 11171
rect 2776 11137 2810 11171
rect 2844 11137 2878 11171
rect 2912 11137 2946 11171
rect 2980 11137 3014 11171
rect 3048 11137 3082 11171
rect 3116 11137 3150 11171
rect 3184 11137 3218 11171
rect 3252 11137 3286 11171
rect 3320 11137 3354 11171
rect 3388 11137 3422 11171
rect 3456 11137 3574 11171
rect 2352 11069 2386 11137
rect 2352 11001 2386 11035
rect 3540 11069 3574 11137
rect 3540 11001 3574 11035
rect 2352 10933 2386 10967
rect 2352 10865 2386 10899
rect 2352 10797 2386 10831
rect 2352 10729 2386 10763
rect 3540 10933 3574 10967
rect 3540 10865 3574 10899
rect 3540 10797 3574 10831
rect 3540 10729 3574 10763
rect 2352 10627 2386 10695
rect 3540 10627 3574 10695
rect 2352 10593 2470 10627
rect 2504 10593 2538 10627
rect 2572 10593 2606 10627
rect 2640 10593 2674 10627
rect 2708 10593 2742 10627
rect 2776 10593 2810 10627
rect 2844 10593 2878 10627
rect 2912 10593 2946 10627
rect 2980 10593 3014 10627
rect 3048 10593 3082 10627
rect 3116 10593 3150 10627
rect 3184 10593 3218 10627
rect 3252 10593 3286 10627
rect 3320 10593 3354 10627
rect 3388 10593 3422 10627
rect 3456 10593 3574 10627
rect 3873 11137 3991 11171
rect 4025 11137 4059 11171
rect 4093 11137 4127 11171
rect 4161 11137 4195 11171
rect 4229 11137 4263 11171
rect 4297 11137 4331 11171
rect 4365 11137 4399 11171
rect 4433 11137 4467 11171
rect 4501 11137 4535 11171
rect 4569 11137 4603 11171
rect 4637 11137 4671 11171
rect 4705 11137 4739 11171
rect 4773 11137 4807 11171
rect 4841 11137 4875 11171
rect 4909 11137 4943 11171
rect 4977 11137 5095 11171
rect 3873 11069 3907 11137
rect 3873 11001 3907 11035
rect 5061 11069 5095 11137
rect 5061 11001 5095 11035
rect 3873 10933 3907 10967
rect 3873 10865 3907 10899
rect 3873 10797 3907 10831
rect 3873 10729 3907 10763
rect 5061 10933 5095 10967
rect 5061 10865 5095 10899
rect 5061 10797 5095 10831
rect 5061 10729 5095 10763
rect 3873 10627 3907 10695
rect 5061 10627 5095 10695
rect 3873 10593 3991 10627
rect 4025 10593 4059 10627
rect 4093 10593 4127 10627
rect 4161 10593 4195 10627
rect 4229 10593 4263 10627
rect 4297 10593 4331 10627
rect 4365 10593 4399 10627
rect 4433 10593 4467 10627
rect 4501 10593 4535 10627
rect 4569 10593 4603 10627
rect 4637 10593 4671 10627
rect 4705 10593 4739 10627
rect 4773 10593 4807 10627
rect 4841 10593 4875 10627
rect 4909 10593 4943 10627
rect 4977 10593 5095 10627
rect 199 9846 317 9880
rect 351 9846 385 9880
rect 419 9846 453 9880
rect 487 9846 521 9880
rect 555 9846 589 9880
rect 623 9846 657 9880
rect 691 9846 725 9880
rect 759 9846 793 9880
rect 827 9846 861 9880
rect 895 9846 929 9880
rect 963 9846 997 9880
rect 1031 9846 1065 9880
rect 1099 9846 1133 9880
rect 1167 9846 1201 9880
rect 1235 9846 1269 9880
rect 1303 9846 1421 9880
rect 199 9778 233 9846
rect 199 9710 233 9744
rect 1387 9778 1421 9846
rect 1387 9710 1421 9744
rect 199 9642 233 9676
rect 199 9574 233 9608
rect 199 9506 233 9540
rect 199 9438 233 9472
rect 1387 9642 1421 9676
rect 1387 9574 1421 9608
rect 1387 9506 1421 9540
rect 1387 9438 1421 9472
rect 199 9336 233 9404
rect 1387 9336 1421 9404
rect 199 9302 317 9336
rect 351 9302 385 9336
rect 419 9302 453 9336
rect 487 9302 521 9336
rect 555 9302 589 9336
rect 623 9302 657 9336
rect 691 9302 725 9336
rect 759 9302 793 9336
rect 827 9302 861 9336
rect 895 9302 929 9336
rect 963 9302 997 9336
rect 1031 9302 1065 9336
rect 1099 9302 1133 9336
rect 1167 9302 1201 9336
rect 1235 9302 1269 9336
rect 1303 9302 1421 9336
rect 2352 9850 2470 9884
rect 2504 9850 2538 9884
rect 2572 9850 2606 9884
rect 2640 9850 2674 9884
rect 2708 9850 2742 9884
rect 2776 9850 2810 9884
rect 2844 9850 2878 9884
rect 2912 9850 2946 9884
rect 2980 9850 3014 9884
rect 3048 9850 3082 9884
rect 3116 9850 3150 9884
rect 3184 9850 3218 9884
rect 3252 9850 3286 9884
rect 3320 9850 3354 9884
rect 3388 9850 3422 9884
rect 3456 9850 3574 9884
rect 2352 9782 2386 9850
rect 2352 9714 2386 9748
rect 3540 9782 3574 9850
rect 3540 9714 3574 9748
rect 2352 9646 2386 9680
rect 2352 9578 2386 9612
rect 2352 9510 2386 9544
rect 2352 9442 2386 9476
rect 3540 9646 3574 9680
rect 3540 9578 3574 9612
rect 3540 9510 3574 9544
rect 3540 9442 3574 9476
rect 2352 9340 2386 9408
rect 3540 9340 3574 9408
rect 2352 9306 2470 9340
rect 2504 9306 2538 9340
rect 2572 9306 2606 9340
rect 2640 9306 2674 9340
rect 2708 9306 2742 9340
rect 2776 9306 2810 9340
rect 2844 9306 2878 9340
rect 2912 9306 2946 9340
rect 2980 9306 3014 9340
rect 3048 9306 3082 9340
rect 3116 9306 3150 9340
rect 3184 9306 3218 9340
rect 3252 9306 3286 9340
rect 3320 9306 3354 9340
rect 3388 9306 3422 9340
rect 3456 9306 3574 9340
rect 3873 9850 3991 9884
rect 4025 9850 4059 9884
rect 4093 9850 4127 9884
rect 4161 9850 4195 9884
rect 4229 9850 4263 9884
rect 4297 9850 4331 9884
rect 4365 9850 4399 9884
rect 4433 9850 4467 9884
rect 4501 9850 4535 9884
rect 4569 9850 4603 9884
rect 4637 9850 4671 9884
rect 4705 9850 4739 9884
rect 4773 9850 4807 9884
rect 4841 9850 4875 9884
rect 4909 9850 4943 9884
rect 4977 9850 5095 9884
rect 3873 9782 3907 9850
rect 3873 9714 3907 9748
rect 5061 9782 5095 9850
rect 5061 9714 5095 9748
rect 3873 9646 3907 9680
rect 3873 9578 3907 9612
rect 3873 9510 3907 9544
rect 3873 9442 3907 9476
rect 5061 9646 5095 9680
rect 5061 9578 5095 9612
rect 5061 9510 5095 9544
rect 5061 9442 5095 9476
rect 3873 9340 3907 9408
rect 5061 9340 5095 9408
rect 3873 9306 3991 9340
rect 4025 9306 4059 9340
rect 4093 9306 4127 9340
rect 4161 9306 4195 9340
rect 4229 9306 4263 9340
rect 4297 9306 4331 9340
rect 4365 9306 4399 9340
rect 4433 9306 4467 9340
rect 4501 9306 4535 9340
rect 4569 9306 4603 9340
rect 4637 9306 4671 9340
rect 4705 9306 4739 9340
rect 4773 9306 4807 9340
rect 4841 9306 4875 9340
rect 4909 9306 4943 9340
rect 4977 9306 5095 9340
rect 199 8559 317 8593
rect 351 8559 385 8593
rect 419 8559 453 8593
rect 487 8559 521 8593
rect 555 8559 589 8593
rect 623 8559 657 8593
rect 691 8559 725 8593
rect 759 8559 793 8593
rect 827 8559 861 8593
rect 895 8559 929 8593
rect 963 8559 997 8593
rect 1031 8559 1065 8593
rect 1099 8559 1133 8593
rect 1167 8559 1201 8593
rect 1235 8559 1269 8593
rect 1303 8559 1421 8593
rect 199 8491 233 8559
rect 199 8423 233 8457
rect 1387 8491 1421 8559
rect 1387 8423 1421 8457
rect 199 8355 233 8389
rect 199 8287 233 8321
rect 199 8219 233 8253
rect 199 8151 233 8185
rect 1387 8355 1421 8389
rect 1387 8287 1421 8321
rect 1387 8219 1421 8253
rect 1387 8151 1421 8185
rect 199 8049 233 8117
rect 1387 8049 1421 8117
rect 199 8015 317 8049
rect 351 8015 385 8049
rect 419 8015 453 8049
rect 487 8015 521 8049
rect 555 8015 589 8049
rect 623 8015 657 8049
rect 691 8015 725 8049
rect 759 8015 793 8049
rect 827 8015 861 8049
rect 895 8015 929 8049
rect 963 8015 997 8049
rect 1031 8015 1065 8049
rect 1099 8015 1133 8049
rect 1167 8015 1201 8049
rect 1235 8015 1269 8049
rect 1303 8015 1421 8049
rect 2352 8563 2470 8597
rect 2504 8563 2538 8597
rect 2572 8563 2606 8597
rect 2640 8563 2674 8597
rect 2708 8563 2742 8597
rect 2776 8563 2810 8597
rect 2844 8563 2878 8597
rect 2912 8563 2946 8597
rect 2980 8563 3014 8597
rect 3048 8563 3082 8597
rect 3116 8563 3150 8597
rect 3184 8563 3218 8597
rect 3252 8563 3286 8597
rect 3320 8563 3354 8597
rect 3388 8563 3422 8597
rect 3456 8563 3574 8597
rect 2352 8495 2386 8563
rect 2352 8427 2386 8461
rect 3540 8495 3574 8563
rect 3540 8427 3574 8461
rect 2352 8359 2386 8393
rect 2352 8291 2386 8325
rect 2352 8223 2386 8257
rect 2352 8155 2386 8189
rect 3540 8359 3574 8393
rect 3540 8291 3574 8325
rect 3540 8223 3574 8257
rect 3540 8155 3574 8189
rect 2352 8053 2386 8121
rect 3540 8053 3574 8121
rect 2352 8019 2470 8053
rect 2504 8019 2538 8053
rect 2572 8019 2606 8053
rect 2640 8019 2674 8053
rect 2708 8019 2742 8053
rect 2776 8019 2810 8053
rect 2844 8019 2878 8053
rect 2912 8019 2946 8053
rect 2980 8019 3014 8053
rect 3048 8019 3082 8053
rect 3116 8019 3150 8053
rect 3184 8019 3218 8053
rect 3252 8019 3286 8053
rect 3320 8019 3354 8053
rect 3388 8019 3422 8053
rect 3456 8019 3574 8053
rect 3873 8563 3991 8597
rect 4025 8563 4059 8597
rect 4093 8563 4127 8597
rect 4161 8563 4195 8597
rect 4229 8563 4263 8597
rect 4297 8563 4331 8597
rect 4365 8563 4399 8597
rect 4433 8563 4467 8597
rect 4501 8563 4535 8597
rect 4569 8563 4603 8597
rect 4637 8563 4671 8597
rect 4705 8563 4739 8597
rect 4773 8563 4807 8597
rect 4841 8563 4875 8597
rect 4909 8563 4943 8597
rect 4977 8563 5095 8597
rect 3873 8495 3907 8563
rect 3873 8427 3907 8461
rect 5061 8495 5095 8563
rect 5061 8427 5095 8461
rect 3873 8359 3907 8393
rect 3873 8291 3907 8325
rect 3873 8223 3907 8257
rect 3873 8155 3907 8189
rect 5061 8359 5095 8393
rect 5061 8291 5095 8325
rect 5061 8223 5095 8257
rect 5061 8155 5095 8189
rect 3873 8053 3907 8121
rect 5061 8053 5095 8121
rect 3873 8019 3991 8053
rect 4025 8019 4059 8053
rect 4093 8019 4127 8053
rect 4161 8019 4195 8053
rect 4229 8019 4263 8053
rect 4297 8019 4331 8053
rect 4365 8019 4399 8053
rect 4433 8019 4467 8053
rect 4501 8019 4535 8053
rect 4569 8019 4603 8053
rect 4637 8019 4671 8053
rect 4705 8019 4739 8053
rect 4773 8019 4807 8053
rect 4841 8019 4875 8053
rect 4909 8019 4943 8053
rect 4977 8019 5095 8053
rect 199 7272 317 7306
rect 351 7272 385 7306
rect 419 7272 453 7306
rect 487 7272 521 7306
rect 555 7272 589 7306
rect 623 7272 657 7306
rect 691 7272 725 7306
rect 759 7272 793 7306
rect 827 7272 861 7306
rect 895 7272 929 7306
rect 963 7272 997 7306
rect 1031 7272 1065 7306
rect 1099 7272 1133 7306
rect 1167 7272 1201 7306
rect 1235 7272 1269 7306
rect 1303 7272 1421 7306
rect 199 7204 233 7272
rect 199 7136 233 7170
rect 1387 7204 1421 7272
rect 1387 7136 1421 7170
rect 199 7068 233 7102
rect 199 7000 233 7034
rect 199 6932 233 6966
rect 199 6864 233 6898
rect 1387 7068 1421 7102
rect 1387 7000 1421 7034
rect 1387 6932 1421 6966
rect 1387 6864 1421 6898
rect 199 6762 233 6830
rect 1387 6762 1421 6830
rect 199 6728 317 6762
rect 351 6728 385 6762
rect 419 6728 453 6762
rect 487 6728 521 6762
rect 555 6728 589 6762
rect 623 6728 657 6762
rect 691 6728 725 6762
rect 759 6728 793 6762
rect 827 6728 861 6762
rect 895 6728 929 6762
rect 963 6728 997 6762
rect 1031 6728 1065 6762
rect 1099 6728 1133 6762
rect 1167 6728 1201 6762
rect 1235 6728 1269 6762
rect 1303 6728 1421 6762
rect 2352 7276 2470 7310
rect 2504 7276 2538 7310
rect 2572 7276 2606 7310
rect 2640 7276 2674 7310
rect 2708 7276 2742 7310
rect 2776 7276 2810 7310
rect 2844 7276 2878 7310
rect 2912 7276 2946 7310
rect 2980 7276 3014 7310
rect 3048 7276 3082 7310
rect 3116 7276 3150 7310
rect 3184 7276 3218 7310
rect 3252 7276 3286 7310
rect 3320 7276 3354 7310
rect 3388 7276 3422 7310
rect 3456 7276 3574 7310
rect 2352 7208 2386 7276
rect 2352 7140 2386 7174
rect 3540 7208 3574 7276
rect 3540 7140 3574 7174
rect 2352 7072 2386 7106
rect 2352 7004 2386 7038
rect 2352 6936 2386 6970
rect 2352 6868 2386 6902
rect 3540 7072 3574 7106
rect 3540 7004 3574 7038
rect 3540 6936 3574 6970
rect 3540 6868 3574 6902
rect 2352 6766 2386 6834
rect 3540 6766 3574 6834
rect 2352 6732 2470 6766
rect 2504 6732 2538 6766
rect 2572 6732 2606 6766
rect 2640 6732 2674 6766
rect 2708 6732 2742 6766
rect 2776 6732 2810 6766
rect 2844 6732 2878 6766
rect 2912 6732 2946 6766
rect 2980 6732 3014 6766
rect 3048 6732 3082 6766
rect 3116 6732 3150 6766
rect 3184 6732 3218 6766
rect 3252 6732 3286 6766
rect 3320 6732 3354 6766
rect 3388 6732 3422 6766
rect 3456 6732 3574 6766
rect 3873 7276 3991 7310
rect 4025 7276 4059 7310
rect 4093 7276 4127 7310
rect 4161 7276 4195 7310
rect 4229 7276 4263 7310
rect 4297 7276 4331 7310
rect 4365 7276 4399 7310
rect 4433 7276 4467 7310
rect 4501 7276 4535 7310
rect 4569 7276 4603 7310
rect 4637 7276 4671 7310
rect 4705 7276 4739 7310
rect 4773 7276 4807 7310
rect 4841 7276 4875 7310
rect 4909 7276 4943 7310
rect 4977 7276 5095 7310
rect 3873 7208 3907 7276
rect 3873 7140 3907 7174
rect 5061 7208 5095 7276
rect 5061 7140 5095 7174
rect 3873 7072 3907 7106
rect 3873 7004 3907 7038
rect 3873 6936 3907 6970
rect 3873 6868 3907 6902
rect 5061 7072 5095 7106
rect 5061 7004 5095 7038
rect 5061 6936 5095 6970
rect 5061 6868 5095 6902
rect 3873 6766 3907 6834
rect 5061 6766 5095 6834
rect 3873 6732 3991 6766
rect 4025 6732 4059 6766
rect 4093 6732 4127 6766
rect 4161 6732 4195 6766
rect 4229 6732 4263 6766
rect 4297 6732 4331 6766
rect 4365 6732 4399 6766
rect 4433 6732 4467 6766
rect 4501 6732 4535 6766
rect 4569 6732 4603 6766
rect 4637 6732 4671 6766
rect 4705 6732 4739 6766
rect 4773 6732 4807 6766
rect 4841 6732 4875 6766
rect 4909 6732 4943 6766
rect 4977 6732 5095 6766
rect 199 5985 317 6019
rect 351 5985 385 6019
rect 419 5985 453 6019
rect 487 5985 521 6019
rect 555 5985 589 6019
rect 623 5985 657 6019
rect 691 5985 725 6019
rect 759 5985 793 6019
rect 827 5985 861 6019
rect 895 5985 929 6019
rect 963 5985 997 6019
rect 1031 5985 1065 6019
rect 1099 5985 1133 6019
rect 1167 5985 1201 6019
rect 1235 5985 1269 6019
rect 1303 5985 1421 6019
rect 199 5917 233 5985
rect 199 5849 233 5883
rect 1387 5917 1421 5985
rect 1387 5849 1421 5883
rect 199 5781 233 5815
rect 199 5713 233 5747
rect 199 5645 233 5679
rect 199 5577 233 5611
rect 1387 5781 1421 5815
rect 1387 5713 1421 5747
rect 1387 5645 1421 5679
rect 1387 5577 1421 5611
rect 199 5475 233 5543
rect 1387 5475 1421 5543
rect 199 5441 317 5475
rect 351 5441 385 5475
rect 419 5441 453 5475
rect 487 5441 521 5475
rect 555 5441 589 5475
rect 623 5441 657 5475
rect 691 5441 725 5475
rect 759 5441 793 5475
rect 827 5441 861 5475
rect 895 5441 929 5475
rect 963 5441 997 5475
rect 1031 5441 1065 5475
rect 1099 5441 1133 5475
rect 1167 5441 1201 5475
rect 1235 5441 1269 5475
rect 1303 5441 1421 5475
rect 2352 5989 2470 6023
rect 2504 5989 2538 6023
rect 2572 5989 2606 6023
rect 2640 5989 2674 6023
rect 2708 5989 2742 6023
rect 2776 5989 2810 6023
rect 2844 5989 2878 6023
rect 2912 5989 2946 6023
rect 2980 5989 3014 6023
rect 3048 5989 3082 6023
rect 3116 5989 3150 6023
rect 3184 5989 3218 6023
rect 3252 5989 3286 6023
rect 3320 5989 3354 6023
rect 3388 5989 3422 6023
rect 3456 5989 3574 6023
rect 2352 5921 2386 5989
rect 2352 5853 2386 5887
rect 3540 5921 3574 5989
rect 3540 5853 3574 5887
rect 2352 5785 2386 5819
rect 2352 5717 2386 5751
rect 2352 5649 2386 5683
rect 2352 5581 2386 5615
rect 3540 5785 3574 5819
rect 3540 5717 3574 5751
rect 3540 5649 3574 5683
rect 3540 5581 3574 5615
rect 2352 5479 2386 5547
rect 3540 5479 3574 5547
rect 2352 5445 2470 5479
rect 2504 5445 2538 5479
rect 2572 5445 2606 5479
rect 2640 5445 2674 5479
rect 2708 5445 2742 5479
rect 2776 5445 2810 5479
rect 2844 5445 2878 5479
rect 2912 5445 2946 5479
rect 2980 5445 3014 5479
rect 3048 5445 3082 5479
rect 3116 5445 3150 5479
rect 3184 5445 3218 5479
rect 3252 5445 3286 5479
rect 3320 5445 3354 5479
rect 3388 5445 3422 5479
rect 3456 5445 3574 5479
rect 3873 5989 3991 6023
rect 4025 5989 4059 6023
rect 4093 5989 4127 6023
rect 4161 5989 4195 6023
rect 4229 5989 4263 6023
rect 4297 5989 4331 6023
rect 4365 5989 4399 6023
rect 4433 5989 4467 6023
rect 4501 5989 4535 6023
rect 4569 5989 4603 6023
rect 4637 5989 4671 6023
rect 4705 5989 4739 6023
rect 4773 5989 4807 6023
rect 4841 5989 4875 6023
rect 4909 5989 4943 6023
rect 4977 5989 5095 6023
rect 3873 5921 3907 5989
rect 3873 5853 3907 5887
rect 5061 5921 5095 5989
rect 5061 5853 5095 5887
rect 3873 5785 3907 5819
rect 3873 5717 3907 5751
rect 3873 5649 3907 5683
rect 3873 5581 3907 5615
rect 5061 5785 5095 5819
rect 5061 5717 5095 5751
rect 5061 5649 5095 5683
rect 5061 5581 5095 5615
rect 3873 5479 3907 5547
rect 5061 5479 5095 5547
rect 3873 5445 3991 5479
rect 4025 5445 4059 5479
rect 4093 5445 4127 5479
rect 4161 5445 4195 5479
rect 4229 5445 4263 5479
rect 4297 5445 4331 5479
rect 4365 5445 4399 5479
rect 4433 5445 4467 5479
rect 4501 5445 4535 5479
rect 4569 5445 4603 5479
rect 4637 5445 4671 5479
rect 4705 5445 4739 5479
rect 4773 5445 4807 5479
rect 4841 5445 4875 5479
rect 4909 5445 4943 5479
rect 4977 5445 5095 5479
rect 199 4698 317 4732
rect 351 4698 385 4732
rect 419 4698 453 4732
rect 487 4698 521 4732
rect 555 4698 589 4732
rect 623 4698 657 4732
rect 691 4698 725 4732
rect 759 4698 793 4732
rect 827 4698 861 4732
rect 895 4698 929 4732
rect 963 4698 997 4732
rect 1031 4698 1065 4732
rect 1099 4698 1133 4732
rect 1167 4698 1201 4732
rect 1235 4698 1269 4732
rect 1303 4698 1421 4732
rect 199 4630 233 4698
rect 199 4562 233 4596
rect 1387 4630 1421 4698
rect 1387 4562 1421 4596
rect 199 4494 233 4528
rect 199 4426 233 4460
rect 199 4358 233 4392
rect 199 4290 233 4324
rect 1387 4494 1421 4528
rect 1387 4426 1421 4460
rect 1387 4358 1421 4392
rect 1387 4290 1421 4324
rect 199 4188 233 4256
rect 1387 4188 1421 4256
rect 199 4154 317 4188
rect 351 4154 385 4188
rect 419 4154 453 4188
rect 487 4154 521 4188
rect 555 4154 589 4188
rect 623 4154 657 4188
rect 691 4154 725 4188
rect 759 4154 793 4188
rect 827 4154 861 4188
rect 895 4154 929 4188
rect 963 4154 997 4188
rect 1031 4154 1065 4188
rect 1099 4154 1133 4188
rect 1167 4154 1201 4188
rect 1235 4154 1269 4188
rect 1303 4154 1421 4188
rect 2352 4702 2470 4736
rect 2504 4702 2538 4736
rect 2572 4702 2606 4736
rect 2640 4702 2674 4736
rect 2708 4702 2742 4736
rect 2776 4702 2810 4736
rect 2844 4702 2878 4736
rect 2912 4702 2946 4736
rect 2980 4702 3014 4736
rect 3048 4702 3082 4736
rect 3116 4702 3150 4736
rect 3184 4702 3218 4736
rect 3252 4702 3286 4736
rect 3320 4702 3354 4736
rect 3388 4702 3422 4736
rect 3456 4702 3574 4736
rect 2352 4634 2386 4702
rect 2352 4566 2386 4600
rect 3540 4634 3574 4702
rect 3540 4566 3574 4600
rect 2352 4498 2386 4532
rect 2352 4430 2386 4464
rect 2352 4362 2386 4396
rect 2352 4294 2386 4328
rect 3540 4498 3574 4532
rect 3540 4430 3574 4464
rect 3540 4362 3574 4396
rect 3540 4294 3574 4328
rect 2352 4192 2386 4260
rect 3540 4192 3574 4260
rect 2352 4158 2470 4192
rect 2504 4158 2538 4192
rect 2572 4158 2606 4192
rect 2640 4158 2674 4192
rect 2708 4158 2742 4192
rect 2776 4158 2810 4192
rect 2844 4158 2878 4192
rect 2912 4158 2946 4192
rect 2980 4158 3014 4192
rect 3048 4158 3082 4192
rect 3116 4158 3150 4192
rect 3184 4158 3218 4192
rect 3252 4158 3286 4192
rect 3320 4158 3354 4192
rect 3388 4158 3422 4192
rect 3456 4158 3574 4192
rect 3873 4702 3991 4736
rect 4025 4702 4059 4736
rect 4093 4702 4127 4736
rect 4161 4702 4195 4736
rect 4229 4702 4263 4736
rect 4297 4702 4331 4736
rect 4365 4702 4399 4736
rect 4433 4702 4467 4736
rect 4501 4702 4535 4736
rect 4569 4702 4603 4736
rect 4637 4702 4671 4736
rect 4705 4702 4739 4736
rect 4773 4702 4807 4736
rect 4841 4702 4875 4736
rect 4909 4702 4943 4736
rect 4977 4702 5095 4736
rect 3873 4634 3907 4702
rect 3873 4566 3907 4600
rect 5061 4634 5095 4702
rect 5061 4566 5095 4600
rect 3873 4498 3907 4532
rect 3873 4430 3907 4464
rect 3873 4362 3907 4396
rect 3873 4294 3907 4328
rect 5061 4498 5095 4532
rect 5061 4430 5095 4464
rect 5061 4362 5095 4396
rect 5061 4294 5095 4328
rect 3873 4192 3907 4260
rect 5061 4192 5095 4260
rect 3873 4158 3991 4192
rect 4025 4158 4059 4192
rect 4093 4158 4127 4192
rect 4161 4158 4195 4192
rect 4229 4158 4263 4192
rect 4297 4158 4331 4192
rect 4365 4158 4399 4192
rect 4433 4158 4467 4192
rect 4501 4158 4535 4192
rect 4569 4158 4603 4192
rect 4637 4158 4671 4192
rect 4705 4158 4739 4192
rect 4773 4158 4807 4192
rect 4841 4158 4875 4192
rect 4909 4158 4943 4192
rect 4977 4158 5095 4192
rect 199 3411 317 3445
rect 351 3411 385 3445
rect 419 3411 453 3445
rect 487 3411 521 3445
rect 555 3411 589 3445
rect 623 3411 657 3445
rect 691 3411 725 3445
rect 759 3411 793 3445
rect 827 3411 861 3445
rect 895 3411 929 3445
rect 963 3411 997 3445
rect 1031 3411 1065 3445
rect 1099 3411 1133 3445
rect 1167 3411 1201 3445
rect 1235 3411 1269 3445
rect 1303 3411 1421 3445
rect 199 3343 233 3411
rect 199 3275 233 3309
rect 1387 3343 1421 3411
rect 1387 3275 1421 3309
rect 199 3207 233 3241
rect 199 3139 233 3173
rect 199 3071 233 3105
rect 199 3003 233 3037
rect 1387 3207 1421 3241
rect 1387 3139 1421 3173
rect 1387 3071 1421 3105
rect 1387 3003 1421 3037
rect 199 2901 233 2969
rect 1387 2901 1421 2969
rect 199 2867 317 2901
rect 351 2867 385 2901
rect 419 2867 453 2901
rect 487 2867 521 2901
rect 555 2867 589 2901
rect 623 2867 657 2901
rect 691 2867 725 2901
rect 759 2867 793 2901
rect 827 2867 861 2901
rect 895 2867 929 2901
rect 963 2867 997 2901
rect 1031 2867 1065 2901
rect 1099 2867 1133 2901
rect 1167 2867 1201 2901
rect 1235 2867 1269 2901
rect 1303 2867 1421 2901
rect 2352 3415 2470 3449
rect 2504 3415 2538 3449
rect 2572 3415 2606 3449
rect 2640 3415 2674 3449
rect 2708 3415 2742 3449
rect 2776 3415 2810 3449
rect 2844 3415 2878 3449
rect 2912 3415 2946 3449
rect 2980 3415 3014 3449
rect 3048 3415 3082 3449
rect 3116 3415 3150 3449
rect 3184 3415 3218 3449
rect 3252 3415 3286 3449
rect 3320 3415 3354 3449
rect 3388 3415 3422 3449
rect 3456 3415 3574 3449
rect 2352 3347 2386 3415
rect 2352 3279 2386 3313
rect 3540 3347 3574 3415
rect 3540 3279 3574 3313
rect 2352 3211 2386 3245
rect 2352 3143 2386 3177
rect 2352 3075 2386 3109
rect 2352 3007 2386 3041
rect 3540 3211 3574 3245
rect 3540 3143 3574 3177
rect 3540 3075 3574 3109
rect 3540 3007 3574 3041
rect 2352 2905 2386 2973
rect 3540 2905 3574 2973
rect 2352 2871 2470 2905
rect 2504 2871 2538 2905
rect 2572 2871 2606 2905
rect 2640 2871 2674 2905
rect 2708 2871 2742 2905
rect 2776 2871 2810 2905
rect 2844 2871 2878 2905
rect 2912 2871 2946 2905
rect 2980 2871 3014 2905
rect 3048 2871 3082 2905
rect 3116 2871 3150 2905
rect 3184 2871 3218 2905
rect 3252 2871 3286 2905
rect 3320 2871 3354 2905
rect 3388 2871 3422 2905
rect 3456 2871 3574 2905
rect 3873 3415 3991 3449
rect 4025 3415 4059 3449
rect 4093 3415 4127 3449
rect 4161 3415 4195 3449
rect 4229 3415 4263 3449
rect 4297 3415 4331 3449
rect 4365 3415 4399 3449
rect 4433 3415 4467 3449
rect 4501 3415 4535 3449
rect 4569 3415 4603 3449
rect 4637 3415 4671 3449
rect 4705 3415 4739 3449
rect 4773 3415 4807 3449
rect 4841 3415 4875 3449
rect 4909 3415 4943 3449
rect 4977 3415 5095 3449
rect 3873 3347 3907 3415
rect 3873 3279 3907 3313
rect 5061 3347 5095 3415
rect 5061 3279 5095 3313
rect 3873 3211 3907 3245
rect 3873 3143 3907 3177
rect 3873 3075 3907 3109
rect 3873 3007 3907 3041
rect 5061 3211 5095 3245
rect 5061 3143 5095 3177
rect 5061 3075 5095 3109
rect 5061 3007 5095 3041
rect 3873 2905 3907 2973
rect 5061 2905 5095 2973
rect 3873 2871 3991 2905
rect 4025 2871 4059 2905
rect 4093 2871 4127 2905
rect 4161 2871 4195 2905
rect 4229 2871 4263 2905
rect 4297 2871 4331 2905
rect 4365 2871 4399 2905
rect 4433 2871 4467 2905
rect 4501 2871 4535 2905
rect 4569 2871 4603 2905
rect 4637 2871 4671 2905
rect 4705 2871 4739 2905
rect 4773 2871 4807 2905
rect 4841 2871 4875 2905
rect 4909 2871 4943 2905
rect 4977 2871 5095 2905
rect 199 2124 317 2158
rect 351 2124 385 2158
rect 419 2124 453 2158
rect 487 2124 521 2158
rect 555 2124 589 2158
rect 623 2124 657 2158
rect 691 2124 725 2158
rect 759 2124 793 2158
rect 827 2124 861 2158
rect 895 2124 929 2158
rect 963 2124 997 2158
rect 1031 2124 1065 2158
rect 1099 2124 1133 2158
rect 1167 2124 1201 2158
rect 1235 2124 1269 2158
rect 1303 2124 1421 2158
rect 199 2056 233 2124
rect 199 1988 233 2022
rect 1387 2056 1421 2124
rect 1387 1988 1421 2022
rect 199 1920 233 1954
rect 199 1852 233 1886
rect 199 1784 233 1818
rect 199 1716 233 1750
rect 1387 1920 1421 1954
rect 1387 1852 1421 1886
rect 1387 1784 1421 1818
rect 1387 1716 1421 1750
rect 199 1614 233 1682
rect 1387 1614 1421 1682
rect 199 1580 317 1614
rect 351 1580 385 1614
rect 419 1580 453 1614
rect 487 1580 521 1614
rect 555 1580 589 1614
rect 623 1580 657 1614
rect 691 1580 725 1614
rect 759 1580 793 1614
rect 827 1580 861 1614
rect 895 1580 929 1614
rect 963 1580 997 1614
rect 1031 1580 1065 1614
rect 1099 1580 1133 1614
rect 1167 1580 1201 1614
rect 1235 1580 1269 1614
rect 1303 1580 1421 1614
rect 2352 2128 2470 2162
rect 2504 2128 2538 2162
rect 2572 2128 2606 2162
rect 2640 2128 2674 2162
rect 2708 2128 2742 2162
rect 2776 2128 2810 2162
rect 2844 2128 2878 2162
rect 2912 2128 2946 2162
rect 2980 2128 3014 2162
rect 3048 2128 3082 2162
rect 3116 2128 3150 2162
rect 3184 2128 3218 2162
rect 3252 2128 3286 2162
rect 3320 2128 3354 2162
rect 3388 2128 3422 2162
rect 3456 2128 3574 2162
rect 2352 2060 2386 2128
rect 2352 1992 2386 2026
rect 3540 2060 3574 2128
rect 3540 1992 3574 2026
rect 2352 1924 2386 1958
rect 2352 1856 2386 1890
rect 2352 1788 2386 1822
rect 2352 1720 2386 1754
rect 3540 1924 3574 1958
rect 3540 1856 3574 1890
rect 3540 1788 3574 1822
rect 3540 1720 3574 1754
rect 2352 1618 2386 1686
rect 3540 1618 3574 1686
rect 2352 1584 2470 1618
rect 2504 1584 2538 1618
rect 2572 1584 2606 1618
rect 2640 1584 2674 1618
rect 2708 1584 2742 1618
rect 2776 1584 2810 1618
rect 2844 1584 2878 1618
rect 2912 1584 2946 1618
rect 2980 1584 3014 1618
rect 3048 1584 3082 1618
rect 3116 1584 3150 1618
rect 3184 1584 3218 1618
rect 3252 1584 3286 1618
rect 3320 1584 3354 1618
rect 3388 1584 3422 1618
rect 3456 1584 3574 1618
rect 3873 2128 3991 2162
rect 4025 2128 4059 2162
rect 4093 2128 4127 2162
rect 4161 2128 4195 2162
rect 4229 2128 4263 2162
rect 4297 2128 4331 2162
rect 4365 2128 4399 2162
rect 4433 2128 4467 2162
rect 4501 2128 4535 2162
rect 4569 2128 4603 2162
rect 4637 2128 4671 2162
rect 4705 2128 4739 2162
rect 4773 2128 4807 2162
rect 4841 2128 4875 2162
rect 4909 2128 4943 2162
rect 4977 2128 5095 2162
rect 3873 2060 3907 2128
rect 3873 1992 3907 2026
rect 5061 2060 5095 2128
rect 5061 1992 5095 2026
rect 3873 1924 3907 1958
rect 3873 1856 3907 1890
rect 3873 1788 3907 1822
rect 3873 1720 3907 1754
rect 5061 1924 5095 1958
rect 5061 1856 5095 1890
rect 5061 1788 5095 1822
rect 5061 1720 5095 1754
rect 3873 1618 3907 1686
rect 5061 1618 5095 1686
rect 3873 1584 3991 1618
rect 4025 1584 4059 1618
rect 4093 1584 4127 1618
rect 4161 1584 4195 1618
rect 4229 1584 4263 1618
rect 4297 1584 4331 1618
rect 4365 1584 4399 1618
rect 4433 1584 4467 1618
rect 4501 1584 4535 1618
rect 4569 1584 4603 1618
rect 4637 1584 4671 1618
rect 4705 1584 4739 1618
rect 4773 1584 4807 1618
rect 4841 1584 4875 1618
rect 4909 1584 4943 1618
rect 4977 1584 5095 1618
<< psubdiffcont >>
rect 317 41369 351 41403
rect 385 41369 419 41403
rect 453 41369 487 41403
rect 521 41369 555 41403
rect 589 41369 623 41403
rect 657 41369 691 41403
rect 725 41369 759 41403
rect 793 41369 827 41403
rect 861 41369 895 41403
rect 929 41369 963 41403
rect 997 41369 1031 41403
rect 1065 41369 1099 41403
rect 1133 41369 1167 41403
rect 1201 41369 1235 41403
rect 1269 41369 1303 41403
rect 199 41259 233 41293
rect 199 41191 233 41225
rect 1387 41259 1421 41293
rect 1387 41191 1421 41225
rect 199 41123 233 41157
rect 1387 41123 1421 41157
rect 317 41013 351 41047
rect 385 41013 419 41047
rect 453 41013 487 41047
rect 521 41013 555 41047
rect 589 41013 623 41047
rect 657 41013 691 41047
rect 725 41013 759 41047
rect 793 41013 827 41047
rect 861 41013 895 41047
rect 929 41013 963 41047
rect 997 41013 1031 41047
rect 1065 41013 1099 41047
rect 1133 41013 1167 41047
rect 1201 41013 1235 41047
rect 1269 41013 1303 41047
rect 2470 41373 2504 41407
rect 2538 41373 2572 41407
rect 2606 41373 2640 41407
rect 2674 41373 2708 41407
rect 2742 41373 2776 41407
rect 2810 41373 2844 41407
rect 2878 41373 2912 41407
rect 2946 41373 2980 41407
rect 3014 41373 3048 41407
rect 3082 41373 3116 41407
rect 3150 41373 3184 41407
rect 3218 41373 3252 41407
rect 3286 41373 3320 41407
rect 3354 41373 3388 41407
rect 3422 41373 3456 41407
rect 2352 41263 2386 41297
rect 3991 41373 4025 41407
rect 4059 41373 4093 41407
rect 4127 41373 4161 41407
rect 4195 41373 4229 41407
rect 4263 41373 4297 41407
rect 4331 41373 4365 41407
rect 4399 41373 4433 41407
rect 4467 41373 4501 41407
rect 4535 41373 4569 41407
rect 4603 41373 4637 41407
rect 4671 41373 4705 41407
rect 4739 41373 4773 41407
rect 4807 41373 4841 41407
rect 4875 41373 4909 41407
rect 4943 41373 4977 41407
rect 2352 41195 2386 41229
rect 3540 41263 3574 41297
rect 3540 41195 3574 41229
rect 3873 41263 3907 41297
rect 2352 41127 2386 41161
rect 3873 41195 3907 41229
rect 3540 41127 3574 41161
rect 2470 41017 2504 41051
rect 2538 41017 2572 41051
rect 2606 41017 2640 41051
rect 2674 41017 2708 41051
rect 2742 41017 2776 41051
rect 2810 41017 2844 41051
rect 2878 41017 2912 41051
rect 2946 41017 2980 41051
rect 3014 41017 3048 41051
rect 3082 41017 3116 41051
rect 3150 41017 3184 41051
rect 3218 41017 3252 41051
rect 3286 41017 3320 41051
rect 3354 41017 3388 41051
rect 3422 41017 3456 41051
rect 5061 41263 5095 41297
rect 5061 41195 5095 41229
rect 3873 41127 3907 41161
rect 5061 41127 5095 41161
rect 3991 41017 4025 41051
rect 4059 41017 4093 41051
rect 4127 41017 4161 41051
rect 4195 41017 4229 41051
rect 4263 41017 4297 41051
rect 4331 41017 4365 41051
rect 4399 41017 4433 41051
rect 4467 41017 4501 41051
rect 4535 41017 4569 41051
rect 4603 41017 4637 41051
rect 4671 41017 4705 41051
rect 4739 41017 4773 41051
rect 4807 41017 4841 41051
rect 4875 41017 4909 41051
rect 4943 41017 4977 41051
rect 317 40082 351 40116
rect 385 40082 419 40116
rect 453 40082 487 40116
rect 521 40082 555 40116
rect 589 40082 623 40116
rect 657 40082 691 40116
rect 725 40082 759 40116
rect 793 40082 827 40116
rect 861 40082 895 40116
rect 929 40082 963 40116
rect 997 40082 1031 40116
rect 1065 40082 1099 40116
rect 1133 40082 1167 40116
rect 1201 40082 1235 40116
rect 1269 40082 1303 40116
rect 199 39972 233 40006
rect 199 39904 233 39938
rect 1387 39972 1421 40006
rect 1387 39904 1421 39938
rect 199 39836 233 39870
rect 1387 39836 1421 39870
rect 317 39726 351 39760
rect 385 39726 419 39760
rect 453 39726 487 39760
rect 521 39726 555 39760
rect 589 39726 623 39760
rect 657 39726 691 39760
rect 725 39726 759 39760
rect 793 39726 827 39760
rect 861 39726 895 39760
rect 929 39726 963 39760
rect 997 39726 1031 39760
rect 1065 39726 1099 39760
rect 1133 39726 1167 39760
rect 1201 39726 1235 39760
rect 1269 39726 1303 39760
rect 2470 40086 2504 40120
rect 2538 40086 2572 40120
rect 2606 40086 2640 40120
rect 2674 40086 2708 40120
rect 2742 40086 2776 40120
rect 2810 40086 2844 40120
rect 2878 40086 2912 40120
rect 2946 40086 2980 40120
rect 3014 40086 3048 40120
rect 3082 40086 3116 40120
rect 3150 40086 3184 40120
rect 3218 40086 3252 40120
rect 3286 40086 3320 40120
rect 3354 40086 3388 40120
rect 3422 40086 3456 40120
rect 2352 39976 2386 40010
rect 3991 40086 4025 40120
rect 4059 40086 4093 40120
rect 4127 40086 4161 40120
rect 4195 40086 4229 40120
rect 4263 40086 4297 40120
rect 4331 40086 4365 40120
rect 4399 40086 4433 40120
rect 4467 40086 4501 40120
rect 4535 40086 4569 40120
rect 4603 40086 4637 40120
rect 4671 40086 4705 40120
rect 4739 40086 4773 40120
rect 4807 40086 4841 40120
rect 4875 40086 4909 40120
rect 4943 40086 4977 40120
rect 2352 39908 2386 39942
rect 3540 39976 3574 40010
rect 3540 39908 3574 39942
rect 3873 39976 3907 40010
rect 2352 39840 2386 39874
rect 3873 39908 3907 39942
rect 3540 39840 3574 39874
rect 2470 39730 2504 39764
rect 2538 39730 2572 39764
rect 2606 39730 2640 39764
rect 2674 39730 2708 39764
rect 2742 39730 2776 39764
rect 2810 39730 2844 39764
rect 2878 39730 2912 39764
rect 2946 39730 2980 39764
rect 3014 39730 3048 39764
rect 3082 39730 3116 39764
rect 3150 39730 3184 39764
rect 3218 39730 3252 39764
rect 3286 39730 3320 39764
rect 3354 39730 3388 39764
rect 3422 39730 3456 39764
rect 5061 39976 5095 40010
rect 5061 39908 5095 39942
rect 3873 39840 3907 39874
rect 5061 39840 5095 39874
rect 3991 39730 4025 39764
rect 4059 39730 4093 39764
rect 4127 39730 4161 39764
rect 4195 39730 4229 39764
rect 4263 39730 4297 39764
rect 4331 39730 4365 39764
rect 4399 39730 4433 39764
rect 4467 39730 4501 39764
rect 4535 39730 4569 39764
rect 4603 39730 4637 39764
rect 4671 39730 4705 39764
rect 4739 39730 4773 39764
rect 4807 39730 4841 39764
rect 4875 39730 4909 39764
rect 4943 39730 4977 39764
rect 317 38795 351 38829
rect 385 38795 419 38829
rect 453 38795 487 38829
rect 521 38795 555 38829
rect 589 38795 623 38829
rect 657 38795 691 38829
rect 725 38795 759 38829
rect 793 38795 827 38829
rect 861 38795 895 38829
rect 929 38795 963 38829
rect 997 38795 1031 38829
rect 1065 38795 1099 38829
rect 1133 38795 1167 38829
rect 1201 38795 1235 38829
rect 1269 38795 1303 38829
rect 199 38685 233 38719
rect 199 38617 233 38651
rect 1387 38685 1421 38719
rect 1387 38617 1421 38651
rect 199 38549 233 38583
rect 1387 38549 1421 38583
rect 317 38439 351 38473
rect 385 38439 419 38473
rect 453 38439 487 38473
rect 521 38439 555 38473
rect 589 38439 623 38473
rect 657 38439 691 38473
rect 725 38439 759 38473
rect 793 38439 827 38473
rect 861 38439 895 38473
rect 929 38439 963 38473
rect 997 38439 1031 38473
rect 1065 38439 1099 38473
rect 1133 38439 1167 38473
rect 1201 38439 1235 38473
rect 1269 38439 1303 38473
rect 2470 38799 2504 38833
rect 2538 38799 2572 38833
rect 2606 38799 2640 38833
rect 2674 38799 2708 38833
rect 2742 38799 2776 38833
rect 2810 38799 2844 38833
rect 2878 38799 2912 38833
rect 2946 38799 2980 38833
rect 3014 38799 3048 38833
rect 3082 38799 3116 38833
rect 3150 38799 3184 38833
rect 3218 38799 3252 38833
rect 3286 38799 3320 38833
rect 3354 38799 3388 38833
rect 3422 38799 3456 38833
rect 2352 38689 2386 38723
rect 3991 38799 4025 38833
rect 4059 38799 4093 38833
rect 4127 38799 4161 38833
rect 4195 38799 4229 38833
rect 4263 38799 4297 38833
rect 4331 38799 4365 38833
rect 4399 38799 4433 38833
rect 4467 38799 4501 38833
rect 4535 38799 4569 38833
rect 4603 38799 4637 38833
rect 4671 38799 4705 38833
rect 4739 38799 4773 38833
rect 4807 38799 4841 38833
rect 4875 38799 4909 38833
rect 4943 38799 4977 38833
rect 2352 38621 2386 38655
rect 3540 38689 3574 38723
rect 3540 38621 3574 38655
rect 3873 38689 3907 38723
rect 2352 38553 2386 38587
rect 3873 38621 3907 38655
rect 3540 38553 3574 38587
rect 2470 38443 2504 38477
rect 2538 38443 2572 38477
rect 2606 38443 2640 38477
rect 2674 38443 2708 38477
rect 2742 38443 2776 38477
rect 2810 38443 2844 38477
rect 2878 38443 2912 38477
rect 2946 38443 2980 38477
rect 3014 38443 3048 38477
rect 3082 38443 3116 38477
rect 3150 38443 3184 38477
rect 3218 38443 3252 38477
rect 3286 38443 3320 38477
rect 3354 38443 3388 38477
rect 3422 38443 3456 38477
rect 5061 38689 5095 38723
rect 5061 38621 5095 38655
rect 3873 38553 3907 38587
rect 5061 38553 5095 38587
rect 3991 38443 4025 38477
rect 4059 38443 4093 38477
rect 4127 38443 4161 38477
rect 4195 38443 4229 38477
rect 4263 38443 4297 38477
rect 4331 38443 4365 38477
rect 4399 38443 4433 38477
rect 4467 38443 4501 38477
rect 4535 38443 4569 38477
rect 4603 38443 4637 38477
rect 4671 38443 4705 38477
rect 4739 38443 4773 38477
rect 4807 38443 4841 38477
rect 4875 38443 4909 38477
rect 4943 38443 4977 38477
rect 317 37508 351 37542
rect 385 37508 419 37542
rect 453 37508 487 37542
rect 521 37508 555 37542
rect 589 37508 623 37542
rect 657 37508 691 37542
rect 725 37508 759 37542
rect 793 37508 827 37542
rect 861 37508 895 37542
rect 929 37508 963 37542
rect 997 37508 1031 37542
rect 1065 37508 1099 37542
rect 1133 37508 1167 37542
rect 1201 37508 1235 37542
rect 1269 37508 1303 37542
rect 199 37398 233 37432
rect 199 37330 233 37364
rect 1387 37398 1421 37432
rect 1387 37330 1421 37364
rect 199 37262 233 37296
rect 1387 37262 1421 37296
rect 317 37152 351 37186
rect 385 37152 419 37186
rect 453 37152 487 37186
rect 521 37152 555 37186
rect 589 37152 623 37186
rect 657 37152 691 37186
rect 725 37152 759 37186
rect 793 37152 827 37186
rect 861 37152 895 37186
rect 929 37152 963 37186
rect 997 37152 1031 37186
rect 1065 37152 1099 37186
rect 1133 37152 1167 37186
rect 1201 37152 1235 37186
rect 1269 37152 1303 37186
rect 2470 37512 2504 37546
rect 2538 37512 2572 37546
rect 2606 37512 2640 37546
rect 2674 37512 2708 37546
rect 2742 37512 2776 37546
rect 2810 37512 2844 37546
rect 2878 37512 2912 37546
rect 2946 37512 2980 37546
rect 3014 37512 3048 37546
rect 3082 37512 3116 37546
rect 3150 37512 3184 37546
rect 3218 37512 3252 37546
rect 3286 37512 3320 37546
rect 3354 37512 3388 37546
rect 3422 37512 3456 37546
rect 2352 37402 2386 37436
rect 3991 37512 4025 37546
rect 4059 37512 4093 37546
rect 4127 37512 4161 37546
rect 4195 37512 4229 37546
rect 4263 37512 4297 37546
rect 4331 37512 4365 37546
rect 4399 37512 4433 37546
rect 4467 37512 4501 37546
rect 4535 37512 4569 37546
rect 4603 37512 4637 37546
rect 4671 37512 4705 37546
rect 4739 37512 4773 37546
rect 4807 37512 4841 37546
rect 4875 37512 4909 37546
rect 4943 37512 4977 37546
rect 2352 37334 2386 37368
rect 3540 37402 3574 37436
rect 3540 37334 3574 37368
rect 3873 37402 3907 37436
rect 2352 37266 2386 37300
rect 3873 37334 3907 37368
rect 3540 37266 3574 37300
rect 2470 37156 2504 37190
rect 2538 37156 2572 37190
rect 2606 37156 2640 37190
rect 2674 37156 2708 37190
rect 2742 37156 2776 37190
rect 2810 37156 2844 37190
rect 2878 37156 2912 37190
rect 2946 37156 2980 37190
rect 3014 37156 3048 37190
rect 3082 37156 3116 37190
rect 3150 37156 3184 37190
rect 3218 37156 3252 37190
rect 3286 37156 3320 37190
rect 3354 37156 3388 37190
rect 3422 37156 3456 37190
rect 5061 37402 5095 37436
rect 5061 37334 5095 37368
rect 3873 37266 3907 37300
rect 5061 37266 5095 37300
rect 3991 37156 4025 37190
rect 4059 37156 4093 37190
rect 4127 37156 4161 37190
rect 4195 37156 4229 37190
rect 4263 37156 4297 37190
rect 4331 37156 4365 37190
rect 4399 37156 4433 37190
rect 4467 37156 4501 37190
rect 4535 37156 4569 37190
rect 4603 37156 4637 37190
rect 4671 37156 4705 37190
rect 4739 37156 4773 37190
rect 4807 37156 4841 37190
rect 4875 37156 4909 37190
rect 4943 37156 4977 37190
rect 317 36221 351 36255
rect 385 36221 419 36255
rect 453 36221 487 36255
rect 521 36221 555 36255
rect 589 36221 623 36255
rect 657 36221 691 36255
rect 725 36221 759 36255
rect 793 36221 827 36255
rect 861 36221 895 36255
rect 929 36221 963 36255
rect 997 36221 1031 36255
rect 1065 36221 1099 36255
rect 1133 36221 1167 36255
rect 1201 36221 1235 36255
rect 1269 36221 1303 36255
rect 199 36111 233 36145
rect 199 36043 233 36077
rect 1387 36111 1421 36145
rect 1387 36043 1421 36077
rect 199 35975 233 36009
rect 1387 35975 1421 36009
rect 317 35865 351 35899
rect 385 35865 419 35899
rect 453 35865 487 35899
rect 521 35865 555 35899
rect 589 35865 623 35899
rect 657 35865 691 35899
rect 725 35865 759 35899
rect 793 35865 827 35899
rect 861 35865 895 35899
rect 929 35865 963 35899
rect 997 35865 1031 35899
rect 1065 35865 1099 35899
rect 1133 35865 1167 35899
rect 1201 35865 1235 35899
rect 1269 35865 1303 35899
rect 2470 36225 2504 36259
rect 2538 36225 2572 36259
rect 2606 36225 2640 36259
rect 2674 36225 2708 36259
rect 2742 36225 2776 36259
rect 2810 36225 2844 36259
rect 2878 36225 2912 36259
rect 2946 36225 2980 36259
rect 3014 36225 3048 36259
rect 3082 36225 3116 36259
rect 3150 36225 3184 36259
rect 3218 36225 3252 36259
rect 3286 36225 3320 36259
rect 3354 36225 3388 36259
rect 3422 36225 3456 36259
rect 2352 36115 2386 36149
rect 3991 36225 4025 36259
rect 4059 36225 4093 36259
rect 4127 36225 4161 36259
rect 4195 36225 4229 36259
rect 4263 36225 4297 36259
rect 4331 36225 4365 36259
rect 4399 36225 4433 36259
rect 4467 36225 4501 36259
rect 4535 36225 4569 36259
rect 4603 36225 4637 36259
rect 4671 36225 4705 36259
rect 4739 36225 4773 36259
rect 4807 36225 4841 36259
rect 4875 36225 4909 36259
rect 4943 36225 4977 36259
rect 2352 36047 2386 36081
rect 3540 36115 3574 36149
rect 3540 36047 3574 36081
rect 3873 36115 3907 36149
rect 2352 35979 2386 36013
rect 3873 36047 3907 36081
rect 3540 35979 3574 36013
rect 2470 35869 2504 35903
rect 2538 35869 2572 35903
rect 2606 35869 2640 35903
rect 2674 35869 2708 35903
rect 2742 35869 2776 35903
rect 2810 35869 2844 35903
rect 2878 35869 2912 35903
rect 2946 35869 2980 35903
rect 3014 35869 3048 35903
rect 3082 35869 3116 35903
rect 3150 35869 3184 35903
rect 3218 35869 3252 35903
rect 3286 35869 3320 35903
rect 3354 35869 3388 35903
rect 3422 35869 3456 35903
rect 5061 36115 5095 36149
rect 5061 36047 5095 36081
rect 3873 35979 3907 36013
rect 5061 35979 5095 36013
rect 3991 35869 4025 35903
rect 4059 35869 4093 35903
rect 4127 35869 4161 35903
rect 4195 35869 4229 35903
rect 4263 35869 4297 35903
rect 4331 35869 4365 35903
rect 4399 35869 4433 35903
rect 4467 35869 4501 35903
rect 4535 35869 4569 35903
rect 4603 35869 4637 35903
rect 4671 35869 4705 35903
rect 4739 35869 4773 35903
rect 4807 35869 4841 35903
rect 4875 35869 4909 35903
rect 4943 35869 4977 35903
rect 317 34934 351 34968
rect 385 34934 419 34968
rect 453 34934 487 34968
rect 521 34934 555 34968
rect 589 34934 623 34968
rect 657 34934 691 34968
rect 725 34934 759 34968
rect 793 34934 827 34968
rect 861 34934 895 34968
rect 929 34934 963 34968
rect 997 34934 1031 34968
rect 1065 34934 1099 34968
rect 1133 34934 1167 34968
rect 1201 34934 1235 34968
rect 1269 34934 1303 34968
rect 199 34824 233 34858
rect 199 34756 233 34790
rect 1387 34824 1421 34858
rect 1387 34756 1421 34790
rect 199 34688 233 34722
rect 1387 34688 1421 34722
rect 317 34578 351 34612
rect 385 34578 419 34612
rect 453 34578 487 34612
rect 521 34578 555 34612
rect 589 34578 623 34612
rect 657 34578 691 34612
rect 725 34578 759 34612
rect 793 34578 827 34612
rect 861 34578 895 34612
rect 929 34578 963 34612
rect 997 34578 1031 34612
rect 1065 34578 1099 34612
rect 1133 34578 1167 34612
rect 1201 34578 1235 34612
rect 1269 34578 1303 34612
rect 2470 34938 2504 34972
rect 2538 34938 2572 34972
rect 2606 34938 2640 34972
rect 2674 34938 2708 34972
rect 2742 34938 2776 34972
rect 2810 34938 2844 34972
rect 2878 34938 2912 34972
rect 2946 34938 2980 34972
rect 3014 34938 3048 34972
rect 3082 34938 3116 34972
rect 3150 34938 3184 34972
rect 3218 34938 3252 34972
rect 3286 34938 3320 34972
rect 3354 34938 3388 34972
rect 3422 34938 3456 34972
rect 2352 34828 2386 34862
rect 3991 34938 4025 34972
rect 4059 34938 4093 34972
rect 4127 34938 4161 34972
rect 4195 34938 4229 34972
rect 4263 34938 4297 34972
rect 4331 34938 4365 34972
rect 4399 34938 4433 34972
rect 4467 34938 4501 34972
rect 4535 34938 4569 34972
rect 4603 34938 4637 34972
rect 4671 34938 4705 34972
rect 4739 34938 4773 34972
rect 4807 34938 4841 34972
rect 4875 34938 4909 34972
rect 4943 34938 4977 34972
rect 2352 34760 2386 34794
rect 3540 34828 3574 34862
rect 3540 34760 3574 34794
rect 3873 34828 3907 34862
rect 2352 34692 2386 34726
rect 3873 34760 3907 34794
rect 3540 34692 3574 34726
rect 2470 34582 2504 34616
rect 2538 34582 2572 34616
rect 2606 34582 2640 34616
rect 2674 34582 2708 34616
rect 2742 34582 2776 34616
rect 2810 34582 2844 34616
rect 2878 34582 2912 34616
rect 2946 34582 2980 34616
rect 3014 34582 3048 34616
rect 3082 34582 3116 34616
rect 3150 34582 3184 34616
rect 3218 34582 3252 34616
rect 3286 34582 3320 34616
rect 3354 34582 3388 34616
rect 3422 34582 3456 34616
rect 5061 34828 5095 34862
rect 5061 34760 5095 34794
rect 3873 34692 3907 34726
rect 5061 34692 5095 34726
rect 3991 34582 4025 34616
rect 4059 34582 4093 34616
rect 4127 34582 4161 34616
rect 4195 34582 4229 34616
rect 4263 34582 4297 34616
rect 4331 34582 4365 34616
rect 4399 34582 4433 34616
rect 4467 34582 4501 34616
rect 4535 34582 4569 34616
rect 4603 34582 4637 34616
rect 4671 34582 4705 34616
rect 4739 34582 4773 34616
rect 4807 34582 4841 34616
rect 4875 34582 4909 34616
rect 4943 34582 4977 34616
rect 317 33647 351 33681
rect 385 33647 419 33681
rect 453 33647 487 33681
rect 521 33647 555 33681
rect 589 33647 623 33681
rect 657 33647 691 33681
rect 725 33647 759 33681
rect 793 33647 827 33681
rect 861 33647 895 33681
rect 929 33647 963 33681
rect 997 33647 1031 33681
rect 1065 33647 1099 33681
rect 1133 33647 1167 33681
rect 1201 33647 1235 33681
rect 1269 33647 1303 33681
rect 199 33537 233 33571
rect 199 33469 233 33503
rect 1387 33537 1421 33571
rect 1387 33469 1421 33503
rect 199 33401 233 33435
rect 1387 33401 1421 33435
rect 317 33291 351 33325
rect 385 33291 419 33325
rect 453 33291 487 33325
rect 521 33291 555 33325
rect 589 33291 623 33325
rect 657 33291 691 33325
rect 725 33291 759 33325
rect 793 33291 827 33325
rect 861 33291 895 33325
rect 929 33291 963 33325
rect 997 33291 1031 33325
rect 1065 33291 1099 33325
rect 1133 33291 1167 33325
rect 1201 33291 1235 33325
rect 1269 33291 1303 33325
rect 2470 33651 2504 33685
rect 2538 33651 2572 33685
rect 2606 33651 2640 33685
rect 2674 33651 2708 33685
rect 2742 33651 2776 33685
rect 2810 33651 2844 33685
rect 2878 33651 2912 33685
rect 2946 33651 2980 33685
rect 3014 33651 3048 33685
rect 3082 33651 3116 33685
rect 3150 33651 3184 33685
rect 3218 33651 3252 33685
rect 3286 33651 3320 33685
rect 3354 33651 3388 33685
rect 3422 33651 3456 33685
rect 2352 33541 2386 33575
rect 3991 33651 4025 33685
rect 4059 33651 4093 33685
rect 4127 33651 4161 33685
rect 4195 33651 4229 33685
rect 4263 33651 4297 33685
rect 4331 33651 4365 33685
rect 4399 33651 4433 33685
rect 4467 33651 4501 33685
rect 4535 33651 4569 33685
rect 4603 33651 4637 33685
rect 4671 33651 4705 33685
rect 4739 33651 4773 33685
rect 4807 33651 4841 33685
rect 4875 33651 4909 33685
rect 4943 33651 4977 33685
rect 2352 33473 2386 33507
rect 3540 33541 3574 33575
rect 3540 33473 3574 33507
rect 3873 33541 3907 33575
rect 2352 33405 2386 33439
rect 3873 33473 3907 33507
rect 3540 33405 3574 33439
rect 2470 33295 2504 33329
rect 2538 33295 2572 33329
rect 2606 33295 2640 33329
rect 2674 33295 2708 33329
rect 2742 33295 2776 33329
rect 2810 33295 2844 33329
rect 2878 33295 2912 33329
rect 2946 33295 2980 33329
rect 3014 33295 3048 33329
rect 3082 33295 3116 33329
rect 3150 33295 3184 33329
rect 3218 33295 3252 33329
rect 3286 33295 3320 33329
rect 3354 33295 3388 33329
rect 3422 33295 3456 33329
rect 5061 33541 5095 33575
rect 5061 33473 5095 33507
rect 3873 33405 3907 33439
rect 5061 33405 5095 33439
rect 3991 33295 4025 33329
rect 4059 33295 4093 33329
rect 4127 33295 4161 33329
rect 4195 33295 4229 33329
rect 4263 33295 4297 33329
rect 4331 33295 4365 33329
rect 4399 33295 4433 33329
rect 4467 33295 4501 33329
rect 4535 33295 4569 33329
rect 4603 33295 4637 33329
rect 4671 33295 4705 33329
rect 4739 33295 4773 33329
rect 4807 33295 4841 33329
rect 4875 33295 4909 33329
rect 4943 33295 4977 33329
rect 317 32360 351 32394
rect 385 32360 419 32394
rect 453 32360 487 32394
rect 521 32360 555 32394
rect 589 32360 623 32394
rect 657 32360 691 32394
rect 725 32360 759 32394
rect 793 32360 827 32394
rect 861 32360 895 32394
rect 929 32360 963 32394
rect 997 32360 1031 32394
rect 1065 32360 1099 32394
rect 1133 32360 1167 32394
rect 1201 32360 1235 32394
rect 1269 32360 1303 32394
rect 199 32250 233 32284
rect 199 32182 233 32216
rect 1387 32250 1421 32284
rect 1387 32182 1421 32216
rect 199 32114 233 32148
rect 1387 32114 1421 32148
rect 317 32004 351 32038
rect 385 32004 419 32038
rect 453 32004 487 32038
rect 521 32004 555 32038
rect 589 32004 623 32038
rect 657 32004 691 32038
rect 725 32004 759 32038
rect 793 32004 827 32038
rect 861 32004 895 32038
rect 929 32004 963 32038
rect 997 32004 1031 32038
rect 1065 32004 1099 32038
rect 1133 32004 1167 32038
rect 1201 32004 1235 32038
rect 1269 32004 1303 32038
rect 2470 32364 2504 32398
rect 2538 32364 2572 32398
rect 2606 32364 2640 32398
rect 2674 32364 2708 32398
rect 2742 32364 2776 32398
rect 2810 32364 2844 32398
rect 2878 32364 2912 32398
rect 2946 32364 2980 32398
rect 3014 32364 3048 32398
rect 3082 32364 3116 32398
rect 3150 32364 3184 32398
rect 3218 32364 3252 32398
rect 3286 32364 3320 32398
rect 3354 32364 3388 32398
rect 3422 32364 3456 32398
rect 2352 32254 2386 32288
rect 3991 32364 4025 32398
rect 4059 32364 4093 32398
rect 4127 32364 4161 32398
rect 4195 32364 4229 32398
rect 4263 32364 4297 32398
rect 4331 32364 4365 32398
rect 4399 32364 4433 32398
rect 4467 32364 4501 32398
rect 4535 32364 4569 32398
rect 4603 32364 4637 32398
rect 4671 32364 4705 32398
rect 4739 32364 4773 32398
rect 4807 32364 4841 32398
rect 4875 32364 4909 32398
rect 4943 32364 4977 32398
rect 2352 32186 2386 32220
rect 3540 32254 3574 32288
rect 3540 32186 3574 32220
rect 3873 32254 3907 32288
rect 2352 32118 2386 32152
rect 3873 32186 3907 32220
rect 3540 32118 3574 32152
rect 2470 32008 2504 32042
rect 2538 32008 2572 32042
rect 2606 32008 2640 32042
rect 2674 32008 2708 32042
rect 2742 32008 2776 32042
rect 2810 32008 2844 32042
rect 2878 32008 2912 32042
rect 2946 32008 2980 32042
rect 3014 32008 3048 32042
rect 3082 32008 3116 32042
rect 3150 32008 3184 32042
rect 3218 32008 3252 32042
rect 3286 32008 3320 32042
rect 3354 32008 3388 32042
rect 3422 32008 3456 32042
rect 5061 32254 5095 32288
rect 5061 32186 5095 32220
rect 3873 32118 3907 32152
rect 5061 32118 5095 32152
rect 3991 32008 4025 32042
rect 4059 32008 4093 32042
rect 4127 32008 4161 32042
rect 4195 32008 4229 32042
rect 4263 32008 4297 32042
rect 4331 32008 4365 32042
rect 4399 32008 4433 32042
rect 4467 32008 4501 32042
rect 4535 32008 4569 32042
rect 4603 32008 4637 32042
rect 4671 32008 4705 32042
rect 4739 32008 4773 32042
rect 4807 32008 4841 32042
rect 4875 32008 4909 32042
rect 4943 32008 4977 32042
rect 317 31073 351 31107
rect 385 31073 419 31107
rect 453 31073 487 31107
rect 521 31073 555 31107
rect 589 31073 623 31107
rect 657 31073 691 31107
rect 725 31073 759 31107
rect 793 31073 827 31107
rect 861 31073 895 31107
rect 929 31073 963 31107
rect 997 31073 1031 31107
rect 1065 31073 1099 31107
rect 1133 31073 1167 31107
rect 1201 31073 1235 31107
rect 1269 31073 1303 31107
rect 199 30963 233 30997
rect 199 30895 233 30929
rect 1387 30963 1421 30997
rect 1387 30895 1421 30929
rect 199 30827 233 30861
rect 1387 30827 1421 30861
rect 317 30717 351 30751
rect 385 30717 419 30751
rect 453 30717 487 30751
rect 521 30717 555 30751
rect 589 30717 623 30751
rect 657 30717 691 30751
rect 725 30717 759 30751
rect 793 30717 827 30751
rect 861 30717 895 30751
rect 929 30717 963 30751
rect 997 30717 1031 30751
rect 1065 30717 1099 30751
rect 1133 30717 1167 30751
rect 1201 30717 1235 30751
rect 1269 30717 1303 30751
rect 2470 31077 2504 31111
rect 2538 31077 2572 31111
rect 2606 31077 2640 31111
rect 2674 31077 2708 31111
rect 2742 31077 2776 31111
rect 2810 31077 2844 31111
rect 2878 31077 2912 31111
rect 2946 31077 2980 31111
rect 3014 31077 3048 31111
rect 3082 31077 3116 31111
rect 3150 31077 3184 31111
rect 3218 31077 3252 31111
rect 3286 31077 3320 31111
rect 3354 31077 3388 31111
rect 3422 31077 3456 31111
rect 2352 30967 2386 31001
rect 3991 31077 4025 31111
rect 4059 31077 4093 31111
rect 4127 31077 4161 31111
rect 4195 31077 4229 31111
rect 4263 31077 4297 31111
rect 4331 31077 4365 31111
rect 4399 31077 4433 31111
rect 4467 31077 4501 31111
rect 4535 31077 4569 31111
rect 4603 31077 4637 31111
rect 4671 31077 4705 31111
rect 4739 31077 4773 31111
rect 4807 31077 4841 31111
rect 4875 31077 4909 31111
rect 4943 31077 4977 31111
rect 2352 30899 2386 30933
rect 3540 30967 3574 31001
rect 3540 30899 3574 30933
rect 3873 30967 3907 31001
rect 2352 30831 2386 30865
rect 3873 30899 3907 30933
rect 3540 30831 3574 30865
rect 2470 30721 2504 30755
rect 2538 30721 2572 30755
rect 2606 30721 2640 30755
rect 2674 30721 2708 30755
rect 2742 30721 2776 30755
rect 2810 30721 2844 30755
rect 2878 30721 2912 30755
rect 2946 30721 2980 30755
rect 3014 30721 3048 30755
rect 3082 30721 3116 30755
rect 3150 30721 3184 30755
rect 3218 30721 3252 30755
rect 3286 30721 3320 30755
rect 3354 30721 3388 30755
rect 3422 30721 3456 30755
rect 5061 30967 5095 31001
rect 5061 30899 5095 30933
rect 3873 30831 3907 30865
rect 5061 30831 5095 30865
rect 3991 30721 4025 30755
rect 4059 30721 4093 30755
rect 4127 30721 4161 30755
rect 4195 30721 4229 30755
rect 4263 30721 4297 30755
rect 4331 30721 4365 30755
rect 4399 30721 4433 30755
rect 4467 30721 4501 30755
rect 4535 30721 4569 30755
rect 4603 30721 4637 30755
rect 4671 30721 4705 30755
rect 4739 30721 4773 30755
rect 4807 30721 4841 30755
rect 4875 30721 4909 30755
rect 4943 30721 4977 30755
rect 317 29786 351 29820
rect 385 29786 419 29820
rect 453 29786 487 29820
rect 521 29786 555 29820
rect 589 29786 623 29820
rect 657 29786 691 29820
rect 725 29786 759 29820
rect 793 29786 827 29820
rect 861 29786 895 29820
rect 929 29786 963 29820
rect 997 29786 1031 29820
rect 1065 29786 1099 29820
rect 1133 29786 1167 29820
rect 1201 29786 1235 29820
rect 1269 29786 1303 29820
rect 199 29676 233 29710
rect 199 29608 233 29642
rect 1387 29676 1421 29710
rect 1387 29608 1421 29642
rect 199 29540 233 29574
rect 1387 29540 1421 29574
rect 317 29430 351 29464
rect 385 29430 419 29464
rect 453 29430 487 29464
rect 521 29430 555 29464
rect 589 29430 623 29464
rect 657 29430 691 29464
rect 725 29430 759 29464
rect 793 29430 827 29464
rect 861 29430 895 29464
rect 929 29430 963 29464
rect 997 29430 1031 29464
rect 1065 29430 1099 29464
rect 1133 29430 1167 29464
rect 1201 29430 1235 29464
rect 1269 29430 1303 29464
rect 2470 29790 2504 29824
rect 2538 29790 2572 29824
rect 2606 29790 2640 29824
rect 2674 29790 2708 29824
rect 2742 29790 2776 29824
rect 2810 29790 2844 29824
rect 2878 29790 2912 29824
rect 2946 29790 2980 29824
rect 3014 29790 3048 29824
rect 3082 29790 3116 29824
rect 3150 29790 3184 29824
rect 3218 29790 3252 29824
rect 3286 29790 3320 29824
rect 3354 29790 3388 29824
rect 3422 29790 3456 29824
rect 2352 29680 2386 29714
rect 3991 29790 4025 29824
rect 4059 29790 4093 29824
rect 4127 29790 4161 29824
rect 4195 29790 4229 29824
rect 4263 29790 4297 29824
rect 4331 29790 4365 29824
rect 4399 29790 4433 29824
rect 4467 29790 4501 29824
rect 4535 29790 4569 29824
rect 4603 29790 4637 29824
rect 4671 29790 4705 29824
rect 4739 29790 4773 29824
rect 4807 29790 4841 29824
rect 4875 29790 4909 29824
rect 4943 29790 4977 29824
rect 2352 29612 2386 29646
rect 3540 29680 3574 29714
rect 3540 29612 3574 29646
rect 3873 29680 3907 29714
rect 2352 29544 2386 29578
rect 3873 29612 3907 29646
rect 3540 29544 3574 29578
rect 2470 29434 2504 29468
rect 2538 29434 2572 29468
rect 2606 29434 2640 29468
rect 2674 29434 2708 29468
rect 2742 29434 2776 29468
rect 2810 29434 2844 29468
rect 2878 29434 2912 29468
rect 2946 29434 2980 29468
rect 3014 29434 3048 29468
rect 3082 29434 3116 29468
rect 3150 29434 3184 29468
rect 3218 29434 3252 29468
rect 3286 29434 3320 29468
rect 3354 29434 3388 29468
rect 3422 29434 3456 29468
rect 5061 29680 5095 29714
rect 5061 29612 5095 29646
rect 3873 29544 3907 29578
rect 5061 29544 5095 29578
rect 3991 29434 4025 29468
rect 4059 29434 4093 29468
rect 4127 29434 4161 29468
rect 4195 29434 4229 29468
rect 4263 29434 4297 29468
rect 4331 29434 4365 29468
rect 4399 29434 4433 29468
rect 4467 29434 4501 29468
rect 4535 29434 4569 29468
rect 4603 29434 4637 29468
rect 4671 29434 4705 29468
rect 4739 29434 4773 29468
rect 4807 29434 4841 29468
rect 4875 29434 4909 29468
rect 4943 29434 4977 29468
rect 317 28499 351 28533
rect 385 28499 419 28533
rect 453 28499 487 28533
rect 521 28499 555 28533
rect 589 28499 623 28533
rect 657 28499 691 28533
rect 725 28499 759 28533
rect 793 28499 827 28533
rect 861 28499 895 28533
rect 929 28499 963 28533
rect 997 28499 1031 28533
rect 1065 28499 1099 28533
rect 1133 28499 1167 28533
rect 1201 28499 1235 28533
rect 1269 28499 1303 28533
rect 199 28389 233 28423
rect 199 28321 233 28355
rect 1387 28389 1421 28423
rect 1387 28321 1421 28355
rect 199 28253 233 28287
rect 1387 28253 1421 28287
rect 317 28143 351 28177
rect 385 28143 419 28177
rect 453 28143 487 28177
rect 521 28143 555 28177
rect 589 28143 623 28177
rect 657 28143 691 28177
rect 725 28143 759 28177
rect 793 28143 827 28177
rect 861 28143 895 28177
rect 929 28143 963 28177
rect 997 28143 1031 28177
rect 1065 28143 1099 28177
rect 1133 28143 1167 28177
rect 1201 28143 1235 28177
rect 1269 28143 1303 28177
rect 2470 28503 2504 28537
rect 2538 28503 2572 28537
rect 2606 28503 2640 28537
rect 2674 28503 2708 28537
rect 2742 28503 2776 28537
rect 2810 28503 2844 28537
rect 2878 28503 2912 28537
rect 2946 28503 2980 28537
rect 3014 28503 3048 28537
rect 3082 28503 3116 28537
rect 3150 28503 3184 28537
rect 3218 28503 3252 28537
rect 3286 28503 3320 28537
rect 3354 28503 3388 28537
rect 3422 28503 3456 28537
rect 2352 28393 2386 28427
rect 3991 28503 4025 28537
rect 4059 28503 4093 28537
rect 4127 28503 4161 28537
rect 4195 28503 4229 28537
rect 4263 28503 4297 28537
rect 4331 28503 4365 28537
rect 4399 28503 4433 28537
rect 4467 28503 4501 28537
rect 4535 28503 4569 28537
rect 4603 28503 4637 28537
rect 4671 28503 4705 28537
rect 4739 28503 4773 28537
rect 4807 28503 4841 28537
rect 4875 28503 4909 28537
rect 4943 28503 4977 28537
rect 2352 28325 2386 28359
rect 3540 28393 3574 28427
rect 3540 28325 3574 28359
rect 3873 28393 3907 28427
rect 2352 28257 2386 28291
rect 3873 28325 3907 28359
rect 3540 28257 3574 28291
rect 2470 28147 2504 28181
rect 2538 28147 2572 28181
rect 2606 28147 2640 28181
rect 2674 28147 2708 28181
rect 2742 28147 2776 28181
rect 2810 28147 2844 28181
rect 2878 28147 2912 28181
rect 2946 28147 2980 28181
rect 3014 28147 3048 28181
rect 3082 28147 3116 28181
rect 3150 28147 3184 28181
rect 3218 28147 3252 28181
rect 3286 28147 3320 28181
rect 3354 28147 3388 28181
rect 3422 28147 3456 28181
rect 5061 28393 5095 28427
rect 5061 28325 5095 28359
rect 3873 28257 3907 28291
rect 5061 28257 5095 28291
rect 3991 28147 4025 28181
rect 4059 28147 4093 28181
rect 4127 28147 4161 28181
rect 4195 28147 4229 28181
rect 4263 28147 4297 28181
rect 4331 28147 4365 28181
rect 4399 28147 4433 28181
rect 4467 28147 4501 28181
rect 4535 28147 4569 28181
rect 4603 28147 4637 28181
rect 4671 28147 4705 28181
rect 4739 28147 4773 28181
rect 4807 28147 4841 28181
rect 4875 28147 4909 28181
rect 4943 28147 4977 28181
rect 317 27212 351 27246
rect 385 27212 419 27246
rect 453 27212 487 27246
rect 521 27212 555 27246
rect 589 27212 623 27246
rect 657 27212 691 27246
rect 725 27212 759 27246
rect 793 27212 827 27246
rect 861 27212 895 27246
rect 929 27212 963 27246
rect 997 27212 1031 27246
rect 1065 27212 1099 27246
rect 1133 27212 1167 27246
rect 1201 27212 1235 27246
rect 1269 27212 1303 27246
rect 199 27102 233 27136
rect 199 27034 233 27068
rect 1387 27102 1421 27136
rect 1387 27034 1421 27068
rect 199 26966 233 27000
rect 1387 26966 1421 27000
rect 317 26856 351 26890
rect 385 26856 419 26890
rect 453 26856 487 26890
rect 521 26856 555 26890
rect 589 26856 623 26890
rect 657 26856 691 26890
rect 725 26856 759 26890
rect 793 26856 827 26890
rect 861 26856 895 26890
rect 929 26856 963 26890
rect 997 26856 1031 26890
rect 1065 26856 1099 26890
rect 1133 26856 1167 26890
rect 1201 26856 1235 26890
rect 1269 26856 1303 26890
rect 2470 27216 2504 27250
rect 2538 27216 2572 27250
rect 2606 27216 2640 27250
rect 2674 27216 2708 27250
rect 2742 27216 2776 27250
rect 2810 27216 2844 27250
rect 2878 27216 2912 27250
rect 2946 27216 2980 27250
rect 3014 27216 3048 27250
rect 3082 27216 3116 27250
rect 3150 27216 3184 27250
rect 3218 27216 3252 27250
rect 3286 27216 3320 27250
rect 3354 27216 3388 27250
rect 3422 27216 3456 27250
rect 2352 27106 2386 27140
rect 3991 27216 4025 27250
rect 4059 27216 4093 27250
rect 4127 27216 4161 27250
rect 4195 27216 4229 27250
rect 4263 27216 4297 27250
rect 4331 27216 4365 27250
rect 4399 27216 4433 27250
rect 4467 27216 4501 27250
rect 4535 27216 4569 27250
rect 4603 27216 4637 27250
rect 4671 27216 4705 27250
rect 4739 27216 4773 27250
rect 4807 27216 4841 27250
rect 4875 27216 4909 27250
rect 4943 27216 4977 27250
rect 2352 27038 2386 27072
rect 3540 27106 3574 27140
rect 3540 27038 3574 27072
rect 3873 27106 3907 27140
rect 2352 26970 2386 27004
rect 3873 27038 3907 27072
rect 3540 26970 3574 27004
rect 2470 26860 2504 26894
rect 2538 26860 2572 26894
rect 2606 26860 2640 26894
rect 2674 26860 2708 26894
rect 2742 26860 2776 26894
rect 2810 26860 2844 26894
rect 2878 26860 2912 26894
rect 2946 26860 2980 26894
rect 3014 26860 3048 26894
rect 3082 26860 3116 26894
rect 3150 26860 3184 26894
rect 3218 26860 3252 26894
rect 3286 26860 3320 26894
rect 3354 26860 3388 26894
rect 3422 26860 3456 26894
rect 5061 27106 5095 27140
rect 5061 27038 5095 27072
rect 3873 26970 3907 27004
rect 5061 26970 5095 27004
rect 3991 26860 4025 26894
rect 4059 26860 4093 26894
rect 4127 26860 4161 26894
rect 4195 26860 4229 26894
rect 4263 26860 4297 26894
rect 4331 26860 4365 26894
rect 4399 26860 4433 26894
rect 4467 26860 4501 26894
rect 4535 26860 4569 26894
rect 4603 26860 4637 26894
rect 4671 26860 4705 26894
rect 4739 26860 4773 26894
rect 4807 26860 4841 26894
rect 4875 26860 4909 26894
rect 4943 26860 4977 26894
rect 317 25925 351 25959
rect 385 25925 419 25959
rect 453 25925 487 25959
rect 521 25925 555 25959
rect 589 25925 623 25959
rect 657 25925 691 25959
rect 725 25925 759 25959
rect 793 25925 827 25959
rect 861 25925 895 25959
rect 929 25925 963 25959
rect 997 25925 1031 25959
rect 1065 25925 1099 25959
rect 1133 25925 1167 25959
rect 1201 25925 1235 25959
rect 1269 25925 1303 25959
rect 199 25815 233 25849
rect 199 25747 233 25781
rect 1387 25815 1421 25849
rect 1387 25747 1421 25781
rect 199 25679 233 25713
rect 1387 25679 1421 25713
rect 317 25569 351 25603
rect 385 25569 419 25603
rect 453 25569 487 25603
rect 521 25569 555 25603
rect 589 25569 623 25603
rect 657 25569 691 25603
rect 725 25569 759 25603
rect 793 25569 827 25603
rect 861 25569 895 25603
rect 929 25569 963 25603
rect 997 25569 1031 25603
rect 1065 25569 1099 25603
rect 1133 25569 1167 25603
rect 1201 25569 1235 25603
rect 1269 25569 1303 25603
rect 2470 25929 2504 25963
rect 2538 25929 2572 25963
rect 2606 25929 2640 25963
rect 2674 25929 2708 25963
rect 2742 25929 2776 25963
rect 2810 25929 2844 25963
rect 2878 25929 2912 25963
rect 2946 25929 2980 25963
rect 3014 25929 3048 25963
rect 3082 25929 3116 25963
rect 3150 25929 3184 25963
rect 3218 25929 3252 25963
rect 3286 25929 3320 25963
rect 3354 25929 3388 25963
rect 3422 25929 3456 25963
rect 2352 25819 2386 25853
rect 3991 25929 4025 25963
rect 4059 25929 4093 25963
rect 4127 25929 4161 25963
rect 4195 25929 4229 25963
rect 4263 25929 4297 25963
rect 4331 25929 4365 25963
rect 4399 25929 4433 25963
rect 4467 25929 4501 25963
rect 4535 25929 4569 25963
rect 4603 25929 4637 25963
rect 4671 25929 4705 25963
rect 4739 25929 4773 25963
rect 4807 25929 4841 25963
rect 4875 25929 4909 25963
rect 4943 25929 4977 25963
rect 2352 25751 2386 25785
rect 3540 25819 3574 25853
rect 3540 25751 3574 25785
rect 3873 25819 3907 25853
rect 2352 25683 2386 25717
rect 3873 25751 3907 25785
rect 3540 25683 3574 25717
rect 2470 25573 2504 25607
rect 2538 25573 2572 25607
rect 2606 25573 2640 25607
rect 2674 25573 2708 25607
rect 2742 25573 2776 25607
rect 2810 25573 2844 25607
rect 2878 25573 2912 25607
rect 2946 25573 2980 25607
rect 3014 25573 3048 25607
rect 3082 25573 3116 25607
rect 3150 25573 3184 25607
rect 3218 25573 3252 25607
rect 3286 25573 3320 25607
rect 3354 25573 3388 25607
rect 3422 25573 3456 25607
rect 5061 25819 5095 25853
rect 5061 25751 5095 25785
rect 3873 25683 3907 25717
rect 5061 25683 5095 25717
rect 3991 25573 4025 25607
rect 4059 25573 4093 25607
rect 4127 25573 4161 25607
rect 4195 25573 4229 25607
rect 4263 25573 4297 25607
rect 4331 25573 4365 25607
rect 4399 25573 4433 25607
rect 4467 25573 4501 25607
rect 4535 25573 4569 25607
rect 4603 25573 4637 25607
rect 4671 25573 4705 25607
rect 4739 25573 4773 25607
rect 4807 25573 4841 25607
rect 4875 25573 4909 25607
rect 4943 25573 4977 25607
rect 317 24638 351 24672
rect 385 24638 419 24672
rect 453 24638 487 24672
rect 521 24638 555 24672
rect 589 24638 623 24672
rect 657 24638 691 24672
rect 725 24638 759 24672
rect 793 24638 827 24672
rect 861 24638 895 24672
rect 929 24638 963 24672
rect 997 24638 1031 24672
rect 1065 24638 1099 24672
rect 1133 24638 1167 24672
rect 1201 24638 1235 24672
rect 1269 24638 1303 24672
rect 199 24528 233 24562
rect 199 24460 233 24494
rect 1387 24528 1421 24562
rect 1387 24460 1421 24494
rect 199 24392 233 24426
rect 1387 24392 1421 24426
rect 317 24282 351 24316
rect 385 24282 419 24316
rect 453 24282 487 24316
rect 521 24282 555 24316
rect 589 24282 623 24316
rect 657 24282 691 24316
rect 725 24282 759 24316
rect 793 24282 827 24316
rect 861 24282 895 24316
rect 929 24282 963 24316
rect 997 24282 1031 24316
rect 1065 24282 1099 24316
rect 1133 24282 1167 24316
rect 1201 24282 1235 24316
rect 1269 24282 1303 24316
rect 2470 24642 2504 24676
rect 2538 24642 2572 24676
rect 2606 24642 2640 24676
rect 2674 24642 2708 24676
rect 2742 24642 2776 24676
rect 2810 24642 2844 24676
rect 2878 24642 2912 24676
rect 2946 24642 2980 24676
rect 3014 24642 3048 24676
rect 3082 24642 3116 24676
rect 3150 24642 3184 24676
rect 3218 24642 3252 24676
rect 3286 24642 3320 24676
rect 3354 24642 3388 24676
rect 3422 24642 3456 24676
rect 2352 24532 2386 24566
rect 3991 24642 4025 24676
rect 4059 24642 4093 24676
rect 4127 24642 4161 24676
rect 4195 24642 4229 24676
rect 4263 24642 4297 24676
rect 4331 24642 4365 24676
rect 4399 24642 4433 24676
rect 4467 24642 4501 24676
rect 4535 24642 4569 24676
rect 4603 24642 4637 24676
rect 4671 24642 4705 24676
rect 4739 24642 4773 24676
rect 4807 24642 4841 24676
rect 4875 24642 4909 24676
rect 4943 24642 4977 24676
rect 2352 24464 2386 24498
rect 3540 24532 3574 24566
rect 3540 24464 3574 24498
rect 3873 24532 3907 24566
rect 2352 24396 2386 24430
rect 3873 24464 3907 24498
rect 3540 24396 3574 24430
rect 2470 24286 2504 24320
rect 2538 24286 2572 24320
rect 2606 24286 2640 24320
rect 2674 24286 2708 24320
rect 2742 24286 2776 24320
rect 2810 24286 2844 24320
rect 2878 24286 2912 24320
rect 2946 24286 2980 24320
rect 3014 24286 3048 24320
rect 3082 24286 3116 24320
rect 3150 24286 3184 24320
rect 3218 24286 3252 24320
rect 3286 24286 3320 24320
rect 3354 24286 3388 24320
rect 3422 24286 3456 24320
rect 5061 24532 5095 24566
rect 5061 24464 5095 24498
rect 3873 24396 3907 24430
rect 5061 24396 5095 24430
rect 3991 24286 4025 24320
rect 4059 24286 4093 24320
rect 4127 24286 4161 24320
rect 4195 24286 4229 24320
rect 4263 24286 4297 24320
rect 4331 24286 4365 24320
rect 4399 24286 4433 24320
rect 4467 24286 4501 24320
rect 4535 24286 4569 24320
rect 4603 24286 4637 24320
rect 4671 24286 4705 24320
rect 4739 24286 4773 24320
rect 4807 24286 4841 24320
rect 4875 24286 4909 24320
rect 4943 24286 4977 24320
rect 317 23351 351 23385
rect 385 23351 419 23385
rect 453 23351 487 23385
rect 521 23351 555 23385
rect 589 23351 623 23385
rect 657 23351 691 23385
rect 725 23351 759 23385
rect 793 23351 827 23385
rect 861 23351 895 23385
rect 929 23351 963 23385
rect 997 23351 1031 23385
rect 1065 23351 1099 23385
rect 1133 23351 1167 23385
rect 1201 23351 1235 23385
rect 1269 23351 1303 23385
rect 199 23241 233 23275
rect 199 23173 233 23207
rect 1387 23241 1421 23275
rect 1387 23173 1421 23207
rect 199 23105 233 23139
rect 1387 23105 1421 23139
rect 317 22995 351 23029
rect 385 22995 419 23029
rect 453 22995 487 23029
rect 521 22995 555 23029
rect 589 22995 623 23029
rect 657 22995 691 23029
rect 725 22995 759 23029
rect 793 22995 827 23029
rect 861 22995 895 23029
rect 929 22995 963 23029
rect 997 22995 1031 23029
rect 1065 22995 1099 23029
rect 1133 22995 1167 23029
rect 1201 22995 1235 23029
rect 1269 22995 1303 23029
rect 2470 23355 2504 23389
rect 2538 23355 2572 23389
rect 2606 23355 2640 23389
rect 2674 23355 2708 23389
rect 2742 23355 2776 23389
rect 2810 23355 2844 23389
rect 2878 23355 2912 23389
rect 2946 23355 2980 23389
rect 3014 23355 3048 23389
rect 3082 23355 3116 23389
rect 3150 23355 3184 23389
rect 3218 23355 3252 23389
rect 3286 23355 3320 23389
rect 3354 23355 3388 23389
rect 3422 23355 3456 23389
rect 2352 23245 2386 23279
rect 3991 23355 4025 23389
rect 4059 23355 4093 23389
rect 4127 23355 4161 23389
rect 4195 23355 4229 23389
rect 4263 23355 4297 23389
rect 4331 23355 4365 23389
rect 4399 23355 4433 23389
rect 4467 23355 4501 23389
rect 4535 23355 4569 23389
rect 4603 23355 4637 23389
rect 4671 23355 4705 23389
rect 4739 23355 4773 23389
rect 4807 23355 4841 23389
rect 4875 23355 4909 23389
rect 4943 23355 4977 23389
rect 2352 23177 2386 23211
rect 3540 23245 3574 23279
rect 3540 23177 3574 23211
rect 3873 23245 3907 23279
rect 2352 23109 2386 23143
rect 3873 23177 3907 23211
rect 3540 23109 3574 23143
rect 2470 22999 2504 23033
rect 2538 22999 2572 23033
rect 2606 22999 2640 23033
rect 2674 22999 2708 23033
rect 2742 22999 2776 23033
rect 2810 22999 2844 23033
rect 2878 22999 2912 23033
rect 2946 22999 2980 23033
rect 3014 22999 3048 23033
rect 3082 22999 3116 23033
rect 3150 22999 3184 23033
rect 3218 22999 3252 23033
rect 3286 22999 3320 23033
rect 3354 22999 3388 23033
rect 3422 22999 3456 23033
rect 5061 23245 5095 23279
rect 5061 23177 5095 23211
rect 3873 23109 3907 23143
rect 5061 23109 5095 23143
rect 3991 22999 4025 23033
rect 4059 22999 4093 23033
rect 4127 22999 4161 23033
rect 4195 22999 4229 23033
rect 4263 22999 4297 23033
rect 4331 22999 4365 23033
rect 4399 22999 4433 23033
rect 4467 22999 4501 23033
rect 4535 22999 4569 23033
rect 4603 22999 4637 23033
rect 4671 22999 4705 23033
rect 4739 22999 4773 23033
rect 4807 22999 4841 23033
rect 4875 22999 4909 23033
rect 4943 22999 4977 23033
rect 317 22064 351 22098
rect 385 22064 419 22098
rect 453 22064 487 22098
rect 521 22064 555 22098
rect 589 22064 623 22098
rect 657 22064 691 22098
rect 725 22064 759 22098
rect 793 22064 827 22098
rect 861 22064 895 22098
rect 929 22064 963 22098
rect 997 22064 1031 22098
rect 1065 22064 1099 22098
rect 1133 22064 1167 22098
rect 1201 22064 1235 22098
rect 1269 22064 1303 22098
rect 199 21954 233 21988
rect 199 21886 233 21920
rect 1387 21954 1421 21988
rect 1387 21886 1421 21920
rect 199 21818 233 21852
rect 1387 21818 1421 21852
rect 317 21708 351 21742
rect 385 21708 419 21742
rect 453 21708 487 21742
rect 521 21708 555 21742
rect 589 21708 623 21742
rect 657 21708 691 21742
rect 725 21708 759 21742
rect 793 21708 827 21742
rect 861 21708 895 21742
rect 929 21708 963 21742
rect 997 21708 1031 21742
rect 1065 21708 1099 21742
rect 1133 21708 1167 21742
rect 1201 21708 1235 21742
rect 1269 21708 1303 21742
rect 2470 22068 2504 22102
rect 2538 22068 2572 22102
rect 2606 22068 2640 22102
rect 2674 22068 2708 22102
rect 2742 22068 2776 22102
rect 2810 22068 2844 22102
rect 2878 22068 2912 22102
rect 2946 22068 2980 22102
rect 3014 22068 3048 22102
rect 3082 22068 3116 22102
rect 3150 22068 3184 22102
rect 3218 22068 3252 22102
rect 3286 22068 3320 22102
rect 3354 22068 3388 22102
rect 3422 22068 3456 22102
rect 2352 21958 2386 21992
rect 3991 22068 4025 22102
rect 4059 22068 4093 22102
rect 4127 22068 4161 22102
rect 4195 22068 4229 22102
rect 4263 22068 4297 22102
rect 4331 22068 4365 22102
rect 4399 22068 4433 22102
rect 4467 22068 4501 22102
rect 4535 22068 4569 22102
rect 4603 22068 4637 22102
rect 4671 22068 4705 22102
rect 4739 22068 4773 22102
rect 4807 22068 4841 22102
rect 4875 22068 4909 22102
rect 4943 22068 4977 22102
rect 2352 21890 2386 21924
rect 3540 21958 3574 21992
rect 3540 21890 3574 21924
rect 3873 21958 3907 21992
rect 2352 21822 2386 21856
rect 3873 21890 3907 21924
rect 3540 21822 3574 21856
rect 2470 21712 2504 21746
rect 2538 21712 2572 21746
rect 2606 21712 2640 21746
rect 2674 21712 2708 21746
rect 2742 21712 2776 21746
rect 2810 21712 2844 21746
rect 2878 21712 2912 21746
rect 2946 21712 2980 21746
rect 3014 21712 3048 21746
rect 3082 21712 3116 21746
rect 3150 21712 3184 21746
rect 3218 21712 3252 21746
rect 3286 21712 3320 21746
rect 3354 21712 3388 21746
rect 3422 21712 3456 21746
rect 5061 21958 5095 21992
rect 5061 21890 5095 21924
rect 3873 21822 3907 21856
rect 5061 21822 5095 21856
rect 3991 21712 4025 21746
rect 4059 21712 4093 21746
rect 4127 21712 4161 21746
rect 4195 21712 4229 21746
rect 4263 21712 4297 21746
rect 4331 21712 4365 21746
rect 4399 21712 4433 21746
rect 4467 21712 4501 21746
rect 4535 21712 4569 21746
rect 4603 21712 4637 21746
rect 4671 21712 4705 21746
rect 4739 21712 4773 21746
rect 4807 21712 4841 21746
rect 4875 21712 4909 21746
rect 4943 21712 4977 21746
rect 317 20777 351 20811
rect 385 20777 419 20811
rect 453 20777 487 20811
rect 521 20777 555 20811
rect 589 20777 623 20811
rect 657 20777 691 20811
rect 725 20777 759 20811
rect 793 20777 827 20811
rect 861 20777 895 20811
rect 929 20777 963 20811
rect 997 20777 1031 20811
rect 1065 20777 1099 20811
rect 1133 20777 1167 20811
rect 1201 20777 1235 20811
rect 1269 20777 1303 20811
rect 199 20667 233 20701
rect 199 20599 233 20633
rect 1387 20667 1421 20701
rect 1387 20599 1421 20633
rect 199 20531 233 20565
rect 1387 20531 1421 20565
rect 317 20421 351 20455
rect 385 20421 419 20455
rect 453 20421 487 20455
rect 521 20421 555 20455
rect 589 20421 623 20455
rect 657 20421 691 20455
rect 725 20421 759 20455
rect 793 20421 827 20455
rect 861 20421 895 20455
rect 929 20421 963 20455
rect 997 20421 1031 20455
rect 1065 20421 1099 20455
rect 1133 20421 1167 20455
rect 1201 20421 1235 20455
rect 1269 20421 1303 20455
rect 2470 20781 2504 20815
rect 2538 20781 2572 20815
rect 2606 20781 2640 20815
rect 2674 20781 2708 20815
rect 2742 20781 2776 20815
rect 2810 20781 2844 20815
rect 2878 20781 2912 20815
rect 2946 20781 2980 20815
rect 3014 20781 3048 20815
rect 3082 20781 3116 20815
rect 3150 20781 3184 20815
rect 3218 20781 3252 20815
rect 3286 20781 3320 20815
rect 3354 20781 3388 20815
rect 3422 20781 3456 20815
rect 2352 20671 2386 20705
rect 3991 20781 4025 20815
rect 4059 20781 4093 20815
rect 4127 20781 4161 20815
rect 4195 20781 4229 20815
rect 4263 20781 4297 20815
rect 4331 20781 4365 20815
rect 4399 20781 4433 20815
rect 4467 20781 4501 20815
rect 4535 20781 4569 20815
rect 4603 20781 4637 20815
rect 4671 20781 4705 20815
rect 4739 20781 4773 20815
rect 4807 20781 4841 20815
rect 4875 20781 4909 20815
rect 4943 20781 4977 20815
rect 2352 20603 2386 20637
rect 3540 20671 3574 20705
rect 3540 20603 3574 20637
rect 3873 20671 3907 20705
rect 2352 20535 2386 20569
rect 3873 20603 3907 20637
rect 3540 20535 3574 20569
rect 2470 20425 2504 20459
rect 2538 20425 2572 20459
rect 2606 20425 2640 20459
rect 2674 20425 2708 20459
rect 2742 20425 2776 20459
rect 2810 20425 2844 20459
rect 2878 20425 2912 20459
rect 2946 20425 2980 20459
rect 3014 20425 3048 20459
rect 3082 20425 3116 20459
rect 3150 20425 3184 20459
rect 3218 20425 3252 20459
rect 3286 20425 3320 20459
rect 3354 20425 3388 20459
rect 3422 20425 3456 20459
rect 5061 20671 5095 20705
rect 5061 20603 5095 20637
rect 3873 20535 3907 20569
rect 5061 20535 5095 20569
rect 3991 20425 4025 20459
rect 4059 20425 4093 20459
rect 4127 20425 4161 20459
rect 4195 20425 4229 20459
rect 4263 20425 4297 20459
rect 4331 20425 4365 20459
rect 4399 20425 4433 20459
rect 4467 20425 4501 20459
rect 4535 20425 4569 20459
rect 4603 20425 4637 20459
rect 4671 20425 4705 20459
rect 4739 20425 4773 20459
rect 4807 20425 4841 20459
rect 4875 20425 4909 20459
rect 4943 20425 4977 20459
rect 317 19490 351 19524
rect 385 19490 419 19524
rect 453 19490 487 19524
rect 521 19490 555 19524
rect 589 19490 623 19524
rect 657 19490 691 19524
rect 725 19490 759 19524
rect 793 19490 827 19524
rect 861 19490 895 19524
rect 929 19490 963 19524
rect 997 19490 1031 19524
rect 1065 19490 1099 19524
rect 1133 19490 1167 19524
rect 1201 19490 1235 19524
rect 1269 19490 1303 19524
rect 199 19380 233 19414
rect 199 19312 233 19346
rect 1387 19380 1421 19414
rect 1387 19312 1421 19346
rect 199 19244 233 19278
rect 1387 19244 1421 19278
rect 317 19134 351 19168
rect 385 19134 419 19168
rect 453 19134 487 19168
rect 521 19134 555 19168
rect 589 19134 623 19168
rect 657 19134 691 19168
rect 725 19134 759 19168
rect 793 19134 827 19168
rect 861 19134 895 19168
rect 929 19134 963 19168
rect 997 19134 1031 19168
rect 1065 19134 1099 19168
rect 1133 19134 1167 19168
rect 1201 19134 1235 19168
rect 1269 19134 1303 19168
rect 2470 19494 2504 19528
rect 2538 19494 2572 19528
rect 2606 19494 2640 19528
rect 2674 19494 2708 19528
rect 2742 19494 2776 19528
rect 2810 19494 2844 19528
rect 2878 19494 2912 19528
rect 2946 19494 2980 19528
rect 3014 19494 3048 19528
rect 3082 19494 3116 19528
rect 3150 19494 3184 19528
rect 3218 19494 3252 19528
rect 3286 19494 3320 19528
rect 3354 19494 3388 19528
rect 3422 19494 3456 19528
rect 2352 19384 2386 19418
rect 3991 19494 4025 19528
rect 4059 19494 4093 19528
rect 4127 19494 4161 19528
rect 4195 19494 4229 19528
rect 4263 19494 4297 19528
rect 4331 19494 4365 19528
rect 4399 19494 4433 19528
rect 4467 19494 4501 19528
rect 4535 19494 4569 19528
rect 4603 19494 4637 19528
rect 4671 19494 4705 19528
rect 4739 19494 4773 19528
rect 4807 19494 4841 19528
rect 4875 19494 4909 19528
rect 4943 19494 4977 19528
rect 2352 19316 2386 19350
rect 3540 19384 3574 19418
rect 3540 19316 3574 19350
rect 3873 19384 3907 19418
rect 2352 19248 2386 19282
rect 3873 19316 3907 19350
rect 3540 19248 3574 19282
rect 2470 19138 2504 19172
rect 2538 19138 2572 19172
rect 2606 19138 2640 19172
rect 2674 19138 2708 19172
rect 2742 19138 2776 19172
rect 2810 19138 2844 19172
rect 2878 19138 2912 19172
rect 2946 19138 2980 19172
rect 3014 19138 3048 19172
rect 3082 19138 3116 19172
rect 3150 19138 3184 19172
rect 3218 19138 3252 19172
rect 3286 19138 3320 19172
rect 3354 19138 3388 19172
rect 3422 19138 3456 19172
rect 5061 19384 5095 19418
rect 5061 19316 5095 19350
rect 3873 19248 3907 19282
rect 5061 19248 5095 19282
rect 3991 19138 4025 19172
rect 4059 19138 4093 19172
rect 4127 19138 4161 19172
rect 4195 19138 4229 19172
rect 4263 19138 4297 19172
rect 4331 19138 4365 19172
rect 4399 19138 4433 19172
rect 4467 19138 4501 19172
rect 4535 19138 4569 19172
rect 4603 19138 4637 19172
rect 4671 19138 4705 19172
rect 4739 19138 4773 19172
rect 4807 19138 4841 19172
rect 4875 19138 4909 19172
rect 4943 19138 4977 19172
rect 317 18203 351 18237
rect 385 18203 419 18237
rect 453 18203 487 18237
rect 521 18203 555 18237
rect 589 18203 623 18237
rect 657 18203 691 18237
rect 725 18203 759 18237
rect 793 18203 827 18237
rect 861 18203 895 18237
rect 929 18203 963 18237
rect 997 18203 1031 18237
rect 1065 18203 1099 18237
rect 1133 18203 1167 18237
rect 1201 18203 1235 18237
rect 1269 18203 1303 18237
rect 199 18093 233 18127
rect 199 18025 233 18059
rect 1387 18093 1421 18127
rect 1387 18025 1421 18059
rect 199 17957 233 17991
rect 1387 17957 1421 17991
rect 317 17847 351 17881
rect 385 17847 419 17881
rect 453 17847 487 17881
rect 521 17847 555 17881
rect 589 17847 623 17881
rect 657 17847 691 17881
rect 725 17847 759 17881
rect 793 17847 827 17881
rect 861 17847 895 17881
rect 929 17847 963 17881
rect 997 17847 1031 17881
rect 1065 17847 1099 17881
rect 1133 17847 1167 17881
rect 1201 17847 1235 17881
rect 1269 17847 1303 17881
rect 2470 18207 2504 18241
rect 2538 18207 2572 18241
rect 2606 18207 2640 18241
rect 2674 18207 2708 18241
rect 2742 18207 2776 18241
rect 2810 18207 2844 18241
rect 2878 18207 2912 18241
rect 2946 18207 2980 18241
rect 3014 18207 3048 18241
rect 3082 18207 3116 18241
rect 3150 18207 3184 18241
rect 3218 18207 3252 18241
rect 3286 18207 3320 18241
rect 3354 18207 3388 18241
rect 3422 18207 3456 18241
rect 2352 18097 2386 18131
rect 3991 18207 4025 18241
rect 4059 18207 4093 18241
rect 4127 18207 4161 18241
rect 4195 18207 4229 18241
rect 4263 18207 4297 18241
rect 4331 18207 4365 18241
rect 4399 18207 4433 18241
rect 4467 18207 4501 18241
rect 4535 18207 4569 18241
rect 4603 18207 4637 18241
rect 4671 18207 4705 18241
rect 4739 18207 4773 18241
rect 4807 18207 4841 18241
rect 4875 18207 4909 18241
rect 4943 18207 4977 18241
rect 2352 18029 2386 18063
rect 3540 18097 3574 18131
rect 3540 18029 3574 18063
rect 3873 18097 3907 18131
rect 2352 17961 2386 17995
rect 3873 18029 3907 18063
rect 3540 17961 3574 17995
rect 2470 17851 2504 17885
rect 2538 17851 2572 17885
rect 2606 17851 2640 17885
rect 2674 17851 2708 17885
rect 2742 17851 2776 17885
rect 2810 17851 2844 17885
rect 2878 17851 2912 17885
rect 2946 17851 2980 17885
rect 3014 17851 3048 17885
rect 3082 17851 3116 17885
rect 3150 17851 3184 17885
rect 3218 17851 3252 17885
rect 3286 17851 3320 17885
rect 3354 17851 3388 17885
rect 3422 17851 3456 17885
rect 5061 18097 5095 18131
rect 5061 18029 5095 18063
rect 3873 17961 3907 17995
rect 5061 17961 5095 17995
rect 3991 17851 4025 17885
rect 4059 17851 4093 17885
rect 4127 17851 4161 17885
rect 4195 17851 4229 17885
rect 4263 17851 4297 17885
rect 4331 17851 4365 17885
rect 4399 17851 4433 17885
rect 4467 17851 4501 17885
rect 4535 17851 4569 17885
rect 4603 17851 4637 17885
rect 4671 17851 4705 17885
rect 4739 17851 4773 17885
rect 4807 17851 4841 17885
rect 4875 17851 4909 17885
rect 4943 17851 4977 17885
rect 317 16916 351 16950
rect 385 16916 419 16950
rect 453 16916 487 16950
rect 521 16916 555 16950
rect 589 16916 623 16950
rect 657 16916 691 16950
rect 725 16916 759 16950
rect 793 16916 827 16950
rect 861 16916 895 16950
rect 929 16916 963 16950
rect 997 16916 1031 16950
rect 1065 16916 1099 16950
rect 1133 16916 1167 16950
rect 1201 16916 1235 16950
rect 1269 16916 1303 16950
rect 199 16806 233 16840
rect 199 16738 233 16772
rect 1387 16806 1421 16840
rect 1387 16738 1421 16772
rect 199 16670 233 16704
rect 1387 16670 1421 16704
rect 317 16560 351 16594
rect 385 16560 419 16594
rect 453 16560 487 16594
rect 521 16560 555 16594
rect 589 16560 623 16594
rect 657 16560 691 16594
rect 725 16560 759 16594
rect 793 16560 827 16594
rect 861 16560 895 16594
rect 929 16560 963 16594
rect 997 16560 1031 16594
rect 1065 16560 1099 16594
rect 1133 16560 1167 16594
rect 1201 16560 1235 16594
rect 1269 16560 1303 16594
rect 2470 16920 2504 16954
rect 2538 16920 2572 16954
rect 2606 16920 2640 16954
rect 2674 16920 2708 16954
rect 2742 16920 2776 16954
rect 2810 16920 2844 16954
rect 2878 16920 2912 16954
rect 2946 16920 2980 16954
rect 3014 16920 3048 16954
rect 3082 16920 3116 16954
rect 3150 16920 3184 16954
rect 3218 16920 3252 16954
rect 3286 16920 3320 16954
rect 3354 16920 3388 16954
rect 3422 16920 3456 16954
rect 2352 16810 2386 16844
rect 3991 16920 4025 16954
rect 4059 16920 4093 16954
rect 4127 16920 4161 16954
rect 4195 16920 4229 16954
rect 4263 16920 4297 16954
rect 4331 16920 4365 16954
rect 4399 16920 4433 16954
rect 4467 16920 4501 16954
rect 4535 16920 4569 16954
rect 4603 16920 4637 16954
rect 4671 16920 4705 16954
rect 4739 16920 4773 16954
rect 4807 16920 4841 16954
rect 4875 16920 4909 16954
rect 4943 16920 4977 16954
rect 2352 16742 2386 16776
rect 3540 16810 3574 16844
rect 3540 16742 3574 16776
rect 3873 16810 3907 16844
rect 2352 16674 2386 16708
rect 3873 16742 3907 16776
rect 3540 16674 3574 16708
rect 2470 16564 2504 16598
rect 2538 16564 2572 16598
rect 2606 16564 2640 16598
rect 2674 16564 2708 16598
rect 2742 16564 2776 16598
rect 2810 16564 2844 16598
rect 2878 16564 2912 16598
rect 2946 16564 2980 16598
rect 3014 16564 3048 16598
rect 3082 16564 3116 16598
rect 3150 16564 3184 16598
rect 3218 16564 3252 16598
rect 3286 16564 3320 16598
rect 3354 16564 3388 16598
rect 3422 16564 3456 16598
rect 5061 16810 5095 16844
rect 5061 16742 5095 16776
rect 3873 16674 3907 16708
rect 5061 16674 5095 16708
rect 3991 16564 4025 16598
rect 4059 16564 4093 16598
rect 4127 16564 4161 16598
rect 4195 16564 4229 16598
rect 4263 16564 4297 16598
rect 4331 16564 4365 16598
rect 4399 16564 4433 16598
rect 4467 16564 4501 16598
rect 4535 16564 4569 16598
rect 4603 16564 4637 16598
rect 4671 16564 4705 16598
rect 4739 16564 4773 16598
rect 4807 16564 4841 16598
rect 4875 16564 4909 16598
rect 4943 16564 4977 16598
rect 317 15629 351 15663
rect 385 15629 419 15663
rect 453 15629 487 15663
rect 521 15629 555 15663
rect 589 15629 623 15663
rect 657 15629 691 15663
rect 725 15629 759 15663
rect 793 15629 827 15663
rect 861 15629 895 15663
rect 929 15629 963 15663
rect 997 15629 1031 15663
rect 1065 15629 1099 15663
rect 1133 15629 1167 15663
rect 1201 15629 1235 15663
rect 1269 15629 1303 15663
rect 199 15519 233 15553
rect 199 15451 233 15485
rect 1387 15519 1421 15553
rect 1387 15451 1421 15485
rect 199 15383 233 15417
rect 1387 15383 1421 15417
rect 317 15273 351 15307
rect 385 15273 419 15307
rect 453 15273 487 15307
rect 521 15273 555 15307
rect 589 15273 623 15307
rect 657 15273 691 15307
rect 725 15273 759 15307
rect 793 15273 827 15307
rect 861 15273 895 15307
rect 929 15273 963 15307
rect 997 15273 1031 15307
rect 1065 15273 1099 15307
rect 1133 15273 1167 15307
rect 1201 15273 1235 15307
rect 1269 15273 1303 15307
rect 2470 15633 2504 15667
rect 2538 15633 2572 15667
rect 2606 15633 2640 15667
rect 2674 15633 2708 15667
rect 2742 15633 2776 15667
rect 2810 15633 2844 15667
rect 2878 15633 2912 15667
rect 2946 15633 2980 15667
rect 3014 15633 3048 15667
rect 3082 15633 3116 15667
rect 3150 15633 3184 15667
rect 3218 15633 3252 15667
rect 3286 15633 3320 15667
rect 3354 15633 3388 15667
rect 3422 15633 3456 15667
rect 2352 15523 2386 15557
rect 3991 15633 4025 15667
rect 4059 15633 4093 15667
rect 4127 15633 4161 15667
rect 4195 15633 4229 15667
rect 4263 15633 4297 15667
rect 4331 15633 4365 15667
rect 4399 15633 4433 15667
rect 4467 15633 4501 15667
rect 4535 15633 4569 15667
rect 4603 15633 4637 15667
rect 4671 15633 4705 15667
rect 4739 15633 4773 15667
rect 4807 15633 4841 15667
rect 4875 15633 4909 15667
rect 4943 15633 4977 15667
rect 2352 15455 2386 15489
rect 3540 15523 3574 15557
rect 3540 15455 3574 15489
rect 3873 15523 3907 15557
rect 2352 15387 2386 15421
rect 3873 15455 3907 15489
rect 3540 15387 3574 15421
rect 2470 15277 2504 15311
rect 2538 15277 2572 15311
rect 2606 15277 2640 15311
rect 2674 15277 2708 15311
rect 2742 15277 2776 15311
rect 2810 15277 2844 15311
rect 2878 15277 2912 15311
rect 2946 15277 2980 15311
rect 3014 15277 3048 15311
rect 3082 15277 3116 15311
rect 3150 15277 3184 15311
rect 3218 15277 3252 15311
rect 3286 15277 3320 15311
rect 3354 15277 3388 15311
rect 3422 15277 3456 15311
rect 5061 15523 5095 15557
rect 5061 15455 5095 15489
rect 3873 15387 3907 15421
rect 5061 15387 5095 15421
rect 3991 15277 4025 15311
rect 4059 15277 4093 15311
rect 4127 15277 4161 15311
rect 4195 15277 4229 15311
rect 4263 15277 4297 15311
rect 4331 15277 4365 15311
rect 4399 15277 4433 15311
rect 4467 15277 4501 15311
rect 4535 15277 4569 15311
rect 4603 15277 4637 15311
rect 4671 15277 4705 15311
rect 4739 15277 4773 15311
rect 4807 15277 4841 15311
rect 4875 15277 4909 15311
rect 4943 15277 4977 15311
rect 317 14342 351 14376
rect 385 14342 419 14376
rect 453 14342 487 14376
rect 521 14342 555 14376
rect 589 14342 623 14376
rect 657 14342 691 14376
rect 725 14342 759 14376
rect 793 14342 827 14376
rect 861 14342 895 14376
rect 929 14342 963 14376
rect 997 14342 1031 14376
rect 1065 14342 1099 14376
rect 1133 14342 1167 14376
rect 1201 14342 1235 14376
rect 1269 14342 1303 14376
rect 199 14232 233 14266
rect 199 14164 233 14198
rect 1387 14232 1421 14266
rect 1387 14164 1421 14198
rect 199 14096 233 14130
rect 1387 14096 1421 14130
rect 317 13986 351 14020
rect 385 13986 419 14020
rect 453 13986 487 14020
rect 521 13986 555 14020
rect 589 13986 623 14020
rect 657 13986 691 14020
rect 725 13986 759 14020
rect 793 13986 827 14020
rect 861 13986 895 14020
rect 929 13986 963 14020
rect 997 13986 1031 14020
rect 1065 13986 1099 14020
rect 1133 13986 1167 14020
rect 1201 13986 1235 14020
rect 1269 13986 1303 14020
rect 2470 14346 2504 14380
rect 2538 14346 2572 14380
rect 2606 14346 2640 14380
rect 2674 14346 2708 14380
rect 2742 14346 2776 14380
rect 2810 14346 2844 14380
rect 2878 14346 2912 14380
rect 2946 14346 2980 14380
rect 3014 14346 3048 14380
rect 3082 14346 3116 14380
rect 3150 14346 3184 14380
rect 3218 14346 3252 14380
rect 3286 14346 3320 14380
rect 3354 14346 3388 14380
rect 3422 14346 3456 14380
rect 2352 14236 2386 14270
rect 3991 14346 4025 14380
rect 4059 14346 4093 14380
rect 4127 14346 4161 14380
rect 4195 14346 4229 14380
rect 4263 14346 4297 14380
rect 4331 14346 4365 14380
rect 4399 14346 4433 14380
rect 4467 14346 4501 14380
rect 4535 14346 4569 14380
rect 4603 14346 4637 14380
rect 4671 14346 4705 14380
rect 4739 14346 4773 14380
rect 4807 14346 4841 14380
rect 4875 14346 4909 14380
rect 4943 14346 4977 14380
rect 2352 14168 2386 14202
rect 3540 14236 3574 14270
rect 3540 14168 3574 14202
rect 3873 14236 3907 14270
rect 2352 14100 2386 14134
rect 3873 14168 3907 14202
rect 3540 14100 3574 14134
rect 2470 13990 2504 14024
rect 2538 13990 2572 14024
rect 2606 13990 2640 14024
rect 2674 13990 2708 14024
rect 2742 13990 2776 14024
rect 2810 13990 2844 14024
rect 2878 13990 2912 14024
rect 2946 13990 2980 14024
rect 3014 13990 3048 14024
rect 3082 13990 3116 14024
rect 3150 13990 3184 14024
rect 3218 13990 3252 14024
rect 3286 13990 3320 14024
rect 3354 13990 3388 14024
rect 3422 13990 3456 14024
rect 5061 14236 5095 14270
rect 5061 14168 5095 14202
rect 3873 14100 3907 14134
rect 5061 14100 5095 14134
rect 3991 13990 4025 14024
rect 4059 13990 4093 14024
rect 4127 13990 4161 14024
rect 4195 13990 4229 14024
rect 4263 13990 4297 14024
rect 4331 13990 4365 14024
rect 4399 13990 4433 14024
rect 4467 13990 4501 14024
rect 4535 13990 4569 14024
rect 4603 13990 4637 14024
rect 4671 13990 4705 14024
rect 4739 13990 4773 14024
rect 4807 13990 4841 14024
rect 4875 13990 4909 14024
rect 4943 13990 4977 14024
rect 317 13055 351 13089
rect 385 13055 419 13089
rect 453 13055 487 13089
rect 521 13055 555 13089
rect 589 13055 623 13089
rect 657 13055 691 13089
rect 725 13055 759 13089
rect 793 13055 827 13089
rect 861 13055 895 13089
rect 929 13055 963 13089
rect 997 13055 1031 13089
rect 1065 13055 1099 13089
rect 1133 13055 1167 13089
rect 1201 13055 1235 13089
rect 1269 13055 1303 13089
rect 199 12945 233 12979
rect 199 12877 233 12911
rect 1387 12945 1421 12979
rect 1387 12877 1421 12911
rect 199 12809 233 12843
rect 1387 12809 1421 12843
rect 317 12699 351 12733
rect 385 12699 419 12733
rect 453 12699 487 12733
rect 521 12699 555 12733
rect 589 12699 623 12733
rect 657 12699 691 12733
rect 725 12699 759 12733
rect 793 12699 827 12733
rect 861 12699 895 12733
rect 929 12699 963 12733
rect 997 12699 1031 12733
rect 1065 12699 1099 12733
rect 1133 12699 1167 12733
rect 1201 12699 1235 12733
rect 1269 12699 1303 12733
rect 2470 13059 2504 13093
rect 2538 13059 2572 13093
rect 2606 13059 2640 13093
rect 2674 13059 2708 13093
rect 2742 13059 2776 13093
rect 2810 13059 2844 13093
rect 2878 13059 2912 13093
rect 2946 13059 2980 13093
rect 3014 13059 3048 13093
rect 3082 13059 3116 13093
rect 3150 13059 3184 13093
rect 3218 13059 3252 13093
rect 3286 13059 3320 13093
rect 3354 13059 3388 13093
rect 3422 13059 3456 13093
rect 2352 12949 2386 12983
rect 3991 13059 4025 13093
rect 4059 13059 4093 13093
rect 4127 13059 4161 13093
rect 4195 13059 4229 13093
rect 4263 13059 4297 13093
rect 4331 13059 4365 13093
rect 4399 13059 4433 13093
rect 4467 13059 4501 13093
rect 4535 13059 4569 13093
rect 4603 13059 4637 13093
rect 4671 13059 4705 13093
rect 4739 13059 4773 13093
rect 4807 13059 4841 13093
rect 4875 13059 4909 13093
rect 4943 13059 4977 13093
rect 2352 12881 2386 12915
rect 3540 12949 3574 12983
rect 3540 12881 3574 12915
rect 3873 12949 3907 12983
rect 2352 12813 2386 12847
rect 3873 12881 3907 12915
rect 3540 12813 3574 12847
rect 2470 12703 2504 12737
rect 2538 12703 2572 12737
rect 2606 12703 2640 12737
rect 2674 12703 2708 12737
rect 2742 12703 2776 12737
rect 2810 12703 2844 12737
rect 2878 12703 2912 12737
rect 2946 12703 2980 12737
rect 3014 12703 3048 12737
rect 3082 12703 3116 12737
rect 3150 12703 3184 12737
rect 3218 12703 3252 12737
rect 3286 12703 3320 12737
rect 3354 12703 3388 12737
rect 3422 12703 3456 12737
rect 5061 12949 5095 12983
rect 5061 12881 5095 12915
rect 3873 12813 3907 12847
rect 5061 12813 5095 12847
rect 3991 12703 4025 12737
rect 4059 12703 4093 12737
rect 4127 12703 4161 12737
rect 4195 12703 4229 12737
rect 4263 12703 4297 12737
rect 4331 12703 4365 12737
rect 4399 12703 4433 12737
rect 4467 12703 4501 12737
rect 4535 12703 4569 12737
rect 4603 12703 4637 12737
rect 4671 12703 4705 12737
rect 4739 12703 4773 12737
rect 4807 12703 4841 12737
rect 4875 12703 4909 12737
rect 4943 12703 4977 12737
rect 317 11768 351 11802
rect 385 11768 419 11802
rect 453 11768 487 11802
rect 521 11768 555 11802
rect 589 11768 623 11802
rect 657 11768 691 11802
rect 725 11768 759 11802
rect 793 11768 827 11802
rect 861 11768 895 11802
rect 929 11768 963 11802
rect 997 11768 1031 11802
rect 1065 11768 1099 11802
rect 1133 11768 1167 11802
rect 1201 11768 1235 11802
rect 1269 11768 1303 11802
rect 199 11658 233 11692
rect 199 11590 233 11624
rect 1387 11658 1421 11692
rect 1387 11590 1421 11624
rect 199 11522 233 11556
rect 1387 11522 1421 11556
rect 317 11412 351 11446
rect 385 11412 419 11446
rect 453 11412 487 11446
rect 521 11412 555 11446
rect 589 11412 623 11446
rect 657 11412 691 11446
rect 725 11412 759 11446
rect 793 11412 827 11446
rect 861 11412 895 11446
rect 929 11412 963 11446
rect 997 11412 1031 11446
rect 1065 11412 1099 11446
rect 1133 11412 1167 11446
rect 1201 11412 1235 11446
rect 1269 11412 1303 11446
rect 2470 11772 2504 11806
rect 2538 11772 2572 11806
rect 2606 11772 2640 11806
rect 2674 11772 2708 11806
rect 2742 11772 2776 11806
rect 2810 11772 2844 11806
rect 2878 11772 2912 11806
rect 2946 11772 2980 11806
rect 3014 11772 3048 11806
rect 3082 11772 3116 11806
rect 3150 11772 3184 11806
rect 3218 11772 3252 11806
rect 3286 11772 3320 11806
rect 3354 11772 3388 11806
rect 3422 11772 3456 11806
rect 2352 11662 2386 11696
rect 3991 11772 4025 11806
rect 4059 11772 4093 11806
rect 4127 11772 4161 11806
rect 4195 11772 4229 11806
rect 4263 11772 4297 11806
rect 4331 11772 4365 11806
rect 4399 11772 4433 11806
rect 4467 11772 4501 11806
rect 4535 11772 4569 11806
rect 4603 11772 4637 11806
rect 4671 11772 4705 11806
rect 4739 11772 4773 11806
rect 4807 11772 4841 11806
rect 4875 11772 4909 11806
rect 4943 11772 4977 11806
rect 2352 11594 2386 11628
rect 3540 11662 3574 11696
rect 3540 11594 3574 11628
rect 3873 11662 3907 11696
rect 2352 11526 2386 11560
rect 3873 11594 3907 11628
rect 3540 11526 3574 11560
rect 2470 11416 2504 11450
rect 2538 11416 2572 11450
rect 2606 11416 2640 11450
rect 2674 11416 2708 11450
rect 2742 11416 2776 11450
rect 2810 11416 2844 11450
rect 2878 11416 2912 11450
rect 2946 11416 2980 11450
rect 3014 11416 3048 11450
rect 3082 11416 3116 11450
rect 3150 11416 3184 11450
rect 3218 11416 3252 11450
rect 3286 11416 3320 11450
rect 3354 11416 3388 11450
rect 3422 11416 3456 11450
rect 5061 11662 5095 11696
rect 5061 11594 5095 11628
rect 3873 11526 3907 11560
rect 5061 11526 5095 11560
rect 3991 11416 4025 11450
rect 4059 11416 4093 11450
rect 4127 11416 4161 11450
rect 4195 11416 4229 11450
rect 4263 11416 4297 11450
rect 4331 11416 4365 11450
rect 4399 11416 4433 11450
rect 4467 11416 4501 11450
rect 4535 11416 4569 11450
rect 4603 11416 4637 11450
rect 4671 11416 4705 11450
rect 4739 11416 4773 11450
rect 4807 11416 4841 11450
rect 4875 11416 4909 11450
rect 4943 11416 4977 11450
rect 317 10481 351 10515
rect 385 10481 419 10515
rect 453 10481 487 10515
rect 521 10481 555 10515
rect 589 10481 623 10515
rect 657 10481 691 10515
rect 725 10481 759 10515
rect 793 10481 827 10515
rect 861 10481 895 10515
rect 929 10481 963 10515
rect 997 10481 1031 10515
rect 1065 10481 1099 10515
rect 1133 10481 1167 10515
rect 1201 10481 1235 10515
rect 1269 10481 1303 10515
rect 199 10371 233 10405
rect 199 10303 233 10337
rect 1387 10371 1421 10405
rect 1387 10303 1421 10337
rect 199 10235 233 10269
rect 1387 10235 1421 10269
rect 317 10125 351 10159
rect 385 10125 419 10159
rect 453 10125 487 10159
rect 521 10125 555 10159
rect 589 10125 623 10159
rect 657 10125 691 10159
rect 725 10125 759 10159
rect 793 10125 827 10159
rect 861 10125 895 10159
rect 929 10125 963 10159
rect 997 10125 1031 10159
rect 1065 10125 1099 10159
rect 1133 10125 1167 10159
rect 1201 10125 1235 10159
rect 1269 10125 1303 10159
rect 2470 10485 2504 10519
rect 2538 10485 2572 10519
rect 2606 10485 2640 10519
rect 2674 10485 2708 10519
rect 2742 10485 2776 10519
rect 2810 10485 2844 10519
rect 2878 10485 2912 10519
rect 2946 10485 2980 10519
rect 3014 10485 3048 10519
rect 3082 10485 3116 10519
rect 3150 10485 3184 10519
rect 3218 10485 3252 10519
rect 3286 10485 3320 10519
rect 3354 10485 3388 10519
rect 3422 10485 3456 10519
rect 2352 10375 2386 10409
rect 3991 10485 4025 10519
rect 4059 10485 4093 10519
rect 4127 10485 4161 10519
rect 4195 10485 4229 10519
rect 4263 10485 4297 10519
rect 4331 10485 4365 10519
rect 4399 10485 4433 10519
rect 4467 10485 4501 10519
rect 4535 10485 4569 10519
rect 4603 10485 4637 10519
rect 4671 10485 4705 10519
rect 4739 10485 4773 10519
rect 4807 10485 4841 10519
rect 4875 10485 4909 10519
rect 4943 10485 4977 10519
rect 2352 10307 2386 10341
rect 3540 10375 3574 10409
rect 3540 10307 3574 10341
rect 3873 10375 3907 10409
rect 2352 10239 2386 10273
rect 3873 10307 3907 10341
rect 3540 10239 3574 10273
rect 2470 10129 2504 10163
rect 2538 10129 2572 10163
rect 2606 10129 2640 10163
rect 2674 10129 2708 10163
rect 2742 10129 2776 10163
rect 2810 10129 2844 10163
rect 2878 10129 2912 10163
rect 2946 10129 2980 10163
rect 3014 10129 3048 10163
rect 3082 10129 3116 10163
rect 3150 10129 3184 10163
rect 3218 10129 3252 10163
rect 3286 10129 3320 10163
rect 3354 10129 3388 10163
rect 3422 10129 3456 10163
rect 5061 10375 5095 10409
rect 5061 10307 5095 10341
rect 3873 10239 3907 10273
rect 5061 10239 5095 10273
rect 3991 10129 4025 10163
rect 4059 10129 4093 10163
rect 4127 10129 4161 10163
rect 4195 10129 4229 10163
rect 4263 10129 4297 10163
rect 4331 10129 4365 10163
rect 4399 10129 4433 10163
rect 4467 10129 4501 10163
rect 4535 10129 4569 10163
rect 4603 10129 4637 10163
rect 4671 10129 4705 10163
rect 4739 10129 4773 10163
rect 4807 10129 4841 10163
rect 4875 10129 4909 10163
rect 4943 10129 4977 10163
rect 317 9194 351 9228
rect 385 9194 419 9228
rect 453 9194 487 9228
rect 521 9194 555 9228
rect 589 9194 623 9228
rect 657 9194 691 9228
rect 725 9194 759 9228
rect 793 9194 827 9228
rect 861 9194 895 9228
rect 929 9194 963 9228
rect 997 9194 1031 9228
rect 1065 9194 1099 9228
rect 1133 9194 1167 9228
rect 1201 9194 1235 9228
rect 1269 9194 1303 9228
rect 199 9084 233 9118
rect 199 9016 233 9050
rect 1387 9084 1421 9118
rect 1387 9016 1421 9050
rect 199 8948 233 8982
rect 1387 8948 1421 8982
rect 317 8838 351 8872
rect 385 8838 419 8872
rect 453 8838 487 8872
rect 521 8838 555 8872
rect 589 8838 623 8872
rect 657 8838 691 8872
rect 725 8838 759 8872
rect 793 8838 827 8872
rect 861 8838 895 8872
rect 929 8838 963 8872
rect 997 8838 1031 8872
rect 1065 8838 1099 8872
rect 1133 8838 1167 8872
rect 1201 8838 1235 8872
rect 1269 8838 1303 8872
rect 2470 9198 2504 9232
rect 2538 9198 2572 9232
rect 2606 9198 2640 9232
rect 2674 9198 2708 9232
rect 2742 9198 2776 9232
rect 2810 9198 2844 9232
rect 2878 9198 2912 9232
rect 2946 9198 2980 9232
rect 3014 9198 3048 9232
rect 3082 9198 3116 9232
rect 3150 9198 3184 9232
rect 3218 9198 3252 9232
rect 3286 9198 3320 9232
rect 3354 9198 3388 9232
rect 3422 9198 3456 9232
rect 2352 9088 2386 9122
rect 3991 9198 4025 9232
rect 4059 9198 4093 9232
rect 4127 9198 4161 9232
rect 4195 9198 4229 9232
rect 4263 9198 4297 9232
rect 4331 9198 4365 9232
rect 4399 9198 4433 9232
rect 4467 9198 4501 9232
rect 4535 9198 4569 9232
rect 4603 9198 4637 9232
rect 4671 9198 4705 9232
rect 4739 9198 4773 9232
rect 4807 9198 4841 9232
rect 4875 9198 4909 9232
rect 4943 9198 4977 9232
rect 2352 9020 2386 9054
rect 3540 9088 3574 9122
rect 3540 9020 3574 9054
rect 3873 9088 3907 9122
rect 2352 8952 2386 8986
rect 3873 9020 3907 9054
rect 3540 8952 3574 8986
rect 2470 8842 2504 8876
rect 2538 8842 2572 8876
rect 2606 8842 2640 8876
rect 2674 8842 2708 8876
rect 2742 8842 2776 8876
rect 2810 8842 2844 8876
rect 2878 8842 2912 8876
rect 2946 8842 2980 8876
rect 3014 8842 3048 8876
rect 3082 8842 3116 8876
rect 3150 8842 3184 8876
rect 3218 8842 3252 8876
rect 3286 8842 3320 8876
rect 3354 8842 3388 8876
rect 3422 8842 3456 8876
rect 5061 9088 5095 9122
rect 5061 9020 5095 9054
rect 3873 8952 3907 8986
rect 5061 8952 5095 8986
rect 3991 8842 4025 8876
rect 4059 8842 4093 8876
rect 4127 8842 4161 8876
rect 4195 8842 4229 8876
rect 4263 8842 4297 8876
rect 4331 8842 4365 8876
rect 4399 8842 4433 8876
rect 4467 8842 4501 8876
rect 4535 8842 4569 8876
rect 4603 8842 4637 8876
rect 4671 8842 4705 8876
rect 4739 8842 4773 8876
rect 4807 8842 4841 8876
rect 4875 8842 4909 8876
rect 4943 8842 4977 8876
rect 317 7907 351 7941
rect 385 7907 419 7941
rect 453 7907 487 7941
rect 521 7907 555 7941
rect 589 7907 623 7941
rect 657 7907 691 7941
rect 725 7907 759 7941
rect 793 7907 827 7941
rect 861 7907 895 7941
rect 929 7907 963 7941
rect 997 7907 1031 7941
rect 1065 7907 1099 7941
rect 1133 7907 1167 7941
rect 1201 7907 1235 7941
rect 1269 7907 1303 7941
rect 199 7797 233 7831
rect 199 7729 233 7763
rect 1387 7797 1421 7831
rect 1387 7729 1421 7763
rect 199 7661 233 7695
rect 1387 7661 1421 7695
rect 317 7551 351 7585
rect 385 7551 419 7585
rect 453 7551 487 7585
rect 521 7551 555 7585
rect 589 7551 623 7585
rect 657 7551 691 7585
rect 725 7551 759 7585
rect 793 7551 827 7585
rect 861 7551 895 7585
rect 929 7551 963 7585
rect 997 7551 1031 7585
rect 1065 7551 1099 7585
rect 1133 7551 1167 7585
rect 1201 7551 1235 7585
rect 1269 7551 1303 7585
rect 2470 7911 2504 7945
rect 2538 7911 2572 7945
rect 2606 7911 2640 7945
rect 2674 7911 2708 7945
rect 2742 7911 2776 7945
rect 2810 7911 2844 7945
rect 2878 7911 2912 7945
rect 2946 7911 2980 7945
rect 3014 7911 3048 7945
rect 3082 7911 3116 7945
rect 3150 7911 3184 7945
rect 3218 7911 3252 7945
rect 3286 7911 3320 7945
rect 3354 7911 3388 7945
rect 3422 7911 3456 7945
rect 2352 7801 2386 7835
rect 3991 7911 4025 7945
rect 4059 7911 4093 7945
rect 4127 7911 4161 7945
rect 4195 7911 4229 7945
rect 4263 7911 4297 7945
rect 4331 7911 4365 7945
rect 4399 7911 4433 7945
rect 4467 7911 4501 7945
rect 4535 7911 4569 7945
rect 4603 7911 4637 7945
rect 4671 7911 4705 7945
rect 4739 7911 4773 7945
rect 4807 7911 4841 7945
rect 4875 7911 4909 7945
rect 4943 7911 4977 7945
rect 2352 7733 2386 7767
rect 3540 7801 3574 7835
rect 3540 7733 3574 7767
rect 3873 7801 3907 7835
rect 2352 7665 2386 7699
rect 3873 7733 3907 7767
rect 3540 7665 3574 7699
rect 2470 7555 2504 7589
rect 2538 7555 2572 7589
rect 2606 7555 2640 7589
rect 2674 7555 2708 7589
rect 2742 7555 2776 7589
rect 2810 7555 2844 7589
rect 2878 7555 2912 7589
rect 2946 7555 2980 7589
rect 3014 7555 3048 7589
rect 3082 7555 3116 7589
rect 3150 7555 3184 7589
rect 3218 7555 3252 7589
rect 3286 7555 3320 7589
rect 3354 7555 3388 7589
rect 3422 7555 3456 7589
rect 5061 7801 5095 7835
rect 5061 7733 5095 7767
rect 3873 7665 3907 7699
rect 5061 7665 5095 7699
rect 3991 7555 4025 7589
rect 4059 7555 4093 7589
rect 4127 7555 4161 7589
rect 4195 7555 4229 7589
rect 4263 7555 4297 7589
rect 4331 7555 4365 7589
rect 4399 7555 4433 7589
rect 4467 7555 4501 7589
rect 4535 7555 4569 7589
rect 4603 7555 4637 7589
rect 4671 7555 4705 7589
rect 4739 7555 4773 7589
rect 4807 7555 4841 7589
rect 4875 7555 4909 7589
rect 4943 7555 4977 7589
rect 317 6620 351 6654
rect 385 6620 419 6654
rect 453 6620 487 6654
rect 521 6620 555 6654
rect 589 6620 623 6654
rect 657 6620 691 6654
rect 725 6620 759 6654
rect 793 6620 827 6654
rect 861 6620 895 6654
rect 929 6620 963 6654
rect 997 6620 1031 6654
rect 1065 6620 1099 6654
rect 1133 6620 1167 6654
rect 1201 6620 1235 6654
rect 1269 6620 1303 6654
rect 199 6510 233 6544
rect 199 6442 233 6476
rect 1387 6510 1421 6544
rect 1387 6442 1421 6476
rect 199 6374 233 6408
rect 1387 6374 1421 6408
rect 317 6264 351 6298
rect 385 6264 419 6298
rect 453 6264 487 6298
rect 521 6264 555 6298
rect 589 6264 623 6298
rect 657 6264 691 6298
rect 725 6264 759 6298
rect 793 6264 827 6298
rect 861 6264 895 6298
rect 929 6264 963 6298
rect 997 6264 1031 6298
rect 1065 6264 1099 6298
rect 1133 6264 1167 6298
rect 1201 6264 1235 6298
rect 1269 6264 1303 6298
rect 2470 6624 2504 6658
rect 2538 6624 2572 6658
rect 2606 6624 2640 6658
rect 2674 6624 2708 6658
rect 2742 6624 2776 6658
rect 2810 6624 2844 6658
rect 2878 6624 2912 6658
rect 2946 6624 2980 6658
rect 3014 6624 3048 6658
rect 3082 6624 3116 6658
rect 3150 6624 3184 6658
rect 3218 6624 3252 6658
rect 3286 6624 3320 6658
rect 3354 6624 3388 6658
rect 3422 6624 3456 6658
rect 2352 6514 2386 6548
rect 3991 6624 4025 6658
rect 4059 6624 4093 6658
rect 4127 6624 4161 6658
rect 4195 6624 4229 6658
rect 4263 6624 4297 6658
rect 4331 6624 4365 6658
rect 4399 6624 4433 6658
rect 4467 6624 4501 6658
rect 4535 6624 4569 6658
rect 4603 6624 4637 6658
rect 4671 6624 4705 6658
rect 4739 6624 4773 6658
rect 4807 6624 4841 6658
rect 4875 6624 4909 6658
rect 4943 6624 4977 6658
rect 2352 6446 2386 6480
rect 3540 6514 3574 6548
rect 3540 6446 3574 6480
rect 3873 6514 3907 6548
rect 2352 6378 2386 6412
rect 3873 6446 3907 6480
rect 3540 6378 3574 6412
rect 2470 6268 2504 6302
rect 2538 6268 2572 6302
rect 2606 6268 2640 6302
rect 2674 6268 2708 6302
rect 2742 6268 2776 6302
rect 2810 6268 2844 6302
rect 2878 6268 2912 6302
rect 2946 6268 2980 6302
rect 3014 6268 3048 6302
rect 3082 6268 3116 6302
rect 3150 6268 3184 6302
rect 3218 6268 3252 6302
rect 3286 6268 3320 6302
rect 3354 6268 3388 6302
rect 3422 6268 3456 6302
rect 5061 6514 5095 6548
rect 5061 6446 5095 6480
rect 3873 6378 3907 6412
rect 5061 6378 5095 6412
rect 3991 6268 4025 6302
rect 4059 6268 4093 6302
rect 4127 6268 4161 6302
rect 4195 6268 4229 6302
rect 4263 6268 4297 6302
rect 4331 6268 4365 6302
rect 4399 6268 4433 6302
rect 4467 6268 4501 6302
rect 4535 6268 4569 6302
rect 4603 6268 4637 6302
rect 4671 6268 4705 6302
rect 4739 6268 4773 6302
rect 4807 6268 4841 6302
rect 4875 6268 4909 6302
rect 4943 6268 4977 6302
rect 317 5333 351 5367
rect 385 5333 419 5367
rect 453 5333 487 5367
rect 521 5333 555 5367
rect 589 5333 623 5367
rect 657 5333 691 5367
rect 725 5333 759 5367
rect 793 5333 827 5367
rect 861 5333 895 5367
rect 929 5333 963 5367
rect 997 5333 1031 5367
rect 1065 5333 1099 5367
rect 1133 5333 1167 5367
rect 1201 5333 1235 5367
rect 1269 5333 1303 5367
rect 199 5223 233 5257
rect 199 5155 233 5189
rect 1387 5223 1421 5257
rect 1387 5155 1421 5189
rect 199 5087 233 5121
rect 1387 5087 1421 5121
rect 317 4977 351 5011
rect 385 4977 419 5011
rect 453 4977 487 5011
rect 521 4977 555 5011
rect 589 4977 623 5011
rect 657 4977 691 5011
rect 725 4977 759 5011
rect 793 4977 827 5011
rect 861 4977 895 5011
rect 929 4977 963 5011
rect 997 4977 1031 5011
rect 1065 4977 1099 5011
rect 1133 4977 1167 5011
rect 1201 4977 1235 5011
rect 1269 4977 1303 5011
rect 2470 5337 2504 5371
rect 2538 5337 2572 5371
rect 2606 5337 2640 5371
rect 2674 5337 2708 5371
rect 2742 5337 2776 5371
rect 2810 5337 2844 5371
rect 2878 5337 2912 5371
rect 2946 5337 2980 5371
rect 3014 5337 3048 5371
rect 3082 5337 3116 5371
rect 3150 5337 3184 5371
rect 3218 5337 3252 5371
rect 3286 5337 3320 5371
rect 3354 5337 3388 5371
rect 3422 5337 3456 5371
rect 2352 5227 2386 5261
rect 3991 5337 4025 5371
rect 4059 5337 4093 5371
rect 4127 5337 4161 5371
rect 4195 5337 4229 5371
rect 4263 5337 4297 5371
rect 4331 5337 4365 5371
rect 4399 5337 4433 5371
rect 4467 5337 4501 5371
rect 4535 5337 4569 5371
rect 4603 5337 4637 5371
rect 4671 5337 4705 5371
rect 4739 5337 4773 5371
rect 4807 5337 4841 5371
rect 4875 5337 4909 5371
rect 4943 5337 4977 5371
rect 2352 5159 2386 5193
rect 3540 5227 3574 5261
rect 3540 5159 3574 5193
rect 3873 5227 3907 5261
rect 2352 5091 2386 5125
rect 3873 5159 3907 5193
rect 3540 5091 3574 5125
rect 2470 4981 2504 5015
rect 2538 4981 2572 5015
rect 2606 4981 2640 5015
rect 2674 4981 2708 5015
rect 2742 4981 2776 5015
rect 2810 4981 2844 5015
rect 2878 4981 2912 5015
rect 2946 4981 2980 5015
rect 3014 4981 3048 5015
rect 3082 4981 3116 5015
rect 3150 4981 3184 5015
rect 3218 4981 3252 5015
rect 3286 4981 3320 5015
rect 3354 4981 3388 5015
rect 3422 4981 3456 5015
rect 5061 5227 5095 5261
rect 5061 5159 5095 5193
rect 3873 5091 3907 5125
rect 5061 5091 5095 5125
rect 3991 4981 4025 5015
rect 4059 4981 4093 5015
rect 4127 4981 4161 5015
rect 4195 4981 4229 5015
rect 4263 4981 4297 5015
rect 4331 4981 4365 5015
rect 4399 4981 4433 5015
rect 4467 4981 4501 5015
rect 4535 4981 4569 5015
rect 4603 4981 4637 5015
rect 4671 4981 4705 5015
rect 4739 4981 4773 5015
rect 4807 4981 4841 5015
rect 4875 4981 4909 5015
rect 4943 4981 4977 5015
rect 317 4046 351 4080
rect 385 4046 419 4080
rect 453 4046 487 4080
rect 521 4046 555 4080
rect 589 4046 623 4080
rect 657 4046 691 4080
rect 725 4046 759 4080
rect 793 4046 827 4080
rect 861 4046 895 4080
rect 929 4046 963 4080
rect 997 4046 1031 4080
rect 1065 4046 1099 4080
rect 1133 4046 1167 4080
rect 1201 4046 1235 4080
rect 1269 4046 1303 4080
rect 199 3936 233 3970
rect 199 3868 233 3902
rect 1387 3936 1421 3970
rect 1387 3868 1421 3902
rect 199 3800 233 3834
rect 1387 3800 1421 3834
rect 317 3690 351 3724
rect 385 3690 419 3724
rect 453 3690 487 3724
rect 521 3690 555 3724
rect 589 3690 623 3724
rect 657 3690 691 3724
rect 725 3690 759 3724
rect 793 3690 827 3724
rect 861 3690 895 3724
rect 929 3690 963 3724
rect 997 3690 1031 3724
rect 1065 3690 1099 3724
rect 1133 3690 1167 3724
rect 1201 3690 1235 3724
rect 1269 3690 1303 3724
rect 2470 4050 2504 4084
rect 2538 4050 2572 4084
rect 2606 4050 2640 4084
rect 2674 4050 2708 4084
rect 2742 4050 2776 4084
rect 2810 4050 2844 4084
rect 2878 4050 2912 4084
rect 2946 4050 2980 4084
rect 3014 4050 3048 4084
rect 3082 4050 3116 4084
rect 3150 4050 3184 4084
rect 3218 4050 3252 4084
rect 3286 4050 3320 4084
rect 3354 4050 3388 4084
rect 3422 4050 3456 4084
rect 2352 3940 2386 3974
rect 3991 4050 4025 4084
rect 4059 4050 4093 4084
rect 4127 4050 4161 4084
rect 4195 4050 4229 4084
rect 4263 4050 4297 4084
rect 4331 4050 4365 4084
rect 4399 4050 4433 4084
rect 4467 4050 4501 4084
rect 4535 4050 4569 4084
rect 4603 4050 4637 4084
rect 4671 4050 4705 4084
rect 4739 4050 4773 4084
rect 4807 4050 4841 4084
rect 4875 4050 4909 4084
rect 4943 4050 4977 4084
rect 2352 3872 2386 3906
rect 3540 3940 3574 3974
rect 3540 3872 3574 3906
rect 3873 3940 3907 3974
rect 2352 3804 2386 3838
rect 3873 3872 3907 3906
rect 3540 3804 3574 3838
rect 2470 3694 2504 3728
rect 2538 3694 2572 3728
rect 2606 3694 2640 3728
rect 2674 3694 2708 3728
rect 2742 3694 2776 3728
rect 2810 3694 2844 3728
rect 2878 3694 2912 3728
rect 2946 3694 2980 3728
rect 3014 3694 3048 3728
rect 3082 3694 3116 3728
rect 3150 3694 3184 3728
rect 3218 3694 3252 3728
rect 3286 3694 3320 3728
rect 3354 3694 3388 3728
rect 3422 3694 3456 3728
rect 5061 3940 5095 3974
rect 5061 3872 5095 3906
rect 3873 3804 3907 3838
rect 5061 3804 5095 3838
rect 3991 3694 4025 3728
rect 4059 3694 4093 3728
rect 4127 3694 4161 3728
rect 4195 3694 4229 3728
rect 4263 3694 4297 3728
rect 4331 3694 4365 3728
rect 4399 3694 4433 3728
rect 4467 3694 4501 3728
rect 4535 3694 4569 3728
rect 4603 3694 4637 3728
rect 4671 3694 4705 3728
rect 4739 3694 4773 3728
rect 4807 3694 4841 3728
rect 4875 3694 4909 3728
rect 4943 3694 4977 3728
rect 317 2759 351 2793
rect 385 2759 419 2793
rect 453 2759 487 2793
rect 521 2759 555 2793
rect 589 2759 623 2793
rect 657 2759 691 2793
rect 725 2759 759 2793
rect 793 2759 827 2793
rect 861 2759 895 2793
rect 929 2759 963 2793
rect 997 2759 1031 2793
rect 1065 2759 1099 2793
rect 1133 2759 1167 2793
rect 1201 2759 1235 2793
rect 1269 2759 1303 2793
rect 199 2649 233 2683
rect 199 2581 233 2615
rect 1387 2649 1421 2683
rect 1387 2581 1421 2615
rect 199 2513 233 2547
rect 1387 2513 1421 2547
rect 317 2403 351 2437
rect 385 2403 419 2437
rect 453 2403 487 2437
rect 521 2403 555 2437
rect 589 2403 623 2437
rect 657 2403 691 2437
rect 725 2403 759 2437
rect 793 2403 827 2437
rect 861 2403 895 2437
rect 929 2403 963 2437
rect 997 2403 1031 2437
rect 1065 2403 1099 2437
rect 1133 2403 1167 2437
rect 1201 2403 1235 2437
rect 1269 2403 1303 2437
rect 2470 2763 2504 2797
rect 2538 2763 2572 2797
rect 2606 2763 2640 2797
rect 2674 2763 2708 2797
rect 2742 2763 2776 2797
rect 2810 2763 2844 2797
rect 2878 2763 2912 2797
rect 2946 2763 2980 2797
rect 3014 2763 3048 2797
rect 3082 2763 3116 2797
rect 3150 2763 3184 2797
rect 3218 2763 3252 2797
rect 3286 2763 3320 2797
rect 3354 2763 3388 2797
rect 3422 2763 3456 2797
rect 2352 2653 2386 2687
rect 3991 2763 4025 2797
rect 4059 2763 4093 2797
rect 4127 2763 4161 2797
rect 4195 2763 4229 2797
rect 4263 2763 4297 2797
rect 4331 2763 4365 2797
rect 4399 2763 4433 2797
rect 4467 2763 4501 2797
rect 4535 2763 4569 2797
rect 4603 2763 4637 2797
rect 4671 2763 4705 2797
rect 4739 2763 4773 2797
rect 4807 2763 4841 2797
rect 4875 2763 4909 2797
rect 4943 2763 4977 2797
rect 2352 2585 2386 2619
rect 3540 2653 3574 2687
rect 3540 2585 3574 2619
rect 3873 2653 3907 2687
rect 2352 2517 2386 2551
rect 3873 2585 3907 2619
rect 3540 2517 3574 2551
rect 2470 2407 2504 2441
rect 2538 2407 2572 2441
rect 2606 2407 2640 2441
rect 2674 2407 2708 2441
rect 2742 2407 2776 2441
rect 2810 2407 2844 2441
rect 2878 2407 2912 2441
rect 2946 2407 2980 2441
rect 3014 2407 3048 2441
rect 3082 2407 3116 2441
rect 3150 2407 3184 2441
rect 3218 2407 3252 2441
rect 3286 2407 3320 2441
rect 3354 2407 3388 2441
rect 3422 2407 3456 2441
rect 5061 2653 5095 2687
rect 5061 2585 5095 2619
rect 3873 2517 3907 2551
rect 5061 2517 5095 2551
rect 3991 2407 4025 2441
rect 4059 2407 4093 2441
rect 4127 2407 4161 2441
rect 4195 2407 4229 2441
rect 4263 2407 4297 2441
rect 4331 2407 4365 2441
rect 4399 2407 4433 2441
rect 4467 2407 4501 2441
rect 4535 2407 4569 2441
rect 4603 2407 4637 2441
rect 4671 2407 4705 2441
rect 4739 2407 4773 2441
rect 4807 2407 4841 2441
rect 4875 2407 4909 2441
rect 4943 2407 4977 2441
rect 317 1472 351 1506
rect 385 1472 419 1506
rect 453 1472 487 1506
rect 521 1472 555 1506
rect 589 1472 623 1506
rect 657 1472 691 1506
rect 725 1472 759 1506
rect 793 1472 827 1506
rect 861 1472 895 1506
rect 929 1472 963 1506
rect 997 1472 1031 1506
rect 1065 1472 1099 1506
rect 1133 1472 1167 1506
rect 1201 1472 1235 1506
rect 1269 1472 1303 1506
rect 199 1362 233 1396
rect 199 1294 233 1328
rect 1387 1362 1421 1396
rect 1387 1294 1421 1328
rect 199 1226 233 1260
rect 1387 1226 1421 1260
rect 317 1116 351 1150
rect 385 1116 419 1150
rect 453 1116 487 1150
rect 521 1116 555 1150
rect 589 1116 623 1150
rect 657 1116 691 1150
rect 725 1116 759 1150
rect 793 1116 827 1150
rect 861 1116 895 1150
rect 929 1116 963 1150
rect 997 1116 1031 1150
rect 1065 1116 1099 1150
rect 1133 1116 1167 1150
rect 1201 1116 1235 1150
rect 1269 1116 1303 1150
rect 2470 1476 2504 1510
rect 2538 1476 2572 1510
rect 2606 1476 2640 1510
rect 2674 1476 2708 1510
rect 2742 1476 2776 1510
rect 2810 1476 2844 1510
rect 2878 1476 2912 1510
rect 2946 1476 2980 1510
rect 3014 1476 3048 1510
rect 3082 1476 3116 1510
rect 3150 1476 3184 1510
rect 3218 1476 3252 1510
rect 3286 1476 3320 1510
rect 3354 1476 3388 1510
rect 3422 1476 3456 1510
rect 2352 1366 2386 1400
rect 3991 1476 4025 1510
rect 4059 1476 4093 1510
rect 4127 1476 4161 1510
rect 4195 1476 4229 1510
rect 4263 1476 4297 1510
rect 4331 1476 4365 1510
rect 4399 1476 4433 1510
rect 4467 1476 4501 1510
rect 4535 1476 4569 1510
rect 4603 1476 4637 1510
rect 4671 1476 4705 1510
rect 4739 1476 4773 1510
rect 4807 1476 4841 1510
rect 4875 1476 4909 1510
rect 4943 1476 4977 1510
rect 2352 1298 2386 1332
rect 3540 1366 3574 1400
rect 3540 1298 3574 1332
rect 3873 1366 3907 1400
rect 2352 1230 2386 1264
rect 3873 1298 3907 1332
rect 3540 1230 3574 1264
rect 2470 1120 2504 1154
rect 2538 1120 2572 1154
rect 2606 1120 2640 1154
rect 2674 1120 2708 1154
rect 2742 1120 2776 1154
rect 2810 1120 2844 1154
rect 2878 1120 2912 1154
rect 2946 1120 2980 1154
rect 3014 1120 3048 1154
rect 3082 1120 3116 1154
rect 3150 1120 3184 1154
rect 3218 1120 3252 1154
rect 3286 1120 3320 1154
rect 3354 1120 3388 1154
rect 3422 1120 3456 1154
rect 5061 1366 5095 1400
rect 5061 1298 5095 1332
rect 3873 1230 3907 1264
rect 5061 1230 5095 1264
rect 3991 1120 4025 1154
rect 4059 1120 4093 1154
rect 4127 1120 4161 1154
rect 4195 1120 4229 1154
rect 4263 1120 4297 1154
rect 4331 1120 4365 1154
rect 4399 1120 4433 1154
rect 4467 1120 4501 1154
rect 4535 1120 4569 1154
rect 4603 1120 4637 1154
rect 4671 1120 4705 1154
rect 4739 1120 4773 1154
rect 4807 1120 4841 1154
rect 4875 1120 4909 1154
rect 4943 1120 4977 1154
<< nsubdiffcont >>
rect 317 42021 351 42055
rect 385 42021 419 42055
rect 453 42021 487 42055
rect 521 42021 555 42055
rect 589 42021 623 42055
rect 657 42021 691 42055
rect 725 42021 759 42055
rect 793 42021 827 42055
rect 861 42021 895 42055
rect 929 42021 963 42055
rect 997 42021 1031 42055
rect 1065 42021 1099 42055
rect 1133 42021 1167 42055
rect 1201 42021 1235 42055
rect 1269 42021 1303 42055
rect 199 41919 233 41953
rect 1387 41919 1421 41953
rect 199 41851 233 41885
rect 199 41783 233 41817
rect 199 41715 233 41749
rect 199 41647 233 41681
rect 199 41579 233 41613
rect 1387 41851 1421 41885
rect 1387 41783 1421 41817
rect 1387 41715 1421 41749
rect 1387 41647 1421 41681
rect 1387 41579 1421 41613
rect 317 41477 351 41511
rect 385 41477 419 41511
rect 453 41477 487 41511
rect 521 41477 555 41511
rect 589 41477 623 41511
rect 657 41477 691 41511
rect 725 41477 759 41511
rect 793 41477 827 41511
rect 861 41477 895 41511
rect 929 41477 963 41511
rect 997 41477 1031 41511
rect 1065 41477 1099 41511
rect 1133 41477 1167 41511
rect 1201 41477 1235 41511
rect 1269 41477 1303 41511
rect 2470 42025 2504 42059
rect 2538 42025 2572 42059
rect 2606 42025 2640 42059
rect 2674 42025 2708 42059
rect 2742 42025 2776 42059
rect 2810 42025 2844 42059
rect 2878 42025 2912 42059
rect 2946 42025 2980 42059
rect 3014 42025 3048 42059
rect 3082 42025 3116 42059
rect 3150 42025 3184 42059
rect 3218 42025 3252 42059
rect 3286 42025 3320 42059
rect 3354 42025 3388 42059
rect 3422 42025 3456 42059
rect 2352 41923 2386 41957
rect 3540 41923 3574 41957
rect 2352 41855 2386 41889
rect 2352 41787 2386 41821
rect 2352 41719 2386 41753
rect 2352 41651 2386 41685
rect 2352 41583 2386 41617
rect 3540 41855 3574 41889
rect 3540 41787 3574 41821
rect 3540 41719 3574 41753
rect 3540 41651 3574 41685
rect 3540 41583 3574 41617
rect 2470 41481 2504 41515
rect 2538 41481 2572 41515
rect 2606 41481 2640 41515
rect 2674 41481 2708 41515
rect 2742 41481 2776 41515
rect 2810 41481 2844 41515
rect 2878 41481 2912 41515
rect 2946 41481 2980 41515
rect 3014 41481 3048 41515
rect 3082 41481 3116 41515
rect 3150 41481 3184 41515
rect 3218 41481 3252 41515
rect 3286 41481 3320 41515
rect 3354 41481 3388 41515
rect 3422 41481 3456 41515
rect 3991 42025 4025 42059
rect 4059 42025 4093 42059
rect 4127 42025 4161 42059
rect 4195 42025 4229 42059
rect 4263 42025 4297 42059
rect 4331 42025 4365 42059
rect 4399 42025 4433 42059
rect 4467 42025 4501 42059
rect 4535 42025 4569 42059
rect 4603 42025 4637 42059
rect 4671 42025 4705 42059
rect 4739 42025 4773 42059
rect 4807 42025 4841 42059
rect 4875 42025 4909 42059
rect 4943 42025 4977 42059
rect 3873 41923 3907 41957
rect 5061 41923 5095 41957
rect 3873 41855 3907 41889
rect 3873 41787 3907 41821
rect 3873 41719 3907 41753
rect 3873 41651 3907 41685
rect 3873 41583 3907 41617
rect 5061 41855 5095 41889
rect 5061 41787 5095 41821
rect 5061 41719 5095 41753
rect 5061 41651 5095 41685
rect 5061 41583 5095 41617
rect 3991 41481 4025 41515
rect 4059 41481 4093 41515
rect 4127 41481 4161 41515
rect 4195 41481 4229 41515
rect 4263 41481 4297 41515
rect 4331 41481 4365 41515
rect 4399 41481 4433 41515
rect 4467 41481 4501 41515
rect 4535 41481 4569 41515
rect 4603 41481 4637 41515
rect 4671 41481 4705 41515
rect 4739 41481 4773 41515
rect 4807 41481 4841 41515
rect 4875 41481 4909 41515
rect 4943 41481 4977 41515
rect 317 40734 351 40768
rect 385 40734 419 40768
rect 453 40734 487 40768
rect 521 40734 555 40768
rect 589 40734 623 40768
rect 657 40734 691 40768
rect 725 40734 759 40768
rect 793 40734 827 40768
rect 861 40734 895 40768
rect 929 40734 963 40768
rect 997 40734 1031 40768
rect 1065 40734 1099 40768
rect 1133 40734 1167 40768
rect 1201 40734 1235 40768
rect 1269 40734 1303 40768
rect 199 40632 233 40666
rect 1387 40632 1421 40666
rect 199 40564 233 40598
rect 199 40496 233 40530
rect 199 40428 233 40462
rect 199 40360 233 40394
rect 199 40292 233 40326
rect 1387 40564 1421 40598
rect 1387 40496 1421 40530
rect 1387 40428 1421 40462
rect 1387 40360 1421 40394
rect 1387 40292 1421 40326
rect 317 40190 351 40224
rect 385 40190 419 40224
rect 453 40190 487 40224
rect 521 40190 555 40224
rect 589 40190 623 40224
rect 657 40190 691 40224
rect 725 40190 759 40224
rect 793 40190 827 40224
rect 861 40190 895 40224
rect 929 40190 963 40224
rect 997 40190 1031 40224
rect 1065 40190 1099 40224
rect 1133 40190 1167 40224
rect 1201 40190 1235 40224
rect 1269 40190 1303 40224
rect 2470 40738 2504 40772
rect 2538 40738 2572 40772
rect 2606 40738 2640 40772
rect 2674 40738 2708 40772
rect 2742 40738 2776 40772
rect 2810 40738 2844 40772
rect 2878 40738 2912 40772
rect 2946 40738 2980 40772
rect 3014 40738 3048 40772
rect 3082 40738 3116 40772
rect 3150 40738 3184 40772
rect 3218 40738 3252 40772
rect 3286 40738 3320 40772
rect 3354 40738 3388 40772
rect 3422 40738 3456 40772
rect 2352 40636 2386 40670
rect 3540 40636 3574 40670
rect 2352 40568 2386 40602
rect 2352 40500 2386 40534
rect 2352 40432 2386 40466
rect 2352 40364 2386 40398
rect 2352 40296 2386 40330
rect 3540 40568 3574 40602
rect 3540 40500 3574 40534
rect 3540 40432 3574 40466
rect 3540 40364 3574 40398
rect 3540 40296 3574 40330
rect 2470 40194 2504 40228
rect 2538 40194 2572 40228
rect 2606 40194 2640 40228
rect 2674 40194 2708 40228
rect 2742 40194 2776 40228
rect 2810 40194 2844 40228
rect 2878 40194 2912 40228
rect 2946 40194 2980 40228
rect 3014 40194 3048 40228
rect 3082 40194 3116 40228
rect 3150 40194 3184 40228
rect 3218 40194 3252 40228
rect 3286 40194 3320 40228
rect 3354 40194 3388 40228
rect 3422 40194 3456 40228
rect 3991 40738 4025 40772
rect 4059 40738 4093 40772
rect 4127 40738 4161 40772
rect 4195 40738 4229 40772
rect 4263 40738 4297 40772
rect 4331 40738 4365 40772
rect 4399 40738 4433 40772
rect 4467 40738 4501 40772
rect 4535 40738 4569 40772
rect 4603 40738 4637 40772
rect 4671 40738 4705 40772
rect 4739 40738 4773 40772
rect 4807 40738 4841 40772
rect 4875 40738 4909 40772
rect 4943 40738 4977 40772
rect 3873 40636 3907 40670
rect 5061 40636 5095 40670
rect 3873 40568 3907 40602
rect 3873 40500 3907 40534
rect 3873 40432 3907 40466
rect 3873 40364 3907 40398
rect 3873 40296 3907 40330
rect 5061 40568 5095 40602
rect 5061 40500 5095 40534
rect 5061 40432 5095 40466
rect 5061 40364 5095 40398
rect 5061 40296 5095 40330
rect 3991 40194 4025 40228
rect 4059 40194 4093 40228
rect 4127 40194 4161 40228
rect 4195 40194 4229 40228
rect 4263 40194 4297 40228
rect 4331 40194 4365 40228
rect 4399 40194 4433 40228
rect 4467 40194 4501 40228
rect 4535 40194 4569 40228
rect 4603 40194 4637 40228
rect 4671 40194 4705 40228
rect 4739 40194 4773 40228
rect 4807 40194 4841 40228
rect 4875 40194 4909 40228
rect 4943 40194 4977 40228
rect 317 39447 351 39481
rect 385 39447 419 39481
rect 453 39447 487 39481
rect 521 39447 555 39481
rect 589 39447 623 39481
rect 657 39447 691 39481
rect 725 39447 759 39481
rect 793 39447 827 39481
rect 861 39447 895 39481
rect 929 39447 963 39481
rect 997 39447 1031 39481
rect 1065 39447 1099 39481
rect 1133 39447 1167 39481
rect 1201 39447 1235 39481
rect 1269 39447 1303 39481
rect 199 39345 233 39379
rect 1387 39345 1421 39379
rect 199 39277 233 39311
rect 199 39209 233 39243
rect 199 39141 233 39175
rect 199 39073 233 39107
rect 199 39005 233 39039
rect 1387 39277 1421 39311
rect 1387 39209 1421 39243
rect 1387 39141 1421 39175
rect 1387 39073 1421 39107
rect 1387 39005 1421 39039
rect 317 38903 351 38937
rect 385 38903 419 38937
rect 453 38903 487 38937
rect 521 38903 555 38937
rect 589 38903 623 38937
rect 657 38903 691 38937
rect 725 38903 759 38937
rect 793 38903 827 38937
rect 861 38903 895 38937
rect 929 38903 963 38937
rect 997 38903 1031 38937
rect 1065 38903 1099 38937
rect 1133 38903 1167 38937
rect 1201 38903 1235 38937
rect 1269 38903 1303 38937
rect 2470 39451 2504 39485
rect 2538 39451 2572 39485
rect 2606 39451 2640 39485
rect 2674 39451 2708 39485
rect 2742 39451 2776 39485
rect 2810 39451 2844 39485
rect 2878 39451 2912 39485
rect 2946 39451 2980 39485
rect 3014 39451 3048 39485
rect 3082 39451 3116 39485
rect 3150 39451 3184 39485
rect 3218 39451 3252 39485
rect 3286 39451 3320 39485
rect 3354 39451 3388 39485
rect 3422 39451 3456 39485
rect 2352 39349 2386 39383
rect 3540 39349 3574 39383
rect 2352 39281 2386 39315
rect 2352 39213 2386 39247
rect 2352 39145 2386 39179
rect 2352 39077 2386 39111
rect 2352 39009 2386 39043
rect 3540 39281 3574 39315
rect 3540 39213 3574 39247
rect 3540 39145 3574 39179
rect 3540 39077 3574 39111
rect 3540 39009 3574 39043
rect 2470 38907 2504 38941
rect 2538 38907 2572 38941
rect 2606 38907 2640 38941
rect 2674 38907 2708 38941
rect 2742 38907 2776 38941
rect 2810 38907 2844 38941
rect 2878 38907 2912 38941
rect 2946 38907 2980 38941
rect 3014 38907 3048 38941
rect 3082 38907 3116 38941
rect 3150 38907 3184 38941
rect 3218 38907 3252 38941
rect 3286 38907 3320 38941
rect 3354 38907 3388 38941
rect 3422 38907 3456 38941
rect 3991 39451 4025 39485
rect 4059 39451 4093 39485
rect 4127 39451 4161 39485
rect 4195 39451 4229 39485
rect 4263 39451 4297 39485
rect 4331 39451 4365 39485
rect 4399 39451 4433 39485
rect 4467 39451 4501 39485
rect 4535 39451 4569 39485
rect 4603 39451 4637 39485
rect 4671 39451 4705 39485
rect 4739 39451 4773 39485
rect 4807 39451 4841 39485
rect 4875 39451 4909 39485
rect 4943 39451 4977 39485
rect 3873 39349 3907 39383
rect 5061 39349 5095 39383
rect 3873 39281 3907 39315
rect 3873 39213 3907 39247
rect 3873 39145 3907 39179
rect 3873 39077 3907 39111
rect 3873 39009 3907 39043
rect 5061 39281 5095 39315
rect 5061 39213 5095 39247
rect 5061 39145 5095 39179
rect 5061 39077 5095 39111
rect 5061 39009 5095 39043
rect 3991 38907 4025 38941
rect 4059 38907 4093 38941
rect 4127 38907 4161 38941
rect 4195 38907 4229 38941
rect 4263 38907 4297 38941
rect 4331 38907 4365 38941
rect 4399 38907 4433 38941
rect 4467 38907 4501 38941
rect 4535 38907 4569 38941
rect 4603 38907 4637 38941
rect 4671 38907 4705 38941
rect 4739 38907 4773 38941
rect 4807 38907 4841 38941
rect 4875 38907 4909 38941
rect 4943 38907 4977 38941
rect 317 38160 351 38194
rect 385 38160 419 38194
rect 453 38160 487 38194
rect 521 38160 555 38194
rect 589 38160 623 38194
rect 657 38160 691 38194
rect 725 38160 759 38194
rect 793 38160 827 38194
rect 861 38160 895 38194
rect 929 38160 963 38194
rect 997 38160 1031 38194
rect 1065 38160 1099 38194
rect 1133 38160 1167 38194
rect 1201 38160 1235 38194
rect 1269 38160 1303 38194
rect 199 38058 233 38092
rect 1387 38058 1421 38092
rect 199 37990 233 38024
rect 199 37922 233 37956
rect 199 37854 233 37888
rect 199 37786 233 37820
rect 199 37718 233 37752
rect 1387 37990 1421 38024
rect 1387 37922 1421 37956
rect 1387 37854 1421 37888
rect 1387 37786 1421 37820
rect 1387 37718 1421 37752
rect 317 37616 351 37650
rect 385 37616 419 37650
rect 453 37616 487 37650
rect 521 37616 555 37650
rect 589 37616 623 37650
rect 657 37616 691 37650
rect 725 37616 759 37650
rect 793 37616 827 37650
rect 861 37616 895 37650
rect 929 37616 963 37650
rect 997 37616 1031 37650
rect 1065 37616 1099 37650
rect 1133 37616 1167 37650
rect 1201 37616 1235 37650
rect 1269 37616 1303 37650
rect 2470 38164 2504 38198
rect 2538 38164 2572 38198
rect 2606 38164 2640 38198
rect 2674 38164 2708 38198
rect 2742 38164 2776 38198
rect 2810 38164 2844 38198
rect 2878 38164 2912 38198
rect 2946 38164 2980 38198
rect 3014 38164 3048 38198
rect 3082 38164 3116 38198
rect 3150 38164 3184 38198
rect 3218 38164 3252 38198
rect 3286 38164 3320 38198
rect 3354 38164 3388 38198
rect 3422 38164 3456 38198
rect 2352 38062 2386 38096
rect 3540 38062 3574 38096
rect 2352 37994 2386 38028
rect 2352 37926 2386 37960
rect 2352 37858 2386 37892
rect 2352 37790 2386 37824
rect 2352 37722 2386 37756
rect 3540 37994 3574 38028
rect 3540 37926 3574 37960
rect 3540 37858 3574 37892
rect 3540 37790 3574 37824
rect 3540 37722 3574 37756
rect 2470 37620 2504 37654
rect 2538 37620 2572 37654
rect 2606 37620 2640 37654
rect 2674 37620 2708 37654
rect 2742 37620 2776 37654
rect 2810 37620 2844 37654
rect 2878 37620 2912 37654
rect 2946 37620 2980 37654
rect 3014 37620 3048 37654
rect 3082 37620 3116 37654
rect 3150 37620 3184 37654
rect 3218 37620 3252 37654
rect 3286 37620 3320 37654
rect 3354 37620 3388 37654
rect 3422 37620 3456 37654
rect 3991 38164 4025 38198
rect 4059 38164 4093 38198
rect 4127 38164 4161 38198
rect 4195 38164 4229 38198
rect 4263 38164 4297 38198
rect 4331 38164 4365 38198
rect 4399 38164 4433 38198
rect 4467 38164 4501 38198
rect 4535 38164 4569 38198
rect 4603 38164 4637 38198
rect 4671 38164 4705 38198
rect 4739 38164 4773 38198
rect 4807 38164 4841 38198
rect 4875 38164 4909 38198
rect 4943 38164 4977 38198
rect 3873 38062 3907 38096
rect 5061 38062 5095 38096
rect 3873 37994 3907 38028
rect 3873 37926 3907 37960
rect 3873 37858 3907 37892
rect 3873 37790 3907 37824
rect 3873 37722 3907 37756
rect 5061 37994 5095 38028
rect 5061 37926 5095 37960
rect 5061 37858 5095 37892
rect 5061 37790 5095 37824
rect 5061 37722 5095 37756
rect 3991 37620 4025 37654
rect 4059 37620 4093 37654
rect 4127 37620 4161 37654
rect 4195 37620 4229 37654
rect 4263 37620 4297 37654
rect 4331 37620 4365 37654
rect 4399 37620 4433 37654
rect 4467 37620 4501 37654
rect 4535 37620 4569 37654
rect 4603 37620 4637 37654
rect 4671 37620 4705 37654
rect 4739 37620 4773 37654
rect 4807 37620 4841 37654
rect 4875 37620 4909 37654
rect 4943 37620 4977 37654
rect 317 36873 351 36907
rect 385 36873 419 36907
rect 453 36873 487 36907
rect 521 36873 555 36907
rect 589 36873 623 36907
rect 657 36873 691 36907
rect 725 36873 759 36907
rect 793 36873 827 36907
rect 861 36873 895 36907
rect 929 36873 963 36907
rect 997 36873 1031 36907
rect 1065 36873 1099 36907
rect 1133 36873 1167 36907
rect 1201 36873 1235 36907
rect 1269 36873 1303 36907
rect 199 36771 233 36805
rect 1387 36771 1421 36805
rect 199 36703 233 36737
rect 199 36635 233 36669
rect 199 36567 233 36601
rect 199 36499 233 36533
rect 199 36431 233 36465
rect 1387 36703 1421 36737
rect 1387 36635 1421 36669
rect 1387 36567 1421 36601
rect 1387 36499 1421 36533
rect 1387 36431 1421 36465
rect 317 36329 351 36363
rect 385 36329 419 36363
rect 453 36329 487 36363
rect 521 36329 555 36363
rect 589 36329 623 36363
rect 657 36329 691 36363
rect 725 36329 759 36363
rect 793 36329 827 36363
rect 861 36329 895 36363
rect 929 36329 963 36363
rect 997 36329 1031 36363
rect 1065 36329 1099 36363
rect 1133 36329 1167 36363
rect 1201 36329 1235 36363
rect 1269 36329 1303 36363
rect 2470 36877 2504 36911
rect 2538 36877 2572 36911
rect 2606 36877 2640 36911
rect 2674 36877 2708 36911
rect 2742 36877 2776 36911
rect 2810 36877 2844 36911
rect 2878 36877 2912 36911
rect 2946 36877 2980 36911
rect 3014 36877 3048 36911
rect 3082 36877 3116 36911
rect 3150 36877 3184 36911
rect 3218 36877 3252 36911
rect 3286 36877 3320 36911
rect 3354 36877 3388 36911
rect 3422 36877 3456 36911
rect 2352 36775 2386 36809
rect 3540 36775 3574 36809
rect 2352 36707 2386 36741
rect 2352 36639 2386 36673
rect 2352 36571 2386 36605
rect 2352 36503 2386 36537
rect 2352 36435 2386 36469
rect 3540 36707 3574 36741
rect 3540 36639 3574 36673
rect 3540 36571 3574 36605
rect 3540 36503 3574 36537
rect 3540 36435 3574 36469
rect 2470 36333 2504 36367
rect 2538 36333 2572 36367
rect 2606 36333 2640 36367
rect 2674 36333 2708 36367
rect 2742 36333 2776 36367
rect 2810 36333 2844 36367
rect 2878 36333 2912 36367
rect 2946 36333 2980 36367
rect 3014 36333 3048 36367
rect 3082 36333 3116 36367
rect 3150 36333 3184 36367
rect 3218 36333 3252 36367
rect 3286 36333 3320 36367
rect 3354 36333 3388 36367
rect 3422 36333 3456 36367
rect 3991 36877 4025 36911
rect 4059 36877 4093 36911
rect 4127 36877 4161 36911
rect 4195 36877 4229 36911
rect 4263 36877 4297 36911
rect 4331 36877 4365 36911
rect 4399 36877 4433 36911
rect 4467 36877 4501 36911
rect 4535 36877 4569 36911
rect 4603 36877 4637 36911
rect 4671 36877 4705 36911
rect 4739 36877 4773 36911
rect 4807 36877 4841 36911
rect 4875 36877 4909 36911
rect 4943 36877 4977 36911
rect 3873 36775 3907 36809
rect 5061 36775 5095 36809
rect 3873 36707 3907 36741
rect 3873 36639 3907 36673
rect 3873 36571 3907 36605
rect 3873 36503 3907 36537
rect 3873 36435 3907 36469
rect 5061 36707 5095 36741
rect 5061 36639 5095 36673
rect 5061 36571 5095 36605
rect 5061 36503 5095 36537
rect 5061 36435 5095 36469
rect 3991 36333 4025 36367
rect 4059 36333 4093 36367
rect 4127 36333 4161 36367
rect 4195 36333 4229 36367
rect 4263 36333 4297 36367
rect 4331 36333 4365 36367
rect 4399 36333 4433 36367
rect 4467 36333 4501 36367
rect 4535 36333 4569 36367
rect 4603 36333 4637 36367
rect 4671 36333 4705 36367
rect 4739 36333 4773 36367
rect 4807 36333 4841 36367
rect 4875 36333 4909 36367
rect 4943 36333 4977 36367
rect 317 35586 351 35620
rect 385 35586 419 35620
rect 453 35586 487 35620
rect 521 35586 555 35620
rect 589 35586 623 35620
rect 657 35586 691 35620
rect 725 35586 759 35620
rect 793 35586 827 35620
rect 861 35586 895 35620
rect 929 35586 963 35620
rect 997 35586 1031 35620
rect 1065 35586 1099 35620
rect 1133 35586 1167 35620
rect 1201 35586 1235 35620
rect 1269 35586 1303 35620
rect 199 35484 233 35518
rect 1387 35484 1421 35518
rect 199 35416 233 35450
rect 199 35348 233 35382
rect 199 35280 233 35314
rect 199 35212 233 35246
rect 199 35144 233 35178
rect 1387 35416 1421 35450
rect 1387 35348 1421 35382
rect 1387 35280 1421 35314
rect 1387 35212 1421 35246
rect 1387 35144 1421 35178
rect 317 35042 351 35076
rect 385 35042 419 35076
rect 453 35042 487 35076
rect 521 35042 555 35076
rect 589 35042 623 35076
rect 657 35042 691 35076
rect 725 35042 759 35076
rect 793 35042 827 35076
rect 861 35042 895 35076
rect 929 35042 963 35076
rect 997 35042 1031 35076
rect 1065 35042 1099 35076
rect 1133 35042 1167 35076
rect 1201 35042 1235 35076
rect 1269 35042 1303 35076
rect 2470 35590 2504 35624
rect 2538 35590 2572 35624
rect 2606 35590 2640 35624
rect 2674 35590 2708 35624
rect 2742 35590 2776 35624
rect 2810 35590 2844 35624
rect 2878 35590 2912 35624
rect 2946 35590 2980 35624
rect 3014 35590 3048 35624
rect 3082 35590 3116 35624
rect 3150 35590 3184 35624
rect 3218 35590 3252 35624
rect 3286 35590 3320 35624
rect 3354 35590 3388 35624
rect 3422 35590 3456 35624
rect 2352 35488 2386 35522
rect 3540 35488 3574 35522
rect 2352 35420 2386 35454
rect 2352 35352 2386 35386
rect 2352 35284 2386 35318
rect 2352 35216 2386 35250
rect 2352 35148 2386 35182
rect 3540 35420 3574 35454
rect 3540 35352 3574 35386
rect 3540 35284 3574 35318
rect 3540 35216 3574 35250
rect 3540 35148 3574 35182
rect 2470 35046 2504 35080
rect 2538 35046 2572 35080
rect 2606 35046 2640 35080
rect 2674 35046 2708 35080
rect 2742 35046 2776 35080
rect 2810 35046 2844 35080
rect 2878 35046 2912 35080
rect 2946 35046 2980 35080
rect 3014 35046 3048 35080
rect 3082 35046 3116 35080
rect 3150 35046 3184 35080
rect 3218 35046 3252 35080
rect 3286 35046 3320 35080
rect 3354 35046 3388 35080
rect 3422 35046 3456 35080
rect 3991 35590 4025 35624
rect 4059 35590 4093 35624
rect 4127 35590 4161 35624
rect 4195 35590 4229 35624
rect 4263 35590 4297 35624
rect 4331 35590 4365 35624
rect 4399 35590 4433 35624
rect 4467 35590 4501 35624
rect 4535 35590 4569 35624
rect 4603 35590 4637 35624
rect 4671 35590 4705 35624
rect 4739 35590 4773 35624
rect 4807 35590 4841 35624
rect 4875 35590 4909 35624
rect 4943 35590 4977 35624
rect 3873 35488 3907 35522
rect 5061 35488 5095 35522
rect 3873 35420 3907 35454
rect 3873 35352 3907 35386
rect 3873 35284 3907 35318
rect 3873 35216 3907 35250
rect 3873 35148 3907 35182
rect 5061 35420 5095 35454
rect 5061 35352 5095 35386
rect 5061 35284 5095 35318
rect 5061 35216 5095 35250
rect 5061 35148 5095 35182
rect 3991 35046 4025 35080
rect 4059 35046 4093 35080
rect 4127 35046 4161 35080
rect 4195 35046 4229 35080
rect 4263 35046 4297 35080
rect 4331 35046 4365 35080
rect 4399 35046 4433 35080
rect 4467 35046 4501 35080
rect 4535 35046 4569 35080
rect 4603 35046 4637 35080
rect 4671 35046 4705 35080
rect 4739 35046 4773 35080
rect 4807 35046 4841 35080
rect 4875 35046 4909 35080
rect 4943 35046 4977 35080
rect 317 34299 351 34333
rect 385 34299 419 34333
rect 453 34299 487 34333
rect 521 34299 555 34333
rect 589 34299 623 34333
rect 657 34299 691 34333
rect 725 34299 759 34333
rect 793 34299 827 34333
rect 861 34299 895 34333
rect 929 34299 963 34333
rect 997 34299 1031 34333
rect 1065 34299 1099 34333
rect 1133 34299 1167 34333
rect 1201 34299 1235 34333
rect 1269 34299 1303 34333
rect 199 34197 233 34231
rect 1387 34197 1421 34231
rect 199 34129 233 34163
rect 199 34061 233 34095
rect 199 33993 233 34027
rect 199 33925 233 33959
rect 199 33857 233 33891
rect 1387 34129 1421 34163
rect 1387 34061 1421 34095
rect 1387 33993 1421 34027
rect 1387 33925 1421 33959
rect 1387 33857 1421 33891
rect 317 33755 351 33789
rect 385 33755 419 33789
rect 453 33755 487 33789
rect 521 33755 555 33789
rect 589 33755 623 33789
rect 657 33755 691 33789
rect 725 33755 759 33789
rect 793 33755 827 33789
rect 861 33755 895 33789
rect 929 33755 963 33789
rect 997 33755 1031 33789
rect 1065 33755 1099 33789
rect 1133 33755 1167 33789
rect 1201 33755 1235 33789
rect 1269 33755 1303 33789
rect 2470 34303 2504 34337
rect 2538 34303 2572 34337
rect 2606 34303 2640 34337
rect 2674 34303 2708 34337
rect 2742 34303 2776 34337
rect 2810 34303 2844 34337
rect 2878 34303 2912 34337
rect 2946 34303 2980 34337
rect 3014 34303 3048 34337
rect 3082 34303 3116 34337
rect 3150 34303 3184 34337
rect 3218 34303 3252 34337
rect 3286 34303 3320 34337
rect 3354 34303 3388 34337
rect 3422 34303 3456 34337
rect 2352 34201 2386 34235
rect 3540 34201 3574 34235
rect 2352 34133 2386 34167
rect 2352 34065 2386 34099
rect 2352 33997 2386 34031
rect 2352 33929 2386 33963
rect 2352 33861 2386 33895
rect 3540 34133 3574 34167
rect 3540 34065 3574 34099
rect 3540 33997 3574 34031
rect 3540 33929 3574 33963
rect 3540 33861 3574 33895
rect 2470 33759 2504 33793
rect 2538 33759 2572 33793
rect 2606 33759 2640 33793
rect 2674 33759 2708 33793
rect 2742 33759 2776 33793
rect 2810 33759 2844 33793
rect 2878 33759 2912 33793
rect 2946 33759 2980 33793
rect 3014 33759 3048 33793
rect 3082 33759 3116 33793
rect 3150 33759 3184 33793
rect 3218 33759 3252 33793
rect 3286 33759 3320 33793
rect 3354 33759 3388 33793
rect 3422 33759 3456 33793
rect 3991 34303 4025 34337
rect 4059 34303 4093 34337
rect 4127 34303 4161 34337
rect 4195 34303 4229 34337
rect 4263 34303 4297 34337
rect 4331 34303 4365 34337
rect 4399 34303 4433 34337
rect 4467 34303 4501 34337
rect 4535 34303 4569 34337
rect 4603 34303 4637 34337
rect 4671 34303 4705 34337
rect 4739 34303 4773 34337
rect 4807 34303 4841 34337
rect 4875 34303 4909 34337
rect 4943 34303 4977 34337
rect 3873 34201 3907 34235
rect 5061 34201 5095 34235
rect 3873 34133 3907 34167
rect 3873 34065 3907 34099
rect 3873 33997 3907 34031
rect 3873 33929 3907 33963
rect 3873 33861 3907 33895
rect 5061 34133 5095 34167
rect 5061 34065 5095 34099
rect 5061 33997 5095 34031
rect 5061 33929 5095 33963
rect 5061 33861 5095 33895
rect 3991 33759 4025 33793
rect 4059 33759 4093 33793
rect 4127 33759 4161 33793
rect 4195 33759 4229 33793
rect 4263 33759 4297 33793
rect 4331 33759 4365 33793
rect 4399 33759 4433 33793
rect 4467 33759 4501 33793
rect 4535 33759 4569 33793
rect 4603 33759 4637 33793
rect 4671 33759 4705 33793
rect 4739 33759 4773 33793
rect 4807 33759 4841 33793
rect 4875 33759 4909 33793
rect 4943 33759 4977 33793
rect 317 33012 351 33046
rect 385 33012 419 33046
rect 453 33012 487 33046
rect 521 33012 555 33046
rect 589 33012 623 33046
rect 657 33012 691 33046
rect 725 33012 759 33046
rect 793 33012 827 33046
rect 861 33012 895 33046
rect 929 33012 963 33046
rect 997 33012 1031 33046
rect 1065 33012 1099 33046
rect 1133 33012 1167 33046
rect 1201 33012 1235 33046
rect 1269 33012 1303 33046
rect 199 32910 233 32944
rect 1387 32910 1421 32944
rect 199 32842 233 32876
rect 199 32774 233 32808
rect 199 32706 233 32740
rect 199 32638 233 32672
rect 199 32570 233 32604
rect 1387 32842 1421 32876
rect 1387 32774 1421 32808
rect 1387 32706 1421 32740
rect 1387 32638 1421 32672
rect 1387 32570 1421 32604
rect 317 32468 351 32502
rect 385 32468 419 32502
rect 453 32468 487 32502
rect 521 32468 555 32502
rect 589 32468 623 32502
rect 657 32468 691 32502
rect 725 32468 759 32502
rect 793 32468 827 32502
rect 861 32468 895 32502
rect 929 32468 963 32502
rect 997 32468 1031 32502
rect 1065 32468 1099 32502
rect 1133 32468 1167 32502
rect 1201 32468 1235 32502
rect 1269 32468 1303 32502
rect 2470 33016 2504 33050
rect 2538 33016 2572 33050
rect 2606 33016 2640 33050
rect 2674 33016 2708 33050
rect 2742 33016 2776 33050
rect 2810 33016 2844 33050
rect 2878 33016 2912 33050
rect 2946 33016 2980 33050
rect 3014 33016 3048 33050
rect 3082 33016 3116 33050
rect 3150 33016 3184 33050
rect 3218 33016 3252 33050
rect 3286 33016 3320 33050
rect 3354 33016 3388 33050
rect 3422 33016 3456 33050
rect 2352 32914 2386 32948
rect 3540 32914 3574 32948
rect 2352 32846 2386 32880
rect 2352 32778 2386 32812
rect 2352 32710 2386 32744
rect 2352 32642 2386 32676
rect 2352 32574 2386 32608
rect 3540 32846 3574 32880
rect 3540 32778 3574 32812
rect 3540 32710 3574 32744
rect 3540 32642 3574 32676
rect 3540 32574 3574 32608
rect 2470 32472 2504 32506
rect 2538 32472 2572 32506
rect 2606 32472 2640 32506
rect 2674 32472 2708 32506
rect 2742 32472 2776 32506
rect 2810 32472 2844 32506
rect 2878 32472 2912 32506
rect 2946 32472 2980 32506
rect 3014 32472 3048 32506
rect 3082 32472 3116 32506
rect 3150 32472 3184 32506
rect 3218 32472 3252 32506
rect 3286 32472 3320 32506
rect 3354 32472 3388 32506
rect 3422 32472 3456 32506
rect 3991 33016 4025 33050
rect 4059 33016 4093 33050
rect 4127 33016 4161 33050
rect 4195 33016 4229 33050
rect 4263 33016 4297 33050
rect 4331 33016 4365 33050
rect 4399 33016 4433 33050
rect 4467 33016 4501 33050
rect 4535 33016 4569 33050
rect 4603 33016 4637 33050
rect 4671 33016 4705 33050
rect 4739 33016 4773 33050
rect 4807 33016 4841 33050
rect 4875 33016 4909 33050
rect 4943 33016 4977 33050
rect 3873 32914 3907 32948
rect 5061 32914 5095 32948
rect 3873 32846 3907 32880
rect 3873 32778 3907 32812
rect 3873 32710 3907 32744
rect 3873 32642 3907 32676
rect 3873 32574 3907 32608
rect 5061 32846 5095 32880
rect 5061 32778 5095 32812
rect 5061 32710 5095 32744
rect 5061 32642 5095 32676
rect 5061 32574 5095 32608
rect 3991 32472 4025 32506
rect 4059 32472 4093 32506
rect 4127 32472 4161 32506
rect 4195 32472 4229 32506
rect 4263 32472 4297 32506
rect 4331 32472 4365 32506
rect 4399 32472 4433 32506
rect 4467 32472 4501 32506
rect 4535 32472 4569 32506
rect 4603 32472 4637 32506
rect 4671 32472 4705 32506
rect 4739 32472 4773 32506
rect 4807 32472 4841 32506
rect 4875 32472 4909 32506
rect 4943 32472 4977 32506
rect 317 31725 351 31759
rect 385 31725 419 31759
rect 453 31725 487 31759
rect 521 31725 555 31759
rect 589 31725 623 31759
rect 657 31725 691 31759
rect 725 31725 759 31759
rect 793 31725 827 31759
rect 861 31725 895 31759
rect 929 31725 963 31759
rect 997 31725 1031 31759
rect 1065 31725 1099 31759
rect 1133 31725 1167 31759
rect 1201 31725 1235 31759
rect 1269 31725 1303 31759
rect 199 31623 233 31657
rect 1387 31623 1421 31657
rect 199 31555 233 31589
rect 199 31487 233 31521
rect 199 31419 233 31453
rect 199 31351 233 31385
rect 199 31283 233 31317
rect 1387 31555 1421 31589
rect 1387 31487 1421 31521
rect 1387 31419 1421 31453
rect 1387 31351 1421 31385
rect 1387 31283 1421 31317
rect 317 31181 351 31215
rect 385 31181 419 31215
rect 453 31181 487 31215
rect 521 31181 555 31215
rect 589 31181 623 31215
rect 657 31181 691 31215
rect 725 31181 759 31215
rect 793 31181 827 31215
rect 861 31181 895 31215
rect 929 31181 963 31215
rect 997 31181 1031 31215
rect 1065 31181 1099 31215
rect 1133 31181 1167 31215
rect 1201 31181 1235 31215
rect 1269 31181 1303 31215
rect 2470 31729 2504 31763
rect 2538 31729 2572 31763
rect 2606 31729 2640 31763
rect 2674 31729 2708 31763
rect 2742 31729 2776 31763
rect 2810 31729 2844 31763
rect 2878 31729 2912 31763
rect 2946 31729 2980 31763
rect 3014 31729 3048 31763
rect 3082 31729 3116 31763
rect 3150 31729 3184 31763
rect 3218 31729 3252 31763
rect 3286 31729 3320 31763
rect 3354 31729 3388 31763
rect 3422 31729 3456 31763
rect 2352 31627 2386 31661
rect 3540 31627 3574 31661
rect 2352 31559 2386 31593
rect 2352 31491 2386 31525
rect 2352 31423 2386 31457
rect 2352 31355 2386 31389
rect 2352 31287 2386 31321
rect 3540 31559 3574 31593
rect 3540 31491 3574 31525
rect 3540 31423 3574 31457
rect 3540 31355 3574 31389
rect 3540 31287 3574 31321
rect 2470 31185 2504 31219
rect 2538 31185 2572 31219
rect 2606 31185 2640 31219
rect 2674 31185 2708 31219
rect 2742 31185 2776 31219
rect 2810 31185 2844 31219
rect 2878 31185 2912 31219
rect 2946 31185 2980 31219
rect 3014 31185 3048 31219
rect 3082 31185 3116 31219
rect 3150 31185 3184 31219
rect 3218 31185 3252 31219
rect 3286 31185 3320 31219
rect 3354 31185 3388 31219
rect 3422 31185 3456 31219
rect 3991 31729 4025 31763
rect 4059 31729 4093 31763
rect 4127 31729 4161 31763
rect 4195 31729 4229 31763
rect 4263 31729 4297 31763
rect 4331 31729 4365 31763
rect 4399 31729 4433 31763
rect 4467 31729 4501 31763
rect 4535 31729 4569 31763
rect 4603 31729 4637 31763
rect 4671 31729 4705 31763
rect 4739 31729 4773 31763
rect 4807 31729 4841 31763
rect 4875 31729 4909 31763
rect 4943 31729 4977 31763
rect 3873 31627 3907 31661
rect 5061 31627 5095 31661
rect 3873 31559 3907 31593
rect 3873 31491 3907 31525
rect 3873 31423 3907 31457
rect 3873 31355 3907 31389
rect 3873 31287 3907 31321
rect 5061 31559 5095 31593
rect 5061 31491 5095 31525
rect 5061 31423 5095 31457
rect 5061 31355 5095 31389
rect 5061 31287 5095 31321
rect 3991 31185 4025 31219
rect 4059 31185 4093 31219
rect 4127 31185 4161 31219
rect 4195 31185 4229 31219
rect 4263 31185 4297 31219
rect 4331 31185 4365 31219
rect 4399 31185 4433 31219
rect 4467 31185 4501 31219
rect 4535 31185 4569 31219
rect 4603 31185 4637 31219
rect 4671 31185 4705 31219
rect 4739 31185 4773 31219
rect 4807 31185 4841 31219
rect 4875 31185 4909 31219
rect 4943 31185 4977 31219
rect 317 30438 351 30472
rect 385 30438 419 30472
rect 453 30438 487 30472
rect 521 30438 555 30472
rect 589 30438 623 30472
rect 657 30438 691 30472
rect 725 30438 759 30472
rect 793 30438 827 30472
rect 861 30438 895 30472
rect 929 30438 963 30472
rect 997 30438 1031 30472
rect 1065 30438 1099 30472
rect 1133 30438 1167 30472
rect 1201 30438 1235 30472
rect 1269 30438 1303 30472
rect 199 30336 233 30370
rect 1387 30336 1421 30370
rect 199 30268 233 30302
rect 199 30200 233 30234
rect 199 30132 233 30166
rect 199 30064 233 30098
rect 199 29996 233 30030
rect 1387 30268 1421 30302
rect 1387 30200 1421 30234
rect 1387 30132 1421 30166
rect 1387 30064 1421 30098
rect 1387 29996 1421 30030
rect 317 29894 351 29928
rect 385 29894 419 29928
rect 453 29894 487 29928
rect 521 29894 555 29928
rect 589 29894 623 29928
rect 657 29894 691 29928
rect 725 29894 759 29928
rect 793 29894 827 29928
rect 861 29894 895 29928
rect 929 29894 963 29928
rect 997 29894 1031 29928
rect 1065 29894 1099 29928
rect 1133 29894 1167 29928
rect 1201 29894 1235 29928
rect 1269 29894 1303 29928
rect 2470 30442 2504 30476
rect 2538 30442 2572 30476
rect 2606 30442 2640 30476
rect 2674 30442 2708 30476
rect 2742 30442 2776 30476
rect 2810 30442 2844 30476
rect 2878 30442 2912 30476
rect 2946 30442 2980 30476
rect 3014 30442 3048 30476
rect 3082 30442 3116 30476
rect 3150 30442 3184 30476
rect 3218 30442 3252 30476
rect 3286 30442 3320 30476
rect 3354 30442 3388 30476
rect 3422 30442 3456 30476
rect 2352 30340 2386 30374
rect 3540 30340 3574 30374
rect 2352 30272 2386 30306
rect 2352 30204 2386 30238
rect 2352 30136 2386 30170
rect 2352 30068 2386 30102
rect 2352 30000 2386 30034
rect 3540 30272 3574 30306
rect 3540 30204 3574 30238
rect 3540 30136 3574 30170
rect 3540 30068 3574 30102
rect 3540 30000 3574 30034
rect 2470 29898 2504 29932
rect 2538 29898 2572 29932
rect 2606 29898 2640 29932
rect 2674 29898 2708 29932
rect 2742 29898 2776 29932
rect 2810 29898 2844 29932
rect 2878 29898 2912 29932
rect 2946 29898 2980 29932
rect 3014 29898 3048 29932
rect 3082 29898 3116 29932
rect 3150 29898 3184 29932
rect 3218 29898 3252 29932
rect 3286 29898 3320 29932
rect 3354 29898 3388 29932
rect 3422 29898 3456 29932
rect 3991 30442 4025 30476
rect 4059 30442 4093 30476
rect 4127 30442 4161 30476
rect 4195 30442 4229 30476
rect 4263 30442 4297 30476
rect 4331 30442 4365 30476
rect 4399 30442 4433 30476
rect 4467 30442 4501 30476
rect 4535 30442 4569 30476
rect 4603 30442 4637 30476
rect 4671 30442 4705 30476
rect 4739 30442 4773 30476
rect 4807 30442 4841 30476
rect 4875 30442 4909 30476
rect 4943 30442 4977 30476
rect 3873 30340 3907 30374
rect 5061 30340 5095 30374
rect 3873 30272 3907 30306
rect 3873 30204 3907 30238
rect 3873 30136 3907 30170
rect 3873 30068 3907 30102
rect 3873 30000 3907 30034
rect 5061 30272 5095 30306
rect 5061 30204 5095 30238
rect 5061 30136 5095 30170
rect 5061 30068 5095 30102
rect 5061 30000 5095 30034
rect 3991 29898 4025 29932
rect 4059 29898 4093 29932
rect 4127 29898 4161 29932
rect 4195 29898 4229 29932
rect 4263 29898 4297 29932
rect 4331 29898 4365 29932
rect 4399 29898 4433 29932
rect 4467 29898 4501 29932
rect 4535 29898 4569 29932
rect 4603 29898 4637 29932
rect 4671 29898 4705 29932
rect 4739 29898 4773 29932
rect 4807 29898 4841 29932
rect 4875 29898 4909 29932
rect 4943 29898 4977 29932
rect 317 29151 351 29185
rect 385 29151 419 29185
rect 453 29151 487 29185
rect 521 29151 555 29185
rect 589 29151 623 29185
rect 657 29151 691 29185
rect 725 29151 759 29185
rect 793 29151 827 29185
rect 861 29151 895 29185
rect 929 29151 963 29185
rect 997 29151 1031 29185
rect 1065 29151 1099 29185
rect 1133 29151 1167 29185
rect 1201 29151 1235 29185
rect 1269 29151 1303 29185
rect 199 29049 233 29083
rect 1387 29049 1421 29083
rect 199 28981 233 29015
rect 199 28913 233 28947
rect 199 28845 233 28879
rect 199 28777 233 28811
rect 199 28709 233 28743
rect 1387 28981 1421 29015
rect 1387 28913 1421 28947
rect 1387 28845 1421 28879
rect 1387 28777 1421 28811
rect 1387 28709 1421 28743
rect 317 28607 351 28641
rect 385 28607 419 28641
rect 453 28607 487 28641
rect 521 28607 555 28641
rect 589 28607 623 28641
rect 657 28607 691 28641
rect 725 28607 759 28641
rect 793 28607 827 28641
rect 861 28607 895 28641
rect 929 28607 963 28641
rect 997 28607 1031 28641
rect 1065 28607 1099 28641
rect 1133 28607 1167 28641
rect 1201 28607 1235 28641
rect 1269 28607 1303 28641
rect 2470 29155 2504 29189
rect 2538 29155 2572 29189
rect 2606 29155 2640 29189
rect 2674 29155 2708 29189
rect 2742 29155 2776 29189
rect 2810 29155 2844 29189
rect 2878 29155 2912 29189
rect 2946 29155 2980 29189
rect 3014 29155 3048 29189
rect 3082 29155 3116 29189
rect 3150 29155 3184 29189
rect 3218 29155 3252 29189
rect 3286 29155 3320 29189
rect 3354 29155 3388 29189
rect 3422 29155 3456 29189
rect 2352 29053 2386 29087
rect 3540 29053 3574 29087
rect 2352 28985 2386 29019
rect 2352 28917 2386 28951
rect 2352 28849 2386 28883
rect 2352 28781 2386 28815
rect 2352 28713 2386 28747
rect 3540 28985 3574 29019
rect 3540 28917 3574 28951
rect 3540 28849 3574 28883
rect 3540 28781 3574 28815
rect 3540 28713 3574 28747
rect 2470 28611 2504 28645
rect 2538 28611 2572 28645
rect 2606 28611 2640 28645
rect 2674 28611 2708 28645
rect 2742 28611 2776 28645
rect 2810 28611 2844 28645
rect 2878 28611 2912 28645
rect 2946 28611 2980 28645
rect 3014 28611 3048 28645
rect 3082 28611 3116 28645
rect 3150 28611 3184 28645
rect 3218 28611 3252 28645
rect 3286 28611 3320 28645
rect 3354 28611 3388 28645
rect 3422 28611 3456 28645
rect 3991 29155 4025 29189
rect 4059 29155 4093 29189
rect 4127 29155 4161 29189
rect 4195 29155 4229 29189
rect 4263 29155 4297 29189
rect 4331 29155 4365 29189
rect 4399 29155 4433 29189
rect 4467 29155 4501 29189
rect 4535 29155 4569 29189
rect 4603 29155 4637 29189
rect 4671 29155 4705 29189
rect 4739 29155 4773 29189
rect 4807 29155 4841 29189
rect 4875 29155 4909 29189
rect 4943 29155 4977 29189
rect 3873 29053 3907 29087
rect 5061 29053 5095 29087
rect 3873 28985 3907 29019
rect 3873 28917 3907 28951
rect 3873 28849 3907 28883
rect 3873 28781 3907 28815
rect 3873 28713 3907 28747
rect 5061 28985 5095 29019
rect 5061 28917 5095 28951
rect 5061 28849 5095 28883
rect 5061 28781 5095 28815
rect 5061 28713 5095 28747
rect 3991 28611 4025 28645
rect 4059 28611 4093 28645
rect 4127 28611 4161 28645
rect 4195 28611 4229 28645
rect 4263 28611 4297 28645
rect 4331 28611 4365 28645
rect 4399 28611 4433 28645
rect 4467 28611 4501 28645
rect 4535 28611 4569 28645
rect 4603 28611 4637 28645
rect 4671 28611 4705 28645
rect 4739 28611 4773 28645
rect 4807 28611 4841 28645
rect 4875 28611 4909 28645
rect 4943 28611 4977 28645
rect 317 27864 351 27898
rect 385 27864 419 27898
rect 453 27864 487 27898
rect 521 27864 555 27898
rect 589 27864 623 27898
rect 657 27864 691 27898
rect 725 27864 759 27898
rect 793 27864 827 27898
rect 861 27864 895 27898
rect 929 27864 963 27898
rect 997 27864 1031 27898
rect 1065 27864 1099 27898
rect 1133 27864 1167 27898
rect 1201 27864 1235 27898
rect 1269 27864 1303 27898
rect 199 27762 233 27796
rect 1387 27762 1421 27796
rect 199 27694 233 27728
rect 199 27626 233 27660
rect 199 27558 233 27592
rect 199 27490 233 27524
rect 199 27422 233 27456
rect 1387 27694 1421 27728
rect 1387 27626 1421 27660
rect 1387 27558 1421 27592
rect 1387 27490 1421 27524
rect 1387 27422 1421 27456
rect 317 27320 351 27354
rect 385 27320 419 27354
rect 453 27320 487 27354
rect 521 27320 555 27354
rect 589 27320 623 27354
rect 657 27320 691 27354
rect 725 27320 759 27354
rect 793 27320 827 27354
rect 861 27320 895 27354
rect 929 27320 963 27354
rect 997 27320 1031 27354
rect 1065 27320 1099 27354
rect 1133 27320 1167 27354
rect 1201 27320 1235 27354
rect 1269 27320 1303 27354
rect 2470 27868 2504 27902
rect 2538 27868 2572 27902
rect 2606 27868 2640 27902
rect 2674 27868 2708 27902
rect 2742 27868 2776 27902
rect 2810 27868 2844 27902
rect 2878 27868 2912 27902
rect 2946 27868 2980 27902
rect 3014 27868 3048 27902
rect 3082 27868 3116 27902
rect 3150 27868 3184 27902
rect 3218 27868 3252 27902
rect 3286 27868 3320 27902
rect 3354 27868 3388 27902
rect 3422 27868 3456 27902
rect 2352 27766 2386 27800
rect 3540 27766 3574 27800
rect 2352 27698 2386 27732
rect 2352 27630 2386 27664
rect 2352 27562 2386 27596
rect 2352 27494 2386 27528
rect 2352 27426 2386 27460
rect 3540 27698 3574 27732
rect 3540 27630 3574 27664
rect 3540 27562 3574 27596
rect 3540 27494 3574 27528
rect 3540 27426 3574 27460
rect 2470 27324 2504 27358
rect 2538 27324 2572 27358
rect 2606 27324 2640 27358
rect 2674 27324 2708 27358
rect 2742 27324 2776 27358
rect 2810 27324 2844 27358
rect 2878 27324 2912 27358
rect 2946 27324 2980 27358
rect 3014 27324 3048 27358
rect 3082 27324 3116 27358
rect 3150 27324 3184 27358
rect 3218 27324 3252 27358
rect 3286 27324 3320 27358
rect 3354 27324 3388 27358
rect 3422 27324 3456 27358
rect 3991 27868 4025 27902
rect 4059 27868 4093 27902
rect 4127 27868 4161 27902
rect 4195 27868 4229 27902
rect 4263 27868 4297 27902
rect 4331 27868 4365 27902
rect 4399 27868 4433 27902
rect 4467 27868 4501 27902
rect 4535 27868 4569 27902
rect 4603 27868 4637 27902
rect 4671 27868 4705 27902
rect 4739 27868 4773 27902
rect 4807 27868 4841 27902
rect 4875 27868 4909 27902
rect 4943 27868 4977 27902
rect 3873 27766 3907 27800
rect 5061 27766 5095 27800
rect 3873 27698 3907 27732
rect 3873 27630 3907 27664
rect 3873 27562 3907 27596
rect 3873 27494 3907 27528
rect 3873 27426 3907 27460
rect 5061 27698 5095 27732
rect 5061 27630 5095 27664
rect 5061 27562 5095 27596
rect 5061 27494 5095 27528
rect 5061 27426 5095 27460
rect 3991 27324 4025 27358
rect 4059 27324 4093 27358
rect 4127 27324 4161 27358
rect 4195 27324 4229 27358
rect 4263 27324 4297 27358
rect 4331 27324 4365 27358
rect 4399 27324 4433 27358
rect 4467 27324 4501 27358
rect 4535 27324 4569 27358
rect 4603 27324 4637 27358
rect 4671 27324 4705 27358
rect 4739 27324 4773 27358
rect 4807 27324 4841 27358
rect 4875 27324 4909 27358
rect 4943 27324 4977 27358
rect 317 26577 351 26611
rect 385 26577 419 26611
rect 453 26577 487 26611
rect 521 26577 555 26611
rect 589 26577 623 26611
rect 657 26577 691 26611
rect 725 26577 759 26611
rect 793 26577 827 26611
rect 861 26577 895 26611
rect 929 26577 963 26611
rect 997 26577 1031 26611
rect 1065 26577 1099 26611
rect 1133 26577 1167 26611
rect 1201 26577 1235 26611
rect 1269 26577 1303 26611
rect 199 26475 233 26509
rect 1387 26475 1421 26509
rect 199 26407 233 26441
rect 199 26339 233 26373
rect 199 26271 233 26305
rect 199 26203 233 26237
rect 199 26135 233 26169
rect 1387 26407 1421 26441
rect 1387 26339 1421 26373
rect 1387 26271 1421 26305
rect 1387 26203 1421 26237
rect 1387 26135 1421 26169
rect 317 26033 351 26067
rect 385 26033 419 26067
rect 453 26033 487 26067
rect 521 26033 555 26067
rect 589 26033 623 26067
rect 657 26033 691 26067
rect 725 26033 759 26067
rect 793 26033 827 26067
rect 861 26033 895 26067
rect 929 26033 963 26067
rect 997 26033 1031 26067
rect 1065 26033 1099 26067
rect 1133 26033 1167 26067
rect 1201 26033 1235 26067
rect 1269 26033 1303 26067
rect 2470 26581 2504 26615
rect 2538 26581 2572 26615
rect 2606 26581 2640 26615
rect 2674 26581 2708 26615
rect 2742 26581 2776 26615
rect 2810 26581 2844 26615
rect 2878 26581 2912 26615
rect 2946 26581 2980 26615
rect 3014 26581 3048 26615
rect 3082 26581 3116 26615
rect 3150 26581 3184 26615
rect 3218 26581 3252 26615
rect 3286 26581 3320 26615
rect 3354 26581 3388 26615
rect 3422 26581 3456 26615
rect 2352 26479 2386 26513
rect 3540 26479 3574 26513
rect 2352 26411 2386 26445
rect 2352 26343 2386 26377
rect 2352 26275 2386 26309
rect 2352 26207 2386 26241
rect 2352 26139 2386 26173
rect 3540 26411 3574 26445
rect 3540 26343 3574 26377
rect 3540 26275 3574 26309
rect 3540 26207 3574 26241
rect 3540 26139 3574 26173
rect 2470 26037 2504 26071
rect 2538 26037 2572 26071
rect 2606 26037 2640 26071
rect 2674 26037 2708 26071
rect 2742 26037 2776 26071
rect 2810 26037 2844 26071
rect 2878 26037 2912 26071
rect 2946 26037 2980 26071
rect 3014 26037 3048 26071
rect 3082 26037 3116 26071
rect 3150 26037 3184 26071
rect 3218 26037 3252 26071
rect 3286 26037 3320 26071
rect 3354 26037 3388 26071
rect 3422 26037 3456 26071
rect 3991 26581 4025 26615
rect 4059 26581 4093 26615
rect 4127 26581 4161 26615
rect 4195 26581 4229 26615
rect 4263 26581 4297 26615
rect 4331 26581 4365 26615
rect 4399 26581 4433 26615
rect 4467 26581 4501 26615
rect 4535 26581 4569 26615
rect 4603 26581 4637 26615
rect 4671 26581 4705 26615
rect 4739 26581 4773 26615
rect 4807 26581 4841 26615
rect 4875 26581 4909 26615
rect 4943 26581 4977 26615
rect 3873 26479 3907 26513
rect 5061 26479 5095 26513
rect 3873 26411 3907 26445
rect 3873 26343 3907 26377
rect 3873 26275 3907 26309
rect 3873 26207 3907 26241
rect 3873 26139 3907 26173
rect 5061 26411 5095 26445
rect 5061 26343 5095 26377
rect 5061 26275 5095 26309
rect 5061 26207 5095 26241
rect 5061 26139 5095 26173
rect 3991 26037 4025 26071
rect 4059 26037 4093 26071
rect 4127 26037 4161 26071
rect 4195 26037 4229 26071
rect 4263 26037 4297 26071
rect 4331 26037 4365 26071
rect 4399 26037 4433 26071
rect 4467 26037 4501 26071
rect 4535 26037 4569 26071
rect 4603 26037 4637 26071
rect 4671 26037 4705 26071
rect 4739 26037 4773 26071
rect 4807 26037 4841 26071
rect 4875 26037 4909 26071
rect 4943 26037 4977 26071
rect 317 25290 351 25324
rect 385 25290 419 25324
rect 453 25290 487 25324
rect 521 25290 555 25324
rect 589 25290 623 25324
rect 657 25290 691 25324
rect 725 25290 759 25324
rect 793 25290 827 25324
rect 861 25290 895 25324
rect 929 25290 963 25324
rect 997 25290 1031 25324
rect 1065 25290 1099 25324
rect 1133 25290 1167 25324
rect 1201 25290 1235 25324
rect 1269 25290 1303 25324
rect 199 25188 233 25222
rect 1387 25188 1421 25222
rect 199 25120 233 25154
rect 199 25052 233 25086
rect 199 24984 233 25018
rect 199 24916 233 24950
rect 199 24848 233 24882
rect 1387 25120 1421 25154
rect 1387 25052 1421 25086
rect 1387 24984 1421 25018
rect 1387 24916 1421 24950
rect 1387 24848 1421 24882
rect 317 24746 351 24780
rect 385 24746 419 24780
rect 453 24746 487 24780
rect 521 24746 555 24780
rect 589 24746 623 24780
rect 657 24746 691 24780
rect 725 24746 759 24780
rect 793 24746 827 24780
rect 861 24746 895 24780
rect 929 24746 963 24780
rect 997 24746 1031 24780
rect 1065 24746 1099 24780
rect 1133 24746 1167 24780
rect 1201 24746 1235 24780
rect 1269 24746 1303 24780
rect 2470 25294 2504 25328
rect 2538 25294 2572 25328
rect 2606 25294 2640 25328
rect 2674 25294 2708 25328
rect 2742 25294 2776 25328
rect 2810 25294 2844 25328
rect 2878 25294 2912 25328
rect 2946 25294 2980 25328
rect 3014 25294 3048 25328
rect 3082 25294 3116 25328
rect 3150 25294 3184 25328
rect 3218 25294 3252 25328
rect 3286 25294 3320 25328
rect 3354 25294 3388 25328
rect 3422 25294 3456 25328
rect 2352 25192 2386 25226
rect 3540 25192 3574 25226
rect 2352 25124 2386 25158
rect 2352 25056 2386 25090
rect 2352 24988 2386 25022
rect 2352 24920 2386 24954
rect 2352 24852 2386 24886
rect 3540 25124 3574 25158
rect 3540 25056 3574 25090
rect 3540 24988 3574 25022
rect 3540 24920 3574 24954
rect 3540 24852 3574 24886
rect 2470 24750 2504 24784
rect 2538 24750 2572 24784
rect 2606 24750 2640 24784
rect 2674 24750 2708 24784
rect 2742 24750 2776 24784
rect 2810 24750 2844 24784
rect 2878 24750 2912 24784
rect 2946 24750 2980 24784
rect 3014 24750 3048 24784
rect 3082 24750 3116 24784
rect 3150 24750 3184 24784
rect 3218 24750 3252 24784
rect 3286 24750 3320 24784
rect 3354 24750 3388 24784
rect 3422 24750 3456 24784
rect 3991 25294 4025 25328
rect 4059 25294 4093 25328
rect 4127 25294 4161 25328
rect 4195 25294 4229 25328
rect 4263 25294 4297 25328
rect 4331 25294 4365 25328
rect 4399 25294 4433 25328
rect 4467 25294 4501 25328
rect 4535 25294 4569 25328
rect 4603 25294 4637 25328
rect 4671 25294 4705 25328
rect 4739 25294 4773 25328
rect 4807 25294 4841 25328
rect 4875 25294 4909 25328
rect 4943 25294 4977 25328
rect 3873 25192 3907 25226
rect 5061 25192 5095 25226
rect 3873 25124 3907 25158
rect 3873 25056 3907 25090
rect 3873 24988 3907 25022
rect 3873 24920 3907 24954
rect 3873 24852 3907 24886
rect 5061 25124 5095 25158
rect 5061 25056 5095 25090
rect 5061 24988 5095 25022
rect 5061 24920 5095 24954
rect 5061 24852 5095 24886
rect 3991 24750 4025 24784
rect 4059 24750 4093 24784
rect 4127 24750 4161 24784
rect 4195 24750 4229 24784
rect 4263 24750 4297 24784
rect 4331 24750 4365 24784
rect 4399 24750 4433 24784
rect 4467 24750 4501 24784
rect 4535 24750 4569 24784
rect 4603 24750 4637 24784
rect 4671 24750 4705 24784
rect 4739 24750 4773 24784
rect 4807 24750 4841 24784
rect 4875 24750 4909 24784
rect 4943 24750 4977 24784
rect 317 24003 351 24037
rect 385 24003 419 24037
rect 453 24003 487 24037
rect 521 24003 555 24037
rect 589 24003 623 24037
rect 657 24003 691 24037
rect 725 24003 759 24037
rect 793 24003 827 24037
rect 861 24003 895 24037
rect 929 24003 963 24037
rect 997 24003 1031 24037
rect 1065 24003 1099 24037
rect 1133 24003 1167 24037
rect 1201 24003 1235 24037
rect 1269 24003 1303 24037
rect 199 23901 233 23935
rect 1387 23901 1421 23935
rect 199 23833 233 23867
rect 199 23765 233 23799
rect 199 23697 233 23731
rect 199 23629 233 23663
rect 199 23561 233 23595
rect 1387 23833 1421 23867
rect 1387 23765 1421 23799
rect 1387 23697 1421 23731
rect 1387 23629 1421 23663
rect 1387 23561 1421 23595
rect 317 23459 351 23493
rect 385 23459 419 23493
rect 453 23459 487 23493
rect 521 23459 555 23493
rect 589 23459 623 23493
rect 657 23459 691 23493
rect 725 23459 759 23493
rect 793 23459 827 23493
rect 861 23459 895 23493
rect 929 23459 963 23493
rect 997 23459 1031 23493
rect 1065 23459 1099 23493
rect 1133 23459 1167 23493
rect 1201 23459 1235 23493
rect 1269 23459 1303 23493
rect 2470 24007 2504 24041
rect 2538 24007 2572 24041
rect 2606 24007 2640 24041
rect 2674 24007 2708 24041
rect 2742 24007 2776 24041
rect 2810 24007 2844 24041
rect 2878 24007 2912 24041
rect 2946 24007 2980 24041
rect 3014 24007 3048 24041
rect 3082 24007 3116 24041
rect 3150 24007 3184 24041
rect 3218 24007 3252 24041
rect 3286 24007 3320 24041
rect 3354 24007 3388 24041
rect 3422 24007 3456 24041
rect 2352 23905 2386 23939
rect 3540 23905 3574 23939
rect 2352 23837 2386 23871
rect 2352 23769 2386 23803
rect 2352 23701 2386 23735
rect 2352 23633 2386 23667
rect 2352 23565 2386 23599
rect 3540 23837 3574 23871
rect 3540 23769 3574 23803
rect 3540 23701 3574 23735
rect 3540 23633 3574 23667
rect 3540 23565 3574 23599
rect 2470 23463 2504 23497
rect 2538 23463 2572 23497
rect 2606 23463 2640 23497
rect 2674 23463 2708 23497
rect 2742 23463 2776 23497
rect 2810 23463 2844 23497
rect 2878 23463 2912 23497
rect 2946 23463 2980 23497
rect 3014 23463 3048 23497
rect 3082 23463 3116 23497
rect 3150 23463 3184 23497
rect 3218 23463 3252 23497
rect 3286 23463 3320 23497
rect 3354 23463 3388 23497
rect 3422 23463 3456 23497
rect 3991 24007 4025 24041
rect 4059 24007 4093 24041
rect 4127 24007 4161 24041
rect 4195 24007 4229 24041
rect 4263 24007 4297 24041
rect 4331 24007 4365 24041
rect 4399 24007 4433 24041
rect 4467 24007 4501 24041
rect 4535 24007 4569 24041
rect 4603 24007 4637 24041
rect 4671 24007 4705 24041
rect 4739 24007 4773 24041
rect 4807 24007 4841 24041
rect 4875 24007 4909 24041
rect 4943 24007 4977 24041
rect 3873 23905 3907 23939
rect 5061 23905 5095 23939
rect 3873 23837 3907 23871
rect 3873 23769 3907 23803
rect 3873 23701 3907 23735
rect 3873 23633 3907 23667
rect 3873 23565 3907 23599
rect 5061 23837 5095 23871
rect 5061 23769 5095 23803
rect 5061 23701 5095 23735
rect 5061 23633 5095 23667
rect 5061 23565 5095 23599
rect 3991 23463 4025 23497
rect 4059 23463 4093 23497
rect 4127 23463 4161 23497
rect 4195 23463 4229 23497
rect 4263 23463 4297 23497
rect 4331 23463 4365 23497
rect 4399 23463 4433 23497
rect 4467 23463 4501 23497
rect 4535 23463 4569 23497
rect 4603 23463 4637 23497
rect 4671 23463 4705 23497
rect 4739 23463 4773 23497
rect 4807 23463 4841 23497
rect 4875 23463 4909 23497
rect 4943 23463 4977 23497
rect 317 22716 351 22750
rect 385 22716 419 22750
rect 453 22716 487 22750
rect 521 22716 555 22750
rect 589 22716 623 22750
rect 657 22716 691 22750
rect 725 22716 759 22750
rect 793 22716 827 22750
rect 861 22716 895 22750
rect 929 22716 963 22750
rect 997 22716 1031 22750
rect 1065 22716 1099 22750
rect 1133 22716 1167 22750
rect 1201 22716 1235 22750
rect 1269 22716 1303 22750
rect 199 22614 233 22648
rect 1387 22614 1421 22648
rect 199 22546 233 22580
rect 199 22478 233 22512
rect 199 22410 233 22444
rect 199 22342 233 22376
rect 199 22274 233 22308
rect 1387 22546 1421 22580
rect 1387 22478 1421 22512
rect 1387 22410 1421 22444
rect 1387 22342 1421 22376
rect 1387 22274 1421 22308
rect 317 22172 351 22206
rect 385 22172 419 22206
rect 453 22172 487 22206
rect 521 22172 555 22206
rect 589 22172 623 22206
rect 657 22172 691 22206
rect 725 22172 759 22206
rect 793 22172 827 22206
rect 861 22172 895 22206
rect 929 22172 963 22206
rect 997 22172 1031 22206
rect 1065 22172 1099 22206
rect 1133 22172 1167 22206
rect 1201 22172 1235 22206
rect 1269 22172 1303 22206
rect 2470 22720 2504 22754
rect 2538 22720 2572 22754
rect 2606 22720 2640 22754
rect 2674 22720 2708 22754
rect 2742 22720 2776 22754
rect 2810 22720 2844 22754
rect 2878 22720 2912 22754
rect 2946 22720 2980 22754
rect 3014 22720 3048 22754
rect 3082 22720 3116 22754
rect 3150 22720 3184 22754
rect 3218 22720 3252 22754
rect 3286 22720 3320 22754
rect 3354 22720 3388 22754
rect 3422 22720 3456 22754
rect 2352 22618 2386 22652
rect 3540 22618 3574 22652
rect 2352 22550 2386 22584
rect 2352 22482 2386 22516
rect 2352 22414 2386 22448
rect 2352 22346 2386 22380
rect 2352 22278 2386 22312
rect 3540 22550 3574 22584
rect 3540 22482 3574 22516
rect 3540 22414 3574 22448
rect 3540 22346 3574 22380
rect 3540 22278 3574 22312
rect 2470 22176 2504 22210
rect 2538 22176 2572 22210
rect 2606 22176 2640 22210
rect 2674 22176 2708 22210
rect 2742 22176 2776 22210
rect 2810 22176 2844 22210
rect 2878 22176 2912 22210
rect 2946 22176 2980 22210
rect 3014 22176 3048 22210
rect 3082 22176 3116 22210
rect 3150 22176 3184 22210
rect 3218 22176 3252 22210
rect 3286 22176 3320 22210
rect 3354 22176 3388 22210
rect 3422 22176 3456 22210
rect 3991 22720 4025 22754
rect 4059 22720 4093 22754
rect 4127 22720 4161 22754
rect 4195 22720 4229 22754
rect 4263 22720 4297 22754
rect 4331 22720 4365 22754
rect 4399 22720 4433 22754
rect 4467 22720 4501 22754
rect 4535 22720 4569 22754
rect 4603 22720 4637 22754
rect 4671 22720 4705 22754
rect 4739 22720 4773 22754
rect 4807 22720 4841 22754
rect 4875 22720 4909 22754
rect 4943 22720 4977 22754
rect 3873 22618 3907 22652
rect 5061 22618 5095 22652
rect 3873 22550 3907 22584
rect 3873 22482 3907 22516
rect 3873 22414 3907 22448
rect 3873 22346 3907 22380
rect 3873 22278 3907 22312
rect 5061 22550 5095 22584
rect 5061 22482 5095 22516
rect 5061 22414 5095 22448
rect 5061 22346 5095 22380
rect 5061 22278 5095 22312
rect 3991 22176 4025 22210
rect 4059 22176 4093 22210
rect 4127 22176 4161 22210
rect 4195 22176 4229 22210
rect 4263 22176 4297 22210
rect 4331 22176 4365 22210
rect 4399 22176 4433 22210
rect 4467 22176 4501 22210
rect 4535 22176 4569 22210
rect 4603 22176 4637 22210
rect 4671 22176 4705 22210
rect 4739 22176 4773 22210
rect 4807 22176 4841 22210
rect 4875 22176 4909 22210
rect 4943 22176 4977 22210
rect 317 21429 351 21463
rect 385 21429 419 21463
rect 453 21429 487 21463
rect 521 21429 555 21463
rect 589 21429 623 21463
rect 657 21429 691 21463
rect 725 21429 759 21463
rect 793 21429 827 21463
rect 861 21429 895 21463
rect 929 21429 963 21463
rect 997 21429 1031 21463
rect 1065 21429 1099 21463
rect 1133 21429 1167 21463
rect 1201 21429 1235 21463
rect 1269 21429 1303 21463
rect 199 21327 233 21361
rect 1387 21327 1421 21361
rect 199 21259 233 21293
rect 199 21191 233 21225
rect 199 21123 233 21157
rect 199 21055 233 21089
rect 199 20987 233 21021
rect 1387 21259 1421 21293
rect 1387 21191 1421 21225
rect 1387 21123 1421 21157
rect 1387 21055 1421 21089
rect 1387 20987 1421 21021
rect 317 20885 351 20919
rect 385 20885 419 20919
rect 453 20885 487 20919
rect 521 20885 555 20919
rect 589 20885 623 20919
rect 657 20885 691 20919
rect 725 20885 759 20919
rect 793 20885 827 20919
rect 861 20885 895 20919
rect 929 20885 963 20919
rect 997 20885 1031 20919
rect 1065 20885 1099 20919
rect 1133 20885 1167 20919
rect 1201 20885 1235 20919
rect 1269 20885 1303 20919
rect 2470 21433 2504 21467
rect 2538 21433 2572 21467
rect 2606 21433 2640 21467
rect 2674 21433 2708 21467
rect 2742 21433 2776 21467
rect 2810 21433 2844 21467
rect 2878 21433 2912 21467
rect 2946 21433 2980 21467
rect 3014 21433 3048 21467
rect 3082 21433 3116 21467
rect 3150 21433 3184 21467
rect 3218 21433 3252 21467
rect 3286 21433 3320 21467
rect 3354 21433 3388 21467
rect 3422 21433 3456 21467
rect 2352 21331 2386 21365
rect 3540 21331 3574 21365
rect 2352 21263 2386 21297
rect 2352 21195 2386 21229
rect 2352 21127 2386 21161
rect 2352 21059 2386 21093
rect 2352 20991 2386 21025
rect 3540 21263 3574 21297
rect 3540 21195 3574 21229
rect 3540 21127 3574 21161
rect 3540 21059 3574 21093
rect 3540 20991 3574 21025
rect 2470 20889 2504 20923
rect 2538 20889 2572 20923
rect 2606 20889 2640 20923
rect 2674 20889 2708 20923
rect 2742 20889 2776 20923
rect 2810 20889 2844 20923
rect 2878 20889 2912 20923
rect 2946 20889 2980 20923
rect 3014 20889 3048 20923
rect 3082 20889 3116 20923
rect 3150 20889 3184 20923
rect 3218 20889 3252 20923
rect 3286 20889 3320 20923
rect 3354 20889 3388 20923
rect 3422 20889 3456 20923
rect 3991 21433 4025 21467
rect 4059 21433 4093 21467
rect 4127 21433 4161 21467
rect 4195 21433 4229 21467
rect 4263 21433 4297 21467
rect 4331 21433 4365 21467
rect 4399 21433 4433 21467
rect 4467 21433 4501 21467
rect 4535 21433 4569 21467
rect 4603 21433 4637 21467
rect 4671 21433 4705 21467
rect 4739 21433 4773 21467
rect 4807 21433 4841 21467
rect 4875 21433 4909 21467
rect 4943 21433 4977 21467
rect 3873 21331 3907 21365
rect 5061 21331 5095 21365
rect 3873 21263 3907 21297
rect 3873 21195 3907 21229
rect 3873 21127 3907 21161
rect 3873 21059 3907 21093
rect 3873 20991 3907 21025
rect 5061 21263 5095 21297
rect 5061 21195 5095 21229
rect 5061 21127 5095 21161
rect 5061 21059 5095 21093
rect 5061 20991 5095 21025
rect 3991 20889 4025 20923
rect 4059 20889 4093 20923
rect 4127 20889 4161 20923
rect 4195 20889 4229 20923
rect 4263 20889 4297 20923
rect 4331 20889 4365 20923
rect 4399 20889 4433 20923
rect 4467 20889 4501 20923
rect 4535 20889 4569 20923
rect 4603 20889 4637 20923
rect 4671 20889 4705 20923
rect 4739 20889 4773 20923
rect 4807 20889 4841 20923
rect 4875 20889 4909 20923
rect 4943 20889 4977 20923
rect 317 20142 351 20176
rect 385 20142 419 20176
rect 453 20142 487 20176
rect 521 20142 555 20176
rect 589 20142 623 20176
rect 657 20142 691 20176
rect 725 20142 759 20176
rect 793 20142 827 20176
rect 861 20142 895 20176
rect 929 20142 963 20176
rect 997 20142 1031 20176
rect 1065 20142 1099 20176
rect 1133 20142 1167 20176
rect 1201 20142 1235 20176
rect 1269 20142 1303 20176
rect 199 20040 233 20074
rect 1387 20040 1421 20074
rect 199 19972 233 20006
rect 199 19904 233 19938
rect 199 19836 233 19870
rect 199 19768 233 19802
rect 199 19700 233 19734
rect 1387 19972 1421 20006
rect 1387 19904 1421 19938
rect 1387 19836 1421 19870
rect 1387 19768 1421 19802
rect 1387 19700 1421 19734
rect 317 19598 351 19632
rect 385 19598 419 19632
rect 453 19598 487 19632
rect 521 19598 555 19632
rect 589 19598 623 19632
rect 657 19598 691 19632
rect 725 19598 759 19632
rect 793 19598 827 19632
rect 861 19598 895 19632
rect 929 19598 963 19632
rect 997 19598 1031 19632
rect 1065 19598 1099 19632
rect 1133 19598 1167 19632
rect 1201 19598 1235 19632
rect 1269 19598 1303 19632
rect 2470 20146 2504 20180
rect 2538 20146 2572 20180
rect 2606 20146 2640 20180
rect 2674 20146 2708 20180
rect 2742 20146 2776 20180
rect 2810 20146 2844 20180
rect 2878 20146 2912 20180
rect 2946 20146 2980 20180
rect 3014 20146 3048 20180
rect 3082 20146 3116 20180
rect 3150 20146 3184 20180
rect 3218 20146 3252 20180
rect 3286 20146 3320 20180
rect 3354 20146 3388 20180
rect 3422 20146 3456 20180
rect 2352 20044 2386 20078
rect 3540 20044 3574 20078
rect 2352 19976 2386 20010
rect 2352 19908 2386 19942
rect 2352 19840 2386 19874
rect 2352 19772 2386 19806
rect 2352 19704 2386 19738
rect 3540 19976 3574 20010
rect 3540 19908 3574 19942
rect 3540 19840 3574 19874
rect 3540 19772 3574 19806
rect 3540 19704 3574 19738
rect 2470 19602 2504 19636
rect 2538 19602 2572 19636
rect 2606 19602 2640 19636
rect 2674 19602 2708 19636
rect 2742 19602 2776 19636
rect 2810 19602 2844 19636
rect 2878 19602 2912 19636
rect 2946 19602 2980 19636
rect 3014 19602 3048 19636
rect 3082 19602 3116 19636
rect 3150 19602 3184 19636
rect 3218 19602 3252 19636
rect 3286 19602 3320 19636
rect 3354 19602 3388 19636
rect 3422 19602 3456 19636
rect 3991 20146 4025 20180
rect 4059 20146 4093 20180
rect 4127 20146 4161 20180
rect 4195 20146 4229 20180
rect 4263 20146 4297 20180
rect 4331 20146 4365 20180
rect 4399 20146 4433 20180
rect 4467 20146 4501 20180
rect 4535 20146 4569 20180
rect 4603 20146 4637 20180
rect 4671 20146 4705 20180
rect 4739 20146 4773 20180
rect 4807 20146 4841 20180
rect 4875 20146 4909 20180
rect 4943 20146 4977 20180
rect 3873 20044 3907 20078
rect 5061 20044 5095 20078
rect 3873 19976 3907 20010
rect 3873 19908 3907 19942
rect 3873 19840 3907 19874
rect 3873 19772 3907 19806
rect 3873 19704 3907 19738
rect 5061 19976 5095 20010
rect 5061 19908 5095 19942
rect 5061 19840 5095 19874
rect 5061 19772 5095 19806
rect 5061 19704 5095 19738
rect 3991 19602 4025 19636
rect 4059 19602 4093 19636
rect 4127 19602 4161 19636
rect 4195 19602 4229 19636
rect 4263 19602 4297 19636
rect 4331 19602 4365 19636
rect 4399 19602 4433 19636
rect 4467 19602 4501 19636
rect 4535 19602 4569 19636
rect 4603 19602 4637 19636
rect 4671 19602 4705 19636
rect 4739 19602 4773 19636
rect 4807 19602 4841 19636
rect 4875 19602 4909 19636
rect 4943 19602 4977 19636
rect 317 18855 351 18889
rect 385 18855 419 18889
rect 453 18855 487 18889
rect 521 18855 555 18889
rect 589 18855 623 18889
rect 657 18855 691 18889
rect 725 18855 759 18889
rect 793 18855 827 18889
rect 861 18855 895 18889
rect 929 18855 963 18889
rect 997 18855 1031 18889
rect 1065 18855 1099 18889
rect 1133 18855 1167 18889
rect 1201 18855 1235 18889
rect 1269 18855 1303 18889
rect 199 18753 233 18787
rect 1387 18753 1421 18787
rect 199 18685 233 18719
rect 199 18617 233 18651
rect 199 18549 233 18583
rect 199 18481 233 18515
rect 199 18413 233 18447
rect 1387 18685 1421 18719
rect 1387 18617 1421 18651
rect 1387 18549 1421 18583
rect 1387 18481 1421 18515
rect 1387 18413 1421 18447
rect 317 18311 351 18345
rect 385 18311 419 18345
rect 453 18311 487 18345
rect 521 18311 555 18345
rect 589 18311 623 18345
rect 657 18311 691 18345
rect 725 18311 759 18345
rect 793 18311 827 18345
rect 861 18311 895 18345
rect 929 18311 963 18345
rect 997 18311 1031 18345
rect 1065 18311 1099 18345
rect 1133 18311 1167 18345
rect 1201 18311 1235 18345
rect 1269 18311 1303 18345
rect 2470 18859 2504 18893
rect 2538 18859 2572 18893
rect 2606 18859 2640 18893
rect 2674 18859 2708 18893
rect 2742 18859 2776 18893
rect 2810 18859 2844 18893
rect 2878 18859 2912 18893
rect 2946 18859 2980 18893
rect 3014 18859 3048 18893
rect 3082 18859 3116 18893
rect 3150 18859 3184 18893
rect 3218 18859 3252 18893
rect 3286 18859 3320 18893
rect 3354 18859 3388 18893
rect 3422 18859 3456 18893
rect 2352 18757 2386 18791
rect 3540 18757 3574 18791
rect 2352 18689 2386 18723
rect 2352 18621 2386 18655
rect 2352 18553 2386 18587
rect 2352 18485 2386 18519
rect 2352 18417 2386 18451
rect 3540 18689 3574 18723
rect 3540 18621 3574 18655
rect 3540 18553 3574 18587
rect 3540 18485 3574 18519
rect 3540 18417 3574 18451
rect 2470 18315 2504 18349
rect 2538 18315 2572 18349
rect 2606 18315 2640 18349
rect 2674 18315 2708 18349
rect 2742 18315 2776 18349
rect 2810 18315 2844 18349
rect 2878 18315 2912 18349
rect 2946 18315 2980 18349
rect 3014 18315 3048 18349
rect 3082 18315 3116 18349
rect 3150 18315 3184 18349
rect 3218 18315 3252 18349
rect 3286 18315 3320 18349
rect 3354 18315 3388 18349
rect 3422 18315 3456 18349
rect 3991 18859 4025 18893
rect 4059 18859 4093 18893
rect 4127 18859 4161 18893
rect 4195 18859 4229 18893
rect 4263 18859 4297 18893
rect 4331 18859 4365 18893
rect 4399 18859 4433 18893
rect 4467 18859 4501 18893
rect 4535 18859 4569 18893
rect 4603 18859 4637 18893
rect 4671 18859 4705 18893
rect 4739 18859 4773 18893
rect 4807 18859 4841 18893
rect 4875 18859 4909 18893
rect 4943 18859 4977 18893
rect 3873 18757 3907 18791
rect 5061 18757 5095 18791
rect 3873 18689 3907 18723
rect 3873 18621 3907 18655
rect 3873 18553 3907 18587
rect 3873 18485 3907 18519
rect 3873 18417 3907 18451
rect 5061 18689 5095 18723
rect 5061 18621 5095 18655
rect 5061 18553 5095 18587
rect 5061 18485 5095 18519
rect 5061 18417 5095 18451
rect 3991 18315 4025 18349
rect 4059 18315 4093 18349
rect 4127 18315 4161 18349
rect 4195 18315 4229 18349
rect 4263 18315 4297 18349
rect 4331 18315 4365 18349
rect 4399 18315 4433 18349
rect 4467 18315 4501 18349
rect 4535 18315 4569 18349
rect 4603 18315 4637 18349
rect 4671 18315 4705 18349
rect 4739 18315 4773 18349
rect 4807 18315 4841 18349
rect 4875 18315 4909 18349
rect 4943 18315 4977 18349
rect 317 17568 351 17602
rect 385 17568 419 17602
rect 453 17568 487 17602
rect 521 17568 555 17602
rect 589 17568 623 17602
rect 657 17568 691 17602
rect 725 17568 759 17602
rect 793 17568 827 17602
rect 861 17568 895 17602
rect 929 17568 963 17602
rect 997 17568 1031 17602
rect 1065 17568 1099 17602
rect 1133 17568 1167 17602
rect 1201 17568 1235 17602
rect 1269 17568 1303 17602
rect 199 17466 233 17500
rect 1387 17466 1421 17500
rect 199 17398 233 17432
rect 199 17330 233 17364
rect 199 17262 233 17296
rect 199 17194 233 17228
rect 199 17126 233 17160
rect 1387 17398 1421 17432
rect 1387 17330 1421 17364
rect 1387 17262 1421 17296
rect 1387 17194 1421 17228
rect 1387 17126 1421 17160
rect 317 17024 351 17058
rect 385 17024 419 17058
rect 453 17024 487 17058
rect 521 17024 555 17058
rect 589 17024 623 17058
rect 657 17024 691 17058
rect 725 17024 759 17058
rect 793 17024 827 17058
rect 861 17024 895 17058
rect 929 17024 963 17058
rect 997 17024 1031 17058
rect 1065 17024 1099 17058
rect 1133 17024 1167 17058
rect 1201 17024 1235 17058
rect 1269 17024 1303 17058
rect 2470 17572 2504 17606
rect 2538 17572 2572 17606
rect 2606 17572 2640 17606
rect 2674 17572 2708 17606
rect 2742 17572 2776 17606
rect 2810 17572 2844 17606
rect 2878 17572 2912 17606
rect 2946 17572 2980 17606
rect 3014 17572 3048 17606
rect 3082 17572 3116 17606
rect 3150 17572 3184 17606
rect 3218 17572 3252 17606
rect 3286 17572 3320 17606
rect 3354 17572 3388 17606
rect 3422 17572 3456 17606
rect 2352 17470 2386 17504
rect 3540 17470 3574 17504
rect 2352 17402 2386 17436
rect 2352 17334 2386 17368
rect 2352 17266 2386 17300
rect 2352 17198 2386 17232
rect 2352 17130 2386 17164
rect 3540 17402 3574 17436
rect 3540 17334 3574 17368
rect 3540 17266 3574 17300
rect 3540 17198 3574 17232
rect 3540 17130 3574 17164
rect 2470 17028 2504 17062
rect 2538 17028 2572 17062
rect 2606 17028 2640 17062
rect 2674 17028 2708 17062
rect 2742 17028 2776 17062
rect 2810 17028 2844 17062
rect 2878 17028 2912 17062
rect 2946 17028 2980 17062
rect 3014 17028 3048 17062
rect 3082 17028 3116 17062
rect 3150 17028 3184 17062
rect 3218 17028 3252 17062
rect 3286 17028 3320 17062
rect 3354 17028 3388 17062
rect 3422 17028 3456 17062
rect 3991 17572 4025 17606
rect 4059 17572 4093 17606
rect 4127 17572 4161 17606
rect 4195 17572 4229 17606
rect 4263 17572 4297 17606
rect 4331 17572 4365 17606
rect 4399 17572 4433 17606
rect 4467 17572 4501 17606
rect 4535 17572 4569 17606
rect 4603 17572 4637 17606
rect 4671 17572 4705 17606
rect 4739 17572 4773 17606
rect 4807 17572 4841 17606
rect 4875 17572 4909 17606
rect 4943 17572 4977 17606
rect 3873 17470 3907 17504
rect 5061 17470 5095 17504
rect 3873 17402 3907 17436
rect 3873 17334 3907 17368
rect 3873 17266 3907 17300
rect 3873 17198 3907 17232
rect 3873 17130 3907 17164
rect 5061 17402 5095 17436
rect 5061 17334 5095 17368
rect 5061 17266 5095 17300
rect 5061 17198 5095 17232
rect 5061 17130 5095 17164
rect 3991 17028 4025 17062
rect 4059 17028 4093 17062
rect 4127 17028 4161 17062
rect 4195 17028 4229 17062
rect 4263 17028 4297 17062
rect 4331 17028 4365 17062
rect 4399 17028 4433 17062
rect 4467 17028 4501 17062
rect 4535 17028 4569 17062
rect 4603 17028 4637 17062
rect 4671 17028 4705 17062
rect 4739 17028 4773 17062
rect 4807 17028 4841 17062
rect 4875 17028 4909 17062
rect 4943 17028 4977 17062
rect 317 16281 351 16315
rect 385 16281 419 16315
rect 453 16281 487 16315
rect 521 16281 555 16315
rect 589 16281 623 16315
rect 657 16281 691 16315
rect 725 16281 759 16315
rect 793 16281 827 16315
rect 861 16281 895 16315
rect 929 16281 963 16315
rect 997 16281 1031 16315
rect 1065 16281 1099 16315
rect 1133 16281 1167 16315
rect 1201 16281 1235 16315
rect 1269 16281 1303 16315
rect 199 16179 233 16213
rect 1387 16179 1421 16213
rect 199 16111 233 16145
rect 199 16043 233 16077
rect 199 15975 233 16009
rect 199 15907 233 15941
rect 199 15839 233 15873
rect 1387 16111 1421 16145
rect 1387 16043 1421 16077
rect 1387 15975 1421 16009
rect 1387 15907 1421 15941
rect 1387 15839 1421 15873
rect 317 15737 351 15771
rect 385 15737 419 15771
rect 453 15737 487 15771
rect 521 15737 555 15771
rect 589 15737 623 15771
rect 657 15737 691 15771
rect 725 15737 759 15771
rect 793 15737 827 15771
rect 861 15737 895 15771
rect 929 15737 963 15771
rect 997 15737 1031 15771
rect 1065 15737 1099 15771
rect 1133 15737 1167 15771
rect 1201 15737 1235 15771
rect 1269 15737 1303 15771
rect 2470 16285 2504 16319
rect 2538 16285 2572 16319
rect 2606 16285 2640 16319
rect 2674 16285 2708 16319
rect 2742 16285 2776 16319
rect 2810 16285 2844 16319
rect 2878 16285 2912 16319
rect 2946 16285 2980 16319
rect 3014 16285 3048 16319
rect 3082 16285 3116 16319
rect 3150 16285 3184 16319
rect 3218 16285 3252 16319
rect 3286 16285 3320 16319
rect 3354 16285 3388 16319
rect 3422 16285 3456 16319
rect 2352 16183 2386 16217
rect 3540 16183 3574 16217
rect 2352 16115 2386 16149
rect 2352 16047 2386 16081
rect 2352 15979 2386 16013
rect 2352 15911 2386 15945
rect 2352 15843 2386 15877
rect 3540 16115 3574 16149
rect 3540 16047 3574 16081
rect 3540 15979 3574 16013
rect 3540 15911 3574 15945
rect 3540 15843 3574 15877
rect 2470 15741 2504 15775
rect 2538 15741 2572 15775
rect 2606 15741 2640 15775
rect 2674 15741 2708 15775
rect 2742 15741 2776 15775
rect 2810 15741 2844 15775
rect 2878 15741 2912 15775
rect 2946 15741 2980 15775
rect 3014 15741 3048 15775
rect 3082 15741 3116 15775
rect 3150 15741 3184 15775
rect 3218 15741 3252 15775
rect 3286 15741 3320 15775
rect 3354 15741 3388 15775
rect 3422 15741 3456 15775
rect 3991 16285 4025 16319
rect 4059 16285 4093 16319
rect 4127 16285 4161 16319
rect 4195 16285 4229 16319
rect 4263 16285 4297 16319
rect 4331 16285 4365 16319
rect 4399 16285 4433 16319
rect 4467 16285 4501 16319
rect 4535 16285 4569 16319
rect 4603 16285 4637 16319
rect 4671 16285 4705 16319
rect 4739 16285 4773 16319
rect 4807 16285 4841 16319
rect 4875 16285 4909 16319
rect 4943 16285 4977 16319
rect 3873 16183 3907 16217
rect 5061 16183 5095 16217
rect 3873 16115 3907 16149
rect 3873 16047 3907 16081
rect 3873 15979 3907 16013
rect 3873 15911 3907 15945
rect 3873 15843 3907 15877
rect 5061 16115 5095 16149
rect 5061 16047 5095 16081
rect 5061 15979 5095 16013
rect 5061 15911 5095 15945
rect 5061 15843 5095 15877
rect 3991 15741 4025 15775
rect 4059 15741 4093 15775
rect 4127 15741 4161 15775
rect 4195 15741 4229 15775
rect 4263 15741 4297 15775
rect 4331 15741 4365 15775
rect 4399 15741 4433 15775
rect 4467 15741 4501 15775
rect 4535 15741 4569 15775
rect 4603 15741 4637 15775
rect 4671 15741 4705 15775
rect 4739 15741 4773 15775
rect 4807 15741 4841 15775
rect 4875 15741 4909 15775
rect 4943 15741 4977 15775
rect 317 14994 351 15028
rect 385 14994 419 15028
rect 453 14994 487 15028
rect 521 14994 555 15028
rect 589 14994 623 15028
rect 657 14994 691 15028
rect 725 14994 759 15028
rect 793 14994 827 15028
rect 861 14994 895 15028
rect 929 14994 963 15028
rect 997 14994 1031 15028
rect 1065 14994 1099 15028
rect 1133 14994 1167 15028
rect 1201 14994 1235 15028
rect 1269 14994 1303 15028
rect 199 14892 233 14926
rect 1387 14892 1421 14926
rect 199 14824 233 14858
rect 199 14756 233 14790
rect 199 14688 233 14722
rect 199 14620 233 14654
rect 199 14552 233 14586
rect 1387 14824 1421 14858
rect 1387 14756 1421 14790
rect 1387 14688 1421 14722
rect 1387 14620 1421 14654
rect 1387 14552 1421 14586
rect 317 14450 351 14484
rect 385 14450 419 14484
rect 453 14450 487 14484
rect 521 14450 555 14484
rect 589 14450 623 14484
rect 657 14450 691 14484
rect 725 14450 759 14484
rect 793 14450 827 14484
rect 861 14450 895 14484
rect 929 14450 963 14484
rect 997 14450 1031 14484
rect 1065 14450 1099 14484
rect 1133 14450 1167 14484
rect 1201 14450 1235 14484
rect 1269 14450 1303 14484
rect 2470 14998 2504 15032
rect 2538 14998 2572 15032
rect 2606 14998 2640 15032
rect 2674 14998 2708 15032
rect 2742 14998 2776 15032
rect 2810 14998 2844 15032
rect 2878 14998 2912 15032
rect 2946 14998 2980 15032
rect 3014 14998 3048 15032
rect 3082 14998 3116 15032
rect 3150 14998 3184 15032
rect 3218 14998 3252 15032
rect 3286 14998 3320 15032
rect 3354 14998 3388 15032
rect 3422 14998 3456 15032
rect 2352 14896 2386 14930
rect 3540 14896 3574 14930
rect 2352 14828 2386 14862
rect 2352 14760 2386 14794
rect 2352 14692 2386 14726
rect 2352 14624 2386 14658
rect 2352 14556 2386 14590
rect 3540 14828 3574 14862
rect 3540 14760 3574 14794
rect 3540 14692 3574 14726
rect 3540 14624 3574 14658
rect 3540 14556 3574 14590
rect 2470 14454 2504 14488
rect 2538 14454 2572 14488
rect 2606 14454 2640 14488
rect 2674 14454 2708 14488
rect 2742 14454 2776 14488
rect 2810 14454 2844 14488
rect 2878 14454 2912 14488
rect 2946 14454 2980 14488
rect 3014 14454 3048 14488
rect 3082 14454 3116 14488
rect 3150 14454 3184 14488
rect 3218 14454 3252 14488
rect 3286 14454 3320 14488
rect 3354 14454 3388 14488
rect 3422 14454 3456 14488
rect 3991 14998 4025 15032
rect 4059 14998 4093 15032
rect 4127 14998 4161 15032
rect 4195 14998 4229 15032
rect 4263 14998 4297 15032
rect 4331 14998 4365 15032
rect 4399 14998 4433 15032
rect 4467 14998 4501 15032
rect 4535 14998 4569 15032
rect 4603 14998 4637 15032
rect 4671 14998 4705 15032
rect 4739 14998 4773 15032
rect 4807 14998 4841 15032
rect 4875 14998 4909 15032
rect 4943 14998 4977 15032
rect 3873 14896 3907 14930
rect 5061 14896 5095 14930
rect 3873 14828 3907 14862
rect 3873 14760 3907 14794
rect 3873 14692 3907 14726
rect 3873 14624 3907 14658
rect 3873 14556 3907 14590
rect 5061 14828 5095 14862
rect 5061 14760 5095 14794
rect 5061 14692 5095 14726
rect 5061 14624 5095 14658
rect 5061 14556 5095 14590
rect 3991 14454 4025 14488
rect 4059 14454 4093 14488
rect 4127 14454 4161 14488
rect 4195 14454 4229 14488
rect 4263 14454 4297 14488
rect 4331 14454 4365 14488
rect 4399 14454 4433 14488
rect 4467 14454 4501 14488
rect 4535 14454 4569 14488
rect 4603 14454 4637 14488
rect 4671 14454 4705 14488
rect 4739 14454 4773 14488
rect 4807 14454 4841 14488
rect 4875 14454 4909 14488
rect 4943 14454 4977 14488
rect 317 13707 351 13741
rect 385 13707 419 13741
rect 453 13707 487 13741
rect 521 13707 555 13741
rect 589 13707 623 13741
rect 657 13707 691 13741
rect 725 13707 759 13741
rect 793 13707 827 13741
rect 861 13707 895 13741
rect 929 13707 963 13741
rect 997 13707 1031 13741
rect 1065 13707 1099 13741
rect 1133 13707 1167 13741
rect 1201 13707 1235 13741
rect 1269 13707 1303 13741
rect 199 13605 233 13639
rect 1387 13605 1421 13639
rect 199 13537 233 13571
rect 199 13469 233 13503
rect 199 13401 233 13435
rect 199 13333 233 13367
rect 199 13265 233 13299
rect 1387 13537 1421 13571
rect 1387 13469 1421 13503
rect 1387 13401 1421 13435
rect 1387 13333 1421 13367
rect 1387 13265 1421 13299
rect 317 13163 351 13197
rect 385 13163 419 13197
rect 453 13163 487 13197
rect 521 13163 555 13197
rect 589 13163 623 13197
rect 657 13163 691 13197
rect 725 13163 759 13197
rect 793 13163 827 13197
rect 861 13163 895 13197
rect 929 13163 963 13197
rect 997 13163 1031 13197
rect 1065 13163 1099 13197
rect 1133 13163 1167 13197
rect 1201 13163 1235 13197
rect 1269 13163 1303 13197
rect 2470 13711 2504 13745
rect 2538 13711 2572 13745
rect 2606 13711 2640 13745
rect 2674 13711 2708 13745
rect 2742 13711 2776 13745
rect 2810 13711 2844 13745
rect 2878 13711 2912 13745
rect 2946 13711 2980 13745
rect 3014 13711 3048 13745
rect 3082 13711 3116 13745
rect 3150 13711 3184 13745
rect 3218 13711 3252 13745
rect 3286 13711 3320 13745
rect 3354 13711 3388 13745
rect 3422 13711 3456 13745
rect 2352 13609 2386 13643
rect 3540 13609 3574 13643
rect 2352 13541 2386 13575
rect 2352 13473 2386 13507
rect 2352 13405 2386 13439
rect 2352 13337 2386 13371
rect 2352 13269 2386 13303
rect 3540 13541 3574 13575
rect 3540 13473 3574 13507
rect 3540 13405 3574 13439
rect 3540 13337 3574 13371
rect 3540 13269 3574 13303
rect 2470 13167 2504 13201
rect 2538 13167 2572 13201
rect 2606 13167 2640 13201
rect 2674 13167 2708 13201
rect 2742 13167 2776 13201
rect 2810 13167 2844 13201
rect 2878 13167 2912 13201
rect 2946 13167 2980 13201
rect 3014 13167 3048 13201
rect 3082 13167 3116 13201
rect 3150 13167 3184 13201
rect 3218 13167 3252 13201
rect 3286 13167 3320 13201
rect 3354 13167 3388 13201
rect 3422 13167 3456 13201
rect 3991 13711 4025 13745
rect 4059 13711 4093 13745
rect 4127 13711 4161 13745
rect 4195 13711 4229 13745
rect 4263 13711 4297 13745
rect 4331 13711 4365 13745
rect 4399 13711 4433 13745
rect 4467 13711 4501 13745
rect 4535 13711 4569 13745
rect 4603 13711 4637 13745
rect 4671 13711 4705 13745
rect 4739 13711 4773 13745
rect 4807 13711 4841 13745
rect 4875 13711 4909 13745
rect 4943 13711 4977 13745
rect 3873 13609 3907 13643
rect 5061 13609 5095 13643
rect 3873 13541 3907 13575
rect 3873 13473 3907 13507
rect 3873 13405 3907 13439
rect 3873 13337 3907 13371
rect 3873 13269 3907 13303
rect 5061 13541 5095 13575
rect 5061 13473 5095 13507
rect 5061 13405 5095 13439
rect 5061 13337 5095 13371
rect 5061 13269 5095 13303
rect 3991 13167 4025 13201
rect 4059 13167 4093 13201
rect 4127 13167 4161 13201
rect 4195 13167 4229 13201
rect 4263 13167 4297 13201
rect 4331 13167 4365 13201
rect 4399 13167 4433 13201
rect 4467 13167 4501 13201
rect 4535 13167 4569 13201
rect 4603 13167 4637 13201
rect 4671 13167 4705 13201
rect 4739 13167 4773 13201
rect 4807 13167 4841 13201
rect 4875 13167 4909 13201
rect 4943 13167 4977 13201
rect 317 12420 351 12454
rect 385 12420 419 12454
rect 453 12420 487 12454
rect 521 12420 555 12454
rect 589 12420 623 12454
rect 657 12420 691 12454
rect 725 12420 759 12454
rect 793 12420 827 12454
rect 861 12420 895 12454
rect 929 12420 963 12454
rect 997 12420 1031 12454
rect 1065 12420 1099 12454
rect 1133 12420 1167 12454
rect 1201 12420 1235 12454
rect 1269 12420 1303 12454
rect 199 12318 233 12352
rect 1387 12318 1421 12352
rect 199 12250 233 12284
rect 199 12182 233 12216
rect 199 12114 233 12148
rect 199 12046 233 12080
rect 199 11978 233 12012
rect 1387 12250 1421 12284
rect 1387 12182 1421 12216
rect 1387 12114 1421 12148
rect 1387 12046 1421 12080
rect 1387 11978 1421 12012
rect 317 11876 351 11910
rect 385 11876 419 11910
rect 453 11876 487 11910
rect 521 11876 555 11910
rect 589 11876 623 11910
rect 657 11876 691 11910
rect 725 11876 759 11910
rect 793 11876 827 11910
rect 861 11876 895 11910
rect 929 11876 963 11910
rect 997 11876 1031 11910
rect 1065 11876 1099 11910
rect 1133 11876 1167 11910
rect 1201 11876 1235 11910
rect 1269 11876 1303 11910
rect 2470 12424 2504 12458
rect 2538 12424 2572 12458
rect 2606 12424 2640 12458
rect 2674 12424 2708 12458
rect 2742 12424 2776 12458
rect 2810 12424 2844 12458
rect 2878 12424 2912 12458
rect 2946 12424 2980 12458
rect 3014 12424 3048 12458
rect 3082 12424 3116 12458
rect 3150 12424 3184 12458
rect 3218 12424 3252 12458
rect 3286 12424 3320 12458
rect 3354 12424 3388 12458
rect 3422 12424 3456 12458
rect 2352 12322 2386 12356
rect 3540 12322 3574 12356
rect 2352 12254 2386 12288
rect 2352 12186 2386 12220
rect 2352 12118 2386 12152
rect 2352 12050 2386 12084
rect 2352 11982 2386 12016
rect 3540 12254 3574 12288
rect 3540 12186 3574 12220
rect 3540 12118 3574 12152
rect 3540 12050 3574 12084
rect 3540 11982 3574 12016
rect 2470 11880 2504 11914
rect 2538 11880 2572 11914
rect 2606 11880 2640 11914
rect 2674 11880 2708 11914
rect 2742 11880 2776 11914
rect 2810 11880 2844 11914
rect 2878 11880 2912 11914
rect 2946 11880 2980 11914
rect 3014 11880 3048 11914
rect 3082 11880 3116 11914
rect 3150 11880 3184 11914
rect 3218 11880 3252 11914
rect 3286 11880 3320 11914
rect 3354 11880 3388 11914
rect 3422 11880 3456 11914
rect 3991 12424 4025 12458
rect 4059 12424 4093 12458
rect 4127 12424 4161 12458
rect 4195 12424 4229 12458
rect 4263 12424 4297 12458
rect 4331 12424 4365 12458
rect 4399 12424 4433 12458
rect 4467 12424 4501 12458
rect 4535 12424 4569 12458
rect 4603 12424 4637 12458
rect 4671 12424 4705 12458
rect 4739 12424 4773 12458
rect 4807 12424 4841 12458
rect 4875 12424 4909 12458
rect 4943 12424 4977 12458
rect 3873 12322 3907 12356
rect 5061 12322 5095 12356
rect 3873 12254 3907 12288
rect 3873 12186 3907 12220
rect 3873 12118 3907 12152
rect 3873 12050 3907 12084
rect 3873 11982 3907 12016
rect 5061 12254 5095 12288
rect 5061 12186 5095 12220
rect 5061 12118 5095 12152
rect 5061 12050 5095 12084
rect 5061 11982 5095 12016
rect 3991 11880 4025 11914
rect 4059 11880 4093 11914
rect 4127 11880 4161 11914
rect 4195 11880 4229 11914
rect 4263 11880 4297 11914
rect 4331 11880 4365 11914
rect 4399 11880 4433 11914
rect 4467 11880 4501 11914
rect 4535 11880 4569 11914
rect 4603 11880 4637 11914
rect 4671 11880 4705 11914
rect 4739 11880 4773 11914
rect 4807 11880 4841 11914
rect 4875 11880 4909 11914
rect 4943 11880 4977 11914
rect 317 11133 351 11167
rect 385 11133 419 11167
rect 453 11133 487 11167
rect 521 11133 555 11167
rect 589 11133 623 11167
rect 657 11133 691 11167
rect 725 11133 759 11167
rect 793 11133 827 11167
rect 861 11133 895 11167
rect 929 11133 963 11167
rect 997 11133 1031 11167
rect 1065 11133 1099 11167
rect 1133 11133 1167 11167
rect 1201 11133 1235 11167
rect 1269 11133 1303 11167
rect 199 11031 233 11065
rect 1387 11031 1421 11065
rect 199 10963 233 10997
rect 199 10895 233 10929
rect 199 10827 233 10861
rect 199 10759 233 10793
rect 199 10691 233 10725
rect 1387 10963 1421 10997
rect 1387 10895 1421 10929
rect 1387 10827 1421 10861
rect 1387 10759 1421 10793
rect 1387 10691 1421 10725
rect 317 10589 351 10623
rect 385 10589 419 10623
rect 453 10589 487 10623
rect 521 10589 555 10623
rect 589 10589 623 10623
rect 657 10589 691 10623
rect 725 10589 759 10623
rect 793 10589 827 10623
rect 861 10589 895 10623
rect 929 10589 963 10623
rect 997 10589 1031 10623
rect 1065 10589 1099 10623
rect 1133 10589 1167 10623
rect 1201 10589 1235 10623
rect 1269 10589 1303 10623
rect 2470 11137 2504 11171
rect 2538 11137 2572 11171
rect 2606 11137 2640 11171
rect 2674 11137 2708 11171
rect 2742 11137 2776 11171
rect 2810 11137 2844 11171
rect 2878 11137 2912 11171
rect 2946 11137 2980 11171
rect 3014 11137 3048 11171
rect 3082 11137 3116 11171
rect 3150 11137 3184 11171
rect 3218 11137 3252 11171
rect 3286 11137 3320 11171
rect 3354 11137 3388 11171
rect 3422 11137 3456 11171
rect 2352 11035 2386 11069
rect 3540 11035 3574 11069
rect 2352 10967 2386 11001
rect 2352 10899 2386 10933
rect 2352 10831 2386 10865
rect 2352 10763 2386 10797
rect 2352 10695 2386 10729
rect 3540 10967 3574 11001
rect 3540 10899 3574 10933
rect 3540 10831 3574 10865
rect 3540 10763 3574 10797
rect 3540 10695 3574 10729
rect 2470 10593 2504 10627
rect 2538 10593 2572 10627
rect 2606 10593 2640 10627
rect 2674 10593 2708 10627
rect 2742 10593 2776 10627
rect 2810 10593 2844 10627
rect 2878 10593 2912 10627
rect 2946 10593 2980 10627
rect 3014 10593 3048 10627
rect 3082 10593 3116 10627
rect 3150 10593 3184 10627
rect 3218 10593 3252 10627
rect 3286 10593 3320 10627
rect 3354 10593 3388 10627
rect 3422 10593 3456 10627
rect 3991 11137 4025 11171
rect 4059 11137 4093 11171
rect 4127 11137 4161 11171
rect 4195 11137 4229 11171
rect 4263 11137 4297 11171
rect 4331 11137 4365 11171
rect 4399 11137 4433 11171
rect 4467 11137 4501 11171
rect 4535 11137 4569 11171
rect 4603 11137 4637 11171
rect 4671 11137 4705 11171
rect 4739 11137 4773 11171
rect 4807 11137 4841 11171
rect 4875 11137 4909 11171
rect 4943 11137 4977 11171
rect 3873 11035 3907 11069
rect 5061 11035 5095 11069
rect 3873 10967 3907 11001
rect 3873 10899 3907 10933
rect 3873 10831 3907 10865
rect 3873 10763 3907 10797
rect 3873 10695 3907 10729
rect 5061 10967 5095 11001
rect 5061 10899 5095 10933
rect 5061 10831 5095 10865
rect 5061 10763 5095 10797
rect 5061 10695 5095 10729
rect 3991 10593 4025 10627
rect 4059 10593 4093 10627
rect 4127 10593 4161 10627
rect 4195 10593 4229 10627
rect 4263 10593 4297 10627
rect 4331 10593 4365 10627
rect 4399 10593 4433 10627
rect 4467 10593 4501 10627
rect 4535 10593 4569 10627
rect 4603 10593 4637 10627
rect 4671 10593 4705 10627
rect 4739 10593 4773 10627
rect 4807 10593 4841 10627
rect 4875 10593 4909 10627
rect 4943 10593 4977 10627
rect 317 9846 351 9880
rect 385 9846 419 9880
rect 453 9846 487 9880
rect 521 9846 555 9880
rect 589 9846 623 9880
rect 657 9846 691 9880
rect 725 9846 759 9880
rect 793 9846 827 9880
rect 861 9846 895 9880
rect 929 9846 963 9880
rect 997 9846 1031 9880
rect 1065 9846 1099 9880
rect 1133 9846 1167 9880
rect 1201 9846 1235 9880
rect 1269 9846 1303 9880
rect 199 9744 233 9778
rect 1387 9744 1421 9778
rect 199 9676 233 9710
rect 199 9608 233 9642
rect 199 9540 233 9574
rect 199 9472 233 9506
rect 199 9404 233 9438
rect 1387 9676 1421 9710
rect 1387 9608 1421 9642
rect 1387 9540 1421 9574
rect 1387 9472 1421 9506
rect 1387 9404 1421 9438
rect 317 9302 351 9336
rect 385 9302 419 9336
rect 453 9302 487 9336
rect 521 9302 555 9336
rect 589 9302 623 9336
rect 657 9302 691 9336
rect 725 9302 759 9336
rect 793 9302 827 9336
rect 861 9302 895 9336
rect 929 9302 963 9336
rect 997 9302 1031 9336
rect 1065 9302 1099 9336
rect 1133 9302 1167 9336
rect 1201 9302 1235 9336
rect 1269 9302 1303 9336
rect 2470 9850 2504 9884
rect 2538 9850 2572 9884
rect 2606 9850 2640 9884
rect 2674 9850 2708 9884
rect 2742 9850 2776 9884
rect 2810 9850 2844 9884
rect 2878 9850 2912 9884
rect 2946 9850 2980 9884
rect 3014 9850 3048 9884
rect 3082 9850 3116 9884
rect 3150 9850 3184 9884
rect 3218 9850 3252 9884
rect 3286 9850 3320 9884
rect 3354 9850 3388 9884
rect 3422 9850 3456 9884
rect 2352 9748 2386 9782
rect 3540 9748 3574 9782
rect 2352 9680 2386 9714
rect 2352 9612 2386 9646
rect 2352 9544 2386 9578
rect 2352 9476 2386 9510
rect 2352 9408 2386 9442
rect 3540 9680 3574 9714
rect 3540 9612 3574 9646
rect 3540 9544 3574 9578
rect 3540 9476 3574 9510
rect 3540 9408 3574 9442
rect 2470 9306 2504 9340
rect 2538 9306 2572 9340
rect 2606 9306 2640 9340
rect 2674 9306 2708 9340
rect 2742 9306 2776 9340
rect 2810 9306 2844 9340
rect 2878 9306 2912 9340
rect 2946 9306 2980 9340
rect 3014 9306 3048 9340
rect 3082 9306 3116 9340
rect 3150 9306 3184 9340
rect 3218 9306 3252 9340
rect 3286 9306 3320 9340
rect 3354 9306 3388 9340
rect 3422 9306 3456 9340
rect 3991 9850 4025 9884
rect 4059 9850 4093 9884
rect 4127 9850 4161 9884
rect 4195 9850 4229 9884
rect 4263 9850 4297 9884
rect 4331 9850 4365 9884
rect 4399 9850 4433 9884
rect 4467 9850 4501 9884
rect 4535 9850 4569 9884
rect 4603 9850 4637 9884
rect 4671 9850 4705 9884
rect 4739 9850 4773 9884
rect 4807 9850 4841 9884
rect 4875 9850 4909 9884
rect 4943 9850 4977 9884
rect 3873 9748 3907 9782
rect 5061 9748 5095 9782
rect 3873 9680 3907 9714
rect 3873 9612 3907 9646
rect 3873 9544 3907 9578
rect 3873 9476 3907 9510
rect 3873 9408 3907 9442
rect 5061 9680 5095 9714
rect 5061 9612 5095 9646
rect 5061 9544 5095 9578
rect 5061 9476 5095 9510
rect 5061 9408 5095 9442
rect 3991 9306 4025 9340
rect 4059 9306 4093 9340
rect 4127 9306 4161 9340
rect 4195 9306 4229 9340
rect 4263 9306 4297 9340
rect 4331 9306 4365 9340
rect 4399 9306 4433 9340
rect 4467 9306 4501 9340
rect 4535 9306 4569 9340
rect 4603 9306 4637 9340
rect 4671 9306 4705 9340
rect 4739 9306 4773 9340
rect 4807 9306 4841 9340
rect 4875 9306 4909 9340
rect 4943 9306 4977 9340
rect 317 8559 351 8593
rect 385 8559 419 8593
rect 453 8559 487 8593
rect 521 8559 555 8593
rect 589 8559 623 8593
rect 657 8559 691 8593
rect 725 8559 759 8593
rect 793 8559 827 8593
rect 861 8559 895 8593
rect 929 8559 963 8593
rect 997 8559 1031 8593
rect 1065 8559 1099 8593
rect 1133 8559 1167 8593
rect 1201 8559 1235 8593
rect 1269 8559 1303 8593
rect 199 8457 233 8491
rect 1387 8457 1421 8491
rect 199 8389 233 8423
rect 199 8321 233 8355
rect 199 8253 233 8287
rect 199 8185 233 8219
rect 199 8117 233 8151
rect 1387 8389 1421 8423
rect 1387 8321 1421 8355
rect 1387 8253 1421 8287
rect 1387 8185 1421 8219
rect 1387 8117 1421 8151
rect 317 8015 351 8049
rect 385 8015 419 8049
rect 453 8015 487 8049
rect 521 8015 555 8049
rect 589 8015 623 8049
rect 657 8015 691 8049
rect 725 8015 759 8049
rect 793 8015 827 8049
rect 861 8015 895 8049
rect 929 8015 963 8049
rect 997 8015 1031 8049
rect 1065 8015 1099 8049
rect 1133 8015 1167 8049
rect 1201 8015 1235 8049
rect 1269 8015 1303 8049
rect 2470 8563 2504 8597
rect 2538 8563 2572 8597
rect 2606 8563 2640 8597
rect 2674 8563 2708 8597
rect 2742 8563 2776 8597
rect 2810 8563 2844 8597
rect 2878 8563 2912 8597
rect 2946 8563 2980 8597
rect 3014 8563 3048 8597
rect 3082 8563 3116 8597
rect 3150 8563 3184 8597
rect 3218 8563 3252 8597
rect 3286 8563 3320 8597
rect 3354 8563 3388 8597
rect 3422 8563 3456 8597
rect 2352 8461 2386 8495
rect 3540 8461 3574 8495
rect 2352 8393 2386 8427
rect 2352 8325 2386 8359
rect 2352 8257 2386 8291
rect 2352 8189 2386 8223
rect 2352 8121 2386 8155
rect 3540 8393 3574 8427
rect 3540 8325 3574 8359
rect 3540 8257 3574 8291
rect 3540 8189 3574 8223
rect 3540 8121 3574 8155
rect 2470 8019 2504 8053
rect 2538 8019 2572 8053
rect 2606 8019 2640 8053
rect 2674 8019 2708 8053
rect 2742 8019 2776 8053
rect 2810 8019 2844 8053
rect 2878 8019 2912 8053
rect 2946 8019 2980 8053
rect 3014 8019 3048 8053
rect 3082 8019 3116 8053
rect 3150 8019 3184 8053
rect 3218 8019 3252 8053
rect 3286 8019 3320 8053
rect 3354 8019 3388 8053
rect 3422 8019 3456 8053
rect 3991 8563 4025 8597
rect 4059 8563 4093 8597
rect 4127 8563 4161 8597
rect 4195 8563 4229 8597
rect 4263 8563 4297 8597
rect 4331 8563 4365 8597
rect 4399 8563 4433 8597
rect 4467 8563 4501 8597
rect 4535 8563 4569 8597
rect 4603 8563 4637 8597
rect 4671 8563 4705 8597
rect 4739 8563 4773 8597
rect 4807 8563 4841 8597
rect 4875 8563 4909 8597
rect 4943 8563 4977 8597
rect 3873 8461 3907 8495
rect 5061 8461 5095 8495
rect 3873 8393 3907 8427
rect 3873 8325 3907 8359
rect 3873 8257 3907 8291
rect 3873 8189 3907 8223
rect 3873 8121 3907 8155
rect 5061 8393 5095 8427
rect 5061 8325 5095 8359
rect 5061 8257 5095 8291
rect 5061 8189 5095 8223
rect 5061 8121 5095 8155
rect 3991 8019 4025 8053
rect 4059 8019 4093 8053
rect 4127 8019 4161 8053
rect 4195 8019 4229 8053
rect 4263 8019 4297 8053
rect 4331 8019 4365 8053
rect 4399 8019 4433 8053
rect 4467 8019 4501 8053
rect 4535 8019 4569 8053
rect 4603 8019 4637 8053
rect 4671 8019 4705 8053
rect 4739 8019 4773 8053
rect 4807 8019 4841 8053
rect 4875 8019 4909 8053
rect 4943 8019 4977 8053
rect 317 7272 351 7306
rect 385 7272 419 7306
rect 453 7272 487 7306
rect 521 7272 555 7306
rect 589 7272 623 7306
rect 657 7272 691 7306
rect 725 7272 759 7306
rect 793 7272 827 7306
rect 861 7272 895 7306
rect 929 7272 963 7306
rect 997 7272 1031 7306
rect 1065 7272 1099 7306
rect 1133 7272 1167 7306
rect 1201 7272 1235 7306
rect 1269 7272 1303 7306
rect 199 7170 233 7204
rect 1387 7170 1421 7204
rect 199 7102 233 7136
rect 199 7034 233 7068
rect 199 6966 233 7000
rect 199 6898 233 6932
rect 199 6830 233 6864
rect 1387 7102 1421 7136
rect 1387 7034 1421 7068
rect 1387 6966 1421 7000
rect 1387 6898 1421 6932
rect 1387 6830 1421 6864
rect 317 6728 351 6762
rect 385 6728 419 6762
rect 453 6728 487 6762
rect 521 6728 555 6762
rect 589 6728 623 6762
rect 657 6728 691 6762
rect 725 6728 759 6762
rect 793 6728 827 6762
rect 861 6728 895 6762
rect 929 6728 963 6762
rect 997 6728 1031 6762
rect 1065 6728 1099 6762
rect 1133 6728 1167 6762
rect 1201 6728 1235 6762
rect 1269 6728 1303 6762
rect 2470 7276 2504 7310
rect 2538 7276 2572 7310
rect 2606 7276 2640 7310
rect 2674 7276 2708 7310
rect 2742 7276 2776 7310
rect 2810 7276 2844 7310
rect 2878 7276 2912 7310
rect 2946 7276 2980 7310
rect 3014 7276 3048 7310
rect 3082 7276 3116 7310
rect 3150 7276 3184 7310
rect 3218 7276 3252 7310
rect 3286 7276 3320 7310
rect 3354 7276 3388 7310
rect 3422 7276 3456 7310
rect 2352 7174 2386 7208
rect 3540 7174 3574 7208
rect 2352 7106 2386 7140
rect 2352 7038 2386 7072
rect 2352 6970 2386 7004
rect 2352 6902 2386 6936
rect 2352 6834 2386 6868
rect 3540 7106 3574 7140
rect 3540 7038 3574 7072
rect 3540 6970 3574 7004
rect 3540 6902 3574 6936
rect 3540 6834 3574 6868
rect 2470 6732 2504 6766
rect 2538 6732 2572 6766
rect 2606 6732 2640 6766
rect 2674 6732 2708 6766
rect 2742 6732 2776 6766
rect 2810 6732 2844 6766
rect 2878 6732 2912 6766
rect 2946 6732 2980 6766
rect 3014 6732 3048 6766
rect 3082 6732 3116 6766
rect 3150 6732 3184 6766
rect 3218 6732 3252 6766
rect 3286 6732 3320 6766
rect 3354 6732 3388 6766
rect 3422 6732 3456 6766
rect 3991 7276 4025 7310
rect 4059 7276 4093 7310
rect 4127 7276 4161 7310
rect 4195 7276 4229 7310
rect 4263 7276 4297 7310
rect 4331 7276 4365 7310
rect 4399 7276 4433 7310
rect 4467 7276 4501 7310
rect 4535 7276 4569 7310
rect 4603 7276 4637 7310
rect 4671 7276 4705 7310
rect 4739 7276 4773 7310
rect 4807 7276 4841 7310
rect 4875 7276 4909 7310
rect 4943 7276 4977 7310
rect 3873 7174 3907 7208
rect 5061 7174 5095 7208
rect 3873 7106 3907 7140
rect 3873 7038 3907 7072
rect 3873 6970 3907 7004
rect 3873 6902 3907 6936
rect 3873 6834 3907 6868
rect 5061 7106 5095 7140
rect 5061 7038 5095 7072
rect 5061 6970 5095 7004
rect 5061 6902 5095 6936
rect 5061 6834 5095 6868
rect 3991 6732 4025 6766
rect 4059 6732 4093 6766
rect 4127 6732 4161 6766
rect 4195 6732 4229 6766
rect 4263 6732 4297 6766
rect 4331 6732 4365 6766
rect 4399 6732 4433 6766
rect 4467 6732 4501 6766
rect 4535 6732 4569 6766
rect 4603 6732 4637 6766
rect 4671 6732 4705 6766
rect 4739 6732 4773 6766
rect 4807 6732 4841 6766
rect 4875 6732 4909 6766
rect 4943 6732 4977 6766
rect 317 5985 351 6019
rect 385 5985 419 6019
rect 453 5985 487 6019
rect 521 5985 555 6019
rect 589 5985 623 6019
rect 657 5985 691 6019
rect 725 5985 759 6019
rect 793 5985 827 6019
rect 861 5985 895 6019
rect 929 5985 963 6019
rect 997 5985 1031 6019
rect 1065 5985 1099 6019
rect 1133 5985 1167 6019
rect 1201 5985 1235 6019
rect 1269 5985 1303 6019
rect 199 5883 233 5917
rect 1387 5883 1421 5917
rect 199 5815 233 5849
rect 199 5747 233 5781
rect 199 5679 233 5713
rect 199 5611 233 5645
rect 199 5543 233 5577
rect 1387 5815 1421 5849
rect 1387 5747 1421 5781
rect 1387 5679 1421 5713
rect 1387 5611 1421 5645
rect 1387 5543 1421 5577
rect 317 5441 351 5475
rect 385 5441 419 5475
rect 453 5441 487 5475
rect 521 5441 555 5475
rect 589 5441 623 5475
rect 657 5441 691 5475
rect 725 5441 759 5475
rect 793 5441 827 5475
rect 861 5441 895 5475
rect 929 5441 963 5475
rect 997 5441 1031 5475
rect 1065 5441 1099 5475
rect 1133 5441 1167 5475
rect 1201 5441 1235 5475
rect 1269 5441 1303 5475
rect 2470 5989 2504 6023
rect 2538 5989 2572 6023
rect 2606 5989 2640 6023
rect 2674 5989 2708 6023
rect 2742 5989 2776 6023
rect 2810 5989 2844 6023
rect 2878 5989 2912 6023
rect 2946 5989 2980 6023
rect 3014 5989 3048 6023
rect 3082 5989 3116 6023
rect 3150 5989 3184 6023
rect 3218 5989 3252 6023
rect 3286 5989 3320 6023
rect 3354 5989 3388 6023
rect 3422 5989 3456 6023
rect 2352 5887 2386 5921
rect 3540 5887 3574 5921
rect 2352 5819 2386 5853
rect 2352 5751 2386 5785
rect 2352 5683 2386 5717
rect 2352 5615 2386 5649
rect 2352 5547 2386 5581
rect 3540 5819 3574 5853
rect 3540 5751 3574 5785
rect 3540 5683 3574 5717
rect 3540 5615 3574 5649
rect 3540 5547 3574 5581
rect 2470 5445 2504 5479
rect 2538 5445 2572 5479
rect 2606 5445 2640 5479
rect 2674 5445 2708 5479
rect 2742 5445 2776 5479
rect 2810 5445 2844 5479
rect 2878 5445 2912 5479
rect 2946 5445 2980 5479
rect 3014 5445 3048 5479
rect 3082 5445 3116 5479
rect 3150 5445 3184 5479
rect 3218 5445 3252 5479
rect 3286 5445 3320 5479
rect 3354 5445 3388 5479
rect 3422 5445 3456 5479
rect 3991 5989 4025 6023
rect 4059 5989 4093 6023
rect 4127 5989 4161 6023
rect 4195 5989 4229 6023
rect 4263 5989 4297 6023
rect 4331 5989 4365 6023
rect 4399 5989 4433 6023
rect 4467 5989 4501 6023
rect 4535 5989 4569 6023
rect 4603 5989 4637 6023
rect 4671 5989 4705 6023
rect 4739 5989 4773 6023
rect 4807 5989 4841 6023
rect 4875 5989 4909 6023
rect 4943 5989 4977 6023
rect 3873 5887 3907 5921
rect 5061 5887 5095 5921
rect 3873 5819 3907 5853
rect 3873 5751 3907 5785
rect 3873 5683 3907 5717
rect 3873 5615 3907 5649
rect 3873 5547 3907 5581
rect 5061 5819 5095 5853
rect 5061 5751 5095 5785
rect 5061 5683 5095 5717
rect 5061 5615 5095 5649
rect 5061 5547 5095 5581
rect 3991 5445 4025 5479
rect 4059 5445 4093 5479
rect 4127 5445 4161 5479
rect 4195 5445 4229 5479
rect 4263 5445 4297 5479
rect 4331 5445 4365 5479
rect 4399 5445 4433 5479
rect 4467 5445 4501 5479
rect 4535 5445 4569 5479
rect 4603 5445 4637 5479
rect 4671 5445 4705 5479
rect 4739 5445 4773 5479
rect 4807 5445 4841 5479
rect 4875 5445 4909 5479
rect 4943 5445 4977 5479
rect 317 4698 351 4732
rect 385 4698 419 4732
rect 453 4698 487 4732
rect 521 4698 555 4732
rect 589 4698 623 4732
rect 657 4698 691 4732
rect 725 4698 759 4732
rect 793 4698 827 4732
rect 861 4698 895 4732
rect 929 4698 963 4732
rect 997 4698 1031 4732
rect 1065 4698 1099 4732
rect 1133 4698 1167 4732
rect 1201 4698 1235 4732
rect 1269 4698 1303 4732
rect 199 4596 233 4630
rect 1387 4596 1421 4630
rect 199 4528 233 4562
rect 199 4460 233 4494
rect 199 4392 233 4426
rect 199 4324 233 4358
rect 199 4256 233 4290
rect 1387 4528 1421 4562
rect 1387 4460 1421 4494
rect 1387 4392 1421 4426
rect 1387 4324 1421 4358
rect 1387 4256 1421 4290
rect 317 4154 351 4188
rect 385 4154 419 4188
rect 453 4154 487 4188
rect 521 4154 555 4188
rect 589 4154 623 4188
rect 657 4154 691 4188
rect 725 4154 759 4188
rect 793 4154 827 4188
rect 861 4154 895 4188
rect 929 4154 963 4188
rect 997 4154 1031 4188
rect 1065 4154 1099 4188
rect 1133 4154 1167 4188
rect 1201 4154 1235 4188
rect 1269 4154 1303 4188
rect 2470 4702 2504 4736
rect 2538 4702 2572 4736
rect 2606 4702 2640 4736
rect 2674 4702 2708 4736
rect 2742 4702 2776 4736
rect 2810 4702 2844 4736
rect 2878 4702 2912 4736
rect 2946 4702 2980 4736
rect 3014 4702 3048 4736
rect 3082 4702 3116 4736
rect 3150 4702 3184 4736
rect 3218 4702 3252 4736
rect 3286 4702 3320 4736
rect 3354 4702 3388 4736
rect 3422 4702 3456 4736
rect 2352 4600 2386 4634
rect 3540 4600 3574 4634
rect 2352 4532 2386 4566
rect 2352 4464 2386 4498
rect 2352 4396 2386 4430
rect 2352 4328 2386 4362
rect 2352 4260 2386 4294
rect 3540 4532 3574 4566
rect 3540 4464 3574 4498
rect 3540 4396 3574 4430
rect 3540 4328 3574 4362
rect 3540 4260 3574 4294
rect 2470 4158 2504 4192
rect 2538 4158 2572 4192
rect 2606 4158 2640 4192
rect 2674 4158 2708 4192
rect 2742 4158 2776 4192
rect 2810 4158 2844 4192
rect 2878 4158 2912 4192
rect 2946 4158 2980 4192
rect 3014 4158 3048 4192
rect 3082 4158 3116 4192
rect 3150 4158 3184 4192
rect 3218 4158 3252 4192
rect 3286 4158 3320 4192
rect 3354 4158 3388 4192
rect 3422 4158 3456 4192
rect 3991 4702 4025 4736
rect 4059 4702 4093 4736
rect 4127 4702 4161 4736
rect 4195 4702 4229 4736
rect 4263 4702 4297 4736
rect 4331 4702 4365 4736
rect 4399 4702 4433 4736
rect 4467 4702 4501 4736
rect 4535 4702 4569 4736
rect 4603 4702 4637 4736
rect 4671 4702 4705 4736
rect 4739 4702 4773 4736
rect 4807 4702 4841 4736
rect 4875 4702 4909 4736
rect 4943 4702 4977 4736
rect 3873 4600 3907 4634
rect 5061 4600 5095 4634
rect 3873 4532 3907 4566
rect 3873 4464 3907 4498
rect 3873 4396 3907 4430
rect 3873 4328 3907 4362
rect 3873 4260 3907 4294
rect 5061 4532 5095 4566
rect 5061 4464 5095 4498
rect 5061 4396 5095 4430
rect 5061 4328 5095 4362
rect 5061 4260 5095 4294
rect 3991 4158 4025 4192
rect 4059 4158 4093 4192
rect 4127 4158 4161 4192
rect 4195 4158 4229 4192
rect 4263 4158 4297 4192
rect 4331 4158 4365 4192
rect 4399 4158 4433 4192
rect 4467 4158 4501 4192
rect 4535 4158 4569 4192
rect 4603 4158 4637 4192
rect 4671 4158 4705 4192
rect 4739 4158 4773 4192
rect 4807 4158 4841 4192
rect 4875 4158 4909 4192
rect 4943 4158 4977 4192
rect 317 3411 351 3445
rect 385 3411 419 3445
rect 453 3411 487 3445
rect 521 3411 555 3445
rect 589 3411 623 3445
rect 657 3411 691 3445
rect 725 3411 759 3445
rect 793 3411 827 3445
rect 861 3411 895 3445
rect 929 3411 963 3445
rect 997 3411 1031 3445
rect 1065 3411 1099 3445
rect 1133 3411 1167 3445
rect 1201 3411 1235 3445
rect 1269 3411 1303 3445
rect 199 3309 233 3343
rect 1387 3309 1421 3343
rect 199 3241 233 3275
rect 199 3173 233 3207
rect 199 3105 233 3139
rect 199 3037 233 3071
rect 199 2969 233 3003
rect 1387 3241 1421 3275
rect 1387 3173 1421 3207
rect 1387 3105 1421 3139
rect 1387 3037 1421 3071
rect 1387 2969 1421 3003
rect 317 2867 351 2901
rect 385 2867 419 2901
rect 453 2867 487 2901
rect 521 2867 555 2901
rect 589 2867 623 2901
rect 657 2867 691 2901
rect 725 2867 759 2901
rect 793 2867 827 2901
rect 861 2867 895 2901
rect 929 2867 963 2901
rect 997 2867 1031 2901
rect 1065 2867 1099 2901
rect 1133 2867 1167 2901
rect 1201 2867 1235 2901
rect 1269 2867 1303 2901
rect 2470 3415 2504 3449
rect 2538 3415 2572 3449
rect 2606 3415 2640 3449
rect 2674 3415 2708 3449
rect 2742 3415 2776 3449
rect 2810 3415 2844 3449
rect 2878 3415 2912 3449
rect 2946 3415 2980 3449
rect 3014 3415 3048 3449
rect 3082 3415 3116 3449
rect 3150 3415 3184 3449
rect 3218 3415 3252 3449
rect 3286 3415 3320 3449
rect 3354 3415 3388 3449
rect 3422 3415 3456 3449
rect 2352 3313 2386 3347
rect 3540 3313 3574 3347
rect 2352 3245 2386 3279
rect 2352 3177 2386 3211
rect 2352 3109 2386 3143
rect 2352 3041 2386 3075
rect 2352 2973 2386 3007
rect 3540 3245 3574 3279
rect 3540 3177 3574 3211
rect 3540 3109 3574 3143
rect 3540 3041 3574 3075
rect 3540 2973 3574 3007
rect 2470 2871 2504 2905
rect 2538 2871 2572 2905
rect 2606 2871 2640 2905
rect 2674 2871 2708 2905
rect 2742 2871 2776 2905
rect 2810 2871 2844 2905
rect 2878 2871 2912 2905
rect 2946 2871 2980 2905
rect 3014 2871 3048 2905
rect 3082 2871 3116 2905
rect 3150 2871 3184 2905
rect 3218 2871 3252 2905
rect 3286 2871 3320 2905
rect 3354 2871 3388 2905
rect 3422 2871 3456 2905
rect 3991 3415 4025 3449
rect 4059 3415 4093 3449
rect 4127 3415 4161 3449
rect 4195 3415 4229 3449
rect 4263 3415 4297 3449
rect 4331 3415 4365 3449
rect 4399 3415 4433 3449
rect 4467 3415 4501 3449
rect 4535 3415 4569 3449
rect 4603 3415 4637 3449
rect 4671 3415 4705 3449
rect 4739 3415 4773 3449
rect 4807 3415 4841 3449
rect 4875 3415 4909 3449
rect 4943 3415 4977 3449
rect 3873 3313 3907 3347
rect 5061 3313 5095 3347
rect 3873 3245 3907 3279
rect 3873 3177 3907 3211
rect 3873 3109 3907 3143
rect 3873 3041 3907 3075
rect 3873 2973 3907 3007
rect 5061 3245 5095 3279
rect 5061 3177 5095 3211
rect 5061 3109 5095 3143
rect 5061 3041 5095 3075
rect 5061 2973 5095 3007
rect 3991 2871 4025 2905
rect 4059 2871 4093 2905
rect 4127 2871 4161 2905
rect 4195 2871 4229 2905
rect 4263 2871 4297 2905
rect 4331 2871 4365 2905
rect 4399 2871 4433 2905
rect 4467 2871 4501 2905
rect 4535 2871 4569 2905
rect 4603 2871 4637 2905
rect 4671 2871 4705 2905
rect 4739 2871 4773 2905
rect 4807 2871 4841 2905
rect 4875 2871 4909 2905
rect 4943 2871 4977 2905
rect 317 2124 351 2158
rect 385 2124 419 2158
rect 453 2124 487 2158
rect 521 2124 555 2158
rect 589 2124 623 2158
rect 657 2124 691 2158
rect 725 2124 759 2158
rect 793 2124 827 2158
rect 861 2124 895 2158
rect 929 2124 963 2158
rect 997 2124 1031 2158
rect 1065 2124 1099 2158
rect 1133 2124 1167 2158
rect 1201 2124 1235 2158
rect 1269 2124 1303 2158
rect 199 2022 233 2056
rect 1387 2022 1421 2056
rect 199 1954 233 1988
rect 199 1886 233 1920
rect 199 1818 233 1852
rect 199 1750 233 1784
rect 199 1682 233 1716
rect 1387 1954 1421 1988
rect 1387 1886 1421 1920
rect 1387 1818 1421 1852
rect 1387 1750 1421 1784
rect 1387 1682 1421 1716
rect 317 1580 351 1614
rect 385 1580 419 1614
rect 453 1580 487 1614
rect 521 1580 555 1614
rect 589 1580 623 1614
rect 657 1580 691 1614
rect 725 1580 759 1614
rect 793 1580 827 1614
rect 861 1580 895 1614
rect 929 1580 963 1614
rect 997 1580 1031 1614
rect 1065 1580 1099 1614
rect 1133 1580 1167 1614
rect 1201 1580 1235 1614
rect 1269 1580 1303 1614
rect 2470 2128 2504 2162
rect 2538 2128 2572 2162
rect 2606 2128 2640 2162
rect 2674 2128 2708 2162
rect 2742 2128 2776 2162
rect 2810 2128 2844 2162
rect 2878 2128 2912 2162
rect 2946 2128 2980 2162
rect 3014 2128 3048 2162
rect 3082 2128 3116 2162
rect 3150 2128 3184 2162
rect 3218 2128 3252 2162
rect 3286 2128 3320 2162
rect 3354 2128 3388 2162
rect 3422 2128 3456 2162
rect 2352 2026 2386 2060
rect 3540 2026 3574 2060
rect 2352 1958 2386 1992
rect 2352 1890 2386 1924
rect 2352 1822 2386 1856
rect 2352 1754 2386 1788
rect 2352 1686 2386 1720
rect 3540 1958 3574 1992
rect 3540 1890 3574 1924
rect 3540 1822 3574 1856
rect 3540 1754 3574 1788
rect 3540 1686 3574 1720
rect 2470 1584 2504 1618
rect 2538 1584 2572 1618
rect 2606 1584 2640 1618
rect 2674 1584 2708 1618
rect 2742 1584 2776 1618
rect 2810 1584 2844 1618
rect 2878 1584 2912 1618
rect 2946 1584 2980 1618
rect 3014 1584 3048 1618
rect 3082 1584 3116 1618
rect 3150 1584 3184 1618
rect 3218 1584 3252 1618
rect 3286 1584 3320 1618
rect 3354 1584 3388 1618
rect 3422 1584 3456 1618
rect 3991 2128 4025 2162
rect 4059 2128 4093 2162
rect 4127 2128 4161 2162
rect 4195 2128 4229 2162
rect 4263 2128 4297 2162
rect 4331 2128 4365 2162
rect 4399 2128 4433 2162
rect 4467 2128 4501 2162
rect 4535 2128 4569 2162
rect 4603 2128 4637 2162
rect 4671 2128 4705 2162
rect 4739 2128 4773 2162
rect 4807 2128 4841 2162
rect 4875 2128 4909 2162
rect 4943 2128 4977 2162
rect 3873 2026 3907 2060
rect 5061 2026 5095 2060
rect 3873 1958 3907 1992
rect 3873 1890 3907 1924
rect 3873 1822 3907 1856
rect 3873 1754 3907 1788
rect 3873 1686 3907 1720
rect 5061 1958 5095 1992
rect 5061 1890 5095 1924
rect 5061 1822 5095 1856
rect 5061 1754 5095 1788
rect 5061 1686 5095 1720
rect 3991 1584 4025 1618
rect 4059 1584 4093 1618
rect 4127 1584 4161 1618
rect 4195 1584 4229 1618
rect 4263 1584 4297 1618
rect 4331 1584 4365 1618
rect 4399 1584 4433 1618
rect 4467 1584 4501 1618
rect 4535 1584 4569 1618
rect 4603 1584 4637 1618
rect 4671 1584 4705 1618
rect 4739 1584 4773 1618
rect 4807 1584 4841 1618
rect 4875 1584 4909 1618
rect 4943 1584 4977 1618
<< poly >>
rect 297 41953 1323 41969
rect 297 41919 313 41953
rect 347 41919 505 41953
rect 539 41919 697 41953
rect 731 41919 889 41953
rect 923 41919 1081 41953
rect 1115 41919 1273 41953
rect 1307 41919 1323 41953
rect 297 41903 1323 41919
rect 363 41871 393 41903
rect 459 41871 489 41903
rect 555 41871 585 41903
rect 651 41871 681 41903
rect 747 41871 777 41903
rect 843 41871 873 41903
rect 939 41871 969 41903
rect 1035 41871 1065 41903
rect 1131 41871 1161 41903
rect 1227 41871 1257 41903
rect 363 41573 393 41599
rect 459 41573 489 41599
rect 555 41573 585 41599
rect 651 41573 681 41599
rect 747 41573 777 41599
rect 843 41573 873 41599
rect 939 41573 969 41599
rect 1035 41573 1065 41599
rect 1131 41573 1161 41599
rect 1227 41573 1257 41599
rect 2450 41957 3476 41973
rect 2450 41923 2466 41957
rect 2500 41923 2658 41957
rect 2692 41923 2850 41957
rect 2884 41923 3042 41957
rect 3076 41923 3234 41957
rect 3268 41923 3426 41957
rect 3460 41923 3476 41957
rect 2450 41907 3476 41923
rect 2516 41875 2546 41907
rect 2612 41875 2642 41907
rect 2708 41875 2738 41907
rect 2804 41875 2834 41907
rect 2900 41875 2930 41907
rect 2996 41875 3026 41907
rect 3092 41875 3122 41907
rect 3188 41875 3218 41907
rect 3284 41875 3314 41907
rect 3380 41875 3410 41907
rect 2516 41577 2546 41603
rect 2612 41577 2642 41603
rect 2708 41577 2738 41603
rect 2804 41577 2834 41603
rect 2900 41577 2930 41603
rect 2996 41577 3026 41603
rect 3092 41577 3122 41603
rect 3188 41577 3218 41603
rect 3284 41577 3314 41603
rect 3380 41577 3410 41603
rect 3971 41957 4997 41973
rect 3971 41923 3987 41957
rect 4021 41923 4179 41957
rect 4213 41923 4371 41957
rect 4405 41923 4563 41957
rect 4597 41923 4755 41957
rect 4789 41923 4947 41957
rect 4981 41923 4997 41957
rect 3971 41907 4997 41923
rect 4037 41875 4067 41907
rect 4133 41875 4163 41907
rect 4229 41875 4259 41907
rect 4325 41875 4355 41907
rect 4421 41875 4451 41907
rect 4517 41875 4547 41907
rect 4613 41875 4643 41907
rect 4709 41875 4739 41907
rect 4805 41875 4835 41907
rect 4901 41875 4931 41907
rect 5400 41662 5430 41688
rect 4037 41577 4067 41603
rect 4133 41577 4163 41603
rect 4229 41577 4259 41603
rect 4325 41577 4355 41603
rect 4421 41577 4451 41603
rect 4517 41577 4547 41603
rect 4613 41577 4643 41603
rect 4709 41577 4739 41603
rect 4805 41577 4835 41603
rect 4901 41577 4931 41603
rect 5400 41430 5430 41462
rect 5400 41414 5486 41430
rect 363 41291 393 41317
rect 459 41291 489 41317
rect 555 41291 585 41317
rect 651 41291 681 41317
rect 747 41291 777 41317
rect 843 41291 873 41317
rect 939 41291 969 41317
rect 1035 41291 1065 41317
rect 1131 41291 1161 41317
rect 1227 41291 1257 41317
rect 363 41165 393 41187
rect 459 41165 489 41187
rect 555 41165 585 41187
rect 651 41165 681 41187
rect 747 41165 777 41187
rect 843 41165 873 41187
rect 939 41165 969 41187
rect 1035 41165 1065 41187
rect 1131 41165 1161 41187
rect 1227 41165 1257 41187
rect 297 41145 1323 41165
rect 297 41111 313 41145
rect 347 41111 505 41145
rect 539 41111 697 41145
rect 731 41111 889 41145
rect 923 41111 1081 41145
rect 1115 41111 1273 41145
rect 1307 41111 1323 41145
rect 297 41099 1323 41111
rect 2516 41295 2546 41321
rect 2612 41295 2642 41321
rect 2708 41295 2738 41321
rect 2804 41295 2834 41321
rect 2900 41295 2930 41321
rect 2996 41295 3026 41321
rect 3092 41295 3122 41321
rect 3188 41295 3218 41321
rect 3284 41295 3314 41321
rect 3380 41295 3410 41321
rect 3675 41371 3741 41387
rect 3675 41337 3691 41371
rect 3725 41337 3741 41371
rect 3675 41321 3741 41337
rect 3693 41299 3723 41321
rect 4037 41295 4067 41321
rect 4133 41295 4163 41321
rect 4229 41295 4259 41321
rect 4325 41295 4355 41321
rect 4421 41295 4451 41321
rect 4517 41295 4547 41321
rect 4613 41295 4643 41321
rect 4709 41295 4739 41321
rect 4805 41295 4835 41321
rect 4901 41295 4931 41321
rect 5400 41380 5436 41414
rect 5470 41380 5486 41414
rect 5400 41364 5486 41380
rect 5400 41342 5430 41364
rect 2516 41169 2546 41191
rect 2612 41169 2642 41191
rect 2708 41169 2738 41191
rect 2804 41169 2834 41191
rect 2900 41169 2930 41191
rect 2996 41169 3026 41191
rect 3092 41169 3122 41191
rect 3188 41169 3218 41191
rect 3284 41169 3314 41191
rect 3380 41169 3410 41191
rect 2450 41149 3476 41169
rect 2450 41115 2466 41149
rect 2500 41115 2658 41149
rect 2692 41115 2850 41149
rect 2884 41115 3042 41149
rect 3076 41115 3234 41149
rect 3268 41115 3426 41149
rect 3460 41115 3476 41149
rect 2450 41103 3476 41115
rect 3693 41173 3723 41199
rect 4037 41169 4067 41191
rect 4133 41169 4163 41191
rect 4229 41169 4259 41191
rect 4325 41169 4355 41191
rect 4421 41169 4451 41191
rect 4517 41169 4547 41191
rect 4613 41169 4643 41191
rect 4709 41169 4739 41191
rect 4805 41169 4835 41191
rect 4901 41169 4931 41191
rect 3971 41149 4997 41169
rect 3971 41115 3987 41149
rect 4021 41115 4179 41149
rect 4213 41115 4371 41149
rect 4405 41115 4563 41149
rect 4597 41115 4755 41149
rect 4789 41115 4947 41149
rect 4981 41115 4997 41149
rect 3971 41103 4997 41115
rect 5400 41186 5430 41212
rect 297 40666 1323 40682
rect 297 40632 313 40666
rect 347 40632 505 40666
rect 539 40632 697 40666
rect 731 40632 889 40666
rect 923 40632 1081 40666
rect 1115 40632 1273 40666
rect 1307 40632 1323 40666
rect 297 40616 1323 40632
rect 363 40584 393 40616
rect 459 40584 489 40616
rect 555 40584 585 40616
rect 651 40584 681 40616
rect 747 40584 777 40616
rect 843 40584 873 40616
rect 939 40584 969 40616
rect 1035 40584 1065 40616
rect 1131 40584 1161 40616
rect 1227 40584 1257 40616
rect 363 40286 393 40312
rect 459 40286 489 40312
rect 555 40286 585 40312
rect 651 40286 681 40312
rect 747 40286 777 40312
rect 843 40286 873 40312
rect 939 40286 969 40312
rect 1035 40286 1065 40312
rect 1131 40286 1161 40312
rect 1227 40286 1257 40312
rect 2450 40670 3476 40686
rect 2450 40636 2466 40670
rect 2500 40636 2658 40670
rect 2692 40636 2850 40670
rect 2884 40636 3042 40670
rect 3076 40636 3234 40670
rect 3268 40636 3426 40670
rect 3460 40636 3476 40670
rect 2450 40620 3476 40636
rect 2516 40588 2546 40620
rect 2612 40588 2642 40620
rect 2708 40588 2738 40620
rect 2804 40588 2834 40620
rect 2900 40588 2930 40620
rect 2996 40588 3026 40620
rect 3092 40588 3122 40620
rect 3188 40588 3218 40620
rect 3284 40588 3314 40620
rect 3380 40588 3410 40620
rect 2516 40290 2546 40316
rect 2612 40290 2642 40316
rect 2708 40290 2738 40316
rect 2804 40290 2834 40316
rect 2900 40290 2930 40316
rect 2996 40290 3026 40316
rect 3092 40290 3122 40316
rect 3188 40290 3218 40316
rect 3284 40290 3314 40316
rect 3380 40290 3410 40316
rect 3971 40670 4997 40686
rect 3971 40636 3987 40670
rect 4021 40636 4179 40670
rect 4213 40636 4371 40670
rect 4405 40636 4563 40670
rect 4597 40636 4755 40670
rect 4789 40636 4947 40670
rect 4981 40636 4997 40670
rect 3971 40620 4997 40636
rect 4037 40588 4067 40620
rect 4133 40588 4163 40620
rect 4229 40588 4259 40620
rect 4325 40588 4355 40620
rect 4421 40588 4451 40620
rect 4517 40588 4547 40620
rect 4613 40588 4643 40620
rect 4709 40588 4739 40620
rect 4805 40588 4835 40620
rect 4901 40588 4931 40620
rect 5400 40375 5430 40401
rect 4037 40290 4067 40316
rect 4133 40290 4163 40316
rect 4229 40290 4259 40316
rect 4325 40290 4355 40316
rect 4421 40290 4451 40316
rect 4517 40290 4547 40316
rect 4613 40290 4643 40316
rect 4709 40290 4739 40316
rect 4805 40290 4835 40316
rect 4901 40290 4931 40316
rect 5400 40143 5430 40175
rect 5400 40127 5486 40143
rect 363 40004 393 40030
rect 459 40004 489 40030
rect 555 40004 585 40030
rect 651 40004 681 40030
rect 747 40004 777 40030
rect 843 40004 873 40030
rect 939 40004 969 40030
rect 1035 40004 1065 40030
rect 1131 40004 1161 40030
rect 1227 40004 1257 40030
rect 363 39878 393 39900
rect 459 39878 489 39900
rect 555 39878 585 39900
rect 651 39878 681 39900
rect 747 39878 777 39900
rect 843 39878 873 39900
rect 939 39878 969 39900
rect 1035 39878 1065 39900
rect 1131 39878 1161 39900
rect 1227 39878 1257 39900
rect 297 39858 1323 39878
rect 297 39824 313 39858
rect 347 39824 505 39858
rect 539 39824 697 39858
rect 731 39824 889 39858
rect 923 39824 1081 39858
rect 1115 39824 1273 39858
rect 1307 39824 1323 39858
rect 297 39812 1323 39824
rect 2516 40008 2546 40034
rect 2612 40008 2642 40034
rect 2708 40008 2738 40034
rect 2804 40008 2834 40034
rect 2900 40008 2930 40034
rect 2996 40008 3026 40034
rect 3092 40008 3122 40034
rect 3188 40008 3218 40034
rect 3284 40008 3314 40034
rect 3380 40008 3410 40034
rect 3675 40084 3741 40100
rect 3675 40050 3691 40084
rect 3725 40050 3741 40084
rect 3675 40034 3741 40050
rect 3693 40012 3723 40034
rect 4037 40008 4067 40034
rect 4133 40008 4163 40034
rect 4229 40008 4259 40034
rect 4325 40008 4355 40034
rect 4421 40008 4451 40034
rect 4517 40008 4547 40034
rect 4613 40008 4643 40034
rect 4709 40008 4739 40034
rect 4805 40008 4835 40034
rect 4901 40008 4931 40034
rect 5400 40093 5436 40127
rect 5470 40093 5486 40127
rect 5400 40077 5486 40093
rect 5400 40055 5430 40077
rect 2516 39882 2546 39904
rect 2612 39882 2642 39904
rect 2708 39882 2738 39904
rect 2804 39882 2834 39904
rect 2900 39882 2930 39904
rect 2996 39882 3026 39904
rect 3092 39882 3122 39904
rect 3188 39882 3218 39904
rect 3284 39882 3314 39904
rect 3380 39882 3410 39904
rect 2450 39862 3476 39882
rect 2450 39828 2466 39862
rect 2500 39828 2658 39862
rect 2692 39828 2850 39862
rect 2884 39828 3042 39862
rect 3076 39828 3234 39862
rect 3268 39828 3426 39862
rect 3460 39828 3476 39862
rect 2450 39816 3476 39828
rect 3693 39886 3723 39912
rect 4037 39882 4067 39904
rect 4133 39882 4163 39904
rect 4229 39882 4259 39904
rect 4325 39882 4355 39904
rect 4421 39882 4451 39904
rect 4517 39882 4547 39904
rect 4613 39882 4643 39904
rect 4709 39882 4739 39904
rect 4805 39882 4835 39904
rect 4901 39882 4931 39904
rect 3971 39862 4997 39882
rect 3971 39828 3987 39862
rect 4021 39828 4179 39862
rect 4213 39828 4371 39862
rect 4405 39828 4563 39862
rect 4597 39828 4755 39862
rect 4789 39828 4947 39862
rect 4981 39828 4997 39862
rect 3971 39816 4997 39828
rect 5400 39899 5430 39925
rect 297 39379 1323 39395
rect 297 39345 313 39379
rect 347 39345 505 39379
rect 539 39345 697 39379
rect 731 39345 889 39379
rect 923 39345 1081 39379
rect 1115 39345 1273 39379
rect 1307 39345 1323 39379
rect 297 39329 1323 39345
rect 363 39297 393 39329
rect 459 39297 489 39329
rect 555 39297 585 39329
rect 651 39297 681 39329
rect 747 39297 777 39329
rect 843 39297 873 39329
rect 939 39297 969 39329
rect 1035 39297 1065 39329
rect 1131 39297 1161 39329
rect 1227 39297 1257 39329
rect 363 38999 393 39025
rect 459 38999 489 39025
rect 555 38999 585 39025
rect 651 38999 681 39025
rect 747 38999 777 39025
rect 843 38999 873 39025
rect 939 38999 969 39025
rect 1035 38999 1065 39025
rect 1131 38999 1161 39025
rect 1227 38999 1257 39025
rect 2450 39383 3476 39399
rect 2450 39349 2466 39383
rect 2500 39349 2658 39383
rect 2692 39349 2850 39383
rect 2884 39349 3042 39383
rect 3076 39349 3234 39383
rect 3268 39349 3426 39383
rect 3460 39349 3476 39383
rect 2450 39333 3476 39349
rect 2516 39301 2546 39333
rect 2612 39301 2642 39333
rect 2708 39301 2738 39333
rect 2804 39301 2834 39333
rect 2900 39301 2930 39333
rect 2996 39301 3026 39333
rect 3092 39301 3122 39333
rect 3188 39301 3218 39333
rect 3284 39301 3314 39333
rect 3380 39301 3410 39333
rect 2516 39003 2546 39029
rect 2612 39003 2642 39029
rect 2708 39003 2738 39029
rect 2804 39003 2834 39029
rect 2900 39003 2930 39029
rect 2996 39003 3026 39029
rect 3092 39003 3122 39029
rect 3188 39003 3218 39029
rect 3284 39003 3314 39029
rect 3380 39003 3410 39029
rect 3971 39383 4997 39399
rect 3971 39349 3987 39383
rect 4021 39349 4179 39383
rect 4213 39349 4371 39383
rect 4405 39349 4563 39383
rect 4597 39349 4755 39383
rect 4789 39349 4947 39383
rect 4981 39349 4997 39383
rect 3971 39333 4997 39349
rect 4037 39301 4067 39333
rect 4133 39301 4163 39333
rect 4229 39301 4259 39333
rect 4325 39301 4355 39333
rect 4421 39301 4451 39333
rect 4517 39301 4547 39333
rect 4613 39301 4643 39333
rect 4709 39301 4739 39333
rect 4805 39301 4835 39333
rect 4901 39301 4931 39333
rect 5400 39088 5430 39114
rect 4037 39003 4067 39029
rect 4133 39003 4163 39029
rect 4229 39003 4259 39029
rect 4325 39003 4355 39029
rect 4421 39003 4451 39029
rect 4517 39003 4547 39029
rect 4613 39003 4643 39029
rect 4709 39003 4739 39029
rect 4805 39003 4835 39029
rect 4901 39003 4931 39029
rect 5400 38856 5430 38888
rect 5400 38840 5486 38856
rect 363 38717 393 38743
rect 459 38717 489 38743
rect 555 38717 585 38743
rect 651 38717 681 38743
rect 747 38717 777 38743
rect 843 38717 873 38743
rect 939 38717 969 38743
rect 1035 38717 1065 38743
rect 1131 38717 1161 38743
rect 1227 38717 1257 38743
rect 363 38591 393 38613
rect 459 38591 489 38613
rect 555 38591 585 38613
rect 651 38591 681 38613
rect 747 38591 777 38613
rect 843 38591 873 38613
rect 939 38591 969 38613
rect 1035 38591 1065 38613
rect 1131 38591 1161 38613
rect 1227 38591 1257 38613
rect 297 38571 1323 38591
rect 297 38537 313 38571
rect 347 38537 505 38571
rect 539 38537 697 38571
rect 731 38537 889 38571
rect 923 38537 1081 38571
rect 1115 38537 1273 38571
rect 1307 38537 1323 38571
rect 297 38525 1323 38537
rect 2516 38721 2546 38747
rect 2612 38721 2642 38747
rect 2708 38721 2738 38747
rect 2804 38721 2834 38747
rect 2900 38721 2930 38747
rect 2996 38721 3026 38747
rect 3092 38721 3122 38747
rect 3188 38721 3218 38747
rect 3284 38721 3314 38747
rect 3380 38721 3410 38747
rect 3675 38797 3741 38813
rect 3675 38763 3691 38797
rect 3725 38763 3741 38797
rect 3675 38747 3741 38763
rect 3693 38725 3723 38747
rect 4037 38721 4067 38747
rect 4133 38721 4163 38747
rect 4229 38721 4259 38747
rect 4325 38721 4355 38747
rect 4421 38721 4451 38747
rect 4517 38721 4547 38747
rect 4613 38721 4643 38747
rect 4709 38721 4739 38747
rect 4805 38721 4835 38747
rect 4901 38721 4931 38747
rect 5400 38806 5436 38840
rect 5470 38806 5486 38840
rect 5400 38790 5486 38806
rect 5400 38768 5430 38790
rect 2516 38595 2546 38617
rect 2612 38595 2642 38617
rect 2708 38595 2738 38617
rect 2804 38595 2834 38617
rect 2900 38595 2930 38617
rect 2996 38595 3026 38617
rect 3092 38595 3122 38617
rect 3188 38595 3218 38617
rect 3284 38595 3314 38617
rect 3380 38595 3410 38617
rect 2450 38575 3476 38595
rect 2450 38541 2466 38575
rect 2500 38541 2658 38575
rect 2692 38541 2850 38575
rect 2884 38541 3042 38575
rect 3076 38541 3234 38575
rect 3268 38541 3426 38575
rect 3460 38541 3476 38575
rect 2450 38529 3476 38541
rect 3693 38599 3723 38625
rect 4037 38595 4067 38617
rect 4133 38595 4163 38617
rect 4229 38595 4259 38617
rect 4325 38595 4355 38617
rect 4421 38595 4451 38617
rect 4517 38595 4547 38617
rect 4613 38595 4643 38617
rect 4709 38595 4739 38617
rect 4805 38595 4835 38617
rect 4901 38595 4931 38617
rect 3971 38575 4997 38595
rect 3971 38541 3987 38575
rect 4021 38541 4179 38575
rect 4213 38541 4371 38575
rect 4405 38541 4563 38575
rect 4597 38541 4755 38575
rect 4789 38541 4947 38575
rect 4981 38541 4997 38575
rect 3971 38529 4997 38541
rect 5400 38612 5430 38638
rect 297 38092 1323 38108
rect 297 38058 313 38092
rect 347 38058 505 38092
rect 539 38058 697 38092
rect 731 38058 889 38092
rect 923 38058 1081 38092
rect 1115 38058 1273 38092
rect 1307 38058 1323 38092
rect 297 38042 1323 38058
rect 363 38010 393 38042
rect 459 38010 489 38042
rect 555 38010 585 38042
rect 651 38010 681 38042
rect 747 38010 777 38042
rect 843 38010 873 38042
rect 939 38010 969 38042
rect 1035 38010 1065 38042
rect 1131 38010 1161 38042
rect 1227 38010 1257 38042
rect 363 37712 393 37738
rect 459 37712 489 37738
rect 555 37712 585 37738
rect 651 37712 681 37738
rect 747 37712 777 37738
rect 843 37712 873 37738
rect 939 37712 969 37738
rect 1035 37712 1065 37738
rect 1131 37712 1161 37738
rect 1227 37712 1257 37738
rect 2450 38096 3476 38112
rect 2450 38062 2466 38096
rect 2500 38062 2658 38096
rect 2692 38062 2850 38096
rect 2884 38062 3042 38096
rect 3076 38062 3234 38096
rect 3268 38062 3426 38096
rect 3460 38062 3476 38096
rect 2450 38046 3476 38062
rect 2516 38014 2546 38046
rect 2612 38014 2642 38046
rect 2708 38014 2738 38046
rect 2804 38014 2834 38046
rect 2900 38014 2930 38046
rect 2996 38014 3026 38046
rect 3092 38014 3122 38046
rect 3188 38014 3218 38046
rect 3284 38014 3314 38046
rect 3380 38014 3410 38046
rect 2516 37716 2546 37742
rect 2612 37716 2642 37742
rect 2708 37716 2738 37742
rect 2804 37716 2834 37742
rect 2900 37716 2930 37742
rect 2996 37716 3026 37742
rect 3092 37716 3122 37742
rect 3188 37716 3218 37742
rect 3284 37716 3314 37742
rect 3380 37716 3410 37742
rect 3971 38096 4997 38112
rect 3971 38062 3987 38096
rect 4021 38062 4179 38096
rect 4213 38062 4371 38096
rect 4405 38062 4563 38096
rect 4597 38062 4755 38096
rect 4789 38062 4947 38096
rect 4981 38062 4997 38096
rect 3971 38046 4997 38062
rect 4037 38014 4067 38046
rect 4133 38014 4163 38046
rect 4229 38014 4259 38046
rect 4325 38014 4355 38046
rect 4421 38014 4451 38046
rect 4517 38014 4547 38046
rect 4613 38014 4643 38046
rect 4709 38014 4739 38046
rect 4805 38014 4835 38046
rect 4901 38014 4931 38046
rect 5400 37801 5430 37827
rect 4037 37716 4067 37742
rect 4133 37716 4163 37742
rect 4229 37716 4259 37742
rect 4325 37716 4355 37742
rect 4421 37716 4451 37742
rect 4517 37716 4547 37742
rect 4613 37716 4643 37742
rect 4709 37716 4739 37742
rect 4805 37716 4835 37742
rect 4901 37716 4931 37742
rect 5400 37569 5430 37601
rect 5400 37553 5486 37569
rect 363 37430 393 37456
rect 459 37430 489 37456
rect 555 37430 585 37456
rect 651 37430 681 37456
rect 747 37430 777 37456
rect 843 37430 873 37456
rect 939 37430 969 37456
rect 1035 37430 1065 37456
rect 1131 37430 1161 37456
rect 1227 37430 1257 37456
rect 363 37304 393 37326
rect 459 37304 489 37326
rect 555 37304 585 37326
rect 651 37304 681 37326
rect 747 37304 777 37326
rect 843 37304 873 37326
rect 939 37304 969 37326
rect 1035 37304 1065 37326
rect 1131 37304 1161 37326
rect 1227 37304 1257 37326
rect 297 37284 1323 37304
rect 297 37250 313 37284
rect 347 37250 505 37284
rect 539 37250 697 37284
rect 731 37250 889 37284
rect 923 37250 1081 37284
rect 1115 37250 1273 37284
rect 1307 37250 1323 37284
rect 297 37238 1323 37250
rect 2516 37434 2546 37460
rect 2612 37434 2642 37460
rect 2708 37434 2738 37460
rect 2804 37434 2834 37460
rect 2900 37434 2930 37460
rect 2996 37434 3026 37460
rect 3092 37434 3122 37460
rect 3188 37434 3218 37460
rect 3284 37434 3314 37460
rect 3380 37434 3410 37460
rect 3675 37510 3741 37526
rect 3675 37476 3691 37510
rect 3725 37476 3741 37510
rect 3675 37460 3741 37476
rect 3693 37438 3723 37460
rect 4037 37434 4067 37460
rect 4133 37434 4163 37460
rect 4229 37434 4259 37460
rect 4325 37434 4355 37460
rect 4421 37434 4451 37460
rect 4517 37434 4547 37460
rect 4613 37434 4643 37460
rect 4709 37434 4739 37460
rect 4805 37434 4835 37460
rect 4901 37434 4931 37460
rect 5400 37519 5436 37553
rect 5470 37519 5486 37553
rect 5400 37503 5486 37519
rect 5400 37481 5430 37503
rect 2516 37308 2546 37330
rect 2612 37308 2642 37330
rect 2708 37308 2738 37330
rect 2804 37308 2834 37330
rect 2900 37308 2930 37330
rect 2996 37308 3026 37330
rect 3092 37308 3122 37330
rect 3188 37308 3218 37330
rect 3284 37308 3314 37330
rect 3380 37308 3410 37330
rect 2450 37288 3476 37308
rect 2450 37254 2466 37288
rect 2500 37254 2658 37288
rect 2692 37254 2850 37288
rect 2884 37254 3042 37288
rect 3076 37254 3234 37288
rect 3268 37254 3426 37288
rect 3460 37254 3476 37288
rect 2450 37242 3476 37254
rect 3693 37312 3723 37338
rect 4037 37308 4067 37330
rect 4133 37308 4163 37330
rect 4229 37308 4259 37330
rect 4325 37308 4355 37330
rect 4421 37308 4451 37330
rect 4517 37308 4547 37330
rect 4613 37308 4643 37330
rect 4709 37308 4739 37330
rect 4805 37308 4835 37330
rect 4901 37308 4931 37330
rect 3971 37288 4997 37308
rect 3971 37254 3987 37288
rect 4021 37254 4179 37288
rect 4213 37254 4371 37288
rect 4405 37254 4563 37288
rect 4597 37254 4755 37288
rect 4789 37254 4947 37288
rect 4981 37254 4997 37288
rect 3971 37242 4997 37254
rect 5400 37325 5430 37351
rect 297 36805 1323 36821
rect 297 36771 313 36805
rect 347 36771 505 36805
rect 539 36771 697 36805
rect 731 36771 889 36805
rect 923 36771 1081 36805
rect 1115 36771 1273 36805
rect 1307 36771 1323 36805
rect 297 36755 1323 36771
rect 363 36723 393 36755
rect 459 36723 489 36755
rect 555 36723 585 36755
rect 651 36723 681 36755
rect 747 36723 777 36755
rect 843 36723 873 36755
rect 939 36723 969 36755
rect 1035 36723 1065 36755
rect 1131 36723 1161 36755
rect 1227 36723 1257 36755
rect 363 36425 393 36451
rect 459 36425 489 36451
rect 555 36425 585 36451
rect 651 36425 681 36451
rect 747 36425 777 36451
rect 843 36425 873 36451
rect 939 36425 969 36451
rect 1035 36425 1065 36451
rect 1131 36425 1161 36451
rect 1227 36425 1257 36451
rect 2450 36809 3476 36825
rect 2450 36775 2466 36809
rect 2500 36775 2658 36809
rect 2692 36775 2850 36809
rect 2884 36775 3042 36809
rect 3076 36775 3234 36809
rect 3268 36775 3426 36809
rect 3460 36775 3476 36809
rect 2450 36759 3476 36775
rect 2516 36727 2546 36759
rect 2612 36727 2642 36759
rect 2708 36727 2738 36759
rect 2804 36727 2834 36759
rect 2900 36727 2930 36759
rect 2996 36727 3026 36759
rect 3092 36727 3122 36759
rect 3188 36727 3218 36759
rect 3284 36727 3314 36759
rect 3380 36727 3410 36759
rect 2516 36429 2546 36455
rect 2612 36429 2642 36455
rect 2708 36429 2738 36455
rect 2804 36429 2834 36455
rect 2900 36429 2930 36455
rect 2996 36429 3026 36455
rect 3092 36429 3122 36455
rect 3188 36429 3218 36455
rect 3284 36429 3314 36455
rect 3380 36429 3410 36455
rect 3971 36809 4997 36825
rect 3971 36775 3987 36809
rect 4021 36775 4179 36809
rect 4213 36775 4371 36809
rect 4405 36775 4563 36809
rect 4597 36775 4755 36809
rect 4789 36775 4947 36809
rect 4981 36775 4997 36809
rect 3971 36759 4997 36775
rect 4037 36727 4067 36759
rect 4133 36727 4163 36759
rect 4229 36727 4259 36759
rect 4325 36727 4355 36759
rect 4421 36727 4451 36759
rect 4517 36727 4547 36759
rect 4613 36727 4643 36759
rect 4709 36727 4739 36759
rect 4805 36727 4835 36759
rect 4901 36727 4931 36759
rect 5400 36514 5430 36540
rect 4037 36429 4067 36455
rect 4133 36429 4163 36455
rect 4229 36429 4259 36455
rect 4325 36429 4355 36455
rect 4421 36429 4451 36455
rect 4517 36429 4547 36455
rect 4613 36429 4643 36455
rect 4709 36429 4739 36455
rect 4805 36429 4835 36455
rect 4901 36429 4931 36455
rect 5400 36282 5430 36314
rect 5400 36266 5486 36282
rect 363 36143 393 36169
rect 459 36143 489 36169
rect 555 36143 585 36169
rect 651 36143 681 36169
rect 747 36143 777 36169
rect 843 36143 873 36169
rect 939 36143 969 36169
rect 1035 36143 1065 36169
rect 1131 36143 1161 36169
rect 1227 36143 1257 36169
rect 363 36017 393 36039
rect 459 36017 489 36039
rect 555 36017 585 36039
rect 651 36017 681 36039
rect 747 36017 777 36039
rect 843 36017 873 36039
rect 939 36017 969 36039
rect 1035 36017 1065 36039
rect 1131 36017 1161 36039
rect 1227 36017 1257 36039
rect 297 35997 1323 36017
rect 297 35963 313 35997
rect 347 35963 505 35997
rect 539 35963 697 35997
rect 731 35963 889 35997
rect 923 35963 1081 35997
rect 1115 35963 1273 35997
rect 1307 35963 1323 35997
rect 297 35951 1323 35963
rect 2516 36147 2546 36173
rect 2612 36147 2642 36173
rect 2708 36147 2738 36173
rect 2804 36147 2834 36173
rect 2900 36147 2930 36173
rect 2996 36147 3026 36173
rect 3092 36147 3122 36173
rect 3188 36147 3218 36173
rect 3284 36147 3314 36173
rect 3380 36147 3410 36173
rect 3675 36223 3741 36239
rect 3675 36189 3691 36223
rect 3725 36189 3741 36223
rect 3675 36173 3741 36189
rect 3693 36151 3723 36173
rect 4037 36147 4067 36173
rect 4133 36147 4163 36173
rect 4229 36147 4259 36173
rect 4325 36147 4355 36173
rect 4421 36147 4451 36173
rect 4517 36147 4547 36173
rect 4613 36147 4643 36173
rect 4709 36147 4739 36173
rect 4805 36147 4835 36173
rect 4901 36147 4931 36173
rect 5400 36232 5436 36266
rect 5470 36232 5486 36266
rect 5400 36216 5486 36232
rect 5400 36194 5430 36216
rect 2516 36021 2546 36043
rect 2612 36021 2642 36043
rect 2708 36021 2738 36043
rect 2804 36021 2834 36043
rect 2900 36021 2930 36043
rect 2996 36021 3026 36043
rect 3092 36021 3122 36043
rect 3188 36021 3218 36043
rect 3284 36021 3314 36043
rect 3380 36021 3410 36043
rect 2450 36001 3476 36021
rect 2450 35967 2466 36001
rect 2500 35967 2658 36001
rect 2692 35967 2850 36001
rect 2884 35967 3042 36001
rect 3076 35967 3234 36001
rect 3268 35967 3426 36001
rect 3460 35967 3476 36001
rect 2450 35955 3476 35967
rect 3693 36025 3723 36051
rect 4037 36021 4067 36043
rect 4133 36021 4163 36043
rect 4229 36021 4259 36043
rect 4325 36021 4355 36043
rect 4421 36021 4451 36043
rect 4517 36021 4547 36043
rect 4613 36021 4643 36043
rect 4709 36021 4739 36043
rect 4805 36021 4835 36043
rect 4901 36021 4931 36043
rect 3971 36001 4997 36021
rect 3971 35967 3987 36001
rect 4021 35967 4179 36001
rect 4213 35967 4371 36001
rect 4405 35967 4563 36001
rect 4597 35967 4755 36001
rect 4789 35967 4947 36001
rect 4981 35967 4997 36001
rect 3971 35955 4997 35967
rect 5400 36038 5430 36064
rect 297 35518 1323 35534
rect 297 35484 313 35518
rect 347 35484 505 35518
rect 539 35484 697 35518
rect 731 35484 889 35518
rect 923 35484 1081 35518
rect 1115 35484 1273 35518
rect 1307 35484 1323 35518
rect 297 35468 1323 35484
rect 363 35436 393 35468
rect 459 35436 489 35468
rect 555 35436 585 35468
rect 651 35436 681 35468
rect 747 35436 777 35468
rect 843 35436 873 35468
rect 939 35436 969 35468
rect 1035 35436 1065 35468
rect 1131 35436 1161 35468
rect 1227 35436 1257 35468
rect 363 35138 393 35164
rect 459 35138 489 35164
rect 555 35138 585 35164
rect 651 35138 681 35164
rect 747 35138 777 35164
rect 843 35138 873 35164
rect 939 35138 969 35164
rect 1035 35138 1065 35164
rect 1131 35138 1161 35164
rect 1227 35138 1257 35164
rect 2450 35522 3476 35538
rect 2450 35488 2466 35522
rect 2500 35488 2658 35522
rect 2692 35488 2850 35522
rect 2884 35488 3042 35522
rect 3076 35488 3234 35522
rect 3268 35488 3426 35522
rect 3460 35488 3476 35522
rect 2450 35472 3476 35488
rect 2516 35440 2546 35472
rect 2612 35440 2642 35472
rect 2708 35440 2738 35472
rect 2804 35440 2834 35472
rect 2900 35440 2930 35472
rect 2996 35440 3026 35472
rect 3092 35440 3122 35472
rect 3188 35440 3218 35472
rect 3284 35440 3314 35472
rect 3380 35440 3410 35472
rect 2516 35142 2546 35168
rect 2612 35142 2642 35168
rect 2708 35142 2738 35168
rect 2804 35142 2834 35168
rect 2900 35142 2930 35168
rect 2996 35142 3026 35168
rect 3092 35142 3122 35168
rect 3188 35142 3218 35168
rect 3284 35142 3314 35168
rect 3380 35142 3410 35168
rect 3971 35522 4997 35538
rect 3971 35488 3987 35522
rect 4021 35488 4179 35522
rect 4213 35488 4371 35522
rect 4405 35488 4563 35522
rect 4597 35488 4755 35522
rect 4789 35488 4947 35522
rect 4981 35488 4997 35522
rect 3971 35472 4997 35488
rect 4037 35440 4067 35472
rect 4133 35440 4163 35472
rect 4229 35440 4259 35472
rect 4325 35440 4355 35472
rect 4421 35440 4451 35472
rect 4517 35440 4547 35472
rect 4613 35440 4643 35472
rect 4709 35440 4739 35472
rect 4805 35440 4835 35472
rect 4901 35440 4931 35472
rect 5400 35227 5430 35253
rect 4037 35142 4067 35168
rect 4133 35142 4163 35168
rect 4229 35142 4259 35168
rect 4325 35142 4355 35168
rect 4421 35142 4451 35168
rect 4517 35142 4547 35168
rect 4613 35142 4643 35168
rect 4709 35142 4739 35168
rect 4805 35142 4835 35168
rect 4901 35142 4931 35168
rect 5400 34995 5430 35027
rect 5400 34979 5486 34995
rect 363 34856 393 34882
rect 459 34856 489 34882
rect 555 34856 585 34882
rect 651 34856 681 34882
rect 747 34856 777 34882
rect 843 34856 873 34882
rect 939 34856 969 34882
rect 1035 34856 1065 34882
rect 1131 34856 1161 34882
rect 1227 34856 1257 34882
rect 363 34730 393 34752
rect 459 34730 489 34752
rect 555 34730 585 34752
rect 651 34730 681 34752
rect 747 34730 777 34752
rect 843 34730 873 34752
rect 939 34730 969 34752
rect 1035 34730 1065 34752
rect 1131 34730 1161 34752
rect 1227 34730 1257 34752
rect 297 34710 1323 34730
rect 297 34676 313 34710
rect 347 34676 505 34710
rect 539 34676 697 34710
rect 731 34676 889 34710
rect 923 34676 1081 34710
rect 1115 34676 1273 34710
rect 1307 34676 1323 34710
rect 297 34664 1323 34676
rect 2516 34860 2546 34886
rect 2612 34860 2642 34886
rect 2708 34860 2738 34886
rect 2804 34860 2834 34886
rect 2900 34860 2930 34886
rect 2996 34860 3026 34886
rect 3092 34860 3122 34886
rect 3188 34860 3218 34886
rect 3284 34860 3314 34886
rect 3380 34860 3410 34886
rect 3675 34936 3741 34952
rect 3675 34902 3691 34936
rect 3725 34902 3741 34936
rect 3675 34886 3741 34902
rect 3693 34864 3723 34886
rect 4037 34860 4067 34886
rect 4133 34860 4163 34886
rect 4229 34860 4259 34886
rect 4325 34860 4355 34886
rect 4421 34860 4451 34886
rect 4517 34860 4547 34886
rect 4613 34860 4643 34886
rect 4709 34860 4739 34886
rect 4805 34860 4835 34886
rect 4901 34860 4931 34886
rect 5400 34945 5436 34979
rect 5470 34945 5486 34979
rect 5400 34929 5486 34945
rect 5400 34907 5430 34929
rect 2516 34734 2546 34756
rect 2612 34734 2642 34756
rect 2708 34734 2738 34756
rect 2804 34734 2834 34756
rect 2900 34734 2930 34756
rect 2996 34734 3026 34756
rect 3092 34734 3122 34756
rect 3188 34734 3218 34756
rect 3284 34734 3314 34756
rect 3380 34734 3410 34756
rect 2450 34714 3476 34734
rect 2450 34680 2466 34714
rect 2500 34680 2658 34714
rect 2692 34680 2850 34714
rect 2884 34680 3042 34714
rect 3076 34680 3234 34714
rect 3268 34680 3426 34714
rect 3460 34680 3476 34714
rect 2450 34668 3476 34680
rect 3693 34738 3723 34764
rect 4037 34734 4067 34756
rect 4133 34734 4163 34756
rect 4229 34734 4259 34756
rect 4325 34734 4355 34756
rect 4421 34734 4451 34756
rect 4517 34734 4547 34756
rect 4613 34734 4643 34756
rect 4709 34734 4739 34756
rect 4805 34734 4835 34756
rect 4901 34734 4931 34756
rect 3971 34714 4997 34734
rect 3971 34680 3987 34714
rect 4021 34680 4179 34714
rect 4213 34680 4371 34714
rect 4405 34680 4563 34714
rect 4597 34680 4755 34714
rect 4789 34680 4947 34714
rect 4981 34680 4997 34714
rect 3971 34668 4997 34680
rect 5400 34751 5430 34777
rect 297 34231 1323 34247
rect 297 34197 313 34231
rect 347 34197 505 34231
rect 539 34197 697 34231
rect 731 34197 889 34231
rect 923 34197 1081 34231
rect 1115 34197 1273 34231
rect 1307 34197 1323 34231
rect 297 34181 1323 34197
rect 363 34149 393 34181
rect 459 34149 489 34181
rect 555 34149 585 34181
rect 651 34149 681 34181
rect 747 34149 777 34181
rect 843 34149 873 34181
rect 939 34149 969 34181
rect 1035 34149 1065 34181
rect 1131 34149 1161 34181
rect 1227 34149 1257 34181
rect 363 33851 393 33877
rect 459 33851 489 33877
rect 555 33851 585 33877
rect 651 33851 681 33877
rect 747 33851 777 33877
rect 843 33851 873 33877
rect 939 33851 969 33877
rect 1035 33851 1065 33877
rect 1131 33851 1161 33877
rect 1227 33851 1257 33877
rect 2450 34235 3476 34251
rect 2450 34201 2466 34235
rect 2500 34201 2658 34235
rect 2692 34201 2850 34235
rect 2884 34201 3042 34235
rect 3076 34201 3234 34235
rect 3268 34201 3426 34235
rect 3460 34201 3476 34235
rect 2450 34185 3476 34201
rect 2516 34153 2546 34185
rect 2612 34153 2642 34185
rect 2708 34153 2738 34185
rect 2804 34153 2834 34185
rect 2900 34153 2930 34185
rect 2996 34153 3026 34185
rect 3092 34153 3122 34185
rect 3188 34153 3218 34185
rect 3284 34153 3314 34185
rect 3380 34153 3410 34185
rect 2516 33855 2546 33881
rect 2612 33855 2642 33881
rect 2708 33855 2738 33881
rect 2804 33855 2834 33881
rect 2900 33855 2930 33881
rect 2996 33855 3026 33881
rect 3092 33855 3122 33881
rect 3188 33855 3218 33881
rect 3284 33855 3314 33881
rect 3380 33855 3410 33881
rect 3971 34235 4997 34251
rect 3971 34201 3987 34235
rect 4021 34201 4179 34235
rect 4213 34201 4371 34235
rect 4405 34201 4563 34235
rect 4597 34201 4755 34235
rect 4789 34201 4947 34235
rect 4981 34201 4997 34235
rect 3971 34185 4997 34201
rect 4037 34153 4067 34185
rect 4133 34153 4163 34185
rect 4229 34153 4259 34185
rect 4325 34153 4355 34185
rect 4421 34153 4451 34185
rect 4517 34153 4547 34185
rect 4613 34153 4643 34185
rect 4709 34153 4739 34185
rect 4805 34153 4835 34185
rect 4901 34153 4931 34185
rect 5400 33940 5430 33966
rect 4037 33855 4067 33881
rect 4133 33855 4163 33881
rect 4229 33855 4259 33881
rect 4325 33855 4355 33881
rect 4421 33855 4451 33881
rect 4517 33855 4547 33881
rect 4613 33855 4643 33881
rect 4709 33855 4739 33881
rect 4805 33855 4835 33881
rect 4901 33855 4931 33881
rect 5400 33708 5430 33740
rect 5400 33692 5486 33708
rect 363 33569 393 33595
rect 459 33569 489 33595
rect 555 33569 585 33595
rect 651 33569 681 33595
rect 747 33569 777 33595
rect 843 33569 873 33595
rect 939 33569 969 33595
rect 1035 33569 1065 33595
rect 1131 33569 1161 33595
rect 1227 33569 1257 33595
rect 363 33443 393 33465
rect 459 33443 489 33465
rect 555 33443 585 33465
rect 651 33443 681 33465
rect 747 33443 777 33465
rect 843 33443 873 33465
rect 939 33443 969 33465
rect 1035 33443 1065 33465
rect 1131 33443 1161 33465
rect 1227 33443 1257 33465
rect 297 33423 1323 33443
rect 297 33389 313 33423
rect 347 33389 505 33423
rect 539 33389 697 33423
rect 731 33389 889 33423
rect 923 33389 1081 33423
rect 1115 33389 1273 33423
rect 1307 33389 1323 33423
rect 297 33377 1323 33389
rect 2516 33573 2546 33599
rect 2612 33573 2642 33599
rect 2708 33573 2738 33599
rect 2804 33573 2834 33599
rect 2900 33573 2930 33599
rect 2996 33573 3026 33599
rect 3092 33573 3122 33599
rect 3188 33573 3218 33599
rect 3284 33573 3314 33599
rect 3380 33573 3410 33599
rect 3675 33649 3741 33665
rect 3675 33615 3691 33649
rect 3725 33615 3741 33649
rect 3675 33599 3741 33615
rect 3693 33577 3723 33599
rect 4037 33573 4067 33599
rect 4133 33573 4163 33599
rect 4229 33573 4259 33599
rect 4325 33573 4355 33599
rect 4421 33573 4451 33599
rect 4517 33573 4547 33599
rect 4613 33573 4643 33599
rect 4709 33573 4739 33599
rect 4805 33573 4835 33599
rect 4901 33573 4931 33599
rect 5400 33658 5436 33692
rect 5470 33658 5486 33692
rect 5400 33642 5486 33658
rect 5400 33620 5430 33642
rect 2516 33447 2546 33469
rect 2612 33447 2642 33469
rect 2708 33447 2738 33469
rect 2804 33447 2834 33469
rect 2900 33447 2930 33469
rect 2996 33447 3026 33469
rect 3092 33447 3122 33469
rect 3188 33447 3218 33469
rect 3284 33447 3314 33469
rect 3380 33447 3410 33469
rect 2450 33427 3476 33447
rect 2450 33393 2466 33427
rect 2500 33393 2658 33427
rect 2692 33393 2850 33427
rect 2884 33393 3042 33427
rect 3076 33393 3234 33427
rect 3268 33393 3426 33427
rect 3460 33393 3476 33427
rect 2450 33381 3476 33393
rect 3693 33451 3723 33477
rect 4037 33447 4067 33469
rect 4133 33447 4163 33469
rect 4229 33447 4259 33469
rect 4325 33447 4355 33469
rect 4421 33447 4451 33469
rect 4517 33447 4547 33469
rect 4613 33447 4643 33469
rect 4709 33447 4739 33469
rect 4805 33447 4835 33469
rect 4901 33447 4931 33469
rect 3971 33427 4997 33447
rect 3971 33393 3987 33427
rect 4021 33393 4179 33427
rect 4213 33393 4371 33427
rect 4405 33393 4563 33427
rect 4597 33393 4755 33427
rect 4789 33393 4947 33427
rect 4981 33393 4997 33427
rect 3971 33381 4997 33393
rect 5400 33464 5430 33490
rect 297 32944 1323 32960
rect 297 32910 313 32944
rect 347 32910 505 32944
rect 539 32910 697 32944
rect 731 32910 889 32944
rect 923 32910 1081 32944
rect 1115 32910 1273 32944
rect 1307 32910 1323 32944
rect 297 32894 1323 32910
rect 363 32862 393 32894
rect 459 32862 489 32894
rect 555 32862 585 32894
rect 651 32862 681 32894
rect 747 32862 777 32894
rect 843 32862 873 32894
rect 939 32862 969 32894
rect 1035 32862 1065 32894
rect 1131 32862 1161 32894
rect 1227 32862 1257 32894
rect 363 32564 393 32590
rect 459 32564 489 32590
rect 555 32564 585 32590
rect 651 32564 681 32590
rect 747 32564 777 32590
rect 843 32564 873 32590
rect 939 32564 969 32590
rect 1035 32564 1065 32590
rect 1131 32564 1161 32590
rect 1227 32564 1257 32590
rect 2450 32948 3476 32964
rect 2450 32914 2466 32948
rect 2500 32914 2658 32948
rect 2692 32914 2850 32948
rect 2884 32914 3042 32948
rect 3076 32914 3234 32948
rect 3268 32914 3426 32948
rect 3460 32914 3476 32948
rect 2450 32898 3476 32914
rect 2516 32866 2546 32898
rect 2612 32866 2642 32898
rect 2708 32866 2738 32898
rect 2804 32866 2834 32898
rect 2900 32866 2930 32898
rect 2996 32866 3026 32898
rect 3092 32866 3122 32898
rect 3188 32866 3218 32898
rect 3284 32866 3314 32898
rect 3380 32866 3410 32898
rect 2516 32568 2546 32594
rect 2612 32568 2642 32594
rect 2708 32568 2738 32594
rect 2804 32568 2834 32594
rect 2900 32568 2930 32594
rect 2996 32568 3026 32594
rect 3092 32568 3122 32594
rect 3188 32568 3218 32594
rect 3284 32568 3314 32594
rect 3380 32568 3410 32594
rect 3971 32948 4997 32964
rect 3971 32914 3987 32948
rect 4021 32914 4179 32948
rect 4213 32914 4371 32948
rect 4405 32914 4563 32948
rect 4597 32914 4755 32948
rect 4789 32914 4947 32948
rect 4981 32914 4997 32948
rect 3971 32898 4997 32914
rect 4037 32866 4067 32898
rect 4133 32866 4163 32898
rect 4229 32866 4259 32898
rect 4325 32866 4355 32898
rect 4421 32866 4451 32898
rect 4517 32866 4547 32898
rect 4613 32866 4643 32898
rect 4709 32866 4739 32898
rect 4805 32866 4835 32898
rect 4901 32866 4931 32898
rect 5400 32653 5430 32679
rect 4037 32568 4067 32594
rect 4133 32568 4163 32594
rect 4229 32568 4259 32594
rect 4325 32568 4355 32594
rect 4421 32568 4451 32594
rect 4517 32568 4547 32594
rect 4613 32568 4643 32594
rect 4709 32568 4739 32594
rect 4805 32568 4835 32594
rect 4901 32568 4931 32594
rect 5400 32421 5430 32453
rect 5400 32405 5486 32421
rect 363 32282 393 32308
rect 459 32282 489 32308
rect 555 32282 585 32308
rect 651 32282 681 32308
rect 747 32282 777 32308
rect 843 32282 873 32308
rect 939 32282 969 32308
rect 1035 32282 1065 32308
rect 1131 32282 1161 32308
rect 1227 32282 1257 32308
rect 363 32156 393 32178
rect 459 32156 489 32178
rect 555 32156 585 32178
rect 651 32156 681 32178
rect 747 32156 777 32178
rect 843 32156 873 32178
rect 939 32156 969 32178
rect 1035 32156 1065 32178
rect 1131 32156 1161 32178
rect 1227 32156 1257 32178
rect 297 32136 1323 32156
rect 297 32102 313 32136
rect 347 32102 505 32136
rect 539 32102 697 32136
rect 731 32102 889 32136
rect 923 32102 1081 32136
rect 1115 32102 1273 32136
rect 1307 32102 1323 32136
rect 297 32090 1323 32102
rect 2516 32286 2546 32312
rect 2612 32286 2642 32312
rect 2708 32286 2738 32312
rect 2804 32286 2834 32312
rect 2900 32286 2930 32312
rect 2996 32286 3026 32312
rect 3092 32286 3122 32312
rect 3188 32286 3218 32312
rect 3284 32286 3314 32312
rect 3380 32286 3410 32312
rect 3675 32362 3741 32378
rect 3675 32328 3691 32362
rect 3725 32328 3741 32362
rect 3675 32312 3741 32328
rect 3693 32290 3723 32312
rect 4037 32286 4067 32312
rect 4133 32286 4163 32312
rect 4229 32286 4259 32312
rect 4325 32286 4355 32312
rect 4421 32286 4451 32312
rect 4517 32286 4547 32312
rect 4613 32286 4643 32312
rect 4709 32286 4739 32312
rect 4805 32286 4835 32312
rect 4901 32286 4931 32312
rect 5400 32371 5436 32405
rect 5470 32371 5486 32405
rect 5400 32355 5486 32371
rect 5400 32333 5430 32355
rect 2516 32160 2546 32182
rect 2612 32160 2642 32182
rect 2708 32160 2738 32182
rect 2804 32160 2834 32182
rect 2900 32160 2930 32182
rect 2996 32160 3026 32182
rect 3092 32160 3122 32182
rect 3188 32160 3218 32182
rect 3284 32160 3314 32182
rect 3380 32160 3410 32182
rect 2450 32140 3476 32160
rect 2450 32106 2466 32140
rect 2500 32106 2658 32140
rect 2692 32106 2850 32140
rect 2884 32106 3042 32140
rect 3076 32106 3234 32140
rect 3268 32106 3426 32140
rect 3460 32106 3476 32140
rect 2450 32094 3476 32106
rect 3693 32164 3723 32190
rect 4037 32160 4067 32182
rect 4133 32160 4163 32182
rect 4229 32160 4259 32182
rect 4325 32160 4355 32182
rect 4421 32160 4451 32182
rect 4517 32160 4547 32182
rect 4613 32160 4643 32182
rect 4709 32160 4739 32182
rect 4805 32160 4835 32182
rect 4901 32160 4931 32182
rect 3971 32140 4997 32160
rect 3971 32106 3987 32140
rect 4021 32106 4179 32140
rect 4213 32106 4371 32140
rect 4405 32106 4563 32140
rect 4597 32106 4755 32140
rect 4789 32106 4947 32140
rect 4981 32106 4997 32140
rect 3971 32094 4997 32106
rect 5400 32177 5430 32203
rect 297 31657 1323 31673
rect 297 31623 313 31657
rect 347 31623 505 31657
rect 539 31623 697 31657
rect 731 31623 889 31657
rect 923 31623 1081 31657
rect 1115 31623 1273 31657
rect 1307 31623 1323 31657
rect 297 31607 1323 31623
rect 363 31575 393 31607
rect 459 31575 489 31607
rect 555 31575 585 31607
rect 651 31575 681 31607
rect 747 31575 777 31607
rect 843 31575 873 31607
rect 939 31575 969 31607
rect 1035 31575 1065 31607
rect 1131 31575 1161 31607
rect 1227 31575 1257 31607
rect 363 31277 393 31303
rect 459 31277 489 31303
rect 555 31277 585 31303
rect 651 31277 681 31303
rect 747 31277 777 31303
rect 843 31277 873 31303
rect 939 31277 969 31303
rect 1035 31277 1065 31303
rect 1131 31277 1161 31303
rect 1227 31277 1257 31303
rect 2450 31661 3476 31677
rect 2450 31627 2466 31661
rect 2500 31627 2658 31661
rect 2692 31627 2850 31661
rect 2884 31627 3042 31661
rect 3076 31627 3234 31661
rect 3268 31627 3426 31661
rect 3460 31627 3476 31661
rect 2450 31611 3476 31627
rect 2516 31579 2546 31611
rect 2612 31579 2642 31611
rect 2708 31579 2738 31611
rect 2804 31579 2834 31611
rect 2900 31579 2930 31611
rect 2996 31579 3026 31611
rect 3092 31579 3122 31611
rect 3188 31579 3218 31611
rect 3284 31579 3314 31611
rect 3380 31579 3410 31611
rect 2516 31281 2546 31307
rect 2612 31281 2642 31307
rect 2708 31281 2738 31307
rect 2804 31281 2834 31307
rect 2900 31281 2930 31307
rect 2996 31281 3026 31307
rect 3092 31281 3122 31307
rect 3188 31281 3218 31307
rect 3284 31281 3314 31307
rect 3380 31281 3410 31307
rect 3971 31661 4997 31677
rect 3971 31627 3987 31661
rect 4021 31627 4179 31661
rect 4213 31627 4371 31661
rect 4405 31627 4563 31661
rect 4597 31627 4755 31661
rect 4789 31627 4947 31661
rect 4981 31627 4997 31661
rect 3971 31611 4997 31627
rect 4037 31579 4067 31611
rect 4133 31579 4163 31611
rect 4229 31579 4259 31611
rect 4325 31579 4355 31611
rect 4421 31579 4451 31611
rect 4517 31579 4547 31611
rect 4613 31579 4643 31611
rect 4709 31579 4739 31611
rect 4805 31579 4835 31611
rect 4901 31579 4931 31611
rect 5400 31366 5430 31392
rect 4037 31281 4067 31307
rect 4133 31281 4163 31307
rect 4229 31281 4259 31307
rect 4325 31281 4355 31307
rect 4421 31281 4451 31307
rect 4517 31281 4547 31307
rect 4613 31281 4643 31307
rect 4709 31281 4739 31307
rect 4805 31281 4835 31307
rect 4901 31281 4931 31307
rect 5400 31134 5430 31166
rect 5400 31118 5486 31134
rect 363 30995 393 31021
rect 459 30995 489 31021
rect 555 30995 585 31021
rect 651 30995 681 31021
rect 747 30995 777 31021
rect 843 30995 873 31021
rect 939 30995 969 31021
rect 1035 30995 1065 31021
rect 1131 30995 1161 31021
rect 1227 30995 1257 31021
rect 363 30869 393 30891
rect 459 30869 489 30891
rect 555 30869 585 30891
rect 651 30869 681 30891
rect 747 30869 777 30891
rect 843 30869 873 30891
rect 939 30869 969 30891
rect 1035 30869 1065 30891
rect 1131 30869 1161 30891
rect 1227 30869 1257 30891
rect 297 30849 1323 30869
rect 297 30815 313 30849
rect 347 30815 505 30849
rect 539 30815 697 30849
rect 731 30815 889 30849
rect 923 30815 1081 30849
rect 1115 30815 1273 30849
rect 1307 30815 1323 30849
rect 297 30803 1323 30815
rect 2516 30999 2546 31025
rect 2612 30999 2642 31025
rect 2708 30999 2738 31025
rect 2804 30999 2834 31025
rect 2900 30999 2930 31025
rect 2996 30999 3026 31025
rect 3092 30999 3122 31025
rect 3188 30999 3218 31025
rect 3284 30999 3314 31025
rect 3380 30999 3410 31025
rect 3675 31075 3741 31091
rect 3675 31041 3691 31075
rect 3725 31041 3741 31075
rect 3675 31025 3741 31041
rect 3693 31003 3723 31025
rect 4037 30999 4067 31025
rect 4133 30999 4163 31025
rect 4229 30999 4259 31025
rect 4325 30999 4355 31025
rect 4421 30999 4451 31025
rect 4517 30999 4547 31025
rect 4613 30999 4643 31025
rect 4709 30999 4739 31025
rect 4805 30999 4835 31025
rect 4901 30999 4931 31025
rect 5400 31084 5436 31118
rect 5470 31084 5486 31118
rect 5400 31068 5486 31084
rect 5400 31046 5430 31068
rect 2516 30873 2546 30895
rect 2612 30873 2642 30895
rect 2708 30873 2738 30895
rect 2804 30873 2834 30895
rect 2900 30873 2930 30895
rect 2996 30873 3026 30895
rect 3092 30873 3122 30895
rect 3188 30873 3218 30895
rect 3284 30873 3314 30895
rect 3380 30873 3410 30895
rect 2450 30853 3476 30873
rect 2450 30819 2466 30853
rect 2500 30819 2658 30853
rect 2692 30819 2850 30853
rect 2884 30819 3042 30853
rect 3076 30819 3234 30853
rect 3268 30819 3426 30853
rect 3460 30819 3476 30853
rect 2450 30807 3476 30819
rect 3693 30877 3723 30903
rect 4037 30873 4067 30895
rect 4133 30873 4163 30895
rect 4229 30873 4259 30895
rect 4325 30873 4355 30895
rect 4421 30873 4451 30895
rect 4517 30873 4547 30895
rect 4613 30873 4643 30895
rect 4709 30873 4739 30895
rect 4805 30873 4835 30895
rect 4901 30873 4931 30895
rect 3971 30853 4997 30873
rect 3971 30819 3987 30853
rect 4021 30819 4179 30853
rect 4213 30819 4371 30853
rect 4405 30819 4563 30853
rect 4597 30819 4755 30853
rect 4789 30819 4947 30853
rect 4981 30819 4997 30853
rect 3971 30807 4997 30819
rect 5400 30890 5430 30916
rect 297 30370 1323 30386
rect 297 30336 313 30370
rect 347 30336 505 30370
rect 539 30336 697 30370
rect 731 30336 889 30370
rect 923 30336 1081 30370
rect 1115 30336 1273 30370
rect 1307 30336 1323 30370
rect 297 30320 1323 30336
rect 363 30288 393 30320
rect 459 30288 489 30320
rect 555 30288 585 30320
rect 651 30288 681 30320
rect 747 30288 777 30320
rect 843 30288 873 30320
rect 939 30288 969 30320
rect 1035 30288 1065 30320
rect 1131 30288 1161 30320
rect 1227 30288 1257 30320
rect 363 29990 393 30016
rect 459 29990 489 30016
rect 555 29990 585 30016
rect 651 29990 681 30016
rect 747 29990 777 30016
rect 843 29990 873 30016
rect 939 29990 969 30016
rect 1035 29990 1065 30016
rect 1131 29990 1161 30016
rect 1227 29990 1257 30016
rect 2450 30374 3476 30390
rect 2450 30340 2466 30374
rect 2500 30340 2658 30374
rect 2692 30340 2850 30374
rect 2884 30340 3042 30374
rect 3076 30340 3234 30374
rect 3268 30340 3426 30374
rect 3460 30340 3476 30374
rect 2450 30324 3476 30340
rect 2516 30292 2546 30324
rect 2612 30292 2642 30324
rect 2708 30292 2738 30324
rect 2804 30292 2834 30324
rect 2900 30292 2930 30324
rect 2996 30292 3026 30324
rect 3092 30292 3122 30324
rect 3188 30292 3218 30324
rect 3284 30292 3314 30324
rect 3380 30292 3410 30324
rect 2516 29994 2546 30020
rect 2612 29994 2642 30020
rect 2708 29994 2738 30020
rect 2804 29994 2834 30020
rect 2900 29994 2930 30020
rect 2996 29994 3026 30020
rect 3092 29994 3122 30020
rect 3188 29994 3218 30020
rect 3284 29994 3314 30020
rect 3380 29994 3410 30020
rect 3971 30374 4997 30390
rect 3971 30340 3987 30374
rect 4021 30340 4179 30374
rect 4213 30340 4371 30374
rect 4405 30340 4563 30374
rect 4597 30340 4755 30374
rect 4789 30340 4947 30374
rect 4981 30340 4997 30374
rect 3971 30324 4997 30340
rect 4037 30292 4067 30324
rect 4133 30292 4163 30324
rect 4229 30292 4259 30324
rect 4325 30292 4355 30324
rect 4421 30292 4451 30324
rect 4517 30292 4547 30324
rect 4613 30292 4643 30324
rect 4709 30292 4739 30324
rect 4805 30292 4835 30324
rect 4901 30292 4931 30324
rect 5400 30079 5430 30105
rect 4037 29994 4067 30020
rect 4133 29994 4163 30020
rect 4229 29994 4259 30020
rect 4325 29994 4355 30020
rect 4421 29994 4451 30020
rect 4517 29994 4547 30020
rect 4613 29994 4643 30020
rect 4709 29994 4739 30020
rect 4805 29994 4835 30020
rect 4901 29994 4931 30020
rect 5400 29847 5430 29879
rect 5400 29831 5486 29847
rect 363 29708 393 29734
rect 459 29708 489 29734
rect 555 29708 585 29734
rect 651 29708 681 29734
rect 747 29708 777 29734
rect 843 29708 873 29734
rect 939 29708 969 29734
rect 1035 29708 1065 29734
rect 1131 29708 1161 29734
rect 1227 29708 1257 29734
rect 363 29582 393 29604
rect 459 29582 489 29604
rect 555 29582 585 29604
rect 651 29582 681 29604
rect 747 29582 777 29604
rect 843 29582 873 29604
rect 939 29582 969 29604
rect 1035 29582 1065 29604
rect 1131 29582 1161 29604
rect 1227 29582 1257 29604
rect 297 29562 1323 29582
rect 297 29528 313 29562
rect 347 29528 505 29562
rect 539 29528 697 29562
rect 731 29528 889 29562
rect 923 29528 1081 29562
rect 1115 29528 1273 29562
rect 1307 29528 1323 29562
rect 297 29516 1323 29528
rect 2516 29712 2546 29738
rect 2612 29712 2642 29738
rect 2708 29712 2738 29738
rect 2804 29712 2834 29738
rect 2900 29712 2930 29738
rect 2996 29712 3026 29738
rect 3092 29712 3122 29738
rect 3188 29712 3218 29738
rect 3284 29712 3314 29738
rect 3380 29712 3410 29738
rect 3675 29788 3741 29804
rect 3675 29754 3691 29788
rect 3725 29754 3741 29788
rect 3675 29738 3741 29754
rect 3693 29716 3723 29738
rect 4037 29712 4067 29738
rect 4133 29712 4163 29738
rect 4229 29712 4259 29738
rect 4325 29712 4355 29738
rect 4421 29712 4451 29738
rect 4517 29712 4547 29738
rect 4613 29712 4643 29738
rect 4709 29712 4739 29738
rect 4805 29712 4835 29738
rect 4901 29712 4931 29738
rect 5400 29797 5436 29831
rect 5470 29797 5486 29831
rect 5400 29781 5486 29797
rect 5400 29759 5430 29781
rect 2516 29586 2546 29608
rect 2612 29586 2642 29608
rect 2708 29586 2738 29608
rect 2804 29586 2834 29608
rect 2900 29586 2930 29608
rect 2996 29586 3026 29608
rect 3092 29586 3122 29608
rect 3188 29586 3218 29608
rect 3284 29586 3314 29608
rect 3380 29586 3410 29608
rect 2450 29566 3476 29586
rect 2450 29532 2466 29566
rect 2500 29532 2658 29566
rect 2692 29532 2850 29566
rect 2884 29532 3042 29566
rect 3076 29532 3234 29566
rect 3268 29532 3426 29566
rect 3460 29532 3476 29566
rect 2450 29520 3476 29532
rect 3693 29590 3723 29616
rect 4037 29586 4067 29608
rect 4133 29586 4163 29608
rect 4229 29586 4259 29608
rect 4325 29586 4355 29608
rect 4421 29586 4451 29608
rect 4517 29586 4547 29608
rect 4613 29586 4643 29608
rect 4709 29586 4739 29608
rect 4805 29586 4835 29608
rect 4901 29586 4931 29608
rect 3971 29566 4997 29586
rect 3971 29532 3987 29566
rect 4021 29532 4179 29566
rect 4213 29532 4371 29566
rect 4405 29532 4563 29566
rect 4597 29532 4755 29566
rect 4789 29532 4947 29566
rect 4981 29532 4997 29566
rect 3971 29520 4997 29532
rect 5400 29603 5430 29629
rect 297 29083 1323 29099
rect 297 29049 313 29083
rect 347 29049 505 29083
rect 539 29049 697 29083
rect 731 29049 889 29083
rect 923 29049 1081 29083
rect 1115 29049 1273 29083
rect 1307 29049 1323 29083
rect 297 29033 1323 29049
rect 363 29001 393 29033
rect 459 29001 489 29033
rect 555 29001 585 29033
rect 651 29001 681 29033
rect 747 29001 777 29033
rect 843 29001 873 29033
rect 939 29001 969 29033
rect 1035 29001 1065 29033
rect 1131 29001 1161 29033
rect 1227 29001 1257 29033
rect 363 28703 393 28729
rect 459 28703 489 28729
rect 555 28703 585 28729
rect 651 28703 681 28729
rect 747 28703 777 28729
rect 843 28703 873 28729
rect 939 28703 969 28729
rect 1035 28703 1065 28729
rect 1131 28703 1161 28729
rect 1227 28703 1257 28729
rect 2450 29087 3476 29103
rect 2450 29053 2466 29087
rect 2500 29053 2658 29087
rect 2692 29053 2850 29087
rect 2884 29053 3042 29087
rect 3076 29053 3234 29087
rect 3268 29053 3426 29087
rect 3460 29053 3476 29087
rect 2450 29037 3476 29053
rect 2516 29005 2546 29037
rect 2612 29005 2642 29037
rect 2708 29005 2738 29037
rect 2804 29005 2834 29037
rect 2900 29005 2930 29037
rect 2996 29005 3026 29037
rect 3092 29005 3122 29037
rect 3188 29005 3218 29037
rect 3284 29005 3314 29037
rect 3380 29005 3410 29037
rect 2516 28707 2546 28733
rect 2612 28707 2642 28733
rect 2708 28707 2738 28733
rect 2804 28707 2834 28733
rect 2900 28707 2930 28733
rect 2996 28707 3026 28733
rect 3092 28707 3122 28733
rect 3188 28707 3218 28733
rect 3284 28707 3314 28733
rect 3380 28707 3410 28733
rect 3971 29087 4997 29103
rect 3971 29053 3987 29087
rect 4021 29053 4179 29087
rect 4213 29053 4371 29087
rect 4405 29053 4563 29087
rect 4597 29053 4755 29087
rect 4789 29053 4947 29087
rect 4981 29053 4997 29087
rect 3971 29037 4997 29053
rect 4037 29005 4067 29037
rect 4133 29005 4163 29037
rect 4229 29005 4259 29037
rect 4325 29005 4355 29037
rect 4421 29005 4451 29037
rect 4517 29005 4547 29037
rect 4613 29005 4643 29037
rect 4709 29005 4739 29037
rect 4805 29005 4835 29037
rect 4901 29005 4931 29037
rect 5400 28792 5430 28818
rect 4037 28707 4067 28733
rect 4133 28707 4163 28733
rect 4229 28707 4259 28733
rect 4325 28707 4355 28733
rect 4421 28707 4451 28733
rect 4517 28707 4547 28733
rect 4613 28707 4643 28733
rect 4709 28707 4739 28733
rect 4805 28707 4835 28733
rect 4901 28707 4931 28733
rect 5400 28560 5430 28592
rect 5400 28544 5486 28560
rect 363 28421 393 28447
rect 459 28421 489 28447
rect 555 28421 585 28447
rect 651 28421 681 28447
rect 747 28421 777 28447
rect 843 28421 873 28447
rect 939 28421 969 28447
rect 1035 28421 1065 28447
rect 1131 28421 1161 28447
rect 1227 28421 1257 28447
rect 363 28295 393 28317
rect 459 28295 489 28317
rect 555 28295 585 28317
rect 651 28295 681 28317
rect 747 28295 777 28317
rect 843 28295 873 28317
rect 939 28295 969 28317
rect 1035 28295 1065 28317
rect 1131 28295 1161 28317
rect 1227 28295 1257 28317
rect 297 28275 1323 28295
rect 297 28241 313 28275
rect 347 28241 505 28275
rect 539 28241 697 28275
rect 731 28241 889 28275
rect 923 28241 1081 28275
rect 1115 28241 1273 28275
rect 1307 28241 1323 28275
rect 297 28229 1323 28241
rect 2516 28425 2546 28451
rect 2612 28425 2642 28451
rect 2708 28425 2738 28451
rect 2804 28425 2834 28451
rect 2900 28425 2930 28451
rect 2996 28425 3026 28451
rect 3092 28425 3122 28451
rect 3188 28425 3218 28451
rect 3284 28425 3314 28451
rect 3380 28425 3410 28451
rect 3675 28501 3741 28517
rect 3675 28467 3691 28501
rect 3725 28467 3741 28501
rect 3675 28451 3741 28467
rect 3693 28429 3723 28451
rect 4037 28425 4067 28451
rect 4133 28425 4163 28451
rect 4229 28425 4259 28451
rect 4325 28425 4355 28451
rect 4421 28425 4451 28451
rect 4517 28425 4547 28451
rect 4613 28425 4643 28451
rect 4709 28425 4739 28451
rect 4805 28425 4835 28451
rect 4901 28425 4931 28451
rect 5400 28510 5436 28544
rect 5470 28510 5486 28544
rect 5400 28494 5486 28510
rect 5400 28472 5430 28494
rect 2516 28299 2546 28321
rect 2612 28299 2642 28321
rect 2708 28299 2738 28321
rect 2804 28299 2834 28321
rect 2900 28299 2930 28321
rect 2996 28299 3026 28321
rect 3092 28299 3122 28321
rect 3188 28299 3218 28321
rect 3284 28299 3314 28321
rect 3380 28299 3410 28321
rect 2450 28279 3476 28299
rect 2450 28245 2466 28279
rect 2500 28245 2658 28279
rect 2692 28245 2850 28279
rect 2884 28245 3042 28279
rect 3076 28245 3234 28279
rect 3268 28245 3426 28279
rect 3460 28245 3476 28279
rect 2450 28233 3476 28245
rect 3693 28303 3723 28329
rect 4037 28299 4067 28321
rect 4133 28299 4163 28321
rect 4229 28299 4259 28321
rect 4325 28299 4355 28321
rect 4421 28299 4451 28321
rect 4517 28299 4547 28321
rect 4613 28299 4643 28321
rect 4709 28299 4739 28321
rect 4805 28299 4835 28321
rect 4901 28299 4931 28321
rect 3971 28279 4997 28299
rect 3971 28245 3987 28279
rect 4021 28245 4179 28279
rect 4213 28245 4371 28279
rect 4405 28245 4563 28279
rect 4597 28245 4755 28279
rect 4789 28245 4947 28279
rect 4981 28245 4997 28279
rect 3971 28233 4997 28245
rect 5400 28316 5430 28342
rect 297 27796 1323 27812
rect 297 27762 313 27796
rect 347 27762 505 27796
rect 539 27762 697 27796
rect 731 27762 889 27796
rect 923 27762 1081 27796
rect 1115 27762 1273 27796
rect 1307 27762 1323 27796
rect 297 27746 1323 27762
rect 363 27714 393 27746
rect 459 27714 489 27746
rect 555 27714 585 27746
rect 651 27714 681 27746
rect 747 27714 777 27746
rect 843 27714 873 27746
rect 939 27714 969 27746
rect 1035 27714 1065 27746
rect 1131 27714 1161 27746
rect 1227 27714 1257 27746
rect 363 27416 393 27442
rect 459 27416 489 27442
rect 555 27416 585 27442
rect 651 27416 681 27442
rect 747 27416 777 27442
rect 843 27416 873 27442
rect 939 27416 969 27442
rect 1035 27416 1065 27442
rect 1131 27416 1161 27442
rect 1227 27416 1257 27442
rect 2450 27800 3476 27816
rect 2450 27766 2466 27800
rect 2500 27766 2658 27800
rect 2692 27766 2850 27800
rect 2884 27766 3042 27800
rect 3076 27766 3234 27800
rect 3268 27766 3426 27800
rect 3460 27766 3476 27800
rect 2450 27750 3476 27766
rect 2516 27718 2546 27750
rect 2612 27718 2642 27750
rect 2708 27718 2738 27750
rect 2804 27718 2834 27750
rect 2900 27718 2930 27750
rect 2996 27718 3026 27750
rect 3092 27718 3122 27750
rect 3188 27718 3218 27750
rect 3284 27718 3314 27750
rect 3380 27718 3410 27750
rect 2516 27420 2546 27446
rect 2612 27420 2642 27446
rect 2708 27420 2738 27446
rect 2804 27420 2834 27446
rect 2900 27420 2930 27446
rect 2996 27420 3026 27446
rect 3092 27420 3122 27446
rect 3188 27420 3218 27446
rect 3284 27420 3314 27446
rect 3380 27420 3410 27446
rect 3971 27800 4997 27816
rect 3971 27766 3987 27800
rect 4021 27766 4179 27800
rect 4213 27766 4371 27800
rect 4405 27766 4563 27800
rect 4597 27766 4755 27800
rect 4789 27766 4947 27800
rect 4981 27766 4997 27800
rect 3971 27750 4997 27766
rect 4037 27718 4067 27750
rect 4133 27718 4163 27750
rect 4229 27718 4259 27750
rect 4325 27718 4355 27750
rect 4421 27718 4451 27750
rect 4517 27718 4547 27750
rect 4613 27718 4643 27750
rect 4709 27718 4739 27750
rect 4805 27718 4835 27750
rect 4901 27718 4931 27750
rect 5400 27505 5430 27531
rect 4037 27420 4067 27446
rect 4133 27420 4163 27446
rect 4229 27420 4259 27446
rect 4325 27420 4355 27446
rect 4421 27420 4451 27446
rect 4517 27420 4547 27446
rect 4613 27420 4643 27446
rect 4709 27420 4739 27446
rect 4805 27420 4835 27446
rect 4901 27420 4931 27446
rect 5400 27273 5430 27305
rect 5400 27257 5486 27273
rect 363 27134 393 27160
rect 459 27134 489 27160
rect 555 27134 585 27160
rect 651 27134 681 27160
rect 747 27134 777 27160
rect 843 27134 873 27160
rect 939 27134 969 27160
rect 1035 27134 1065 27160
rect 1131 27134 1161 27160
rect 1227 27134 1257 27160
rect 363 27008 393 27030
rect 459 27008 489 27030
rect 555 27008 585 27030
rect 651 27008 681 27030
rect 747 27008 777 27030
rect 843 27008 873 27030
rect 939 27008 969 27030
rect 1035 27008 1065 27030
rect 1131 27008 1161 27030
rect 1227 27008 1257 27030
rect 297 26988 1323 27008
rect 297 26954 313 26988
rect 347 26954 505 26988
rect 539 26954 697 26988
rect 731 26954 889 26988
rect 923 26954 1081 26988
rect 1115 26954 1273 26988
rect 1307 26954 1323 26988
rect 297 26942 1323 26954
rect 2516 27138 2546 27164
rect 2612 27138 2642 27164
rect 2708 27138 2738 27164
rect 2804 27138 2834 27164
rect 2900 27138 2930 27164
rect 2996 27138 3026 27164
rect 3092 27138 3122 27164
rect 3188 27138 3218 27164
rect 3284 27138 3314 27164
rect 3380 27138 3410 27164
rect 3675 27214 3741 27230
rect 3675 27180 3691 27214
rect 3725 27180 3741 27214
rect 3675 27164 3741 27180
rect 3693 27142 3723 27164
rect 4037 27138 4067 27164
rect 4133 27138 4163 27164
rect 4229 27138 4259 27164
rect 4325 27138 4355 27164
rect 4421 27138 4451 27164
rect 4517 27138 4547 27164
rect 4613 27138 4643 27164
rect 4709 27138 4739 27164
rect 4805 27138 4835 27164
rect 4901 27138 4931 27164
rect 5400 27223 5436 27257
rect 5470 27223 5486 27257
rect 5400 27207 5486 27223
rect 5400 27185 5430 27207
rect 2516 27012 2546 27034
rect 2612 27012 2642 27034
rect 2708 27012 2738 27034
rect 2804 27012 2834 27034
rect 2900 27012 2930 27034
rect 2996 27012 3026 27034
rect 3092 27012 3122 27034
rect 3188 27012 3218 27034
rect 3284 27012 3314 27034
rect 3380 27012 3410 27034
rect 2450 26992 3476 27012
rect 2450 26958 2466 26992
rect 2500 26958 2658 26992
rect 2692 26958 2850 26992
rect 2884 26958 3042 26992
rect 3076 26958 3234 26992
rect 3268 26958 3426 26992
rect 3460 26958 3476 26992
rect 2450 26946 3476 26958
rect 3693 27016 3723 27042
rect 4037 27012 4067 27034
rect 4133 27012 4163 27034
rect 4229 27012 4259 27034
rect 4325 27012 4355 27034
rect 4421 27012 4451 27034
rect 4517 27012 4547 27034
rect 4613 27012 4643 27034
rect 4709 27012 4739 27034
rect 4805 27012 4835 27034
rect 4901 27012 4931 27034
rect 3971 26992 4997 27012
rect 3971 26958 3987 26992
rect 4021 26958 4179 26992
rect 4213 26958 4371 26992
rect 4405 26958 4563 26992
rect 4597 26958 4755 26992
rect 4789 26958 4947 26992
rect 4981 26958 4997 26992
rect 3971 26946 4997 26958
rect 5400 27029 5430 27055
rect 297 26509 1323 26525
rect 297 26475 313 26509
rect 347 26475 505 26509
rect 539 26475 697 26509
rect 731 26475 889 26509
rect 923 26475 1081 26509
rect 1115 26475 1273 26509
rect 1307 26475 1323 26509
rect 297 26459 1323 26475
rect 363 26427 393 26459
rect 459 26427 489 26459
rect 555 26427 585 26459
rect 651 26427 681 26459
rect 747 26427 777 26459
rect 843 26427 873 26459
rect 939 26427 969 26459
rect 1035 26427 1065 26459
rect 1131 26427 1161 26459
rect 1227 26427 1257 26459
rect 363 26129 393 26155
rect 459 26129 489 26155
rect 555 26129 585 26155
rect 651 26129 681 26155
rect 747 26129 777 26155
rect 843 26129 873 26155
rect 939 26129 969 26155
rect 1035 26129 1065 26155
rect 1131 26129 1161 26155
rect 1227 26129 1257 26155
rect 2450 26513 3476 26529
rect 2450 26479 2466 26513
rect 2500 26479 2658 26513
rect 2692 26479 2850 26513
rect 2884 26479 3042 26513
rect 3076 26479 3234 26513
rect 3268 26479 3426 26513
rect 3460 26479 3476 26513
rect 2450 26463 3476 26479
rect 2516 26431 2546 26463
rect 2612 26431 2642 26463
rect 2708 26431 2738 26463
rect 2804 26431 2834 26463
rect 2900 26431 2930 26463
rect 2996 26431 3026 26463
rect 3092 26431 3122 26463
rect 3188 26431 3218 26463
rect 3284 26431 3314 26463
rect 3380 26431 3410 26463
rect 2516 26133 2546 26159
rect 2612 26133 2642 26159
rect 2708 26133 2738 26159
rect 2804 26133 2834 26159
rect 2900 26133 2930 26159
rect 2996 26133 3026 26159
rect 3092 26133 3122 26159
rect 3188 26133 3218 26159
rect 3284 26133 3314 26159
rect 3380 26133 3410 26159
rect 3971 26513 4997 26529
rect 3971 26479 3987 26513
rect 4021 26479 4179 26513
rect 4213 26479 4371 26513
rect 4405 26479 4563 26513
rect 4597 26479 4755 26513
rect 4789 26479 4947 26513
rect 4981 26479 4997 26513
rect 3971 26463 4997 26479
rect 4037 26431 4067 26463
rect 4133 26431 4163 26463
rect 4229 26431 4259 26463
rect 4325 26431 4355 26463
rect 4421 26431 4451 26463
rect 4517 26431 4547 26463
rect 4613 26431 4643 26463
rect 4709 26431 4739 26463
rect 4805 26431 4835 26463
rect 4901 26431 4931 26463
rect 5400 26218 5430 26244
rect 4037 26133 4067 26159
rect 4133 26133 4163 26159
rect 4229 26133 4259 26159
rect 4325 26133 4355 26159
rect 4421 26133 4451 26159
rect 4517 26133 4547 26159
rect 4613 26133 4643 26159
rect 4709 26133 4739 26159
rect 4805 26133 4835 26159
rect 4901 26133 4931 26159
rect 5400 25986 5430 26018
rect 5400 25970 5486 25986
rect 363 25847 393 25873
rect 459 25847 489 25873
rect 555 25847 585 25873
rect 651 25847 681 25873
rect 747 25847 777 25873
rect 843 25847 873 25873
rect 939 25847 969 25873
rect 1035 25847 1065 25873
rect 1131 25847 1161 25873
rect 1227 25847 1257 25873
rect 363 25721 393 25743
rect 459 25721 489 25743
rect 555 25721 585 25743
rect 651 25721 681 25743
rect 747 25721 777 25743
rect 843 25721 873 25743
rect 939 25721 969 25743
rect 1035 25721 1065 25743
rect 1131 25721 1161 25743
rect 1227 25721 1257 25743
rect 297 25701 1323 25721
rect 297 25667 313 25701
rect 347 25667 505 25701
rect 539 25667 697 25701
rect 731 25667 889 25701
rect 923 25667 1081 25701
rect 1115 25667 1273 25701
rect 1307 25667 1323 25701
rect 297 25655 1323 25667
rect 2516 25851 2546 25877
rect 2612 25851 2642 25877
rect 2708 25851 2738 25877
rect 2804 25851 2834 25877
rect 2900 25851 2930 25877
rect 2996 25851 3026 25877
rect 3092 25851 3122 25877
rect 3188 25851 3218 25877
rect 3284 25851 3314 25877
rect 3380 25851 3410 25877
rect 3675 25927 3741 25943
rect 3675 25893 3691 25927
rect 3725 25893 3741 25927
rect 3675 25877 3741 25893
rect 3693 25855 3723 25877
rect 4037 25851 4067 25877
rect 4133 25851 4163 25877
rect 4229 25851 4259 25877
rect 4325 25851 4355 25877
rect 4421 25851 4451 25877
rect 4517 25851 4547 25877
rect 4613 25851 4643 25877
rect 4709 25851 4739 25877
rect 4805 25851 4835 25877
rect 4901 25851 4931 25877
rect 5400 25936 5436 25970
rect 5470 25936 5486 25970
rect 5400 25920 5486 25936
rect 5400 25898 5430 25920
rect 2516 25725 2546 25747
rect 2612 25725 2642 25747
rect 2708 25725 2738 25747
rect 2804 25725 2834 25747
rect 2900 25725 2930 25747
rect 2996 25725 3026 25747
rect 3092 25725 3122 25747
rect 3188 25725 3218 25747
rect 3284 25725 3314 25747
rect 3380 25725 3410 25747
rect 2450 25705 3476 25725
rect 2450 25671 2466 25705
rect 2500 25671 2658 25705
rect 2692 25671 2850 25705
rect 2884 25671 3042 25705
rect 3076 25671 3234 25705
rect 3268 25671 3426 25705
rect 3460 25671 3476 25705
rect 2450 25659 3476 25671
rect 3693 25729 3723 25755
rect 4037 25725 4067 25747
rect 4133 25725 4163 25747
rect 4229 25725 4259 25747
rect 4325 25725 4355 25747
rect 4421 25725 4451 25747
rect 4517 25725 4547 25747
rect 4613 25725 4643 25747
rect 4709 25725 4739 25747
rect 4805 25725 4835 25747
rect 4901 25725 4931 25747
rect 3971 25705 4997 25725
rect 3971 25671 3987 25705
rect 4021 25671 4179 25705
rect 4213 25671 4371 25705
rect 4405 25671 4563 25705
rect 4597 25671 4755 25705
rect 4789 25671 4947 25705
rect 4981 25671 4997 25705
rect 3971 25659 4997 25671
rect 5400 25742 5430 25768
rect 297 25222 1323 25238
rect 297 25188 313 25222
rect 347 25188 505 25222
rect 539 25188 697 25222
rect 731 25188 889 25222
rect 923 25188 1081 25222
rect 1115 25188 1273 25222
rect 1307 25188 1323 25222
rect 297 25172 1323 25188
rect 363 25140 393 25172
rect 459 25140 489 25172
rect 555 25140 585 25172
rect 651 25140 681 25172
rect 747 25140 777 25172
rect 843 25140 873 25172
rect 939 25140 969 25172
rect 1035 25140 1065 25172
rect 1131 25140 1161 25172
rect 1227 25140 1257 25172
rect 363 24842 393 24868
rect 459 24842 489 24868
rect 555 24842 585 24868
rect 651 24842 681 24868
rect 747 24842 777 24868
rect 843 24842 873 24868
rect 939 24842 969 24868
rect 1035 24842 1065 24868
rect 1131 24842 1161 24868
rect 1227 24842 1257 24868
rect 2450 25226 3476 25242
rect 2450 25192 2466 25226
rect 2500 25192 2658 25226
rect 2692 25192 2850 25226
rect 2884 25192 3042 25226
rect 3076 25192 3234 25226
rect 3268 25192 3426 25226
rect 3460 25192 3476 25226
rect 2450 25176 3476 25192
rect 2516 25144 2546 25176
rect 2612 25144 2642 25176
rect 2708 25144 2738 25176
rect 2804 25144 2834 25176
rect 2900 25144 2930 25176
rect 2996 25144 3026 25176
rect 3092 25144 3122 25176
rect 3188 25144 3218 25176
rect 3284 25144 3314 25176
rect 3380 25144 3410 25176
rect 2516 24846 2546 24872
rect 2612 24846 2642 24872
rect 2708 24846 2738 24872
rect 2804 24846 2834 24872
rect 2900 24846 2930 24872
rect 2996 24846 3026 24872
rect 3092 24846 3122 24872
rect 3188 24846 3218 24872
rect 3284 24846 3314 24872
rect 3380 24846 3410 24872
rect 3971 25226 4997 25242
rect 3971 25192 3987 25226
rect 4021 25192 4179 25226
rect 4213 25192 4371 25226
rect 4405 25192 4563 25226
rect 4597 25192 4755 25226
rect 4789 25192 4947 25226
rect 4981 25192 4997 25226
rect 3971 25176 4997 25192
rect 4037 25144 4067 25176
rect 4133 25144 4163 25176
rect 4229 25144 4259 25176
rect 4325 25144 4355 25176
rect 4421 25144 4451 25176
rect 4517 25144 4547 25176
rect 4613 25144 4643 25176
rect 4709 25144 4739 25176
rect 4805 25144 4835 25176
rect 4901 25144 4931 25176
rect 5400 24931 5430 24957
rect 4037 24846 4067 24872
rect 4133 24846 4163 24872
rect 4229 24846 4259 24872
rect 4325 24846 4355 24872
rect 4421 24846 4451 24872
rect 4517 24846 4547 24872
rect 4613 24846 4643 24872
rect 4709 24846 4739 24872
rect 4805 24846 4835 24872
rect 4901 24846 4931 24872
rect 5400 24699 5430 24731
rect 5400 24683 5486 24699
rect 363 24560 393 24586
rect 459 24560 489 24586
rect 555 24560 585 24586
rect 651 24560 681 24586
rect 747 24560 777 24586
rect 843 24560 873 24586
rect 939 24560 969 24586
rect 1035 24560 1065 24586
rect 1131 24560 1161 24586
rect 1227 24560 1257 24586
rect 363 24434 393 24456
rect 459 24434 489 24456
rect 555 24434 585 24456
rect 651 24434 681 24456
rect 747 24434 777 24456
rect 843 24434 873 24456
rect 939 24434 969 24456
rect 1035 24434 1065 24456
rect 1131 24434 1161 24456
rect 1227 24434 1257 24456
rect 297 24414 1323 24434
rect 297 24380 313 24414
rect 347 24380 505 24414
rect 539 24380 697 24414
rect 731 24380 889 24414
rect 923 24380 1081 24414
rect 1115 24380 1273 24414
rect 1307 24380 1323 24414
rect 297 24368 1323 24380
rect 2516 24564 2546 24590
rect 2612 24564 2642 24590
rect 2708 24564 2738 24590
rect 2804 24564 2834 24590
rect 2900 24564 2930 24590
rect 2996 24564 3026 24590
rect 3092 24564 3122 24590
rect 3188 24564 3218 24590
rect 3284 24564 3314 24590
rect 3380 24564 3410 24590
rect 3675 24640 3741 24656
rect 3675 24606 3691 24640
rect 3725 24606 3741 24640
rect 3675 24590 3741 24606
rect 3693 24568 3723 24590
rect 4037 24564 4067 24590
rect 4133 24564 4163 24590
rect 4229 24564 4259 24590
rect 4325 24564 4355 24590
rect 4421 24564 4451 24590
rect 4517 24564 4547 24590
rect 4613 24564 4643 24590
rect 4709 24564 4739 24590
rect 4805 24564 4835 24590
rect 4901 24564 4931 24590
rect 5400 24649 5436 24683
rect 5470 24649 5486 24683
rect 5400 24633 5486 24649
rect 5400 24611 5430 24633
rect 2516 24438 2546 24460
rect 2612 24438 2642 24460
rect 2708 24438 2738 24460
rect 2804 24438 2834 24460
rect 2900 24438 2930 24460
rect 2996 24438 3026 24460
rect 3092 24438 3122 24460
rect 3188 24438 3218 24460
rect 3284 24438 3314 24460
rect 3380 24438 3410 24460
rect 2450 24418 3476 24438
rect 2450 24384 2466 24418
rect 2500 24384 2658 24418
rect 2692 24384 2850 24418
rect 2884 24384 3042 24418
rect 3076 24384 3234 24418
rect 3268 24384 3426 24418
rect 3460 24384 3476 24418
rect 2450 24372 3476 24384
rect 3693 24442 3723 24468
rect 4037 24438 4067 24460
rect 4133 24438 4163 24460
rect 4229 24438 4259 24460
rect 4325 24438 4355 24460
rect 4421 24438 4451 24460
rect 4517 24438 4547 24460
rect 4613 24438 4643 24460
rect 4709 24438 4739 24460
rect 4805 24438 4835 24460
rect 4901 24438 4931 24460
rect 3971 24418 4997 24438
rect 3971 24384 3987 24418
rect 4021 24384 4179 24418
rect 4213 24384 4371 24418
rect 4405 24384 4563 24418
rect 4597 24384 4755 24418
rect 4789 24384 4947 24418
rect 4981 24384 4997 24418
rect 3971 24372 4997 24384
rect 5400 24455 5430 24481
rect 297 23935 1323 23951
rect 297 23901 313 23935
rect 347 23901 505 23935
rect 539 23901 697 23935
rect 731 23901 889 23935
rect 923 23901 1081 23935
rect 1115 23901 1273 23935
rect 1307 23901 1323 23935
rect 297 23885 1323 23901
rect 363 23853 393 23885
rect 459 23853 489 23885
rect 555 23853 585 23885
rect 651 23853 681 23885
rect 747 23853 777 23885
rect 843 23853 873 23885
rect 939 23853 969 23885
rect 1035 23853 1065 23885
rect 1131 23853 1161 23885
rect 1227 23853 1257 23885
rect 363 23555 393 23581
rect 459 23555 489 23581
rect 555 23555 585 23581
rect 651 23555 681 23581
rect 747 23555 777 23581
rect 843 23555 873 23581
rect 939 23555 969 23581
rect 1035 23555 1065 23581
rect 1131 23555 1161 23581
rect 1227 23555 1257 23581
rect 2450 23939 3476 23955
rect 2450 23905 2466 23939
rect 2500 23905 2658 23939
rect 2692 23905 2850 23939
rect 2884 23905 3042 23939
rect 3076 23905 3234 23939
rect 3268 23905 3426 23939
rect 3460 23905 3476 23939
rect 2450 23889 3476 23905
rect 2516 23857 2546 23889
rect 2612 23857 2642 23889
rect 2708 23857 2738 23889
rect 2804 23857 2834 23889
rect 2900 23857 2930 23889
rect 2996 23857 3026 23889
rect 3092 23857 3122 23889
rect 3188 23857 3218 23889
rect 3284 23857 3314 23889
rect 3380 23857 3410 23889
rect 2516 23559 2546 23585
rect 2612 23559 2642 23585
rect 2708 23559 2738 23585
rect 2804 23559 2834 23585
rect 2900 23559 2930 23585
rect 2996 23559 3026 23585
rect 3092 23559 3122 23585
rect 3188 23559 3218 23585
rect 3284 23559 3314 23585
rect 3380 23559 3410 23585
rect 3971 23939 4997 23955
rect 3971 23905 3987 23939
rect 4021 23905 4179 23939
rect 4213 23905 4371 23939
rect 4405 23905 4563 23939
rect 4597 23905 4755 23939
rect 4789 23905 4947 23939
rect 4981 23905 4997 23939
rect 3971 23889 4997 23905
rect 4037 23857 4067 23889
rect 4133 23857 4163 23889
rect 4229 23857 4259 23889
rect 4325 23857 4355 23889
rect 4421 23857 4451 23889
rect 4517 23857 4547 23889
rect 4613 23857 4643 23889
rect 4709 23857 4739 23889
rect 4805 23857 4835 23889
rect 4901 23857 4931 23889
rect 5400 23644 5430 23670
rect 4037 23559 4067 23585
rect 4133 23559 4163 23585
rect 4229 23559 4259 23585
rect 4325 23559 4355 23585
rect 4421 23559 4451 23585
rect 4517 23559 4547 23585
rect 4613 23559 4643 23585
rect 4709 23559 4739 23585
rect 4805 23559 4835 23585
rect 4901 23559 4931 23585
rect 5400 23412 5430 23444
rect 5400 23396 5486 23412
rect 363 23273 393 23299
rect 459 23273 489 23299
rect 555 23273 585 23299
rect 651 23273 681 23299
rect 747 23273 777 23299
rect 843 23273 873 23299
rect 939 23273 969 23299
rect 1035 23273 1065 23299
rect 1131 23273 1161 23299
rect 1227 23273 1257 23299
rect 363 23147 393 23169
rect 459 23147 489 23169
rect 555 23147 585 23169
rect 651 23147 681 23169
rect 747 23147 777 23169
rect 843 23147 873 23169
rect 939 23147 969 23169
rect 1035 23147 1065 23169
rect 1131 23147 1161 23169
rect 1227 23147 1257 23169
rect 297 23127 1323 23147
rect 297 23093 313 23127
rect 347 23093 505 23127
rect 539 23093 697 23127
rect 731 23093 889 23127
rect 923 23093 1081 23127
rect 1115 23093 1273 23127
rect 1307 23093 1323 23127
rect 297 23081 1323 23093
rect 2516 23277 2546 23303
rect 2612 23277 2642 23303
rect 2708 23277 2738 23303
rect 2804 23277 2834 23303
rect 2900 23277 2930 23303
rect 2996 23277 3026 23303
rect 3092 23277 3122 23303
rect 3188 23277 3218 23303
rect 3284 23277 3314 23303
rect 3380 23277 3410 23303
rect 3675 23353 3741 23369
rect 3675 23319 3691 23353
rect 3725 23319 3741 23353
rect 3675 23303 3741 23319
rect 3693 23281 3723 23303
rect 4037 23277 4067 23303
rect 4133 23277 4163 23303
rect 4229 23277 4259 23303
rect 4325 23277 4355 23303
rect 4421 23277 4451 23303
rect 4517 23277 4547 23303
rect 4613 23277 4643 23303
rect 4709 23277 4739 23303
rect 4805 23277 4835 23303
rect 4901 23277 4931 23303
rect 5400 23362 5436 23396
rect 5470 23362 5486 23396
rect 5400 23346 5486 23362
rect 5400 23324 5430 23346
rect 2516 23151 2546 23173
rect 2612 23151 2642 23173
rect 2708 23151 2738 23173
rect 2804 23151 2834 23173
rect 2900 23151 2930 23173
rect 2996 23151 3026 23173
rect 3092 23151 3122 23173
rect 3188 23151 3218 23173
rect 3284 23151 3314 23173
rect 3380 23151 3410 23173
rect 2450 23131 3476 23151
rect 2450 23097 2466 23131
rect 2500 23097 2658 23131
rect 2692 23097 2850 23131
rect 2884 23097 3042 23131
rect 3076 23097 3234 23131
rect 3268 23097 3426 23131
rect 3460 23097 3476 23131
rect 2450 23085 3476 23097
rect 3693 23155 3723 23181
rect 4037 23151 4067 23173
rect 4133 23151 4163 23173
rect 4229 23151 4259 23173
rect 4325 23151 4355 23173
rect 4421 23151 4451 23173
rect 4517 23151 4547 23173
rect 4613 23151 4643 23173
rect 4709 23151 4739 23173
rect 4805 23151 4835 23173
rect 4901 23151 4931 23173
rect 3971 23131 4997 23151
rect 3971 23097 3987 23131
rect 4021 23097 4179 23131
rect 4213 23097 4371 23131
rect 4405 23097 4563 23131
rect 4597 23097 4755 23131
rect 4789 23097 4947 23131
rect 4981 23097 4997 23131
rect 3971 23085 4997 23097
rect 5400 23168 5430 23194
rect 297 22648 1323 22664
rect 297 22614 313 22648
rect 347 22614 505 22648
rect 539 22614 697 22648
rect 731 22614 889 22648
rect 923 22614 1081 22648
rect 1115 22614 1273 22648
rect 1307 22614 1323 22648
rect 297 22598 1323 22614
rect 363 22566 393 22598
rect 459 22566 489 22598
rect 555 22566 585 22598
rect 651 22566 681 22598
rect 747 22566 777 22598
rect 843 22566 873 22598
rect 939 22566 969 22598
rect 1035 22566 1065 22598
rect 1131 22566 1161 22598
rect 1227 22566 1257 22598
rect 363 22268 393 22294
rect 459 22268 489 22294
rect 555 22268 585 22294
rect 651 22268 681 22294
rect 747 22268 777 22294
rect 843 22268 873 22294
rect 939 22268 969 22294
rect 1035 22268 1065 22294
rect 1131 22268 1161 22294
rect 1227 22268 1257 22294
rect 2450 22652 3476 22668
rect 2450 22618 2466 22652
rect 2500 22618 2658 22652
rect 2692 22618 2850 22652
rect 2884 22618 3042 22652
rect 3076 22618 3234 22652
rect 3268 22618 3426 22652
rect 3460 22618 3476 22652
rect 2450 22602 3476 22618
rect 2516 22570 2546 22602
rect 2612 22570 2642 22602
rect 2708 22570 2738 22602
rect 2804 22570 2834 22602
rect 2900 22570 2930 22602
rect 2996 22570 3026 22602
rect 3092 22570 3122 22602
rect 3188 22570 3218 22602
rect 3284 22570 3314 22602
rect 3380 22570 3410 22602
rect 2516 22272 2546 22298
rect 2612 22272 2642 22298
rect 2708 22272 2738 22298
rect 2804 22272 2834 22298
rect 2900 22272 2930 22298
rect 2996 22272 3026 22298
rect 3092 22272 3122 22298
rect 3188 22272 3218 22298
rect 3284 22272 3314 22298
rect 3380 22272 3410 22298
rect 3971 22652 4997 22668
rect 3971 22618 3987 22652
rect 4021 22618 4179 22652
rect 4213 22618 4371 22652
rect 4405 22618 4563 22652
rect 4597 22618 4755 22652
rect 4789 22618 4947 22652
rect 4981 22618 4997 22652
rect 3971 22602 4997 22618
rect 4037 22570 4067 22602
rect 4133 22570 4163 22602
rect 4229 22570 4259 22602
rect 4325 22570 4355 22602
rect 4421 22570 4451 22602
rect 4517 22570 4547 22602
rect 4613 22570 4643 22602
rect 4709 22570 4739 22602
rect 4805 22570 4835 22602
rect 4901 22570 4931 22602
rect 5400 22357 5430 22383
rect 4037 22272 4067 22298
rect 4133 22272 4163 22298
rect 4229 22272 4259 22298
rect 4325 22272 4355 22298
rect 4421 22272 4451 22298
rect 4517 22272 4547 22298
rect 4613 22272 4643 22298
rect 4709 22272 4739 22298
rect 4805 22272 4835 22298
rect 4901 22272 4931 22298
rect 5400 22125 5430 22157
rect 5400 22109 5486 22125
rect 363 21986 393 22012
rect 459 21986 489 22012
rect 555 21986 585 22012
rect 651 21986 681 22012
rect 747 21986 777 22012
rect 843 21986 873 22012
rect 939 21986 969 22012
rect 1035 21986 1065 22012
rect 1131 21986 1161 22012
rect 1227 21986 1257 22012
rect 363 21860 393 21882
rect 459 21860 489 21882
rect 555 21860 585 21882
rect 651 21860 681 21882
rect 747 21860 777 21882
rect 843 21860 873 21882
rect 939 21860 969 21882
rect 1035 21860 1065 21882
rect 1131 21860 1161 21882
rect 1227 21860 1257 21882
rect 297 21840 1323 21860
rect 297 21806 313 21840
rect 347 21806 505 21840
rect 539 21806 697 21840
rect 731 21806 889 21840
rect 923 21806 1081 21840
rect 1115 21806 1273 21840
rect 1307 21806 1323 21840
rect 297 21794 1323 21806
rect 2516 21990 2546 22016
rect 2612 21990 2642 22016
rect 2708 21990 2738 22016
rect 2804 21990 2834 22016
rect 2900 21990 2930 22016
rect 2996 21990 3026 22016
rect 3092 21990 3122 22016
rect 3188 21990 3218 22016
rect 3284 21990 3314 22016
rect 3380 21990 3410 22016
rect 3675 22066 3741 22082
rect 3675 22032 3691 22066
rect 3725 22032 3741 22066
rect 3675 22016 3741 22032
rect 3693 21994 3723 22016
rect 4037 21990 4067 22016
rect 4133 21990 4163 22016
rect 4229 21990 4259 22016
rect 4325 21990 4355 22016
rect 4421 21990 4451 22016
rect 4517 21990 4547 22016
rect 4613 21990 4643 22016
rect 4709 21990 4739 22016
rect 4805 21990 4835 22016
rect 4901 21990 4931 22016
rect 5400 22075 5436 22109
rect 5470 22075 5486 22109
rect 5400 22059 5486 22075
rect 5400 22037 5430 22059
rect 2516 21864 2546 21886
rect 2612 21864 2642 21886
rect 2708 21864 2738 21886
rect 2804 21864 2834 21886
rect 2900 21864 2930 21886
rect 2996 21864 3026 21886
rect 3092 21864 3122 21886
rect 3188 21864 3218 21886
rect 3284 21864 3314 21886
rect 3380 21864 3410 21886
rect 2450 21844 3476 21864
rect 2450 21810 2466 21844
rect 2500 21810 2658 21844
rect 2692 21810 2850 21844
rect 2884 21810 3042 21844
rect 3076 21810 3234 21844
rect 3268 21810 3426 21844
rect 3460 21810 3476 21844
rect 2450 21798 3476 21810
rect 3693 21868 3723 21894
rect 4037 21864 4067 21886
rect 4133 21864 4163 21886
rect 4229 21864 4259 21886
rect 4325 21864 4355 21886
rect 4421 21864 4451 21886
rect 4517 21864 4547 21886
rect 4613 21864 4643 21886
rect 4709 21864 4739 21886
rect 4805 21864 4835 21886
rect 4901 21864 4931 21886
rect 3971 21844 4997 21864
rect 3971 21810 3987 21844
rect 4021 21810 4179 21844
rect 4213 21810 4371 21844
rect 4405 21810 4563 21844
rect 4597 21810 4755 21844
rect 4789 21810 4947 21844
rect 4981 21810 4997 21844
rect 3971 21798 4997 21810
rect 5400 21881 5430 21907
rect 297 21361 1323 21377
rect 297 21327 313 21361
rect 347 21327 505 21361
rect 539 21327 697 21361
rect 731 21327 889 21361
rect 923 21327 1081 21361
rect 1115 21327 1273 21361
rect 1307 21327 1323 21361
rect 297 21311 1323 21327
rect 363 21279 393 21311
rect 459 21279 489 21311
rect 555 21279 585 21311
rect 651 21279 681 21311
rect 747 21279 777 21311
rect 843 21279 873 21311
rect 939 21279 969 21311
rect 1035 21279 1065 21311
rect 1131 21279 1161 21311
rect 1227 21279 1257 21311
rect 363 20981 393 21007
rect 459 20981 489 21007
rect 555 20981 585 21007
rect 651 20981 681 21007
rect 747 20981 777 21007
rect 843 20981 873 21007
rect 939 20981 969 21007
rect 1035 20981 1065 21007
rect 1131 20981 1161 21007
rect 1227 20981 1257 21007
rect 2450 21365 3476 21381
rect 2450 21331 2466 21365
rect 2500 21331 2658 21365
rect 2692 21331 2850 21365
rect 2884 21331 3042 21365
rect 3076 21331 3234 21365
rect 3268 21331 3426 21365
rect 3460 21331 3476 21365
rect 2450 21315 3476 21331
rect 2516 21283 2546 21315
rect 2612 21283 2642 21315
rect 2708 21283 2738 21315
rect 2804 21283 2834 21315
rect 2900 21283 2930 21315
rect 2996 21283 3026 21315
rect 3092 21283 3122 21315
rect 3188 21283 3218 21315
rect 3284 21283 3314 21315
rect 3380 21283 3410 21315
rect 2516 20985 2546 21011
rect 2612 20985 2642 21011
rect 2708 20985 2738 21011
rect 2804 20985 2834 21011
rect 2900 20985 2930 21011
rect 2996 20985 3026 21011
rect 3092 20985 3122 21011
rect 3188 20985 3218 21011
rect 3284 20985 3314 21011
rect 3380 20985 3410 21011
rect 3971 21365 4997 21381
rect 3971 21331 3987 21365
rect 4021 21331 4179 21365
rect 4213 21331 4371 21365
rect 4405 21331 4563 21365
rect 4597 21331 4755 21365
rect 4789 21331 4947 21365
rect 4981 21331 4997 21365
rect 3971 21315 4997 21331
rect 4037 21283 4067 21315
rect 4133 21283 4163 21315
rect 4229 21283 4259 21315
rect 4325 21283 4355 21315
rect 4421 21283 4451 21315
rect 4517 21283 4547 21315
rect 4613 21283 4643 21315
rect 4709 21283 4739 21315
rect 4805 21283 4835 21315
rect 4901 21283 4931 21315
rect 5400 21070 5430 21096
rect 4037 20985 4067 21011
rect 4133 20985 4163 21011
rect 4229 20985 4259 21011
rect 4325 20985 4355 21011
rect 4421 20985 4451 21011
rect 4517 20985 4547 21011
rect 4613 20985 4643 21011
rect 4709 20985 4739 21011
rect 4805 20985 4835 21011
rect 4901 20985 4931 21011
rect 5400 20838 5430 20870
rect 5400 20822 5486 20838
rect 363 20699 393 20725
rect 459 20699 489 20725
rect 555 20699 585 20725
rect 651 20699 681 20725
rect 747 20699 777 20725
rect 843 20699 873 20725
rect 939 20699 969 20725
rect 1035 20699 1065 20725
rect 1131 20699 1161 20725
rect 1227 20699 1257 20725
rect 363 20573 393 20595
rect 459 20573 489 20595
rect 555 20573 585 20595
rect 651 20573 681 20595
rect 747 20573 777 20595
rect 843 20573 873 20595
rect 939 20573 969 20595
rect 1035 20573 1065 20595
rect 1131 20573 1161 20595
rect 1227 20573 1257 20595
rect 297 20553 1323 20573
rect 297 20519 313 20553
rect 347 20519 505 20553
rect 539 20519 697 20553
rect 731 20519 889 20553
rect 923 20519 1081 20553
rect 1115 20519 1273 20553
rect 1307 20519 1323 20553
rect 297 20507 1323 20519
rect 2516 20703 2546 20729
rect 2612 20703 2642 20729
rect 2708 20703 2738 20729
rect 2804 20703 2834 20729
rect 2900 20703 2930 20729
rect 2996 20703 3026 20729
rect 3092 20703 3122 20729
rect 3188 20703 3218 20729
rect 3284 20703 3314 20729
rect 3380 20703 3410 20729
rect 3675 20779 3741 20795
rect 3675 20745 3691 20779
rect 3725 20745 3741 20779
rect 3675 20729 3741 20745
rect 3693 20707 3723 20729
rect 4037 20703 4067 20729
rect 4133 20703 4163 20729
rect 4229 20703 4259 20729
rect 4325 20703 4355 20729
rect 4421 20703 4451 20729
rect 4517 20703 4547 20729
rect 4613 20703 4643 20729
rect 4709 20703 4739 20729
rect 4805 20703 4835 20729
rect 4901 20703 4931 20729
rect 5400 20788 5436 20822
rect 5470 20788 5486 20822
rect 5400 20772 5486 20788
rect 5400 20750 5430 20772
rect 2516 20577 2546 20599
rect 2612 20577 2642 20599
rect 2708 20577 2738 20599
rect 2804 20577 2834 20599
rect 2900 20577 2930 20599
rect 2996 20577 3026 20599
rect 3092 20577 3122 20599
rect 3188 20577 3218 20599
rect 3284 20577 3314 20599
rect 3380 20577 3410 20599
rect 2450 20557 3476 20577
rect 2450 20523 2466 20557
rect 2500 20523 2658 20557
rect 2692 20523 2850 20557
rect 2884 20523 3042 20557
rect 3076 20523 3234 20557
rect 3268 20523 3426 20557
rect 3460 20523 3476 20557
rect 2450 20511 3476 20523
rect 3693 20581 3723 20607
rect 4037 20577 4067 20599
rect 4133 20577 4163 20599
rect 4229 20577 4259 20599
rect 4325 20577 4355 20599
rect 4421 20577 4451 20599
rect 4517 20577 4547 20599
rect 4613 20577 4643 20599
rect 4709 20577 4739 20599
rect 4805 20577 4835 20599
rect 4901 20577 4931 20599
rect 3971 20557 4997 20577
rect 3971 20523 3987 20557
rect 4021 20523 4179 20557
rect 4213 20523 4371 20557
rect 4405 20523 4563 20557
rect 4597 20523 4755 20557
rect 4789 20523 4947 20557
rect 4981 20523 4997 20557
rect 3971 20511 4997 20523
rect 5400 20594 5430 20620
rect 297 20074 1323 20090
rect 297 20040 313 20074
rect 347 20040 505 20074
rect 539 20040 697 20074
rect 731 20040 889 20074
rect 923 20040 1081 20074
rect 1115 20040 1273 20074
rect 1307 20040 1323 20074
rect 297 20024 1323 20040
rect 363 19992 393 20024
rect 459 19992 489 20024
rect 555 19992 585 20024
rect 651 19992 681 20024
rect 747 19992 777 20024
rect 843 19992 873 20024
rect 939 19992 969 20024
rect 1035 19992 1065 20024
rect 1131 19992 1161 20024
rect 1227 19992 1257 20024
rect 363 19694 393 19720
rect 459 19694 489 19720
rect 555 19694 585 19720
rect 651 19694 681 19720
rect 747 19694 777 19720
rect 843 19694 873 19720
rect 939 19694 969 19720
rect 1035 19694 1065 19720
rect 1131 19694 1161 19720
rect 1227 19694 1257 19720
rect 2450 20078 3476 20094
rect 2450 20044 2466 20078
rect 2500 20044 2658 20078
rect 2692 20044 2850 20078
rect 2884 20044 3042 20078
rect 3076 20044 3234 20078
rect 3268 20044 3426 20078
rect 3460 20044 3476 20078
rect 2450 20028 3476 20044
rect 2516 19996 2546 20028
rect 2612 19996 2642 20028
rect 2708 19996 2738 20028
rect 2804 19996 2834 20028
rect 2900 19996 2930 20028
rect 2996 19996 3026 20028
rect 3092 19996 3122 20028
rect 3188 19996 3218 20028
rect 3284 19996 3314 20028
rect 3380 19996 3410 20028
rect 2516 19698 2546 19724
rect 2612 19698 2642 19724
rect 2708 19698 2738 19724
rect 2804 19698 2834 19724
rect 2900 19698 2930 19724
rect 2996 19698 3026 19724
rect 3092 19698 3122 19724
rect 3188 19698 3218 19724
rect 3284 19698 3314 19724
rect 3380 19698 3410 19724
rect 3971 20078 4997 20094
rect 3971 20044 3987 20078
rect 4021 20044 4179 20078
rect 4213 20044 4371 20078
rect 4405 20044 4563 20078
rect 4597 20044 4755 20078
rect 4789 20044 4947 20078
rect 4981 20044 4997 20078
rect 3971 20028 4997 20044
rect 4037 19996 4067 20028
rect 4133 19996 4163 20028
rect 4229 19996 4259 20028
rect 4325 19996 4355 20028
rect 4421 19996 4451 20028
rect 4517 19996 4547 20028
rect 4613 19996 4643 20028
rect 4709 19996 4739 20028
rect 4805 19996 4835 20028
rect 4901 19996 4931 20028
rect 5400 19783 5430 19809
rect 4037 19698 4067 19724
rect 4133 19698 4163 19724
rect 4229 19698 4259 19724
rect 4325 19698 4355 19724
rect 4421 19698 4451 19724
rect 4517 19698 4547 19724
rect 4613 19698 4643 19724
rect 4709 19698 4739 19724
rect 4805 19698 4835 19724
rect 4901 19698 4931 19724
rect 5400 19551 5430 19583
rect 5400 19535 5486 19551
rect 363 19412 393 19438
rect 459 19412 489 19438
rect 555 19412 585 19438
rect 651 19412 681 19438
rect 747 19412 777 19438
rect 843 19412 873 19438
rect 939 19412 969 19438
rect 1035 19412 1065 19438
rect 1131 19412 1161 19438
rect 1227 19412 1257 19438
rect 363 19286 393 19308
rect 459 19286 489 19308
rect 555 19286 585 19308
rect 651 19286 681 19308
rect 747 19286 777 19308
rect 843 19286 873 19308
rect 939 19286 969 19308
rect 1035 19286 1065 19308
rect 1131 19286 1161 19308
rect 1227 19286 1257 19308
rect 297 19266 1323 19286
rect 297 19232 313 19266
rect 347 19232 505 19266
rect 539 19232 697 19266
rect 731 19232 889 19266
rect 923 19232 1081 19266
rect 1115 19232 1273 19266
rect 1307 19232 1323 19266
rect 297 19220 1323 19232
rect 2516 19416 2546 19442
rect 2612 19416 2642 19442
rect 2708 19416 2738 19442
rect 2804 19416 2834 19442
rect 2900 19416 2930 19442
rect 2996 19416 3026 19442
rect 3092 19416 3122 19442
rect 3188 19416 3218 19442
rect 3284 19416 3314 19442
rect 3380 19416 3410 19442
rect 3675 19492 3741 19508
rect 3675 19458 3691 19492
rect 3725 19458 3741 19492
rect 3675 19442 3741 19458
rect 3693 19420 3723 19442
rect 4037 19416 4067 19442
rect 4133 19416 4163 19442
rect 4229 19416 4259 19442
rect 4325 19416 4355 19442
rect 4421 19416 4451 19442
rect 4517 19416 4547 19442
rect 4613 19416 4643 19442
rect 4709 19416 4739 19442
rect 4805 19416 4835 19442
rect 4901 19416 4931 19442
rect 5400 19501 5436 19535
rect 5470 19501 5486 19535
rect 5400 19485 5486 19501
rect 5400 19463 5430 19485
rect 2516 19290 2546 19312
rect 2612 19290 2642 19312
rect 2708 19290 2738 19312
rect 2804 19290 2834 19312
rect 2900 19290 2930 19312
rect 2996 19290 3026 19312
rect 3092 19290 3122 19312
rect 3188 19290 3218 19312
rect 3284 19290 3314 19312
rect 3380 19290 3410 19312
rect 2450 19270 3476 19290
rect 2450 19236 2466 19270
rect 2500 19236 2658 19270
rect 2692 19236 2850 19270
rect 2884 19236 3042 19270
rect 3076 19236 3234 19270
rect 3268 19236 3426 19270
rect 3460 19236 3476 19270
rect 2450 19224 3476 19236
rect 3693 19294 3723 19320
rect 4037 19290 4067 19312
rect 4133 19290 4163 19312
rect 4229 19290 4259 19312
rect 4325 19290 4355 19312
rect 4421 19290 4451 19312
rect 4517 19290 4547 19312
rect 4613 19290 4643 19312
rect 4709 19290 4739 19312
rect 4805 19290 4835 19312
rect 4901 19290 4931 19312
rect 3971 19270 4997 19290
rect 3971 19236 3987 19270
rect 4021 19236 4179 19270
rect 4213 19236 4371 19270
rect 4405 19236 4563 19270
rect 4597 19236 4755 19270
rect 4789 19236 4947 19270
rect 4981 19236 4997 19270
rect 3971 19224 4997 19236
rect 5400 19307 5430 19333
rect 297 18787 1323 18803
rect 297 18753 313 18787
rect 347 18753 505 18787
rect 539 18753 697 18787
rect 731 18753 889 18787
rect 923 18753 1081 18787
rect 1115 18753 1273 18787
rect 1307 18753 1323 18787
rect 297 18737 1323 18753
rect 363 18705 393 18737
rect 459 18705 489 18737
rect 555 18705 585 18737
rect 651 18705 681 18737
rect 747 18705 777 18737
rect 843 18705 873 18737
rect 939 18705 969 18737
rect 1035 18705 1065 18737
rect 1131 18705 1161 18737
rect 1227 18705 1257 18737
rect 363 18407 393 18433
rect 459 18407 489 18433
rect 555 18407 585 18433
rect 651 18407 681 18433
rect 747 18407 777 18433
rect 843 18407 873 18433
rect 939 18407 969 18433
rect 1035 18407 1065 18433
rect 1131 18407 1161 18433
rect 1227 18407 1257 18433
rect 2450 18791 3476 18807
rect 2450 18757 2466 18791
rect 2500 18757 2658 18791
rect 2692 18757 2850 18791
rect 2884 18757 3042 18791
rect 3076 18757 3234 18791
rect 3268 18757 3426 18791
rect 3460 18757 3476 18791
rect 2450 18741 3476 18757
rect 2516 18709 2546 18741
rect 2612 18709 2642 18741
rect 2708 18709 2738 18741
rect 2804 18709 2834 18741
rect 2900 18709 2930 18741
rect 2996 18709 3026 18741
rect 3092 18709 3122 18741
rect 3188 18709 3218 18741
rect 3284 18709 3314 18741
rect 3380 18709 3410 18741
rect 2516 18411 2546 18437
rect 2612 18411 2642 18437
rect 2708 18411 2738 18437
rect 2804 18411 2834 18437
rect 2900 18411 2930 18437
rect 2996 18411 3026 18437
rect 3092 18411 3122 18437
rect 3188 18411 3218 18437
rect 3284 18411 3314 18437
rect 3380 18411 3410 18437
rect 3971 18791 4997 18807
rect 3971 18757 3987 18791
rect 4021 18757 4179 18791
rect 4213 18757 4371 18791
rect 4405 18757 4563 18791
rect 4597 18757 4755 18791
rect 4789 18757 4947 18791
rect 4981 18757 4997 18791
rect 3971 18741 4997 18757
rect 4037 18709 4067 18741
rect 4133 18709 4163 18741
rect 4229 18709 4259 18741
rect 4325 18709 4355 18741
rect 4421 18709 4451 18741
rect 4517 18709 4547 18741
rect 4613 18709 4643 18741
rect 4709 18709 4739 18741
rect 4805 18709 4835 18741
rect 4901 18709 4931 18741
rect 5400 18496 5430 18522
rect 4037 18411 4067 18437
rect 4133 18411 4163 18437
rect 4229 18411 4259 18437
rect 4325 18411 4355 18437
rect 4421 18411 4451 18437
rect 4517 18411 4547 18437
rect 4613 18411 4643 18437
rect 4709 18411 4739 18437
rect 4805 18411 4835 18437
rect 4901 18411 4931 18437
rect 5400 18264 5430 18296
rect 5400 18248 5486 18264
rect 363 18125 393 18151
rect 459 18125 489 18151
rect 555 18125 585 18151
rect 651 18125 681 18151
rect 747 18125 777 18151
rect 843 18125 873 18151
rect 939 18125 969 18151
rect 1035 18125 1065 18151
rect 1131 18125 1161 18151
rect 1227 18125 1257 18151
rect 363 17999 393 18021
rect 459 17999 489 18021
rect 555 17999 585 18021
rect 651 17999 681 18021
rect 747 17999 777 18021
rect 843 17999 873 18021
rect 939 17999 969 18021
rect 1035 17999 1065 18021
rect 1131 17999 1161 18021
rect 1227 17999 1257 18021
rect 297 17979 1323 17999
rect 297 17945 313 17979
rect 347 17945 505 17979
rect 539 17945 697 17979
rect 731 17945 889 17979
rect 923 17945 1081 17979
rect 1115 17945 1273 17979
rect 1307 17945 1323 17979
rect 297 17933 1323 17945
rect 2516 18129 2546 18155
rect 2612 18129 2642 18155
rect 2708 18129 2738 18155
rect 2804 18129 2834 18155
rect 2900 18129 2930 18155
rect 2996 18129 3026 18155
rect 3092 18129 3122 18155
rect 3188 18129 3218 18155
rect 3284 18129 3314 18155
rect 3380 18129 3410 18155
rect 3675 18205 3741 18221
rect 3675 18171 3691 18205
rect 3725 18171 3741 18205
rect 3675 18155 3741 18171
rect 3693 18133 3723 18155
rect 4037 18129 4067 18155
rect 4133 18129 4163 18155
rect 4229 18129 4259 18155
rect 4325 18129 4355 18155
rect 4421 18129 4451 18155
rect 4517 18129 4547 18155
rect 4613 18129 4643 18155
rect 4709 18129 4739 18155
rect 4805 18129 4835 18155
rect 4901 18129 4931 18155
rect 5400 18214 5436 18248
rect 5470 18214 5486 18248
rect 5400 18198 5486 18214
rect 5400 18176 5430 18198
rect 2516 18003 2546 18025
rect 2612 18003 2642 18025
rect 2708 18003 2738 18025
rect 2804 18003 2834 18025
rect 2900 18003 2930 18025
rect 2996 18003 3026 18025
rect 3092 18003 3122 18025
rect 3188 18003 3218 18025
rect 3284 18003 3314 18025
rect 3380 18003 3410 18025
rect 2450 17983 3476 18003
rect 2450 17949 2466 17983
rect 2500 17949 2658 17983
rect 2692 17949 2850 17983
rect 2884 17949 3042 17983
rect 3076 17949 3234 17983
rect 3268 17949 3426 17983
rect 3460 17949 3476 17983
rect 2450 17937 3476 17949
rect 3693 18007 3723 18033
rect 4037 18003 4067 18025
rect 4133 18003 4163 18025
rect 4229 18003 4259 18025
rect 4325 18003 4355 18025
rect 4421 18003 4451 18025
rect 4517 18003 4547 18025
rect 4613 18003 4643 18025
rect 4709 18003 4739 18025
rect 4805 18003 4835 18025
rect 4901 18003 4931 18025
rect 3971 17983 4997 18003
rect 3971 17949 3987 17983
rect 4021 17949 4179 17983
rect 4213 17949 4371 17983
rect 4405 17949 4563 17983
rect 4597 17949 4755 17983
rect 4789 17949 4947 17983
rect 4981 17949 4997 17983
rect 3971 17937 4997 17949
rect 5400 18020 5430 18046
rect 297 17500 1323 17516
rect 297 17466 313 17500
rect 347 17466 505 17500
rect 539 17466 697 17500
rect 731 17466 889 17500
rect 923 17466 1081 17500
rect 1115 17466 1273 17500
rect 1307 17466 1323 17500
rect 297 17450 1323 17466
rect 363 17418 393 17450
rect 459 17418 489 17450
rect 555 17418 585 17450
rect 651 17418 681 17450
rect 747 17418 777 17450
rect 843 17418 873 17450
rect 939 17418 969 17450
rect 1035 17418 1065 17450
rect 1131 17418 1161 17450
rect 1227 17418 1257 17450
rect 363 17120 393 17146
rect 459 17120 489 17146
rect 555 17120 585 17146
rect 651 17120 681 17146
rect 747 17120 777 17146
rect 843 17120 873 17146
rect 939 17120 969 17146
rect 1035 17120 1065 17146
rect 1131 17120 1161 17146
rect 1227 17120 1257 17146
rect 2450 17504 3476 17520
rect 2450 17470 2466 17504
rect 2500 17470 2658 17504
rect 2692 17470 2850 17504
rect 2884 17470 3042 17504
rect 3076 17470 3234 17504
rect 3268 17470 3426 17504
rect 3460 17470 3476 17504
rect 2450 17454 3476 17470
rect 2516 17422 2546 17454
rect 2612 17422 2642 17454
rect 2708 17422 2738 17454
rect 2804 17422 2834 17454
rect 2900 17422 2930 17454
rect 2996 17422 3026 17454
rect 3092 17422 3122 17454
rect 3188 17422 3218 17454
rect 3284 17422 3314 17454
rect 3380 17422 3410 17454
rect 2516 17124 2546 17150
rect 2612 17124 2642 17150
rect 2708 17124 2738 17150
rect 2804 17124 2834 17150
rect 2900 17124 2930 17150
rect 2996 17124 3026 17150
rect 3092 17124 3122 17150
rect 3188 17124 3218 17150
rect 3284 17124 3314 17150
rect 3380 17124 3410 17150
rect 3971 17504 4997 17520
rect 3971 17470 3987 17504
rect 4021 17470 4179 17504
rect 4213 17470 4371 17504
rect 4405 17470 4563 17504
rect 4597 17470 4755 17504
rect 4789 17470 4947 17504
rect 4981 17470 4997 17504
rect 3971 17454 4997 17470
rect 4037 17422 4067 17454
rect 4133 17422 4163 17454
rect 4229 17422 4259 17454
rect 4325 17422 4355 17454
rect 4421 17422 4451 17454
rect 4517 17422 4547 17454
rect 4613 17422 4643 17454
rect 4709 17422 4739 17454
rect 4805 17422 4835 17454
rect 4901 17422 4931 17454
rect 5400 17209 5430 17235
rect 4037 17124 4067 17150
rect 4133 17124 4163 17150
rect 4229 17124 4259 17150
rect 4325 17124 4355 17150
rect 4421 17124 4451 17150
rect 4517 17124 4547 17150
rect 4613 17124 4643 17150
rect 4709 17124 4739 17150
rect 4805 17124 4835 17150
rect 4901 17124 4931 17150
rect 5400 16977 5430 17009
rect 5400 16961 5486 16977
rect 363 16838 393 16864
rect 459 16838 489 16864
rect 555 16838 585 16864
rect 651 16838 681 16864
rect 747 16838 777 16864
rect 843 16838 873 16864
rect 939 16838 969 16864
rect 1035 16838 1065 16864
rect 1131 16838 1161 16864
rect 1227 16838 1257 16864
rect 363 16712 393 16734
rect 459 16712 489 16734
rect 555 16712 585 16734
rect 651 16712 681 16734
rect 747 16712 777 16734
rect 843 16712 873 16734
rect 939 16712 969 16734
rect 1035 16712 1065 16734
rect 1131 16712 1161 16734
rect 1227 16712 1257 16734
rect 297 16692 1323 16712
rect 297 16658 313 16692
rect 347 16658 505 16692
rect 539 16658 697 16692
rect 731 16658 889 16692
rect 923 16658 1081 16692
rect 1115 16658 1273 16692
rect 1307 16658 1323 16692
rect 297 16646 1323 16658
rect 2516 16842 2546 16868
rect 2612 16842 2642 16868
rect 2708 16842 2738 16868
rect 2804 16842 2834 16868
rect 2900 16842 2930 16868
rect 2996 16842 3026 16868
rect 3092 16842 3122 16868
rect 3188 16842 3218 16868
rect 3284 16842 3314 16868
rect 3380 16842 3410 16868
rect 3675 16918 3741 16934
rect 3675 16884 3691 16918
rect 3725 16884 3741 16918
rect 3675 16868 3741 16884
rect 3693 16846 3723 16868
rect 4037 16842 4067 16868
rect 4133 16842 4163 16868
rect 4229 16842 4259 16868
rect 4325 16842 4355 16868
rect 4421 16842 4451 16868
rect 4517 16842 4547 16868
rect 4613 16842 4643 16868
rect 4709 16842 4739 16868
rect 4805 16842 4835 16868
rect 4901 16842 4931 16868
rect 5400 16927 5436 16961
rect 5470 16927 5486 16961
rect 5400 16911 5486 16927
rect 5400 16889 5430 16911
rect 2516 16716 2546 16738
rect 2612 16716 2642 16738
rect 2708 16716 2738 16738
rect 2804 16716 2834 16738
rect 2900 16716 2930 16738
rect 2996 16716 3026 16738
rect 3092 16716 3122 16738
rect 3188 16716 3218 16738
rect 3284 16716 3314 16738
rect 3380 16716 3410 16738
rect 2450 16696 3476 16716
rect 2450 16662 2466 16696
rect 2500 16662 2658 16696
rect 2692 16662 2850 16696
rect 2884 16662 3042 16696
rect 3076 16662 3234 16696
rect 3268 16662 3426 16696
rect 3460 16662 3476 16696
rect 2450 16650 3476 16662
rect 3693 16720 3723 16746
rect 4037 16716 4067 16738
rect 4133 16716 4163 16738
rect 4229 16716 4259 16738
rect 4325 16716 4355 16738
rect 4421 16716 4451 16738
rect 4517 16716 4547 16738
rect 4613 16716 4643 16738
rect 4709 16716 4739 16738
rect 4805 16716 4835 16738
rect 4901 16716 4931 16738
rect 3971 16696 4997 16716
rect 3971 16662 3987 16696
rect 4021 16662 4179 16696
rect 4213 16662 4371 16696
rect 4405 16662 4563 16696
rect 4597 16662 4755 16696
rect 4789 16662 4947 16696
rect 4981 16662 4997 16696
rect 3971 16650 4997 16662
rect 5400 16733 5430 16759
rect 297 16213 1323 16229
rect 297 16179 313 16213
rect 347 16179 505 16213
rect 539 16179 697 16213
rect 731 16179 889 16213
rect 923 16179 1081 16213
rect 1115 16179 1273 16213
rect 1307 16179 1323 16213
rect 297 16163 1323 16179
rect 363 16131 393 16163
rect 459 16131 489 16163
rect 555 16131 585 16163
rect 651 16131 681 16163
rect 747 16131 777 16163
rect 843 16131 873 16163
rect 939 16131 969 16163
rect 1035 16131 1065 16163
rect 1131 16131 1161 16163
rect 1227 16131 1257 16163
rect 363 15833 393 15859
rect 459 15833 489 15859
rect 555 15833 585 15859
rect 651 15833 681 15859
rect 747 15833 777 15859
rect 843 15833 873 15859
rect 939 15833 969 15859
rect 1035 15833 1065 15859
rect 1131 15833 1161 15859
rect 1227 15833 1257 15859
rect 2450 16217 3476 16233
rect 2450 16183 2466 16217
rect 2500 16183 2658 16217
rect 2692 16183 2850 16217
rect 2884 16183 3042 16217
rect 3076 16183 3234 16217
rect 3268 16183 3426 16217
rect 3460 16183 3476 16217
rect 2450 16167 3476 16183
rect 2516 16135 2546 16167
rect 2612 16135 2642 16167
rect 2708 16135 2738 16167
rect 2804 16135 2834 16167
rect 2900 16135 2930 16167
rect 2996 16135 3026 16167
rect 3092 16135 3122 16167
rect 3188 16135 3218 16167
rect 3284 16135 3314 16167
rect 3380 16135 3410 16167
rect 2516 15837 2546 15863
rect 2612 15837 2642 15863
rect 2708 15837 2738 15863
rect 2804 15837 2834 15863
rect 2900 15837 2930 15863
rect 2996 15837 3026 15863
rect 3092 15837 3122 15863
rect 3188 15837 3218 15863
rect 3284 15837 3314 15863
rect 3380 15837 3410 15863
rect 3971 16217 4997 16233
rect 3971 16183 3987 16217
rect 4021 16183 4179 16217
rect 4213 16183 4371 16217
rect 4405 16183 4563 16217
rect 4597 16183 4755 16217
rect 4789 16183 4947 16217
rect 4981 16183 4997 16217
rect 3971 16167 4997 16183
rect 4037 16135 4067 16167
rect 4133 16135 4163 16167
rect 4229 16135 4259 16167
rect 4325 16135 4355 16167
rect 4421 16135 4451 16167
rect 4517 16135 4547 16167
rect 4613 16135 4643 16167
rect 4709 16135 4739 16167
rect 4805 16135 4835 16167
rect 4901 16135 4931 16167
rect 5400 15922 5430 15948
rect 4037 15837 4067 15863
rect 4133 15837 4163 15863
rect 4229 15837 4259 15863
rect 4325 15837 4355 15863
rect 4421 15837 4451 15863
rect 4517 15837 4547 15863
rect 4613 15837 4643 15863
rect 4709 15837 4739 15863
rect 4805 15837 4835 15863
rect 4901 15837 4931 15863
rect 5400 15690 5430 15722
rect 5400 15674 5486 15690
rect 363 15551 393 15577
rect 459 15551 489 15577
rect 555 15551 585 15577
rect 651 15551 681 15577
rect 747 15551 777 15577
rect 843 15551 873 15577
rect 939 15551 969 15577
rect 1035 15551 1065 15577
rect 1131 15551 1161 15577
rect 1227 15551 1257 15577
rect 363 15425 393 15447
rect 459 15425 489 15447
rect 555 15425 585 15447
rect 651 15425 681 15447
rect 747 15425 777 15447
rect 843 15425 873 15447
rect 939 15425 969 15447
rect 1035 15425 1065 15447
rect 1131 15425 1161 15447
rect 1227 15425 1257 15447
rect 297 15405 1323 15425
rect 297 15371 313 15405
rect 347 15371 505 15405
rect 539 15371 697 15405
rect 731 15371 889 15405
rect 923 15371 1081 15405
rect 1115 15371 1273 15405
rect 1307 15371 1323 15405
rect 297 15359 1323 15371
rect 2516 15555 2546 15581
rect 2612 15555 2642 15581
rect 2708 15555 2738 15581
rect 2804 15555 2834 15581
rect 2900 15555 2930 15581
rect 2996 15555 3026 15581
rect 3092 15555 3122 15581
rect 3188 15555 3218 15581
rect 3284 15555 3314 15581
rect 3380 15555 3410 15581
rect 3675 15631 3741 15647
rect 3675 15597 3691 15631
rect 3725 15597 3741 15631
rect 3675 15581 3741 15597
rect 3693 15559 3723 15581
rect 4037 15555 4067 15581
rect 4133 15555 4163 15581
rect 4229 15555 4259 15581
rect 4325 15555 4355 15581
rect 4421 15555 4451 15581
rect 4517 15555 4547 15581
rect 4613 15555 4643 15581
rect 4709 15555 4739 15581
rect 4805 15555 4835 15581
rect 4901 15555 4931 15581
rect 5400 15640 5436 15674
rect 5470 15640 5486 15674
rect 5400 15624 5486 15640
rect 5400 15602 5430 15624
rect 2516 15429 2546 15451
rect 2612 15429 2642 15451
rect 2708 15429 2738 15451
rect 2804 15429 2834 15451
rect 2900 15429 2930 15451
rect 2996 15429 3026 15451
rect 3092 15429 3122 15451
rect 3188 15429 3218 15451
rect 3284 15429 3314 15451
rect 3380 15429 3410 15451
rect 2450 15409 3476 15429
rect 2450 15375 2466 15409
rect 2500 15375 2658 15409
rect 2692 15375 2850 15409
rect 2884 15375 3042 15409
rect 3076 15375 3234 15409
rect 3268 15375 3426 15409
rect 3460 15375 3476 15409
rect 2450 15363 3476 15375
rect 3693 15433 3723 15459
rect 4037 15429 4067 15451
rect 4133 15429 4163 15451
rect 4229 15429 4259 15451
rect 4325 15429 4355 15451
rect 4421 15429 4451 15451
rect 4517 15429 4547 15451
rect 4613 15429 4643 15451
rect 4709 15429 4739 15451
rect 4805 15429 4835 15451
rect 4901 15429 4931 15451
rect 3971 15409 4997 15429
rect 3971 15375 3987 15409
rect 4021 15375 4179 15409
rect 4213 15375 4371 15409
rect 4405 15375 4563 15409
rect 4597 15375 4755 15409
rect 4789 15375 4947 15409
rect 4981 15375 4997 15409
rect 3971 15363 4997 15375
rect 5400 15446 5430 15472
rect 297 14926 1323 14942
rect 297 14892 313 14926
rect 347 14892 505 14926
rect 539 14892 697 14926
rect 731 14892 889 14926
rect 923 14892 1081 14926
rect 1115 14892 1273 14926
rect 1307 14892 1323 14926
rect 297 14876 1323 14892
rect 363 14844 393 14876
rect 459 14844 489 14876
rect 555 14844 585 14876
rect 651 14844 681 14876
rect 747 14844 777 14876
rect 843 14844 873 14876
rect 939 14844 969 14876
rect 1035 14844 1065 14876
rect 1131 14844 1161 14876
rect 1227 14844 1257 14876
rect 363 14546 393 14572
rect 459 14546 489 14572
rect 555 14546 585 14572
rect 651 14546 681 14572
rect 747 14546 777 14572
rect 843 14546 873 14572
rect 939 14546 969 14572
rect 1035 14546 1065 14572
rect 1131 14546 1161 14572
rect 1227 14546 1257 14572
rect 2450 14930 3476 14946
rect 2450 14896 2466 14930
rect 2500 14896 2658 14930
rect 2692 14896 2850 14930
rect 2884 14896 3042 14930
rect 3076 14896 3234 14930
rect 3268 14896 3426 14930
rect 3460 14896 3476 14930
rect 2450 14880 3476 14896
rect 2516 14848 2546 14880
rect 2612 14848 2642 14880
rect 2708 14848 2738 14880
rect 2804 14848 2834 14880
rect 2900 14848 2930 14880
rect 2996 14848 3026 14880
rect 3092 14848 3122 14880
rect 3188 14848 3218 14880
rect 3284 14848 3314 14880
rect 3380 14848 3410 14880
rect 2516 14550 2546 14576
rect 2612 14550 2642 14576
rect 2708 14550 2738 14576
rect 2804 14550 2834 14576
rect 2900 14550 2930 14576
rect 2996 14550 3026 14576
rect 3092 14550 3122 14576
rect 3188 14550 3218 14576
rect 3284 14550 3314 14576
rect 3380 14550 3410 14576
rect 3971 14930 4997 14946
rect 3971 14896 3987 14930
rect 4021 14896 4179 14930
rect 4213 14896 4371 14930
rect 4405 14896 4563 14930
rect 4597 14896 4755 14930
rect 4789 14896 4947 14930
rect 4981 14896 4997 14930
rect 3971 14880 4997 14896
rect 4037 14848 4067 14880
rect 4133 14848 4163 14880
rect 4229 14848 4259 14880
rect 4325 14848 4355 14880
rect 4421 14848 4451 14880
rect 4517 14848 4547 14880
rect 4613 14848 4643 14880
rect 4709 14848 4739 14880
rect 4805 14848 4835 14880
rect 4901 14848 4931 14880
rect 5400 14635 5430 14661
rect 4037 14550 4067 14576
rect 4133 14550 4163 14576
rect 4229 14550 4259 14576
rect 4325 14550 4355 14576
rect 4421 14550 4451 14576
rect 4517 14550 4547 14576
rect 4613 14550 4643 14576
rect 4709 14550 4739 14576
rect 4805 14550 4835 14576
rect 4901 14550 4931 14576
rect 5400 14403 5430 14435
rect 5400 14387 5486 14403
rect 363 14264 393 14290
rect 459 14264 489 14290
rect 555 14264 585 14290
rect 651 14264 681 14290
rect 747 14264 777 14290
rect 843 14264 873 14290
rect 939 14264 969 14290
rect 1035 14264 1065 14290
rect 1131 14264 1161 14290
rect 1227 14264 1257 14290
rect 363 14138 393 14160
rect 459 14138 489 14160
rect 555 14138 585 14160
rect 651 14138 681 14160
rect 747 14138 777 14160
rect 843 14138 873 14160
rect 939 14138 969 14160
rect 1035 14138 1065 14160
rect 1131 14138 1161 14160
rect 1227 14138 1257 14160
rect 297 14118 1323 14138
rect 297 14084 313 14118
rect 347 14084 505 14118
rect 539 14084 697 14118
rect 731 14084 889 14118
rect 923 14084 1081 14118
rect 1115 14084 1273 14118
rect 1307 14084 1323 14118
rect 297 14072 1323 14084
rect 2516 14268 2546 14294
rect 2612 14268 2642 14294
rect 2708 14268 2738 14294
rect 2804 14268 2834 14294
rect 2900 14268 2930 14294
rect 2996 14268 3026 14294
rect 3092 14268 3122 14294
rect 3188 14268 3218 14294
rect 3284 14268 3314 14294
rect 3380 14268 3410 14294
rect 3675 14344 3741 14360
rect 3675 14310 3691 14344
rect 3725 14310 3741 14344
rect 3675 14294 3741 14310
rect 3693 14272 3723 14294
rect 4037 14268 4067 14294
rect 4133 14268 4163 14294
rect 4229 14268 4259 14294
rect 4325 14268 4355 14294
rect 4421 14268 4451 14294
rect 4517 14268 4547 14294
rect 4613 14268 4643 14294
rect 4709 14268 4739 14294
rect 4805 14268 4835 14294
rect 4901 14268 4931 14294
rect 5400 14353 5436 14387
rect 5470 14353 5486 14387
rect 5400 14337 5486 14353
rect 5400 14315 5430 14337
rect 2516 14142 2546 14164
rect 2612 14142 2642 14164
rect 2708 14142 2738 14164
rect 2804 14142 2834 14164
rect 2900 14142 2930 14164
rect 2996 14142 3026 14164
rect 3092 14142 3122 14164
rect 3188 14142 3218 14164
rect 3284 14142 3314 14164
rect 3380 14142 3410 14164
rect 2450 14122 3476 14142
rect 2450 14088 2466 14122
rect 2500 14088 2658 14122
rect 2692 14088 2850 14122
rect 2884 14088 3042 14122
rect 3076 14088 3234 14122
rect 3268 14088 3426 14122
rect 3460 14088 3476 14122
rect 2450 14076 3476 14088
rect 3693 14146 3723 14172
rect 4037 14142 4067 14164
rect 4133 14142 4163 14164
rect 4229 14142 4259 14164
rect 4325 14142 4355 14164
rect 4421 14142 4451 14164
rect 4517 14142 4547 14164
rect 4613 14142 4643 14164
rect 4709 14142 4739 14164
rect 4805 14142 4835 14164
rect 4901 14142 4931 14164
rect 3971 14122 4997 14142
rect 3971 14088 3987 14122
rect 4021 14088 4179 14122
rect 4213 14088 4371 14122
rect 4405 14088 4563 14122
rect 4597 14088 4755 14122
rect 4789 14088 4947 14122
rect 4981 14088 4997 14122
rect 3971 14076 4997 14088
rect 5400 14159 5430 14185
rect 297 13639 1323 13655
rect 297 13605 313 13639
rect 347 13605 505 13639
rect 539 13605 697 13639
rect 731 13605 889 13639
rect 923 13605 1081 13639
rect 1115 13605 1273 13639
rect 1307 13605 1323 13639
rect 297 13589 1323 13605
rect 363 13557 393 13589
rect 459 13557 489 13589
rect 555 13557 585 13589
rect 651 13557 681 13589
rect 747 13557 777 13589
rect 843 13557 873 13589
rect 939 13557 969 13589
rect 1035 13557 1065 13589
rect 1131 13557 1161 13589
rect 1227 13557 1257 13589
rect 363 13259 393 13285
rect 459 13259 489 13285
rect 555 13259 585 13285
rect 651 13259 681 13285
rect 747 13259 777 13285
rect 843 13259 873 13285
rect 939 13259 969 13285
rect 1035 13259 1065 13285
rect 1131 13259 1161 13285
rect 1227 13259 1257 13285
rect 2450 13643 3476 13659
rect 2450 13609 2466 13643
rect 2500 13609 2658 13643
rect 2692 13609 2850 13643
rect 2884 13609 3042 13643
rect 3076 13609 3234 13643
rect 3268 13609 3426 13643
rect 3460 13609 3476 13643
rect 2450 13593 3476 13609
rect 2516 13561 2546 13593
rect 2612 13561 2642 13593
rect 2708 13561 2738 13593
rect 2804 13561 2834 13593
rect 2900 13561 2930 13593
rect 2996 13561 3026 13593
rect 3092 13561 3122 13593
rect 3188 13561 3218 13593
rect 3284 13561 3314 13593
rect 3380 13561 3410 13593
rect 2516 13263 2546 13289
rect 2612 13263 2642 13289
rect 2708 13263 2738 13289
rect 2804 13263 2834 13289
rect 2900 13263 2930 13289
rect 2996 13263 3026 13289
rect 3092 13263 3122 13289
rect 3188 13263 3218 13289
rect 3284 13263 3314 13289
rect 3380 13263 3410 13289
rect 3971 13643 4997 13659
rect 3971 13609 3987 13643
rect 4021 13609 4179 13643
rect 4213 13609 4371 13643
rect 4405 13609 4563 13643
rect 4597 13609 4755 13643
rect 4789 13609 4947 13643
rect 4981 13609 4997 13643
rect 3971 13593 4997 13609
rect 4037 13561 4067 13593
rect 4133 13561 4163 13593
rect 4229 13561 4259 13593
rect 4325 13561 4355 13593
rect 4421 13561 4451 13593
rect 4517 13561 4547 13593
rect 4613 13561 4643 13593
rect 4709 13561 4739 13593
rect 4805 13561 4835 13593
rect 4901 13561 4931 13593
rect 5400 13348 5430 13374
rect 4037 13263 4067 13289
rect 4133 13263 4163 13289
rect 4229 13263 4259 13289
rect 4325 13263 4355 13289
rect 4421 13263 4451 13289
rect 4517 13263 4547 13289
rect 4613 13263 4643 13289
rect 4709 13263 4739 13289
rect 4805 13263 4835 13289
rect 4901 13263 4931 13289
rect 5400 13116 5430 13148
rect 5400 13100 5486 13116
rect 363 12977 393 13003
rect 459 12977 489 13003
rect 555 12977 585 13003
rect 651 12977 681 13003
rect 747 12977 777 13003
rect 843 12977 873 13003
rect 939 12977 969 13003
rect 1035 12977 1065 13003
rect 1131 12977 1161 13003
rect 1227 12977 1257 13003
rect 363 12851 393 12873
rect 459 12851 489 12873
rect 555 12851 585 12873
rect 651 12851 681 12873
rect 747 12851 777 12873
rect 843 12851 873 12873
rect 939 12851 969 12873
rect 1035 12851 1065 12873
rect 1131 12851 1161 12873
rect 1227 12851 1257 12873
rect 297 12831 1323 12851
rect 297 12797 313 12831
rect 347 12797 505 12831
rect 539 12797 697 12831
rect 731 12797 889 12831
rect 923 12797 1081 12831
rect 1115 12797 1273 12831
rect 1307 12797 1323 12831
rect 297 12785 1323 12797
rect 2516 12981 2546 13007
rect 2612 12981 2642 13007
rect 2708 12981 2738 13007
rect 2804 12981 2834 13007
rect 2900 12981 2930 13007
rect 2996 12981 3026 13007
rect 3092 12981 3122 13007
rect 3188 12981 3218 13007
rect 3284 12981 3314 13007
rect 3380 12981 3410 13007
rect 3675 13057 3741 13073
rect 3675 13023 3691 13057
rect 3725 13023 3741 13057
rect 3675 13007 3741 13023
rect 3693 12985 3723 13007
rect 4037 12981 4067 13007
rect 4133 12981 4163 13007
rect 4229 12981 4259 13007
rect 4325 12981 4355 13007
rect 4421 12981 4451 13007
rect 4517 12981 4547 13007
rect 4613 12981 4643 13007
rect 4709 12981 4739 13007
rect 4805 12981 4835 13007
rect 4901 12981 4931 13007
rect 5400 13066 5436 13100
rect 5470 13066 5486 13100
rect 5400 13050 5486 13066
rect 5400 13028 5430 13050
rect 2516 12855 2546 12877
rect 2612 12855 2642 12877
rect 2708 12855 2738 12877
rect 2804 12855 2834 12877
rect 2900 12855 2930 12877
rect 2996 12855 3026 12877
rect 3092 12855 3122 12877
rect 3188 12855 3218 12877
rect 3284 12855 3314 12877
rect 3380 12855 3410 12877
rect 2450 12835 3476 12855
rect 2450 12801 2466 12835
rect 2500 12801 2658 12835
rect 2692 12801 2850 12835
rect 2884 12801 3042 12835
rect 3076 12801 3234 12835
rect 3268 12801 3426 12835
rect 3460 12801 3476 12835
rect 2450 12789 3476 12801
rect 3693 12859 3723 12885
rect 4037 12855 4067 12877
rect 4133 12855 4163 12877
rect 4229 12855 4259 12877
rect 4325 12855 4355 12877
rect 4421 12855 4451 12877
rect 4517 12855 4547 12877
rect 4613 12855 4643 12877
rect 4709 12855 4739 12877
rect 4805 12855 4835 12877
rect 4901 12855 4931 12877
rect 3971 12835 4997 12855
rect 3971 12801 3987 12835
rect 4021 12801 4179 12835
rect 4213 12801 4371 12835
rect 4405 12801 4563 12835
rect 4597 12801 4755 12835
rect 4789 12801 4947 12835
rect 4981 12801 4997 12835
rect 3971 12789 4997 12801
rect 5400 12872 5430 12898
rect 297 12352 1323 12368
rect 297 12318 313 12352
rect 347 12318 505 12352
rect 539 12318 697 12352
rect 731 12318 889 12352
rect 923 12318 1081 12352
rect 1115 12318 1273 12352
rect 1307 12318 1323 12352
rect 297 12302 1323 12318
rect 363 12270 393 12302
rect 459 12270 489 12302
rect 555 12270 585 12302
rect 651 12270 681 12302
rect 747 12270 777 12302
rect 843 12270 873 12302
rect 939 12270 969 12302
rect 1035 12270 1065 12302
rect 1131 12270 1161 12302
rect 1227 12270 1257 12302
rect 363 11972 393 11998
rect 459 11972 489 11998
rect 555 11972 585 11998
rect 651 11972 681 11998
rect 747 11972 777 11998
rect 843 11972 873 11998
rect 939 11972 969 11998
rect 1035 11972 1065 11998
rect 1131 11972 1161 11998
rect 1227 11972 1257 11998
rect 2450 12356 3476 12372
rect 2450 12322 2466 12356
rect 2500 12322 2658 12356
rect 2692 12322 2850 12356
rect 2884 12322 3042 12356
rect 3076 12322 3234 12356
rect 3268 12322 3426 12356
rect 3460 12322 3476 12356
rect 2450 12306 3476 12322
rect 2516 12274 2546 12306
rect 2612 12274 2642 12306
rect 2708 12274 2738 12306
rect 2804 12274 2834 12306
rect 2900 12274 2930 12306
rect 2996 12274 3026 12306
rect 3092 12274 3122 12306
rect 3188 12274 3218 12306
rect 3284 12274 3314 12306
rect 3380 12274 3410 12306
rect 2516 11976 2546 12002
rect 2612 11976 2642 12002
rect 2708 11976 2738 12002
rect 2804 11976 2834 12002
rect 2900 11976 2930 12002
rect 2996 11976 3026 12002
rect 3092 11976 3122 12002
rect 3188 11976 3218 12002
rect 3284 11976 3314 12002
rect 3380 11976 3410 12002
rect 3971 12356 4997 12372
rect 3971 12322 3987 12356
rect 4021 12322 4179 12356
rect 4213 12322 4371 12356
rect 4405 12322 4563 12356
rect 4597 12322 4755 12356
rect 4789 12322 4947 12356
rect 4981 12322 4997 12356
rect 3971 12306 4997 12322
rect 4037 12274 4067 12306
rect 4133 12274 4163 12306
rect 4229 12274 4259 12306
rect 4325 12274 4355 12306
rect 4421 12274 4451 12306
rect 4517 12274 4547 12306
rect 4613 12274 4643 12306
rect 4709 12274 4739 12306
rect 4805 12274 4835 12306
rect 4901 12274 4931 12306
rect 5400 12061 5430 12087
rect 4037 11976 4067 12002
rect 4133 11976 4163 12002
rect 4229 11976 4259 12002
rect 4325 11976 4355 12002
rect 4421 11976 4451 12002
rect 4517 11976 4547 12002
rect 4613 11976 4643 12002
rect 4709 11976 4739 12002
rect 4805 11976 4835 12002
rect 4901 11976 4931 12002
rect 5400 11829 5430 11861
rect 5400 11813 5486 11829
rect 363 11690 393 11716
rect 459 11690 489 11716
rect 555 11690 585 11716
rect 651 11690 681 11716
rect 747 11690 777 11716
rect 843 11690 873 11716
rect 939 11690 969 11716
rect 1035 11690 1065 11716
rect 1131 11690 1161 11716
rect 1227 11690 1257 11716
rect 363 11564 393 11586
rect 459 11564 489 11586
rect 555 11564 585 11586
rect 651 11564 681 11586
rect 747 11564 777 11586
rect 843 11564 873 11586
rect 939 11564 969 11586
rect 1035 11564 1065 11586
rect 1131 11564 1161 11586
rect 1227 11564 1257 11586
rect 297 11544 1323 11564
rect 297 11510 313 11544
rect 347 11510 505 11544
rect 539 11510 697 11544
rect 731 11510 889 11544
rect 923 11510 1081 11544
rect 1115 11510 1273 11544
rect 1307 11510 1323 11544
rect 297 11498 1323 11510
rect 2516 11694 2546 11720
rect 2612 11694 2642 11720
rect 2708 11694 2738 11720
rect 2804 11694 2834 11720
rect 2900 11694 2930 11720
rect 2996 11694 3026 11720
rect 3092 11694 3122 11720
rect 3188 11694 3218 11720
rect 3284 11694 3314 11720
rect 3380 11694 3410 11720
rect 3675 11770 3741 11786
rect 3675 11736 3691 11770
rect 3725 11736 3741 11770
rect 3675 11720 3741 11736
rect 3693 11698 3723 11720
rect 4037 11694 4067 11720
rect 4133 11694 4163 11720
rect 4229 11694 4259 11720
rect 4325 11694 4355 11720
rect 4421 11694 4451 11720
rect 4517 11694 4547 11720
rect 4613 11694 4643 11720
rect 4709 11694 4739 11720
rect 4805 11694 4835 11720
rect 4901 11694 4931 11720
rect 5400 11779 5436 11813
rect 5470 11779 5486 11813
rect 5400 11763 5486 11779
rect 5400 11741 5430 11763
rect 2516 11568 2546 11590
rect 2612 11568 2642 11590
rect 2708 11568 2738 11590
rect 2804 11568 2834 11590
rect 2900 11568 2930 11590
rect 2996 11568 3026 11590
rect 3092 11568 3122 11590
rect 3188 11568 3218 11590
rect 3284 11568 3314 11590
rect 3380 11568 3410 11590
rect 2450 11548 3476 11568
rect 2450 11514 2466 11548
rect 2500 11514 2658 11548
rect 2692 11514 2850 11548
rect 2884 11514 3042 11548
rect 3076 11514 3234 11548
rect 3268 11514 3426 11548
rect 3460 11514 3476 11548
rect 2450 11502 3476 11514
rect 3693 11572 3723 11598
rect 4037 11568 4067 11590
rect 4133 11568 4163 11590
rect 4229 11568 4259 11590
rect 4325 11568 4355 11590
rect 4421 11568 4451 11590
rect 4517 11568 4547 11590
rect 4613 11568 4643 11590
rect 4709 11568 4739 11590
rect 4805 11568 4835 11590
rect 4901 11568 4931 11590
rect 3971 11548 4997 11568
rect 3971 11514 3987 11548
rect 4021 11514 4179 11548
rect 4213 11514 4371 11548
rect 4405 11514 4563 11548
rect 4597 11514 4755 11548
rect 4789 11514 4947 11548
rect 4981 11514 4997 11548
rect 3971 11502 4997 11514
rect 5400 11585 5430 11611
rect 297 11065 1323 11081
rect 297 11031 313 11065
rect 347 11031 505 11065
rect 539 11031 697 11065
rect 731 11031 889 11065
rect 923 11031 1081 11065
rect 1115 11031 1273 11065
rect 1307 11031 1323 11065
rect 297 11015 1323 11031
rect 363 10983 393 11015
rect 459 10983 489 11015
rect 555 10983 585 11015
rect 651 10983 681 11015
rect 747 10983 777 11015
rect 843 10983 873 11015
rect 939 10983 969 11015
rect 1035 10983 1065 11015
rect 1131 10983 1161 11015
rect 1227 10983 1257 11015
rect 363 10685 393 10711
rect 459 10685 489 10711
rect 555 10685 585 10711
rect 651 10685 681 10711
rect 747 10685 777 10711
rect 843 10685 873 10711
rect 939 10685 969 10711
rect 1035 10685 1065 10711
rect 1131 10685 1161 10711
rect 1227 10685 1257 10711
rect 2450 11069 3476 11085
rect 2450 11035 2466 11069
rect 2500 11035 2658 11069
rect 2692 11035 2850 11069
rect 2884 11035 3042 11069
rect 3076 11035 3234 11069
rect 3268 11035 3426 11069
rect 3460 11035 3476 11069
rect 2450 11019 3476 11035
rect 2516 10987 2546 11019
rect 2612 10987 2642 11019
rect 2708 10987 2738 11019
rect 2804 10987 2834 11019
rect 2900 10987 2930 11019
rect 2996 10987 3026 11019
rect 3092 10987 3122 11019
rect 3188 10987 3218 11019
rect 3284 10987 3314 11019
rect 3380 10987 3410 11019
rect 2516 10689 2546 10715
rect 2612 10689 2642 10715
rect 2708 10689 2738 10715
rect 2804 10689 2834 10715
rect 2900 10689 2930 10715
rect 2996 10689 3026 10715
rect 3092 10689 3122 10715
rect 3188 10689 3218 10715
rect 3284 10689 3314 10715
rect 3380 10689 3410 10715
rect 3971 11069 4997 11085
rect 3971 11035 3987 11069
rect 4021 11035 4179 11069
rect 4213 11035 4371 11069
rect 4405 11035 4563 11069
rect 4597 11035 4755 11069
rect 4789 11035 4947 11069
rect 4981 11035 4997 11069
rect 3971 11019 4997 11035
rect 4037 10987 4067 11019
rect 4133 10987 4163 11019
rect 4229 10987 4259 11019
rect 4325 10987 4355 11019
rect 4421 10987 4451 11019
rect 4517 10987 4547 11019
rect 4613 10987 4643 11019
rect 4709 10987 4739 11019
rect 4805 10987 4835 11019
rect 4901 10987 4931 11019
rect 5400 10774 5430 10800
rect 4037 10689 4067 10715
rect 4133 10689 4163 10715
rect 4229 10689 4259 10715
rect 4325 10689 4355 10715
rect 4421 10689 4451 10715
rect 4517 10689 4547 10715
rect 4613 10689 4643 10715
rect 4709 10689 4739 10715
rect 4805 10689 4835 10715
rect 4901 10689 4931 10715
rect 5400 10542 5430 10574
rect 5400 10526 5486 10542
rect 363 10403 393 10429
rect 459 10403 489 10429
rect 555 10403 585 10429
rect 651 10403 681 10429
rect 747 10403 777 10429
rect 843 10403 873 10429
rect 939 10403 969 10429
rect 1035 10403 1065 10429
rect 1131 10403 1161 10429
rect 1227 10403 1257 10429
rect 363 10277 393 10299
rect 459 10277 489 10299
rect 555 10277 585 10299
rect 651 10277 681 10299
rect 747 10277 777 10299
rect 843 10277 873 10299
rect 939 10277 969 10299
rect 1035 10277 1065 10299
rect 1131 10277 1161 10299
rect 1227 10277 1257 10299
rect 297 10257 1323 10277
rect 297 10223 313 10257
rect 347 10223 505 10257
rect 539 10223 697 10257
rect 731 10223 889 10257
rect 923 10223 1081 10257
rect 1115 10223 1273 10257
rect 1307 10223 1323 10257
rect 297 10211 1323 10223
rect 2516 10407 2546 10433
rect 2612 10407 2642 10433
rect 2708 10407 2738 10433
rect 2804 10407 2834 10433
rect 2900 10407 2930 10433
rect 2996 10407 3026 10433
rect 3092 10407 3122 10433
rect 3188 10407 3218 10433
rect 3284 10407 3314 10433
rect 3380 10407 3410 10433
rect 3675 10483 3741 10499
rect 3675 10449 3691 10483
rect 3725 10449 3741 10483
rect 3675 10433 3741 10449
rect 3693 10411 3723 10433
rect 4037 10407 4067 10433
rect 4133 10407 4163 10433
rect 4229 10407 4259 10433
rect 4325 10407 4355 10433
rect 4421 10407 4451 10433
rect 4517 10407 4547 10433
rect 4613 10407 4643 10433
rect 4709 10407 4739 10433
rect 4805 10407 4835 10433
rect 4901 10407 4931 10433
rect 5400 10492 5436 10526
rect 5470 10492 5486 10526
rect 5400 10476 5486 10492
rect 5400 10454 5430 10476
rect 2516 10281 2546 10303
rect 2612 10281 2642 10303
rect 2708 10281 2738 10303
rect 2804 10281 2834 10303
rect 2900 10281 2930 10303
rect 2996 10281 3026 10303
rect 3092 10281 3122 10303
rect 3188 10281 3218 10303
rect 3284 10281 3314 10303
rect 3380 10281 3410 10303
rect 2450 10261 3476 10281
rect 2450 10227 2466 10261
rect 2500 10227 2658 10261
rect 2692 10227 2850 10261
rect 2884 10227 3042 10261
rect 3076 10227 3234 10261
rect 3268 10227 3426 10261
rect 3460 10227 3476 10261
rect 2450 10215 3476 10227
rect 3693 10285 3723 10311
rect 4037 10281 4067 10303
rect 4133 10281 4163 10303
rect 4229 10281 4259 10303
rect 4325 10281 4355 10303
rect 4421 10281 4451 10303
rect 4517 10281 4547 10303
rect 4613 10281 4643 10303
rect 4709 10281 4739 10303
rect 4805 10281 4835 10303
rect 4901 10281 4931 10303
rect 3971 10261 4997 10281
rect 3971 10227 3987 10261
rect 4021 10227 4179 10261
rect 4213 10227 4371 10261
rect 4405 10227 4563 10261
rect 4597 10227 4755 10261
rect 4789 10227 4947 10261
rect 4981 10227 4997 10261
rect 3971 10215 4997 10227
rect 5400 10298 5430 10324
rect 297 9778 1323 9794
rect 297 9744 313 9778
rect 347 9744 505 9778
rect 539 9744 697 9778
rect 731 9744 889 9778
rect 923 9744 1081 9778
rect 1115 9744 1273 9778
rect 1307 9744 1323 9778
rect 297 9728 1323 9744
rect 363 9696 393 9728
rect 459 9696 489 9728
rect 555 9696 585 9728
rect 651 9696 681 9728
rect 747 9696 777 9728
rect 843 9696 873 9728
rect 939 9696 969 9728
rect 1035 9696 1065 9728
rect 1131 9696 1161 9728
rect 1227 9696 1257 9728
rect 363 9398 393 9424
rect 459 9398 489 9424
rect 555 9398 585 9424
rect 651 9398 681 9424
rect 747 9398 777 9424
rect 843 9398 873 9424
rect 939 9398 969 9424
rect 1035 9398 1065 9424
rect 1131 9398 1161 9424
rect 1227 9398 1257 9424
rect 2450 9782 3476 9798
rect 2450 9748 2466 9782
rect 2500 9748 2658 9782
rect 2692 9748 2850 9782
rect 2884 9748 3042 9782
rect 3076 9748 3234 9782
rect 3268 9748 3426 9782
rect 3460 9748 3476 9782
rect 2450 9732 3476 9748
rect 2516 9700 2546 9732
rect 2612 9700 2642 9732
rect 2708 9700 2738 9732
rect 2804 9700 2834 9732
rect 2900 9700 2930 9732
rect 2996 9700 3026 9732
rect 3092 9700 3122 9732
rect 3188 9700 3218 9732
rect 3284 9700 3314 9732
rect 3380 9700 3410 9732
rect 2516 9402 2546 9428
rect 2612 9402 2642 9428
rect 2708 9402 2738 9428
rect 2804 9402 2834 9428
rect 2900 9402 2930 9428
rect 2996 9402 3026 9428
rect 3092 9402 3122 9428
rect 3188 9402 3218 9428
rect 3284 9402 3314 9428
rect 3380 9402 3410 9428
rect 3971 9782 4997 9798
rect 3971 9748 3987 9782
rect 4021 9748 4179 9782
rect 4213 9748 4371 9782
rect 4405 9748 4563 9782
rect 4597 9748 4755 9782
rect 4789 9748 4947 9782
rect 4981 9748 4997 9782
rect 3971 9732 4997 9748
rect 4037 9700 4067 9732
rect 4133 9700 4163 9732
rect 4229 9700 4259 9732
rect 4325 9700 4355 9732
rect 4421 9700 4451 9732
rect 4517 9700 4547 9732
rect 4613 9700 4643 9732
rect 4709 9700 4739 9732
rect 4805 9700 4835 9732
rect 4901 9700 4931 9732
rect 5400 9487 5430 9513
rect 4037 9402 4067 9428
rect 4133 9402 4163 9428
rect 4229 9402 4259 9428
rect 4325 9402 4355 9428
rect 4421 9402 4451 9428
rect 4517 9402 4547 9428
rect 4613 9402 4643 9428
rect 4709 9402 4739 9428
rect 4805 9402 4835 9428
rect 4901 9402 4931 9428
rect 5400 9255 5430 9287
rect 5400 9239 5486 9255
rect 363 9116 393 9142
rect 459 9116 489 9142
rect 555 9116 585 9142
rect 651 9116 681 9142
rect 747 9116 777 9142
rect 843 9116 873 9142
rect 939 9116 969 9142
rect 1035 9116 1065 9142
rect 1131 9116 1161 9142
rect 1227 9116 1257 9142
rect 363 8990 393 9012
rect 459 8990 489 9012
rect 555 8990 585 9012
rect 651 8990 681 9012
rect 747 8990 777 9012
rect 843 8990 873 9012
rect 939 8990 969 9012
rect 1035 8990 1065 9012
rect 1131 8990 1161 9012
rect 1227 8990 1257 9012
rect 297 8970 1323 8990
rect 297 8936 313 8970
rect 347 8936 505 8970
rect 539 8936 697 8970
rect 731 8936 889 8970
rect 923 8936 1081 8970
rect 1115 8936 1273 8970
rect 1307 8936 1323 8970
rect 297 8924 1323 8936
rect 2516 9120 2546 9146
rect 2612 9120 2642 9146
rect 2708 9120 2738 9146
rect 2804 9120 2834 9146
rect 2900 9120 2930 9146
rect 2996 9120 3026 9146
rect 3092 9120 3122 9146
rect 3188 9120 3218 9146
rect 3284 9120 3314 9146
rect 3380 9120 3410 9146
rect 3675 9196 3741 9212
rect 3675 9162 3691 9196
rect 3725 9162 3741 9196
rect 3675 9146 3741 9162
rect 3693 9124 3723 9146
rect 4037 9120 4067 9146
rect 4133 9120 4163 9146
rect 4229 9120 4259 9146
rect 4325 9120 4355 9146
rect 4421 9120 4451 9146
rect 4517 9120 4547 9146
rect 4613 9120 4643 9146
rect 4709 9120 4739 9146
rect 4805 9120 4835 9146
rect 4901 9120 4931 9146
rect 5400 9205 5436 9239
rect 5470 9205 5486 9239
rect 5400 9189 5486 9205
rect 5400 9167 5430 9189
rect 2516 8994 2546 9016
rect 2612 8994 2642 9016
rect 2708 8994 2738 9016
rect 2804 8994 2834 9016
rect 2900 8994 2930 9016
rect 2996 8994 3026 9016
rect 3092 8994 3122 9016
rect 3188 8994 3218 9016
rect 3284 8994 3314 9016
rect 3380 8994 3410 9016
rect 2450 8974 3476 8994
rect 2450 8940 2466 8974
rect 2500 8940 2658 8974
rect 2692 8940 2850 8974
rect 2884 8940 3042 8974
rect 3076 8940 3234 8974
rect 3268 8940 3426 8974
rect 3460 8940 3476 8974
rect 2450 8928 3476 8940
rect 3693 8998 3723 9024
rect 4037 8994 4067 9016
rect 4133 8994 4163 9016
rect 4229 8994 4259 9016
rect 4325 8994 4355 9016
rect 4421 8994 4451 9016
rect 4517 8994 4547 9016
rect 4613 8994 4643 9016
rect 4709 8994 4739 9016
rect 4805 8994 4835 9016
rect 4901 8994 4931 9016
rect 3971 8974 4997 8994
rect 3971 8940 3987 8974
rect 4021 8940 4179 8974
rect 4213 8940 4371 8974
rect 4405 8940 4563 8974
rect 4597 8940 4755 8974
rect 4789 8940 4947 8974
rect 4981 8940 4997 8974
rect 3971 8928 4997 8940
rect 5400 9011 5430 9037
rect 297 8491 1323 8507
rect 297 8457 313 8491
rect 347 8457 505 8491
rect 539 8457 697 8491
rect 731 8457 889 8491
rect 923 8457 1081 8491
rect 1115 8457 1273 8491
rect 1307 8457 1323 8491
rect 297 8441 1323 8457
rect 363 8409 393 8441
rect 459 8409 489 8441
rect 555 8409 585 8441
rect 651 8409 681 8441
rect 747 8409 777 8441
rect 843 8409 873 8441
rect 939 8409 969 8441
rect 1035 8409 1065 8441
rect 1131 8409 1161 8441
rect 1227 8409 1257 8441
rect 363 8111 393 8137
rect 459 8111 489 8137
rect 555 8111 585 8137
rect 651 8111 681 8137
rect 747 8111 777 8137
rect 843 8111 873 8137
rect 939 8111 969 8137
rect 1035 8111 1065 8137
rect 1131 8111 1161 8137
rect 1227 8111 1257 8137
rect 2450 8495 3476 8511
rect 2450 8461 2466 8495
rect 2500 8461 2658 8495
rect 2692 8461 2850 8495
rect 2884 8461 3042 8495
rect 3076 8461 3234 8495
rect 3268 8461 3426 8495
rect 3460 8461 3476 8495
rect 2450 8445 3476 8461
rect 2516 8413 2546 8445
rect 2612 8413 2642 8445
rect 2708 8413 2738 8445
rect 2804 8413 2834 8445
rect 2900 8413 2930 8445
rect 2996 8413 3026 8445
rect 3092 8413 3122 8445
rect 3188 8413 3218 8445
rect 3284 8413 3314 8445
rect 3380 8413 3410 8445
rect 2516 8115 2546 8141
rect 2612 8115 2642 8141
rect 2708 8115 2738 8141
rect 2804 8115 2834 8141
rect 2900 8115 2930 8141
rect 2996 8115 3026 8141
rect 3092 8115 3122 8141
rect 3188 8115 3218 8141
rect 3284 8115 3314 8141
rect 3380 8115 3410 8141
rect 3971 8495 4997 8511
rect 3971 8461 3987 8495
rect 4021 8461 4179 8495
rect 4213 8461 4371 8495
rect 4405 8461 4563 8495
rect 4597 8461 4755 8495
rect 4789 8461 4947 8495
rect 4981 8461 4997 8495
rect 3971 8445 4997 8461
rect 4037 8413 4067 8445
rect 4133 8413 4163 8445
rect 4229 8413 4259 8445
rect 4325 8413 4355 8445
rect 4421 8413 4451 8445
rect 4517 8413 4547 8445
rect 4613 8413 4643 8445
rect 4709 8413 4739 8445
rect 4805 8413 4835 8445
rect 4901 8413 4931 8445
rect 5400 8200 5430 8226
rect 4037 8115 4067 8141
rect 4133 8115 4163 8141
rect 4229 8115 4259 8141
rect 4325 8115 4355 8141
rect 4421 8115 4451 8141
rect 4517 8115 4547 8141
rect 4613 8115 4643 8141
rect 4709 8115 4739 8141
rect 4805 8115 4835 8141
rect 4901 8115 4931 8141
rect 5400 7968 5430 8000
rect 5400 7952 5486 7968
rect 363 7829 393 7855
rect 459 7829 489 7855
rect 555 7829 585 7855
rect 651 7829 681 7855
rect 747 7829 777 7855
rect 843 7829 873 7855
rect 939 7829 969 7855
rect 1035 7829 1065 7855
rect 1131 7829 1161 7855
rect 1227 7829 1257 7855
rect 363 7703 393 7725
rect 459 7703 489 7725
rect 555 7703 585 7725
rect 651 7703 681 7725
rect 747 7703 777 7725
rect 843 7703 873 7725
rect 939 7703 969 7725
rect 1035 7703 1065 7725
rect 1131 7703 1161 7725
rect 1227 7703 1257 7725
rect 297 7683 1323 7703
rect 297 7649 313 7683
rect 347 7649 505 7683
rect 539 7649 697 7683
rect 731 7649 889 7683
rect 923 7649 1081 7683
rect 1115 7649 1273 7683
rect 1307 7649 1323 7683
rect 297 7637 1323 7649
rect 2516 7833 2546 7859
rect 2612 7833 2642 7859
rect 2708 7833 2738 7859
rect 2804 7833 2834 7859
rect 2900 7833 2930 7859
rect 2996 7833 3026 7859
rect 3092 7833 3122 7859
rect 3188 7833 3218 7859
rect 3284 7833 3314 7859
rect 3380 7833 3410 7859
rect 3675 7909 3741 7925
rect 3675 7875 3691 7909
rect 3725 7875 3741 7909
rect 3675 7859 3741 7875
rect 3693 7837 3723 7859
rect 4037 7833 4067 7859
rect 4133 7833 4163 7859
rect 4229 7833 4259 7859
rect 4325 7833 4355 7859
rect 4421 7833 4451 7859
rect 4517 7833 4547 7859
rect 4613 7833 4643 7859
rect 4709 7833 4739 7859
rect 4805 7833 4835 7859
rect 4901 7833 4931 7859
rect 5400 7918 5436 7952
rect 5470 7918 5486 7952
rect 5400 7902 5486 7918
rect 5400 7880 5430 7902
rect 2516 7707 2546 7729
rect 2612 7707 2642 7729
rect 2708 7707 2738 7729
rect 2804 7707 2834 7729
rect 2900 7707 2930 7729
rect 2996 7707 3026 7729
rect 3092 7707 3122 7729
rect 3188 7707 3218 7729
rect 3284 7707 3314 7729
rect 3380 7707 3410 7729
rect 2450 7687 3476 7707
rect 2450 7653 2466 7687
rect 2500 7653 2658 7687
rect 2692 7653 2850 7687
rect 2884 7653 3042 7687
rect 3076 7653 3234 7687
rect 3268 7653 3426 7687
rect 3460 7653 3476 7687
rect 2450 7641 3476 7653
rect 3693 7711 3723 7737
rect 4037 7707 4067 7729
rect 4133 7707 4163 7729
rect 4229 7707 4259 7729
rect 4325 7707 4355 7729
rect 4421 7707 4451 7729
rect 4517 7707 4547 7729
rect 4613 7707 4643 7729
rect 4709 7707 4739 7729
rect 4805 7707 4835 7729
rect 4901 7707 4931 7729
rect 3971 7687 4997 7707
rect 3971 7653 3987 7687
rect 4021 7653 4179 7687
rect 4213 7653 4371 7687
rect 4405 7653 4563 7687
rect 4597 7653 4755 7687
rect 4789 7653 4947 7687
rect 4981 7653 4997 7687
rect 3971 7641 4997 7653
rect 5400 7724 5430 7750
rect 297 7204 1323 7220
rect 297 7170 313 7204
rect 347 7170 505 7204
rect 539 7170 697 7204
rect 731 7170 889 7204
rect 923 7170 1081 7204
rect 1115 7170 1273 7204
rect 1307 7170 1323 7204
rect 297 7154 1323 7170
rect 363 7122 393 7154
rect 459 7122 489 7154
rect 555 7122 585 7154
rect 651 7122 681 7154
rect 747 7122 777 7154
rect 843 7122 873 7154
rect 939 7122 969 7154
rect 1035 7122 1065 7154
rect 1131 7122 1161 7154
rect 1227 7122 1257 7154
rect 363 6824 393 6850
rect 459 6824 489 6850
rect 555 6824 585 6850
rect 651 6824 681 6850
rect 747 6824 777 6850
rect 843 6824 873 6850
rect 939 6824 969 6850
rect 1035 6824 1065 6850
rect 1131 6824 1161 6850
rect 1227 6824 1257 6850
rect 2450 7208 3476 7224
rect 2450 7174 2466 7208
rect 2500 7174 2658 7208
rect 2692 7174 2850 7208
rect 2884 7174 3042 7208
rect 3076 7174 3234 7208
rect 3268 7174 3426 7208
rect 3460 7174 3476 7208
rect 2450 7158 3476 7174
rect 2516 7126 2546 7158
rect 2612 7126 2642 7158
rect 2708 7126 2738 7158
rect 2804 7126 2834 7158
rect 2900 7126 2930 7158
rect 2996 7126 3026 7158
rect 3092 7126 3122 7158
rect 3188 7126 3218 7158
rect 3284 7126 3314 7158
rect 3380 7126 3410 7158
rect 2516 6828 2546 6854
rect 2612 6828 2642 6854
rect 2708 6828 2738 6854
rect 2804 6828 2834 6854
rect 2900 6828 2930 6854
rect 2996 6828 3026 6854
rect 3092 6828 3122 6854
rect 3188 6828 3218 6854
rect 3284 6828 3314 6854
rect 3380 6828 3410 6854
rect 3971 7208 4997 7224
rect 3971 7174 3987 7208
rect 4021 7174 4179 7208
rect 4213 7174 4371 7208
rect 4405 7174 4563 7208
rect 4597 7174 4755 7208
rect 4789 7174 4947 7208
rect 4981 7174 4997 7208
rect 3971 7158 4997 7174
rect 4037 7126 4067 7158
rect 4133 7126 4163 7158
rect 4229 7126 4259 7158
rect 4325 7126 4355 7158
rect 4421 7126 4451 7158
rect 4517 7126 4547 7158
rect 4613 7126 4643 7158
rect 4709 7126 4739 7158
rect 4805 7126 4835 7158
rect 4901 7126 4931 7158
rect 5400 6913 5430 6939
rect 4037 6828 4067 6854
rect 4133 6828 4163 6854
rect 4229 6828 4259 6854
rect 4325 6828 4355 6854
rect 4421 6828 4451 6854
rect 4517 6828 4547 6854
rect 4613 6828 4643 6854
rect 4709 6828 4739 6854
rect 4805 6828 4835 6854
rect 4901 6828 4931 6854
rect 5400 6681 5430 6713
rect 5400 6665 5486 6681
rect 363 6542 393 6568
rect 459 6542 489 6568
rect 555 6542 585 6568
rect 651 6542 681 6568
rect 747 6542 777 6568
rect 843 6542 873 6568
rect 939 6542 969 6568
rect 1035 6542 1065 6568
rect 1131 6542 1161 6568
rect 1227 6542 1257 6568
rect 363 6416 393 6438
rect 459 6416 489 6438
rect 555 6416 585 6438
rect 651 6416 681 6438
rect 747 6416 777 6438
rect 843 6416 873 6438
rect 939 6416 969 6438
rect 1035 6416 1065 6438
rect 1131 6416 1161 6438
rect 1227 6416 1257 6438
rect 297 6396 1323 6416
rect 297 6362 313 6396
rect 347 6362 505 6396
rect 539 6362 697 6396
rect 731 6362 889 6396
rect 923 6362 1081 6396
rect 1115 6362 1273 6396
rect 1307 6362 1323 6396
rect 297 6350 1323 6362
rect 2516 6546 2546 6572
rect 2612 6546 2642 6572
rect 2708 6546 2738 6572
rect 2804 6546 2834 6572
rect 2900 6546 2930 6572
rect 2996 6546 3026 6572
rect 3092 6546 3122 6572
rect 3188 6546 3218 6572
rect 3284 6546 3314 6572
rect 3380 6546 3410 6572
rect 3675 6622 3741 6638
rect 3675 6588 3691 6622
rect 3725 6588 3741 6622
rect 3675 6572 3741 6588
rect 3693 6550 3723 6572
rect 4037 6546 4067 6572
rect 4133 6546 4163 6572
rect 4229 6546 4259 6572
rect 4325 6546 4355 6572
rect 4421 6546 4451 6572
rect 4517 6546 4547 6572
rect 4613 6546 4643 6572
rect 4709 6546 4739 6572
rect 4805 6546 4835 6572
rect 4901 6546 4931 6572
rect 5400 6631 5436 6665
rect 5470 6631 5486 6665
rect 5400 6615 5486 6631
rect 5400 6593 5430 6615
rect 2516 6420 2546 6442
rect 2612 6420 2642 6442
rect 2708 6420 2738 6442
rect 2804 6420 2834 6442
rect 2900 6420 2930 6442
rect 2996 6420 3026 6442
rect 3092 6420 3122 6442
rect 3188 6420 3218 6442
rect 3284 6420 3314 6442
rect 3380 6420 3410 6442
rect 2450 6400 3476 6420
rect 2450 6366 2466 6400
rect 2500 6366 2658 6400
rect 2692 6366 2850 6400
rect 2884 6366 3042 6400
rect 3076 6366 3234 6400
rect 3268 6366 3426 6400
rect 3460 6366 3476 6400
rect 2450 6354 3476 6366
rect 3693 6424 3723 6450
rect 4037 6420 4067 6442
rect 4133 6420 4163 6442
rect 4229 6420 4259 6442
rect 4325 6420 4355 6442
rect 4421 6420 4451 6442
rect 4517 6420 4547 6442
rect 4613 6420 4643 6442
rect 4709 6420 4739 6442
rect 4805 6420 4835 6442
rect 4901 6420 4931 6442
rect 3971 6400 4997 6420
rect 3971 6366 3987 6400
rect 4021 6366 4179 6400
rect 4213 6366 4371 6400
rect 4405 6366 4563 6400
rect 4597 6366 4755 6400
rect 4789 6366 4947 6400
rect 4981 6366 4997 6400
rect 3971 6354 4997 6366
rect 5400 6437 5430 6463
rect 297 5917 1323 5933
rect 297 5883 313 5917
rect 347 5883 505 5917
rect 539 5883 697 5917
rect 731 5883 889 5917
rect 923 5883 1081 5917
rect 1115 5883 1273 5917
rect 1307 5883 1323 5917
rect 297 5867 1323 5883
rect 363 5835 393 5867
rect 459 5835 489 5867
rect 555 5835 585 5867
rect 651 5835 681 5867
rect 747 5835 777 5867
rect 843 5835 873 5867
rect 939 5835 969 5867
rect 1035 5835 1065 5867
rect 1131 5835 1161 5867
rect 1227 5835 1257 5867
rect 363 5537 393 5563
rect 459 5537 489 5563
rect 555 5537 585 5563
rect 651 5537 681 5563
rect 747 5537 777 5563
rect 843 5537 873 5563
rect 939 5537 969 5563
rect 1035 5537 1065 5563
rect 1131 5537 1161 5563
rect 1227 5537 1257 5563
rect 2450 5921 3476 5937
rect 2450 5887 2466 5921
rect 2500 5887 2658 5921
rect 2692 5887 2850 5921
rect 2884 5887 3042 5921
rect 3076 5887 3234 5921
rect 3268 5887 3426 5921
rect 3460 5887 3476 5921
rect 2450 5871 3476 5887
rect 2516 5839 2546 5871
rect 2612 5839 2642 5871
rect 2708 5839 2738 5871
rect 2804 5839 2834 5871
rect 2900 5839 2930 5871
rect 2996 5839 3026 5871
rect 3092 5839 3122 5871
rect 3188 5839 3218 5871
rect 3284 5839 3314 5871
rect 3380 5839 3410 5871
rect 2516 5541 2546 5567
rect 2612 5541 2642 5567
rect 2708 5541 2738 5567
rect 2804 5541 2834 5567
rect 2900 5541 2930 5567
rect 2996 5541 3026 5567
rect 3092 5541 3122 5567
rect 3188 5541 3218 5567
rect 3284 5541 3314 5567
rect 3380 5541 3410 5567
rect 3971 5921 4997 5937
rect 3971 5887 3987 5921
rect 4021 5887 4179 5921
rect 4213 5887 4371 5921
rect 4405 5887 4563 5921
rect 4597 5887 4755 5921
rect 4789 5887 4947 5921
rect 4981 5887 4997 5921
rect 3971 5871 4997 5887
rect 4037 5839 4067 5871
rect 4133 5839 4163 5871
rect 4229 5839 4259 5871
rect 4325 5839 4355 5871
rect 4421 5839 4451 5871
rect 4517 5839 4547 5871
rect 4613 5839 4643 5871
rect 4709 5839 4739 5871
rect 4805 5839 4835 5871
rect 4901 5839 4931 5871
rect 5400 5626 5430 5652
rect 4037 5541 4067 5567
rect 4133 5541 4163 5567
rect 4229 5541 4259 5567
rect 4325 5541 4355 5567
rect 4421 5541 4451 5567
rect 4517 5541 4547 5567
rect 4613 5541 4643 5567
rect 4709 5541 4739 5567
rect 4805 5541 4835 5567
rect 4901 5541 4931 5567
rect 5400 5394 5430 5426
rect 5400 5378 5486 5394
rect 363 5255 393 5281
rect 459 5255 489 5281
rect 555 5255 585 5281
rect 651 5255 681 5281
rect 747 5255 777 5281
rect 843 5255 873 5281
rect 939 5255 969 5281
rect 1035 5255 1065 5281
rect 1131 5255 1161 5281
rect 1227 5255 1257 5281
rect 363 5129 393 5151
rect 459 5129 489 5151
rect 555 5129 585 5151
rect 651 5129 681 5151
rect 747 5129 777 5151
rect 843 5129 873 5151
rect 939 5129 969 5151
rect 1035 5129 1065 5151
rect 1131 5129 1161 5151
rect 1227 5129 1257 5151
rect 297 5109 1323 5129
rect 297 5075 313 5109
rect 347 5075 505 5109
rect 539 5075 697 5109
rect 731 5075 889 5109
rect 923 5075 1081 5109
rect 1115 5075 1273 5109
rect 1307 5075 1323 5109
rect 297 5063 1323 5075
rect 2516 5259 2546 5285
rect 2612 5259 2642 5285
rect 2708 5259 2738 5285
rect 2804 5259 2834 5285
rect 2900 5259 2930 5285
rect 2996 5259 3026 5285
rect 3092 5259 3122 5285
rect 3188 5259 3218 5285
rect 3284 5259 3314 5285
rect 3380 5259 3410 5285
rect 3675 5335 3741 5351
rect 3675 5301 3691 5335
rect 3725 5301 3741 5335
rect 3675 5285 3741 5301
rect 3693 5263 3723 5285
rect 4037 5259 4067 5285
rect 4133 5259 4163 5285
rect 4229 5259 4259 5285
rect 4325 5259 4355 5285
rect 4421 5259 4451 5285
rect 4517 5259 4547 5285
rect 4613 5259 4643 5285
rect 4709 5259 4739 5285
rect 4805 5259 4835 5285
rect 4901 5259 4931 5285
rect 5400 5344 5436 5378
rect 5470 5344 5486 5378
rect 5400 5328 5486 5344
rect 5400 5306 5430 5328
rect 2516 5133 2546 5155
rect 2612 5133 2642 5155
rect 2708 5133 2738 5155
rect 2804 5133 2834 5155
rect 2900 5133 2930 5155
rect 2996 5133 3026 5155
rect 3092 5133 3122 5155
rect 3188 5133 3218 5155
rect 3284 5133 3314 5155
rect 3380 5133 3410 5155
rect 2450 5113 3476 5133
rect 2450 5079 2466 5113
rect 2500 5079 2658 5113
rect 2692 5079 2850 5113
rect 2884 5079 3042 5113
rect 3076 5079 3234 5113
rect 3268 5079 3426 5113
rect 3460 5079 3476 5113
rect 2450 5067 3476 5079
rect 3693 5137 3723 5163
rect 4037 5133 4067 5155
rect 4133 5133 4163 5155
rect 4229 5133 4259 5155
rect 4325 5133 4355 5155
rect 4421 5133 4451 5155
rect 4517 5133 4547 5155
rect 4613 5133 4643 5155
rect 4709 5133 4739 5155
rect 4805 5133 4835 5155
rect 4901 5133 4931 5155
rect 3971 5113 4997 5133
rect 3971 5079 3987 5113
rect 4021 5079 4179 5113
rect 4213 5079 4371 5113
rect 4405 5079 4563 5113
rect 4597 5079 4755 5113
rect 4789 5079 4947 5113
rect 4981 5079 4997 5113
rect 3971 5067 4997 5079
rect 5400 5150 5430 5176
rect 297 4630 1323 4646
rect 297 4596 313 4630
rect 347 4596 505 4630
rect 539 4596 697 4630
rect 731 4596 889 4630
rect 923 4596 1081 4630
rect 1115 4596 1273 4630
rect 1307 4596 1323 4630
rect 297 4580 1323 4596
rect 363 4548 393 4580
rect 459 4548 489 4580
rect 555 4548 585 4580
rect 651 4548 681 4580
rect 747 4548 777 4580
rect 843 4548 873 4580
rect 939 4548 969 4580
rect 1035 4548 1065 4580
rect 1131 4548 1161 4580
rect 1227 4548 1257 4580
rect 363 4250 393 4276
rect 459 4250 489 4276
rect 555 4250 585 4276
rect 651 4250 681 4276
rect 747 4250 777 4276
rect 843 4250 873 4276
rect 939 4250 969 4276
rect 1035 4250 1065 4276
rect 1131 4250 1161 4276
rect 1227 4250 1257 4276
rect 2450 4634 3476 4650
rect 2450 4600 2466 4634
rect 2500 4600 2658 4634
rect 2692 4600 2850 4634
rect 2884 4600 3042 4634
rect 3076 4600 3234 4634
rect 3268 4600 3426 4634
rect 3460 4600 3476 4634
rect 2450 4584 3476 4600
rect 2516 4552 2546 4584
rect 2612 4552 2642 4584
rect 2708 4552 2738 4584
rect 2804 4552 2834 4584
rect 2900 4552 2930 4584
rect 2996 4552 3026 4584
rect 3092 4552 3122 4584
rect 3188 4552 3218 4584
rect 3284 4552 3314 4584
rect 3380 4552 3410 4584
rect 2516 4254 2546 4280
rect 2612 4254 2642 4280
rect 2708 4254 2738 4280
rect 2804 4254 2834 4280
rect 2900 4254 2930 4280
rect 2996 4254 3026 4280
rect 3092 4254 3122 4280
rect 3188 4254 3218 4280
rect 3284 4254 3314 4280
rect 3380 4254 3410 4280
rect 3971 4634 4997 4650
rect 3971 4600 3987 4634
rect 4021 4600 4179 4634
rect 4213 4600 4371 4634
rect 4405 4600 4563 4634
rect 4597 4600 4755 4634
rect 4789 4600 4947 4634
rect 4981 4600 4997 4634
rect 3971 4584 4997 4600
rect 4037 4552 4067 4584
rect 4133 4552 4163 4584
rect 4229 4552 4259 4584
rect 4325 4552 4355 4584
rect 4421 4552 4451 4584
rect 4517 4552 4547 4584
rect 4613 4552 4643 4584
rect 4709 4552 4739 4584
rect 4805 4552 4835 4584
rect 4901 4552 4931 4584
rect 5400 4339 5430 4365
rect 4037 4254 4067 4280
rect 4133 4254 4163 4280
rect 4229 4254 4259 4280
rect 4325 4254 4355 4280
rect 4421 4254 4451 4280
rect 4517 4254 4547 4280
rect 4613 4254 4643 4280
rect 4709 4254 4739 4280
rect 4805 4254 4835 4280
rect 4901 4254 4931 4280
rect 5400 4107 5430 4139
rect 5400 4091 5486 4107
rect 363 3968 393 3994
rect 459 3968 489 3994
rect 555 3968 585 3994
rect 651 3968 681 3994
rect 747 3968 777 3994
rect 843 3968 873 3994
rect 939 3968 969 3994
rect 1035 3968 1065 3994
rect 1131 3968 1161 3994
rect 1227 3968 1257 3994
rect 363 3842 393 3864
rect 459 3842 489 3864
rect 555 3842 585 3864
rect 651 3842 681 3864
rect 747 3842 777 3864
rect 843 3842 873 3864
rect 939 3842 969 3864
rect 1035 3842 1065 3864
rect 1131 3842 1161 3864
rect 1227 3842 1257 3864
rect 297 3822 1323 3842
rect 297 3788 313 3822
rect 347 3788 505 3822
rect 539 3788 697 3822
rect 731 3788 889 3822
rect 923 3788 1081 3822
rect 1115 3788 1273 3822
rect 1307 3788 1323 3822
rect 297 3776 1323 3788
rect 2516 3972 2546 3998
rect 2612 3972 2642 3998
rect 2708 3972 2738 3998
rect 2804 3972 2834 3998
rect 2900 3972 2930 3998
rect 2996 3972 3026 3998
rect 3092 3972 3122 3998
rect 3188 3972 3218 3998
rect 3284 3972 3314 3998
rect 3380 3972 3410 3998
rect 3675 4048 3741 4064
rect 3675 4014 3691 4048
rect 3725 4014 3741 4048
rect 3675 3998 3741 4014
rect 3693 3976 3723 3998
rect 4037 3972 4067 3998
rect 4133 3972 4163 3998
rect 4229 3972 4259 3998
rect 4325 3972 4355 3998
rect 4421 3972 4451 3998
rect 4517 3972 4547 3998
rect 4613 3972 4643 3998
rect 4709 3972 4739 3998
rect 4805 3972 4835 3998
rect 4901 3972 4931 3998
rect 5400 4057 5436 4091
rect 5470 4057 5486 4091
rect 5400 4041 5486 4057
rect 5400 4019 5430 4041
rect 2516 3846 2546 3868
rect 2612 3846 2642 3868
rect 2708 3846 2738 3868
rect 2804 3846 2834 3868
rect 2900 3846 2930 3868
rect 2996 3846 3026 3868
rect 3092 3846 3122 3868
rect 3188 3846 3218 3868
rect 3284 3846 3314 3868
rect 3380 3846 3410 3868
rect 2450 3826 3476 3846
rect 2450 3792 2466 3826
rect 2500 3792 2658 3826
rect 2692 3792 2850 3826
rect 2884 3792 3042 3826
rect 3076 3792 3234 3826
rect 3268 3792 3426 3826
rect 3460 3792 3476 3826
rect 2450 3780 3476 3792
rect 3693 3850 3723 3876
rect 4037 3846 4067 3868
rect 4133 3846 4163 3868
rect 4229 3846 4259 3868
rect 4325 3846 4355 3868
rect 4421 3846 4451 3868
rect 4517 3846 4547 3868
rect 4613 3846 4643 3868
rect 4709 3846 4739 3868
rect 4805 3846 4835 3868
rect 4901 3846 4931 3868
rect 3971 3826 4997 3846
rect 3971 3792 3987 3826
rect 4021 3792 4179 3826
rect 4213 3792 4371 3826
rect 4405 3792 4563 3826
rect 4597 3792 4755 3826
rect 4789 3792 4947 3826
rect 4981 3792 4997 3826
rect 3971 3780 4997 3792
rect 5400 3863 5430 3889
rect 297 3343 1323 3359
rect 297 3309 313 3343
rect 347 3309 505 3343
rect 539 3309 697 3343
rect 731 3309 889 3343
rect 923 3309 1081 3343
rect 1115 3309 1273 3343
rect 1307 3309 1323 3343
rect 297 3293 1323 3309
rect 363 3261 393 3293
rect 459 3261 489 3293
rect 555 3261 585 3293
rect 651 3261 681 3293
rect 747 3261 777 3293
rect 843 3261 873 3293
rect 939 3261 969 3293
rect 1035 3261 1065 3293
rect 1131 3261 1161 3293
rect 1227 3261 1257 3293
rect 363 2963 393 2989
rect 459 2963 489 2989
rect 555 2963 585 2989
rect 651 2963 681 2989
rect 747 2963 777 2989
rect 843 2963 873 2989
rect 939 2963 969 2989
rect 1035 2963 1065 2989
rect 1131 2963 1161 2989
rect 1227 2963 1257 2989
rect 2450 3347 3476 3363
rect 2450 3313 2466 3347
rect 2500 3313 2658 3347
rect 2692 3313 2850 3347
rect 2884 3313 3042 3347
rect 3076 3313 3234 3347
rect 3268 3313 3426 3347
rect 3460 3313 3476 3347
rect 2450 3297 3476 3313
rect 2516 3265 2546 3297
rect 2612 3265 2642 3297
rect 2708 3265 2738 3297
rect 2804 3265 2834 3297
rect 2900 3265 2930 3297
rect 2996 3265 3026 3297
rect 3092 3265 3122 3297
rect 3188 3265 3218 3297
rect 3284 3265 3314 3297
rect 3380 3265 3410 3297
rect 2516 2967 2546 2993
rect 2612 2967 2642 2993
rect 2708 2967 2738 2993
rect 2804 2967 2834 2993
rect 2900 2967 2930 2993
rect 2996 2967 3026 2993
rect 3092 2967 3122 2993
rect 3188 2967 3218 2993
rect 3284 2967 3314 2993
rect 3380 2967 3410 2993
rect 3971 3347 4997 3363
rect 3971 3313 3987 3347
rect 4021 3313 4179 3347
rect 4213 3313 4371 3347
rect 4405 3313 4563 3347
rect 4597 3313 4755 3347
rect 4789 3313 4947 3347
rect 4981 3313 4997 3347
rect 3971 3297 4997 3313
rect 4037 3265 4067 3297
rect 4133 3265 4163 3297
rect 4229 3265 4259 3297
rect 4325 3265 4355 3297
rect 4421 3265 4451 3297
rect 4517 3265 4547 3297
rect 4613 3265 4643 3297
rect 4709 3265 4739 3297
rect 4805 3265 4835 3297
rect 4901 3265 4931 3297
rect 5400 3052 5430 3078
rect 4037 2967 4067 2993
rect 4133 2967 4163 2993
rect 4229 2967 4259 2993
rect 4325 2967 4355 2993
rect 4421 2967 4451 2993
rect 4517 2967 4547 2993
rect 4613 2967 4643 2993
rect 4709 2967 4739 2993
rect 4805 2967 4835 2993
rect 4901 2967 4931 2993
rect 5400 2820 5430 2852
rect 5400 2804 5486 2820
rect 363 2681 393 2707
rect 459 2681 489 2707
rect 555 2681 585 2707
rect 651 2681 681 2707
rect 747 2681 777 2707
rect 843 2681 873 2707
rect 939 2681 969 2707
rect 1035 2681 1065 2707
rect 1131 2681 1161 2707
rect 1227 2681 1257 2707
rect 363 2555 393 2577
rect 459 2555 489 2577
rect 555 2555 585 2577
rect 651 2555 681 2577
rect 747 2555 777 2577
rect 843 2555 873 2577
rect 939 2555 969 2577
rect 1035 2555 1065 2577
rect 1131 2555 1161 2577
rect 1227 2555 1257 2577
rect 297 2535 1323 2555
rect 297 2501 313 2535
rect 347 2501 505 2535
rect 539 2501 697 2535
rect 731 2501 889 2535
rect 923 2501 1081 2535
rect 1115 2501 1273 2535
rect 1307 2501 1323 2535
rect 297 2489 1323 2501
rect 2516 2685 2546 2711
rect 2612 2685 2642 2711
rect 2708 2685 2738 2711
rect 2804 2685 2834 2711
rect 2900 2685 2930 2711
rect 2996 2685 3026 2711
rect 3092 2685 3122 2711
rect 3188 2685 3218 2711
rect 3284 2685 3314 2711
rect 3380 2685 3410 2711
rect 3675 2761 3741 2777
rect 3675 2727 3691 2761
rect 3725 2727 3741 2761
rect 3675 2711 3741 2727
rect 3693 2689 3723 2711
rect 4037 2685 4067 2711
rect 4133 2685 4163 2711
rect 4229 2685 4259 2711
rect 4325 2685 4355 2711
rect 4421 2685 4451 2711
rect 4517 2685 4547 2711
rect 4613 2685 4643 2711
rect 4709 2685 4739 2711
rect 4805 2685 4835 2711
rect 4901 2685 4931 2711
rect 5400 2770 5436 2804
rect 5470 2770 5486 2804
rect 5400 2754 5486 2770
rect 5400 2732 5430 2754
rect 2516 2559 2546 2581
rect 2612 2559 2642 2581
rect 2708 2559 2738 2581
rect 2804 2559 2834 2581
rect 2900 2559 2930 2581
rect 2996 2559 3026 2581
rect 3092 2559 3122 2581
rect 3188 2559 3218 2581
rect 3284 2559 3314 2581
rect 3380 2559 3410 2581
rect 2450 2539 3476 2559
rect 2450 2505 2466 2539
rect 2500 2505 2658 2539
rect 2692 2505 2850 2539
rect 2884 2505 3042 2539
rect 3076 2505 3234 2539
rect 3268 2505 3426 2539
rect 3460 2505 3476 2539
rect 2450 2493 3476 2505
rect 3693 2563 3723 2589
rect 4037 2559 4067 2581
rect 4133 2559 4163 2581
rect 4229 2559 4259 2581
rect 4325 2559 4355 2581
rect 4421 2559 4451 2581
rect 4517 2559 4547 2581
rect 4613 2559 4643 2581
rect 4709 2559 4739 2581
rect 4805 2559 4835 2581
rect 4901 2559 4931 2581
rect 3971 2539 4997 2559
rect 3971 2505 3987 2539
rect 4021 2505 4179 2539
rect 4213 2505 4371 2539
rect 4405 2505 4563 2539
rect 4597 2505 4755 2539
rect 4789 2505 4947 2539
rect 4981 2505 4997 2539
rect 3971 2493 4997 2505
rect 5400 2576 5430 2602
rect 297 2056 1323 2072
rect 297 2022 313 2056
rect 347 2022 505 2056
rect 539 2022 697 2056
rect 731 2022 889 2056
rect 923 2022 1081 2056
rect 1115 2022 1273 2056
rect 1307 2022 1323 2056
rect 297 2006 1323 2022
rect 363 1974 393 2006
rect 459 1974 489 2006
rect 555 1974 585 2006
rect 651 1974 681 2006
rect 747 1974 777 2006
rect 843 1974 873 2006
rect 939 1974 969 2006
rect 1035 1974 1065 2006
rect 1131 1974 1161 2006
rect 1227 1974 1257 2006
rect 363 1676 393 1702
rect 459 1676 489 1702
rect 555 1676 585 1702
rect 651 1676 681 1702
rect 747 1676 777 1702
rect 843 1676 873 1702
rect 939 1676 969 1702
rect 1035 1676 1065 1702
rect 1131 1676 1161 1702
rect 1227 1676 1257 1702
rect 2450 2060 3476 2076
rect 2450 2026 2466 2060
rect 2500 2026 2658 2060
rect 2692 2026 2850 2060
rect 2884 2026 3042 2060
rect 3076 2026 3234 2060
rect 3268 2026 3426 2060
rect 3460 2026 3476 2060
rect 2450 2010 3476 2026
rect 2516 1978 2546 2010
rect 2612 1978 2642 2010
rect 2708 1978 2738 2010
rect 2804 1978 2834 2010
rect 2900 1978 2930 2010
rect 2996 1978 3026 2010
rect 3092 1978 3122 2010
rect 3188 1978 3218 2010
rect 3284 1978 3314 2010
rect 3380 1978 3410 2010
rect 2516 1680 2546 1706
rect 2612 1680 2642 1706
rect 2708 1680 2738 1706
rect 2804 1680 2834 1706
rect 2900 1680 2930 1706
rect 2996 1680 3026 1706
rect 3092 1680 3122 1706
rect 3188 1680 3218 1706
rect 3284 1680 3314 1706
rect 3380 1680 3410 1706
rect 3971 2060 4997 2076
rect 3971 2026 3987 2060
rect 4021 2026 4179 2060
rect 4213 2026 4371 2060
rect 4405 2026 4563 2060
rect 4597 2026 4755 2060
rect 4789 2026 4947 2060
rect 4981 2026 4997 2060
rect 3971 2010 4997 2026
rect 4037 1978 4067 2010
rect 4133 1978 4163 2010
rect 4229 1978 4259 2010
rect 4325 1978 4355 2010
rect 4421 1978 4451 2010
rect 4517 1978 4547 2010
rect 4613 1978 4643 2010
rect 4709 1978 4739 2010
rect 4805 1978 4835 2010
rect 4901 1978 4931 2010
rect 5400 1765 5430 1791
rect 4037 1680 4067 1706
rect 4133 1680 4163 1706
rect 4229 1680 4259 1706
rect 4325 1680 4355 1706
rect 4421 1680 4451 1706
rect 4517 1680 4547 1706
rect 4613 1680 4643 1706
rect 4709 1680 4739 1706
rect 4805 1680 4835 1706
rect 4901 1680 4931 1706
rect 5400 1533 5430 1565
rect 5400 1517 5486 1533
rect 363 1394 393 1420
rect 459 1394 489 1420
rect 555 1394 585 1420
rect 651 1394 681 1420
rect 747 1394 777 1420
rect 843 1394 873 1420
rect 939 1394 969 1420
rect 1035 1394 1065 1420
rect 1131 1394 1161 1420
rect 1227 1394 1257 1420
rect 363 1268 393 1290
rect 459 1268 489 1290
rect 555 1268 585 1290
rect 651 1268 681 1290
rect 747 1268 777 1290
rect 843 1268 873 1290
rect 939 1268 969 1290
rect 1035 1268 1065 1290
rect 1131 1268 1161 1290
rect 1227 1268 1257 1290
rect 297 1248 1323 1268
rect 297 1214 313 1248
rect 347 1214 505 1248
rect 539 1214 697 1248
rect 731 1214 889 1248
rect 923 1214 1081 1248
rect 1115 1214 1273 1248
rect 1307 1214 1323 1248
rect 297 1202 1323 1214
rect 2516 1398 2546 1424
rect 2612 1398 2642 1424
rect 2708 1398 2738 1424
rect 2804 1398 2834 1424
rect 2900 1398 2930 1424
rect 2996 1398 3026 1424
rect 3092 1398 3122 1424
rect 3188 1398 3218 1424
rect 3284 1398 3314 1424
rect 3380 1398 3410 1424
rect 3675 1474 3741 1490
rect 3675 1440 3691 1474
rect 3725 1440 3741 1474
rect 3675 1424 3741 1440
rect 3693 1402 3723 1424
rect 4037 1398 4067 1424
rect 4133 1398 4163 1424
rect 4229 1398 4259 1424
rect 4325 1398 4355 1424
rect 4421 1398 4451 1424
rect 4517 1398 4547 1424
rect 4613 1398 4643 1424
rect 4709 1398 4739 1424
rect 4805 1398 4835 1424
rect 4901 1398 4931 1424
rect 5400 1483 5436 1517
rect 5470 1483 5486 1517
rect 5400 1467 5486 1483
rect 5400 1445 5430 1467
rect 2516 1272 2546 1294
rect 2612 1272 2642 1294
rect 2708 1272 2738 1294
rect 2804 1272 2834 1294
rect 2900 1272 2930 1294
rect 2996 1272 3026 1294
rect 3092 1272 3122 1294
rect 3188 1272 3218 1294
rect 3284 1272 3314 1294
rect 3380 1272 3410 1294
rect 2450 1252 3476 1272
rect 2450 1218 2466 1252
rect 2500 1218 2658 1252
rect 2692 1218 2850 1252
rect 2884 1218 3042 1252
rect 3076 1218 3234 1252
rect 3268 1218 3426 1252
rect 3460 1218 3476 1252
rect 2450 1206 3476 1218
rect 3693 1276 3723 1302
rect 4037 1272 4067 1294
rect 4133 1272 4163 1294
rect 4229 1272 4259 1294
rect 4325 1272 4355 1294
rect 4421 1272 4451 1294
rect 4517 1272 4547 1294
rect 4613 1272 4643 1294
rect 4709 1272 4739 1294
rect 4805 1272 4835 1294
rect 4901 1272 4931 1294
rect 3971 1252 4997 1272
rect 3971 1218 3987 1252
rect 4021 1218 4179 1252
rect 4213 1218 4371 1252
rect 4405 1218 4563 1252
rect 4597 1218 4755 1252
rect 4789 1218 4947 1252
rect 4981 1218 4997 1252
rect 3971 1206 4997 1218
rect 5400 1289 5430 1315
<< polycont >>
rect 313 41919 347 41953
rect 505 41919 539 41953
rect 697 41919 731 41953
rect 889 41919 923 41953
rect 1081 41919 1115 41953
rect 1273 41919 1307 41953
rect 2466 41923 2500 41957
rect 2658 41923 2692 41957
rect 2850 41923 2884 41957
rect 3042 41923 3076 41957
rect 3234 41923 3268 41957
rect 3426 41923 3460 41957
rect 3987 41923 4021 41957
rect 4179 41923 4213 41957
rect 4371 41923 4405 41957
rect 4563 41923 4597 41957
rect 4755 41923 4789 41957
rect 4947 41923 4981 41957
rect 313 41111 347 41145
rect 505 41111 539 41145
rect 697 41111 731 41145
rect 889 41111 923 41145
rect 1081 41111 1115 41145
rect 1273 41111 1307 41145
rect 3691 41337 3725 41371
rect 5436 41380 5470 41414
rect 2466 41115 2500 41149
rect 2658 41115 2692 41149
rect 2850 41115 2884 41149
rect 3042 41115 3076 41149
rect 3234 41115 3268 41149
rect 3426 41115 3460 41149
rect 3987 41115 4021 41149
rect 4179 41115 4213 41149
rect 4371 41115 4405 41149
rect 4563 41115 4597 41149
rect 4755 41115 4789 41149
rect 4947 41115 4981 41149
rect 313 40632 347 40666
rect 505 40632 539 40666
rect 697 40632 731 40666
rect 889 40632 923 40666
rect 1081 40632 1115 40666
rect 1273 40632 1307 40666
rect 2466 40636 2500 40670
rect 2658 40636 2692 40670
rect 2850 40636 2884 40670
rect 3042 40636 3076 40670
rect 3234 40636 3268 40670
rect 3426 40636 3460 40670
rect 3987 40636 4021 40670
rect 4179 40636 4213 40670
rect 4371 40636 4405 40670
rect 4563 40636 4597 40670
rect 4755 40636 4789 40670
rect 4947 40636 4981 40670
rect 313 39824 347 39858
rect 505 39824 539 39858
rect 697 39824 731 39858
rect 889 39824 923 39858
rect 1081 39824 1115 39858
rect 1273 39824 1307 39858
rect 3691 40050 3725 40084
rect 5436 40093 5470 40127
rect 2466 39828 2500 39862
rect 2658 39828 2692 39862
rect 2850 39828 2884 39862
rect 3042 39828 3076 39862
rect 3234 39828 3268 39862
rect 3426 39828 3460 39862
rect 3987 39828 4021 39862
rect 4179 39828 4213 39862
rect 4371 39828 4405 39862
rect 4563 39828 4597 39862
rect 4755 39828 4789 39862
rect 4947 39828 4981 39862
rect 313 39345 347 39379
rect 505 39345 539 39379
rect 697 39345 731 39379
rect 889 39345 923 39379
rect 1081 39345 1115 39379
rect 1273 39345 1307 39379
rect 2466 39349 2500 39383
rect 2658 39349 2692 39383
rect 2850 39349 2884 39383
rect 3042 39349 3076 39383
rect 3234 39349 3268 39383
rect 3426 39349 3460 39383
rect 3987 39349 4021 39383
rect 4179 39349 4213 39383
rect 4371 39349 4405 39383
rect 4563 39349 4597 39383
rect 4755 39349 4789 39383
rect 4947 39349 4981 39383
rect 313 38537 347 38571
rect 505 38537 539 38571
rect 697 38537 731 38571
rect 889 38537 923 38571
rect 1081 38537 1115 38571
rect 1273 38537 1307 38571
rect 3691 38763 3725 38797
rect 5436 38806 5470 38840
rect 2466 38541 2500 38575
rect 2658 38541 2692 38575
rect 2850 38541 2884 38575
rect 3042 38541 3076 38575
rect 3234 38541 3268 38575
rect 3426 38541 3460 38575
rect 3987 38541 4021 38575
rect 4179 38541 4213 38575
rect 4371 38541 4405 38575
rect 4563 38541 4597 38575
rect 4755 38541 4789 38575
rect 4947 38541 4981 38575
rect 313 38058 347 38092
rect 505 38058 539 38092
rect 697 38058 731 38092
rect 889 38058 923 38092
rect 1081 38058 1115 38092
rect 1273 38058 1307 38092
rect 2466 38062 2500 38096
rect 2658 38062 2692 38096
rect 2850 38062 2884 38096
rect 3042 38062 3076 38096
rect 3234 38062 3268 38096
rect 3426 38062 3460 38096
rect 3987 38062 4021 38096
rect 4179 38062 4213 38096
rect 4371 38062 4405 38096
rect 4563 38062 4597 38096
rect 4755 38062 4789 38096
rect 4947 38062 4981 38096
rect 313 37250 347 37284
rect 505 37250 539 37284
rect 697 37250 731 37284
rect 889 37250 923 37284
rect 1081 37250 1115 37284
rect 1273 37250 1307 37284
rect 3691 37476 3725 37510
rect 5436 37519 5470 37553
rect 2466 37254 2500 37288
rect 2658 37254 2692 37288
rect 2850 37254 2884 37288
rect 3042 37254 3076 37288
rect 3234 37254 3268 37288
rect 3426 37254 3460 37288
rect 3987 37254 4021 37288
rect 4179 37254 4213 37288
rect 4371 37254 4405 37288
rect 4563 37254 4597 37288
rect 4755 37254 4789 37288
rect 4947 37254 4981 37288
rect 313 36771 347 36805
rect 505 36771 539 36805
rect 697 36771 731 36805
rect 889 36771 923 36805
rect 1081 36771 1115 36805
rect 1273 36771 1307 36805
rect 2466 36775 2500 36809
rect 2658 36775 2692 36809
rect 2850 36775 2884 36809
rect 3042 36775 3076 36809
rect 3234 36775 3268 36809
rect 3426 36775 3460 36809
rect 3987 36775 4021 36809
rect 4179 36775 4213 36809
rect 4371 36775 4405 36809
rect 4563 36775 4597 36809
rect 4755 36775 4789 36809
rect 4947 36775 4981 36809
rect 313 35963 347 35997
rect 505 35963 539 35997
rect 697 35963 731 35997
rect 889 35963 923 35997
rect 1081 35963 1115 35997
rect 1273 35963 1307 35997
rect 3691 36189 3725 36223
rect 5436 36232 5470 36266
rect 2466 35967 2500 36001
rect 2658 35967 2692 36001
rect 2850 35967 2884 36001
rect 3042 35967 3076 36001
rect 3234 35967 3268 36001
rect 3426 35967 3460 36001
rect 3987 35967 4021 36001
rect 4179 35967 4213 36001
rect 4371 35967 4405 36001
rect 4563 35967 4597 36001
rect 4755 35967 4789 36001
rect 4947 35967 4981 36001
rect 313 35484 347 35518
rect 505 35484 539 35518
rect 697 35484 731 35518
rect 889 35484 923 35518
rect 1081 35484 1115 35518
rect 1273 35484 1307 35518
rect 2466 35488 2500 35522
rect 2658 35488 2692 35522
rect 2850 35488 2884 35522
rect 3042 35488 3076 35522
rect 3234 35488 3268 35522
rect 3426 35488 3460 35522
rect 3987 35488 4021 35522
rect 4179 35488 4213 35522
rect 4371 35488 4405 35522
rect 4563 35488 4597 35522
rect 4755 35488 4789 35522
rect 4947 35488 4981 35522
rect 313 34676 347 34710
rect 505 34676 539 34710
rect 697 34676 731 34710
rect 889 34676 923 34710
rect 1081 34676 1115 34710
rect 1273 34676 1307 34710
rect 3691 34902 3725 34936
rect 5436 34945 5470 34979
rect 2466 34680 2500 34714
rect 2658 34680 2692 34714
rect 2850 34680 2884 34714
rect 3042 34680 3076 34714
rect 3234 34680 3268 34714
rect 3426 34680 3460 34714
rect 3987 34680 4021 34714
rect 4179 34680 4213 34714
rect 4371 34680 4405 34714
rect 4563 34680 4597 34714
rect 4755 34680 4789 34714
rect 4947 34680 4981 34714
rect 313 34197 347 34231
rect 505 34197 539 34231
rect 697 34197 731 34231
rect 889 34197 923 34231
rect 1081 34197 1115 34231
rect 1273 34197 1307 34231
rect 2466 34201 2500 34235
rect 2658 34201 2692 34235
rect 2850 34201 2884 34235
rect 3042 34201 3076 34235
rect 3234 34201 3268 34235
rect 3426 34201 3460 34235
rect 3987 34201 4021 34235
rect 4179 34201 4213 34235
rect 4371 34201 4405 34235
rect 4563 34201 4597 34235
rect 4755 34201 4789 34235
rect 4947 34201 4981 34235
rect 313 33389 347 33423
rect 505 33389 539 33423
rect 697 33389 731 33423
rect 889 33389 923 33423
rect 1081 33389 1115 33423
rect 1273 33389 1307 33423
rect 3691 33615 3725 33649
rect 5436 33658 5470 33692
rect 2466 33393 2500 33427
rect 2658 33393 2692 33427
rect 2850 33393 2884 33427
rect 3042 33393 3076 33427
rect 3234 33393 3268 33427
rect 3426 33393 3460 33427
rect 3987 33393 4021 33427
rect 4179 33393 4213 33427
rect 4371 33393 4405 33427
rect 4563 33393 4597 33427
rect 4755 33393 4789 33427
rect 4947 33393 4981 33427
rect 313 32910 347 32944
rect 505 32910 539 32944
rect 697 32910 731 32944
rect 889 32910 923 32944
rect 1081 32910 1115 32944
rect 1273 32910 1307 32944
rect 2466 32914 2500 32948
rect 2658 32914 2692 32948
rect 2850 32914 2884 32948
rect 3042 32914 3076 32948
rect 3234 32914 3268 32948
rect 3426 32914 3460 32948
rect 3987 32914 4021 32948
rect 4179 32914 4213 32948
rect 4371 32914 4405 32948
rect 4563 32914 4597 32948
rect 4755 32914 4789 32948
rect 4947 32914 4981 32948
rect 313 32102 347 32136
rect 505 32102 539 32136
rect 697 32102 731 32136
rect 889 32102 923 32136
rect 1081 32102 1115 32136
rect 1273 32102 1307 32136
rect 3691 32328 3725 32362
rect 5436 32371 5470 32405
rect 2466 32106 2500 32140
rect 2658 32106 2692 32140
rect 2850 32106 2884 32140
rect 3042 32106 3076 32140
rect 3234 32106 3268 32140
rect 3426 32106 3460 32140
rect 3987 32106 4021 32140
rect 4179 32106 4213 32140
rect 4371 32106 4405 32140
rect 4563 32106 4597 32140
rect 4755 32106 4789 32140
rect 4947 32106 4981 32140
rect 313 31623 347 31657
rect 505 31623 539 31657
rect 697 31623 731 31657
rect 889 31623 923 31657
rect 1081 31623 1115 31657
rect 1273 31623 1307 31657
rect 2466 31627 2500 31661
rect 2658 31627 2692 31661
rect 2850 31627 2884 31661
rect 3042 31627 3076 31661
rect 3234 31627 3268 31661
rect 3426 31627 3460 31661
rect 3987 31627 4021 31661
rect 4179 31627 4213 31661
rect 4371 31627 4405 31661
rect 4563 31627 4597 31661
rect 4755 31627 4789 31661
rect 4947 31627 4981 31661
rect 313 30815 347 30849
rect 505 30815 539 30849
rect 697 30815 731 30849
rect 889 30815 923 30849
rect 1081 30815 1115 30849
rect 1273 30815 1307 30849
rect 3691 31041 3725 31075
rect 5436 31084 5470 31118
rect 2466 30819 2500 30853
rect 2658 30819 2692 30853
rect 2850 30819 2884 30853
rect 3042 30819 3076 30853
rect 3234 30819 3268 30853
rect 3426 30819 3460 30853
rect 3987 30819 4021 30853
rect 4179 30819 4213 30853
rect 4371 30819 4405 30853
rect 4563 30819 4597 30853
rect 4755 30819 4789 30853
rect 4947 30819 4981 30853
rect 313 30336 347 30370
rect 505 30336 539 30370
rect 697 30336 731 30370
rect 889 30336 923 30370
rect 1081 30336 1115 30370
rect 1273 30336 1307 30370
rect 2466 30340 2500 30374
rect 2658 30340 2692 30374
rect 2850 30340 2884 30374
rect 3042 30340 3076 30374
rect 3234 30340 3268 30374
rect 3426 30340 3460 30374
rect 3987 30340 4021 30374
rect 4179 30340 4213 30374
rect 4371 30340 4405 30374
rect 4563 30340 4597 30374
rect 4755 30340 4789 30374
rect 4947 30340 4981 30374
rect 313 29528 347 29562
rect 505 29528 539 29562
rect 697 29528 731 29562
rect 889 29528 923 29562
rect 1081 29528 1115 29562
rect 1273 29528 1307 29562
rect 3691 29754 3725 29788
rect 5436 29797 5470 29831
rect 2466 29532 2500 29566
rect 2658 29532 2692 29566
rect 2850 29532 2884 29566
rect 3042 29532 3076 29566
rect 3234 29532 3268 29566
rect 3426 29532 3460 29566
rect 3987 29532 4021 29566
rect 4179 29532 4213 29566
rect 4371 29532 4405 29566
rect 4563 29532 4597 29566
rect 4755 29532 4789 29566
rect 4947 29532 4981 29566
rect 313 29049 347 29083
rect 505 29049 539 29083
rect 697 29049 731 29083
rect 889 29049 923 29083
rect 1081 29049 1115 29083
rect 1273 29049 1307 29083
rect 2466 29053 2500 29087
rect 2658 29053 2692 29087
rect 2850 29053 2884 29087
rect 3042 29053 3076 29087
rect 3234 29053 3268 29087
rect 3426 29053 3460 29087
rect 3987 29053 4021 29087
rect 4179 29053 4213 29087
rect 4371 29053 4405 29087
rect 4563 29053 4597 29087
rect 4755 29053 4789 29087
rect 4947 29053 4981 29087
rect 313 28241 347 28275
rect 505 28241 539 28275
rect 697 28241 731 28275
rect 889 28241 923 28275
rect 1081 28241 1115 28275
rect 1273 28241 1307 28275
rect 3691 28467 3725 28501
rect 5436 28510 5470 28544
rect 2466 28245 2500 28279
rect 2658 28245 2692 28279
rect 2850 28245 2884 28279
rect 3042 28245 3076 28279
rect 3234 28245 3268 28279
rect 3426 28245 3460 28279
rect 3987 28245 4021 28279
rect 4179 28245 4213 28279
rect 4371 28245 4405 28279
rect 4563 28245 4597 28279
rect 4755 28245 4789 28279
rect 4947 28245 4981 28279
rect 313 27762 347 27796
rect 505 27762 539 27796
rect 697 27762 731 27796
rect 889 27762 923 27796
rect 1081 27762 1115 27796
rect 1273 27762 1307 27796
rect 2466 27766 2500 27800
rect 2658 27766 2692 27800
rect 2850 27766 2884 27800
rect 3042 27766 3076 27800
rect 3234 27766 3268 27800
rect 3426 27766 3460 27800
rect 3987 27766 4021 27800
rect 4179 27766 4213 27800
rect 4371 27766 4405 27800
rect 4563 27766 4597 27800
rect 4755 27766 4789 27800
rect 4947 27766 4981 27800
rect 313 26954 347 26988
rect 505 26954 539 26988
rect 697 26954 731 26988
rect 889 26954 923 26988
rect 1081 26954 1115 26988
rect 1273 26954 1307 26988
rect 3691 27180 3725 27214
rect 5436 27223 5470 27257
rect 2466 26958 2500 26992
rect 2658 26958 2692 26992
rect 2850 26958 2884 26992
rect 3042 26958 3076 26992
rect 3234 26958 3268 26992
rect 3426 26958 3460 26992
rect 3987 26958 4021 26992
rect 4179 26958 4213 26992
rect 4371 26958 4405 26992
rect 4563 26958 4597 26992
rect 4755 26958 4789 26992
rect 4947 26958 4981 26992
rect 313 26475 347 26509
rect 505 26475 539 26509
rect 697 26475 731 26509
rect 889 26475 923 26509
rect 1081 26475 1115 26509
rect 1273 26475 1307 26509
rect 2466 26479 2500 26513
rect 2658 26479 2692 26513
rect 2850 26479 2884 26513
rect 3042 26479 3076 26513
rect 3234 26479 3268 26513
rect 3426 26479 3460 26513
rect 3987 26479 4021 26513
rect 4179 26479 4213 26513
rect 4371 26479 4405 26513
rect 4563 26479 4597 26513
rect 4755 26479 4789 26513
rect 4947 26479 4981 26513
rect 313 25667 347 25701
rect 505 25667 539 25701
rect 697 25667 731 25701
rect 889 25667 923 25701
rect 1081 25667 1115 25701
rect 1273 25667 1307 25701
rect 3691 25893 3725 25927
rect 5436 25936 5470 25970
rect 2466 25671 2500 25705
rect 2658 25671 2692 25705
rect 2850 25671 2884 25705
rect 3042 25671 3076 25705
rect 3234 25671 3268 25705
rect 3426 25671 3460 25705
rect 3987 25671 4021 25705
rect 4179 25671 4213 25705
rect 4371 25671 4405 25705
rect 4563 25671 4597 25705
rect 4755 25671 4789 25705
rect 4947 25671 4981 25705
rect 313 25188 347 25222
rect 505 25188 539 25222
rect 697 25188 731 25222
rect 889 25188 923 25222
rect 1081 25188 1115 25222
rect 1273 25188 1307 25222
rect 2466 25192 2500 25226
rect 2658 25192 2692 25226
rect 2850 25192 2884 25226
rect 3042 25192 3076 25226
rect 3234 25192 3268 25226
rect 3426 25192 3460 25226
rect 3987 25192 4021 25226
rect 4179 25192 4213 25226
rect 4371 25192 4405 25226
rect 4563 25192 4597 25226
rect 4755 25192 4789 25226
rect 4947 25192 4981 25226
rect 313 24380 347 24414
rect 505 24380 539 24414
rect 697 24380 731 24414
rect 889 24380 923 24414
rect 1081 24380 1115 24414
rect 1273 24380 1307 24414
rect 3691 24606 3725 24640
rect 5436 24649 5470 24683
rect 2466 24384 2500 24418
rect 2658 24384 2692 24418
rect 2850 24384 2884 24418
rect 3042 24384 3076 24418
rect 3234 24384 3268 24418
rect 3426 24384 3460 24418
rect 3987 24384 4021 24418
rect 4179 24384 4213 24418
rect 4371 24384 4405 24418
rect 4563 24384 4597 24418
rect 4755 24384 4789 24418
rect 4947 24384 4981 24418
rect 313 23901 347 23935
rect 505 23901 539 23935
rect 697 23901 731 23935
rect 889 23901 923 23935
rect 1081 23901 1115 23935
rect 1273 23901 1307 23935
rect 2466 23905 2500 23939
rect 2658 23905 2692 23939
rect 2850 23905 2884 23939
rect 3042 23905 3076 23939
rect 3234 23905 3268 23939
rect 3426 23905 3460 23939
rect 3987 23905 4021 23939
rect 4179 23905 4213 23939
rect 4371 23905 4405 23939
rect 4563 23905 4597 23939
rect 4755 23905 4789 23939
rect 4947 23905 4981 23939
rect 313 23093 347 23127
rect 505 23093 539 23127
rect 697 23093 731 23127
rect 889 23093 923 23127
rect 1081 23093 1115 23127
rect 1273 23093 1307 23127
rect 3691 23319 3725 23353
rect 5436 23362 5470 23396
rect 2466 23097 2500 23131
rect 2658 23097 2692 23131
rect 2850 23097 2884 23131
rect 3042 23097 3076 23131
rect 3234 23097 3268 23131
rect 3426 23097 3460 23131
rect 3987 23097 4021 23131
rect 4179 23097 4213 23131
rect 4371 23097 4405 23131
rect 4563 23097 4597 23131
rect 4755 23097 4789 23131
rect 4947 23097 4981 23131
rect 313 22614 347 22648
rect 505 22614 539 22648
rect 697 22614 731 22648
rect 889 22614 923 22648
rect 1081 22614 1115 22648
rect 1273 22614 1307 22648
rect 2466 22618 2500 22652
rect 2658 22618 2692 22652
rect 2850 22618 2884 22652
rect 3042 22618 3076 22652
rect 3234 22618 3268 22652
rect 3426 22618 3460 22652
rect 3987 22618 4021 22652
rect 4179 22618 4213 22652
rect 4371 22618 4405 22652
rect 4563 22618 4597 22652
rect 4755 22618 4789 22652
rect 4947 22618 4981 22652
rect 313 21806 347 21840
rect 505 21806 539 21840
rect 697 21806 731 21840
rect 889 21806 923 21840
rect 1081 21806 1115 21840
rect 1273 21806 1307 21840
rect 3691 22032 3725 22066
rect 5436 22075 5470 22109
rect 2466 21810 2500 21844
rect 2658 21810 2692 21844
rect 2850 21810 2884 21844
rect 3042 21810 3076 21844
rect 3234 21810 3268 21844
rect 3426 21810 3460 21844
rect 3987 21810 4021 21844
rect 4179 21810 4213 21844
rect 4371 21810 4405 21844
rect 4563 21810 4597 21844
rect 4755 21810 4789 21844
rect 4947 21810 4981 21844
rect 313 21327 347 21361
rect 505 21327 539 21361
rect 697 21327 731 21361
rect 889 21327 923 21361
rect 1081 21327 1115 21361
rect 1273 21327 1307 21361
rect 2466 21331 2500 21365
rect 2658 21331 2692 21365
rect 2850 21331 2884 21365
rect 3042 21331 3076 21365
rect 3234 21331 3268 21365
rect 3426 21331 3460 21365
rect 3987 21331 4021 21365
rect 4179 21331 4213 21365
rect 4371 21331 4405 21365
rect 4563 21331 4597 21365
rect 4755 21331 4789 21365
rect 4947 21331 4981 21365
rect 313 20519 347 20553
rect 505 20519 539 20553
rect 697 20519 731 20553
rect 889 20519 923 20553
rect 1081 20519 1115 20553
rect 1273 20519 1307 20553
rect 3691 20745 3725 20779
rect 5436 20788 5470 20822
rect 2466 20523 2500 20557
rect 2658 20523 2692 20557
rect 2850 20523 2884 20557
rect 3042 20523 3076 20557
rect 3234 20523 3268 20557
rect 3426 20523 3460 20557
rect 3987 20523 4021 20557
rect 4179 20523 4213 20557
rect 4371 20523 4405 20557
rect 4563 20523 4597 20557
rect 4755 20523 4789 20557
rect 4947 20523 4981 20557
rect 313 20040 347 20074
rect 505 20040 539 20074
rect 697 20040 731 20074
rect 889 20040 923 20074
rect 1081 20040 1115 20074
rect 1273 20040 1307 20074
rect 2466 20044 2500 20078
rect 2658 20044 2692 20078
rect 2850 20044 2884 20078
rect 3042 20044 3076 20078
rect 3234 20044 3268 20078
rect 3426 20044 3460 20078
rect 3987 20044 4021 20078
rect 4179 20044 4213 20078
rect 4371 20044 4405 20078
rect 4563 20044 4597 20078
rect 4755 20044 4789 20078
rect 4947 20044 4981 20078
rect 313 19232 347 19266
rect 505 19232 539 19266
rect 697 19232 731 19266
rect 889 19232 923 19266
rect 1081 19232 1115 19266
rect 1273 19232 1307 19266
rect 3691 19458 3725 19492
rect 5436 19501 5470 19535
rect 2466 19236 2500 19270
rect 2658 19236 2692 19270
rect 2850 19236 2884 19270
rect 3042 19236 3076 19270
rect 3234 19236 3268 19270
rect 3426 19236 3460 19270
rect 3987 19236 4021 19270
rect 4179 19236 4213 19270
rect 4371 19236 4405 19270
rect 4563 19236 4597 19270
rect 4755 19236 4789 19270
rect 4947 19236 4981 19270
rect 313 18753 347 18787
rect 505 18753 539 18787
rect 697 18753 731 18787
rect 889 18753 923 18787
rect 1081 18753 1115 18787
rect 1273 18753 1307 18787
rect 2466 18757 2500 18791
rect 2658 18757 2692 18791
rect 2850 18757 2884 18791
rect 3042 18757 3076 18791
rect 3234 18757 3268 18791
rect 3426 18757 3460 18791
rect 3987 18757 4021 18791
rect 4179 18757 4213 18791
rect 4371 18757 4405 18791
rect 4563 18757 4597 18791
rect 4755 18757 4789 18791
rect 4947 18757 4981 18791
rect 313 17945 347 17979
rect 505 17945 539 17979
rect 697 17945 731 17979
rect 889 17945 923 17979
rect 1081 17945 1115 17979
rect 1273 17945 1307 17979
rect 3691 18171 3725 18205
rect 5436 18214 5470 18248
rect 2466 17949 2500 17983
rect 2658 17949 2692 17983
rect 2850 17949 2884 17983
rect 3042 17949 3076 17983
rect 3234 17949 3268 17983
rect 3426 17949 3460 17983
rect 3987 17949 4021 17983
rect 4179 17949 4213 17983
rect 4371 17949 4405 17983
rect 4563 17949 4597 17983
rect 4755 17949 4789 17983
rect 4947 17949 4981 17983
rect 313 17466 347 17500
rect 505 17466 539 17500
rect 697 17466 731 17500
rect 889 17466 923 17500
rect 1081 17466 1115 17500
rect 1273 17466 1307 17500
rect 2466 17470 2500 17504
rect 2658 17470 2692 17504
rect 2850 17470 2884 17504
rect 3042 17470 3076 17504
rect 3234 17470 3268 17504
rect 3426 17470 3460 17504
rect 3987 17470 4021 17504
rect 4179 17470 4213 17504
rect 4371 17470 4405 17504
rect 4563 17470 4597 17504
rect 4755 17470 4789 17504
rect 4947 17470 4981 17504
rect 313 16658 347 16692
rect 505 16658 539 16692
rect 697 16658 731 16692
rect 889 16658 923 16692
rect 1081 16658 1115 16692
rect 1273 16658 1307 16692
rect 3691 16884 3725 16918
rect 5436 16927 5470 16961
rect 2466 16662 2500 16696
rect 2658 16662 2692 16696
rect 2850 16662 2884 16696
rect 3042 16662 3076 16696
rect 3234 16662 3268 16696
rect 3426 16662 3460 16696
rect 3987 16662 4021 16696
rect 4179 16662 4213 16696
rect 4371 16662 4405 16696
rect 4563 16662 4597 16696
rect 4755 16662 4789 16696
rect 4947 16662 4981 16696
rect 313 16179 347 16213
rect 505 16179 539 16213
rect 697 16179 731 16213
rect 889 16179 923 16213
rect 1081 16179 1115 16213
rect 1273 16179 1307 16213
rect 2466 16183 2500 16217
rect 2658 16183 2692 16217
rect 2850 16183 2884 16217
rect 3042 16183 3076 16217
rect 3234 16183 3268 16217
rect 3426 16183 3460 16217
rect 3987 16183 4021 16217
rect 4179 16183 4213 16217
rect 4371 16183 4405 16217
rect 4563 16183 4597 16217
rect 4755 16183 4789 16217
rect 4947 16183 4981 16217
rect 313 15371 347 15405
rect 505 15371 539 15405
rect 697 15371 731 15405
rect 889 15371 923 15405
rect 1081 15371 1115 15405
rect 1273 15371 1307 15405
rect 3691 15597 3725 15631
rect 5436 15640 5470 15674
rect 2466 15375 2500 15409
rect 2658 15375 2692 15409
rect 2850 15375 2884 15409
rect 3042 15375 3076 15409
rect 3234 15375 3268 15409
rect 3426 15375 3460 15409
rect 3987 15375 4021 15409
rect 4179 15375 4213 15409
rect 4371 15375 4405 15409
rect 4563 15375 4597 15409
rect 4755 15375 4789 15409
rect 4947 15375 4981 15409
rect 313 14892 347 14926
rect 505 14892 539 14926
rect 697 14892 731 14926
rect 889 14892 923 14926
rect 1081 14892 1115 14926
rect 1273 14892 1307 14926
rect 2466 14896 2500 14930
rect 2658 14896 2692 14930
rect 2850 14896 2884 14930
rect 3042 14896 3076 14930
rect 3234 14896 3268 14930
rect 3426 14896 3460 14930
rect 3987 14896 4021 14930
rect 4179 14896 4213 14930
rect 4371 14896 4405 14930
rect 4563 14896 4597 14930
rect 4755 14896 4789 14930
rect 4947 14896 4981 14930
rect 313 14084 347 14118
rect 505 14084 539 14118
rect 697 14084 731 14118
rect 889 14084 923 14118
rect 1081 14084 1115 14118
rect 1273 14084 1307 14118
rect 3691 14310 3725 14344
rect 5436 14353 5470 14387
rect 2466 14088 2500 14122
rect 2658 14088 2692 14122
rect 2850 14088 2884 14122
rect 3042 14088 3076 14122
rect 3234 14088 3268 14122
rect 3426 14088 3460 14122
rect 3987 14088 4021 14122
rect 4179 14088 4213 14122
rect 4371 14088 4405 14122
rect 4563 14088 4597 14122
rect 4755 14088 4789 14122
rect 4947 14088 4981 14122
rect 313 13605 347 13639
rect 505 13605 539 13639
rect 697 13605 731 13639
rect 889 13605 923 13639
rect 1081 13605 1115 13639
rect 1273 13605 1307 13639
rect 2466 13609 2500 13643
rect 2658 13609 2692 13643
rect 2850 13609 2884 13643
rect 3042 13609 3076 13643
rect 3234 13609 3268 13643
rect 3426 13609 3460 13643
rect 3987 13609 4021 13643
rect 4179 13609 4213 13643
rect 4371 13609 4405 13643
rect 4563 13609 4597 13643
rect 4755 13609 4789 13643
rect 4947 13609 4981 13643
rect 313 12797 347 12831
rect 505 12797 539 12831
rect 697 12797 731 12831
rect 889 12797 923 12831
rect 1081 12797 1115 12831
rect 1273 12797 1307 12831
rect 3691 13023 3725 13057
rect 5436 13066 5470 13100
rect 2466 12801 2500 12835
rect 2658 12801 2692 12835
rect 2850 12801 2884 12835
rect 3042 12801 3076 12835
rect 3234 12801 3268 12835
rect 3426 12801 3460 12835
rect 3987 12801 4021 12835
rect 4179 12801 4213 12835
rect 4371 12801 4405 12835
rect 4563 12801 4597 12835
rect 4755 12801 4789 12835
rect 4947 12801 4981 12835
rect 313 12318 347 12352
rect 505 12318 539 12352
rect 697 12318 731 12352
rect 889 12318 923 12352
rect 1081 12318 1115 12352
rect 1273 12318 1307 12352
rect 2466 12322 2500 12356
rect 2658 12322 2692 12356
rect 2850 12322 2884 12356
rect 3042 12322 3076 12356
rect 3234 12322 3268 12356
rect 3426 12322 3460 12356
rect 3987 12322 4021 12356
rect 4179 12322 4213 12356
rect 4371 12322 4405 12356
rect 4563 12322 4597 12356
rect 4755 12322 4789 12356
rect 4947 12322 4981 12356
rect 313 11510 347 11544
rect 505 11510 539 11544
rect 697 11510 731 11544
rect 889 11510 923 11544
rect 1081 11510 1115 11544
rect 1273 11510 1307 11544
rect 3691 11736 3725 11770
rect 5436 11779 5470 11813
rect 2466 11514 2500 11548
rect 2658 11514 2692 11548
rect 2850 11514 2884 11548
rect 3042 11514 3076 11548
rect 3234 11514 3268 11548
rect 3426 11514 3460 11548
rect 3987 11514 4021 11548
rect 4179 11514 4213 11548
rect 4371 11514 4405 11548
rect 4563 11514 4597 11548
rect 4755 11514 4789 11548
rect 4947 11514 4981 11548
rect 313 11031 347 11065
rect 505 11031 539 11065
rect 697 11031 731 11065
rect 889 11031 923 11065
rect 1081 11031 1115 11065
rect 1273 11031 1307 11065
rect 2466 11035 2500 11069
rect 2658 11035 2692 11069
rect 2850 11035 2884 11069
rect 3042 11035 3076 11069
rect 3234 11035 3268 11069
rect 3426 11035 3460 11069
rect 3987 11035 4021 11069
rect 4179 11035 4213 11069
rect 4371 11035 4405 11069
rect 4563 11035 4597 11069
rect 4755 11035 4789 11069
rect 4947 11035 4981 11069
rect 313 10223 347 10257
rect 505 10223 539 10257
rect 697 10223 731 10257
rect 889 10223 923 10257
rect 1081 10223 1115 10257
rect 1273 10223 1307 10257
rect 3691 10449 3725 10483
rect 5436 10492 5470 10526
rect 2466 10227 2500 10261
rect 2658 10227 2692 10261
rect 2850 10227 2884 10261
rect 3042 10227 3076 10261
rect 3234 10227 3268 10261
rect 3426 10227 3460 10261
rect 3987 10227 4021 10261
rect 4179 10227 4213 10261
rect 4371 10227 4405 10261
rect 4563 10227 4597 10261
rect 4755 10227 4789 10261
rect 4947 10227 4981 10261
rect 313 9744 347 9778
rect 505 9744 539 9778
rect 697 9744 731 9778
rect 889 9744 923 9778
rect 1081 9744 1115 9778
rect 1273 9744 1307 9778
rect 2466 9748 2500 9782
rect 2658 9748 2692 9782
rect 2850 9748 2884 9782
rect 3042 9748 3076 9782
rect 3234 9748 3268 9782
rect 3426 9748 3460 9782
rect 3987 9748 4021 9782
rect 4179 9748 4213 9782
rect 4371 9748 4405 9782
rect 4563 9748 4597 9782
rect 4755 9748 4789 9782
rect 4947 9748 4981 9782
rect 313 8936 347 8970
rect 505 8936 539 8970
rect 697 8936 731 8970
rect 889 8936 923 8970
rect 1081 8936 1115 8970
rect 1273 8936 1307 8970
rect 3691 9162 3725 9196
rect 5436 9205 5470 9239
rect 2466 8940 2500 8974
rect 2658 8940 2692 8974
rect 2850 8940 2884 8974
rect 3042 8940 3076 8974
rect 3234 8940 3268 8974
rect 3426 8940 3460 8974
rect 3987 8940 4021 8974
rect 4179 8940 4213 8974
rect 4371 8940 4405 8974
rect 4563 8940 4597 8974
rect 4755 8940 4789 8974
rect 4947 8940 4981 8974
rect 313 8457 347 8491
rect 505 8457 539 8491
rect 697 8457 731 8491
rect 889 8457 923 8491
rect 1081 8457 1115 8491
rect 1273 8457 1307 8491
rect 2466 8461 2500 8495
rect 2658 8461 2692 8495
rect 2850 8461 2884 8495
rect 3042 8461 3076 8495
rect 3234 8461 3268 8495
rect 3426 8461 3460 8495
rect 3987 8461 4021 8495
rect 4179 8461 4213 8495
rect 4371 8461 4405 8495
rect 4563 8461 4597 8495
rect 4755 8461 4789 8495
rect 4947 8461 4981 8495
rect 313 7649 347 7683
rect 505 7649 539 7683
rect 697 7649 731 7683
rect 889 7649 923 7683
rect 1081 7649 1115 7683
rect 1273 7649 1307 7683
rect 3691 7875 3725 7909
rect 5436 7918 5470 7952
rect 2466 7653 2500 7687
rect 2658 7653 2692 7687
rect 2850 7653 2884 7687
rect 3042 7653 3076 7687
rect 3234 7653 3268 7687
rect 3426 7653 3460 7687
rect 3987 7653 4021 7687
rect 4179 7653 4213 7687
rect 4371 7653 4405 7687
rect 4563 7653 4597 7687
rect 4755 7653 4789 7687
rect 4947 7653 4981 7687
rect 313 7170 347 7204
rect 505 7170 539 7204
rect 697 7170 731 7204
rect 889 7170 923 7204
rect 1081 7170 1115 7204
rect 1273 7170 1307 7204
rect 2466 7174 2500 7208
rect 2658 7174 2692 7208
rect 2850 7174 2884 7208
rect 3042 7174 3076 7208
rect 3234 7174 3268 7208
rect 3426 7174 3460 7208
rect 3987 7174 4021 7208
rect 4179 7174 4213 7208
rect 4371 7174 4405 7208
rect 4563 7174 4597 7208
rect 4755 7174 4789 7208
rect 4947 7174 4981 7208
rect 313 6362 347 6396
rect 505 6362 539 6396
rect 697 6362 731 6396
rect 889 6362 923 6396
rect 1081 6362 1115 6396
rect 1273 6362 1307 6396
rect 3691 6588 3725 6622
rect 5436 6631 5470 6665
rect 2466 6366 2500 6400
rect 2658 6366 2692 6400
rect 2850 6366 2884 6400
rect 3042 6366 3076 6400
rect 3234 6366 3268 6400
rect 3426 6366 3460 6400
rect 3987 6366 4021 6400
rect 4179 6366 4213 6400
rect 4371 6366 4405 6400
rect 4563 6366 4597 6400
rect 4755 6366 4789 6400
rect 4947 6366 4981 6400
rect 313 5883 347 5917
rect 505 5883 539 5917
rect 697 5883 731 5917
rect 889 5883 923 5917
rect 1081 5883 1115 5917
rect 1273 5883 1307 5917
rect 2466 5887 2500 5921
rect 2658 5887 2692 5921
rect 2850 5887 2884 5921
rect 3042 5887 3076 5921
rect 3234 5887 3268 5921
rect 3426 5887 3460 5921
rect 3987 5887 4021 5921
rect 4179 5887 4213 5921
rect 4371 5887 4405 5921
rect 4563 5887 4597 5921
rect 4755 5887 4789 5921
rect 4947 5887 4981 5921
rect 313 5075 347 5109
rect 505 5075 539 5109
rect 697 5075 731 5109
rect 889 5075 923 5109
rect 1081 5075 1115 5109
rect 1273 5075 1307 5109
rect 3691 5301 3725 5335
rect 5436 5344 5470 5378
rect 2466 5079 2500 5113
rect 2658 5079 2692 5113
rect 2850 5079 2884 5113
rect 3042 5079 3076 5113
rect 3234 5079 3268 5113
rect 3426 5079 3460 5113
rect 3987 5079 4021 5113
rect 4179 5079 4213 5113
rect 4371 5079 4405 5113
rect 4563 5079 4597 5113
rect 4755 5079 4789 5113
rect 4947 5079 4981 5113
rect 313 4596 347 4630
rect 505 4596 539 4630
rect 697 4596 731 4630
rect 889 4596 923 4630
rect 1081 4596 1115 4630
rect 1273 4596 1307 4630
rect 2466 4600 2500 4634
rect 2658 4600 2692 4634
rect 2850 4600 2884 4634
rect 3042 4600 3076 4634
rect 3234 4600 3268 4634
rect 3426 4600 3460 4634
rect 3987 4600 4021 4634
rect 4179 4600 4213 4634
rect 4371 4600 4405 4634
rect 4563 4600 4597 4634
rect 4755 4600 4789 4634
rect 4947 4600 4981 4634
rect 313 3788 347 3822
rect 505 3788 539 3822
rect 697 3788 731 3822
rect 889 3788 923 3822
rect 1081 3788 1115 3822
rect 1273 3788 1307 3822
rect 3691 4014 3725 4048
rect 5436 4057 5470 4091
rect 2466 3792 2500 3826
rect 2658 3792 2692 3826
rect 2850 3792 2884 3826
rect 3042 3792 3076 3826
rect 3234 3792 3268 3826
rect 3426 3792 3460 3826
rect 3987 3792 4021 3826
rect 4179 3792 4213 3826
rect 4371 3792 4405 3826
rect 4563 3792 4597 3826
rect 4755 3792 4789 3826
rect 4947 3792 4981 3826
rect 313 3309 347 3343
rect 505 3309 539 3343
rect 697 3309 731 3343
rect 889 3309 923 3343
rect 1081 3309 1115 3343
rect 1273 3309 1307 3343
rect 2466 3313 2500 3347
rect 2658 3313 2692 3347
rect 2850 3313 2884 3347
rect 3042 3313 3076 3347
rect 3234 3313 3268 3347
rect 3426 3313 3460 3347
rect 3987 3313 4021 3347
rect 4179 3313 4213 3347
rect 4371 3313 4405 3347
rect 4563 3313 4597 3347
rect 4755 3313 4789 3347
rect 4947 3313 4981 3347
rect 313 2501 347 2535
rect 505 2501 539 2535
rect 697 2501 731 2535
rect 889 2501 923 2535
rect 1081 2501 1115 2535
rect 1273 2501 1307 2535
rect 3691 2727 3725 2761
rect 5436 2770 5470 2804
rect 2466 2505 2500 2539
rect 2658 2505 2692 2539
rect 2850 2505 2884 2539
rect 3042 2505 3076 2539
rect 3234 2505 3268 2539
rect 3426 2505 3460 2539
rect 3987 2505 4021 2539
rect 4179 2505 4213 2539
rect 4371 2505 4405 2539
rect 4563 2505 4597 2539
rect 4755 2505 4789 2539
rect 4947 2505 4981 2539
rect 313 2022 347 2056
rect 505 2022 539 2056
rect 697 2022 731 2056
rect 889 2022 923 2056
rect 1081 2022 1115 2056
rect 1273 2022 1307 2056
rect 2466 2026 2500 2060
rect 2658 2026 2692 2060
rect 2850 2026 2884 2060
rect 3042 2026 3076 2060
rect 3234 2026 3268 2060
rect 3426 2026 3460 2060
rect 3987 2026 4021 2060
rect 4179 2026 4213 2060
rect 4371 2026 4405 2060
rect 4563 2026 4597 2060
rect 4755 2026 4789 2060
rect 4947 2026 4981 2060
rect 313 1214 347 1248
rect 505 1214 539 1248
rect 697 1214 731 1248
rect 889 1214 923 1248
rect 1081 1214 1115 1248
rect 1273 1214 1307 1248
rect 3691 1440 3725 1474
rect 5436 1483 5470 1517
rect 2466 1218 2500 1252
rect 2658 1218 2692 1252
rect 2850 1218 2884 1252
rect 3042 1218 3076 1252
rect 3234 1218 3268 1252
rect 3426 1218 3460 1252
rect 3987 1218 4021 1252
rect 4179 1218 4213 1252
rect 4371 1218 4405 1252
rect 4563 1218 4597 1252
rect 4755 1218 4789 1252
rect 4947 1218 4981 1252
<< locali >>
rect 199 42021 317 42055
rect 351 42021 385 42055
rect 419 42021 453 42055
rect 487 42021 521 42055
rect 555 42021 589 42055
rect 623 42021 657 42055
rect 691 42021 725 42055
rect 759 42021 793 42055
rect 827 42021 861 42055
rect 895 42021 929 42055
rect 963 42021 997 42055
rect 1031 42021 1065 42055
rect 1099 42021 1133 42055
rect 1167 42021 1201 42055
rect 1235 42021 1269 42055
rect 1303 42021 1421 42055
rect 199 41953 233 42021
rect 1387 41953 1421 42021
rect 297 41919 313 41953
rect 347 41919 363 41953
rect 489 41919 505 41953
rect 539 41919 555 41953
rect 681 41919 697 41953
rect 731 41919 747 41953
rect 873 41919 889 41953
rect 923 41919 939 41953
rect 1065 41919 1081 41953
rect 1115 41919 1131 41953
rect 1257 41919 1273 41953
rect 1307 41919 1323 41953
rect 199 41885 233 41919
rect 1387 41885 1421 41893
rect 199 41817 233 41851
rect 199 41749 233 41783
rect 199 41681 233 41715
rect 199 41613 233 41647
rect 313 41854 347 41875
rect 313 41786 347 41790
rect 313 41680 347 41684
rect 313 41595 347 41616
rect 409 41854 443 41875
rect 409 41786 443 41790
rect 409 41680 443 41684
rect 409 41595 443 41616
rect 505 41854 539 41875
rect 505 41786 539 41790
rect 505 41680 539 41684
rect 505 41595 539 41616
rect 601 41854 635 41875
rect 601 41786 635 41790
rect 601 41680 635 41684
rect 601 41595 635 41616
rect 697 41854 731 41875
rect 697 41786 731 41790
rect 697 41680 731 41684
rect 697 41595 731 41616
rect 793 41854 827 41875
rect 793 41786 827 41790
rect 793 41680 827 41684
rect 793 41595 827 41616
rect 889 41854 923 41875
rect 889 41786 923 41790
rect 889 41680 923 41684
rect 889 41595 923 41616
rect 985 41854 1019 41875
rect 985 41786 1019 41790
rect 985 41680 1019 41684
rect 985 41595 1019 41616
rect 1081 41854 1115 41875
rect 1081 41786 1115 41790
rect 1081 41680 1115 41684
rect 1081 41595 1115 41616
rect 1177 41854 1211 41875
rect 1177 41786 1211 41790
rect 1177 41680 1211 41684
rect 1177 41595 1211 41616
rect 1273 41854 1307 41875
rect 1273 41786 1307 41790
rect 1273 41680 1307 41684
rect 1273 41595 1307 41616
rect 1387 41817 1421 41821
rect 1387 41711 1421 41715
rect 1387 41639 1421 41647
rect 199 41511 233 41579
rect 1387 41511 1421 41579
rect 199 41477 317 41511
rect 351 41477 385 41511
rect 419 41477 453 41511
rect 487 41477 521 41511
rect 555 41477 589 41511
rect 623 41477 657 41511
rect 691 41477 725 41511
rect 759 41477 793 41511
rect 827 41477 861 41511
rect 895 41477 929 41511
rect 963 41477 997 41511
rect 1031 41477 1065 41511
rect 1099 41477 1133 41511
rect 1167 41477 1201 41511
rect 1235 41477 1269 41511
rect 1303 41477 1421 41511
rect 2352 42025 2470 42059
rect 2504 42025 2538 42059
rect 2572 42025 2606 42059
rect 2640 42025 2674 42059
rect 2708 42025 2742 42059
rect 2776 42025 2810 42059
rect 2844 42025 2878 42059
rect 2912 42025 2946 42059
rect 2980 42025 3014 42059
rect 3048 42025 3082 42059
rect 3116 42025 3150 42059
rect 3184 42025 3218 42059
rect 3252 42025 3286 42059
rect 3320 42025 3354 42059
rect 3388 42025 3422 42059
rect 3456 42025 3574 42059
rect 2352 41957 2386 42025
rect 3540 41957 3574 42025
rect 2450 41923 2466 41957
rect 2500 41923 2516 41957
rect 2642 41923 2658 41957
rect 2692 41923 2708 41957
rect 2834 41923 2850 41957
rect 2884 41923 2900 41957
rect 3026 41923 3042 41957
rect 3076 41923 3092 41957
rect 3218 41923 3234 41957
rect 3268 41923 3284 41957
rect 3410 41923 3426 41957
rect 3460 41923 3476 41957
rect 2352 41889 2386 41923
rect 3540 41889 3574 41897
rect 2352 41821 2386 41855
rect 2352 41753 2386 41787
rect 2352 41685 2386 41719
rect 2352 41617 2386 41651
rect 2466 41858 2500 41879
rect 2466 41790 2500 41794
rect 2466 41684 2500 41688
rect 2466 41599 2500 41620
rect 2562 41858 2596 41879
rect 2562 41790 2596 41794
rect 2562 41684 2596 41688
rect 2562 41599 2596 41620
rect 2658 41858 2692 41879
rect 2658 41790 2692 41794
rect 2658 41684 2692 41688
rect 2658 41599 2692 41620
rect 2754 41858 2788 41879
rect 2754 41790 2788 41794
rect 2754 41684 2788 41688
rect 2754 41599 2788 41620
rect 2850 41858 2884 41879
rect 2850 41790 2884 41794
rect 2850 41684 2884 41688
rect 2850 41599 2884 41620
rect 2946 41858 2980 41879
rect 2946 41790 2980 41794
rect 2946 41684 2980 41688
rect 2946 41599 2980 41620
rect 3042 41858 3076 41879
rect 3042 41790 3076 41794
rect 3042 41684 3076 41688
rect 3042 41599 3076 41620
rect 3138 41858 3172 41879
rect 3138 41790 3172 41794
rect 3138 41684 3172 41688
rect 3138 41599 3172 41620
rect 3234 41858 3268 41879
rect 3234 41790 3268 41794
rect 3234 41684 3268 41688
rect 3234 41599 3268 41620
rect 3330 41858 3364 41879
rect 3330 41790 3364 41794
rect 3330 41684 3364 41688
rect 3330 41599 3364 41620
rect 3426 41858 3460 41879
rect 3426 41790 3460 41794
rect 3426 41684 3460 41688
rect 3426 41599 3460 41620
rect 3540 41821 3574 41825
rect 3540 41715 3574 41719
rect 3540 41643 3574 41651
rect 2352 41515 2386 41583
rect 3540 41515 3574 41583
rect 2352 41481 2470 41515
rect 2504 41481 2538 41515
rect 2572 41481 2606 41515
rect 2640 41481 2674 41515
rect 2708 41481 2742 41515
rect 2776 41481 2810 41515
rect 2844 41481 2878 41515
rect 2912 41481 2946 41515
rect 2980 41481 3014 41515
rect 3048 41481 3082 41515
rect 3116 41481 3150 41515
rect 3184 41481 3218 41515
rect 3252 41481 3286 41515
rect 3320 41481 3354 41515
rect 3388 41481 3422 41515
rect 3456 41481 3574 41515
rect 3873 42025 3991 42059
rect 4025 42025 4059 42059
rect 4093 42025 4127 42059
rect 4161 42025 4195 42059
rect 4229 42025 4263 42059
rect 4297 42025 4331 42059
rect 4365 42025 4399 42059
rect 4433 42025 4467 42059
rect 4501 42025 4535 42059
rect 4569 42025 4603 42059
rect 4637 42025 4671 42059
rect 4705 42025 4739 42059
rect 4773 42025 4807 42059
rect 4841 42025 4875 42059
rect 4909 42025 4943 42059
rect 4977 42025 5095 42059
rect 3873 41957 3907 42025
rect 5061 41957 5095 42025
rect 3971 41923 3987 41957
rect 4021 41923 4037 41957
rect 4163 41923 4179 41957
rect 4213 41923 4229 41957
rect 4355 41923 4371 41957
rect 4405 41923 4421 41957
rect 4547 41923 4563 41957
rect 4597 41923 4613 41957
rect 4739 41923 4755 41957
rect 4789 41923 4805 41957
rect 4931 41923 4947 41957
rect 4981 41923 4997 41957
rect 3873 41889 3907 41923
rect 5061 41889 5095 41897
rect 3873 41821 3907 41855
rect 3873 41753 3907 41787
rect 3873 41685 3907 41719
rect 3873 41617 3907 41651
rect 3987 41858 4021 41879
rect 3987 41790 4021 41794
rect 3987 41684 4021 41688
rect 3987 41599 4021 41620
rect 4083 41858 4117 41879
rect 4083 41790 4117 41794
rect 4083 41684 4117 41688
rect 4083 41599 4117 41620
rect 4179 41858 4213 41879
rect 4179 41790 4213 41794
rect 4179 41684 4213 41688
rect 4179 41599 4213 41620
rect 4275 41858 4309 41879
rect 4275 41790 4309 41794
rect 4275 41684 4309 41688
rect 4275 41599 4309 41620
rect 4371 41858 4405 41879
rect 4371 41790 4405 41794
rect 4371 41684 4405 41688
rect 4371 41599 4405 41620
rect 4467 41858 4501 41879
rect 4467 41790 4501 41794
rect 4467 41684 4501 41688
rect 4467 41599 4501 41620
rect 4563 41858 4597 41879
rect 4563 41790 4597 41794
rect 4563 41684 4597 41688
rect 4563 41599 4597 41620
rect 4659 41858 4693 41879
rect 4659 41790 4693 41794
rect 4659 41684 4693 41688
rect 4659 41599 4693 41620
rect 4755 41858 4789 41879
rect 4755 41790 4789 41794
rect 4755 41684 4789 41688
rect 4755 41599 4789 41620
rect 4851 41858 4885 41879
rect 4851 41790 4885 41794
rect 4851 41684 4885 41688
rect 4851 41599 4885 41620
rect 4947 41858 4981 41879
rect 4947 41790 4981 41794
rect 4947 41684 4981 41688
rect 4947 41599 4981 41620
rect 5061 41821 5095 41825
rect 5061 41715 5095 41719
rect 5274 41692 5303 41726
rect 5337 41692 5395 41726
rect 5429 41692 5487 41726
rect 5521 41692 5550 41726
rect 5061 41643 5095 41651
rect 3873 41515 3907 41583
rect 5061 41515 5095 41583
rect 3873 41481 3991 41515
rect 4025 41481 4059 41515
rect 4093 41481 4127 41515
rect 4161 41481 4195 41515
rect 4229 41481 4263 41515
rect 4297 41481 4331 41515
rect 4365 41481 4399 41515
rect 4433 41481 4467 41515
rect 4501 41481 4535 41515
rect 4569 41481 4603 41515
rect 4637 41481 4671 41515
rect 4705 41481 4739 41515
rect 4773 41481 4807 41515
rect 4841 41481 4875 41515
rect 4909 41481 4943 41515
rect 4977 41481 5095 41515
rect 5340 41650 5406 41658
rect 5340 41616 5356 41650
rect 5390 41616 5406 41650
rect 5340 41582 5406 41616
rect 5340 41548 5356 41582
rect 5390 41548 5406 41582
rect 5340 41514 5406 41548
rect 5340 41480 5356 41514
rect 5390 41480 5406 41514
rect 5340 41462 5406 41480
rect 5440 41650 5482 41692
rect 5474 41616 5482 41650
rect 5440 41582 5482 41616
rect 5474 41548 5482 41582
rect 5440 41514 5482 41548
rect 5474 41480 5482 41514
rect 5440 41464 5482 41480
rect 5340 41412 5386 41462
rect 199 41369 317 41403
rect 351 41369 385 41403
rect 419 41369 453 41403
rect 487 41369 521 41403
rect 555 41369 589 41403
rect 623 41369 657 41403
rect 691 41369 725 41403
rect 759 41369 793 41403
rect 827 41369 861 41403
rect 895 41369 929 41403
rect 963 41369 997 41403
rect 1031 41369 1065 41403
rect 1099 41369 1133 41403
rect 1167 41369 1201 41403
rect 1235 41369 1269 41403
rect 1303 41369 1421 41403
rect 199 41293 233 41369
rect 1387 41298 1421 41369
rect 199 41225 233 41259
rect 199 41157 233 41191
rect 313 41256 347 41295
rect 313 41183 347 41222
rect 409 41256 443 41295
rect 409 41183 443 41222
rect 505 41256 539 41295
rect 505 41183 539 41222
rect 601 41256 635 41295
rect 601 41183 635 41222
rect 697 41256 731 41295
rect 697 41183 731 41222
rect 793 41256 827 41295
rect 793 41183 827 41222
rect 889 41256 923 41295
rect 889 41183 923 41222
rect 985 41256 1019 41295
rect 985 41183 1019 41222
rect 1081 41256 1115 41295
rect 1081 41183 1115 41222
rect 1177 41256 1211 41295
rect 1177 41183 1211 41222
rect 1273 41256 1307 41295
rect 1273 41183 1307 41222
rect 1387 41226 1421 41259
rect 1387 41157 1421 41191
rect 199 41047 233 41123
rect 297 41111 313 41145
rect 347 41111 363 41145
rect 489 41111 505 41145
rect 539 41111 555 41145
rect 681 41111 697 41145
rect 731 41111 747 41145
rect 873 41111 889 41145
rect 923 41111 939 41145
rect 1065 41111 1081 41145
rect 1115 41111 1131 41145
rect 1257 41111 1273 41145
rect 1307 41111 1323 41145
rect 1387 41047 1421 41120
rect 199 41013 317 41047
rect 351 41013 385 41047
rect 419 41013 453 41047
rect 487 41013 521 41047
rect 555 41013 589 41047
rect 623 41013 657 41047
rect 691 41013 725 41047
rect 759 41013 793 41047
rect 827 41013 861 41047
rect 895 41013 929 41047
rect 963 41013 997 41047
rect 1031 41013 1065 41047
rect 1099 41013 1133 41047
rect 1167 41013 1201 41047
rect 1235 41013 1269 41047
rect 1303 41013 1421 41047
rect 2352 41373 2470 41407
rect 2504 41373 2538 41407
rect 2572 41373 2606 41407
rect 2640 41373 2674 41407
rect 2708 41373 2742 41407
rect 2776 41373 2810 41407
rect 2844 41373 2878 41407
rect 2912 41373 2946 41407
rect 2980 41373 3014 41407
rect 3048 41373 3082 41407
rect 3116 41373 3150 41407
rect 3184 41373 3218 41407
rect 3252 41373 3286 41407
rect 3320 41373 3354 41407
rect 3388 41373 3422 41407
rect 3456 41373 3574 41407
rect 2352 41297 2386 41373
rect 3540 41302 3574 41373
rect 3873 41373 3991 41407
rect 4025 41373 4059 41407
rect 4093 41373 4127 41407
rect 4161 41373 4195 41407
rect 4229 41373 4263 41407
rect 4297 41373 4331 41407
rect 4365 41373 4399 41407
rect 4433 41373 4467 41407
rect 4501 41373 4535 41407
rect 4569 41373 4603 41407
rect 4637 41373 4671 41407
rect 4705 41373 4739 41407
rect 4773 41373 4807 41407
rect 4841 41373 4875 41407
rect 4909 41373 4943 41407
rect 4977 41373 5095 41407
rect 3675 41337 3691 41371
rect 3725 41337 3741 41371
rect 2352 41229 2386 41263
rect 2352 41161 2386 41195
rect 2466 41260 2500 41299
rect 2466 41187 2500 41226
rect 2562 41260 2596 41299
rect 2562 41187 2596 41226
rect 2658 41260 2692 41299
rect 2658 41187 2692 41226
rect 2754 41260 2788 41299
rect 2754 41187 2788 41226
rect 2850 41260 2884 41299
rect 2850 41187 2884 41226
rect 2946 41260 2980 41299
rect 2946 41187 2980 41226
rect 3042 41260 3076 41299
rect 3042 41187 3076 41226
rect 3138 41260 3172 41299
rect 3138 41187 3172 41226
rect 3234 41260 3268 41299
rect 3234 41187 3268 41226
rect 3330 41260 3364 41299
rect 3330 41187 3364 41226
rect 3426 41260 3460 41299
rect 3426 41187 3460 41226
rect 3540 41230 3574 41263
rect 3647 41287 3681 41303
rect 3647 41195 3681 41211
rect 3735 41287 3769 41303
rect 3735 41195 3769 41211
rect 3873 41297 3907 41373
rect 5061 41302 5095 41373
rect 3873 41229 3907 41263
rect 3540 41161 3574 41195
rect 2352 41051 2386 41127
rect 2450 41115 2466 41149
rect 2500 41115 2516 41149
rect 2642 41115 2658 41149
rect 2692 41115 2708 41149
rect 2834 41115 2850 41149
rect 2884 41115 2900 41149
rect 3026 41115 3042 41149
rect 3076 41115 3092 41149
rect 3218 41115 3234 41149
rect 3268 41115 3284 41149
rect 3410 41115 3426 41149
rect 3460 41115 3476 41149
rect 3540 41051 3574 41124
rect 2352 41017 2470 41051
rect 2504 41017 2538 41051
rect 2572 41017 2606 41051
rect 2640 41017 2674 41051
rect 2708 41017 2742 41051
rect 2776 41017 2810 41051
rect 2844 41017 2878 41051
rect 2912 41017 2946 41051
rect 2980 41017 3014 41051
rect 3048 41017 3082 41051
rect 3116 41017 3150 41051
rect 3184 41017 3218 41051
rect 3252 41017 3286 41051
rect 3320 41017 3354 41051
rect 3388 41017 3422 41051
rect 3456 41017 3574 41051
rect 3873 41161 3907 41195
rect 3987 41260 4021 41299
rect 3987 41187 4021 41226
rect 4083 41260 4117 41299
rect 4083 41187 4117 41226
rect 4179 41260 4213 41299
rect 4179 41187 4213 41226
rect 4275 41260 4309 41299
rect 4275 41187 4309 41226
rect 4371 41260 4405 41299
rect 4371 41187 4405 41226
rect 4467 41260 4501 41299
rect 4467 41187 4501 41226
rect 4563 41260 4597 41299
rect 4563 41187 4597 41226
rect 4659 41260 4693 41299
rect 4659 41187 4693 41226
rect 4755 41260 4789 41299
rect 4755 41187 4789 41226
rect 4851 41260 4885 41299
rect 4851 41187 4885 41226
rect 4947 41260 4981 41299
rect 4947 41187 4981 41226
rect 5061 41230 5095 41263
rect 5340 41378 5348 41412
rect 5382 41378 5386 41412
rect 5420 41417 5486 41428
rect 5420 41414 5450 41417
rect 5420 41380 5436 41414
rect 5484 41383 5486 41417
rect 5470 41380 5486 41383
rect 5340 41342 5386 41378
rect 5340 41330 5406 41342
rect 5340 41296 5356 41330
rect 5390 41296 5406 41330
rect 5340 41262 5406 41296
rect 5340 41228 5356 41262
rect 5390 41228 5406 41262
rect 5340 41216 5406 41228
rect 5440 41330 5486 41346
rect 5474 41296 5486 41330
rect 5440 41262 5486 41296
rect 5474 41228 5486 41262
rect 5061 41161 5095 41195
rect 5440 41182 5486 41228
rect 3873 41051 3907 41127
rect 3971 41115 3987 41149
rect 4021 41115 4037 41149
rect 4163 41115 4179 41149
rect 4213 41115 4229 41149
rect 4355 41115 4371 41149
rect 4405 41115 4421 41149
rect 4547 41115 4563 41149
rect 4597 41115 4613 41149
rect 4739 41115 4755 41149
rect 4789 41115 4805 41149
rect 4931 41115 4947 41149
rect 4981 41115 4997 41149
rect 5274 41148 5303 41182
rect 5337 41148 5395 41182
rect 5429 41148 5487 41182
rect 5521 41148 5550 41182
rect 5061 41051 5095 41124
rect 3873 41017 3991 41051
rect 4025 41017 4059 41051
rect 4093 41017 4127 41051
rect 4161 41017 4195 41051
rect 4229 41017 4263 41051
rect 4297 41017 4331 41051
rect 4365 41017 4399 41051
rect 4433 41017 4467 41051
rect 4501 41017 4535 41051
rect 4569 41017 4603 41051
rect 4637 41017 4671 41051
rect 4705 41017 4739 41051
rect 4773 41017 4807 41051
rect 4841 41017 4875 41051
rect 4909 41017 4943 41051
rect 4977 41017 5095 41051
rect 199 40734 317 40768
rect 351 40734 385 40768
rect 419 40734 453 40768
rect 487 40734 521 40768
rect 555 40734 589 40768
rect 623 40734 657 40768
rect 691 40734 725 40768
rect 759 40734 793 40768
rect 827 40734 861 40768
rect 895 40734 929 40768
rect 963 40734 997 40768
rect 1031 40734 1065 40768
rect 1099 40734 1133 40768
rect 1167 40734 1201 40768
rect 1235 40734 1269 40768
rect 1303 40734 1421 40768
rect 199 40666 233 40734
rect 1387 40666 1421 40734
rect 297 40632 313 40666
rect 347 40632 363 40666
rect 489 40632 505 40666
rect 539 40632 555 40666
rect 681 40632 697 40666
rect 731 40632 747 40666
rect 873 40632 889 40666
rect 923 40632 939 40666
rect 1065 40632 1081 40666
rect 1115 40632 1131 40666
rect 1257 40632 1273 40666
rect 1307 40632 1323 40666
rect 199 40598 233 40632
rect 1387 40598 1421 40606
rect 199 40530 233 40564
rect 199 40462 233 40496
rect 199 40394 233 40428
rect 199 40326 233 40360
rect 313 40567 347 40588
rect 313 40499 347 40503
rect 313 40393 347 40397
rect 313 40308 347 40329
rect 409 40567 443 40588
rect 409 40499 443 40503
rect 409 40393 443 40397
rect 409 40308 443 40329
rect 505 40567 539 40588
rect 505 40499 539 40503
rect 505 40393 539 40397
rect 505 40308 539 40329
rect 601 40567 635 40588
rect 601 40499 635 40503
rect 601 40393 635 40397
rect 601 40308 635 40329
rect 697 40567 731 40588
rect 697 40499 731 40503
rect 697 40393 731 40397
rect 697 40308 731 40329
rect 793 40567 827 40588
rect 793 40499 827 40503
rect 793 40393 827 40397
rect 793 40308 827 40329
rect 889 40567 923 40588
rect 889 40499 923 40503
rect 889 40393 923 40397
rect 889 40308 923 40329
rect 985 40567 1019 40588
rect 985 40499 1019 40503
rect 985 40393 1019 40397
rect 985 40308 1019 40329
rect 1081 40567 1115 40588
rect 1081 40499 1115 40503
rect 1081 40393 1115 40397
rect 1081 40308 1115 40329
rect 1177 40567 1211 40588
rect 1177 40499 1211 40503
rect 1177 40393 1211 40397
rect 1177 40308 1211 40329
rect 1273 40567 1307 40588
rect 1273 40499 1307 40503
rect 1273 40393 1307 40397
rect 1273 40308 1307 40329
rect 1387 40530 1421 40534
rect 1387 40424 1421 40428
rect 1387 40352 1421 40360
rect 199 40224 233 40292
rect 1387 40224 1421 40292
rect 199 40190 317 40224
rect 351 40190 385 40224
rect 419 40190 453 40224
rect 487 40190 521 40224
rect 555 40190 589 40224
rect 623 40190 657 40224
rect 691 40190 725 40224
rect 759 40190 793 40224
rect 827 40190 861 40224
rect 895 40190 929 40224
rect 963 40190 997 40224
rect 1031 40190 1065 40224
rect 1099 40190 1133 40224
rect 1167 40190 1201 40224
rect 1235 40190 1269 40224
rect 1303 40190 1421 40224
rect 2352 40738 2470 40772
rect 2504 40738 2538 40772
rect 2572 40738 2606 40772
rect 2640 40738 2674 40772
rect 2708 40738 2742 40772
rect 2776 40738 2810 40772
rect 2844 40738 2878 40772
rect 2912 40738 2946 40772
rect 2980 40738 3014 40772
rect 3048 40738 3082 40772
rect 3116 40738 3150 40772
rect 3184 40738 3218 40772
rect 3252 40738 3286 40772
rect 3320 40738 3354 40772
rect 3388 40738 3422 40772
rect 3456 40738 3574 40772
rect 2352 40670 2386 40738
rect 3540 40670 3574 40738
rect 2450 40636 2466 40670
rect 2500 40636 2516 40670
rect 2642 40636 2658 40670
rect 2692 40636 2708 40670
rect 2834 40636 2850 40670
rect 2884 40636 2900 40670
rect 3026 40636 3042 40670
rect 3076 40636 3092 40670
rect 3218 40636 3234 40670
rect 3268 40636 3284 40670
rect 3410 40636 3426 40670
rect 3460 40636 3476 40670
rect 2352 40602 2386 40636
rect 3540 40602 3574 40610
rect 2352 40534 2386 40568
rect 2352 40466 2386 40500
rect 2352 40398 2386 40432
rect 2352 40330 2386 40364
rect 2466 40571 2500 40592
rect 2466 40503 2500 40507
rect 2466 40397 2500 40401
rect 2466 40312 2500 40333
rect 2562 40571 2596 40592
rect 2562 40503 2596 40507
rect 2562 40397 2596 40401
rect 2562 40312 2596 40333
rect 2658 40571 2692 40592
rect 2658 40503 2692 40507
rect 2658 40397 2692 40401
rect 2658 40312 2692 40333
rect 2754 40571 2788 40592
rect 2754 40503 2788 40507
rect 2754 40397 2788 40401
rect 2754 40312 2788 40333
rect 2850 40571 2884 40592
rect 2850 40503 2884 40507
rect 2850 40397 2884 40401
rect 2850 40312 2884 40333
rect 2946 40571 2980 40592
rect 2946 40503 2980 40507
rect 2946 40397 2980 40401
rect 2946 40312 2980 40333
rect 3042 40571 3076 40592
rect 3042 40503 3076 40507
rect 3042 40397 3076 40401
rect 3042 40312 3076 40333
rect 3138 40571 3172 40592
rect 3138 40503 3172 40507
rect 3138 40397 3172 40401
rect 3138 40312 3172 40333
rect 3234 40571 3268 40592
rect 3234 40503 3268 40507
rect 3234 40397 3268 40401
rect 3234 40312 3268 40333
rect 3330 40571 3364 40592
rect 3330 40503 3364 40507
rect 3330 40397 3364 40401
rect 3330 40312 3364 40333
rect 3426 40571 3460 40592
rect 3426 40503 3460 40507
rect 3426 40397 3460 40401
rect 3426 40312 3460 40333
rect 3540 40534 3574 40538
rect 3540 40428 3574 40432
rect 3540 40356 3574 40364
rect 2352 40228 2386 40296
rect 3540 40228 3574 40296
rect 2352 40194 2470 40228
rect 2504 40194 2538 40228
rect 2572 40194 2606 40228
rect 2640 40194 2674 40228
rect 2708 40194 2742 40228
rect 2776 40194 2810 40228
rect 2844 40194 2878 40228
rect 2912 40194 2946 40228
rect 2980 40194 3014 40228
rect 3048 40194 3082 40228
rect 3116 40194 3150 40228
rect 3184 40194 3218 40228
rect 3252 40194 3286 40228
rect 3320 40194 3354 40228
rect 3388 40194 3422 40228
rect 3456 40194 3574 40228
rect 3873 40738 3991 40772
rect 4025 40738 4059 40772
rect 4093 40738 4127 40772
rect 4161 40738 4195 40772
rect 4229 40738 4263 40772
rect 4297 40738 4331 40772
rect 4365 40738 4399 40772
rect 4433 40738 4467 40772
rect 4501 40738 4535 40772
rect 4569 40738 4603 40772
rect 4637 40738 4671 40772
rect 4705 40738 4739 40772
rect 4773 40738 4807 40772
rect 4841 40738 4875 40772
rect 4909 40738 4943 40772
rect 4977 40738 5095 40772
rect 3873 40670 3907 40738
rect 5061 40670 5095 40738
rect 3971 40636 3987 40670
rect 4021 40636 4037 40670
rect 4163 40636 4179 40670
rect 4213 40636 4229 40670
rect 4355 40636 4371 40670
rect 4405 40636 4421 40670
rect 4547 40636 4563 40670
rect 4597 40636 4613 40670
rect 4739 40636 4755 40670
rect 4789 40636 4805 40670
rect 4931 40636 4947 40670
rect 4981 40636 4997 40670
rect 3873 40602 3907 40636
rect 5061 40602 5095 40610
rect 3873 40534 3907 40568
rect 3873 40466 3907 40500
rect 3873 40398 3907 40432
rect 3873 40330 3907 40364
rect 3987 40571 4021 40592
rect 3987 40503 4021 40507
rect 3987 40397 4021 40401
rect 3987 40312 4021 40333
rect 4083 40571 4117 40592
rect 4083 40503 4117 40507
rect 4083 40397 4117 40401
rect 4083 40312 4117 40333
rect 4179 40571 4213 40592
rect 4179 40503 4213 40507
rect 4179 40397 4213 40401
rect 4179 40312 4213 40333
rect 4275 40571 4309 40592
rect 4275 40503 4309 40507
rect 4275 40397 4309 40401
rect 4275 40312 4309 40333
rect 4371 40571 4405 40592
rect 4371 40503 4405 40507
rect 4371 40397 4405 40401
rect 4371 40312 4405 40333
rect 4467 40571 4501 40592
rect 4467 40503 4501 40507
rect 4467 40397 4501 40401
rect 4467 40312 4501 40333
rect 4563 40571 4597 40592
rect 4563 40503 4597 40507
rect 4563 40397 4597 40401
rect 4563 40312 4597 40333
rect 4659 40571 4693 40592
rect 4659 40503 4693 40507
rect 4659 40397 4693 40401
rect 4659 40312 4693 40333
rect 4755 40571 4789 40592
rect 4755 40503 4789 40507
rect 4755 40397 4789 40401
rect 4755 40312 4789 40333
rect 4851 40571 4885 40592
rect 4851 40503 4885 40507
rect 4851 40397 4885 40401
rect 4851 40312 4885 40333
rect 4947 40571 4981 40592
rect 4947 40503 4981 40507
rect 4947 40397 4981 40401
rect 4947 40312 4981 40333
rect 5061 40534 5095 40538
rect 5061 40428 5095 40432
rect 5274 40405 5303 40439
rect 5337 40405 5395 40439
rect 5429 40405 5487 40439
rect 5521 40405 5550 40439
rect 5061 40356 5095 40364
rect 3873 40228 3907 40296
rect 5061 40228 5095 40296
rect 3873 40194 3991 40228
rect 4025 40194 4059 40228
rect 4093 40194 4127 40228
rect 4161 40194 4195 40228
rect 4229 40194 4263 40228
rect 4297 40194 4331 40228
rect 4365 40194 4399 40228
rect 4433 40194 4467 40228
rect 4501 40194 4535 40228
rect 4569 40194 4603 40228
rect 4637 40194 4671 40228
rect 4705 40194 4739 40228
rect 4773 40194 4807 40228
rect 4841 40194 4875 40228
rect 4909 40194 4943 40228
rect 4977 40194 5095 40228
rect 5340 40363 5406 40371
rect 5340 40329 5356 40363
rect 5390 40329 5406 40363
rect 5340 40295 5406 40329
rect 5340 40261 5356 40295
rect 5390 40261 5406 40295
rect 5340 40227 5406 40261
rect 5340 40193 5356 40227
rect 5390 40193 5406 40227
rect 5340 40175 5406 40193
rect 5440 40363 5482 40405
rect 5474 40329 5482 40363
rect 5440 40295 5482 40329
rect 5474 40261 5482 40295
rect 5440 40227 5482 40261
rect 5474 40193 5482 40227
rect 5440 40177 5482 40193
rect 5340 40125 5386 40175
rect 199 40082 317 40116
rect 351 40082 385 40116
rect 419 40082 453 40116
rect 487 40082 521 40116
rect 555 40082 589 40116
rect 623 40082 657 40116
rect 691 40082 725 40116
rect 759 40082 793 40116
rect 827 40082 861 40116
rect 895 40082 929 40116
rect 963 40082 997 40116
rect 1031 40082 1065 40116
rect 1099 40082 1133 40116
rect 1167 40082 1201 40116
rect 1235 40082 1269 40116
rect 1303 40082 1421 40116
rect 199 40006 233 40082
rect 1387 40011 1421 40082
rect 199 39938 233 39972
rect 199 39870 233 39904
rect 313 39969 347 40008
rect 313 39896 347 39935
rect 409 39969 443 40008
rect 409 39896 443 39935
rect 505 39969 539 40008
rect 505 39896 539 39935
rect 601 39969 635 40008
rect 601 39896 635 39935
rect 697 39969 731 40008
rect 697 39896 731 39935
rect 793 39969 827 40008
rect 793 39896 827 39935
rect 889 39969 923 40008
rect 889 39896 923 39935
rect 985 39969 1019 40008
rect 985 39896 1019 39935
rect 1081 39969 1115 40008
rect 1081 39896 1115 39935
rect 1177 39969 1211 40008
rect 1177 39896 1211 39935
rect 1273 39969 1307 40008
rect 1273 39896 1307 39935
rect 1387 39939 1421 39972
rect 1387 39870 1421 39904
rect 199 39760 233 39836
rect 297 39824 313 39858
rect 347 39824 363 39858
rect 489 39824 505 39858
rect 539 39824 555 39858
rect 681 39824 697 39858
rect 731 39824 747 39858
rect 873 39824 889 39858
rect 923 39824 939 39858
rect 1065 39824 1081 39858
rect 1115 39824 1131 39858
rect 1257 39824 1273 39858
rect 1307 39824 1323 39858
rect 1387 39760 1421 39833
rect 199 39726 317 39760
rect 351 39726 385 39760
rect 419 39726 453 39760
rect 487 39726 521 39760
rect 555 39726 589 39760
rect 623 39726 657 39760
rect 691 39726 725 39760
rect 759 39726 793 39760
rect 827 39726 861 39760
rect 895 39726 929 39760
rect 963 39726 997 39760
rect 1031 39726 1065 39760
rect 1099 39726 1133 39760
rect 1167 39726 1201 39760
rect 1235 39726 1269 39760
rect 1303 39726 1421 39760
rect 2352 40086 2470 40120
rect 2504 40086 2538 40120
rect 2572 40086 2606 40120
rect 2640 40086 2674 40120
rect 2708 40086 2742 40120
rect 2776 40086 2810 40120
rect 2844 40086 2878 40120
rect 2912 40086 2946 40120
rect 2980 40086 3014 40120
rect 3048 40086 3082 40120
rect 3116 40086 3150 40120
rect 3184 40086 3218 40120
rect 3252 40086 3286 40120
rect 3320 40086 3354 40120
rect 3388 40086 3422 40120
rect 3456 40086 3574 40120
rect 2352 40010 2386 40086
rect 3540 40015 3574 40086
rect 3873 40086 3991 40120
rect 4025 40086 4059 40120
rect 4093 40086 4127 40120
rect 4161 40086 4195 40120
rect 4229 40086 4263 40120
rect 4297 40086 4331 40120
rect 4365 40086 4399 40120
rect 4433 40086 4467 40120
rect 4501 40086 4535 40120
rect 4569 40086 4603 40120
rect 4637 40086 4671 40120
rect 4705 40086 4739 40120
rect 4773 40086 4807 40120
rect 4841 40086 4875 40120
rect 4909 40086 4943 40120
rect 4977 40086 5095 40120
rect 3675 40050 3691 40084
rect 3725 40050 3741 40084
rect 2352 39942 2386 39976
rect 2352 39874 2386 39908
rect 2466 39973 2500 40012
rect 2466 39900 2500 39939
rect 2562 39973 2596 40012
rect 2562 39900 2596 39939
rect 2658 39973 2692 40012
rect 2658 39900 2692 39939
rect 2754 39973 2788 40012
rect 2754 39900 2788 39939
rect 2850 39973 2884 40012
rect 2850 39900 2884 39939
rect 2946 39973 2980 40012
rect 2946 39900 2980 39939
rect 3042 39973 3076 40012
rect 3042 39900 3076 39939
rect 3138 39973 3172 40012
rect 3138 39900 3172 39939
rect 3234 39973 3268 40012
rect 3234 39900 3268 39939
rect 3330 39973 3364 40012
rect 3330 39900 3364 39939
rect 3426 39973 3460 40012
rect 3426 39900 3460 39939
rect 3540 39943 3574 39976
rect 3647 40000 3681 40016
rect 3647 39908 3681 39924
rect 3735 40000 3769 40016
rect 3735 39908 3769 39924
rect 3873 40010 3907 40086
rect 5061 40015 5095 40086
rect 3873 39942 3907 39976
rect 3540 39874 3574 39908
rect 2352 39764 2386 39840
rect 2450 39828 2466 39862
rect 2500 39828 2516 39862
rect 2642 39828 2658 39862
rect 2692 39828 2708 39862
rect 2834 39828 2850 39862
rect 2884 39828 2900 39862
rect 3026 39828 3042 39862
rect 3076 39828 3092 39862
rect 3218 39828 3234 39862
rect 3268 39828 3284 39862
rect 3410 39828 3426 39862
rect 3460 39828 3476 39862
rect 3540 39764 3574 39837
rect 2352 39730 2470 39764
rect 2504 39730 2538 39764
rect 2572 39730 2606 39764
rect 2640 39730 2674 39764
rect 2708 39730 2742 39764
rect 2776 39730 2810 39764
rect 2844 39730 2878 39764
rect 2912 39730 2946 39764
rect 2980 39730 3014 39764
rect 3048 39730 3082 39764
rect 3116 39730 3150 39764
rect 3184 39730 3218 39764
rect 3252 39730 3286 39764
rect 3320 39730 3354 39764
rect 3388 39730 3422 39764
rect 3456 39730 3574 39764
rect 3873 39874 3907 39908
rect 3987 39973 4021 40012
rect 3987 39900 4021 39939
rect 4083 39973 4117 40012
rect 4083 39900 4117 39939
rect 4179 39973 4213 40012
rect 4179 39900 4213 39939
rect 4275 39973 4309 40012
rect 4275 39900 4309 39939
rect 4371 39973 4405 40012
rect 4371 39900 4405 39939
rect 4467 39973 4501 40012
rect 4467 39900 4501 39939
rect 4563 39973 4597 40012
rect 4563 39900 4597 39939
rect 4659 39973 4693 40012
rect 4659 39900 4693 39939
rect 4755 39973 4789 40012
rect 4755 39900 4789 39939
rect 4851 39973 4885 40012
rect 4851 39900 4885 39939
rect 4947 39973 4981 40012
rect 4947 39900 4981 39939
rect 5061 39943 5095 39976
rect 5340 40091 5348 40125
rect 5382 40091 5386 40125
rect 5420 40130 5486 40141
rect 5420 40127 5450 40130
rect 5420 40093 5436 40127
rect 5484 40096 5486 40130
rect 5470 40093 5486 40096
rect 5340 40055 5386 40091
rect 5340 40043 5406 40055
rect 5340 40009 5356 40043
rect 5390 40009 5406 40043
rect 5340 39975 5406 40009
rect 5340 39941 5356 39975
rect 5390 39941 5406 39975
rect 5340 39929 5406 39941
rect 5440 40043 5486 40059
rect 5474 40009 5486 40043
rect 5440 39975 5486 40009
rect 5474 39941 5486 39975
rect 5061 39874 5095 39908
rect 5440 39895 5486 39941
rect 3873 39764 3907 39840
rect 3971 39828 3987 39862
rect 4021 39828 4037 39862
rect 4163 39828 4179 39862
rect 4213 39828 4229 39862
rect 4355 39828 4371 39862
rect 4405 39828 4421 39862
rect 4547 39828 4563 39862
rect 4597 39828 4613 39862
rect 4739 39828 4755 39862
rect 4789 39828 4805 39862
rect 4931 39828 4947 39862
rect 4981 39828 4997 39862
rect 5274 39861 5303 39895
rect 5337 39861 5395 39895
rect 5429 39861 5487 39895
rect 5521 39861 5550 39895
rect 5061 39764 5095 39837
rect 3873 39730 3991 39764
rect 4025 39730 4059 39764
rect 4093 39730 4127 39764
rect 4161 39730 4195 39764
rect 4229 39730 4263 39764
rect 4297 39730 4331 39764
rect 4365 39730 4399 39764
rect 4433 39730 4467 39764
rect 4501 39730 4535 39764
rect 4569 39730 4603 39764
rect 4637 39730 4671 39764
rect 4705 39730 4739 39764
rect 4773 39730 4807 39764
rect 4841 39730 4875 39764
rect 4909 39730 4943 39764
rect 4977 39730 5095 39764
rect 199 39447 317 39481
rect 351 39447 385 39481
rect 419 39447 453 39481
rect 487 39447 521 39481
rect 555 39447 589 39481
rect 623 39447 657 39481
rect 691 39447 725 39481
rect 759 39447 793 39481
rect 827 39447 861 39481
rect 895 39447 929 39481
rect 963 39447 997 39481
rect 1031 39447 1065 39481
rect 1099 39447 1133 39481
rect 1167 39447 1201 39481
rect 1235 39447 1269 39481
rect 1303 39447 1421 39481
rect 199 39379 233 39447
rect 1387 39379 1421 39447
rect 297 39345 313 39379
rect 347 39345 363 39379
rect 489 39345 505 39379
rect 539 39345 555 39379
rect 681 39345 697 39379
rect 731 39345 747 39379
rect 873 39345 889 39379
rect 923 39345 939 39379
rect 1065 39345 1081 39379
rect 1115 39345 1131 39379
rect 1257 39345 1273 39379
rect 1307 39345 1323 39379
rect 199 39311 233 39345
rect 1387 39311 1421 39319
rect 199 39243 233 39277
rect 199 39175 233 39209
rect 199 39107 233 39141
rect 199 39039 233 39073
rect 313 39280 347 39301
rect 313 39212 347 39216
rect 313 39106 347 39110
rect 313 39021 347 39042
rect 409 39280 443 39301
rect 409 39212 443 39216
rect 409 39106 443 39110
rect 409 39021 443 39042
rect 505 39280 539 39301
rect 505 39212 539 39216
rect 505 39106 539 39110
rect 505 39021 539 39042
rect 601 39280 635 39301
rect 601 39212 635 39216
rect 601 39106 635 39110
rect 601 39021 635 39042
rect 697 39280 731 39301
rect 697 39212 731 39216
rect 697 39106 731 39110
rect 697 39021 731 39042
rect 793 39280 827 39301
rect 793 39212 827 39216
rect 793 39106 827 39110
rect 793 39021 827 39042
rect 889 39280 923 39301
rect 889 39212 923 39216
rect 889 39106 923 39110
rect 889 39021 923 39042
rect 985 39280 1019 39301
rect 985 39212 1019 39216
rect 985 39106 1019 39110
rect 985 39021 1019 39042
rect 1081 39280 1115 39301
rect 1081 39212 1115 39216
rect 1081 39106 1115 39110
rect 1081 39021 1115 39042
rect 1177 39280 1211 39301
rect 1177 39212 1211 39216
rect 1177 39106 1211 39110
rect 1177 39021 1211 39042
rect 1273 39280 1307 39301
rect 1273 39212 1307 39216
rect 1273 39106 1307 39110
rect 1273 39021 1307 39042
rect 1387 39243 1421 39247
rect 1387 39137 1421 39141
rect 1387 39065 1421 39073
rect 199 38937 233 39005
rect 1387 38937 1421 39005
rect 199 38903 317 38937
rect 351 38903 385 38937
rect 419 38903 453 38937
rect 487 38903 521 38937
rect 555 38903 589 38937
rect 623 38903 657 38937
rect 691 38903 725 38937
rect 759 38903 793 38937
rect 827 38903 861 38937
rect 895 38903 929 38937
rect 963 38903 997 38937
rect 1031 38903 1065 38937
rect 1099 38903 1133 38937
rect 1167 38903 1201 38937
rect 1235 38903 1269 38937
rect 1303 38903 1421 38937
rect 2352 39451 2470 39485
rect 2504 39451 2538 39485
rect 2572 39451 2606 39485
rect 2640 39451 2674 39485
rect 2708 39451 2742 39485
rect 2776 39451 2810 39485
rect 2844 39451 2878 39485
rect 2912 39451 2946 39485
rect 2980 39451 3014 39485
rect 3048 39451 3082 39485
rect 3116 39451 3150 39485
rect 3184 39451 3218 39485
rect 3252 39451 3286 39485
rect 3320 39451 3354 39485
rect 3388 39451 3422 39485
rect 3456 39451 3574 39485
rect 2352 39383 2386 39451
rect 3540 39383 3574 39451
rect 2450 39349 2466 39383
rect 2500 39349 2516 39383
rect 2642 39349 2658 39383
rect 2692 39349 2708 39383
rect 2834 39349 2850 39383
rect 2884 39349 2900 39383
rect 3026 39349 3042 39383
rect 3076 39349 3092 39383
rect 3218 39349 3234 39383
rect 3268 39349 3284 39383
rect 3410 39349 3426 39383
rect 3460 39349 3476 39383
rect 2352 39315 2386 39349
rect 3540 39315 3574 39323
rect 2352 39247 2386 39281
rect 2352 39179 2386 39213
rect 2352 39111 2386 39145
rect 2352 39043 2386 39077
rect 2466 39284 2500 39305
rect 2466 39216 2500 39220
rect 2466 39110 2500 39114
rect 2466 39025 2500 39046
rect 2562 39284 2596 39305
rect 2562 39216 2596 39220
rect 2562 39110 2596 39114
rect 2562 39025 2596 39046
rect 2658 39284 2692 39305
rect 2658 39216 2692 39220
rect 2658 39110 2692 39114
rect 2658 39025 2692 39046
rect 2754 39284 2788 39305
rect 2754 39216 2788 39220
rect 2754 39110 2788 39114
rect 2754 39025 2788 39046
rect 2850 39284 2884 39305
rect 2850 39216 2884 39220
rect 2850 39110 2884 39114
rect 2850 39025 2884 39046
rect 2946 39284 2980 39305
rect 2946 39216 2980 39220
rect 2946 39110 2980 39114
rect 2946 39025 2980 39046
rect 3042 39284 3076 39305
rect 3042 39216 3076 39220
rect 3042 39110 3076 39114
rect 3042 39025 3076 39046
rect 3138 39284 3172 39305
rect 3138 39216 3172 39220
rect 3138 39110 3172 39114
rect 3138 39025 3172 39046
rect 3234 39284 3268 39305
rect 3234 39216 3268 39220
rect 3234 39110 3268 39114
rect 3234 39025 3268 39046
rect 3330 39284 3364 39305
rect 3330 39216 3364 39220
rect 3330 39110 3364 39114
rect 3330 39025 3364 39046
rect 3426 39284 3460 39305
rect 3426 39216 3460 39220
rect 3426 39110 3460 39114
rect 3426 39025 3460 39046
rect 3540 39247 3574 39251
rect 3540 39141 3574 39145
rect 3540 39069 3574 39077
rect 2352 38941 2386 39009
rect 3540 38941 3574 39009
rect 2352 38907 2470 38941
rect 2504 38907 2538 38941
rect 2572 38907 2606 38941
rect 2640 38907 2674 38941
rect 2708 38907 2742 38941
rect 2776 38907 2810 38941
rect 2844 38907 2878 38941
rect 2912 38907 2946 38941
rect 2980 38907 3014 38941
rect 3048 38907 3082 38941
rect 3116 38907 3150 38941
rect 3184 38907 3218 38941
rect 3252 38907 3286 38941
rect 3320 38907 3354 38941
rect 3388 38907 3422 38941
rect 3456 38907 3574 38941
rect 3873 39451 3991 39485
rect 4025 39451 4059 39485
rect 4093 39451 4127 39485
rect 4161 39451 4195 39485
rect 4229 39451 4263 39485
rect 4297 39451 4331 39485
rect 4365 39451 4399 39485
rect 4433 39451 4467 39485
rect 4501 39451 4535 39485
rect 4569 39451 4603 39485
rect 4637 39451 4671 39485
rect 4705 39451 4739 39485
rect 4773 39451 4807 39485
rect 4841 39451 4875 39485
rect 4909 39451 4943 39485
rect 4977 39451 5095 39485
rect 3873 39383 3907 39451
rect 5061 39383 5095 39451
rect 3971 39349 3987 39383
rect 4021 39349 4037 39383
rect 4163 39349 4179 39383
rect 4213 39349 4229 39383
rect 4355 39349 4371 39383
rect 4405 39349 4421 39383
rect 4547 39349 4563 39383
rect 4597 39349 4613 39383
rect 4739 39349 4755 39383
rect 4789 39349 4805 39383
rect 4931 39349 4947 39383
rect 4981 39349 4997 39383
rect 3873 39315 3907 39349
rect 5061 39315 5095 39323
rect 3873 39247 3907 39281
rect 3873 39179 3907 39213
rect 3873 39111 3907 39145
rect 3873 39043 3907 39077
rect 3987 39284 4021 39305
rect 3987 39216 4021 39220
rect 3987 39110 4021 39114
rect 3987 39025 4021 39046
rect 4083 39284 4117 39305
rect 4083 39216 4117 39220
rect 4083 39110 4117 39114
rect 4083 39025 4117 39046
rect 4179 39284 4213 39305
rect 4179 39216 4213 39220
rect 4179 39110 4213 39114
rect 4179 39025 4213 39046
rect 4275 39284 4309 39305
rect 4275 39216 4309 39220
rect 4275 39110 4309 39114
rect 4275 39025 4309 39046
rect 4371 39284 4405 39305
rect 4371 39216 4405 39220
rect 4371 39110 4405 39114
rect 4371 39025 4405 39046
rect 4467 39284 4501 39305
rect 4467 39216 4501 39220
rect 4467 39110 4501 39114
rect 4467 39025 4501 39046
rect 4563 39284 4597 39305
rect 4563 39216 4597 39220
rect 4563 39110 4597 39114
rect 4563 39025 4597 39046
rect 4659 39284 4693 39305
rect 4659 39216 4693 39220
rect 4659 39110 4693 39114
rect 4659 39025 4693 39046
rect 4755 39284 4789 39305
rect 4755 39216 4789 39220
rect 4755 39110 4789 39114
rect 4755 39025 4789 39046
rect 4851 39284 4885 39305
rect 4851 39216 4885 39220
rect 4851 39110 4885 39114
rect 4851 39025 4885 39046
rect 4947 39284 4981 39305
rect 4947 39216 4981 39220
rect 4947 39110 4981 39114
rect 4947 39025 4981 39046
rect 5061 39247 5095 39251
rect 5061 39141 5095 39145
rect 5274 39118 5303 39152
rect 5337 39118 5395 39152
rect 5429 39118 5487 39152
rect 5521 39118 5550 39152
rect 5061 39069 5095 39077
rect 3873 38941 3907 39009
rect 5061 38941 5095 39009
rect 3873 38907 3991 38941
rect 4025 38907 4059 38941
rect 4093 38907 4127 38941
rect 4161 38907 4195 38941
rect 4229 38907 4263 38941
rect 4297 38907 4331 38941
rect 4365 38907 4399 38941
rect 4433 38907 4467 38941
rect 4501 38907 4535 38941
rect 4569 38907 4603 38941
rect 4637 38907 4671 38941
rect 4705 38907 4739 38941
rect 4773 38907 4807 38941
rect 4841 38907 4875 38941
rect 4909 38907 4943 38941
rect 4977 38907 5095 38941
rect 5340 39076 5406 39084
rect 5340 39042 5356 39076
rect 5390 39042 5406 39076
rect 5340 39008 5406 39042
rect 5340 38974 5356 39008
rect 5390 38974 5406 39008
rect 5340 38940 5406 38974
rect 5340 38906 5356 38940
rect 5390 38906 5406 38940
rect 5340 38888 5406 38906
rect 5440 39076 5482 39118
rect 5474 39042 5482 39076
rect 5440 39008 5482 39042
rect 5474 38974 5482 39008
rect 5440 38940 5482 38974
rect 5474 38906 5482 38940
rect 5440 38890 5482 38906
rect 5340 38838 5386 38888
rect 199 38795 317 38829
rect 351 38795 385 38829
rect 419 38795 453 38829
rect 487 38795 521 38829
rect 555 38795 589 38829
rect 623 38795 657 38829
rect 691 38795 725 38829
rect 759 38795 793 38829
rect 827 38795 861 38829
rect 895 38795 929 38829
rect 963 38795 997 38829
rect 1031 38795 1065 38829
rect 1099 38795 1133 38829
rect 1167 38795 1201 38829
rect 1235 38795 1269 38829
rect 1303 38795 1421 38829
rect 199 38719 233 38795
rect 1387 38724 1421 38795
rect 199 38651 233 38685
rect 199 38583 233 38617
rect 313 38682 347 38721
rect 313 38609 347 38648
rect 409 38682 443 38721
rect 409 38609 443 38648
rect 505 38682 539 38721
rect 505 38609 539 38648
rect 601 38682 635 38721
rect 601 38609 635 38648
rect 697 38682 731 38721
rect 697 38609 731 38648
rect 793 38682 827 38721
rect 793 38609 827 38648
rect 889 38682 923 38721
rect 889 38609 923 38648
rect 985 38682 1019 38721
rect 985 38609 1019 38648
rect 1081 38682 1115 38721
rect 1081 38609 1115 38648
rect 1177 38682 1211 38721
rect 1177 38609 1211 38648
rect 1273 38682 1307 38721
rect 1273 38609 1307 38648
rect 1387 38652 1421 38685
rect 1387 38583 1421 38617
rect 199 38473 233 38549
rect 297 38537 313 38571
rect 347 38537 363 38571
rect 489 38537 505 38571
rect 539 38537 555 38571
rect 681 38537 697 38571
rect 731 38537 747 38571
rect 873 38537 889 38571
rect 923 38537 939 38571
rect 1065 38537 1081 38571
rect 1115 38537 1131 38571
rect 1257 38537 1273 38571
rect 1307 38537 1323 38571
rect 1387 38473 1421 38546
rect 199 38439 317 38473
rect 351 38439 385 38473
rect 419 38439 453 38473
rect 487 38439 521 38473
rect 555 38439 589 38473
rect 623 38439 657 38473
rect 691 38439 725 38473
rect 759 38439 793 38473
rect 827 38439 861 38473
rect 895 38439 929 38473
rect 963 38439 997 38473
rect 1031 38439 1065 38473
rect 1099 38439 1133 38473
rect 1167 38439 1201 38473
rect 1235 38439 1269 38473
rect 1303 38439 1421 38473
rect 2352 38799 2470 38833
rect 2504 38799 2538 38833
rect 2572 38799 2606 38833
rect 2640 38799 2674 38833
rect 2708 38799 2742 38833
rect 2776 38799 2810 38833
rect 2844 38799 2878 38833
rect 2912 38799 2946 38833
rect 2980 38799 3014 38833
rect 3048 38799 3082 38833
rect 3116 38799 3150 38833
rect 3184 38799 3218 38833
rect 3252 38799 3286 38833
rect 3320 38799 3354 38833
rect 3388 38799 3422 38833
rect 3456 38799 3574 38833
rect 2352 38723 2386 38799
rect 3540 38728 3574 38799
rect 3873 38799 3991 38833
rect 4025 38799 4059 38833
rect 4093 38799 4127 38833
rect 4161 38799 4195 38833
rect 4229 38799 4263 38833
rect 4297 38799 4331 38833
rect 4365 38799 4399 38833
rect 4433 38799 4467 38833
rect 4501 38799 4535 38833
rect 4569 38799 4603 38833
rect 4637 38799 4671 38833
rect 4705 38799 4739 38833
rect 4773 38799 4807 38833
rect 4841 38799 4875 38833
rect 4909 38799 4943 38833
rect 4977 38799 5095 38833
rect 3675 38763 3691 38797
rect 3725 38763 3741 38797
rect 2352 38655 2386 38689
rect 2352 38587 2386 38621
rect 2466 38686 2500 38725
rect 2466 38613 2500 38652
rect 2562 38686 2596 38725
rect 2562 38613 2596 38652
rect 2658 38686 2692 38725
rect 2658 38613 2692 38652
rect 2754 38686 2788 38725
rect 2754 38613 2788 38652
rect 2850 38686 2884 38725
rect 2850 38613 2884 38652
rect 2946 38686 2980 38725
rect 2946 38613 2980 38652
rect 3042 38686 3076 38725
rect 3042 38613 3076 38652
rect 3138 38686 3172 38725
rect 3138 38613 3172 38652
rect 3234 38686 3268 38725
rect 3234 38613 3268 38652
rect 3330 38686 3364 38725
rect 3330 38613 3364 38652
rect 3426 38686 3460 38725
rect 3426 38613 3460 38652
rect 3540 38656 3574 38689
rect 3647 38713 3681 38729
rect 3647 38621 3681 38637
rect 3735 38713 3769 38729
rect 3735 38621 3769 38637
rect 3873 38723 3907 38799
rect 5061 38728 5095 38799
rect 3873 38655 3907 38689
rect 3540 38587 3574 38621
rect 2352 38477 2386 38553
rect 2450 38541 2466 38575
rect 2500 38541 2516 38575
rect 2642 38541 2658 38575
rect 2692 38541 2708 38575
rect 2834 38541 2850 38575
rect 2884 38541 2900 38575
rect 3026 38541 3042 38575
rect 3076 38541 3092 38575
rect 3218 38541 3234 38575
rect 3268 38541 3284 38575
rect 3410 38541 3426 38575
rect 3460 38541 3476 38575
rect 3540 38477 3574 38550
rect 2352 38443 2470 38477
rect 2504 38443 2538 38477
rect 2572 38443 2606 38477
rect 2640 38443 2674 38477
rect 2708 38443 2742 38477
rect 2776 38443 2810 38477
rect 2844 38443 2878 38477
rect 2912 38443 2946 38477
rect 2980 38443 3014 38477
rect 3048 38443 3082 38477
rect 3116 38443 3150 38477
rect 3184 38443 3218 38477
rect 3252 38443 3286 38477
rect 3320 38443 3354 38477
rect 3388 38443 3422 38477
rect 3456 38443 3574 38477
rect 3873 38587 3907 38621
rect 3987 38686 4021 38725
rect 3987 38613 4021 38652
rect 4083 38686 4117 38725
rect 4083 38613 4117 38652
rect 4179 38686 4213 38725
rect 4179 38613 4213 38652
rect 4275 38686 4309 38725
rect 4275 38613 4309 38652
rect 4371 38686 4405 38725
rect 4371 38613 4405 38652
rect 4467 38686 4501 38725
rect 4467 38613 4501 38652
rect 4563 38686 4597 38725
rect 4563 38613 4597 38652
rect 4659 38686 4693 38725
rect 4659 38613 4693 38652
rect 4755 38686 4789 38725
rect 4755 38613 4789 38652
rect 4851 38686 4885 38725
rect 4851 38613 4885 38652
rect 4947 38686 4981 38725
rect 4947 38613 4981 38652
rect 5061 38656 5095 38689
rect 5340 38804 5348 38838
rect 5382 38804 5386 38838
rect 5420 38843 5486 38854
rect 5420 38840 5450 38843
rect 5420 38806 5436 38840
rect 5484 38809 5486 38843
rect 5470 38806 5486 38809
rect 5340 38768 5386 38804
rect 5340 38756 5406 38768
rect 5340 38722 5356 38756
rect 5390 38722 5406 38756
rect 5340 38688 5406 38722
rect 5340 38654 5356 38688
rect 5390 38654 5406 38688
rect 5340 38642 5406 38654
rect 5440 38756 5486 38772
rect 5474 38722 5486 38756
rect 5440 38688 5486 38722
rect 5474 38654 5486 38688
rect 5061 38587 5095 38621
rect 5440 38608 5486 38654
rect 3873 38477 3907 38553
rect 3971 38541 3987 38575
rect 4021 38541 4037 38575
rect 4163 38541 4179 38575
rect 4213 38541 4229 38575
rect 4355 38541 4371 38575
rect 4405 38541 4421 38575
rect 4547 38541 4563 38575
rect 4597 38541 4613 38575
rect 4739 38541 4755 38575
rect 4789 38541 4805 38575
rect 4931 38541 4947 38575
rect 4981 38541 4997 38575
rect 5274 38574 5303 38608
rect 5337 38574 5395 38608
rect 5429 38574 5487 38608
rect 5521 38574 5550 38608
rect 5061 38477 5095 38550
rect 3873 38443 3991 38477
rect 4025 38443 4059 38477
rect 4093 38443 4127 38477
rect 4161 38443 4195 38477
rect 4229 38443 4263 38477
rect 4297 38443 4331 38477
rect 4365 38443 4399 38477
rect 4433 38443 4467 38477
rect 4501 38443 4535 38477
rect 4569 38443 4603 38477
rect 4637 38443 4671 38477
rect 4705 38443 4739 38477
rect 4773 38443 4807 38477
rect 4841 38443 4875 38477
rect 4909 38443 4943 38477
rect 4977 38443 5095 38477
rect 199 38160 317 38194
rect 351 38160 385 38194
rect 419 38160 453 38194
rect 487 38160 521 38194
rect 555 38160 589 38194
rect 623 38160 657 38194
rect 691 38160 725 38194
rect 759 38160 793 38194
rect 827 38160 861 38194
rect 895 38160 929 38194
rect 963 38160 997 38194
rect 1031 38160 1065 38194
rect 1099 38160 1133 38194
rect 1167 38160 1201 38194
rect 1235 38160 1269 38194
rect 1303 38160 1421 38194
rect 199 38092 233 38160
rect 1387 38092 1421 38160
rect 297 38058 313 38092
rect 347 38058 363 38092
rect 489 38058 505 38092
rect 539 38058 555 38092
rect 681 38058 697 38092
rect 731 38058 747 38092
rect 873 38058 889 38092
rect 923 38058 939 38092
rect 1065 38058 1081 38092
rect 1115 38058 1131 38092
rect 1257 38058 1273 38092
rect 1307 38058 1323 38092
rect 199 38024 233 38058
rect 1387 38024 1421 38032
rect 199 37956 233 37990
rect 199 37888 233 37922
rect 199 37820 233 37854
rect 199 37752 233 37786
rect 313 37993 347 38014
rect 313 37925 347 37929
rect 313 37819 347 37823
rect 313 37734 347 37755
rect 409 37993 443 38014
rect 409 37925 443 37929
rect 409 37819 443 37823
rect 409 37734 443 37755
rect 505 37993 539 38014
rect 505 37925 539 37929
rect 505 37819 539 37823
rect 505 37734 539 37755
rect 601 37993 635 38014
rect 601 37925 635 37929
rect 601 37819 635 37823
rect 601 37734 635 37755
rect 697 37993 731 38014
rect 697 37925 731 37929
rect 697 37819 731 37823
rect 697 37734 731 37755
rect 793 37993 827 38014
rect 793 37925 827 37929
rect 793 37819 827 37823
rect 793 37734 827 37755
rect 889 37993 923 38014
rect 889 37925 923 37929
rect 889 37819 923 37823
rect 889 37734 923 37755
rect 985 37993 1019 38014
rect 985 37925 1019 37929
rect 985 37819 1019 37823
rect 985 37734 1019 37755
rect 1081 37993 1115 38014
rect 1081 37925 1115 37929
rect 1081 37819 1115 37823
rect 1081 37734 1115 37755
rect 1177 37993 1211 38014
rect 1177 37925 1211 37929
rect 1177 37819 1211 37823
rect 1177 37734 1211 37755
rect 1273 37993 1307 38014
rect 1273 37925 1307 37929
rect 1273 37819 1307 37823
rect 1273 37734 1307 37755
rect 1387 37956 1421 37960
rect 1387 37850 1421 37854
rect 1387 37778 1421 37786
rect 199 37650 233 37718
rect 1387 37650 1421 37718
rect 199 37616 317 37650
rect 351 37616 385 37650
rect 419 37616 453 37650
rect 487 37616 521 37650
rect 555 37616 589 37650
rect 623 37616 657 37650
rect 691 37616 725 37650
rect 759 37616 793 37650
rect 827 37616 861 37650
rect 895 37616 929 37650
rect 963 37616 997 37650
rect 1031 37616 1065 37650
rect 1099 37616 1133 37650
rect 1167 37616 1201 37650
rect 1235 37616 1269 37650
rect 1303 37616 1421 37650
rect 2352 38164 2470 38198
rect 2504 38164 2538 38198
rect 2572 38164 2606 38198
rect 2640 38164 2674 38198
rect 2708 38164 2742 38198
rect 2776 38164 2810 38198
rect 2844 38164 2878 38198
rect 2912 38164 2946 38198
rect 2980 38164 3014 38198
rect 3048 38164 3082 38198
rect 3116 38164 3150 38198
rect 3184 38164 3218 38198
rect 3252 38164 3286 38198
rect 3320 38164 3354 38198
rect 3388 38164 3422 38198
rect 3456 38164 3574 38198
rect 2352 38096 2386 38164
rect 3540 38096 3574 38164
rect 2450 38062 2466 38096
rect 2500 38062 2516 38096
rect 2642 38062 2658 38096
rect 2692 38062 2708 38096
rect 2834 38062 2850 38096
rect 2884 38062 2900 38096
rect 3026 38062 3042 38096
rect 3076 38062 3092 38096
rect 3218 38062 3234 38096
rect 3268 38062 3284 38096
rect 3410 38062 3426 38096
rect 3460 38062 3476 38096
rect 2352 38028 2386 38062
rect 3540 38028 3574 38036
rect 2352 37960 2386 37994
rect 2352 37892 2386 37926
rect 2352 37824 2386 37858
rect 2352 37756 2386 37790
rect 2466 37997 2500 38018
rect 2466 37929 2500 37933
rect 2466 37823 2500 37827
rect 2466 37738 2500 37759
rect 2562 37997 2596 38018
rect 2562 37929 2596 37933
rect 2562 37823 2596 37827
rect 2562 37738 2596 37759
rect 2658 37997 2692 38018
rect 2658 37929 2692 37933
rect 2658 37823 2692 37827
rect 2658 37738 2692 37759
rect 2754 37997 2788 38018
rect 2754 37929 2788 37933
rect 2754 37823 2788 37827
rect 2754 37738 2788 37759
rect 2850 37997 2884 38018
rect 2850 37929 2884 37933
rect 2850 37823 2884 37827
rect 2850 37738 2884 37759
rect 2946 37997 2980 38018
rect 2946 37929 2980 37933
rect 2946 37823 2980 37827
rect 2946 37738 2980 37759
rect 3042 37997 3076 38018
rect 3042 37929 3076 37933
rect 3042 37823 3076 37827
rect 3042 37738 3076 37759
rect 3138 37997 3172 38018
rect 3138 37929 3172 37933
rect 3138 37823 3172 37827
rect 3138 37738 3172 37759
rect 3234 37997 3268 38018
rect 3234 37929 3268 37933
rect 3234 37823 3268 37827
rect 3234 37738 3268 37759
rect 3330 37997 3364 38018
rect 3330 37929 3364 37933
rect 3330 37823 3364 37827
rect 3330 37738 3364 37759
rect 3426 37997 3460 38018
rect 3426 37929 3460 37933
rect 3426 37823 3460 37827
rect 3426 37738 3460 37759
rect 3540 37960 3574 37964
rect 3540 37854 3574 37858
rect 3540 37782 3574 37790
rect 2352 37654 2386 37722
rect 3540 37654 3574 37722
rect 2352 37620 2470 37654
rect 2504 37620 2538 37654
rect 2572 37620 2606 37654
rect 2640 37620 2674 37654
rect 2708 37620 2742 37654
rect 2776 37620 2810 37654
rect 2844 37620 2878 37654
rect 2912 37620 2946 37654
rect 2980 37620 3014 37654
rect 3048 37620 3082 37654
rect 3116 37620 3150 37654
rect 3184 37620 3218 37654
rect 3252 37620 3286 37654
rect 3320 37620 3354 37654
rect 3388 37620 3422 37654
rect 3456 37620 3574 37654
rect 3873 38164 3991 38198
rect 4025 38164 4059 38198
rect 4093 38164 4127 38198
rect 4161 38164 4195 38198
rect 4229 38164 4263 38198
rect 4297 38164 4331 38198
rect 4365 38164 4399 38198
rect 4433 38164 4467 38198
rect 4501 38164 4535 38198
rect 4569 38164 4603 38198
rect 4637 38164 4671 38198
rect 4705 38164 4739 38198
rect 4773 38164 4807 38198
rect 4841 38164 4875 38198
rect 4909 38164 4943 38198
rect 4977 38164 5095 38198
rect 3873 38096 3907 38164
rect 5061 38096 5095 38164
rect 3971 38062 3987 38096
rect 4021 38062 4037 38096
rect 4163 38062 4179 38096
rect 4213 38062 4229 38096
rect 4355 38062 4371 38096
rect 4405 38062 4421 38096
rect 4547 38062 4563 38096
rect 4597 38062 4613 38096
rect 4739 38062 4755 38096
rect 4789 38062 4805 38096
rect 4931 38062 4947 38096
rect 4981 38062 4997 38096
rect 3873 38028 3907 38062
rect 5061 38028 5095 38036
rect 3873 37960 3907 37994
rect 3873 37892 3907 37926
rect 3873 37824 3907 37858
rect 3873 37756 3907 37790
rect 3987 37997 4021 38018
rect 3987 37929 4021 37933
rect 3987 37823 4021 37827
rect 3987 37738 4021 37759
rect 4083 37997 4117 38018
rect 4083 37929 4117 37933
rect 4083 37823 4117 37827
rect 4083 37738 4117 37759
rect 4179 37997 4213 38018
rect 4179 37929 4213 37933
rect 4179 37823 4213 37827
rect 4179 37738 4213 37759
rect 4275 37997 4309 38018
rect 4275 37929 4309 37933
rect 4275 37823 4309 37827
rect 4275 37738 4309 37759
rect 4371 37997 4405 38018
rect 4371 37929 4405 37933
rect 4371 37823 4405 37827
rect 4371 37738 4405 37759
rect 4467 37997 4501 38018
rect 4467 37929 4501 37933
rect 4467 37823 4501 37827
rect 4467 37738 4501 37759
rect 4563 37997 4597 38018
rect 4563 37929 4597 37933
rect 4563 37823 4597 37827
rect 4563 37738 4597 37759
rect 4659 37997 4693 38018
rect 4659 37929 4693 37933
rect 4659 37823 4693 37827
rect 4659 37738 4693 37759
rect 4755 37997 4789 38018
rect 4755 37929 4789 37933
rect 4755 37823 4789 37827
rect 4755 37738 4789 37759
rect 4851 37997 4885 38018
rect 4851 37929 4885 37933
rect 4851 37823 4885 37827
rect 4851 37738 4885 37759
rect 4947 37997 4981 38018
rect 4947 37929 4981 37933
rect 4947 37823 4981 37827
rect 4947 37738 4981 37759
rect 5061 37960 5095 37964
rect 5061 37854 5095 37858
rect 5274 37831 5303 37865
rect 5337 37831 5395 37865
rect 5429 37831 5487 37865
rect 5521 37831 5550 37865
rect 5061 37782 5095 37790
rect 3873 37654 3907 37722
rect 5061 37654 5095 37722
rect 3873 37620 3991 37654
rect 4025 37620 4059 37654
rect 4093 37620 4127 37654
rect 4161 37620 4195 37654
rect 4229 37620 4263 37654
rect 4297 37620 4331 37654
rect 4365 37620 4399 37654
rect 4433 37620 4467 37654
rect 4501 37620 4535 37654
rect 4569 37620 4603 37654
rect 4637 37620 4671 37654
rect 4705 37620 4739 37654
rect 4773 37620 4807 37654
rect 4841 37620 4875 37654
rect 4909 37620 4943 37654
rect 4977 37620 5095 37654
rect 5340 37789 5406 37797
rect 5340 37755 5356 37789
rect 5390 37755 5406 37789
rect 5340 37721 5406 37755
rect 5340 37687 5356 37721
rect 5390 37687 5406 37721
rect 5340 37653 5406 37687
rect 5340 37619 5356 37653
rect 5390 37619 5406 37653
rect 5340 37601 5406 37619
rect 5440 37789 5482 37831
rect 5474 37755 5482 37789
rect 5440 37721 5482 37755
rect 5474 37687 5482 37721
rect 5440 37653 5482 37687
rect 5474 37619 5482 37653
rect 5440 37603 5482 37619
rect 5340 37551 5386 37601
rect 199 37508 317 37542
rect 351 37508 385 37542
rect 419 37508 453 37542
rect 487 37508 521 37542
rect 555 37508 589 37542
rect 623 37508 657 37542
rect 691 37508 725 37542
rect 759 37508 793 37542
rect 827 37508 861 37542
rect 895 37508 929 37542
rect 963 37508 997 37542
rect 1031 37508 1065 37542
rect 1099 37508 1133 37542
rect 1167 37508 1201 37542
rect 1235 37508 1269 37542
rect 1303 37508 1421 37542
rect 199 37432 233 37508
rect 1387 37437 1421 37508
rect 199 37364 233 37398
rect 199 37296 233 37330
rect 313 37395 347 37434
rect 313 37322 347 37361
rect 409 37395 443 37434
rect 409 37322 443 37361
rect 505 37395 539 37434
rect 505 37322 539 37361
rect 601 37395 635 37434
rect 601 37322 635 37361
rect 697 37395 731 37434
rect 697 37322 731 37361
rect 793 37395 827 37434
rect 793 37322 827 37361
rect 889 37395 923 37434
rect 889 37322 923 37361
rect 985 37395 1019 37434
rect 985 37322 1019 37361
rect 1081 37395 1115 37434
rect 1081 37322 1115 37361
rect 1177 37395 1211 37434
rect 1177 37322 1211 37361
rect 1273 37395 1307 37434
rect 1273 37322 1307 37361
rect 1387 37365 1421 37398
rect 1387 37296 1421 37330
rect 199 37186 233 37262
rect 297 37250 313 37284
rect 347 37250 363 37284
rect 489 37250 505 37284
rect 539 37250 555 37284
rect 681 37250 697 37284
rect 731 37250 747 37284
rect 873 37250 889 37284
rect 923 37250 939 37284
rect 1065 37250 1081 37284
rect 1115 37250 1131 37284
rect 1257 37250 1273 37284
rect 1307 37250 1323 37284
rect 1387 37186 1421 37259
rect 199 37152 317 37186
rect 351 37152 385 37186
rect 419 37152 453 37186
rect 487 37152 521 37186
rect 555 37152 589 37186
rect 623 37152 657 37186
rect 691 37152 725 37186
rect 759 37152 793 37186
rect 827 37152 861 37186
rect 895 37152 929 37186
rect 963 37152 997 37186
rect 1031 37152 1065 37186
rect 1099 37152 1133 37186
rect 1167 37152 1201 37186
rect 1235 37152 1269 37186
rect 1303 37152 1421 37186
rect 2352 37512 2470 37546
rect 2504 37512 2538 37546
rect 2572 37512 2606 37546
rect 2640 37512 2674 37546
rect 2708 37512 2742 37546
rect 2776 37512 2810 37546
rect 2844 37512 2878 37546
rect 2912 37512 2946 37546
rect 2980 37512 3014 37546
rect 3048 37512 3082 37546
rect 3116 37512 3150 37546
rect 3184 37512 3218 37546
rect 3252 37512 3286 37546
rect 3320 37512 3354 37546
rect 3388 37512 3422 37546
rect 3456 37512 3574 37546
rect 2352 37436 2386 37512
rect 3540 37441 3574 37512
rect 3873 37512 3991 37546
rect 4025 37512 4059 37546
rect 4093 37512 4127 37546
rect 4161 37512 4195 37546
rect 4229 37512 4263 37546
rect 4297 37512 4331 37546
rect 4365 37512 4399 37546
rect 4433 37512 4467 37546
rect 4501 37512 4535 37546
rect 4569 37512 4603 37546
rect 4637 37512 4671 37546
rect 4705 37512 4739 37546
rect 4773 37512 4807 37546
rect 4841 37512 4875 37546
rect 4909 37512 4943 37546
rect 4977 37512 5095 37546
rect 3675 37476 3691 37510
rect 3725 37476 3741 37510
rect 2352 37368 2386 37402
rect 2352 37300 2386 37334
rect 2466 37399 2500 37438
rect 2466 37326 2500 37365
rect 2562 37399 2596 37438
rect 2562 37326 2596 37365
rect 2658 37399 2692 37438
rect 2658 37326 2692 37365
rect 2754 37399 2788 37438
rect 2754 37326 2788 37365
rect 2850 37399 2884 37438
rect 2850 37326 2884 37365
rect 2946 37399 2980 37438
rect 2946 37326 2980 37365
rect 3042 37399 3076 37438
rect 3042 37326 3076 37365
rect 3138 37399 3172 37438
rect 3138 37326 3172 37365
rect 3234 37399 3268 37438
rect 3234 37326 3268 37365
rect 3330 37399 3364 37438
rect 3330 37326 3364 37365
rect 3426 37399 3460 37438
rect 3426 37326 3460 37365
rect 3540 37369 3574 37402
rect 3647 37426 3681 37442
rect 3647 37334 3681 37350
rect 3735 37426 3769 37442
rect 3735 37334 3769 37350
rect 3873 37436 3907 37512
rect 5061 37441 5095 37512
rect 3873 37368 3907 37402
rect 3540 37300 3574 37334
rect 2352 37190 2386 37266
rect 2450 37254 2466 37288
rect 2500 37254 2516 37288
rect 2642 37254 2658 37288
rect 2692 37254 2708 37288
rect 2834 37254 2850 37288
rect 2884 37254 2900 37288
rect 3026 37254 3042 37288
rect 3076 37254 3092 37288
rect 3218 37254 3234 37288
rect 3268 37254 3284 37288
rect 3410 37254 3426 37288
rect 3460 37254 3476 37288
rect 3540 37190 3574 37263
rect 2352 37156 2470 37190
rect 2504 37156 2538 37190
rect 2572 37156 2606 37190
rect 2640 37156 2674 37190
rect 2708 37156 2742 37190
rect 2776 37156 2810 37190
rect 2844 37156 2878 37190
rect 2912 37156 2946 37190
rect 2980 37156 3014 37190
rect 3048 37156 3082 37190
rect 3116 37156 3150 37190
rect 3184 37156 3218 37190
rect 3252 37156 3286 37190
rect 3320 37156 3354 37190
rect 3388 37156 3422 37190
rect 3456 37156 3574 37190
rect 3873 37300 3907 37334
rect 3987 37399 4021 37438
rect 3987 37326 4021 37365
rect 4083 37399 4117 37438
rect 4083 37326 4117 37365
rect 4179 37399 4213 37438
rect 4179 37326 4213 37365
rect 4275 37399 4309 37438
rect 4275 37326 4309 37365
rect 4371 37399 4405 37438
rect 4371 37326 4405 37365
rect 4467 37399 4501 37438
rect 4467 37326 4501 37365
rect 4563 37399 4597 37438
rect 4563 37326 4597 37365
rect 4659 37399 4693 37438
rect 4659 37326 4693 37365
rect 4755 37399 4789 37438
rect 4755 37326 4789 37365
rect 4851 37399 4885 37438
rect 4851 37326 4885 37365
rect 4947 37399 4981 37438
rect 4947 37326 4981 37365
rect 5061 37369 5095 37402
rect 5340 37517 5348 37551
rect 5382 37517 5386 37551
rect 5420 37556 5486 37567
rect 5420 37553 5450 37556
rect 5420 37519 5436 37553
rect 5484 37522 5486 37556
rect 5470 37519 5486 37522
rect 5340 37481 5386 37517
rect 5340 37469 5406 37481
rect 5340 37435 5356 37469
rect 5390 37435 5406 37469
rect 5340 37401 5406 37435
rect 5340 37367 5356 37401
rect 5390 37367 5406 37401
rect 5340 37355 5406 37367
rect 5440 37469 5486 37485
rect 5474 37435 5486 37469
rect 5440 37401 5486 37435
rect 5474 37367 5486 37401
rect 5061 37300 5095 37334
rect 5440 37321 5486 37367
rect 3873 37190 3907 37266
rect 3971 37254 3987 37288
rect 4021 37254 4037 37288
rect 4163 37254 4179 37288
rect 4213 37254 4229 37288
rect 4355 37254 4371 37288
rect 4405 37254 4421 37288
rect 4547 37254 4563 37288
rect 4597 37254 4613 37288
rect 4739 37254 4755 37288
rect 4789 37254 4805 37288
rect 4931 37254 4947 37288
rect 4981 37254 4997 37288
rect 5274 37287 5303 37321
rect 5337 37287 5395 37321
rect 5429 37287 5487 37321
rect 5521 37287 5550 37321
rect 5061 37190 5095 37263
rect 3873 37156 3991 37190
rect 4025 37156 4059 37190
rect 4093 37156 4127 37190
rect 4161 37156 4195 37190
rect 4229 37156 4263 37190
rect 4297 37156 4331 37190
rect 4365 37156 4399 37190
rect 4433 37156 4467 37190
rect 4501 37156 4535 37190
rect 4569 37156 4603 37190
rect 4637 37156 4671 37190
rect 4705 37156 4739 37190
rect 4773 37156 4807 37190
rect 4841 37156 4875 37190
rect 4909 37156 4943 37190
rect 4977 37156 5095 37190
rect 199 36873 317 36907
rect 351 36873 385 36907
rect 419 36873 453 36907
rect 487 36873 521 36907
rect 555 36873 589 36907
rect 623 36873 657 36907
rect 691 36873 725 36907
rect 759 36873 793 36907
rect 827 36873 861 36907
rect 895 36873 929 36907
rect 963 36873 997 36907
rect 1031 36873 1065 36907
rect 1099 36873 1133 36907
rect 1167 36873 1201 36907
rect 1235 36873 1269 36907
rect 1303 36873 1421 36907
rect 199 36805 233 36873
rect 1387 36805 1421 36873
rect 297 36771 313 36805
rect 347 36771 363 36805
rect 489 36771 505 36805
rect 539 36771 555 36805
rect 681 36771 697 36805
rect 731 36771 747 36805
rect 873 36771 889 36805
rect 923 36771 939 36805
rect 1065 36771 1081 36805
rect 1115 36771 1131 36805
rect 1257 36771 1273 36805
rect 1307 36771 1323 36805
rect 199 36737 233 36771
rect 1387 36737 1421 36745
rect 199 36669 233 36703
rect 199 36601 233 36635
rect 199 36533 233 36567
rect 199 36465 233 36499
rect 313 36706 347 36727
rect 313 36638 347 36642
rect 313 36532 347 36536
rect 313 36447 347 36468
rect 409 36706 443 36727
rect 409 36638 443 36642
rect 409 36532 443 36536
rect 409 36447 443 36468
rect 505 36706 539 36727
rect 505 36638 539 36642
rect 505 36532 539 36536
rect 505 36447 539 36468
rect 601 36706 635 36727
rect 601 36638 635 36642
rect 601 36532 635 36536
rect 601 36447 635 36468
rect 697 36706 731 36727
rect 697 36638 731 36642
rect 697 36532 731 36536
rect 697 36447 731 36468
rect 793 36706 827 36727
rect 793 36638 827 36642
rect 793 36532 827 36536
rect 793 36447 827 36468
rect 889 36706 923 36727
rect 889 36638 923 36642
rect 889 36532 923 36536
rect 889 36447 923 36468
rect 985 36706 1019 36727
rect 985 36638 1019 36642
rect 985 36532 1019 36536
rect 985 36447 1019 36468
rect 1081 36706 1115 36727
rect 1081 36638 1115 36642
rect 1081 36532 1115 36536
rect 1081 36447 1115 36468
rect 1177 36706 1211 36727
rect 1177 36638 1211 36642
rect 1177 36532 1211 36536
rect 1177 36447 1211 36468
rect 1273 36706 1307 36727
rect 1273 36638 1307 36642
rect 1273 36532 1307 36536
rect 1273 36447 1307 36468
rect 1387 36669 1421 36673
rect 1387 36563 1421 36567
rect 1387 36491 1421 36499
rect 199 36363 233 36431
rect 1387 36363 1421 36431
rect 199 36329 317 36363
rect 351 36329 385 36363
rect 419 36329 453 36363
rect 487 36329 521 36363
rect 555 36329 589 36363
rect 623 36329 657 36363
rect 691 36329 725 36363
rect 759 36329 793 36363
rect 827 36329 861 36363
rect 895 36329 929 36363
rect 963 36329 997 36363
rect 1031 36329 1065 36363
rect 1099 36329 1133 36363
rect 1167 36329 1201 36363
rect 1235 36329 1269 36363
rect 1303 36329 1421 36363
rect 2352 36877 2470 36911
rect 2504 36877 2538 36911
rect 2572 36877 2606 36911
rect 2640 36877 2674 36911
rect 2708 36877 2742 36911
rect 2776 36877 2810 36911
rect 2844 36877 2878 36911
rect 2912 36877 2946 36911
rect 2980 36877 3014 36911
rect 3048 36877 3082 36911
rect 3116 36877 3150 36911
rect 3184 36877 3218 36911
rect 3252 36877 3286 36911
rect 3320 36877 3354 36911
rect 3388 36877 3422 36911
rect 3456 36877 3574 36911
rect 2352 36809 2386 36877
rect 3540 36809 3574 36877
rect 2450 36775 2466 36809
rect 2500 36775 2516 36809
rect 2642 36775 2658 36809
rect 2692 36775 2708 36809
rect 2834 36775 2850 36809
rect 2884 36775 2900 36809
rect 3026 36775 3042 36809
rect 3076 36775 3092 36809
rect 3218 36775 3234 36809
rect 3268 36775 3284 36809
rect 3410 36775 3426 36809
rect 3460 36775 3476 36809
rect 2352 36741 2386 36775
rect 3540 36741 3574 36749
rect 2352 36673 2386 36707
rect 2352 36605 2386 36639
rect 2352 36537 2386 36571
rect 2352 36469 2386 36503
rect 2466 36710 2500 36731
rect 2466 36642 2500 36646
rect 2466 36536 2500 36540
rect 2466 36451 2500 36472
rect 2562 36710 2596 36731
rect 2562 36642 2596 36646
rect 2562 36536 2596 36540
rect 2562 36451 2596 36472
rect 2658 36710 2692 36731
rect 2658 36642 2692 36646
rect 2658 36536 2692 36540
rect 2658 36451 2692 36472
rect 2754 36710 2788 36731
rect 2754 36642 2788 36646
rect 2754 36536 2788 36540
rect 2754 36451 2788 36472
rect 2850 36710 2884 36731
rect 2850 36642 2884 36646
rect 2850 36536 2884 36540
rect 2850 36451 2884 36472
rect 2946 36710 2980 36731
rect 2946 36642 2980 36646
rect 2946 36536 2980 36540
rect 2946 36451 2980 36472
rect 3042 36710 3076 36731
rect 3042 36642 3076 36646
rect 3042 36536 3076 36540
rect 3042 36451 3076 36472
rect 3138 36710 3172 36731
rect 3138 36642 3172 36646
rect 3138 36536 3172 36540
rect 3138 36451 3172 36472
rect 3234 36710 3268 36731
rect 3234 36642 3268 36646
rect 3234 36536 3268 36540
rect 3234 36451 3268 36472
rect 3330 36710 3364 36731
rect 3330 36642 3364 36646
rect 3330 36536 3364 36540
rect 3330 36451 3364 36472
rect 3426 36710 3460 36731
rect 3426 36642 3460 36646
rect 3426 36536 3460 36540
rect 3426 36451 3460 36472
rect 3540 36673 3574 36677
rect 3540 36567 3574 36571
rect 3540 36495 3574 36503
rect 2352 36367 2386 36435
rect 3540 36367 3574 36435
rect 2352 36333 2470 36367
rect 2504 36333 2538 36367
rect 2572 36333 2606 36367
rect 2640 36333 2674 36367
rect 2708 36333 2742 36367
rect 2776 36333 2810 36367
rect 2844 36333 2878 36367
rect 2912 36333 2946 36367
rect 2980 36333 3014 36367
rect 3048 36333 3082 36367
rect 3116 36333 3150 36367
rect 3184 36333 3218 36367
rect 3252 36333 3286 36367
rect 3320 36333 3354 36367
rect 3388 36333 3422 36367
rect 3456 36333 3574 36367
rect 3873 36877 3991 36911
rect 4025 36877 4059 36911
rect 4093 36877 4127 36911
rect 4161 36877 4195 36911
rect 4229 36877 4263 36911
rect 4297 36877 4331 36911
rect 4365 36877 4399 36911
rect 4433 36877 4467 36911
rect 4501 36877 4535 36911
rect 4569 36877 4603 36911
rect 4637 36877 4671 36911
rect 4705 36877 4739 36911
rect 4773 36877 4807 36911
rect 4841 36877 4875 36911
rect 4909 36877 4943 36911
rect 4977 36877 5095 36911
rect 3873 36809 3907 36877
rect 5061 36809 5095 36877
rect 3971 36775 3987 36809
rect 4021 36775 4037 36809
rect 4163 36775 4179 36809
rect 4213 36775 4229 36809
rect 4355 36775 4371 36809
rect 4405 36775 4421 36809
rect 4547 36775 4563 36809
rect 4597 36775 4613 36809
rect 4739 36775 4755 36809
rect 4789 36775 4805 36809
rect 4931 36775 4947 36809
rect 4981 36775 4997 36809
rect 3873 36741 3907 36775
rect 5061 36741 5095 36749
rect 3873 36673 3907 36707
rect 3873 36605 3907 36639
rect 3873 36537 3907 36571
rect 3873 36469 3907 36503
rect 3987 36710 4021 36731
rect 3987 36642 4021 36646
rect 3987 36536 4021 36540
rect 3987 36451 4021 36472
rect 4083 36710 4117 36731
rect 4083 36642 4117 36646
rect 4083 36536 4117 36540
rect 4083 36451 4117 36472
rect 4179 36710 4213 36731
rect 4179 36642 4213 36646
rect 4179 36536 4213 36540
rect 4179 36451 4213 36472
rect 4275 36710 4309 36731
rect 4275 36642 4309 36646
rect 4275 36536 4309 36540
rect 4275 36451 4309 36472
rect 4371 36710 4405 36731
rect 4371 36642 4405 36646
rect 4371 36536 4405 36540
rect 4371 36451 4405 36472
rect 4467 36710 4501 36731
rect 4467 36642 4501 36646
rect 4467 36536 4501 36540
rect 4467 36451 4501 36472
rect 4563 36710 4597 36731
rect 4563 36642 4597 36646
rect 4563 36536 4597 36540
rect 4563 36451 4597 36472
rect 4659 36710 4693 36731
rect 4659 36642 4693 36646
rect 4659 36536 4693 36540
rect 4659 36451 4693 36472
rect 4755 36710 4789 36731
rect 4755 36642 4789 36646
rect 4755 36536 4789 36540
rect 4755 36451 4789 36472
rect 4851 36710 4885 36731
rect 4851 36642 4885 36646
rect 4851 36536 4885 36540
rect 4851 36451 4885 36472
rect 4947 36710 4981 36731
rect 4947 36642 4981 36646
rect 4947 36536 4981 36540
rect 4947 36451 4981 36472
rect 5061 36673 5095 36677
rect 5061 36567 5095 36571
rect 5274 36544 5303 36578
rect 5337 36544 5395 36578
rect 5429 36544 5487 36578
rect 5521 36544 5550 36578
rect 5061 36495 5095 36503
rect 3873 36367 3907 36435
rect 5061 36367 5095 36435
rect 3873 36333 3991 36367
rect 4025 36333 4059 36367
rect 4093 36333 4127 36367
rect 4161 36333 4195 36367
rect 4229 36333 4263 36367
rect 4297 36333 4331 36367
rect 4365 36333 4399 36367
rect 4433 36333 4467 36367
rect 4501 36333 4535 36367
rect 4569 36333 4603 36367
rect 4637 36333 4671 36367
rect 4705 36333 4739 36367
rect 4773 36333 4807 36367
rect 4841 36333 4875 36367
rect 4909 36333 4943 36367
rect 4977 36333 5095 36367
rect 5340 36502 5406 36510
rect 5340 36468 5356 36502
rect 5390 36468 5406 36502
rect 5340 36434 5406 36468
rect 5340 36400 5356 36434
rect 5390 36400 5406 36434
rect 5340 36366 5406 36400
rect 5340 36332 5356 36366
rect 5390 36332 5406 36366
rect 5340 36314 5406 36332
rect 5440 36502 5482 36544
rect 5474 36468 5482 36502
rect 5440 36434 5482 36468
rect 5474 36400 5482 36434
rect 5440 36366 5482 36400
rect 5474 36332 5482 36366
rect 5440 36316 5482 36332
rect 5340 36264 5386 36314
rect 199 36221 317 36255
rect 351 36221 385 36255
rect 419 36221 453 36255
rect 487 36221 521 36255
rect 555 36221 589 36255
rect 623 36221 657 36255
rect 691 36221 725 36255
rect 759 36221 793 36255
rect 827 36221 861 36255
rect 895 36221 929 36255
rect 963 36221 997 36255
rect 1031 36221 1065 36255
rect 1099 36221 1133 36255
rect 1167 36221 1201 36255
rect 1235 36221 1269 36255
rect 1303 36221 1421 36255
rect 199 36145 233 36221
rect 1387 36150 1421 36221
rect 199 36077 233 36111
rect 199 36009 233 36043
rect 313 36108 347 36147
rect 313 36035 347 36074
rect 409 36108 443 36147
rect 409 36035 443 36074
rect 505 36108 539 36147
rect 505 36035 539 36074
rect 601 36108 635 36147
rect 601 36035 635 36074
rect 697 36108 731 36147
rect 697 36035 731 36074
rect 793 36108 827 36147
rect 793 36035 827 36074
rect 889 36108 923 36147
rect 889 36035 923 36074
rect 985 36108 1019 36147
rect 985 36035 1019 36074
rect 1081 36108 1115 36147
rect 1081 36035 1115 36074
rect 1177 36108 1211 36147
rect 1177 36035 1211 36074
rect 1273 36108 1307 36147
rect 1273 36035 1307 36074
rect 1387 36078 1421 36111
rect 1387 36009 1421 36043
rect 199 35899 233 35975
rect 297 35963 313 35997
rect 347 35963 363 35997
rect 489 35963 505 35997
rect 539 35963 555 35997
rect 681 35963 697 35997
rect 731 35963 747 35997
rect 873 35963 889 35997
rect 923 35963 939 35997
rect 1065 35963 1081 35997
rect 1115 35963 1131 35997
rect 1257 35963 1273 35997
rect 1307 35963 1323 35997
rect 1387 35899 1421 35972
rect 199 35865 317 35899
rect 351 35865 385 35899
rect 419 35865 453 35899
rect 487 35865 521 35899
rect 555 35865 589 35899
rect 623 35865 657 35899
rect 691 35865 725 35899
rect 759 35865 793 35899
rect 827 35865 861 35899
rect 895 35865 929 35899
rect 963 35865 997 35899
rect 1031 35865 1065 35899
rect 1099 35865 1133 35899
rect 1167 35865 1201 35899
rect 1235 35865 1269 35899
rect 1303 35865 1421 35899
rect 2352 36225 2470 36259
rect 2504 36225 2538 36259
rect 2572 36225 2606 36259
rect 2640 36225 2674 36259
rect 2708 36225 2742 36259
rect 2776 36225 2810 36259
rect 2844 36225 2878 36259
rect 2912 36225 2946 36259
rect 2980 36225 3014 36259
rect 3048 36225 3082 36259
rect 3116 36225 3150 36259
rect 3184 36225 3218 36259
rect 3252 36225 3286 36259
rect 3320 36225 3354 36259
rect 3388 36225 3422 36259
rect 3456 36225 3574 36259
rect 2352 36149 2386 36225
rect 3540 36154 3574 36225
rect 3873 36225 3991 36259
rect 4025 36225 4059 36259
rect 4093 36225 4127 36259
rect 4161 36225 4195 36259
rect 4229 36225 4263 36259
rect 4297 36225 4331 36259
rect 4365 36225 4399 36259
rect 4433 36225 4467 36259
rect 4501 36225 4535 36259
rect 4569 36225 4603 36259
rect 4637 36225 4671 36259
rect 4705 36225 4739 36259
rect 4773 36225 4807 36259
rect 4841 36225 4875 36259
rect 4909 36225 4943 36259
rect 4977 36225 5095 36259
rect 3675 36189 3691 36223
rect 3725 36189 3741 36223
rect 2352 36081 2386 36115
rect 2352 36013 2386 36047
rect 2466 36112 2500 36151
rect 2466 36039 2500 36078
rect 2562 36112 2596 36151
rect 2562 36039 2596 36078
rect 2658 36112 2692 36151
rect 2658 36039 2692 36078
rect 2754 36112 2788 36151
rect 2754 36039 2788 36078
rect 2850 36112 2884 36151
rect 2850 36039 2884 36078
rect 2946 36112 2980 36151
rect 2946 36039 2980 36078
rect 3042 36112 3076 36151
rect 3042 36039 3076 36078
rect 3138 36112 3172 36151
rect 3138 36039 3172 36078
rect 3234 36112 3268 36151
rect 3234 36039 3268 36078
rect 3330 36112 3364 36151
rect 3330 36039 3364 36078
rect 3426 36112 3460 36151
rect 3426 36039 3460 36078
rect 3540 36082 3574 36115
rect 3647 36139 3681 36155
rect 3647 36047 3681 36063
rect 3735 36139 3769 36155
rect 3735 36047 3769 36063
rect 3873 36149 3907 36225
rect 5061 36154 5095 36225
rect 3873 36081 3907 36115
rect 3540 36013 3574 36047
rect 2352 35903 2386 35979
rect 2450 35967 2466 36001
rect 2500 35967 2516 36001
rect 2642 35967 2658 36001
rect 2692 35967 2708 36001
rect 2834 35967 2850 36001
rect 2884 35967 2900 36001
rect 3026 35967 3042 36001
rect 3076 35967 3092 36001
rect 3218 35967 3234 36001
rect 3268 35967 3284 36001
rect 3410 35967 3426 36001
rect 3460 35967 3476 36001
rect 3540 35903 3574 35976
rect 2352 35869 2470 35903
rect 2504 35869 2538 35903
rect 2572 35869 2606 35903
rect 2640 35869 2674 35903
rect 2708 35869 2742 35903
rect 2776 35869 2810 35903
rect 2844 35869 2878 35903
rect 2912 35869 2946 35903
rect 2980 35869 3014 35903
rect 3048 35869 3082 35903
rect 3116 35869 3150 35903
rect 3184 35869 3218 35903
rect 3252 35869 3286 35903
rect 3320 35869 3354 35903
rect 3388 35869 3422 35903
rect 3456 35869 3574 35903
rect 3873 36013 3907 36047
rect 3987 36112 4021 36151
rect 3987 36039 4021 36078
rect 4083 36112 4117 36151
rect 4083 36039 4117 36078
rect 4179 36112 4213 36151
rect 4179 36039 4213 36078
rect 4275 36112 4309 36151
rect 4275 36039 4309 36078
rect 4371 36112 4405 36151
rect 4371 36039 4405 36078
rect 4467 36112 4501 36151
rect 4467 36039 4501 36078
rect 4563 36112 4597 36151
rect 4563 36039 4597 36078
rect 4659 36112 4693 36151
rect 4659 36039 4693 36078
rect 4755 36112 4789 36151
rect 4755 36039 4789 36078
rect 4851 36112 4885 36151
rect 4851 36039 4885 36078
rect 4947 36112 4981 36151
rect 4947 36039 4981 36078
rect 5061 36082 5095 36115
rect 5340 36230 5348 36264
rect 5382 36230 5386 36264
rect 5420 36269 5486 36280
rect 5420 36266 5450 36269
rect 5420 36232 5436 36266
rect 5484 36235 5486 36269
rect 5470 36232 5486 36235
rect 5340 36194 5386 36230
rect 5340 36182 5406 36194
rect 5340 36148 5356 36182
rect 5390 36148 5406 36182
rect 5340 36114 5406 36148
rect 5340 36080 5356 36114
rect 5390 36080 5406 36114
rect 5340 36068 5406 36080
rect 5440 36182 5486 36198
rect 5474 36148 5486 36182
rect 5440 36114 5486 36148
rect 5474 36080 5486 36114
rect 5061 36013 5095 36047
rect 5440 36034 5486 36080
rect 3873 35903 3907 35979
rect 3971 35967 3987 36001
rect 4021 35967 4037 36001
rect 4163 35967 4179 36001
rect 4213 35967 4229 36001
rect 4355 35967 4371 36001
rect 4405 35967 4421 36001
rect 4547 35967 4563 36001
rect 4597 35967 4613 36001
rect 4739 35967 4755 36001
rect 4789 35967 4805 36001
rect 4931 35967 4947 36001
rect 4981 35967 4997 36001
rect 5274 36000 5303 36034
rect 5337 36000 5395 36034
rect 5429 36000 5487 36034
rect 5521 36000 5550 36034
rect 5061 35903 5095 35976
rect 3873 35869 3991 35903
rect 4025 35869 4059 35903
rect 4093 35869 4127 35903
rect 4161 35869 4195 35903
rect 4229 35869 4263 35903
rect 4297 35869 4331 35903
rect 4365 35869 4399 35903
rect 4433 35869 4467 35903
rect 4501 35869 4535 35903
rect 4569 35869 4603 35903
rect 4637 35869 4671 35903
rect 4705 35869 4739 35903
rect 4773 35869 4807 35903
rect 4841 35869 4875 35903
rect 4909 35869 4943 35903
rect 4977 35869 5095 35903
rect 199 35586 317 35620
rect 351 35586 385 35620
rect 419 35586 453 35620
rect 487 35586 521 35620
rect 555 35586 589 35620
rect 623 35586 657 35620
rect 691 35586 725 35620
rect 759 35586 793 35620
rect 827 35586 861 35620
rect 895 35586 929 35620
rect 963 35586 997 35620
rect 1031 35586 1065 35620
rect 1099 35586 1133 35620
rect 1167 35586 1201 35620
rect 1235 35586 1269 35620
rect 1303 35586 1421 35620
rect 199 35518 233 35586
rect 1387 35518 1421 35586
rect 297 35484 313 35518
rect 347 35484 363 35518
rect 489 35484 505 35518
rect 539 35484 555 35518
rect 681 35484 697 35518
rect 731 35484 747 35518
rect 873 35484 889 35518
rect 923 35484 939 35518
rect 1065 35484 1081 35518
rect 1115 35484 1131 35518
rect 1257 35484 1273 35518
rect 1307 35484 1323 35518
rect 199 35450 233 35484
rect 1387 35450 1421 35458
rect 199 35382 233 35416
rect 199 35314 233 35348
rect 199 35246 233 35280
rect 199 35178 233 35212
rect 313 35419 347 35440
rect 313 35351 347 35355
rect 313 35245 347 35249
rect 313 35160 347 35181
rect 409 35419 443 35440
rect 409 35351 443 35355
rect 409 35245 443 35249
rect 409 35160 443 35181
rect 505 35419 539 35440
rect 505 35351 539 35355
rect 505 35245 539 35249
rect 505 35160 539 35181
rect 601 35419 635 35440
rect 601 35351 635 35355
rect 601 35245 635 35249
rect 601 35160 635 35181
rect 697 35419 731 35440
rect 697 35351 731 35355
rect 697 35245 731 35249
rect 697 35160 731 35181
rect 793 35419 827 35440
rect 793 35351 827 35355
rect 793 35245 827 35249
rect 793 35160 827 35181
rect 889 35419 923 35440
rect 889 35351 923 35355
rect 889 35245 923 35249
rect 889 35160 923 35181
rect 985 35419 1019 35440
rect 985 35351 1019 35355
rect 985 35245 1019 35249
rect 985 35160 1019 35181
rect 1081 35419 1115 35440
rect 1081 35351 1115 35355
rect 1081 35245 1115 35249
rect 1081 35160 1115 35181
rect 1177 35419 1211 35440
rect 1177 35351 1211 35355
rect 1177 35245 1211 35249
rect 1177 35160 1211 35181
rect 1273 35419 1307 35440
rect 1273 35351 1307 35355
rect 1273 35245 1307 35249
rect 1273 35160 1307 35181
rect 1387 35382 1421 35386
rect 1387 35276 1421 35280
rect 1387 35204 1421 35212
rect 199 35076 233 35144
rect 1387 35076 1421 35144
rect 199 35042 317 35076
rect 351 35042 385 35076
rect 419 35042 453 35076
rect 487 35042 521 35076
rect 555 35042 589 35076
rect 623 35042 657 35076
rect 691 35042 725 35076
rect 759 35042 793 35076
rect 827 35042 861 35076
rect 895 35042 929 35076
rect 963 35042 997 35076
rect 1031 35042 1065 35076
rect 1099 35042 1133 35076
rect 1167 35042 1201 35076
rect 1235 35042 1269 35076
rect 1303 35042 1421 35076
rect 2352 35590 2470 35624
rect 2504 35590 2538 35624
rect 2572 35590 2606 35624
rect 2640 35590 2674 35624
rect 2708 35590 2742 35624
rect 2776 35590 2810 35624
rect 2844 35590 2878 35624
rect 2912 35590 2946 35624
rect 2980 35590 3014 35624
rect 3048 35590 3082 35624
rect 3116 35590 3150 35624
rect 3184 35590 3218 35624
rect 3252 35590 3286 35624
rect 3320 35590 3354 35624
rect 3388 35590 3422 35624
rect 3456 35590 3574 35624
rect 2352 35522 2386 35590
rect 3540 35522 3574 35590
rect 2450 35488 2466 35522
rect 2500 35488 2516 35522
rect 2642 35488 2658 35522
rect 2692 35488 2708 35522
rect 2834 35488 2850 35522
rect 2884 35488 2900 35522
rect 3026 35488 3042 35522
rect 3076 35488 3092 35522
rect 3218 35488 3234 35522
rect 3268 35488 3284 35522
rect 3410 35488 3426 35522
rect 3460 35488 3476 35522
rect 2352 35454 2386 35488
rect 3540 35454 3574 35462
rect 2352 35386 2386 35420
rect 2352 35318 2386 35352
rect 2352 35250 2386 35284
rect 2352 35182 2386 35216
rect 2466 35423 2500 35444
rect 2466 35355 2500 35359
rect 2466 35249 2500 35253
rect 2466 35164 2500 35185
rect 2562 35423 2596 35444
rect 2562 35355 2596 35359
rect 2562 35249 2596 35253
rect 2562 35164 2596 35185
rect 2658 35423 2692 35444
rect 2658 35355 2692 35359
rect 2658 35249 2692 35253
rect 2658 35164 2692 35185
rect 2754 35423 2788 35444
rect 2754 35355 2788 35359
rect 2754 35249 2788 35253
rect 2754 35164 2788 35185
rect 2850 35423 2884 35444
rect 2850 35355 2884 35359
rect 2850 35249 2884 35253
rect 2850 35164 2884 35185
rect 2946 35423 2980 35444
rect 2946 35355 2980 35359
rect 2946 35249 2980 35253
rect 2946 35164 2980 35185
rect 3042 35423 3076 35444
rect 3042 35355 3076 35359
rect 3042 35249 3076 35253
rect 3042 35164 3076 35185
rect 3138 35423 3172 35444
rect 3138 35355 3172 35359
rect 3138 35249 3172 35253
rect 3138 35164 3172 35185
rect 3234 35423 3268 35444
rect 3234 35355 3268 35359
rect 3234 35249 3268 35253
rect 3234 35164 3268 35185
rect 3330 35423 3364 35444
rect 3330 35355 3364 35359
rect 3330 35249 3364 35253
rect 3330 35164 3364 35185
rect 3426 35423 3460 35444
rect 3426 35355 3460 35359
rect 3426 35249 3460 35253
rect 3426 35164 3460 35185
rect 3540 35386 3574 35390
rect 3540 35280 3574 35284
rect 3540 35208 3574 35216
rect 2352 35080 2386 35148
rect 3540 35080 3574 35148
rect 2352 35046 2470 35080
rect 2504 35046 2538 35080
rect 2572 35046 2606 35080
rect 2640 35046 2674 35080
rect 2708 35046 2742 35080
rect 2776 35046 2810 35080
rect 2844 35046 2878 35080
rect 2912 35046 2946 35080
rect 2980 35046 3014 35080
rect 3048 35046 3082 35080
rect 3116 35046 3150 35080
rect 3184 35046 3218 35080
rect 3252 35046 3286 35080
rect 3320 35046 3354 35080
rect 3388 35046 3422 35080
rect 3456 35046 3574 35080
rect 3873 35590 3991 35624
rect 4025 35590 4059 35624
rect 4093 35590 4127 35624
rect 4161 35590 4195 35624
rect 4229 35590 4263 35624
rect 4297 35590 4331 35624
rect 4365 35590 4399 35624
rect 4433 35590 4467 35624
rect 4501 35590 4535 35624
rect 4569 35590 4603 35624
rect 4637 35590 4671 35624
rect 4705 35590 4739 35624
rect 4773 35590 4807 35624
rect 4841 35590 4875 35624
rect 4909 35590 4943 35624
rect 4977 35590 5095 35624
rect 3873 35522 3907 35590
rect 5061 35522 5095 35590
rect 3971 35488 3987 35522
rect 4021 35488 4037 35522
rect 4163 35488 4179 35522
rect 4213 35488 4229 35522
rect 4355 35488 4371 35522
rect 4405 35488 4421 35522
rect 4547 35488 4563 35522
rect 4597 35488 4613 35522
rect 4739 35488 4755 35522
rect 4789 35488 4805 35522
rect 4931 35488 4947 35522
rect 4981 35488 4997 35522
rect 3873 35454 3907 35488
rect 5061 35454 5095 35462
rect 3873 35386 3907 35420
rect 3873 35318 3907 35352
rect 3873 35250 3907 35284
rect 3873 35182 3907 35216
rect 3987 35423 4021 35444
rect 3987 35355 4021 35359
rect 3987 35249 4021 35253
rect 3987 35164 4021 35185
rect 4083 35423 4117 35444
rect 4083 35355 4117 35359
rect 4083 35249 4117 35253
rect 4083 35164 4117 35185
rect 4179 35423 4213 35444
rect 4179 35355 4213 35359
rect 4179 35249 4213 35253
rect 4179 35164 4213 35185
rect 4275 35423 4309 35444
rect 4275 35355 4309 35359
rect 4275 35249 4309 35253
rect 4275 35164 4309 35185
rect 4371 35423 4405 35444
rect 4371 35355 4405 35359
rect 4371 35249 4405 35253
rect 4371 35164 4405 35185
rect 4467 35423 4501 35444
rect 4467 35355 4501 35359
rect 4467 35249 4501 35253
rect 4467 35164 4501 35185
rect 4563 35423 4597 35444
rect 4563 35355 4597 35359
rect 4563 35249 4597 35253
rect 4563 35164 4597 35185
rect 4659 35423 4693 35444
rect 4659 35355 4693 35359
rect 4659 35249 4693 35253
rect 4659 35164 4693 35185
rect 4755 35423 4789 35444
rect 4755 35355 4789 35359
rect 4755 35249 4789 35253
rect 4755 35164 4789 35185
rect 4851 35423 4885 35444
rect 4851 35355 4885 35359
rect 4851 35249 4885 35253
rect 4851 35164 4885 35185
rect 4947 35423 4981 35444
rect 4947 35355 4981 35359
rect 4947 35249 4981 35253
rect 4947 35164 4981 35185
rect 5061 35386 5095 35390
rect 5061 35280 5095 35284
rect 5274 35257 5303 35291
rect 5337 35257 5395 35291
rect 5429 35257 5487 35291
rect 5521 35257 5550 35291
rect 5061 35208 5095 35216
rect 3873 35080 3907 35148
rect 5061 35080 5095 35148
rect 3873 35046 3991 35080
rect 4025 35046 4059 35080
rect 4093 35046 4127 35080
rect 4161 35046 4195 35080
rect 4229 35046 4263 35080
rect 4297 35046 4331 35080
rect 4365 35046 4399 35080
rect 4433 35046 4467 35080
rect 4501 35046 4535 35080
rect 4569 35046 4603 35080
rect 4637 35046 4671 35080
rect 4705 35046 4739 35080
rect 4773 35046 4807 35080
rect 4841 35046 4875 35080
rect 4909 35046 4943 35080
rect 4977 35046 5095 35080
rect 5340 35215 5406 35223
rect 5340 35181 5356 35215
rect 5390 35181 5406 35215
rect 5340 35147 5406 35181
rect 5340 35113 5356 35147
rect 5390 35113 5406 35147
rect 5340 35079 5406 35113
rect 5340 35045 5356 35079
rect 5390 35045 5406 35079
rect 5340 35027 5406 35045
rect 5440 35215 5482 35257
rect 5474 35181 5482 35215
rect 5440 35147 5482 35181
rect 5474 35113 5482 35147
rect 5440 35079 5482 35113
rect 5474 35045 5482 35079
rect 5440 35029 5482 35045
rect 5340 34977 5386 35027
rect 199 34934 317 34968
rect 351 34934 385 34968
rect 419 34934 453 34968
rect 487 34934 521 34968
rect 555 34934 589 34968
rect 623 34934 657 34968
rect 691 34934 725 34968
rect 759 34934 793 34968
rect 827 34934 861 34968
rect 895 34934 929 34968
rect 963 34934 997 34968
rect 1031 34934 1065 34968
rect 1099 34934 1133 34968
rect 1167 34934 1201 34968
rect 1235 34934 1269 34968
rect 1303 34934 1421 34968
rect 199 34858 233 34934
rect 1387 34863 1421 34934
rect 199 34790 233 34824
rect 199 34722 233 34756
rect 313 34821 347 34860
rect 313 34748 347 34787
rect 409 34821 443 34860
rect 409 34748 443 34787
rect 505 34821 539 34860
rect 505 34748 539 34787
rect 601 34821 635 34860
rect 601 34748 635 34787
rect 697 34821 731 34860
rect 697 34748 731 34787
rect 793 34821 827 34860
rect 793 34748 827 34787
rect 889 34821 923 34860
rect 889 34748 923 34787
rect 985 34821 1019 34860
rect 985 34748 1019 34787
rect 1081 34821 1115 34860
rect 1081 34748 1115 34787
rect 1177 34821 1211 34860
rect 1177 34748 1211 34787
rect 1273 34821 1307 34860
rect 1273 34748 1307 34787
rect 1387 34791 1421 34824
rect 1387 34722 1421 34756
rect 199 34612 233 34688
rect 297 34676 313 34710
rect 347 34676 363 34710
rect 489 34676 505 34710
rect 539 34676 555 34710
rect 681 34676 697 34710
rect 731 34676 747 34710
rect 873 34676 889 34710
rect 923 34676 939 34710
rect 1065 34676 1081 34710
rect 1115 34676 1131 34710
rect 1257 34676 1273 34710
rect 1307 34676 1323 34710
rect 1387 34612 1421 34685
rect 199 34578 317 34612
rect 351 34578 385 34612
rect 419 34578 453 34612
rect 487 34578 521 34612
rect 555 34578 589 34612
rect 623 34578 657 34612
rect 691 34578 725 34612
rect 759 34578 793 34612
rect 827 34578 861 34612
rect 895 34578 929 34612
rect 963 34578 997 34612
rect 1031 34578 1065 34612
rect 1099 34578 1133 34612
rect 1167 34578 1201 34612
rect 1235 34578 1269 34612
rect 1303 34578 1421 34612
rect 2352 34938 2470 34972
rect 2504 34938 2538 34972
rect 2572 34938 2606 34972
rect 2640 34938 2674 34972
rect 2708 34938 2742 34972
rect 2776 34938 2810 34972
rect 2844 34938 2878 34972
rect 2912 34938 2946 34972
rect 2980 34938 3014 34972
rect 3048 34938 3082 34972
rect 3116 34938 3150 34972
rect 3184 34938 3218 34972
rect 3252 34938 3286 34972
rect 3320 34938 3354 34972
rect 3388 34938 3422 34972
rect 3456 34938 3574 34972
rect 2352 34862 2386 34938
rect 3540 34867 3574 34938
rect 3873 34938 3991 34972
rect 4025 34938 4059 34972
rect 4093 34938 4127 34972
rect 4161 34938 4195 34972
rect 4229 34938 4263 34972
rect 4297 34938 4331 34972
rect 4365 34938 4399 34972
rect 4433 34938 4467 34972
rect 4501 34938 4535 34972
rect 4569 34938 4603 34972
rect 4637 34938 4671 34972
rect 4705 34938 4739 34972
rect 4773 34938 4807 34972
rect 4841 34938 4875 34972
rect 4909 34938 4943 34972
rect 4977 34938 5095 34972
rect 3675 34902 3691 34936
rect 3725 34902 3741 34936
rect 2352 34794 2386 34828
rect 2352 34726 2386 34760
rect 2466 34825 2500 34864
rect 2466 34752 2500 34791
rect 2562 34825 2596 34864
rect 2562 34752 2596 34791
rect 2658 34825 2692 34864
rect 2658 34752 2692 34791
rect 2754 34825 2788 34864
rect 2754 34752 2788 34791
rect 2850 34825 2884 34864
rect 2850 34752 2884 34791
rect 2946 34825 2980 34864
rect 2946 34752 2980 34791
rect 3042 34825 3076 34864
rect 3042 34752 3076 34791
rect 3138 34825 3172 34864
rect 3138 34752 3172 34791
rect 3234 34825 3268 34864
rect 3234 34752 3268 34791
rect 3330 34825 3364 34864
rect 3330 34752 3364 34791
rect 3426 34825 3460 34864
rect 3426 34752 3460 34791
rect 3540 34795 3574 34828
rect 3647 34852 3681 34868
rect 3647 34760 3681 34776
rect 3735 34852 3769 34868
rect 3735 34760 3769 34776
rect 3873 34862 3907 34938
rect 5061 34867 5095 34938
rect 3873 34794 3907 34828
rect 3540 34726 3574 34760
rect 2352 34616 2386 34692
rect 2450 34680 2466 34714
rect 2500 34680 2516 34714
rect 2642 34680 2658 34714
rect 2692 34680 2708 34714
rect 2834 34680 2850 34714
rect 2884 34680 2900 34714
rect 3026 34680 3042 34714
rect 3076 34680 3092 34714
rect 3218 34680 3234 34714
rect 3268 34680 3284 34714
rect 3410 34680 3426 34714
rect 3460 34680 3476 34714
rect 3540 34616 3574 34689
rect 2352 34582 2470 34616
rect 2504 34582 2538 34616
rect 2572 34582 2606 34616
rect 2640 34582 2674 34616
rect 2708 34582 2742 34616
rect 2776 34582 2810 34616
rect 2844 34582 2878 34616
rect 2912 34582 2946 34616
rect 2980 34582 3014 34616
rect 3048 34582 3082 34616
rect 3116 34582 3150 34616
rect 3184 34582 3218 34616
rect 3252 34582 3286 34616
rect 3320 34582 3354 34616
rect 3388 34582 3422 34616
rect 3456 34582 3574 34616
rect 3873 34726 3907 34760
rect 3987 34825 4021 34864
rect 3987 34752 4021 34791
rect 4083 34825 4117 34864
rect 4083 34752 4117 34791
rect 4179 34825 4213 34864
rect 4179 34752 4213 34791
rect 4275 34825 4309 34864
rect 4275 34752 4309 34791
rect 4371 34825 4405 34864
rect 4371 34752 4405 34791
rect 4467 34825 4501 34864
rect 4467 34752 4501 34791
rect 4563 34825 4597 34864
rect 4563 34752 4597 34791
rect 4659 34825 4693 34864
rect 4659 34752 4693 34791
rect 4755 34825 4789 34864
rect 4755 34752 4789 34791
rect 4851 34825 4885 34864
rect 4851 34752 4885 34791
rect 4947 34825 4981 34864
rect 4947 34752 4981 34791
rect 5061 34795 5095 34828
rect 5340 34943 5348 34977
rect 5382 34943 5386 34977
rect 5420 34982 5486 34993
rect 5420 34979 5450 34982
rect 5420 34945 5436 34979
rect 5484 34948 5486 34982
rect 5470 34945 5486 34948
rect 5340 34907 5386 34943
rect 5340 34895 5406 34907
rect 5340 34861 5356 34895
rect 5390 34861 5406 34895
rect 5340 34827 5406 34861
rect 5340 34793 5356 34827
rect 5390 34793 5406 34827
rect 5340 34781 5406 34793
rect 5440 34895 5486 34911
rect 5474 34861 5486 34895
rect 5440 34827 5486 34861
rect 5474 34793 5486 34827
rect 5061 34726 5095 34760
rect 5440 34747 5486 34793
rect 3873 34616 3907 34692
rect 3971 34680 3987 34714
rect 4021 34680 4037 34714
rect 4163 34680 4179 34714
rect 4213 34680 4229 34714
rect 4355 34680 4371 34714
rect 4405 34680 4421 34714
rect 4547 34680 4563 34714
rect 4597 34680 4613 34714
rect 4739 34680 4755 34714
rect 4789 34680 4805 34714
rect 4931 34680 4947 34714
rect 4981 34680 4997 34714
rect 5274 34713 5303 34747
rect 5337 34713 5395 34747
rect 5429 34713 5487 34747
rect 5521 34713 5550 34747
rect 5061 34616 5095 34689
rect 3873 34582 3991 34616
rect 4025 34582 4059 34616
rect 4093 34582 4127 34616
rect 4161 34582 4195 34616
rect 4229 34582 4263 34616
rect 4297 34582 4331 34616
rect 4365 34582 4399 34616
rect 4433 34582 4467 34616
rect 4501 34582 4535 34616
rect 4569 34582 4603 34616
rect 4637 34582 4671 34616
rect 4705 34582 4739 34616
rect 4773 34582 4807 34616
rect 4841 34582 4875 34616
rect 4909 34582 4943 34616
rect 4977 34582 5095 34616
rect 199 34299 317 34333
rect 351 34299 385 34333
rect 419 34299 453 34333
rect 487 34299 521 34333
rect 555 34299 589 34333
rect 623 34299 657 34333
rect 691 34299 725 34333
rect 759 34299 793 34333
rect 827 34299 861 34333
rect 895 34299 929 34333
rect 963 34299 997 34333
rect 1031 34299 1065 34333
rect 1099 34299 1133 34333
rect 1167 34299 1201 34333
rect 1235 34299 1269 34333
rect 1303 34299 1421 34333
rect 199 34231 233 34299
rect 1387 34231 1421 34299
rect 297 34197 313 34231
rect 347 34197 363 34231
rect 489 34197 505 34231
rect 539 34197 555 34231
rect 681 34197 697 34231
rect 731 34197 747 34231
rect 873 34197 889 34231
rect 923 34197 939 34231
rect 1065 34197 1081 34231
rect 1115 34197 1131 34231
rect 1257 34197 1273 34231
rect 1307 34197 1323 34231
rect 199 34163 233 34197
rect 1387 34163 1421 34171
rect 199 34095 233 34129
rect 199 34027 233 34061
rect 199 33959 233 33993
rect 199 33891 233 33925
rect 313 34132 347 34153
rect 313 34064 347 34068
rect 313 33958 347 33962
rect 313 33873 347 33894
rect 409 34132 443 34153
rect 409 34064 443 34068
rect 409 33958 443 33962
rect 409 33873 443 33894
rect 505 34132 539 34153
rect 505 34064 539 34068
rect 505 33958 539 33962
rect 505 33873 539 33894
rect 601 34132 635 34153
rect 601 34064 635 34068
rect 601 33958 635 33962
rect 601 33873 635 33894
rect 697 34132 731 34153
rect 697 34064 731 34068
rect 697 33958 731 33962
rect 697 33873 731 33894
rect 793 34132 827 34153
rect 793 34064 827 34068
rect 793 33958 827 33962
rect 793 33873 827 33894
rect 889 34132 923 34153
rect 889 34064 923 34068
rect 889 33958 923 33962
rect 889 33873 923 33894
rect 985 34132 1019 34153
rect 985 34064 1019 34068
rect 985 33958 1019 33962
rect 985 33873 1019 33894
rect 1081 34132 1115 34153
rect 1081 34064 1115 34068
rect 1081 33958 1115 33962
rect 1081 33873 1115 33894
rect 1177 34132 1211 34153
rect 1177 34064 1211 34068
rect 1177 33958 1211 33962
rect 1177 33873 1211 33894
rect 1273 34132 1307 34153
rect 1273 34064 1307 34068
rect 1273 33958 1307 33962
rect 1273 33873 1307 33894
rect 1387 34095 1421 34099
rect 1387 33989 1421 33993
rect 1387 33917 1421 33925
rect 199 33789 233 33857
rect 1387 33789 1421 33857
rect 199 33755 317 33789
rect 351 33755 385 33789
rect 419 33755 453 33789
rect 487 33755 521 33789
rect 555 33755 589 33789
rect 623 33755 657 33789
rect 691 33755 725 33789
rect 759 33755 793 33789
rect 827 33755 861 33789
rect 895 33755 929 33789
rect 963 33755 997 33789
rect 1031 33755 1065 33789
rect 1099 33755 1133 33789
rect 1167 33755 1201 33789
rect 1235 33755 1269 33789
rect 1303 33755 1421 33789
rect 2352 34303 2470 34337
rect 2504 34303 2538 34337
rect 2572 34303 2606 34337
rect 2640 34303 2674 34337
rect 2708 34303 2742 34337
rect 2776 34303 2810 34337
rect 2844 34303 2878 34337
rect 2912 34303 2946 34337
rect 2980 34303 3014 34337
rect 3048 34303 3082 34337
rect 3116 34303 3150 34337
rect 3184 34303 3218 34337
rect 3252 34303 3286 34337
rect 3320 34303 3354 34337
rect 3388 34303 3422 34337
rect 3456 34303 3574 34337
rect 2352 34235 2386 34303
rect 3540 34235 3574 34303
rect 2450 34201 2466 34235
rect 2500 34201 2516 34235
rect 2642 34201 2658 34235
rect 2692 34201 2708 34235
rect 2834 34201 2850 34235
rect 2884 34201 2900 34235
rect 3026 34201 3042 34235
rect 3076 34201 3092 34235
rect 3218 34201 3234 34235
rect 3268 34201 3284 34235
rect 3410 34201 3426 34235
rect 3460 34201 3476 34235
rect 2352 34167 2386 34201
rect 3540 34167 3574 34175
rect 2352 34099 2386 34133
rect 2352 34031 2386 34065
rect 2352 33963 2386 33997
rect 2352 33895 2386 33929
rect 2466 34136 2500 34157
rect 2466 34068 2500 34072
rect 2466 33962 2500 33966
rect 2466 33877 2500 33898
rect 2562 34136 2596 34157
rect 2562 34068 2596 34072
rect 2562 33962 2596 33966
rect 2562 33877 2596 33898
rect 2658 34136 2692 34157
rect 2658 34068 2692 34072
rect 2658 33962 2692 33966
rect 2658 33877 2692 33898
rect 2754 34136 2788 34157
rect 2754 34068 2788 34072
rect 2754 33962 2788 33966
rect 2754 33877 2788 33898
rect 2850 34136 2884 34157
rect 2850 34068 2884 34072
rect 2850 33962 2884 33966
rect 2850 33877 2884 33898
rect 2946 34136 2980 34157
rect 2946 34068 2980 34072
rect 2946 33962 2980 33966
rect 2946 33877 2980 33898
rect 3042 34136 3076 34157
rect 3042 34068 3076 34072
rect 3042 33962 3076 33966
rect 3042 33877 3076 33898
rect 3138 34136 3172 34157
rect 3138 34068 3172 34072
rect 3138 33962 3172 33966
rect 3138 33877 3172 33898
rect 3234 34136 3268 34157
rect 3234 34068 3268 34072
rect 3234 33962 3268 33966
rect 3234 33877 3268 33898
rect 3330 34136 3364 34157
rect 3330 34068 3364 34072
rect 3330 33962 3364 33966
rect 3330 33877 3364 33898
rect 3426 34136 3460 34157
rect 3426 34068 3460 34072
rect 3426 33962 3460 33966
rect 3426 33877 3460 33898
rect 3540 34099 3574 34103
rect 3540 33993 3574 33997
rect 3540 33921 3574 33929
rect 2352 33793 2386 33861
rect 3540 33793 3574 33861
rect 2352 33759 2470 33793
rect 2504 33759 2538 33793
rect 2572 33759 2606 33793
rect 2640 33759 2674 33793
rect 2708 33759 2742 33793
rect 2776 33759 2810 33793
rect 2844 33759 2878 33793
rect 2912 33759 2946 33793
rect 2980 33759 3014 33793
rect 3048 33759 3082 33793
rect 3116 33759 3150 33793
rect 3184 33759 3218 33793
rect 3252 33759 3286 33793
rect 3320 33759 3354 33793
rect 3388 33759 3422 33793
rect 3456 33759 3574 33793
rect 3873 34303 3991 34337
rect 4025 34303 4059 34337
rect 4093 34303 4127 34337
rect 4161 34303 4195 34337
rect 4229 34303 4263 34337
rect 4297 34303 4331 34337
rect 4365 34303 4399 34337
rect 4433 34303 4467 34337
rect 4501 34303 4535 34337
rect 4569 34303 4603 34337
rect 4637 34303 4671 34337
rect 4705 34303 4739 34337
rect 4773 34303 4807 34337
rect 4841 34303 4875 34337
rect 4909 34303 4943 34337
rect 4977 34303 5095 34337
rect 3873 34235 3907 34303
rect 5061 34235 5095 34303
rect 3971 34201 3987 34235
rect 4021 34201 4037 34235
rect 4163 34201 4179 34235
rect 4213 34201 4229 34235
rect 4355 34201 4371 34235
rect 4405 34201 4421 34235
rect 4547 34201 4563 34235
rect 4597 34201 4613 34235
rect 4739 34201 4755 34235
rect 4789 34201 4805 34235
rect 4931 34201 4947 34235
rect 4981 34201 4997 34235
rect 3873 34167 3907 34201
rect 5061 34167 5095 34175
rect 3873 34099 3907 34133
rect 3873 34031 3907 34065
rect 3873 33963 3907 33997
rect 3873 33895 3907 33929
rect 3987 34136 4021 34157
rect 3987 34068 4021 34072
rect 3987 33962 4021 33966
rect 3987 33877 4021 33898
rect 4083 34136 4117 34157
rect 4083 34068 4117 34072
rect 4083 33962 4117 33966
rect 4083 33877 4117 33898
rect 4179 34136 4213 34157
rect 4179 34068 4213 34072
rect 4179 33962 4213 33966
rect 4179 33877 4213 33898
rect 4275 34136 4309 34157
rect 4275 34068 4309 34072
rect 4275 33962 4309 33966
rect 4275 33877 4309 33898
rect 4371 34136 4405 34157
rect 4371 34068 4405 34072
rect 4371 33962 4405 33966
rect 4371 33877 4405 33898
rect 4467 34136 4501 34157
rect 4467 34068 4501 34072
rect 4467 33962 4501 33966
rect 4467 33877 4501 33898
rect 4563 34136 4597 34157
rect 4563 34068 4597 34072
rect 4563 33962 4597 33966
rect 4563 33877 4597 33898
rect 4659 34136 4693 34157
rect 4659 34068 4693 34072
rect 4659 33962 4693 33966
rect 4659 33877 4693 33898
rect 4755 34136 4789 34157
rect 4755 34068 4789 34072
rect 4755 33962 4789 33966
rect 4755 33877 4789 33898
rect 4851 34136 4885 34157
rect 4851 34068 4885 34072
rect 4851 33962 4885 33966
rect 4851 33877 4885 33898
rect 4947 34136 4981 34157
rect 4947 34068 4981 34072
rect 4947 33962 4981 33966
rect 4947 33877 4981 33898
rect 5061 34099 5095 34103
rect 5061 33993 5095 33997
rect 5274 33970 5303 34004
rect 5337 33970 5395 34004
rect 5429 33970 5487 34004
rect 5521 33970 5550 34004
rect 5061 33921 5095 33929
rect 3873 33793 3907 33861
rect 5061 33793 5095 33861
rect 3873 33759 3991 33793
rect 4025 33759 4059 33793
rect 4093 33759 4127 33793
rect 4161 33759 4195 33793
rect 4229 33759 4263 33793
rect 4297 33759 4331 33793
rect 4365 33759 4399 33793
rect 4433 33759 4467 33793
rect 4501 33759 4535 33793
rect 4569 33759 4603 33793
rect 4637 33759 4671 33793
rect 4705 33759 4739 33793
rect 4773 33759 4807 33793
rect 4841 33759 4875 33793
rect 4909 33759 4943 33793
rect 4977 33759 5095 33793
rect 5340 33928 5406 33936
rect 5340 33894 5356 33928
rect 5390 33894 5406 33928
rect 5340 33860 5406 33894
rect 5340 33826 5356 33860
rect 5390 33826 5406 33860
rect 5340 33792 5406 33826
rect 5340 33758 5356 33792
rect 5390 33758 5406 33792
rect 5340 33740 5406 33758
rect 5440 33928 5482 33970
rect 5474 33894 5482 33928
rect 5440 33860 5482 33894
rect 5474 33826 5482 33860
rect 5440 33792 5482 33826
rect 5474 33758 5482 33792
rect 5440 33742 5482 33758
rect 5340 33690 5386 33740
rect 199 33647 317 33681
rect 351 33647 385 33681
rect 419 33647 453 33681
rect 487 33647 521 33681
rect 555 33647 589 33681
rect 623 33647 657 33681
rect 691 33647 725 33681
rect 759 33647 793 33681
rect 827 33647 861 33681
rect 895 33647 929 33681
rect 963 33647 997 33681
rect 1031 33647 1065 33681
rect 1099 33647 1133 33681
rect 1167 33647 1201 33681
rect 1235 33647 1269 33681
rect 1303 33647 1421 33681
rect 199 33571 233 33647
rect 1387 33576 1421 33647
rect 199 33503 233 33537
rect 199 33435 233 33469
rect 313 33534 347 33573
rect 313 33461 347 33500
rect 409 33534 443 33573
rect 409 33461 443 33500
rect 505 33534 539 33573
rect 505 33461 539 33500
rect 601 33534 635 33573
rect 601 33461 635 33500
rect 697 33534 731 33573
rect 697 33461 731 33500
rect 793 33534 827 33573
rect 793 33461 827 33500
rect 889 33534 923 33573
rect 889 33461 923 33500
rect 985 33534 1019 33573
rect 985 33461 1019 33500
rect 1081 33534 1115 33573
rect 1081 33461 1115 33500
rect 1177 33534 1211 33573
rect 1177 33461 1211 33500
rect 1273 33534 1307 33573
rect 1273 33461 1307 33500
rect 1387 33504 1421 33537
rect 1387 33435 1421 33469
rect 199 33325 233 33401
rect 297 33389 313 33423
rect 347 33389 363 33423
rect 489 33389 505 33423
rect 539 33389 555 33423
rect 681 33389 697 33423
rect 731 33389 747 33423
rect 873 33389 889 33423
rect 923 33389 939 33423
rect 1065 33389 1081 33423
rect 1115 33389 1131 33423
rect 1257 33389 1273 33423
rect 1307 33389 1323 33423
rect 1387 33325 1421 33398
rect 199 33291 317 33325
rect 351 33291 385 33325
rect 419 33291 453 33325
rect 487 33291 521 33325
rect 555 33291 589 33325
rect 623 33291 657 33325
rect 691 33291 725 33325
rect 759 33291 793 33325
rect 827 33291 861 33325
rect 895 33291 929 33325
rect 963 33291 997 33325
rect 1031 33291 1065 33325
rect 1099 33291 1133 33325
rect 1167 33291 1201 33325
rect 1235 33291 1269 33325
rect 1303 33291 1421 33325
rect 2352 33651 2470 33685
rect 2504 33651 2538 33685
rect 2572 33651 2606 33685
rect 2640 33651 2674 33685
rect 2708 33651 2742 33685
rect 2776 33651 2810 33685
rect 2844 33651 2878 33685
rect 2912 33651 2946 33685
rect 2980 33651 3014 33685
rect 3048 33651 3082 33685
rect 3116 33651 3150 33685
rect 3184 33651 3218 33685
rect 3252 33651 3286 33685
rect 3320 33651 3354 33685
rect 3388 33651 3422 33685
rect 3456 33651 3574 33685
rect 2352 33575 2386 33651
rect 3540 33580 3574 33651
rect 3873 33651 3991 33685
rect 4025 33651 4059 33685
rect 4093 33651 4127 33685
rect 4161 33651 4195 33685
rect 4229 33651 4263 33685
rect 4297 33651 4331 33685
rect 4365 33651 4399 33685
rect 4433 33651 4467 33685
rect 4501 33651 4535 33685
rect 4569 33651 4603 33685
rect 4637 33651 4671 33685
rect 4705 33651 4739 33685
rect 4773 33651 4807 33685
rect 4841 33651 4875 33685
rect 4909 33651 4943 33685
rect 4977 33651 5095 33685
rect 3675 33615 3691 33649
rect 3725 33615 3741 33649
rect 2352 33507 2386 33541
rect 2352 33439 2386 33473
rect 2466 33538 2500 33577
rect 2466 33465 2500 33504
rect 2562 33538 2596 33577
rect 2562 33465 2596 33504
rect 2658 33538 2692 33577
rect 2658 33465 2692 33504
rect 2754 33538 2788 33577
rect 2754 33465 2788 33504
rect 2850 33538 2884 33577
rect 2850 33465 2884 33504
rect 2946 33538 2980 33577
rect 2946 33465 2980 33504
rect 3042 33538 3076 33577
rect 3042 33465 3076 33504
rect 3138 33538 3172 33577
rect 3138 33465 3172 33504
rect 3234 33538 3268 33577
rect 3234 33465 3268 33504
rect 3330 33538 3364 33577
rect 3330 33465 3364 33504
rect 3426 33538 3460 33577
rect 3426 33465 3460 33504
rect 3540 33508 3574 33541
rect 3647 33565 3681 33581
rect 3647 33473 3681 33489
rect 3735 33565 3769 33581
rect 3735 33473 3769 33489
rect 3873 33575 3907 33651
rect 5061 33580 5095 33651
rect 3873 33507 3907 33541
rect 3540 33439 3574 33473
rect 2352 33329 2386 33405
rect 2450 33393 2466 33427
rect 2500 33393 2516 33427
rect 2642 33393 2658 33427
rect 2692 33393 2708 33427
rect 2834 33393 2850 33427
rect 2884 33393 2900 33427
rect 3026 33393 3042 33427
rect 3076 33393 3092 33427
rect 3218 33393 3234 33427
rect 3268 33393 3284 33427
rect 3410 33393 3426 33427
rect 3460 33393 3476 33427
rect 3540 33329 3574 33402
rect 2352 33295 2470 33329
rect 2504 33295 2538 33329
rect 2572 33295 2606 33329
rect 2640 33295 2674 33329
rect 2708 33295 2742 33329
rect 2776 33295 2810 33329
rect 2844 33295 2878 33329
rect 2912 33295 2946 33329
rect 2980 33295 3014 33329
rect 3048 33295 3082 33329
rect 3116 33295 3150 33329
rect 3184 33295 3218 33329
rect 3252 33295 3286 33329
rect 3320 33295 3354 33329
rect 3388 33295 3422 33329
rect 3456 33295 3574 33329
rect 3873 33439 3907 33473
rect 3987 33538 4021 33577
rect 3987 33465 4021 33504
rect 4083 33538 4117 33577
rect 4083 33465 4117 33504
rect 4179 33538 4213 33577
rect 4179 33465 4213 33504
rect 4275 33538 4309 33577
rect 4275 33465 4309 33504
rect 4371 33538 4405 33577
rect 4371 33465 4405 33504
rect 4467 33538 4501 33577
rect 4467 33465 4501 33504
rect 4563 33538 4597 33577
rect 4563 33465 4597 33504
rect 4659 33538 4693 33577
rect 4659 33465 4693 33504
rect 4755 33538 4789 33577
rect 4755 33465 4789 33504
rect 4851 33538 4885 33577
rect 4851 33465 4885 33504
rect 4947 33538 4981 33577
rect 4947 33465 4981 33504
rect 5061 33508 5095 33541
rect 5340 33656 5348 33690
rect 5382 33656 5386 33690
rect 5420 33695 5486 33706
rect 5420 33692 5450 33695
rect 5420 33658 5436 33692
rect 5484 33661 5486 33695
rect 5470 33658 5486 33661
rect 5340 33620 5386 33656
rect 5340 33608 5406 33620
rect 5340 33574 5356 33608
rect 5390 33574 5406 33608
rect 5340 33540 5406 33574
rect 5340 33506 5356 33540
rect 5390 33506 5406 33540
rect 5340 33494 5406 33506
rect 5440 33608 5486 33624
rect 5474 33574 5486 33608
rect 5440 33540 5486 33574
rect 5474 33506 5486 33540
rect 5061 33439 5095 33473
rect 5440 33460 5486 33506
rect 3873 33329 3907 33405
rect 3971 33393 3987 33427
rect 4021 33393 4037 33427
rect 4163 33393 4179 33427
rect 4213 33393 4229 33427
rect 4355 33393 4371 33427
rect 4405 33393 4421 33427
rect 4547 33393 4563 33427
rect 4597 33393 4613 33427
rect 4739 33393 4755 33427
rect 4789 33393 4805 33427
rect 4931 33393 4947 33427
rect 4981 33393 4997 33427
rect 5274 33426 5303 33460
rect 5337 33426 5395 33460
rect 5429 33426 5487 33460
rect 5521 33426 5550 33460
rect 5061 33329 5095 33402
rect 3873 33295 3991 33329
rect 4025 33295 4059 33329
rect 4093 33295 4127 33329
rect 4161 33295 4195 33329
rect 4229 33295 4263 33329
rect 4297 33295 4331 33329
rect 4365 33295 4399 33329
rect 4433 33295 4467 33329
rect 4501 33295 4535 33329
rect 4569 33295 4603 33329
rect 4637 33295 4671 33329
rect 4705 33295 4739 33329
rect 4773 33295 4807 33329
rect 4841 33295 4875 33329
rect 4909 33295 4943 33329
rect 4977 33295 5095 33329
rect 199 33012 317 33046
rect 351 33012 385 33046
rect 419 33012 453 33046
rect 487 33012 521 33046
rect 555 33012 589 33046
rect 623 33012 657 33046
rect 691 33012 725 33046
rect 759 33012 793 33046
rect 827 33012 861 33046
rect 895 33012 929 33046
rect 963 33012 997 33046
rect 1031 33012 1065 33046
rect 1099 33012 1133 33046
rect 1167 33012 1201 33046
rect 1235 33012 1269 33046
rect 1303 33012 1421 33046
rect 199 32944 233 33012
rect 1387 32944 1421 33012
rect 297 32910 313 32944
rect 347 32910 363 32944
rect 489 32910 505 32944
rect 539 32910 555 32944
rect 681 32910 697 32944
rect 731 32910 747 32944
rect 873 32910 889 32944
rect 923 32910 939 32944
rect 1065 32910 1081 32944
rect 1115 32910 1131 32944
rect 1257 32910 1273 32944
rect 1307 32910 1323 32944
rect 199 32876 233 32910
rect 1387 32876 1421 32884
rect 199 32808 233 32842
rect 199 32740 233 32774
rect 199 32672 233 32706
rect 199 32604 233 32638
rect 313 32845 347 32866
rect 313 32777 347 32781
rect 313 32671 347 32675
rect 313 32586 347 32607
rect 409 32845 443 32866
rect 409 32777 443 32781
rect 409 32671 443 32675
rect 409 32586 443 32607
rect 505 32845 539 32866
rect 505 32777 539 32781
rect 505 32671 539 32675
rect 505 32586 539 32607
rect 601 32845 635 32866
rect 601 32777 635 32781
rect 601 32671 635 32675
rect 601 32586 635 32607
rect 697 32845 731 32866
rect 697 32777 731 32781
rect 697 32671 731 32675
rect 697 32586 731 32607
rect 793 32845 827 32866
rect 793 32777 827 32781
rect 793 32671 827 32675
rect 793 32586 827 32607
rect 889 32845 923 32866
rect 889 32777 923 32781
rect 889 32671 923 32675
rect 889 32586 923 32607
rect 985 32845 1019 32866
rect 985 32777 1019 32781
rect 985 32671 1019 32675
rect 985 32586 1019 32607
rect 1081 32845 1115 32866
rect 1081 32777 1115 32781
rect 1081 32671 1115 32675
rect 1081 32586 1115 32607
rect 1177 32845 1211 32866
rect 1177 32777 1211 32781
rect 1177 32671 1211 32675
rect 1177 32586 1211 32607
rect 1273 32845 1307 32866
rect 1273 32777 1307 32781
rect 1273 32671 1307 32675
rect 1273 32586 1307 32607
rect 1387 32808 1421 32812
rect 1387 32702 1421 32706
rect 1387 32630 1421 32638
rect 199 32502 233 32570
rect 1387 32502 1421 32570
rect 199 32468 317 32502
rect 351 32468 385 32502
rect 419 32468 453 32502
rect 487 32468 521 32502
rect 555 32468 589 32502
rect 623 32468 657 32502
rect 691 32468 725 32502
rect 759 32468 793 32502
rect 827 32468 861 32502
rect 895 32468 929 32502
rect 963 32468 997 32502
rect 1031 32468 1065 32502
rect 1099 32468 1133 32502
rect 1167 32468 1201 32502
rect 1235 32468 1269 32502
rect 1303 32468 1421 32502
rect 2352 33016 2470 33050
rect 2504 33016 2538 33050
rect 2572 33016 2606 33050
rect 2640 33016 2674 33050
rect 2708 33016 2742 33050
rect 2776 33016 2810 33050
rect 2844 33016 2878 33050
rect 2912 33016 2946 33050
rect 2980 33016 3014 33050
rect 3048 33016 3082 33050
rect 3116 33016 3150 33050
rect 3184 33016 3218 33050
rect 3252 33016 3286 33050
rect 3320 33016 3354 33050
rect 3388 33016 3422 33050
rect 3456 33016 3574 33050
rect 2352 32948 2386 33016
rect 3540 32948 3574 33016
rect 2450 32914 2466 32948
rect 2500 32914 2516 32948
rect 2642 32914 2658 32948
rect 2692 32914 2708 32948
rect 2834 32914 2850 32948
rect 2884 32914 2900 32948
rect 3026 32914 3042 32948
rect 3076 32914 3092 32948
rect 3218 32914 3234 32948
rect 3268 32914 3284 32948
rect 3410 32914 3426 32948
rect 3460 32914 3476 32948
rect 2352 32880 2386 32914
rect 3540 32880 3574 32888
rect 2352 32812 2386 32846
rect 2352 32744 2386 32778
rect 2352 32676 2386 32710
rect 2352 32608 2386 32642
rect 2466 32849 2500 32870
rect 2466 32781 2500 32785
rect 2466 32675 2500 32679
rect 2466 32590 2500 32611
rect 2562 32849 2596 32870
rect 2562 32781 2596 32785
rect 2562 32675 2596 32679
rect 2562 32590 2596 32611
rect 2658 32849 2692 32870
rect 2658 32781 2692 32785
rect 2658 32675 2692 32679
rect 2658 32590 2692 32611
rect 2754 32849 2788 32870
rect 2754 32781 2788 32785
rect 2754 32675 2788 32679
rect 2754 32590 2788 32611
rect 2850 32849 2884 32870
rect 2850 32781 2884 32785
rect 2850 32675 2884 32679
rect 2850 32590 2884 32611
rect 2946 32849 2980 32870
rect 2946 32781 2980 32785
rect 2946 32675 2980 32679
rect 2946 32590 2980 32611
rect 3042 32849 3076 32870
rect 3042 32781 3076 32785
rect 3042 32675 3076 32679
rect 3042 32590 3076 32611
rect 3138 32849 3172 32870
rect 3138 32781 3172 32785
rect 3138 32675 3172 32679
rect 3138 32590 3172 32611
rect 3234 32849 3268 32870
rect 3234 32781 3268 32785
rect 3234 32675 3268 32679
rect 3234 32590 3268 32611
rect 3330 32849 3364 32870
rect 3330 32781 3364 32785
rect 3330 32675 3364 32679
rect 3330 32590 3364 32611
rect 3426 32849 3460 32870
rect 3426 32781 3460 32785
rect 3426 32675 3460 32679
rect 3426 32590 3460 32611
rect 3540 32812 3574 32816
rect 3540 32706 3574 32710
rect 3540 32634 3574 32642
rect 2352 32506 2386 32574
rect 3540 32506 3574 32574
rect 2352 32472 2470 32506
rect 2504 32472 2538 32506
rect 2572 32472 2606 32506
rect 2640 32472 2674 32506
rect 2708 32472 2742 32506
rect 2776 32472 2810 32506
rect 2844 32472 2878 32506
rect 2912 32472 2946 32506
rect 2980 32472 3014 32506
rect 3048 32472 3082 32506
rect 3116 32472 3150 32506
rect 3184 32472 3218 32506
rect 3252 32472 3286 32506
rect 3320 32472 3354 32506
rect 3388 32472 3422 32506
rect 3456 32472 3574 32506
rect 3873 33016 3991 33050
rect 4025 33016 4059 33050
rect 4093 33016 4127 33050
rect 4161 33016 4195 33050
rect 4229 33016 4263 33050
rect 4297 33016 4331 33050
rect 4365 33016 4399 33050
rect 4433 33016 4467 33050
rect 4501 33016 4535 33050
rect 4569 33016 4603 33050
rect 4637 33016 4671 33050
rect 4705 33016 4739 33050
rect 4773 33016 4807 33050
rect 4841 33016 4875 33050
rect 4909 33016 4943 33050
rect 4977 33016 5095 33050
rect 3873 32948 3907 33016
rect 5061 32948 5095 33016
rect 3971 32914 3987 32948
rect 4021 32914 4037 32948
rect 4163 32914 4179 32948
rect 4213 32914 4229 32948
rect 4355 32914 4371 32948
rect 4405 32914 4421 32948
rect 4547 32914 4563 32948
rect 4597 32914 4613 32948
rect 4739 32914 4755 32948
rect 4789 32914 4805 32948
rect 4931 32914 4947 32948
rect 4981 32914 4997 32948
rect 3873 32880 3907 32914
rect 5061 32880 5095 32888
rect 3873 32812 3907 32846
rect 3873 32744 3907 32778
rect 3873 32676 3907 32710
rect 3873 32608 3907 32642
rect 3987 32849 4021 32870
rect 3987 32781 4021 32785
rect 3987 32675 4021 32679
rect 3987 32590 4021 32611
rect 4083 32849 4117 32870
rect 4083 32781 4117 32785
rect 4083 32675 4117 32679
rect 4083 32590 4117 32611
rect 4179 32849 4213 32870
rect 4179 32781 4213 32785
rect 4179 32675 4213 32679
rect 4179 32590 4213 32611
rect 4275 32849 4309 32870
rect 4275 32781 4309 32785
rect 4275 32675 4309 32679
rect 4275 32590 4309 32611
rect 4371 32849 4405 32870
rect 4371 32781 4405 32785
rect 4371 32675 4405 32679
rect 4371 32590 4405 32611
rect 4467 32849 4501 32870
rect 4467 32781 4501 32785
rect 4467 32675 4501 32679
rect 4467 32590 4501 32611
rect 4563 32849 4597 32870
rect 4563 32781 4597 32785
rect 4563 32675 4597 32679
rect 4563 32590 4597 32611
rect 4659 32849 4693 32870
rect 4659 32781 4693 32785
rect 4659 32675 4693 32679
rect 4659 32590 4693 32611
rect 4755 32849 4789 32870
rect 4755 32781 4789 32785
rect 4755 32675 4789 32679
rect 4755 32590 4789 32611
rect 4851 32849 4885 32870
rect 4851 32781 4885 32785
rect 4851 32675 4885 32679
rect 4851 32590 4885 32611
rect 4947 32849 4981 32870
rect 4947 32781 4981 32785
rect 4947 32675 4981 32679
rect 4947 32590 4981 32611
rect 5061 32812 5095 32816
rect 5061 32706 5095 32710
rect 5274 32683 5303 32717
rect 5337 32683 5395 32717
rect 5429 32683 5487 32717
rect 5521 32683 5550 32717
rect 5061 32634 5095 32642
rect 3873 32506 3907 32574
rect 5061 32506 5095 32574
rect 3873 32472 3991 32506
rect 4025 32472 4059 32506
rect 4093 32472 4127 32506
rect 4161 32472 4195 32506
rect 4229 32472 4263 32506
rect 4297 32472 4331 32506
rect 4365 32472 4399 32506
rect 4433 32472 4467 32506
rect 4501 32472 4535 32506
rect 4569 32472 4603 32506
rect 4637 32472 4671 32506
rect 4705 32472 4739 32506
rect 4773 32472 4807 32506
rect 4841 32472 4875 32506
rect 4909 32472 4943 32506
rect 4977 32472 5095 32506
rect 5340 32641 5406 32649
rect 5340 32607 5356 32641
rect 5390 32607 5406 32641
rect 5340 32573 5406 32607
rect 5340 32539 5356 32573
rect 5390 32539 5406 32573
rect 5340 32505 5406 32539
rect 5340 32471 5356 32505
rect 5390 32471 5406 32505
rect 5340 32453 5406 32471
rect 5440 32641 5482 32683
rect 5474 32607 5482 32641
rect 5440 32573 5482 32607
rect 5474 32539 5482 32573
rect 5440 32505 5482 32539
rect 5474 32471 5482 32505
rect 5440 32455 5482 32471
rect 5340 32403 5386 32453
rect 199 32360 317 32394
rect 351 32360 385 32394
rect 419 32360 453 32394
rect 487 32360 521 32394
rect 555 32360 589 32394
rect 623 32360 657 32394
rect 691 32360 725 32394
rect 759 32360 793 32394
rect 827 32360 861 32394
rect 895 32360 929 32394
rect 963 32360 997 32394
rect 1031 32360 1065 32394
rect 1099 32360 1133 32394
rect 1167 32360 1201 32394
rect 1235 32360 1269 32394
rect 1303 32360 1421 32394
rect 199 32284 233 32360
rect 1387 32289 1421 32360
rect 199 32216 233 32250
rect 199 32148 233 32182
rect 313 32247 347 32286
rect 313 32174 347 32213
rect 409 32247 443 32286
rect 409 32174 443 32213
rect 505 32247 539 32286
rect 505 32174 539 32213
rect 601 32247 635 32286
rect 601 32174 635 32213
rect 697 32247 731 32286
rect 697 32174 731 32213
rect 793 32247 827 32286
rect 793 32174 827 32213
rect 889 32247 923 32286
rect 889 32174 923 32213
rect 985 32247 1019 32286
rect 985 32174 1019 32213
rect 1081 32247 1115 32286
rect 1081 32174 1115 32213
rect 1177 32247 1211 32286
rect 1177 32174 1211 32213
rect 1273 32247 1307 32286
rect 1273 32174 1307 32213
rect 1387 32217 1421 32250
rect 1387 32148 1421 32182
rect 199 32038 233 32114
rect 297 32102 313 32136
rect 347 32102 363 32136
rect 489 32102 505 32136
rect 539 32102 555 32136
rect 681 32102 697 32136
rect 731 32102 747 32136
rect 873 32102 889 32136
rect 923 32102 939 32136
rect 1065 32102 1081 32136
rect 1115 32102 1131 32136
rect 1257 32102 1273 32136
rect 1307 32102 1323 32136
rect 1387 32038 1421 32111
rect 199 32004 317 32038
rect 351 32004 385 32038
rect 419 32004 453 32038
rect 487 32004 521 32038
rect 555 32004 589 32038
rect 623 32004 657 32038
rect 691 32004 725 32038
rect 759 32004 793 32038
rect 827 32004 861 32038
rect 895 32004 929 32038
rect 963 32004 997 32038
rect 1031 32004 1065 32038
rect 1099 32004 1133 32038
rect 1167 32004 1201 32038
rect 1235 32004 1269 32038
rect 1303 32004 1421 32038
rect 2352 32364 2470 32398
rect 2504 32364 2538 32398
rect 2572 32364 2606 32398
rect 2640 32364 2674 32398
rect 2708 32364 2742 32398
rect 2776 32364 2810 32398
rect 2844 32364 2878 32398
rect 2912 32364 2946 32398
rect 2980 32364 3014 32398
rect 3048 32364 3082 32398
rect 3116 32364 3150 32398
rect 3184 32364 3218 32398
rect 3252 32364 3286 32398
rect 3320 32364 3354 32398
rect 3388 32364 3422 32398
rect 3456 32364 3574 32398
rect 2352 32288 2386 32364
rect 3540 32293 3574 32364
rect 3873 32364 3991 32398
rect 4025 32364 4059 32398
rect 4093 32364 4127 32398
rect 4161 32364 4195 32398
rect 4229 32364 4263 32398
rect 4297 32364 4331 32398
rect 4365 32364 4399 32398
rect 4433 32364 4467 32398
rect 4501 32364 4535 32398
rect 4569 32364 4603 32398
rect 4637 32364 4671 32398
rect 4705 32364 4739 32398
rect 4773 32364 4807 32398
rect 4841 32364 4875 32398
rect 4909 32364 4943 32398
rect 4977 32364 5095 32398
rect 3675 32328 3691 32362
rect 3725 32328 3741 32362
rect 2352 32220 2386 32254
rect 2352 32152 2386 32186
rect 2466 32251 2500 32290
rect 2466 32178 2500 32217
rect 2562 32251 2596 32290
rect 2562 32178 2596 32217
rect 2658 32251 2692 32290
rect 2658 32178 2692 32217
rect 2754 32251 2788 32290
rect 2754 32178 2788 32217
rect 2850 32251 2884 32290
rect 2850 32178 2884 32217
rect 2946 32251 2980 32290
rect 2946 32178 2980 32217
rect 3042 32251 3076 32290
rect 3042 32178 3076 32217
rect 3138 32251 3172 32290
rect 3138 32178 3172 32217
rect 3234 32251 3268 32290
rect 3234 32178 3268 32217
rect 3330 32251 3364 32290
rect 3330 32178 3364 32217
rect 3426 32251 3460 32290
rect 3426 32178 3460 32217
rect 3540 32221 3574 32254
rect 3647 32278 3681 32294
rect 3647 32186 3681 32202
rect 3735 32278 3769 32294
rect 3735 32186 3769 32202
rect 3873 32288 3907 32364
rect 5061 32293 5095 32364
rect 3873 32220 3907 32254
rect 3540 32152 3574 32186
rect 2352 32042 2386 32118
rect 2450 32106 2466 32140
rect 2500 32106 2516 32140
rect 2642 32106 2658 32140
rect 2692 32106 2708 32140
rect 2834 32106 2850 32140
rect 2884 32106 2900 32140
rect 3026 32106 3042 32140
rect 3076 32106 3092 32140
rect 3218 32106 3234 32140
rect 3268 32106 3284 32140
rect 3410 32106 3426 32140
rect 3460 32106 3476 32140
rect 3540 32042 3574 32115
rect 2352 32008 2470 32042
rect 2504 32008 2538 32042
rect 2572 32008 2606 32042
rect 2640 32008 2674 32042
rect 2708 32008 2742 32042
rect 2776 32008 2810 32042
rect 2844 32008 2878 32042
rect 2912 32008 2946 32042
rect 2980 32008 3014 32042
rect 3048 32008 3082 32042
rect 3116 32008 3150 32042
rect 3184 32008 3218 32042
rect 3252 32008 3286 32042
rect 3320 32008 3354 32042
rect 3388 32008 3422 32042
rect 3456 32008 3574 32042
rect 3873 32152 3907 32186
rect 3987 32251 4021 32290
rect 3987 32178 4021 32217
rect 4083 32251 4117 32290
rect 4083 32178 4117 32217
rect 4179 32251 4213 32290
rect 4179 32178 4213 32217
rect 4275 32251 4309 32290
rect 4275 32178 4309 32217
rect 4371 32251 4405 32290
rect 4371 32178 4405 32217
rect 4467 32251 4501 32290
rect 4467 32178 4501 32217
rect 4563 32251 4597 32290
rect 4563 32178 4597 32217
rect 4659 32251 4693 32290
rect 4659 32178 4693 32217
rect 4755 32251 4789 32290
rect 4755 32178 4789 32217
rect 4851 32251 4885 32290
rect 4851 32178 4885 32217
rect 4947 32251 4981 32290
rect 4947 32178 4981 32217
rect 5061 32221 5095 32254
rect 5340 32369 5348 32403
rect 5382 32369 5386 32403
rect 5420 32408 5486 32419
rect 5420 32405 5450 32408
rect 5420 32371 5436 32405
rect 5484 32374 5486 32408
rect 5470 32371 5486 32374
rect 5340 32333 5386 32369
rect 5340 32321 5406 32333
rect 5340 32287 5356 32321
rect 5390 32287 5406 32321
rect 5340 32253 5406 32287
rect 5340 32219 5356 32253
rect 5390 32219 5406 32253
rect 5340 32207 5406 32219
rect 5440 32321 5486 32337
rect 5474 32287 5486 32321
rect 5440 32253 5486 32287
rect 5474 32219 5486 32253
rect 5061 32152 5095 32186
rect 5440 32173 5486 32219
rect 3873 32042 3907 32118
rect 3971 32106 3987 32140
rect 4021 32106 4037 32140
rect 4163 32106 4179 32140
rect 4213 32106 4229 32140
rect 4355 32106 4371 32140
rect 4405 32106 4421 32140
rect 4547 32106 4563 32140
rect 4597 32106 4613 32140
rect 4739 32106 4755 32140
rect 4789 32106 4805 32140
rect 4931 32106 4947 32140
rect 4981 32106 4997 32140
rect 5274 32139 5303 32173
rect 5337 32139 5395 32173
rect 5429 32139 5487 32173
rect 5521 32139 5550 32173
rect 5061 32042 5095 32115
rect 3873 32008 3991 32042
rect 4025 32008 4059 32042
rect 4093 32008 4127 32042
rect 4161 32008 4195 32042
rect 4229 32008 4263 32042
rect 4297 32008 4331 32042
rect 4365 32008 4399 32042
rect 4433 32008 4467 32042
rect 4501 32008 4535 32042
rect 4569 32008 4603 32042
rect 4637 32008 4671 32042
rect 4705 32008 4739 32042
rect 4773 32008 4807 32042
rect 4841 32008 4875 32042
rect 4909 32008 4943 32042
rect 4977 32008 5095 32042
rect 199 31725 317 31759
rect 351 31725 385 31759
rect 419 31725 453 31759
rect 487 31725 521 31759
rect 555 31725 589 31759
rect 623 31725 657 31759
rect 691 31725 725 31759
rect 759 31725 793 31759
rect 827 31725 861 31759
rect 895 31725 929 31759
rect 963 31725 997 31759
rect 1031 31725 1065 31759
rect 1099 31725 1133 31759
rect 1167 31725 1201 31759
rect 1235 31725 1269 31759
rect 1303 31725 1421 31759
rect 199 31657 233 31725
rect 1387 31657 1421 31725
rect 297 31623 313 31657
rect 347 31623 363 31657
rect 489 31623 505 31657
rect 539 31623 555 31657
rect 681 31623 697 31657
rect 731 31623 747 31657
rect 873 31623 889 31657
rect 923 31623 939 31657
rect 1065 31623 1081 31657
rect 1115 31623 1131 31657
rect 1257 31623 1273 31657
rect 1307 31623 1323 31657
rect 199 31589 233 31623
rect 1387 31589 1421 31597
rect 199 31521 233 31555
rect 199 31453 233 31487
rect 199 31385 233 31419
rect 199 31317 233 31351
rect 313 31558 347 31579
rect 313 31490 347 31494
rect 313 31384 347 31388
rect 313 31299 347 31320
rect 409 31558 443 31579
rect 409 31490 443 31494
rect 409 31384 443 31388
rect 409 31299 443 31320
rect 505 31558 539 31579
rect 505 31490 539 31494
rect 505 31384 539 31388
rect 505 31299 539 31320
rect 601 31558 635 31579
rect 601 31490 635 31494
rect 601 31384 635 31388
rect 601 31299 635 31320
rect 697 31558 731 31579
rect 697 31490 731 31494
rect 697 31384 731 31388
rect 697 31299 731 31320
rect 793 31558 827 31579
rect 793 31490 827 31494
rect 793 31384 827 31388
rect 793 31299 827 31320
rect 889 31558 923 31579
rect 889 31490 923 31494
rect 889 31384 923 31388
rect 889 31299 923 31320
rect 985 31558 1019 31579
rect 985 31490 1019 31494
rect 985 31384 1019 31388
rect 985 31299 1019 31320
rect 1081 31558 1115 31579
rect 1081 31490 1115 31494
rect 1081 31384 1115 31388
rect 1081 31299 1115 31320
rect 1177 31558 1211 31579
rect 1177 31490 1211 31494
rect 1177 31384 1211 31388
rect 1177 31299 1211 31320
rect 1273 31558 1307 31579
rect 1273 31490 1307 31494
rect 1273 31384 1307 31388
rect 1273 31299 1307 31320
rect 1387 31521 1421 31525
rect 1387 31415 1421 31419
rect 1387 31343 1421 31351
rect 199 31215 233 31283
rect 1387 31215 1421 31283
rect 199 31181 317 31215
rect 351 31181 385 31215
rect 419 31181 453 31215
rect 487 31181 521 31215
rect 555 31181 589 31215
rect 623 31181 657 31215
rect 691 31181 725 31215
rect 759 31181 793 31215
rect 827 31181 861 31215
rect 895 31181 929 31215
rect 963 31181 997 31215
rect 1031 31181 1065 31215
rect 1099 31181 1133 31215
rect 1167 31181 1201 31215
rect 1235 31181 1269 31215
rect 1303 31181 1421 31215
rect 2352 31729 2470 31763
rect 2504 31729 2538 31763
rect 2572 31729 2606 31763
rect 2640 31729 2674 31763
rect 2708 31729 2742 31763
rect 2776 31729 2810 31763
rect 2844 31729 2878 31763
rect 2912 31729 2946 31763
rect 2980 31729 3014 31763
rect 3048 31729 3082 31763
rect 3116 31729 3150 31763
rect 3184 31729 3218 31763
rect 3252 31729 3286 31763
rect 3320 31729 3354 31763
rect 3388 31729 3422 31763
rect 3456 31729 3574 31763
rect 2352 31661 2386 31729
rect 3540 31661 3574 31729
rect 2450 31627 2466 31661
rect 2500 31627 2516 31661
rect 2642 31627 2658 31661
rect 2692 31627 2708 31661
rect 2834 31627 2850 31661
rect 2884 31627 2900 31661
rect 3026 31627 3042 31661
rect 3076 31627 3092 31661
rect 3218 31627 3234 31661
rect 3268 31627 3284 31661
rect 3410 31627 3426 31661
rect 3460 31627 3476 31661
rect 2352 31593 2386 31627
rect 3540 31593 3574 31601
rect 2352 31525 2386 31559
rect 2352 31457 2386 31491
rect 2352 31389 2386 31423
rect 2352 31321 2386 31355
rect 2466 31562 2500 31583
rect 2466 31494 2500 31498
rect 2466 31388 2500 31392
rect 2466 31303 2500 31324
rect 2562 31562 2596 31583
rect 2562 31494 2596 31498
rect 2562 31388 2596 31392
rect 2562 31303 2596 31324
rect 2658 31562 2692 31583
rect 2658 31494 2692 31498
rect 2658 31388 2692 31392
rect 2658 31303 2692 31324
rect 2754 31562 2788 31583
rect 2754 31494 2788 31498
rect 2754 31388 2788 31392
rect 2754 31303 2788 31324
rect 2850 31562 2884 31583
rect 2850 31494 2884 31498
rect 2850 31388 2884 31392
rect 2850 31303 2884 31324
rect 2946 31562 2980 31583
rect 2946 31494 2980 31498
rect 2946 31388 2980 31392
rect 2946 31303 2980 31324
rect 3042 31562 3076 31583
rect 3042 31494 3076 31498
rect 3042 31388 3076 31392
rect 3042 31303 3076 31324
rect 3138 31562 3172 31583
rect 3138 31494 3172 31498
rect 3138 31388 3172 31392
rect 3138 31303 3172 31324
rect 3234 31562 3268 31583
rect 3234 31494 3268 31498
rect 3234 31388 3268 31392
rect 3234 31303 3268 31324
rect 3330 31562 3364 31583
rect 3330 31494 3364 31498
rect 3330 31388 3364 31392
rect 3330 31303 3364 31324
rect 3426 31562 3460 31583
rect 3426 31494 3460 31498
rect 3426 31388 3460 31392
rect 3426 31303 3460 31324
rect 3540 31525 3574 31529
rect 3540 31419 3574 31423
rect 3540 31347 3574 31355
rect 2352 31219 2386 31287
rect 3540 31219 3574 31287
rect 2352 31185 2470 31219
rect 2504 31185 2538 31219
rect 2572 31185 2606 31219
rect 2640 31185 2674 31219
rect 2708 31185 2742 31219
rect 2776 31185 2810 31219
rect 2844 31185 2878 31219
rect 2912 31185 2946 31219
rect 2980 31185 3014 31219
rect 3048 31185 3082 31219
rect 3116 31185 3150 31219
rect 3184 31185 3218 31219
rect 3252 31185 3286 31219
rect 3320 31185 3354 31219
rect 3388 31185 3422 31219
rect 3456 31185 3574 31219
rect 3873 31729 3991 31763
rect 4025 31729 4059 31763
rect 4093 31729 4127 31763
rect 4161 31729 4195 31763
rect 4229 31729 4263 31763
rect 4297 31729 4331 31763
rect 4365 31729 4399 31763
rect 4433 31729 4467 31763
rect 4501 31729 4535 31763
rect 4569 31729 4603 31763
rect 4637 31729 4671 31763
rect 4705 31729 4739 31763
rect 4773 31729 4807 31763
rect 4841 31729 4875 31763
rect 4909 31729 4943 31763
rect 4977 31729 5095 31763
rect 3873 31661 3907 31729
rect 5061 31661 5095 31729
rect 3971 31627 3987 31661
rect 4021 31627 4037 31661
rect 4163 31627 4179 31661
rect 4213 31627 4229 31661
rect 4355 31627 4371 31661
rect 4405 31627 4421 31661
rect 4547 31627 4563 31661
rect 4597 31627 4613 31661
rect 4739 31627 4755 31661
rect 4789 31627 4805 31661
rect 4931 31627 4947 31661
rect 4981 31627 4997 31661
rect 3873 31593 3907 31627
rect 5061 31593 5095 31601
rect 3873 31525 3907 31559
rect 3873 31457 3907 31491
rect 3873 31389 3907 31423
rect 3873 31321 3907 31355
rect 3987 31562 4021 31583
rect 3987 31494 4021 31498
rect 3987 31388 4021 31392
rect 3987 31303 4021 31324
rect 4083 31562 4117 31583
rect 4083 31494 4117 31498
rect 4083 31388 4117 31392
rect 4083 31303 4117 31324
rect 4179 31562 4213 31583
rect 4179 31494 4213 31498
rect 4179 31388 4213 31392
rect 4179 31303 4213 31324
rect 4275 31562 4309 31583
rect 4275 31494 4309 31498
rect 4275 31388 4309 31392
rect 4275 31303 4309 31324
rect 4371 31562 4405 31583
rect 4371 31494 4405 31498
rect 4371 31388 4405 31392
rect 4371 31303 4405 31324
rect 4467 31562 4501 31583
rect 4467 31494 4501 31498
rect 4467 31388 4501 31392
rect 4467 31303 4501 31324
rect 4563 31562 4597 31583
rect 4563 31494 4597 31498
rect 4563 31388 4597 31392
rect 4563 31303 4597 31324
rect 4659 31562 4693 31583
rect 4659 31494 4693 31498
rect 4659 31388 4693 31392
rect 4659 31303 4693 31324
rect 4755 31562 4789 31583
rect 4755 31494 4789 31498
rect 4755 31388 4789 31392
rect 4755 31303 4789 31324
rect 4851 31562 4885 31583
rect 4851 31494 4885 31498
rect 4851 31388 4885 31392
rect 4851 31303 4885 31324
rect 4947 31562 4981 31583
rect 4947 31494 4981 31498
rect 4947 31388 4981 31392
rect 4947 31303 4981 31324
rect 5061 31525 5095 31529
rect 5061 31419 5095 31423
rect 5274 31396 5303 31430
rect 5337 31396 5395 31430
rect 5429 31396 5487 31430
rect 5521 31396 5550 31430
rect 5061 31347 5095 31355
rect 3873 31219 3907 31287
rect 5061 31219 5095 31287
rect 3873 31185 3991 31219
rect 4025 31185 4059 31219
rect 4093 31185 4127 31219
rect 4161 31185 4195 31219
rect 4229 31185 4263 31219
rect 4297 31185 4331 31219
rect 4365 31185 4399 31219
rect 4433 31185 4467 31219
rect 4501 31185 4535 31219
rect 4569 31185 4603 31219
rect 4637 31185 4671 31219
rect 4705 31185 4739 31219
rect 4773 31185 4807 31219
rect 4841 31185 4875 31219
rect 4909 31185 4943 31219
rect 4977 31185 5095 31219
rect 5340 31354 5406 31362
rect 5340 31320 5356 31354
rect 5390 31320 5406 31354
rect 5340 31286 5406 31320
rect 5340 31252 5356 31286
rect 5390 31252 5406 31286
rect 5340 31218 5406 31252
rect 5340 31184 5356 31218
rect 5390 31184 5406 31218
rect 5340 31166 5406 31184
rect 5440 31354 5482 31396
rect 5474 31320 5482 31354
rect 5440 31286 5482 31320
rect 5474 31252 5482 31286
rect 5440 31218 5482 31252
rect 5474 31184 5482 31218
rect 5440 31168 5482 31184
rect 5340 31116 5386 31166
rect 199 31073 317 31107
rect 351 31073 385 31107
rect 419 31073 453 31107
rect 487 31073 521 31107
rect 555 31073 589 31107
rect 623 31073 657 31107
rect 691 31073 725 31107
rect 759 31073 793 31107
rect 827 31073 861 31107
rect 895 31073 929 31107
rect 963 31073 997 31107
rect 1031 31073 1065 31107
rect 1099 31073 1133 31107
rect 1167 31073 1201 31107
rect 1235 31073 1269 31107
rect 1303 31073 1421 31107
rect 199 30997 233 31073
rect 1387 31002 1421 31073
rect 199 30929 233 30963
rect 199 30861 233 30895
rect 313 30960 347 30999
rect 313 30887 347 30926
rect 409 30960 443 30999
rect 409 30887 443 30926
rect 505 30960 539 30999
rect 505 30887 539 30926
rect 601 30960 635 30999
rect 601 30887 635 30926
rect 697 30960 731 30999
rect 697 30887 731 30926
rect 793 30960 827 30999
rect 793 30887 827 30926
rect 889 30960 923 30999
rect 889 30887 923 30926
rect 985 30960 1019 30999
rect 985 30887 1019 30926
rect 1081 30960 1115 30999
rect 1081 30887 1115 30926
rect 1177 30960 1211 30999
rect 1177 30887 1211 30926
rect 1273 30960 1307 30999
rect 1273 30887 1307 30926
rect 1387 30930 1421 30963
rect 1387 30861 1421 30895
rect 199 30751 233 30827
rect 297 30815 313 30849
rect 347 30815 363 30849
rect 489 30815 505 30849
rect 539 30815 555 30849
rect 681 30815 697 30849
rect 731 30815 747 30849
rect 873 30815 889 30849
rect 923 30815 939 30849
rect 1065 30815 1081 30849
rect 1115 30815 1131 30849
rect 1257 30815 1273 30849
rect 1307 30815 1323 30849
rect 1387 30751 1421 30824
rect 199 30717 317 30751
rect 351 30717 385 30751
rect 419 30717 453 30751
rect 487 30717 521 30751
rect 555 30717 589 30751
rect 623 30717 657 30751
rect 691 30717 725 30751
rect 759 30717 793 30751
rect 827 30717 861 30751
rect 895 30717 929 30751
rect 963 30717 997 30751
rect 1031 30717 1065 30751
rect 1099 30717 1133 30751
rect 1167 30717 1201 30751
rect 1235 30717 1269 30751
rect 1303 30717 1421 30751
rect 2352 31077 2470 31111
rect 2504 31077 2538 31111
rect 2572 31077 2606 31111
rect 2640 31077 2674 31111
rect 2708 31077 2742 31111
rect 2776 31077 2810 31111
rect 2844 31077 2878 31111
rect 2912 31077 2946 31111
rect 2980 31077 3014 31111
rect 3048 31077 3082 31111
rect 3116 31077 3150 31111
rect 3184 31077 3218 31111
rect 3252 31077 3286 31111
rect 3320 31077 3354 31111
rect 3388 31077 3422 31111
rect 3456 31077 3574 31111
rect 2352 31001 2386 31077
rect 3540 31006 3574 31077
rect 3873 31077 3991 31111
rect 4025 31077 4059 31111
rect 4093 31077 4127 31111
rect 4161 31077 4195 31111
rect 4229 31077 4263 31111
rect 4297 31077 4331 31111
rect 4365 31077 4399 31111
rect 4433 31077 4467 31111
rect 4501 31077 4535 31111
rect 4569 31077 4603 31111
rect 4637 31077 4671 31111
rect 4705 31077 4739 31111
rect 4773 31077 4807 31111
rect 4841 31077 4875 31111
rect 4909 31077 4943 31111
rect 4977 31077 5095 31111
rect 3675 31041 3691 31075
rect 3725 31041 3741 31075
rect 2352 30933 2386 30967
rect 2352 30865 2386 30899
rect 2466 30964 2500 31003
rect 2466 30891 2500 30930
rect 2562 30964 2596 31003
rect 2562 30891 2596 30930
rect 2658 30964 2692 31003
rect 2658 30891 2692 30930
rect 2754 30964 2788 31003
rect 2754 30891 2788 30930
rect 2850 30964 2884 31003
rect 2850 30891 2884 30930
rect 2946 30964 2980 31003
rect 2946 30891 2980 30930
rect 3042 30964 3076 31003
rect 3042 30891 3076 30930
rect 3138 30964 3172 31003
rect 3138 30891 3172 30930
rect 3234 30964 3268 31003
rect 3234 30891 3268 30930
rect 3330 30964 3364 31003
rect 3330 30891 3364 30930
rect 3426 30964 3460 31003
rect 3426 30891 3460 30930
rect 3540 30934 3574 30967
rect 3647 30991 3681 31007
rect 3647 30899 3681 30915
rect 3735 30991 3769 31007
rect 3735 30899 3769 30915
rect 3873 31001 3907 31077
rect 5061 31006 5095 31077
rect 3873 30933 3907 30967
rect 3540 30865 3574 30899
rect 2352 30755 2386 30831
rect 2450 30819 2466 30853
rect 2500 30819 2516 30853
rect 2642 30819 2658 30853
rect 2692 30819 2708 30853
rect 2834 30819 2850 30853
rect 2884 30819 2900 30853
rect 3026 30819 3042 30853
rect 3076 30819 3092 30853
rect 3218 30819 3234 30853
rect 3268 30819 3284 30853
rect 3410 30819 3426 30853
rect 3460 30819 3476 30853
rect 3540 30755 3574 30828
rect 2352 30721 2470 30755
rect 2504 30721 2538 30755
rect 2572 30721 2606 30755
rect 2640 30721 2674 30755
rect 2708 30721 2742 30755
rect 2776 30721 2810 30755
rect 2844 30721 2878 30755
rect 2912 30721 2946 30755
rect 2980 30721 3014 30755
rect 3048 30721 3082 30755
rect 3116 30721 3150 30755
rect 3184 30721 3218 30755
rect 3252 30721 3286 30755
rect 3320 30721 3354 30755
rect 3388 30721 3422 30755
rect 3456 30721 3574 30755
rect 3873 30865 3907 30899
rect 3987 30964 4021 31003
rect 3987 30891 4021 30930
rect 4083 30964 4117 31003
rect 4083 30891 4117 30930
rect 4179 30964 4213 31003
rect 4179 30891 4213 30930
rect 4275 30964 4309 31003
rect 4275 30891 4309 30930
rect 4371 30964 4405 31003
rect 4371 30891 4405 30930
rect 4467 30964 4501 31003
rect 4467 30891 4501 30930
rect 4563 30964 4597 31003
rect 4563 30891 4597 30930
rect 4659 30964 4693 31003
rect 4659 30891 4693 30930
rect 4755 30964 4789 31003
rect 4755 30891 4789 30930
rect 4851 30964 4885 31003
rect 4851 30891 4885 30930
rect 4947 30964 4981 31003
rect 4947 30891 4981 30930
rect 5061 30934 5095 30967
rect 5340 31082 5348 31116
rect 5382 31082 5386 31116
rect 5420 31121 5486 31132
rect 5420 31118 5450 31121
rect 5420 31084 5436 31118
rect 5484 31087 5486 31121
rect 5470 31084 5486 31087
rect 5340 31046 5386 31082
rect 5340 31034 5406 31046
rect 5340 31000 5356 31034
rect 5390 31000 5406 31034
rect 5340 30966 5406 31000
rect 5340 30932 5356 30966
rect 5390 30932 5406 30966
rect 5340 30920 5406 30932
rect 5440 31034 5486 31050
rect 5474 31000 5486 31034
rect 5440 30966 5486 31000
rect 5474 30932 5486 30966
rect 5061 30865 5095 30899
rect 5440 30886 5486 30932
rect 3873 30755 3907 30831
rect 3971 30819 3987 30853
rect 4021 30819 4037 30853
rect 4163 30819 4179 30853
rect 4213 30819 4229 30853
rect 4355 30819 4371 30853
rect 4405 30819 4421 30853
rect 4547 30819 4563 30853
rect 4597 30819 4613 30853
rect 4739 30819 4755 30853
rect 4789 30819 4805 30853
rect 4931 30819 4947 30853
rect 4981 30819 4997 30853
rect 5274 30852 5303 30886
rect 5337 30852 5395 30886
rect 5429 30852 5487 30886
rect 5521 30852 5550 30886
rect 5061 30755 5095 30828
rect 3873 30721 3991 30755
rect 4025 30721 4059 30755
rect 4093 30721 4127 30755
rect 4161 30721 4195 30755
rect 4229 30721 4263 30755
rect 4297 30721 4331 30755
rect 4365 30721 4399 30755
rect 4433 30721 4467 30755
rect 4501 30721 4535 30755
rect 4569 30721 4603 30755
rect 4637 30721 4671 30755
rect 4705 30721 4739 30755
rect 4773 30721 4807 30755
rect 4841 30721 4875 30755
rect 4909 30721 4943 30755
rect 4977 30721 5095 30755
rect 199 30438 317 30472
rect 351 30438 385 30472
rect 419 30438 453 30472
rect 487 30438 521 30472
rect 555 30438 589 30472
rect 623 30438 657 30472
rect 691 30438 725 30472
rect 759 30438 793 30472
rect 827 30438 861 30472
rect 895 30438 929 30472
rect 963 30438 997 30472
rect 1031 30438 1065 30472
rect 1099 30438 1133 30472
rect 1167 30438 1201 30472
rect 1235 30438 1269 30472
rect 1303 30438 1421 30472
rect 199 30370 233 30438
rect 1387 30370 1421 30438
rect 297 30336 313 30370
rect 347 30336 363 30370
rect 489 30336 505 30370
rect 539 30336 555 30370
rect 681 30336 697 30370
rect 731 30336 747 30370
rect 873 30336 889 30370
rect 923 30336 939 30370
rect 1065 30336 1081 30370
rect 1115 30336 1131 30370
rect 1257 30336 1273 30370
rect 1307 30336 1323 30370
rect 199 30302 233 30336
rect 1387 30302 1421 30310
rect 199 30234 233 30268
rect 199 30166 233 30200
rect 199 30098 233 30132
rect 199 30030 233 30064
rect 313 30271 347 30292
rect 313 30203 347 30207
rect 313 30097 347 30101
rect 313 30012 347 30033
rect 409 30271 443 30292
rect 409 30203 443 30207
rect 409 30097 443 30101
rect 409 30012 443 30033
rect 505 30271 539 30292
rect 505 30203 539 30207
rect 505 30097 539 30101
rect 505 30012 539 30033
rect 601 30271 635 30292
rect 601 30203 635 30207
rect 601 30097 635 30101
rect 601 30012 635 30033
rect 697 30271 731 30292
rect 697 30203 731 30207
rect 697 30097 731 30101
rect 697 30012 731 30033
rect 793 30271 827 30292
rect 793 30203 827 30207
rect 793 30097 827 30101
rect 793 30012 827 30033
rect 889 30271 923 30292
rect 889 30203 923 30207
rect 889 30097 923 30101
rect 889 30012 923 30033
rect 985 30271 1019 30292
rect 985 30203 1019 30207
rect 985 30097 1019 30101
rect 985 30012 1019 30033
rect 1081 30271 1115 30292
rect 1081 30203 1115 30207
rect 1081 30097 1115 30101
rect 1081 30012 1115 30033
rect 1177 30271 1211 30292
rect 1177 30203 1211 30207
rect 1177 30097 1211 30101
rect 1177 30012 1211 30033
rect 1273 30271 1307 30292
rect 1273 30203 1307 30207
rect 1273 30097 1307 30101
rect 1273 30012 1307 30033
rect 1387 30234 1421 30238
rect 1387 30128 1421 30132
rect 1387 30056 1421 30064
rect 199 29928 233 29996
rect 1387 29928 1421 29996
rect 199 29894 317 29928
rect 351 29894 385 29928
rect 419 29894 453 29928
rect 487 29894 521 29928
rect 555 29894 589 29928
rect 623 29894 657 29928
rect 691 29894 725 29928
rect 759 29894 793 29928
rect 827 29894 861 29928
rect 895 29894 929 29928
rect 963 29894 997 29928
rect 1031 29894 1065 29928
rect 1099 29894 1133 29928
rect 1167 29894 1201 29928
rect 1235 29894 1269 29928
rect 1303 29894 1421 29928
rect 2352 30442 2470 30476
rect 2504 30442 2538 30476
rect 2572 30442 2606 30476
rect 2640 30442 2674 30476
rect 2708 30442 2742 30476
rect 2776 30442 2810 30476
rect 2844 30442 2878 30476
rect 2912 30442 2946 30476
rect 2980 30442 3014 30476
rect 3048 30442 3082 30476
rect 3116 30442 3150 30476
rect 3184 30442 3218 30476
rect 3252 30442 3286 30476
rect 3320 30442 3354 30476
rect 3388 30442 3422 30476
rect 3456 30442 3574 30476
rect 2352 30374 2386 30442
rect 3540 30374 3574 30442
rect 2450 30340 2466 30374
rect 2500 30340 2516 30374
rect 2642 30340 2658 30374
rect 2692 30340 2708 30374
rect 2834 30340 2850 30374
rect 2884 30340 2900 30374
rect 3026 30340 3042 30374
rect 3076 30340 3092 30374
rect 3218 30340 3234 30374
rect 3268 30340 3284 30374
rect 3410 30340 3426 30374
rect 3460 30340 3476 30374
rect 2352 30306 2386 30340
rect 3540 30306 3574 30314
rect 2352 30238 2386 30272
rect 2352 30170 2386 30204
rect 2352 30102 2386 30136
rect 2352 30034 2386 30068
rect 2466 30275 2500 30296
rect 2466 30207 2500 30211
rect 2466 30101 2500 30105
rect 2466 30016 2500 30037
rect 2562 30275 2596 30296
rect 2562 30207 2596 30211
rect 2562 30101 2596 30105
rect 2562 30016 2596 30037
rect 2658 30275 2692 30296
rect 2658 30207 2692 30211
rect 2658 30101 2692 30105
rect 2658 30016 2692 30037
rect 2754 30275 2788 30296
rect 2754 30207 2788 30211
rect 2754 30101 2788 30105
rect 2754 30016 2788 30037
rect 2850 30275 2884 30296
rect 2850 30207 2884 30211
rect 2850 30101 2884 30105
rect 2850 30016 2884 30037
rect 2946 30275 2980 30296
rect 2946 30207 2980 30211
rect 2946 30101 2980 30105
rect 2946 30016 2980 30037
rect 3042 30275 3076 30296
rect 3042 30207 3076 30211
rect 3042 30101 3076 30105
rect 3042 30016 3076 30037
rect 3138 30275 3172 30296
rect 3138 30207 3172 30211
rect 3138 30101 3172 30105
rect 3138 30016 3172 30037
rect 3234 30275 3268 30296
rect 3234 30207 3268 30211
rect 3234 30101 3268 30105
rect 3234 30016 3268 30037
rect 3330 30275 3364 30296
rect 3330 30207 3364 30211
rect 3330 30101 3364 30105
rect 3330 30016 3364 30037
rect 3426 30275 3460 30296
rect 3426 30207 3460 30211
rect 3426 30101 3460 30105
rect 3426 30016 3460 30037
rect 3540 30238 3574 30242
rect 3540 30132 3574 30136
rect 3540 30060 3574 30068
rect 2352 29932 2386 30000
rect 3540 29932 3574 30000
rect 2352 29898 2470 29932
rect 2504 29898 2538 29932
rect 2572 29898 2606 29932
rect 2640 29898 2674 29932
rect 2708 29898 2742 29932
rect 2776 29898 2810 29932
rect 2844 29898 2878 29932
rect 2912 29898 2946 29932
rect 2980 29898 3014 29932
rect 3048 29898 3082 29932
rect 3116 29898 3150 29932
rect 3184 29898 3218 29932
rect 3252 29898 3286 29932
rect 3320 29898 3354 29932
rect 3388 29898 3422 29932
rect 3456 29898 3574 29932
rect 3873 30442 3991 30476
rect 4025 30442 4059 30476
rect 4093 30442 4127 30476
rect 4161 30442 4195 30476
rect 4229 30442 4263 30476
rect 4297 30442 4331 30476
rect 4365 30442 4399 30476
rect 4433 30442 4467 30476
rect 4501 30442 4535 30476
rect 4569 30442 4603 30476
rect 4637 30442 4671 30476
rect 4705 30442 4739 30476
rect 4773 30442 4807 30476
rect 4841 30442 4875 30476
rect 4909 30442 4943 30476
rect 4977 30442 5095 30476
rect 3873 30374 3907 30442
rect 5061 30374 5095 30442
rect 3971 30340 3987 30374
rect 4021 30340 4037 30374
rect 4163 30340 4179 30374
rect 4213 30340 4229 30374
rect 4355 30340 4371 30374
rect 4405 30340 4421 30374
rect 4547 30340 4563 30374
rect 4597 30340 4613 30374
rect 4739 30340 4755 30374
rect 4789 30340 4805 30374
rect 4931 30340 4947 30374
rect 4981 30340 4997 30374
rect 3873 30306 3907 30340
rect 5061 30306 5095 30314
rect 3873 30238 3907 30272
rect 3873 30170 3907 30204
rect 3873 30102 3907 30136
rect 3873 30034 3907 30068
rect 3987 30275 4021 30296
rect 3987 30207 4021 30211
rect 3987 30101 4021 30105
rect 3987 30016 4021 30037
rect 4083 30275 4117 30296
rect 4083 30207 4117 30211
rect 4083 30101 4117 30105
rect 4083 30016 4117 30037
rect 4179 30275 4213 30296
rect 4179 30207 4213 30211
rect 4179 30101 4213 30105
rect 4179 30016 4213 30037
rect 4275 30275 4309 30296
rect 4275 30207 4309 30211
rect 4275 30101 4309 30105
rect 4275 30016 4309 30037
rect 4371 30275 4405 30296
rect 4371 30207 4405 30211
rect 4371 30101 4405 30105
rect 4371 30016 4405 30037
rect 4467 30275 4501 30296
rect 4467 30207 4501 30211
rect 4467 30101 4501 30105
rect 4467 30016 4501 30037
rect 4563 30275 4597 30296
rect 4563 30207 4597 30211
rect 4563 30101 4597 30105
rect 4563 30016 4597 30037
rect 4659 30275 4693 30296
rect 4659 30207 4693 30211
rect 4659 30101 4693 30105
rect 4659 30016 4693 30037
rect 4755 30275 4789 30296
rect 4755 30207 4789 30211
rect 4755 30101 4789 30105
rect 4755 30016 4789 30037
rect 4851 30275 4885 30296
rect 4851 30207 4885 30211
rect 4851 30101 4885 30105
rect 4851 30016 4885 30037
rect 4947 30275 4981 30296
rect 4947 30207 4981 30211
rect 4947 30101 4981 30105
rect 4947 30016 4981 30037
rect 5061 30238 5095 30242
rect 5061 30132 5095 30136
rect 5274 30109 5303 30143
rect 5337 30109 5395 30143
rect 5429 30109 5487 30143
rect 5521 30109 5550 30143
rect 5061 30060 5095 30068
rect 3873 29932 3907 30000
rect 5061 29932 5095 30000
rect 3873 29898 3991 29932
rect 4025 29898 4059 29932
rect 4093 29898 4127 29932
rect 4161 29898 4195 29932
rect 4229 29898 4263 29932
rect 4297 29898 4331 29932
rect 4365 29898 4399 29932
rect 4433 29898 4467 29932
rect 4501 29898 4535 29932
rect 4569 29898 4603 29932
rect 4637 29898 4671 29932
rect 4705 29898 4739 29932
rect 4773 29898 4807 29932
rect 4841 29898 4875 29932
rect 4909 29898 4943 29932
rect 4977 29898 5095 29932
rect 5340 30067 5406 30075
rect 5340 30033 5356 30067
rect 5390 30033 5406 30067
rect 5340 29999 5406 30033
rect 5340 29965 5356 29999
rect 5390 29965 5406 29999
rect 5340 29931 5406 29965
rect 5340 29897 5356 29931
rect 5390 29897 5406 29931
rect 5340 29879 5406 29897
rect 5440 30067 5482 30109
rect 5474 30033 5482 30067
rect 5440 29999 5482 30033
rect 5474 29965 5482 29999
rect 5440 29931 5482 29965
rect 5474 29897 5482 29931
rect 5440 29881 5482 29897
rect 5340 29829 5386 29879
rect 199 29786 317 29820
rect 351 29786 385 29820
rect 419 29786 453 29820
rect 487 29786 521 29820
rect 555 29786 589 29820
rect 623 29786 657 29820
rect 691 29786 725 29820
rect 759 29786 793 29820
rect 827 29786 861 29820
rect 895 29786 929 29820
rect 963 29786 997 29820
rect 1031 29786 1065 29820
rect 1099 29786 1133 29820
rect 1167 29786 1201 29820
rect 1235 29786 1269 29820
rect 1303 29786 1421 29820
rect 199 29710 233 29786
rect 1387 29715 1421 29786
rect 199 29642 233 29676
rect 199 29574 233 29608
rect 313 29673 347 29712
rect 313 29600 347 29639
rect 409 29673 443 29712
rect 409 29600 443 29639
rect 505 29673 539 29712
rect 505 29600 539 29639
rect 601 29673 635 29712
rect 601 29600 635 29639
rect 697 29673 731 29712
rect 697 29600 731 29639
rect 793 29673 827 29712
rect 793 29600 827 29639
rect 889 29673 923 29712
rect 889 29600 923 29639
rect 985 29673 1019 29712
rect 985 29600 1019 29639
rect 1081 29673 1115 29712
rect 1081 29600 1115 29639
rect 1177 29673 1211 29712
rect 1177 29600 1211 29639
rect 1273 29673 1307 29712
rect 1273 29600 1307 29639
rect 1387 29643 1421 29676
rect 1387 29574 1421 29608
rect 199 29464 233 29540
rect 297 29528 313 29562
rect 347 29528 363 29562
rect 489 29528 505 29562
rect 539 29528 555 29562
rect 681 29528 697 29562
rect 731 29528 747 29562
rect 873 29528 889 29562
rect 923 29528 939 29562
rect 1065 29528 1081 29562
rect 1115 29528 1131 29562
rect 1257 29528 1273 29562
rect 1307 29528 1323 29562
rect 1387 29464 1421 29537
rect 199 29430 317 29464
rect 351 29430 385 29464
rect 419 29430 453 29464
rect 487 29430 521 29464
rect 555 29430 589 29464
rect 623 29430 657 29464
rect 691 29430 725 29464
rect 759 29430 793 29464
rect 827 29430 861 29464
rect 895 29430 929 29464
rect 963 29430 997 29464
rect 1031 29430 1065 29464
rect 1099 29430 1133 29464
rect 1167 29430 1201 29464
rect 1235 29430 1269 29464
rect 1303 29430 1421 29464
rect 2352 29790 2470 29824
rect 2504 29790 2538 29824
rect 2572 29790 2606 29824
rect 2640 29790 2674 29824
rect 2708 29790 2742 29824
rect 2776 29790 2810 29824
rect 2844 29790 2878 29824
rect 2912 29790 2946 29824
rect 2980 29790 3014 29824
rect 3048 29790 3082 29824
rect 3116 29790 3150 29824
rect 3184 29790 3218 29824
rect 3252 29790 3286 29824
rect 3320 29790 3354 29824
rect 3388 29790 3422 29824
rect 3456 29790 3574 29824
rect 2352 29714 2386 29790
rect 3540 29719 3574 29790
rect 3873 29790 3991 29824
rect 4025 29790 4059 29824
rect 4093 29790 4127 29824
rect 4161 29790 4195 29824
rect 4229 29790 4263 29824
rect 4297 29790 4331 29824
rect 4365 29790 4399 29824
rect 4433 29790 4467 29824
rect 4501 29790 4535 29824
rect 4569 29790 4603 29824
rect 4637 29790 4671 29824
rect 4705 29790 4739 29824
rect 4773 29790 4807 29824
rect 4841 29790 4875 29824
rect 4909 29790 4943 29824
rect 4977 29790 5095 29824
rect 3675 29754 3691 29788
rect 3725 29754 3741 29788
rect 2352 29646 2386 29680
rect 2352 29578 2386 29612
rect 2466 29677 2500 29716
rect 2466 29604 2500 29643
rect 2562 29677 2596 29716
rect 2562 29604 2596 29643
rect 2658 29677 2692 29716
rect 2658 29604 2692 29643
rect 2754 29677 2788 29716
rect 2754 29604 2788 29643
rect 2850 29677 2884 29716
rect 2850 29604 2884 29643
rect 2946 29677 2980 29716
rect 2946 29604 2980 29643
rect 3042 29677 3076 29716
rect 3042 29604 3076 29643
rect 3138 29677 3172 29716
rect 3138 29604 3172 29643
rect 3234 29677 3268 29716
rect 3234 29604 3268 29643
rect 3330 29677 3364 29716
rect 3330 29604 3364 29643
rect 3426 29677 3460 29716
rect 3426 29604 3460 29643
rect 3540 29647 3574 29680
rect 3647 29704 3681 29720
rect 3647 29612 3681 29628
rect 3735 29704 3769 29720
rect 3735 29612 3769 29628
rect 3873 29714 3907 29790
rect 5061 29719 5095 29790
rect 3873 29646 3907 29680
rect 3540 29578 3574 29612
rect 2352 29468 2386 29544
rect 2450 29532 2466 29566
rect 2500 29532 2516 29566
rect 2642 29532 2658 29566
rect 2692 29532 2708 29566
rect 2834 29532 2850 29566
rect 2884 29532 2900 29566
rect 3026 29532 3042 29566
rect 3076 29532 3092 29566
rect 3218 29532 3234 29566
rect 3268 29532 3284 29566
rect 3410 29532 3426 29566
rect 3460 29532 3476 29566
rect 3540 29468 3574 29541
rect 2352 29434 2470 29468
rect 2504 29434 2538 29468
rect 2572 29434 2606 29468
rect 2640 29434 2674 29468
rect 2708 29434 2742 29468
rect 2776 29434 2810 29468
rect 2844 29434 2878 29468
rect 2912 29434 2946 29468
rect 2980 29434 3014 29468
rect 3048 29434 3082 29468
rect 3116 29434 3150 29468
rect 3184 29434 3218 29468
rect 3252 29434 3286 29468
rect 3320 29434 3354 29468
rect 3388 29434 3422 29468
rect 3456 29434 3574 29468
rect 3873 29578 3907 29612
rect 3987 29677 4021 29716
rect 3987 29604 4021 29643
rect 4083 29677 4117 29716
rect 4083 29604 4117 29643
rect 4179 29677 4213 29716
rect 4179 29604 4213 29643
rect 4275 29677 4309 29716
rect 4275 29604 4309 29643
rect 4371 29677 4405 29716
rect 4371 29604 4405 29643
rect 4467 29677 4501 29716
rect 4467 29604 4501 29643
rect 4563 29677 4597 29716
rect 4563 29604 4597 29643
rect 4659 29677 4693 29716
rect 4659 29604 4693 29643
rect 4755 29677 4789 29716
rect 4755 29604 4789 29643
rect 4851 29677 4885 29716
rect 4851 29604 4885 29643
rect 4947 29677 4981 29716
rect 4947 29604 4981 29643
rect 5061 29647 5095 29680
rect 5340 29795 5348 29829
rect 5382 29795 5386 29829
rect 5420 29834 5486 29845
rect 5420 29831 5450 29834
rect 5420 29797 5436 29831
rect 5484 29800 5486 29834
rect 5470 29797 5486 29800
rect 5340 29759 5386 29795
rect 5340 29747 5406 29759
rect 5340 29713 5356 29747
rect 5390 29713 5406 29747
rect 5340 29679 5406 29713
rect 5340 29645 5356 29679
rect 5390 29645 5406 29679
rect 5340 29633 5406 29645
rect 5440 29747 5486 29763
rect 5474 29713 5486 29747
rect 5440 29679 5486 29713
rect 5474 29645 5486 29679
rect 5061 29578 5095 29612
rect 5440 29599 5486 29645
rect 3873 29468 3907 29544
rect 3971 29532 3987 29566
rect 4021 29532 4037 29566
rect 4163 29532 4179 29566
rect 4213 29532 4229 29566
rect 4355 29532 4371 29566
rect 4405 29532 4421 29566
rect 4547 29532 4563 29566
rect 4597 29532 4613 29566
rect 4739 29532 4755 29566
rect 4789 29532 4805 29566
rect 4931 29532 4947 29566
rect 4981 29532 4997 29566
rect 5274 29565 5303 29599
rect 5337 29565 5395 29599
rect 5429 29565 5487 29599
rect 5521 29565 5550 29599
rect 5061 29468 5095 29541
rect 3873 29434 3991 29468
rect 4025 29434 4059 29468
rect 4093 29434 4127 29468
rect 4161 29434 4195 29468
rect 4229 29434 4263 29468
rect 4297 29434 4331 29468
rect 4365 29434 4399 29468
rect 4433 29434 4467 29468
rect 4501 29434 4535 29468
rect 4569 29434 4603 29468
rect 4637 29434 4671 29468
rect 4705 29434 4739 29468
rect 4773 29434 4807 29468
rect 4841 29434 4875 29468
rect 4909 29434 4943 29468
rect 4977 29434 5095 29468
rect 199 29151 317 29185
rect 351 29151 385 29185
rect 419 29151 453 29185
rect 487 29151 521 29185
rect 555 29151 589 29185
rect 623 29151 657 29185
rect 691 29151 725 29185
rect 759 29151 793 29185
rect 827 29151 861 29185
rect 895 29151 929 29185
rect 963 29151 997 29185
rect 1031 29151 1065 29185
rect 1099 29151 1133 29185
rect 1167 29151 1201 29185
rect 1235 29151 1269 29185
rect 1303 29151 1421 29185
rect 199 29083 233 29151
rect 1387 29083 1421 29151
rect 297 29049 313 29083
rect 347 29049 363 29083
rect 489 29049 505 29083
rect 539 29049 555 29083
rect 681 29049 697 29083
rect 731 29049 747 29083
rect 873 29049 889 29083
rect 923 29049 939 29083
rect 1065 29049 1081 29083
rect 1115 29049 1131 29083
rect 1257 29049 1273 29083
rect 1307 29049 1323 29083
rect 199 29015 233 29049
rect 1387 29015 1421 29023
rect 199 28947 233 28981
rect 199 28879 233 28913
rect 199 28811 233 28845
rect 199 28743 233 28777
rect 313 28984 347 29005
rect 313 28916 347 28920
rect 313 28810 347 28814
rect 313 28725 347 28746
rect 409 28984 443 29005
rect 409 28916 443 28920
rect 409 28810 443 28814
rect 409 28725 443 28746
rect 505 28984 539 29005
rect 505 28916 539 28920
rect 505 28810 539 28814
rect 505 28725 539 28746
rect 601 28984 635 29005
rect 601 28916 635 28920
rect 601 28810 635 28814
rect 601 28725 635 28746
rect 697 28984 731 29005
rect 697 28916 731 28920
rect 697 28810 731 28814
rect 697 28725 731 28746
rect 793 28984 827 29005
rect 793 28916 827 28920
rect 793 28810 827 28814
rect 793 28725 827 28746
rect 889 28984 923 29005
rect 889 28916 923 28920
rect 889 28810 923 28814
rect 889 28725 923 28746
rect 985 28984 1019 29005
rect 985 28916 1019 28920
rect 985 28810 1019 28814
rect 985 28725 1019 28746
rect 1081 28984 1115 29005
rect 1081 28916 1115 28920
rect 1081 28810 1115 28814
rect 1081 28725 1115 28746
rect 1177 28984 1211 29005
rect 1177 28916 1211 28920
rect 1177 28810 1211 28814
rect 1177 28725 1211 28746
rect 1273 28984 1307 29005
rect 1273 28916 1307 28920
rect 1273 28810 1307 28814
rect 1273 28725 1307 28746
rect 1387 28947 1421 28951
rect 1387 28841 1421 28845
rect 1387 28769 1421 28777
rect 199 28641 233 28709
rect 1387 28641 1421 28709
rect 199 28607 317 28641
rect 351 28607 385 28641
rect 419 28607 453 28641
rect 487 28607 521 28641
rect 555 28607 589 28641
rect 623 28607 657 28641
rect 691 28607 725 28641
rect 759 28607 793 28641
rect 827 28607 861 28641
rect 895 28607 929 28641
rect 963 28607 997 28641
rect 1031 28607 1065 28641
rect 1099 28607 1133 28641
rect 1167 28607 1201 28641
rect 1235 28607 1269 28641
rect 1303 28607 1421 28641
rect 2352 29155 2470 29189
rect 2504 29155 2538 29189
rect 2572 29155 2606 29189
rect 2640 29155 2674 29189
rect 2708 29155 2742 29189
rect 2776 29155 2810 29189
rect 2844 29155 2878 29189
rect 2912 29155 2946 29189
rect 2980 29155 3014 29189
rect 3048 29155 3082 29189
rect 3116 29155 3150 29189
rect 3184 29155 3218 29189
rect 3252 29155 3286 29189
rect 3320 29155 3354 29189
rect 3388 29155 3422 29189
rect 3456 29155 3574 29189
rect 2352 29087 2386 29155
rect 3540 29087 3574 29155
rect 2450 29053 2466 29087
rect 2500 29053 2516 29087
rect 2642 29053 2658 29087
rect 2692 29053 2708 29087
rect 2834 29053 2850 29087
rect 2884 29053 2900 29087
rect 3026 29053 3042 29087
rect 3076 29053 3092 29087
rect 3218 29053 3234 29087
rect 3268 29053 3284 29087
rect 3410 29053 3426 29087
rect 3460 29053 3476 29087
rect 2352 29019 2386 29053
rect 3540 29019 3574 29027
rect 2352 28951 2386 28985
rect 2352 28883 2386 28917
rect 2352 28815 2386 28849
rect 2352 28747 2386 28781
rect 2466 28988 2500 29009
rect 2466 28920 2500 28924
rect 2466 28814 2500 28818
rect 2466 28729 2500 28750
rect 2562 28988 2596 29009
rect 2562 28920 2596 28924
rect 2562 28814 2596 28818
rect 2562 28729 2596 28750
rect 2658 28988 2692 29009
rect 2658 28920 2692 28924
rect 2658 28814 2692 28818
rect 2658 28729 2692 28750
rect 2754 28988 2788 29009
rect 2754 28920 2788 28924
rect 2754 28814 2788 28818
rect 2754 28729 2788 28750
rect 2850 28988 2884 29009
rect 2850 28920 2884 28924
rect 2850 28814 2884 28818
rect 2850 28729 2884 28750
rect 2946 28988 2980 29009
rect 2946 28920 2980 28924
rect 2946 28814 2980 28818
rect 2946 28729 2980 28750
rect 3042 28988 3076 29009
rect 3042 28920 3076 28924
rect 3042 28814 3076 28818
rect 3042 28729 3076 28750
rect 3138 28988 3172 29009
rect 3138 28920 3172 28924
rect 3138 28814 3172 28818
rect 3138 28729 3172 28750
rect 3234 28988 3268 29009
rect 3234 28920 3268 28924
rect 3234 28814 3268 28818
rect 3234 28729 3268 28750
rect 3330 28988 3364 29009
rect 3330 28920 3364 28924
rect 3330 28814 3364 28818
rect 3330 28729 3364 28750
rect 3426 28988 3460 29009
rect 3426 28920 3460 28924
rect 3426 28814 3460 28818
rect 3426 28729 3460 28750
rect 3540 28951 3574 28955
rect 3540 28845 3574 28849
rect 3540 28773 3574 28781
rect 2352 28645 2386 28713
rect 3540 28645 3574 28713
rect 2352 28611 2470 28645
rect 2504 28611 2538 28645
rect 2572 28611 2606 28645
rect 2640 28611 2674 28645
rect 2708 28611 2742 28645
rect 2776 28611 2810 28645
rect 2844 28611 2878 28645
rect 2912 28611 2946 28645
rect 2980 28611 3014 28645
rect 3048 28611 3082 28645
rect 3116 28611 3150 28645
rect 3184 28611 3218 28645
rect 3252 28611 3286 28645
rect 3320 28611 3354 28645
rect 3388 28611 3422 28645
rect 3456 28611 3574 28645
rect 3873 29155 3991 29189
rect 4025 29155 4059 29189
rect 4093 29155 4127 29189
rect 4161 29155 4195 29189
rect 4229 29155 4263 29189
rect 4297 29155 4331 29189
rect 4365 29155 4399 29189
rect 4433 29155 4467 29189
rect 4501 29155 4535 29189
rect 4569 29155 4603 29189
rect 4637 29155 4671 29189
rect 4705 29155 4739 29189
rect 4773 29155 4807 29189
rect 4841 29155 4875 29189
rect 4909 29155 4943 29189
rect 4977 29155 5095 29189
rect 3873 29087 3907 29155
rect 5061 29087 5095 29155
rect 3971 29053 3987 29087
rect 4021 29053 4037 29087
rect 4163 29053 4179 29087
rect 4213 29053 4229 29087
rect 4355 29053 4371 29087
rect 4405 29053 4421 29087
rect 4547 29053 4563 29087
rect 4597 29053 4613 29087
rect 4739 29053 4755 29087
rect 4789 29053 4805 29087
rect 4931 29053 4947 29087
rect 4981 29053 4997 29087
rect 3873 29019 3907 29053
rect 5061 29019 5095 29027
rect 3873 28951 3907 28985
rect 3873 28883 3907 28917
rect 3873 28815 3907 28849
rect 3873 28747 3907 28781
rect 3987 28988 4021 29009
rect 3987 28920 4021 28924
rect 3987 28814 4021 28818
rect 3987 28729 4021 28750
rect 4083 28988 4117 29009
rect 4083 28920 4117 28924
rect 4083 28814 4117 28818
rect 4083 28729 4117 28750
rect 4179 28988 4213 29009
rect 4179 28920 4213 28924
rect 4179 28814 4213 28818
rect 4179 28729 4213 28750
rect 4275 28988 4309 29009
rect 4275 28920 4309 28924
rect 4275 28814 4309 28818
rect 4275 28729 4309 28750
rect 4371 28988 4405 29009
rect 4371 28920 4405 28924
rect 4371 28814 4405 28818
rect 4371 28729 4405 28750
rect 4467 28988 4501 29009
rect 4467 28920 4501 28924
rect 4467 28814 4501 28818
rect 4467 28729 4501 28750
rect 4563 28988 4597 29009
rect 4563 28920 4597 28924
rect 4563 28814 4597 28818
rect 4563 28729 4597 28750
rect 4659 28988 4693 29009
rect 4659 28920 4693 28924
rect 4659 28814 4693 28818
rect 4659 28729 4693 28750
rect 4755 28988 4789 29009
rect 4755 28920 4789 28924
rect 4755 28814 4789 28818
rect 4755 28729 4789 28750
rect 4851 28988 4885 29009
rect 4851 28920 4885 28924
rect 4851 28814 4885 28818
rect 4851 28729 4885 28750
rect 4947 28988 4981 29009
rect 4947 28920 4981 28924
rect 4947 28814 4981 28818
rect 4947 28729 4981 28750
rect 5061 28951 5095 28955
rect 5061 28845 5095 28849
rect 5274 28822 5303 28856
rect 5337 28822 5395 28856
rect 5429 28822 5487 28856
rect 5521 28822 5550 28856
rect 5061 28773 5095 28781
rect 3873 28645 3907 28713
rect 5061 28645 5095 28713
rect 3873 28611 3991 28645
rect 4025 28611 4059 28645
rect 4093 28611 4127 28645
rect 4161 28611 4195 28645
rect 4229 28611 4263 28645
rect 4297 28611 4331 28645
rect 4365 28611 4399 28645
rect 4433 28611 4467 28645
rect 4501 28611 4535 28645
rect 4569 28611 4603 28645
rect 4637 28611 4671 28645
rect 4705 28611 4739 28645
rect 4773 28611 4807 28645
rect 4841 28611 4875 28645
rect 4909 28611 4943 28645
rect 4977 28611 5095 28645
rect 5340 28780 5406 28788
rect 5340 28746 5356 28780
rect 5390 28746 5406 28780
rect 5340 28712 5406 28746
rect 5340 28678 5356 28712
rect 5390 28678 5406 28712
rect 5340 28644 5406 28678
rect 5340 28610 5356 28644
rect 5390 28610 5406 28644
rect 5340 28592 5406 28610
rect 5440 28780 5482 28822
rect 5474 28746 5482 28780
rect 5440 28712 5482 28746
rect 5474 28678 5482 28712
rect 5440 28644 5482 28678
rect 5474 28610 5482 28644
rect 5440 28594 5482 28610
rect 5340 28542 5386 28592
rect 199 28499 317 28533
rect 351 28499 385 28533
rect 419 28499 453 28533
rect 487 28499 521 28533
rect 555 28499 589 28533
rect 623 28499 657 28533
rect 691 28499 725 28533
rect 759 28499 793 28533
rect 827 28499 861 28533
rect 895 28499 929 28533
rect 963 28499 997 28533
rect 1031 28499 1065 28533
rect 1099 28499 1133 28533
rect 1167 28499 1201 28533
rect 1235 28499 1269 28533
rect 1303 28499 1421 28533
rect 199 28423 233 28499
rect 1387 28428 1421 28499
rect 199 28355 233 28389
rect 199 28287 233 28321
rect 313 28386 347 28425
rect 313 28313 347 28352
rect 409 28386 443 28425
rect 409 28313 443 28352
rect 505 28386 539 28425
rect 505 28313 539 28352
rect 601 28386 635 28425
rect 601 28313 635 28352
rect 697 28386 731 28425
rect 697 28313 731 28352
rect 793 28386 827 28425
rect 793 28313 827 28352
rect 889 28386 923 28425
rect 889 28313 923 28352
rect 985 28386 1019 28425
rect 985 28313 1019 28352
rect 1081 28386 1115 28425
rect 1081 28313 1115 28352
rect 1177 28386 1211 28425
rect 1177 28313 1211 28352
rect 1273 28386 1307 28425
rect 1273 28313 1307 28352
rect 1387 28356 1421 28389
rect 1387 28287 1421 28321
rect 199 28177 233 28253
rect 297 28241 313 28275
rect 347 28241 363 28275
rect 489 28241 505 28275
rect 539 28241 555 28275
rect 681 28241 697 28275
rect 731 28241 747 28275
rect 873 28241 889 28275
rect 923 28241 939 28275
rect 1065 28241 1081 28275
rect 1115 28241 1131 28275
rect 1257 28241 1273 28275
rect 1307 28241 1323 28275
rect 1387 28177 1421 28250
rect 199 28143 317 28177
rect 351 28143 385 28177
rect 419 28143 453 28177
rect 487 28143 521 28177
rect 555 28143 589 28177
rect 623 28143 657 28177
rect 691 28143 725 28177
rect 759 28143 793 28177
rect 827 28143 861 28177
rect 895 28143 929 28177
rect 963 28143 997 28177
rect 1031 28143 1065 28177
rect 1099 28143 1133 28177
rect 1167 28143 1201 28177
rect 1235 28143 1269 28177
rect 1303 28143 1421 28177
rect 2352 28503 2470 28537
rect 2504 28503 2538 28537
rect 2572 28503 2606 28537
rect 2640 28503 2674 28537
rect 2708 28503 2742 28537
rect 2776 28503 2810 28537
rect 2844 28503 2878 28537
rect 2912 28503 2946 28537
rect 2980 28503 3014 28537
rect 3048 28503 3082 28537
rect 3116 28503 3150 28537
rect 3184 28503 3218 28537
rect 3252 28503 3286 28537
rect 3320 28503 3354 28537
rect 3388 28503 3422 28537
rect 3456 28503 3574 28537
rect 2352 28427 2386 28503
rect 3540 28432 3574 28503
rect 3873 28503 3991 28537
rect 4025 28503 4059 28537
rect 4093 28503 4127 28537
rect 4161 28503 4195 28537
rect 4229 28503 4263 28537
rect 4297 28503 4331 28537
rect 4365 28503 4399 28537
rect 4433 28503 4467 28537
rect 4501 28503 4535 28537
rect 4569 28503 4603 28537
rect 4637 28503 4671 28537
rect 4705 28503 4739 28537
rect 4773 28503 4807 28537
rect 4841 28503 4875 28537
rect 4909 28503 4943 28537
rect 4977 28503 5095 28537
rect 3675 28467 3691 28501
rect 3725 28467 3741 28501
rect 2352 28359 2386 28393
rect 2352 28291 2386 28325
rect 2466 28390 2500 28429
rect 2466 28317 2500 28356
rect 2562 28390 2596 28429
rect 2562 28317 2596 28356
rect 2658 28390 2692 28429
rect 2658 28317 2692 28356
rect 2754 28390 2788 28429
rect 2754 28317 2788 28356
rect 2850 28390 2884 28429
rect 2850 28317 2884 28356
rect 2946 28390 2980 28429
rect 2946 28317 2980 28356
rect 3042 28390 3076 28429
rect 3042 28317 3076 28356
rect 3138 28390 3172 28429
rect 3138 28317 3172 28356
rect 3234 28390 3268 28429
rect 3234 28317 3268 28356
rect 3330 28390 3364 28429
rect 3330 28317 3364 28356
rect 3426 28390 3460 28429
rect 3426 28317 3460 28356
rect 3540 28360 3574 28393
rect 3647 28417 3681 28433
rect 3647 28325 3681 28341
rect 3735 28417 3769 28433
rect 3735 28325 3769 28341
rect 3873 28427 3907 28503
rect 5061 28432 5095 28503
rect 3873 28359 3907 28393
rect 3540 28291 3574 28325
rect 2352 28181 2386 28257
rect 2450 28245 2466 28279
rect 2500 28245 2516 28279
rect 2642 28245 2658 28279
rect 2692 28245 2708 28279
rect 2834 28245 2850 28279
rect 2884 28245 2900 28279
rect 3026 28245 3042 28279
rect 3076 28245 3092 28279
rect 3218 28245 3234 28279
rect 3268 28245 3284 28279
rect 3410 28245 3426 28279
rect 3460 28245 3476 28279
rect 3540 28181 3574 28254
rect 2352 28147 2470 28181
rect 2504 28147 2538 28181
rect 2572 28147 2606 28181
rect 2640 28147 2674 28181
rect 2708 28147 2742 28181
rect 2776 28147 2810 28181
rect 2844 28147 2878 28181
rect 2912 28147 2946 28181
rect 2980 28147 3014 28181
rect 3048 28147 3082 28181
rect 3116 28147 3150 28181
rect 3184 28147 3218 28181
rect 3252 28147 3286 28181
rect 3320 28147 3354 28181
rect 3388 28147 3422 28181
rect 3456 28147 3574 28181
rect 3873 28291 3907 28325
rect 3987 28390 4021 28429
rect 3987 28317 4021 28356
rect 4083 28390 4117 28429
rect 4083 28317 4117 28356
rect 4179 28390 4213 28429
rect 4179 28317 4213 28356
rect 4275 28390 4309 28429
rect 4275 28317 4309 28356
rect 4371 28390 4405 28429
rect 4371 28317 4405 28356
rect 4467 28390 4501 28429
rect 4467 28317 4501 28356
rect 4563 28390 4597 28429
rect 4563 28317 4597 28356
rect 4659 28390 4693 28429
rect 4659 28317 4693 28356
rect 4755 28390 4789 28429
rect 4755 28317 4789 28356
rect 4851 28390 4885 28429
rect 4851 28317 4885 28356
rect 4947 28390 4981 28429
rect 4947 28317 4981 28356
rect 5061 28360 5095 28393
rect 5340 28508 5348 28542
rect 5382 28508 5386 28542
rect 5420 28547 5486 28558
rect 5420 28544 5450 28547
rect 5420 28510 5436 28544
rect 5484 28513 5486 28547
rect 5470 28510 5486 28513
rect 5340 28472 5386 28508
rect 5340 28460 5406 28472
rect 5340 28426 5356 28460
rect 5390 28426 5406 28460
rect 5340 28392 5406 28426
rect 5340 28358 5356 28392
rect 5390 28358 5406 28392
rect 5340 28346 5406 28358
rect 5440 28460 5486 28476
rect 5474 28426 5486 28460
rect 5440 28392 5486 28426
rect 5474 28358 5486 28392
rect 5061 28291 5095 28325
rect 5440 28312 5486 28358
rect 3873 28181 3907 28257
rect 3971 28245 3987 28279
rect 4021 28245 4037 28279
rect 4163 28245 4179 28279
rect 4213 28245 4229 28279
rect 4355 28245 4371 28279
rect 4405 28245 4421 28279
rect 4547 28245 4563 28279
rect 4597 28245 4613 28279
rect 4739 28245 4755 28279
rect 4789 28245 4805 28279
rect 4931 28245 4947 28279
rect 4981 28245 4997 28279
rect 5274 28278 5303 28312
rect 5337 28278 5395 28312
rect 5429 28278 5487 28312
rect 5521 28278 5550 28312
rect 5061 28181 5095 28254
rect 3873 28147 3991 28181
rect 4025 28147 4059 28181
rect 4093 28147 4127 28181
rect 4161 28147 4195 28181
rect 4229 28147 4263 28181
rect 4297 28147 4331 28181
rect 4365 28147 4399 28181
rect 4433 28147 4467 28181
rect 4501 28147 4535 28181
rect 4569 28147 4603 28181
rect 4637 28147 4671 28181
rect 4705 28147 4739 28181
rect 4773 28147 4807 28181
rect 4841 28147 4875 28181
rect 4909 28147 4943 28181
rect 4977 28147 5095 28181
rect 199 27864 317 27898
rect 351 27864 385 27898
rect 419 27864 453 27898
rect 487 27864 521 27898
rect 555 27864 589 27898
rect 623 27864 657 27898
rect 691 27864 725 27898
rect 759 27864 793 27898
rect 827 27864 861 27898
rect 895 27864 929 27898
rect 963 27864 997 27898
rect 1031 27864 1065 27898
rect 1099 27864 1133 27898
rect 1167 27864 1201 27898
rect 1235 27864 1269 27898
rect 1303 27864 1421 27898
rect 199 27796 233 27864
rect 1387 27796 1421 27864
rect 297 27762 313 27796
rect 347 27762 363 27796
rect 489 27762 505 27796
rect 539 27762 555 27796
rect 681 27762 697 27796
rect 731 27762 747 27796
rect 873 27762 889 27796
rect 923 27762 939 27796
rect 1065 27762 1081 27796
rect 1115 27762 1131 27796
rect 1257 27762 1273 27796
rect 1307 27762 1323 27796
rect 199 27728 233 27762
rect 1387 27728 1421 27736
rect 199 27660 233 27694
rect 199 27592 233 27626
rect 199 27524 233 27558
rect 199 27456 233 27490
rect 313 27697 347 27718
rect 313 27629 347 27633
rect 313 27523 347 27527
rect 313 27438 347 27459
rect 409 27697 443 27718
rect 409 27629 443 27633
rect 409 27523 443 27527
rect 409 27438 443 27459
rect 505 27697 539 27718
rect 505 27629 539 27633
rect 505 27523 539 27527
rect 505 27438 539 27459
rect 601 27697 635 27718
rect 601 27629 635 27633
rect 601 27523 635 27527
rect 601 27438 635 27459
rect 697 27697 731 27718
rect 697 27629 731 27633
rect 697 27523 731 27527
rect 697 27438 731 27459
rect 793 27697 827 27718
rect 793 27629 827 27633
rect 793 27523 827 27527
rect 793 27438 827 27459
rect 889 27697 923 27718
rect 889 27629 923 27633
rect 889 27523 923 27527
rect 889 27438 923 27459
rect 985 27697 1019 27718
rect 985 27629 1019 27633
rect 985 27523 1019 27527
rect 985 27438 1019 27459
rect 1081 27697 1115 27718
rect 1081 27629 1115 27633
rect 1081 27523 1115 27527
rect 1081 27438 1115 27459
rect 1177 27697 1211 27718
rect 1177 27629 1211 27633
rect 1177 27523 1211 27527
rect 1177 27438 1211 27459
rect 1273 27697 1307 27718
rect 1273 27629 1307 27633
rect 1273 27523 1307 27527
rect 1273 27438 1307 27459
rect 1387 27660 1421 27664
rect 1387 27554 1421 27558
rect 1387 27482 1421 27490
rect 199 27354 233 27422
rect 1387 27354 1421 27422
rect 199 27320 317 27354
rect 351 27320 385 27354
rect 419 27320 453 27354
rect 487 27320 521 27354
rect 555 27320 589 27354
rect 623 27320 657 27354
rect 691 27320 725 27354
rect 759 27320 793 27354
rect 827 27320 861 27354
rect 895 27320 929 27354
rect 963 27320 997 27354
rect 1031 27320 1065 27354
rect 1099 27320 1133 27354
rect 1167 27320 1201 27354
rect 1235 27320 1269 27354
rect 1303 27320 1421 27354
rect 2352 27868 2470 27902
rect 2504 27868 2538 27902
rect 2572 27868 2606 27902
rect 2640 27868 2674 27902
rect 2708 27868 2742 27902
rect 2776 27868 2810 27902
rect 2844 27868 2878 27902
rect 2912 27868 2946 27902
rect 2980 27868 3014 27902
rect 3048 27868 3082 27902
rect 3116 27868 3150 27902
rect 3184 27868 3218 27902
rect 3252 27868 3286 27902
rect 3320 27868 3354 27902
rect 3388 27868 3422 27902
rect 3456 27868 3574 27902
rect 2352 27800 2386 27868
rect 3540 27800 3574 27868
rect 2450 27766 2466 27800
rect 2500 27766 2516 27800
rect 2642 27766 2658 27800
rect 2692 27766 2708 27800
rect 2834 27766 2850 27800
rect 2884 27766 2900 27800
rect 3026 27766 3042 27800
rect 3076 27766 3092 27800
rect 3218 27766 3234 27800
rect 3268 27766 3284 27800
rect 3410 27766 3426 27800
rect 3460 27766 3476 27800
rect 2352 27732 2386 27766
rect 3540 27732 3574 27740
rect 2352 27664 2386 27698
rect 2352 27596 2386 27630
rect 2352 27528 2386 27562
rect 2352 27460 2386 27494
rect 2466 27701 2500 27722
rect 2466 27633 2500 27637
rect 2466 27527 2500 27531
rect 2466 27442 2500 27463
rect 2562 27701 2596 27722
rect 2562 27633 2596 27637
rect 2562 27527 2596 27531
rect 2562 27442 2596 27463
rect 2658 27701 2692 27722
rect 2658 27633 2692 27637
rect 2658 27527 2692 27531
rect 2658 27442 2692 27463
rect 2754 27701 2788 27722
rect 2754 27633 2788 27637
rect 2754 27527 2788 27531
rect 2754 27442 2788 27463
rect 2850 27701 2884 27722
rect 2850 27633 2884 27637
rect 2850 27527 2884 27531
rect 2850 27442 2884 27463
rect 2946 27701 2980 27722
rect 2946 27633 2980 27637
rect 2946 27527 2980 27531
rect 2946 27442 2980 27463
rect 3042 27701 3076 27722
rect 3042 27633 3076 27637
rect 3042 27527 3076 27531
rect 3042 27442 3076 27463
rect 3138 27701 3172 27722
rect 3138 27633 3172 27637
rect 3138 27527 3172 27531
rect 3138 27442 3172 27463
rect 3234 27701 3268 27722
rect 3234 27633 3268 27637
rect 3234 27527 3268 27531
rect 3234 27442 3268 27463
rect 3330 27701 3364 27722
rect 3330 27633 3364 27637
rect 3330 27527 3364 27531
rect 3330 27442 3364 27463
rect 3426 27701 3460 27722
rect 3426 27633 3460 27637
rect 3426 27527 3460 27531
rect 3426 27442 3460 27463
rect 3540 27664 3574 27668
rect 3540 27558 3574 27562
rect 3540 27486 3574 27494
rect 2352 27358 2386 27426
rect 3540 27358 3574 27426
rect 2352 27324 2470 27358
rect 2504 27324 2538 27358
rect 2572 27324 2606 27358
rect 2640 27324 2674 27358
rect 2708 27324 2742 27358
rect 2776 27324 2810 27358
rect 2844 27324 2878 27358
rect 2912 27324 2946 27358
rect 2980 27324 3014 27358
rect 3048 27324 3082 27358
rect 3116 27324 3150 27358
rect 3184 27324 3218 27358
rect 3252 27324 3286 27358
rect 3320 27324 3354 27358
rect 3388 27324 3422 27358
rect 3456 27324 3574 27358
rect 3873 27868 3991 27902
rect 4025 27868 4059 27902
rect 4093 27868 4127 27902
rect 4161 27868 4195 27902
rect 4229 27868 4263 27902
rect 4297 27868 4331 27902
rect 4365 27868 4399 27902
rect 4433 27868 4467 27902
rect 4501 27868 4535 27902
rect 4569 27868 4603 27902
rect 4637 27868 4671 27902
rect 4705 27868 4739 27902
rect 4773 27868 4807 27902
rect 4841 27868 4875 27902
rect 4909 27868 4943 27902
rect 4977 27868 5095 27902
rect 3873 27800 3907 27868
rect 5061 27800 5095 27868
rect 3971 27766 3987 27800
rect 4021 27766 4037 27800
rect 4163 27766 4179 27800
rect 4213 27766 4229 27800
rect 4355 27766 4371 27800
rect 4405 27766 4421 27800
rect 4547 27766 4563 27800
rect 4597 27766 4613 27800
rect 4739 27766 4755 27800
rect 4789 27766 4805 27800
rect 4931 27766 4947 27800
rect 4981 27766 4997 27800
rect 3873 27732 3907 27766
rect 5061 27732 5095 27740
rect 3873 27664 3907 27698
rect 3873 27596 3907 27630
rect 3873 27528 3907 27562
rect 3873 27460 3907 27494
rect 3987 27701 4021 27722
rect 3987 27633 4021 27637
rect 3987 27527 4021 27531
rect 3987 27442 4021 27463
rect 4083 27701 4117 27722
rect 4083 27633 4117 27637
rect 4083 27527 4117 27531
rect 4083 27442 4117 27463
rect 4179 27701 4213 27722
rect 4179 27633 4213 27637
rect 4179 27527 4213 27531
rect 4179 27442 4213 27463
rect 4275 27701 4309 27722
rect 4275 27633 4309 27637
rect 4275 27527 4309 27531
rect 4275 27442 4309 27463
rect 4371 27701 4405 27722
rect 4371 27633 4405 27637
rect 4371 27527 4405 27531
rect 4371 27442 4405 27463
rect 4467 27701 4501 27722
rect 4467 27633 4501 27637
rect 4467 27527 4501 27531
rect 4467 27442 4501 27463
rect 4563 27701 4597 27722
rect 4563 27633 4597 27637
rect 4563 27527 4597 27531
rect 4563 27442 4597 27463
rect 4659 27701 4693 27722
rect 4659 27633 4693 27637
rect 4659 27527 4693 27531
rect 4659 27442 4693 27463
rect 4755 27701 4789 27722
rect 4755 27633 4789 27637
rect 4755 27527 4789 27531
rect 4755 27442 4789 27463
rect 4851 27701 4885 27722
rect 4851 27633 4885 27637
rect 4851 27527 4885 27531
rect 4851 27442 4885 27463
rect 4947 27701 4981 27722
rect 4947 27633 4981 27637
rect 4947 27527 4981 27531
rect 4947 27442 4981 27463
rect 5061 27664 5095 27668
rect 5061 27558 5095 27562
rect 5274 27535 5303 27569
rect 5337 27535 5395 27569
rect 5429 27535 5487 27569
rect 5521 27535 5550 27569
rect 5061 27486 5095 27494
rect 3873 27358 3907 27426
rect 5061 27358 5095 27426
rect 3873 27324 3991 27358
rect 4025 27324 4059 27358
rect 4093 27324 4127 27358
rect 4161 27324 4195 27358
rect 4229 27324 4263 27358
rect 4297 27324 4331 27358
rect 4365 27324 4399 27358
rect 4433 27324 4467 27358
rect 4501 27324 4535 27358
rect 4569 27324 4603 27358
rect 4637 27324 4671 27358
rect 4705 27324 4739 27358
rect 4773 27324 4807 27358
rect 4841 27324 4875 27358
rect 4909 27324 4943 27358
rect 4977 27324 5095 27358
rect 5340 27493 5406 27501
rect 5340 27459 5356 27493
rect 5390 27459 5406 27493
rect 5340 27425 5406 27459
rect 5340 27391 5356 27425
rect 5390 27391 5406 27425
rect 5340 27357 5406 27391
rect 5340 27323 5356 27357
rect 5390 27323 5406 27357
rect 5340 27305 5406 27323
rect 5440 27493 5482 27535
rect 5474 27459 5482 27493
rect 5440 27425 5482 27459
rect 5474 27391 5482 27425
rect 5440 27357 5482 27391
rect 5474 27323 5482 27357
rect 5440 27307 5482 27323
rect 5340 27255 5386 27305
rect 199 27212 317 27246
rect 351 27212 385 27246
rect 419 27212 453 27246
rect 487 27212 521 27246
rect 555 27212 589 27246
rect 623 27212 657 27246
rect 691 27212 725 27246
rect 759 27212 793 27246
rect 827 27212 861 27246
rect 895 27212 929 27246
rect 963 27212 997 27246
rect 1031 27212 1065 27246
rect 1099 27212 1133 27246
rect 1167 27212 1201 27246
rect 1235 27212 1269 27246
rect 1303 27212 1421 27246
rect 199 27136 233 27212
rect 1387 27141 1421 27212
rect 199 27068 233 27102
rect 199 27000 233 27034
rect 313 27099 347 27138
rect 313 27026 347 27065
rect 409 27099 443 27138
rect 409 27026 443 27065
rect 505 27099 539 27138
rect 505 27026 539 27065
rect 601 27099 635 27138
rect 601 27026 635 27065
rect 697 27099 731 27138
rect 697 27026 731 27065
rect 793 27099 827 27138
rect 793 27026 827 27065
rect 889 27099 923 27138
rect 889 27026 923 27065
rect 985 27099 1019 27138
rect 985 27026 1019 27065
rect 1081 27099 1115 27138
rect 1081 27026 1115 27065
rect 1177 27099 1211 27138
rect 1177 27026 1211 27065
rect 1273 27099 1307 27138
rect 1273 27026 1307 27065
rect 1387 27069 1421 27102
rect 1387 27000 1421 27034
rect 199 26890 233 26966
rect 297 26954 313 26988
rect 347 26954 363 26988
rect 489 26954 505 26988
rect 539 26954 555 26988
rect 681 26954 697 26988
rect 731 26954 747 26988
rect 873 26954 889 26988
rect 923 26954 939 26988
rect 1065 26954 1081 26988
rect 1115 26954 1131 26988
rect 1257 26954 1273 26988
rect 1307 26954 1323 26988
rect 1387 26890 1421 26963
rect 199 26856 317 26890
rect 351 26856 385 26890
rect 419 26856 453 26890
rect 487 26856 521 26890
rect 555 26856 589 26890
rect 623 26856 657 26890
rect 691 26856 725 26890
rect 759 26856 793 26890
rect 827 26856 861 26890
rect 895 26856 929 26890
rect 963 26856 997 26890
rect 1031 26856 1065 26890
rect 1099 26856 1133 26890
rect 1167 26856 1201 26890
rect 1235 26856 1269 26890
rect 1303 26856 1421 26890
rect 2352 27216 2470 27250
rect 2504 27216 2538 27250
rect 2572 27216 2606 27250
rect 2640 27216 2674 27250
rect 2708 27216 2742 27250
rect 2776 27216 2810 27250
rect 2844 27216 2878 27250
rect 2912 27216 2946 27250
rect 2980 27216 3014 27250
rect 3048 27216 3082 27250
rect 3116 27216 3150 27250
rect 3184 27216 3218 27250
rect 3252 27216 3286 27250
rect 3320 27216 3354 27250
rect 3388 27216 3422 27250
rect 3456 27216 3574 27250
rect 2352 27140 2386 27216
rect 3540 27145 3574 27216
rect 3873 27216 3991 27250
rect 4025 27216 4059 27250
rect 4093 27216 4127 27250
rect 4161 27216 4195 27250
rect 4229 27216 4263 27250
rect 4297 27216 4331 27250
rect 4365 27216 4399 27250
rect 4433 27216 4467 27250
rect 4501 27216 4535 27250
rect 4569 27216 4603 27250
rect 4637 27216 4671 27250
rect 4705 27216 4739 27250
rect 4773 27216 4807 27250
rect 4841 27216 4875 27250
rect 4909 27216 4943 27250
rect 4977 27216 5095 27250
rect 3675 27180 3691 27214
rect 3725 27180 3741 27214
rect 2352 27072 2386 27106
rect 2352 27004 2386 27038
rect 2466 27103 2500 27142
rect 2466 27030 2500 27069
rect 2562 27103 2596 27142
rect 2562 27030 2596 27069
rect 2658 27103 2692 27142
rect 2658 27030 2692 27069
rect 2754 27103 2788 27142
rect 2754 27030 2788 27069
rect 2850 27103 2884 27142
rect 2850 27030 2884 27069
rect 2946 27103 2980 27142
rect 2946 27030 2980 27069
rect 3042 27103 3076 27142
rect 3042 27030 3076 27069
rect 3138 27103 3172 27142
rect 3138 27030 3172 27069
rect 3234 27103 3268 27142
rect 3234 27030 3268 27069
rect 3330 27103 3364 27142
rect 3330 27030 3364 27069
rect 3426 27103 3460 27142
rect 3426 27030 3460 27069
rect 3540 27073 3574 27106
rect 3647 27130 3681 27146
rect 3647 27038 3681 27054
rect 3735 27130 3769 27146
rect 3735 27038 3769 27054
rect 3873 27140 3907 27216
rect 5061 27145 5095 27216
rect 3873 27072 3907 27106
rect 3540 27004 3574 27038
rect 2352 26894 2386 26970
rect 2450 26958 2466 26992
rect 2500 26958 2516 26992
rect 2642 26958 2658 26992
rect 2692 26958 2708 26992
rect 2834 26958 2850 26992
rect 2884 26958 2900 26992
rect 3026 26958 3042 26992
rect 3076 26958 3092 26992
rect 3218 26958 3234 26992
rect 3268 26958 3284 26992
rect 3410 26958 3426 26992
rect 3460 26958 3476 26992
rect 3540 26894 3574 26967
rect 2352 26860 2470 26894
rect 2504 26860 2538 26894
rect 2572 26860 2606 26894
rect 2640 26860 2674 26894
rect 2708 26860 2742 26894
rect 2776 26860 2810 26894
rect 2844 26860 2878 26894
rect 2912 26860 2946 26894
rect 2980 26860 3014 26894
rect 3048 26860 3082 26894
rect 3116 26860 3150 26894
rect 3184 26860 3218 26894
rect 3252 26860 3286 26894
rect 3320 26860 3354 26894
rect 3388 26860 3422 26894
rect 3456 26860 3574 26894
rect 3873 27004 3907 27038
rect 3987 27103 4021 27142
rect 3987 27030 4021 27069
rect 4083 27103 4117 27142
rect 4083 27030 4117 27069
rect 4179 27103 4213 27142
rect 4179 27030 4213 27069
rect 4275 27103 4309 27142
rect 4275 27030 4309 27069
rect 4371 27103 4405 27142
rect 4371 27030 4405 27069
rect 4467 27103 4501 27142
rect 4467 27030 4501 27069
rect 4563 27103 4597 27142
rect 4563 27030 4597 27069
rect 4659 27103 4693 27142
rect 4659 27030 4693 27069
rect 4755 27103 4789 27142
rect 4755 27030 4789 27069
rect 4851 27103 4885 27142
rect 4851 27030 4885 27069
rect 4947 27103 4981 27142
rect 4947 27030 4981 27069
rect 5061 27073 5095 27106
rect 5340 27221 5348 27255
rect 5382 27221 5386 27255
rect 5420 27260 5486 27271
rect 5420 27257 5450 27260
rect 5420 27223 5436 27257
rect 5484 27226 5486 27260
rect 5470 27223 5486 27226
rect 5340 27185 5386 27221
rect 5340 27173 5406 27185
rect 5340 27139 5356 27173
rect 5390 27139 5406 27173
rect 5340 27105 5406 27139
rect 5340 27071 5356 27105
rect 5390 27071 5406 27105
rect 5340 27059 5406 27071
rect 5440 27173 5486 27189
rect 5474 27139 5486 27173
rect 5440 27105 5486 27139
rect 5474 27071 5486 27105
rect 5061 27004 5095 27038
rect 5440 27025 5486 27071
rect 3873 26894 3907 26970
rect 3971 26958 3987 26992
rect 4021 26958 4037 26992
rect 4163 26958 4179 26992
rect 4213 26958 4229 26992
rect 4355 26958 4371 26992
rect 4405 26958 4421 26992
rect 4547 26958 4563 26992
rect 4597 26958 4613 26992
rect 4739 26958 4755 26992
rect 4789 26958 4805 26992
rect 4931 26958 4947 26992
rect 4981 26958 4997 26992
rect 5274 26991 5303 27025
rect 5337 26991 5395 27025
rect 5429 26991 5487 27025
rect 5521 26991 5550 27025
rect 5061 26894 5095 26967
rect 3873 26860 3991 26894
rect 4025 26860 4059 26894
rect 4093 26860 4127 26894
rect 4161 26860 4195 26894
rect 4229 26860 4263 26894
rect 4297 26860 4331 26894
rect 4365 26860 4399 26894
rect 4433 26860 4467 26894
rect 4501 26860 4535 26894
rect 4569 26860 4603 26894
rect 4637 26860 4671 26894
rect 4705 26860 4739 26894
rect 4773 26860 4807 26894
rect 4841 26860 4875 26894
rect 4909 26860 4943 26894
rect 4977 26860 5095 26894
rect 199 26577 317 26611
rect 351 26577 385 26611
rect 419 26577 453 26611
rect 487 26577 521 26611
rect 555 26577 589 26611
rect 623 26577 657 26611
rect 691 26577 725 26611
rect 759 26577 793 26611
rect 827 26577 861 26611
rect 895 26577 929 26611
rect 963 26577 997 26611
rect 1031 26577 1065 26611
rect 1099 26577 1133 26611
rect 1167 26577 1201 26611
rect 1235 26577 1269 26611
rect 1303 26577 1421 26611
rect 199 26509 233 26577
rect 1387 26509 1421 26577
rect 297 26475 313 26509
rect 347 26475 363 26509
rect 489 26475 505 26509
rect 539 26475 555 26509
rect 681 26475 697 26509
rect 731 26475 747 26509
rect 873 26475 889 26509
rect 923 26475 939 26509
rect 1065 26475 1081 26509
rect 1115 26475 1131 26509
rect 1257 26475 1273 26509
rect 1307 26475 1323 26509
rect 199 26441 233 26475
rect 1387 26441 1421 26449
rect 199 26373 233 26407
rect 199 26305 233 26339
rect 199 26237 233 26271
rect 199 26169 233 26203
rect 313 26410 347 26431
rect 313 26342 347 26346
rect 313 26236 347 26240
rect 313 26151 347 26172
rect 409 26410 443 26431
rect 409 26342 443 26346
rect 409 26236 443 26240
rect 409 26151 443 26172
rect 505 26410 539 26431
rect 505 26342 539 26346
rect 505 26236 539 26240
rect 505 26151 539 26172
rect 601 26410 635 26431
rect 601 26342 635 26346
rect 601 26236 635 26240
rect 601 26151 635 26172
rect 697 26410 731 26431
rect 697 26342 731 26346
rect 697 26236 731 26240
rect 697 26151 731 26172
rect 793 26410 827 26431
rect 793 26342 827 26346
rect 793 26236 827 26240
rect 793 26151 827 26172
rect 889 26410 923 26431
rect 889 26342 923 26346
rect 889 26236 923 26240
rect 889 26151 923 26172
rect 985 26410 1019 26431
rect 985 26342 1019 26346
rect 985 26236 1019 26240
rect 985 26151 1019 26172
rect 1081 26410 1115 26431
rect 1081 26342 1115 26346
rect 1081 26236 1115 26240
rect 1081 26151 1115 26172
rect 1177 26410 1211 26431
rect 1177 26342 1211 26346
rect 1177 26236 1211 26240
rect 1177 26151 1211 26172
rect 1273 26410 1307 26431
rect 1273 26342 1307 26346
rect 1273 26236 1307 26240
rect 1273 26151 1307 26172
rect 1387 26373 1421 26377
rect 1387 26267 1421 26271
rect 1387 26195 1421 26203
rect 199 26067 233 26135
rect 1387 26067 1421 26135
rect 199 26033 317 26067
rect 351 26033 385 26067
rect 419 26033 453 26067
rect 487 26033 521 26067
rect 555 26033 589 26067
rect 623 26033 657 26067
rect 691 26033 725 26067
rect 759 26033 793 26067
rect 827 26033 861 26067
rect 895 26033 929 26067
rect 963 26033 997 26067
rect 1031 26033 1065 26067
rect 1099 26033 1133 26067
rect 1167 26033 1201 26067
rect 1235 26033 1269 26067
rect 1303 26033 1421 26067
rect 2352 26581 2470 26615
rect 2504 26581 2538 26615
rect 2572 26581 2606 26615
rect 2640 26581 2674 26615
rect 2708 26581 2742 26615
rect 2776 26581 2810 26615
rect 2844 26581 2878 26615
rect 2912 26581 2946 26615
rect 2980 26581 3014 26615
rect 3048 26581 3082 26615
rect 3116 26581 3150 26615
rect 3184 26581 3218 26615
rect 3252 26581 3286 26615
rect 3320 26581 3354 26615
rect 3388 26581 3422 26615
rect 3456 26581 3574 26615
rect 2352 26513 2386 26581
rect 3540 26513 3574 26581
rect 2450 26479 2466 26513
rect 2500 26479 2516 26513
rect 2642 26479 2658 26513
rect 2692 26479 2708 26513
rect 2834 26479 2850 26513
rect 2884 26479 2900 26513
rect 3026 26479 3042 26513
rect 3076 26479 3092 26513
rect 3218 26479 3234 26513
rect 3268 26479 3284 26513
rect 3410 26479 3426 26513
rect 3460 26479 3476 26513
rect 2352 26445 2386 26479
rect 3540 26445 3574 26453
rect 2352 26377 2386 26411
rect 2352 26309 2386 26343
rect 2352 26241 2386 26275
rect 2352 26173 2386 26207
rect 2466 26414 2500 26435
rect 2466 26346 2500 26350
rect 2466 26240 2500 26244
rect 2466 26155 2500 26176
rect 2562 26414 2596 26435
rect 2562 26346 2596 26350
rect 2562 26240 2596 26244
rect 2562 26155 2596 26176
rect 2658 26414 2692 26435
rect 2658 26346 2692 26350
rect 2658 26240 2692 26244
rect 2658 26155 2692 26176
rect 2754 26414 2788 26435
rect 2754 26346 2788 26350
rect 2754 26240 2788 26244
rect 2754 26155 2788 26176
rect 2850 26414 2884 26435
rect 2850 26346 2884 26350
rect 2850 26240 2884 26244
rect 2850 26155 2884 26176
rect 2946 26414 2980 26435
rect 2946 26346 2980 26350
rect 2946 26240 2980 26244
rect 2946 26155 2980 26176
rect 3042 26414 3076 26435
rect 3042 26346 3076 26350
rect 3042 26240 3076 26244
rect 3042 26155 3076 26176
rect 3138 26414 3172 26435
rect 3138 26346 3172 26350
rect 3138 26240 3172 26244
rect 3138 26155 3172 26176
rect 3234 26414 3268 26435
rect 3234 26346 3268 26350
rect 3234 26240 3268 26244
rect 3234 26155 3268 26176
rect 3330 26414 3364 26435
rect 3330 26346 3364 26350
rect 3330 26240 3364 26244
rect 3330 26155 3364 26176
rect 3426 26414 3460 26435
rect 3426 26346 3460 26350
rect 3426 26240 3460 26244
rect 3426 26155 3460 26176
rect 3540 26377 3574 26381
rect 3540 26271 3574 26275
rect 3540 26199 3574 26207
rect 2352 26071 2386 26139
rect 3540 26071 3574 26139
rect 2352 26037 2470 26071
rect 2504 26037 2538 26071
rect 2572 26037 2606 26071
rect 2640 26037 2674 26071
rect 2708 26037 2742 26071
rect 2776 26037 2810 26071
rect 2844 26037 2878 26071
rect 2912 26037 2946 26071
rect 2980 26037 3014 26071
rect 3048 26037 3082 26071
rect 3116 26037 3150 26071
rect 3184 26037 3218 26071
rect 3252 26037 3286 26071
rect 3320 26037 3354 26071
rect 3388 26037 3422 26071
rect 3456 26037 3574 26071
rect 3873 26581 3991 26615
rect 4025 26581 4059 26615
rect 4093 26581 4127 26615
rect 4161 26581 4195 26615
rect 4229 26581 4263 26615
rect 4297 26581 4331 26615
rect 4365 26581 4399 26615
rect 4433 26581 4467 26615
rect 4501 26581 4535 26615
rect 4569 26581 4603 26615
rect 4637 26581 4671 26615
rect 4705 26581 4739 26615
rect 4773 26581 4807 26615
rect 4841 26581 4875 26615
rect 4909 26581 4943 26615
rect 4977 26581 5095 26615
rect 3873 26513 3907 26581
rect 5061 26513 5095 26581
rect 3971 26479 3987 26513
rect 4021 26479 4037 26513
rect 4163 26479 4179 26513
rect 4213 26479 4229 26513
rect 4355 26479 4371 26513
rect 4405 26479 4421 26513
rect 4547 26479 4563 26513
rect 4597 26479 4613 26513
rect 4739 26479 4755 26513
rect 4789 26479 4805 26513
rect 4931 26479 4947 26513
rect 4981 26479 4997 26513
rect 3873 26445 3907 26479
rect 5061 26445 5095 26453
rect 3873 26377 3907 26411
rect 3873 26309 3907 26343
rect 3873 26241 3907 26275
rect 3873 26173 3907 26207
rect 3987 26414 4021 26435
rect 3987 26346 4021 26350
rect 3987 26240 4021 26244
rect 3987 26155 4021 26176
rect 4083 26414 4117 26435
rect 4083 26346 4117 26350
rect 4083 26240 4117 26244
rect 4083 26155 4117 26176
rect 4179 26414 4213 26435
rect 4179 26346 4213 26350
rect 4179 26240 4213 26244
rect 4179 26155 4213 26176
rect 4275 26414 4309 26435
rect 4275 26346 4309 26350
rect 4275 26240 4309 26244
rect 4275 26155 4309 26176
rect 4371 26414 4405 26435
rect 4371 26346 4405 26350
rect 4371 26240 4405 26244
rect 4371 26155 4405 26176
rect 4467 26414 4501 26435
rect 4467 26346 4501 26350
rect 4467 26240 4501 26244
rect 4467 26155 4501 26176
rect 4563 26414 4597 26435
rect 4563 26346 4597 26350
rect 4563 26240 4597 26244
rect 4563 26155 4597 26176
rect 4659 26414 4693 26435
rect 4659 26346 4693 26350
rect 4659 26240 4693 26244
rect 4659 26155 4693 26176
rect 4755 26414 4789 26435
rect 4755 26346 4789 26350
rect 4755 26240 4789 26244
rect 4755 26155 4789 26176
rect 4851 26414 4885 26435
rect 4851 26346 4885 26350
rect 4851 26240 4885 26244
rect 4851 26155 4885 26176
rect 4947 26414 4981 26435
rect 4947 26346 4981 26350
rect 4947 26240 4981 26244
rect 4947 26155 4981 26176
rect 5061 26377 5095 26381
rect 5061 26271 5095 26275
rect 5274 26248 5303 26282
rect 5337 26248 5395 26282
rect 5429 26248 5487 26282
rect 5521 26248 5550 26282
rect 5061 26199 5095 26207
rect 3873 26071 3907 26139
rect 5061 26071 5095 26139
rect 3873 26037 3991 26071
rect 4025 26037 4059 26071
rect 4093 26037 4127 26071
rect 4161 26037 4195 26071
rect 4229 26037 4263 26071
rect 4297 26037 4331 26071
rect 4365 26037 4399 26071
rect 4433 26037 4467 26071
rect 4501 26037 4535 26071
rect 4569 26037 4603 26071
rect 4637 26037 4671 26071
rect 4705 26037 4739 26071
rect 4773 26037 4807 26071
rect 4841 26037 4875 26071
rect 4909 26037 4943 26071
rect 4977 26037 5095 26071
rect 5340 26206 5406 26214
rect 5340 26172 5356 26206
rect 5390 26172 5406 26206
rect 5340 26138 5406 26172
rect 5340 26104 5356 26138
rect 5390 26104 5406 26138
rect 5340 26070 5406 26104
rect 5340 26036 5356 26070
rect 5390 26036 5406 26070
rect 5340 26018 5406 26036
rect 5440 26206 5482 26248
rect 5474 26172 5482 26206
rect 5440 26138 5482 26172
rect 5474 26104 5482 26138
rect 5440 26070 5482 26104
rect 5474 26036 5482 26070
rect 5440 26020 5482 26036
rect 5340 25968 5386 26018
rect 199 25925 317 25959
rect 351 25925 385 25959
rect 419 25925 453 25959
rect 487 25925 521 25959
rect 555 25925 589 25959
rect 623 25925 657 25959
rect 691 25925 725 25959
rect 759 25925 793 25959
rect 827 25925 861 25959
rect 895 25925 929 25959
rect 963 25925 997 25959
rect 1031 25925 1065 25959
rect 1099 25925 1133 25959
rect 1167 25925 1201 25959
rect 1235 25925 1269 25959
rect 1303 25925 1421 25959
rect 199 25849 233 25925
rect 1387 25854 1421 25925
rect 199 25781 233 25815
rect 199 25713 233 25747
rect 313 25812 347 25851
rect 313 25739 347 25778
rect 409 25812 443 25851
rect 409 25739 443 25778
rect 505 25812 539 25851
rect 505 25739 539 25778
rect 601 25812 635 25851
rect 601 25739 635 25778
rect 697 25812 731 25851
rect 697 25739 731 25778
rect 793 25812 827 25851
rect 793 25739 827 25778
rect 889 25812 923 25851
rect 889 25739 923 25778
rect 985 25812 1019 25851
rect 985 25739 1019 25778
rect 1081 25812 1115 25851
rect 1081 25739 1115 25778
rect 1177 25812 1211 25851
rect 1177 25739 1211 25778
rect 1273 25812 1307 25851
rect 1273 25739 1307 25778
rect 1387 25782 1421 25815
rect 1387 25713 1421 25747
rect 199 25603 233 25679
rect 297 25667 313 25701
rect 347 25667 363 25701
rect 489 25667 505 25701
rect 539 25667 555 25701
rect 681 25667 697 25701
rect 731 25667 747 25701
rect 873 25667 889 25701
rect 923 25667 939 25701
rect 1065 25667 1081 25701
rect 1115 25667 1131 25701
rect 1257 25667 1273 25701
rect 1307 25667 1323 25701
rect 1387 25603 1421 25676
rect 199 25569 317 25603
rect 351 25569 385 25603
rect 419 25569 453 25603
rect 487 25569 521 25603
rect 555 25569 589 25603
rect 623 25569 657 25603
rect 691 25569 725 25603
rect 759 25569 793 25603
rect 827 25569 861 25603
rect 895 25569 929 25603
rect 963 25569 997 25603
rect 1031 25569 1065 25603
rect 1099 25569 1133 25603
rect 1167 25569 1201 25603
rect 1235 25569 1269 25603
rect 1303 25569 1421 25603
rect 2352 25929 2470 25963
rect 2504 25929 2538 25963
rect 2572 25929 2606 25963
rect 2640 25929 2674 25963
rect 2708 25929 2742 25963
rect 2776 25929 2810 25963
rect 2844 25929 2878 25963
rect 2912 25929 2946 25963
rect 2980 25929 3014 25963
rect 3048 25929 3082 25963
rect 3116 25929 3150 25963
rect 3184 25929 3218 25963
rect 3252 25929 3286 25963
rect 3320 25929 3354 25963
rect 3388 25929 3422 25963
rect 3456 25929 3574 25963
rect 2352 25853 2386 25929
rect 3540 25858 3574 25929
rect 3873 25929 3991 25963
rect 4025 25929 4059 25963
rect 4093 25929 4127 25963
rect 4161 25929 4195 25963
rect 4229 25929 4263 25963
rect 4297 25929 4331 25963
rect 4365 25929 4399 25963
rect 4433 25929 4467 25963
rect 4501 25929 4535 25963
rect 4569 25929 4603 25963
rect 4637 25929 4671 25963
rect 4705 25929 4739 25963
rect 4773 25929 4807 25963
rect 4841 25929 4875 25963
rect 4909 25929 4943 25963
rect 4977 25929 5095 25963
rect 3675 25893 3691 25927
rect 3725 25893 3741 25927
rect 2352 25785 2386 25819
rect 2352 25717 2386 25751
rect 2466 25816 2500 25855
rect 2466 25743 2500 25782
rect 2562 25816 2596 25855
rect 2562 25743 2596 25782
rect 2658 25816 2692 25855
rect 2658 25743 2692 25782
rect 2754 25816 2788 25855
rect 2754 25743 2788 25782
rect 2850 25816 2884 25855
rect 2850 25743 2884 25782
rect 2946 25816 2980 25855
rect 2946 25743 2980 25782
rect 3042 25816 3076 25855
rect 3042 25743 3076 25782
rect 3138 25816 3172 25855
rect 3138 25743 3172 25782
rect 3234 25816 3268 25855
rect 3234 25743 3268 25782
rect 3330 25816 3364 25855
rect 3330 25743 3364 25782
rect 3426 25816 3460 25855
rect 3426 25743 3460 25782
rect 3540 25786 3574 25819
rect 3647 25843 3681 25859
rect 3647 25751 3681 25767
rect 3735 25843 3769 25859
rect 3735 25751 3769 25767
rect 3873 25853 3907 25929
rect 5061 25858 5095 25929
rect 3873 25785 3907 25819
rect 3540 25717 3574 25751
rect 2352 25607 2386 25683
rect 2450 25671 2466 25705
rect 2500 25671 2516 25705
rect 2642 25671 2658 25705
rect 2692 25671 2708 25705
rect 2834 25671 2850 25705
rect 2884 25671 2900 25705
rect 3026 25671 3042 25705
rect 3076 25671 3092 25705
rect 3218 25671 3234 25705
rect 3268 25671 3284 25705
rect 3410 25671 3426 25705
rect 3460 25671 3476 25705
rect 3540 25607 3574 25680
rect 2352 25573 2470 25607
rect 2504 25573 2538 25607
rect 2572 25573 2606 25607
rect 2640 25573 2674 25607
rect 2708 25573 2742 25607
rect 2776 25573 2810 25607
rect 2844 25573 2878 25607
rect 2912 25573 2946 25607
rect 2980 25573 3014 25607
rect 3048 25573 3082 25607
rect 3116 25573 3150 25607
rect 3184 25573 3218 25607
rect 3252 25573 3286 25607
rect 3320 25573 3354 25607
rect 3388 25573 3422 25607
rect 3456 25573 3574 25607
rect 3873 25717 3907 25751
rect 3987 25816 4021 25855
rect 3987 25743 4021 25782
rect 4083 25816 4117 25855
rect 4083 25743 4117 25782
rect 4179 25816 4213 25855
rect 4179 25743 4213 25782
rect 4275 25816 4309 25855
rect 4275 25743 4309 25782
rect 4371 25816 4405 25855
rect 4371 25743 4405 25782
rect 4467 25816 4501 25855
rect 4467 25743 4501 25782
rect 4563 25816 4597 25855
rect 4563 25743 4597 25782
rect 4659 25816 4693 25855
rect 4659 25743 4693 25782
rect 4755 25816 4789 25855
rect 4755 25743 4789 25782
rect 4851 25816 4885 25855
rect 4851 25743 4885 25782
rect 4947 25816 4981 25855
rect 4947 25743 4981 25782
rect 5061 25786 5095 25819
rect 5340 25934 5348 25968
rect 5382 25934 5386 25968
rect 5420 25973 5486 25984
rect 5420 25970 5450 25973
rect 5420 25936 5436 25970
rect 5484 25939 5486 25973
rect 5470 25936 5486 25939
rect 5340 25898 5386 25934
rect 5340 25886 5406 25898
rect 5340 25852 5356 25886
rect 5390 25852 5406 25886
rect 5340 25818 5406 25852
rect 5340 25784 5356 25818
rect 5390 25784 5406 25818
rect 5340 25772 5406 25784
rect 5440 25886 5486 25902
rect 5474 25852 5486 25886
rect 5440 25818 5486 25852
rect 5474 25784 5486 25818
rect 5061 25717 5095 25751
rect 5440 25738 5486 25784
rect 3873 25607 3907 25683
rect 3971 25671 3987 25705
rect 4021 25671 4037 25705
rect 4163 25671 4179 25705
rect 4213 25671 4229 25705
rect 4355 25671 4371 25705
rect 4405 25671 4421 25705
rect 4547 25671 4563 25705
rect 4597 25671 4613 25705
rect 4739 25671 4755 25705
rect 4789 25671 4805 25705
rect 4931 25671 4947 25705
rect 4981 25671 4997 25705
rect 5274 25704 5303 25738
rect 5337 25704 5395 25738
rect 5429 25704 5487 25738
rect 5521 25704 5550 25738
rect 5061 25607 5095 25680
rect 3873 25573 3991 25607
rect 4025 25573 4059 25607
rect 4093 25573 4127 25607
rect 4161 25573 4195 25607
rect 4229 25573 4263 25607
rect 4297 25573 4331 25607
rect 4365 25573 4399 25607
rect 4433 25573 4467 25607
rect 4501 25573 4535 25607
rect 4569 25573 4603 25607
rect 4637 25573 4671 25607
rect 4705 25573 4739 25607
rect 4773 25573 4807 25607
rect 4841 25573 4875 25607
rect 4909 25573 4943 25607
rect 4977 25573 5095 25607
rect 199 25290 317 25324
rect 351 25290 385 25324
rect 419 25290 453 25324
rect 487 25290 521 25324
rect 555 25290 589 25324
rect 623 25290 657 25324
rect 691 25290 725 25324
rect 759 25290 793 25324
rect 827 25290 861 25324
rect 895 25290 929 25324
rect 963 25290 997 25324
rect 1031 25290 1065 25324
rect 1099 25290 1133 25324
rect 1167 25290 1201 25324
rect 1235 25290 1269 25324
rect 1303 25290 1421 25324
rect 199 25222 233 25290
rect 1387 25222 1421 25290
rect 297 25188 313 25222
rect 347 25188 363 25222
rect 489 25188 505 25222
rect 539 25188 555 25222
rect 681 25188 697 25222
rect 731 25188 747 25222
rect 873 25188 889 25222
rect 923 25188 939 25222
rect 1065 25188 1081 25222
rect 1115 25188 1131 25222
rect 1257 25188 1273 25222
rect 1307 25188 1323 25222
rect 199 25154 233 25188
rect 1387 25154 1421 25162
rect 199 25086 233 25120
rect 199 25018 233 25052
rect 199 24950 233 24984
rect 199 24882 233 24916
rect 313 25123 347 25144
rect 313 25055 347 25059
rect 313 24949 347 24953
rect 313 24864 347 24885
rect 409 25123 443 25144
rect 409 25055 443 25059
rect 409 24949 443 24953
rect 409 24864 443 24885
rect 505 25123 539 25144
rect 505 25055 539 25059
rect 505 24949 539 24953
rect 505 24864 539 24885
rect 601 25123 635 25144
rect 601 25055 635 25059
rect 601 24949 635 24953
rect 601 24864 635 24885
rect 697 25123 731 25144
rect 697 25055 731 25059
rect 697 24949 731 24953
rect 697 24864 731 24885
rect 793 25123 827 25144
rect 793 25055 827 25059
rect 793 24949 827 24953
rect 793 24864 827 24885
rect 889 25123 923 25144
rect 889 25055 923 25059
rect 889 24949 923 24953
rect 889 24864 923 24885
rect 985 25123 1019 25144
rect 985 25055 1019 25059
rect 985 24949 1019 24953
rect 985 24864 1019 24885
rect 1081 25123 1115 25144
rect 1081 25055 1115 25059
rect 1081 24949 1115 24953
rect 1081 24864 1115 24885
rect 1177 25123 1211 25144
rect 1177 25055 1211 25059
rect 1177 24949 1211 24953
rect 1177 24864 1211 24885
rect 1273 25123 1307 25144
rect 1273 25055 1307 25059
rect 1273 24949 1307 24953
rect 1273 24864 1307 24885
rect 1387 25086 1421 25090
rect 1387 24980 1421 24984
rect 1387 24908 1421 24916
rect 199 24780 233 24848
rect 1387 24780 1421 24848
rect 199 24746 317 24780
rect 351 24746 385 24780
rect 419 24746 453 24780
rect 487 24746 521 24780
rect 555 24746 589 24780
rect 623 24746 657 24780
rect 691 24746 725 24780
rect 759 24746 793 24780
rect 827 24746 861 24780
rect 895 24746 929 24780
rect 963 24746 997 24780
rect 1031 24746 1065 24780
rect 1099 24746 1133 24780
rect 1167 24746 1201 24780
rect 1235 24746 1269 24780
rect 1303 24746 1421 24780
rect 2352 25294 2470 25328
rect 2504 25294 2538 25328
rect 2572 25294 2606 25328
rect 2640 25294 2674 25328
rect 2708 25294 2742 25328
rect 2776 25294 2810 25328
rect 2844 25294 2878 25328
rect 2912 25294 2946 25328
rect 2980 25294 3014 25328
rect 3048 25294 3082 25328
rect 3116 25294 3150 25328
rect 3184 25294 3218 25328
rect 3252 25294 3286 25328
rect 3320 25294 3354 25328
rect 3388 25294 3422 25328
rect 3456 25294 3574 25328
rect 2352 25226 2386 25294
rect 3540 25226 3574 25294
rect 2450 25192 2466 25226
rect 2500 25192 2516 25226
rect 2642 25192 2658 25226
rect 2692 25192 2708 25226
rect 2834 25192 2850 25226
rect 2884 25192 2900 25226
rect 3026 25192 3042 25226
rect 3076 25192 3092 25226
rect 3218 25192 3234 25226
rect 3268 25192 3284 25226
rect 3410 25192 3426 25226
rect 3460 25192 3476 25226
rect 2352 25158 2386 25192
rect 3540 25158 3574 25166
rect 2352 25090 2386 25124
rect 2352 25022 2386 25056
rect 2352 24954 2386 24988
rect 2352 24886 2386 24920
rect 2466 25127 2500 25148
rect 2466 25059 2500 25063
rect 2466 24953 2500 24957
rect 2466 24868 2500 24889
rect 2562 25127 2596 25148
rect 2562 25059 2596 25063
rect 2562 24953 2596 24957
rect 2562 24868 2596 24889
rect 2658 25127 2692 25148
rect 2658 25059 2692 25063
rect 2658 24953 2692 24957
rect 2658 24868 2692 24889
rect 2754 25127 2788 25148
rect 2754 25059 2788 25063
rect 2754 24953 2788 24957
rect 2754 24868 2788 24889
rect 2850 25127 2884 25148
rect 2850 25059 2884 25063
rect 2850 24953 2884 24957
rect 2850 24868 2884 24889
rect 2946 25127 2980 25148
rect 2946 25059 2980 25063
rect 2946 24953 2980 24957
rect 2946 24868 2980 24889
rect 3042 25127 3076 25148
rect 3042 25059 3076 25063
rect 3042 24953 3076 24957
rect 3042 24868 3076 24889
rect 3138 25127 3172 25148
rect 3138 25059 3172 25063
rect 3138 24953 3172 24957
rect 3138 24868 3172 24889
rect 3234 25127 3268 25148
rect 3234 25059 3268 25063
rect 3234 24953 3268 24957
rect 3234 24868 3268 24889
rect 3330 25127 3364 25148
rect 3330 25059 3364 25063
rect 3330 24953 3364 24957
rect 3330 24868 3364 24889
rect 3426 25127 3460 25148
rect 3426 25059 3460 25063
rect 3426 24953 3460 24957
rect 3426 24868 3460 24889
rect 3540 25090 3574 25094
rect 3540 24984 3574 24988
rect 3540 24912 3574 24920
rect 2352 24784 2386 24852
rect 3540 24784 3574 24852
rect 2352 24750 2470 24784
rect 2504 24750 2538 24784
rect 2572 24750 2606 24784
rect 2640 24750 2674 24784
rect 2708 24750 2742 24784
rect 2776 24750 2810 24784
rect 2844 24750 2878 24784
rect 2912 24750 2946 24784
rect 2980 24750 3014 24784
rect 3048 24750 3082 24784
rect 3116 24750 3150 24784
rect 3184 24750 3218 24784
rect 3252 24750 3286 24784
rect 3320 24750 3354 24784
rect 3388 24750 3422 24784
rect 3456 24750 3574 24784
rect 3873 25294 3991 25328
rect 4025 25294 4059 25328
rect 4093 25294 4127 25328
rect 4161 25294 4195 25328
rect 4229 25294 4263 25328
rect 4297 25294 4331 25328
rect 4365 25294 4399 25328
rect 4433 25294 4467 25328
rect 4501 25294 4535 25328
rect 4569 25294 4603 25328
rect 4637 25294 4671 25328
rect 4705 25294 4739 25328
rect 4773 25294 4807 25328
rect 4841 25294 4875 25328
rect 4909 25294 4943 25328
rect 4977 25294 5095 25328
rect 3873 25226 3907 25294
rect 5061 25226 5095 25294
rect 3971 25192 3987 25226
rect 4021 25192 4037 25226
rect 4163 25192 4179 25226
rect 4213 25192 4229 25226
rect 4355 25192 4371 25226
rect 4405 25192 4421 25226
rect 4547 25192 4563 25226
rect 4597 25192 4613 25226
rect 4739 25192 4755 25226
rect 4789 25192 4805 25226
rect 4931 25192 4947 25226
rect 4981 25192 4997 25226
rect 3873 25158 3907 25192
rect 5061 25158 5095 25166
rect 3873 25090 3907 25124
rect 3873 25022 3907 25056
rect 3873 24954 3907 24988
rect 3873 24886 3907 24920
rect 3987 25127 4021 25148
rect 3987 25059 4021 25063
rect 3987 24953 4021 24957
rect 3987 24868 4021 24889
rect 4083 25127 4117 25148
rect 4083 25059 4117 25063
rect 4083 24953 4117 24957
rect 4083 24868 4117 24889
rect 4179 25127 4213 25148
rect 4179 25059 4213 25063
rect 4179 24953 4213 24957
rect 4179 24868 4213 24889
rect 4275 25127 4309 25148
rect 4275 25059 4309 25063
rect 4275 24953 4309 24957
rect 4275 24868 4309 24889
rect 4371 25127 4405 25148
rect 4371 25059 4405 25063
rect 4371 24953 4405 24957
rect 4371 24868 4405 24889
rect 4467 25127 4501 25148
rect 4467 25059 4501 25063
rect 4467 24953 4501 24957
rect 4467 24868 4501 24889
rect 4563 25127 4597 25148
rect 4563 25059 4597 25063
rect 4563 24953 4597 24957
rect 4563 24868 4597 24889
rect 4659 25127 4693 25148
rect 4659 25059 4693 25063
rect 4659 24953 4693 24957
rect 4659 24868 4693 24889
rect 4755 25127 4789 25148
rect 4755 25059 4789 25063
rect 4755 24953 4789 24957
rect 4755 24868 4789 24889
rect 4851 25127 4885 25148
rect 4851 25059 4885 25063
rect 4851 24953 4885 24957
rect 4851 24868 4885 24889
rect 4947 25127 4981 25148
rect 4947 25059 4981 25063
rect 4947 24953 4981 24957
rect 4947 24868 4981 24889
rect 5061 25090 5095 25094
rect 5061 24984 5095 24988
rect 5274 24961 5303 24995
rect 5337 24961 5395 24995
rect 5429 24961 5487 24995
rect 5521 24961 5550 24995
rect 5061 24912 5095 24920
rect 3873 24784 3907 24852
rect 5061 24784 5095 24852
rect 3873 24750 3991 24784
rect 4025 24750 4059 24784
rect 4093 24750 4127 24784
rect 4161 24750 4195 24784
rect 4229 24750 4263 24784
rect 4297 24750 4331 24784
rect 4365 24750 4399 24784
rect 4433 24750 4467 24784
rect 4501 24750 4535 24784
rect 4569 24750 4603 24784
rect 4637 24750 4671 24784
rect 4705 24750 4739 24784
rect 4773 24750 4807 24784
rect 4841 24750 4875 24784
rect 4909 24750 4943 24784
rect 4977 24750 5095 24784
rect 5340 24919 5406 24927
rect 5340 24885 5356 24919
rect 5390 24885 5406 24919
rect 5340 24851 5406 24885
rect 5340 24817 5356 24851
rect 5390 24817 5406 24851
rect 5340 24783 5406 24817
rect 5340 24749 5356 24783
rect 5390 24749 5406 24783
rect 5340 24731 5406 24749
rect 5440 24919 5482 24961
rect 5474 24885 5482 24919
rect 5440 24851 5482 24885
rect 5474 24817 5482 24851
rect 5440 24783 5482 24817
rect 5474 24749 5482 24783
rect 5440 24733 5482 24749
rect 5340 24681 5386 24731
rect 199 24638 317 24672
rect 351 24638 385 24672
rect 419 24638 453 24672
rect 487 24638 521 24672
rect 555 24638 589 24672
rect 623 24638 657 24672
rect 691 24638 725 24672
rect 759 24638 793 24672
rect 827 24638 861 24672
rect 895 24638 929 24672
rect 963 24638 997 24672
rect 1031 24638 1065 24672
rect 1099 24638 1133 24672
rect 1167 24638 1201 24672
rect 1235 24638 1269 24672
rect 1303 24638 1421 24672
rect 199 24562 233 24638
rect 1387 24567 1421 24638
rect 199 24494 233 24528
rect 199 24426 233 24460
rect 313 24525 347 24564
rect 313 24452 347 24491
rect 409 24525 443 24564
rect 409 24452 443 24491
rect 505 24525 539 24564
rect 505 24452 539 24491
rect 601 24525 635 24564
rect 601 24452 635 24491
rect 697 24525 731 24564
rect 697 24452 731 24491
rect 793 24525 827 24564
rect 793 24452 827 24491
rect 889 24525 923 24564
rect 889 24452 923 24491
rect 985 24525 1019 24564
rect 985 24452 1019 24491
rect 1081 24525 1115 24564
rect 1081 24452 1115 24491
rect 1177 24525 1211 24564
rect 1177 24452 1211 24491
rect 1273 24525 1307 24564
rect 1273 24452 1307 24491
rect 1387 24495 1421 24528
rect 1387 24426 1421 24460
rect 199 24316 233 24392
rect 297 24380 313 24414
rect 347 24380 363 24414
rect 489 24380 505 24414
rect 539 24380 555 24414
rect 681 24380 697 24414
rect 731 24380 747 24414
rect 873 24380 889 24414
rect 923 24380 939 24414
rect 1065 24380 1081 24414
rect 1115 24380 1131 24414
rect 1257 24380 1273 24414
rect 1307 24380 1323 24414
rect 1387 24316 1421 24389
rect 199 24282 317 24316
rect 351 24282 385 24316
rect 419 24282 453 24316
rect 487 24282 521 24316
rect 555 24282 589 24316
rect 623 24282 657 24316
rect 691 24282 725 24316
rect 759 24282 793 24316
rect 827 24282 861 24316
rect 895 24282 929 24316
rect 963 24282 997 24316
rect 1031 24282 1065 24316
rect 1099 24282 1133 24316
rect 1167 24282 1201 24316
rect 1235 24282 1269 24316
rect 1303 24282 1421 24316
rect 2352 24642 2470 24676
rect 2504 24642 2538 24676
rect 2572 24642 2606 24676
rect 2640 24642 2674 24676
rect 2708 24642 2742 24676
rect 2776 24642 2810 24676
rect 2844 24642 2878 24676
rect 2912 24642 2946 24676
rect 2980 24642 3014 24676
rect 3048 24642 3082 24676
rect 3116 24642 3150 24676
rect 3184 24642 3218 24676
rect 3252 24642 3286 24676
rect 3320 24642 3354 24676
rect 3388 24642 3422 24676
rect 3456 24642 3574 24676
rect 2352 24566 2386 24642
rect 3540 24571 3574 24642
rect 3873 24642 3991 24676
rect 4025 24642 4059 24676
rect 4093 24642 4127 24676
rect 4161 24642 4195 24676
rect 4229 24642 4263 24676
rect 4297 24642 4331 24676
rect 4365 24642 4399 24676
rect 4433 24642 4467 24676
rect 4501 24642 4535 24676
rect 4569 24642 4603 24676
rect 4637 24642 4671 24676
rect 4705 24642 4739 24676
rect 4773 24642 4807 24676
rect 4841 24642 4875 24676
rect 4909 24642 4943 24676
rect 4977 24642 5095 24676
rect 3675 24606 3691 24640
rect 3725 24606 3741 24640
rect 2352 24498 2386 24532
rect 2352 24430 2386 24464
rect 2466 24529 2500 24568
rect 2466 24456 2500 24495
rect 2562 24529 2596 24568
rect 2562 24456 2596 24495
rect 2658 24529 2692 24568
rect 2658 24456 2692 24495
rect 2754 24529 2788 24568
rect 2754 24456 2788 24495
rect 2850 24529 2884 24568
rect 2850 24456 2884 24495
rect 2946 24529 2980 24568
rect 2946 24456 2980 24495
rect 3042 24529 3076 24568
rect 3042 24456 3076 24495
rect 3138 24529 3172 24568
rect 3138 24456 3172 24495
rect 3234 24529 3268 24568
rect 3234 24456 3268 24495
rect 3330 24529 3364 24568
rect 3330 24456 3364 24495
rect 3426 24529 3460 24568
rect 3426 24456 3460 24495
rect 3540 24499 3574 24532
rect 3647 24556 3681 24572
rect 3647 24464 3681 24480
rect 3735 24556 3769 24572
rect 3735 24464 3769 24480
rect 3873 24566 3907 24642
rect 5061 24571 5095 24642
rect 3873 24498 3907 24532
rect 3540 24430 3574 24464
rect 2352 24320 2386 24396
rect 2450 24384 2466 24418
rect 2500 24384 2516 24418
rect 2642 24384 2658 24418
rect 2692 24384 2708 24418
rect 2834 24384 2850 24418
rect 2884 24384 2900 24418
rect 3026 24384 3042 24418
rect 3076 24384 3092 24418
rect 3218 24384 3234 24418
rect 3268 24384 3284 24418
rect 3410 24384 3426 24418
rect 3460 24384 3476 24418
rect 3540 24320 3574 24393
rect 2352 24286 2470 24320
rect 2504 24286 2538 24320
rect 2572 24286 2606 24320
rect 2640 24286 2674 24320
rect 2708 24286 2742 24320
rect 2776 24286 2810 24320
rect 2844 24286 2878 24320
rect 2912 24286 2946 24320
rect 2980 24286 3014 24320
rect 3048 24286 3082 24320
rect 3116 24286 3150 24320
rect 3184 24286 3218 24320
rect 3252 24286 3286 24320
rect 3320 24286 3354 24320
rect 3388 24286 3422 24320
rect 3456 24286 3574 24320
rect 3873 24430 3907 24464
rect 3987 24529 4021 24568
rect 3987 24456 4021 24495
rect 4083 24529 4117 24568
rect 4083 24456 4117 24495
rect 4179 24529 4213 24568
rect 4179 24456 4213 24495
rect 4275 24529 4309 24568
rect 4275 24456 4309 24495
rect 4371 24529 4405 24568
rect 4371 24456 4405 24495
rect 4467 24529 4501 24568
rect 4467 24456 4501 24495
rect 4563 24529 4597 24568
rect 4563 24456 4597 24495
rect 4659 24529 4693 24568
rect 4659 24456 4693 24495
rect 4755 24529 4789 24568
rect 4755 24456 4789 24495
rect 4851 24529 4885 24568
rect 4851 24456 4885 24495
rect 4947 24529 4981 24568
rect 4947 24456 4981 24495
rect 5061 24499 5095 24532
rect 5340 24647 5348 24681
rect 5382 24647 5386 24681
rect 5420 24686 5486 24697
rect 5420 24683 5450 24686
rect 5420 24649 5436 24683
rect 5484 24652 5486 24686
rect 5470 24649 5486 24652
rect 5340 24611 5386 24647
rect 5340 24599 5406 24611
rect 5340 24565 5356 24599
rect 5390 24565 5406 24599
rect 5340 24531 5406 24565
rect 5340 24497 5356 24531
rect 5390 24497 5406 24531
rect 5340 24485 5406 24497
rect 5440 24599 5486 24615
rect 5474 24565 5486 24599
rect 5440 24531 5486 24565
rect 5474 24497 5486 24531
rect 5061 24430 5095 24464
rect 5440 24451 5486 24497
rect 3873 24320 3907 24396
rect 3971 24384 3987 24418
rect 4021 24384 4037 24418
rect 4163 24384 4179 24418
rect 4213 24384 4229 24418
rect 4355 24384 4371 24418
rect 4405 24384 4421 24418
rect 4547 24384 4563 24418
rect 4597 24384 4613 24418
rect 4739 24384 4755 24418
rect 4789 24384 4805 24418
rect 4931 24384 4947 24418
rect 4981 24384 4997 24418
rect 5274 24417 5303 24451
rect 5337 24417 5395 24451
rect 5429 24417 5487 24451
rect 5521 24417 5550 24451
rect 5061 24320 5095 24393
rect 3873 24286 3991 24320
rect 4025 24286 4059 24320
rect 4093 24286 4127 24320
rect 4161 24286 4195 24320
rect 4229 24286 4263 24320
rect 4297 24286 4331 24320
rect 4365 24286 4399 24320
rect 4433 24286 4467 24320
rect 4501 24286 4535 24320
rect 4569 24286 4603 24320
rect 4637 24286 4671 24320
rect 4705 24286 4739 24320
rect 4773 24286 4807 24320
rect 4841 24286 4875 24320
rect 4909 24286 4943 24320
rect 4977 24286 5095 24320
rect 199 24003 317 24037
rect 351 24003 385 24037
rect 419 24003 453 24037
rect 487 24003 521 24037
rect 555 24003 589 24037
rect 623 24003 657 24037
rect 691 24003 725 24037
rect 759 24003 793 24037
rect 827 24003 861 24037
rect 895 24003 929 24037
rect 963 24003 997 24037
rect 1031 24003 1065 24037
rect 1099 24003 1133 24037
rect 1167 24003 1201 24037
rect 1235 24003 1269 24037
rect 1303 24003 1421 24037
rect 199 23935 233 24003
rect 1387 23935 1421 24003
rect 297 23901 313 23935
rect 347 23901 363 23935
rect 489 23901 505 23935
rect 539 23901 555 23935
rect 681 23901 697 23935
rect 731 23901 747 23935
rect 873 23901 889 23935
rect 923 23901 939 23935
rect 1065 23901 1081 23935
rect 1115 23901 1131 23935
rect 1257 23901 1273 23935
rect 1307 23901 1323 23935
rect 199 23867 233 23901
rect 1387 23867 1421 23875
rect 199 23799 233 23833
rect 199 23731 233 23765
rect 199 23663 233 23697
rect 199 23595 233 23629
rect 313 23836 347 23857
rect 313 23768 347 23772
rect 313 23662 347 23666
rect 313 23577 347 23598
rect 409 23836 443 23857
rect 409 23768 443 23772
rect 409 23662 443 23666
rect 409 23577 443 23598
rect 505 23836 539 23857
rect 505 23768 539 23772
rect 505 23662 539 23666
rect 505 23577 539 23598
rect 601 23836 635 23857
rect 601 23768 635 23772
rect 601 23662 635 23666
rect 601 23577 635 23598
rect 697 23836 731 23857
rect 697 23768 731 23772
rect 697 23662 731 23666
rect 697 23577 731 23598
rect 793 23836 827 23857
rect 793 23768 827 23772
rect 793 23662 827 23666
rect 793 23577 827 23598
rect 889 23836 923 23857
rect 889 23768 923 23772
rect 889 23662 923 23666
rect 889 23577 923 23598
rect 985 23836 1019 23857
rect 985 23768 1019 23772
rect 985 23662 1019 23666
rect 985 23577 1019 23598
rect 1081 23836 1115 23857
rect 1081 23768 1115 23772
rect 1081 23662 1115 23666
rect 1081 23577 1115 23598
rect 1177 23836 1211 23857
rect 1177 23768 1211 23772
rect 1177 23662 1211 23666
rect 1177 23577 1211 23598
rect 1273 23836 1307 23857
rect 1273 23768 1307 23772
rect 1273 23662 1307 23666
rect 1273 23577 1307 23598
rect 1387 23799 1421 23803
rect 1387 23693 1421 23697
rect 1387 23621 1421 23629
rect 199 23493 233 23561
rect 1387 23493 1421 23561
rect 199 23459 317 23493
rect 351 23459 385 23493
rect 419 23459 453 23493
rect 487 23459 521 23493
rect 555 23459 589 23493
rect 623 23459 657 23493
rect 691 23459 725 23493
rect 759 23459 793 23493
rect 827 23459 861 23493
rect 895 23459 929 23493
rect 963 23459 997 23493
rect 1031 23459 1065 23493
rect 1099 23459 1133 23493
rect 1167 23459 1201 23493
rect 1235 23459 1269 23493
rect 1303 23459 1421 23493
rect 2352 24007 2470 24041
rect 2504 24007 2538 24041
rect 2572 24007 2606 24041
rect 2640 24007 2674 24041
rect 2708 24007 2742 24041
rect 2776 24007 2810 24041
rect 2844 24007 2878 24041
rect 2912 24007 2946 24041
rect 2980 24007 3014 24041
rect 3048 24007 3082 24041
rect 3116 24007 3150 24041
rect 3184 24007 3218 24041
rect 3252 24007 3286 24041
rect 3320 24007 3354 24041
rect 3388 24007 3422 24041
rect 3456 24007 3574 24041
rect 2352 23939 2386 24007
rect 3540 23939 3574 24007
rect 2450 23905 2466 23939
rect 2500 23905 2516 23939
rect 2642 23905 2658 23939
rect 2692 23905 2708 23939
rect 2834 23905 2850 23939
rect 2884 23905 2900 23939
rect 3026 23905 3042 23939
rect 3076 23905 3092 23939
rect 3218 23905 3234 23939
rect 3268 23905 3284 23939
rect 3410 23905 3426 23939
rect 3460 23905 3476 23939
rect 2352 23871 2386 23905
rect 3540 23871 3574 23879
rect 2352 23803 2386 23837
rect 2352 23735 2386 23769
rect 2352 23667 2386 23701
rect 2352 23599 2386 23633
rect 2466 23840 2500 23861
rect 2466 23772 2500 23776
rect 2466 23666 2500 23670
rect 2466 23581 2500 23602
rect 2562 23840 2596 23861
rect 2562 23772 2596 23776
rect 2562 23666 2596 23670
rect 2562 23581 2596 23602
rect 2658 23840 2692 23861
rect 2658 23772 2692 23776
rect 2658 23666 2692 23670
rect 2658 23581 2692 23602
rect 2754 23840 2788 23861
rect 2754 23772 2788 23776
rect 2754 23666 2788 23670
rect 2754 23581 2788 23602
rect 2850 23840 2884 23861
rect 2850 23772 2884 23776
rect 2850 23666 2884 23670
rect 2850 23581 2884 23602
rect 2946 23840 2980 23861
rect 2946 23772 2980 23776
rect 2946 23666 2980 23670
rect 2946 23581 2980 23602
rect 3042 23840 3076 23861
rect 3042 23772 3076 23776
rect 3042 23666 3076 23670
rect 3042 23581 3076 23602
rect 3138 23840 3172 23861
rect 3138 23772 3172 23776
rect 3138 23666 3172 23670
rect 3138 23581 3172 23602
rect 3234 23840 3268 23861
rect 3234 23772 3268 23776
rect 3234 23666 3268 23670
rect 3234 23581 3268 23602
rect 3330 23840 3364 23861
rect 3330 23772 3364 23776
rect 3330 23666 3364 23670
rect 3330 23581 3364 23602
rect 3426 23840 3460 23861
rect 3426 23772 3460 23776
rect 3426 23666 3460 23670
rect 3426 23581 3460 23602
rect 3540 23803 3574 23807
rect 3540 23697 3574 23701
rect 3540 23625 3574 23633
rect 2352 23497 2386 23565
rect 3540 23497 3574 23565
rect 2352 23463 2470 23497
rect 2504 23463 2538 23497
rect 2572 23463 2606 23497
rect 2640 23463 2674 23497
rect 2708 23463 2742 23497
rect 2776 23463 2810 23497
rect 2844 23463 2878 23497
rect 2912 23463 2946 23497
rect 2980 23463 3014 23497
rect 3048 23463 3082 23497
rect 3116 23463 3150 23497
rect 3184 23463 3218 23497
rect 3252 23463 3286 23497
rect 3320 23463 3354 23497
rect 3388 23463 3422 23497
rect 3456 23463 3574 23497
rect 3873 24007 3991 24041
rect 4025 24007 4059 24041
rect 4093 24007 4127 24041
rect 4161 24007 4195 24041
rect 4229 24007 4263 24041
rect 4297 24007 4331 24041
rect 4365 24007 4399 24041
rect 4433 24007 4467 24041
rect 4501 24007 4535 24041
rect 4569 24007 4603 24041
rect 4637 24007 4671 24041
rect 4705 24007 4739 24041
rect 4773 24007 4807 24041
rect 4841 24007 4875 24041
rect 4909 24007 4943 24041
rect 4977 24007 5095 24041
rect 3873 23939 3907 24007
rect 5061 23939 5095 24007
rect 3971 23905 3987 23939
rect 4021 23905 4037 23939
rect 4163 23905 4179 23939
rect 4213 23905 4229 23939
rect 4355 23905 4371 23939
rect 4405 23905 4421 23939
rect 4547 23905 4563 23939
rect 4597 23905 4613 23939
rect 4739 23905 4755 23939
rect 4789 23905 4805 23939
rect 4931 23905 4947 23939
rect 4981 23905 4997 23939
rect 3873 23871 3907 23905
rect 5061 23871 5095 23879
rect 3873 23803 3907 23837
rect 3873 23735 3907 23769
rect 3873 23667 3907 23701
rect 3873 23599 3907 23633
rect 3987 23840 4021 23861
rect 3987 23772 4021 23776
rect 3987 23666 4021 23670
rect 3987 23581 4021 23602
rect 4083 23840 4117 23861
rect 4083 23772 4117 23776
rect 4083 23666 4117 23670
rect 4083 23581 4117 23602
rect 4179 23840 4213 23861
rect 4179 23772 4213 23776
rect 4179 23666 4213 23670
rect 4179 23581 4213 23602
rect 4275 23840 4309 23861
rect 4275 23772 4309 23776
rect 4275 23666 4309 23670
rect 4275 23581 4309 23602
rect 4371 23840 4405 23861
rect 4371 23772 4405 23776
rect 4371 23666 4405 23670
rect 4371 23581 4405 23602
rect 4467 23840 4501 23861
rect 4467 23772 4501 23776
rect 4467 23666 4501 23670
rect 4467 23581 4501 23602
rect 4563 23840 4597 23861
rect 4563 23772 4597 23776
rect 4563 23666 4597 23670
rect 4563 23581 4597 23602
rect 4659 23840 4693 23861
rect 4659 23772 4693 23776
rect 4659 23666 4693 23670
rect 4659 23581 4693 23602
rect 4755 23840 4789 23861
rect 4755 23772 4789 23776
rect 4755 23666 4789 23670
rect 4755 23581 4789 23602
rect 4851 23840 4885 23861
rect 4851 23772 4885 23776
rect 4851 23666 4885 23670
rect 4851 23581 4885 23602
rect 4947 23840 4981 23861
rect 4947 23772 4981 23776
rect 4947 23666 4981 23670
rect 4947 23581 4981 23602
rect 5061 23803 5095 23807
rect 5061 23697 5095 23701
rect 5274 23674 5303 23708
rect 5337 23674 5395 23708
rect 5429 23674 5487 23708
rect 5521 23674 5550 23708
rect 5061 23625 5095 23633
rect 3873 23497 3907 23565
rect 5061 23497 5095 23565
rect 3873 23463 3991 23497
rect 4025 23463 4059 23497
rect 4093 23463 4127 23497
rect 4161 23463 4195 23497
rect 4229 23463 4263 23497
rect 4297 23463 4331 23497
rect 4365 23463 4399 23497
rect 4433 23463 4467 23497
rect 4501 23463 4535 23497
rect 4569 23463 4603 23497
rect 4637 23463 4671 23497
rect 4705 23463 4739 23497
rect 4773 23463 4807 23497
rect 4841 23463 4875 23497
rect 4909 23463 4943 23497
rect 4977 23463 5095 23497
rect 5340 23632 5406 23640
rect 5340 23598 5356 23632
rect 5390 23598 5406 23632
rect 5340 23564 5406 23598
rect 5340 23530 5356 23564
rect 5390 23530 5406 23564
rect 5340 23496 5406 23530
rect 5340 23462 5356 23496
rect 5390 23462 5406 23496
rect 5340 23444 5406 23462
rect 5440 23632 5482 23674
rect 5474 23598 5482 23632
rect 5440 23564 5482 23598
rect 5474 23530 5482 23564
rect 5440 23496 5482 23530
rect 5474 23462 5482 23496
rect 5440 23446 5482 23462
rect 5340 23394 5386 23444
rect 199 23351 317 23385
rect 351 23351 385 23385
rect 419 23351 453 23385
rect 487 23351 521 23385
rect 555 23351 589 23385
rect 623 23351 657 23385
rect 691 23351 725 23385
rect 759 23351 793 23385
rect 827 23351 861 23385
rect 895 23351 929 23385
rect 963 23351 997 23385
rect 1031 23351 1065 23385
rect 1099 23351 1133 23385
rect 1167 23351 1201 23385
rect 1235 23351 1269 23385
rect 1303 23351 1421 23385
rect 199 23275 233 23351
rect 1387 23280 1421 23351
rect 199 23207 233 23241
rect 199 23139 233 23173
rect 313 23238 347 23277
rect 313 23165 347 23204
rect 409 23238 443 23277
rect 409 23165 443 23204
rect 505 23238 539 23277
rect 505 23165 539 23204
rect 601 23238 635 23277
rect 601 23165 635 23204
rect 697 23238 731 23277
rect 697 23165 731 23204
rect 793 23238 827 23277
rect 793 23165 827 23204
rect 889 23238 923 23277
rect 889 23165 923 23204
rect 985 23238 1019 23277
rect 985 23165 1019 23204
rect 1081 23238 1115 23277
rect 1081 23165 1115 23204
rect 1177 23238 1211 23277
rect 1177 23165 1211 23204
rect 1273 23238 1307 23277
rect 1273 23165 1307 23204
rect 1387 23208 1421 23241
rect 1387 23139 1421 23173
rect 199 23029 233 23105
rect 297 23093 313 23127
rect 347 23093 363 23127
rect 489 23093 505 23127
rect 539 23093 555 23127
rect 681 23093 697 23127
rect 731 23093 747 23127
rect 873 23093 889 23127
rect 923 23093 939 23127
rect 1065 23093 1081 23127
rect 1115 23093 1131 23127
rect 1257 23093 1273 23127
rect 1307 23093 1323 23127
rect 1387 23029 1421 23102
rect 199 22995 317 23029
rect 351 22995 385 23029
rect 419 22995 453 23029
rect 487 22995 521 23029
rect 555 22995 589 23029
rect 623 22995 657 23029
rect 691 22995 725 23029
rect 759 22995 793 23029
rect 827 22995 861 23029
rect 895 22995 929 23029
rect 963 22995 997 23029
rect 1031 22995 1065 23029
rect 1099 22995 1133 23029
rect 1167 22995 1201 23029
rect 1235 22995 1269 23029
rect 1303 22995 1421 23029
rect 2352 23355 2470 23389
rect 2504 23355 2538 23389
rect 2572 23355 2606 23389
rect 2640 23355 2674 23389
rect 2708 23355 2742 23389
rect 2776 23355 2810 23389
rect 2844 23355 2878 23389
rect 2912 23355 2946 23389
rect 2980 23355 3014 23389
rect 3048 23355 3082 23389
rect 3116 23355 3150 23389
rect 3184 23355 3218 23389
rect 3252 23355 3286 23389
rect 3320 23355 3354 23389
rect 3388 23355 3422 23389
rect 3456 23355 3574 23389
rect 2352 23279 2386 23355
rect 3540 23284 3574 23355
rect 3873 23355 3991 23389
rect 4025 23355 4059 23389
rect 4093 23355 4127 23389
rect 4161 23355 4195 23389
rect 4229 23355 4263 23389
rect 4297 23355 4331 23389
rect 4365 23355 4399 23389
rect 4433 23355 4467 23389
rect 4501 23355 4535 23389
rect 4569 23355 4603 23389
rect 4637 23355 4671 23389
rect 4705 23355 4739 23389
rect 4773 23355 4807 23389
rect 4841 23355 4875 23389
rect 4909 23355 4943 23389
rect 4977 23355 5095 23389
rect 3675 23319 3691 23353
rect 3725 23319 3741 23353
rect 2352 23211 2386 23245
rect 2352 23143 2386 23177
rect 2466 23242 2500 23281
rect 2466 23169 2500 23208
rect 2562 23242 2596 23281
rect 2562 23169 2596 23208
rect 2658 23242 2692 23281
rect 2658 23169 2692 23208
rect 2754 23242 2788 23281
rect 2754 23169 2788 23208
rect 2850 23242 2884 23281
rect 2850 23169 2884 23208
rect 2946 23242 2980 23281
rect 2946 23169 2980 23208
rect 3042 23242 3076 23281
rect 3042 23169 3076 23208
rect 3138 23242 3172 23281
rect 3138 23169 3172 23208
rect 3234 23242 3268 23281
rect 3234 23169 3268 23208
rect 3330 23242 3364 23281
rect 3330 23169 3364 23208
rect 3426 23242 3460 23281
rect 3426 23169 3460 23208
rect 3540 23212 3574 23245
rect 3647 23269 3681 23285
rect 3647 23177 3681 23193
rect 3735 23269 3769 23285
rect 3735 23177 3769 23193
rect 3873 23279 3907 23355
rect 5061 23284 5095 23355
rect 3873 23211 3907 23245
rect 3540 23143 3574 23177
rect 2352 23033 2386 23109
rect 2450 23097 2466 23131
rect 2500 23097 2516 23131
rect 2642 23097 2658 23131
rect 2692 23097 2708 23131
rect 2834 23097 2850 23131
rect 2884 23097 2900 23131
rect 3026 23097 3042 23131
rect 3076 23097 3092 23131
rect 3218 23097 3234 23131
rect 3268 23097 3284 23131
rect 3410 23097 3426 23131
rect 3460 23097 3476 23131
rect 3540 23033 3574 23106
rect 2352 22999 2470 23033
rect 2504 22999 2538 23033
rect 2572 22999 2606 23033
rect 2640 22999 2674 23033
rect 2708 22999 2742 23033
rect 2776 22999 2810 23033
rect 2844 22999 2878 23033
rect 2912 22999 2946 23033
rect 2980 22999 3014 23033
rect 3048 22999 3082 23033
rect 3116 22999 3150 23033
rect 3184 22999 3218 23033
rect 3252 22999 3286 23033
rect 3320 22999 3354 23033
rect 3388 22999 3422 23033
rect 3456 22999 3574 23033
rect 3873 23143 3907 23177
rect 3987 23242 4021 23281
rect 3987 23169 4021 23208
rect 4083 23242 4117 23281
rect 4083 23169 4117 23208
rect 4179 23242 4213 23281
rect 4179 23169 4213 23208
rect 4275 23242 4309 23281
rect 4275 23169 4309 23208
rect 4371 23242 4405 23281
rect 4371 23169 4405 23208
rect 4467 23242 4501 23281
rect 4467 23169 4501 23208
rect 4563 23242 4597 23281
rect 4563 23169 4597 23208
rect 4659 23242 4693 23281
rect 4659 23169 4693 23208
rect 4755 23242 4789 23281
rect 4755 23169 4789 23208
rect 4851 23242 4885 23281
rect 4851 23169 4885 23208
rect 4947 23242 4981 23281
rect 4947 23169 4981 23208
rect 5061 23212 5095 23245
rect 5340 23360 5348 23394
rect 5382 23360 5386 23394
rect 5420 23399 5486 23410
rect 5420 23396 5450 23399
rect 5420 23362 5436 23396
rect 5484 23365 5486 23399
rect 5470 23362 5486 23365
rect 5340 23324 5386 23360
rect 5340 23312 5406 23324
rect 5340 23278 5356 23312
rect 5390 23278 5406 23312
rect 5340 23244 5406 23278
rect 5340 23210 5356 23244
rect 5390 23210 5406 23244
rect 5340 23198 5406 23210
rect 5440 23312 5486 23328
rect 5474 23278 5486 23312
rect 5440 23244 5486 23278
rect 5474 23210 5486 23244
rect 5061 23143 5095 23177
rect 5440 23164 5486 23210
rect 3873 23033 3907 23109
rect 3971 23097 3987 23131
rect 4021 23097 4037 23131
rect 4163 23097 4179 23131
rect 4213 23097 4229 23131
rect 4355 23097 4371 23131
rect 4405 23097 4421 23131
rect 4547 23097 4563 23131
rect 4597 23097 4613 23131
rect 4739 23097 4755 23131
rect 4789 23097 4805 23131
rect 4931 23097 4947 23131
rect 4981 23097 4997 23131
rect 5274 23130 5303 23164
rect 5337 23130 5395 23164
rect 5429 23130 5487 23164
rect 5521 23130 5550 23164
rect 5061 23033 5095 23106
rect 3873 22999 3991 23033
rect 4025 22999 4059 23033
rect 4093 22999 4127 23033
rect 4161 22999 4195 23033
rect 4229 22999 4263 23033
rect 4297 22999 4331 23033
rect 4365 22999 4399 23033
rect 4433 22999 4467 23033
rect 4501 22999 4535 23033
rect 4569 22999 4603 23033
rect 4637 22999 4671 23033
rect 4705 22999 4739 23033
rect 4773 22999 4807 23033
rect 4841 22999 4875 23033
rect 4909 22999 4943 23033
rect 4977 22999 5095 23033
rect 199 22716 317 22750
rect 351 22716 385 22750
rect 419 22716 453 22750
rect 487 22716 521 22750
rect 555 22716 589 22750
rect 623 22716 657 22750
rect 691 22716 725 22750
rect 759 22716 793 22750
rect 827 22716 861 22750
rect 895 22716 929 22750
rect 963 22716 997 22750
rect 1031 22716 1065 22750
rect 1099 22716 1133 22750
rect 1167 22716 1201 22750
rect 1235 22716 1269 22750
rect 1303 22716 1421 22750
rect 199 22648 233 22716
rect 1387 22648 1421 22716
rect 297 22614 313 22648
rect 347 22614 363 22648
rect 489 22614 505 22648
rect 539 22614 555 22648
rect 681 22614 697 22648
rect 731 22614 747 22648
rect 873 22614 889 22648
rect 923 22614 939 22648
rect 1065 22614 1081 22648
rect 1115 22614 1131 22648
rect 1257 22614 1273 22648
rect 1307 22614 1323 22648
rect 199 22580 233 22614
rect 1387 22580 1421 22588
rect 199 22512 233 22546
rect 199 22444 233 22478
rect 199 22376 233 22410
rect 199 22308 233 22342
rect 313 22549 347 22570
rect 313 22481 347 22485
rect 313 22375 347 22379
rect 313 22290 347 22311
rect 409 22549 443 22570
rect 409 22481 443 22485
rect 409 22375 443 22379
rect 409 22290 443 22311
rect 505 22549 539 22570
rect 505 22481 539 22485
rect 505 22375 539 22379
rect 505 22290 539 22311
rect 601 22549 635 22570
rect 601 22481 635 22485
rect 601 22375 635 22379
rect 601 22290 635 22311
rect 697 22549 731 22570
rect 697 22481 731 22485
rect 697 22375 731 22379
rect 697 22290 731 22311
rect 793 22549 827 22570
rect 793 22481 827 22485
rect 793 22375 827 22379
rect 793 22290 827 22311
rect 889 22549 923 22570
rect 889 22481 923 22485
rect 889 22375 923 22379
rect 889 22290 923 22311
rect 985 22549 1019 22570
rect 985 22481 1019 22485
rect 985 22375 1019 22379
rect 985 22290 1019 22311
rect 1081 22549 1115 22570
rect 1081 22481 1115 22485
rect 1081 22375 1115 22379
rect 1081 22290 1115 22311
rect 1177 22549 1211 22570
rect 1177 22481 1211 22485
rect 1177 22375 1211 22379
rect 1177 22290 1211 22311
rect 1273 22549 1307 22570
rect 1273 22481 1307 22485
rect 1273 22375 1307 22379
rect 1273 22290 1307 22311
rect 1387 22512 1421 22516
rect 1387 22406 1421 22410
rect 1387 22334 1421 22342
rect 199 22206 233 22274
rect 1387 22206 1421 22274
rect 199 22172 317 22206
rect 351 22172 385 22206
rect 419 22172 453 22206
rect 487 22172 521 22206
rect 555 22172 589 22206
rect 623 22172 657 22206
rect 691 22172 725 22206
rect 759 22172 793 22206
rect 827 22172 861 22206
rect 895 22172 929 22206
rect 963 22172 997 22206
rect 1031 22172 1065 22206
rect 1099 22172 1133 22206
rect 1167 22172 1201 22206
rect 1235 22172 1269 22206
rect 1303 22172 1421 22206
rect 2352 22720 2470 22754
rect 2504 22720 2538 22754
rect 2572 22720 2606 22754
rect 2640 22720 2674 22754
rect 2708 22720 2742 22754
rect 2776 22720 2810 22754
rect 2844 22720 2878 22754
rect 2912 22720 2946 22754
rect 2980 22720 3014 22754
rect 3048 22720 3082 22754
rect 3116 22720 3150 22754
rect 3184 22720 3218 22754
rect 3252 22720 3286 22754
rect 3320 22720 3354 22754
rect 3388 22720 3422 22754
rect 3456 22720 3574 22754
rect 2352 22652 2386 22720
rect 3540 22652 3574 22720
rect 2450 22618 2466 22652
rect 2500 22618 2516 22652
rect 2642 22618 2658 22652
rect 2692 22618 2708 22652
rect 2834 22618 2850 22652
rect 2884 22618 2900 22652
rect 3026 22618 3042 22652
rect 3076 22618 3092 22652
rect 3218 22618 3234 22652
rect 3268 22618 3284 22652
rect 3410 22618 3426 22652
rect 3460 22618 3476 22652
rect 2352 22584 2386 22618
rect 3540 22584 3574 22592
rect 2352 22516 2386 22550
rect 2352 22448 2386 22482
rect 2352 22380 2386 22414
rect 2352 22312 2386 22346
rect 2466 22553 2500 22574
rect 2466 22485 2500 22489
rect 2466 22379 2500 22383
rect 2466 22294 2500 22315
rect 2562 22553 2596 22574
rect 2562 22485 2596 22489
rect 2562 22379 2596 22383
rect 2562 22294 2596 22315
rect 2658 22553 2692 22574
rect 2658 22485 2692 22489
rect 2658 22379 2692 22383
rect 2658 22294 2692 22315
rect 2754 22553 2788 22574
rect 2754 22485 2788 22489
rect 2754 22379 2788 22383
rect 2754 22294 2788 22315
rect 2850 22553 2884 22574
rect 2850 22485 2884 22489
rect 2850 22379 2884 22383
rect 2850 22294 2884 22315
rect 2946 22553 2980 22574
rect 2946 22485 2980 22489
rect 2946 22379 2980 22383
rect 2946 22294 2980 22315
rect 3042 22553 3076 22574
rect 3042 22485 3076 22489
rect 3042 22379 3076 22383
rect 3042 22294 3076 22315
rect 3138 22553 3172 22574
rect 3138 22485 3172 22489
rect 3138 22379 3172 22383
rect 3138 22294 3172 22315
rect 3234 22553 3268 22574
rect 3234 22485 3268 22489
rect 3234 22379 3268 22383
rect 3234 22294 3268 22315
rect 3330 22553 3364 22574
rect 3330 22485 3364 22489
rect 3330 22379 3364 22383
rect 3330 22294 3364 22315
rect 3426 22553 3460 22574
rect 3426 22485 3460 22489
rect 3426 22379 3460 22383
rect 3426 22294 3460 22315
rect 3540 22516 3574 22520
rect 3540 22410 3574 22414
rect 3540 22338 3574 22346
rect 2352 22210 2386 22278
rect 3540 22210 3574 22278
rect 2352 22176 2470 22210
rect 2504 22176 2538 22210
rect 2572 22176 2606 22210
rect 2640 22176 2674 22210
rect 2708 22176 2742 22210
rect 2776 22176 2810 22210
rect 2844 22176 2878 22210
rect 2912 22176 2946 22210
rect 2980 22176 3014 22210
rect 3048 22176 3082 22210
rect 3116 22176 3150 22210
rect 3184 22176 3218 22210
rect 3252 22176 3286 22210
rect 3320 22176 3354 22210
rect 3388 22176 3422 22210
rect 3456 22176 3574 22210
rect 3873 22720 3991 22754
rect 4025 22720 4059 22754
rect 4093 22720 4127 22754
rect 4161 22720 4195 22754
rect 4229 22720 4263 22754
rect 4297 22720 4331 22754
rect 4365 22720 4399 22754
rect 4433 22720 4467 22754
rect 4501 22720 4535 22754
rect 4569 22720 4603 22754
rect 4637 22720 4671 22754
rect 4705 22720 4739 22754
rect 4773 22720 4807 22754
rect 4841 22720 4875 22754
rect 4909 22720 4943 22754
rect 4977 22720 5095 22754
rect 3873 22652 3907 22720
rect 5061 22652 5095 22720
rect 3971 22618 3987 22652
rect 4021 22618 4037 22652
rect 4163 22618 4179 22652
rect 4213 22618 4229 22652
rect 4355 22618 4371 22652
rect 4405 22618 4421 22652
rect 4547 22618 4563 22652
rect 4597 22618 4613 22652
rect 4739 22618 4755 22652
rect 4789 22618 4805 22652
rect 4931 22618 4947 22652
rect 4981 22618 4997 22652
rect 3873 22584 3907 22618
rect 5061 22584 5095 22592
rect 3873 22516 3907 22550
rect 3873 22448 3907 22482
rect 3873 22380 3907 22414
rect 3873 22312 3907 22346
rect 3987 22553 4021 22574
rect 3987 22485 4021 22489
rect 3987 22379 4021 22383
rect 3987 22294 4021 22315
rect 4083 22553 4117 22574
rect 4083 22485 4117 22489
rect 4083 22379 4117 22383
rect 4083 22294 4117 22315
rect 4179 22553 4213 22574
rect 4179 22485 4213 22489
rect 4179 22379 4213 22383
rect 4179 22294 4213 22315
rect 4275 22553 4309 22574
rect 4275 22485 4309 22489
rect 4275 22379 4309 22383
rect 4275 22294 4309 22315
rect 4371 22553 4405 22574
rect 4371 22485 4405 22489
rect 4371 22379 4405 22383
rect 4371 22294 4405 22315
rect 4467 22553 4501 22574
rect 4467 22485 4501 22489
rect 4467 22379 4501 22383
rect 4467 22294 4501 22315
rect 4563 22553 4597 22574
rect 4563 22485 4597 22489
rect 4563 22379 4597 22383
rect 4563 22294 4597 22315
rect 4659 22553 4693 22574
rect 4659 22485 4693 22489
rect 4659 22379 4693 22383
rect 4659 22294 4693 22315
rect 4755 22553 4789 22574
rect 4755 22485 4789 22489
rect 4755 22379 4789 22383
rect 4755 22294 4789 22315
rect 4851 22553 4885 22574
rect 4851 22485 4885 22489
rect 4851 22379 4885 22383
rect 4851 22294 4885 22315
rect 4947 22553 4981 22574
rect 4947 22485 4981 22489
rect 4947 22379 4981 22383
rect 4947 22294 4981 22315
rect 5061 22516 5095 22520
rect 5061 22410 5095 22414
rect 5274 22387 5303 22421
rect 5337 22387 5395 22421
rect 5429 22387 5487 22421
rect 5521 22387 5550 22421
rect 5061 22338 5095 22346
rect 3873 22210 3907 22278
rect 5061 22210 5095 22278
rect 3873 22176 3991 22210
rect 4025 22176 4059 22210
rect 4093 22176 4127 22210
rect 4161 22176 4195 22210
rect 4229 22176 4263 22210
rect 4297 22176 4331 22210
rect 4365 22176 4399 22210
rect 4433 22176 4467 22210
rect 4501 22176 4535 22210
rect 4569 22176 4603 22210
rect 4637 22176 4671 22210
rect 4705 22176 4739 22210
rect 4773 22176 4807 22210
rect 4841 22176 4875 22210
rect 4909 22176 4943 22210
rect 4977 22176 5095 22210
rect 5340 22345 5406 22353
rect 5340 22311 5356 22345
rect 5390 22311 5406 22345
rect 5340 22277 5406 22311
rect 5340 22243 5356 22277
rect 5390 22243 5406 22277
rect 5340 22209 5406 22243
rect 5340 22175 5356 22209
rect 5390 22175 5406 22209
rect 5340 22157 5406 22175
rect 5440 22345 5482 22387
rect 5474 22311 5482 22345
rect 5440 22277 5482 22311
rect 5474 22243 5482 22277
rect 5440 22209 5482 22243
rect 5474 22175 5482 22209
rect 5440 22159 5482 22175
rect 5340 22107 5386 22157
rect 199 22064 317 22098
rect 351 22064 385 22098
rect 419 22064 453 22098
rect 487 22064 521 22098
rect 555 22064 589 22098
rect 623 22064 657 22098
rect 691 22064 725 22098
rect 759 22064 793 22098
rect 827 22064 861 22098
rect 895 22064 929 22098
rect 963 22064 997 22098
rect 1031 22064 1065 22098
rect 1099 22064 1133 22098
rect 1167 22064 1201 22098
rect 1235 22064 1269 22098
rect 1303 22064 1421 22098
rect 199 21988 233 22064
rect 1387 21993 1421 22064
rect 199 21920 233 21954
rect 199 21852 233 21886
rect 313 21951 347 21990
rect 313 21878 347 21917
rect 409 21951 443 21990
rect 409 21878 443 21917
rect 505 21951 539 21990
rect 505 21878 539 21917
rect 601 21951 635 21990
rect 601 21878 635 21917
rect 697 21951 731 21990
rect 697 21878 731 21917
rect 793 21951 827 21990
rect 793 21878 827 21917
rect 889 21951 923 21990
rect 889 21878 923 21917
rect 985 21951 1019 21990
rect 985 21878 1019 21917
rect 1081 21951 1115 21990
rect 1081 21878 1115 21917
rect 1177 21951 1211 21990
rect 1177 21878 1211 21917
rect 1273 21951 1307 21990
rect 1273 21878 1307 21917
rect 1387 21921 1421 21954
rect 1387 21852 1421 21886
rect 199 21742 233 21818
rect 297 21806 313 21840
rect 347 21806 363 21840
rect 489 21806 505 21840
rect 539 21806 555 21840
rect 681 21806 697 21840
rect 731 21806 747 21840
rect 873 21806 889 21840
rect 923 21806 939 21840
rect 1065 21806 1081 21840
rect 1115 21806 1131 21840
rect 1257 21806 1273 21840
rect 1307 21806 1323 21840
rect 1387 21742 1421 21815
rect 199 21708 317 21742
rect 351 21708 385 21742
rect 419 21708 453 21742
rect 487 21708 521 21742
rect 555 21708 589 21742
rect 623 21708 657 21742
rect 691 21708 725 21742
rect 759 21708 793 21742
rect 827 21708 861 21742
rect 895 21708 929 21742
rect 963 21708 997 21742
rect 1031 21708 1065 21742
rect 1099 21708 1133 21742
rect 1167 21708 1201 21742
rect 1235 21708 1269 21742
rect 1303 21708 1421 21742
rect 2352 22068 2470 22102
rect 2504 22068 2538 22102
rect 2572 22068 2606 22102
rect 2640 22068 2674 22102
rect 2708 22068 2742 22102
rect 2776 22068 2810 22102
rect 2844 22068 2878 22102
rect 2912 22068 2946 22102
rect 2980 22068 3014 22102
rect 3048 22068 3082 22102
rect 3116 22068 3150 22102
rect 3184 22068 3218 22102
rect 3252 22068 3286 22102
rect 3320 22068 3354 22102
rect 3388 22068 3422 22102
rect 3456 22068 3574 22102
rect 2352 21992 2386 22068
rect 3540 21997 3574 22068
rect 3873 22068 3991 22102
rect 4025 22068 4059 22102
rect 4093 22068 4127 22102
rect 4161 22068 4195 22102
rect 4229 22068 4263 22102
rect 4297 22068 4331 22102
rect 4365 22068 4399 22102
rect 4433 22068 4467 22102
rect 4501 22068 4535 22102
rect 4569 22068 4603 22102
rect 4637 22068 4671 22102
rect 4705 22068 4739 22102
rect 4773 22068 4807 22102
rect 4841 22068 4875 22102
rect 4909 22068 4943 22102
rect 4977 22068 5095 22102
rect 3675 22032 3691 22066
rect 3725 22032 3741 22066
rect 2352 21924 2386 21958
rect 2352 21856 2386 21890
rect 2466 21955 2500 21994
rect 2466 21882 2500 21921
rect 2562 21955 2596 21994
rect 2562 21882 2596 21921
rect 2658 21955 2692 21994
rect 2658 21882 2692 21921
rect 2754 21955 2788 21994
rect 2754 21882 2788 21921
rect 2850 21955 2884 21994
rect 2850 21882 2884 21921
rect 2946 21955 2980 21994
rect 2946 21882 2980 21921
rect 3042 21955 3076 21994
rect 3042 21882 3076 21921
rect 3138 21955 3172 21994
rect 3138 21882 3172 21921
rect 3234 21955 3268 21994
rect 3234 21882 3268 21921
rect 3330 21955 3364 21994
rect 3330 21882 3364 21921
rect 3426 21955 3460 21994
rect 3426 21882 3460 21921
rect 3540 21925 3574 21958
rect 3647 21982 3681 21998
rect 3647 21890 3681 21906
rect 3735 21982 3769 21998
rect 3735 21890 3769 21906
rect 3873 21992 3907 22068
rect 5061 21997 5095 22068
rect 3873 21924 3907 21958
rect 3540 21856 3574 21890
rect 2352 21746 2386 21822
rect 2450 21810 2466 21844
rect 2500 21810 2516 21844
rect 2642 21810 2658 21844
rect 2692 21810 2708 21844
rect 2834 21810 2850 21844
rect 2884 21810 2900 21844
rect 3026 21810 3042 21844
rect 3076 21810 3092 21844
rect 3218 21810 3234 21844
rect 3268 21810 3284 21844
rect 3410 21810 3426 21844
rect 3460 21810 3476 21844
rect 3540 21746 3574 21819
rect 2352 21712 2470 21746
rect 2504 21712 2538 21746
rect 2572 21712 2606 21746
rect 2640 21712 2674 21746
rect 2708 21712 2742 21746
rect 2776 21712 2810 21746
rect 2844 21712 2878 21746
rect 2912 21712 2946 21746
rect 2980 21712 3014 21746
rect 3048 21712 3082 21746
rect 3116 21712 3150 21746
rect 3184 21712 3218 21746
rect 3252 21712 3286 21746
rect 3320 21712 3354 21746
rect 3388 21712 3422 21746
rect 3456 21712 3574 21746
rect 3873 21856 3907 21890
rect 3987 21955 4021 21994
rect 3987 21882 4021 21921
rect 4083 21955 4117 21994
rect 4083 21882 4117 21921
rect 4179 21955 4213 21994
rect 4179 21882 4213 21921
rect 4275 21955 4309 21994
rect 4275 21882 4309 21921
rect 4371 21955 4405 21994
rect 4371 21882 4405 21921
rect 4467 21955 4501 21994
rect 4467 21882 4501 21921
rect 4563 21955 4597 21994
rect 4563 21882 4597 21921
rect 4659 21955 4693 21994
rect 4659 21882 4693 21921
rect 4755 21955 4789 21994
rect 4755 21882 4789 21921
rect 4851 21955 4885 21994
rect 4851 21882 4885 21921
rect 4947 21955 4981 21994
rect 4947 21882 4981 21921
rect 5061 21925 5095 21958
rect 5340 22073 5348 22107
rect 5382 22073 5386 22107
rect 5420 22112 5486 22123
rect 5420 22109 5450 22112
rect 5420 22075 5436 22109
rect 5484 22078 5486 22112
rect 5470 22075 5486 22078
rect 5340 22037 5386 22073
rect 5340 22025 5406 22037
rect 5340 21991 5356 22025
rect 5390 21991 5406 22025
rect 5340 21957 5406 21991
rect 5340 21923 5356 21957
rect 5390 21923 5406 21957
rect 5340 21911 5406 21923
rect 5440 22025 5486 22041
rect 5474 21991 5486 22025
rect 5440 21957 5486 21991
rect 5474 21923 5486 21957
rect 5061 21856 5095 21890
rect 5440 21877 5486 21923
rect 3873 21746 3907 21822
rect 3971 21810 3987 21844
rect 4021 21810 4037 21844
rect 4163 21810 4179 21844
rect 4213 21810 4229 21844
rect 4355 21810 4371 21844
rect 4405 21810 4421 21844
rect 4547 21810 4563 21844
rect 4597 21810 4613 21844
rect 4739 21810 4755 21844
rect 4789 21810 4805 21844
rect 4931 21810 4947 21844
rect 4981 21810 4997 21844
rect 5274 21843 5303 21877
rect 5337 21843 5395 21877
rect 5429 21843 5487 21877
rect 5521 21843 5550 21877
rect 5061 21746 5095 21819
rect 3873 21712 3991 21746
rect 4025 21712 4059 21746
rect 4093 21712 4127 21746
rect 4161 21712 4195 21746
rect 4229 21712 4263 21746
rect 4297 21712 4331 21746
rect 4365 21712 4399 21746
rect 4433 21712 4467 21746
rect 4501 21712 4535 21746
rect 4569 21712 4603 21746
rect 4637 21712 4671 21746
rect 4705 21712 4739 21746
rect 4773 21712 4807 21746
rect 4841 21712 4875 21746
rect 4909 21712 4943 21746
rect 4977 21712 5095 21746
rect 199 21429 317 21463
rect 351 21429 385 21463
rect 419 21429 453 21463
rect 487 21429 521 21463
rect 555 21429 589 21463
rect 623 21429 657 21463
rect 691 21429 725 21463
rect 759 21429 793 21463
rect 827 21429 861 21463
rect 895 21429 929 21463
rect 963 21429 997 21463
rect 1031 21429 1065 21463
rect 1099 21429 1133 21463
rect 1167 21429 1201 21463
rect 1235 21429 1269 21463
rect 1303 21429 1421 21463
rect 199 21361 233 21429
rect 1387 21361 1421 21429
rect 297 21327 313 21361
rect 347 21327 363 21361
rect 489 21327 505 21361
rect 539 21327 555 21361
rect 681 21327 697 21361
rect 731 21327 747 21361
rect 873 21327 889 21361
rect 923 21327 939 21361
rect 1065 21327 1081 21361
rect 1115 21327 1131 21361
rect 1257 21327 1273 21361
rect 1307 21327 1323 21361
rect 199 21293 233 21327
rect 1387 21293 1421 21301
rect 199 21225 233 21259
rect 199 21157 233 21191
rect 199 21089 233 21123
rect 199 21021 233 21055
rect 313 21262 347 21283
rect 313 21194 347 21198
rect 313 21088 347 21092
rect 313 21003 347 21024
rect 409 21262 443 21283
rect 409 21194 443 21198
rect 409 21088 443 21092
rect 409 21003 443 21024
rect 505 21262 539 21283
rect 505 21194 539 21198
rect 505 21088 539 21092
rect 505 21003 539 21024
rect 601 21262 635 21283
rect 601 21194 635 21198
rect 601 21088 635 21092
rect 601 21003 635 21024
rect 697 21262 731 21283
rect 697 21194 731 21198
rect 697 21088 731 21092
rect 697 21003 731 21024
rect 793 21262 827 21283
rect 793 21194 827 21198
rect 793 21088 827 21092
rect 793 21003 827 21024
rect 889 21262 923 21283
rect 889 21194 923 21198
rect 889 21088 923 21092
rect 889 21003 923 21024
rect 985 21262 1019 21283
rect 985 21194 1019 21198
rect 985 21088 1019 21092
rect 985 21003 1019 21024
rect 1081 21262 1115 21283
rect 1081 21194 1115 21198
rect 1081 21088 1115 21092
rect 1081 21003 1115 21024
rect 1177 21262 1211 21283
rect 1177 21194 1211 21198
rect 1177 21088 1211 21092
rect 1177 21003 1211 21024
rect 1273 21262 1307 21283
rect 1273 21194 1307 21198
rect 1273 21088 1307 21092
rect 1273 21003 1307 21024
rect 1387 21225 1421 21229
rect 1387 21119 1421 21123
rect 1387 21047 1421 21055
rect 199 20919 233 20987
rect 1387 20919 1421 20987
rect 199 20885 317 20919
rect 351 20885 385 20919
rect 419 20885 453 20919
rect 487 20885 521 20919
rect 555 20885 589 20919
rect 623 20885 657 20919
rect 691 20885 725 20919
rect 759 20885 793 20919
rect 827 20885 861 20919
rect 895 20885 929 20919
rect 963 20885 997 20919
rect 1031 20885 1065 20919
rect 1099 20885 1133 20919
rect 1167 20885 1201 20919
rect 1235 20885 1269 20919
rect 1303 20885 1421 20919
rect 2352 21433 2470 21467
rect 2504 21433 2538 21467
rect 2572 21433 2606 21467
rect 2640 21433 2674 21467
rect 2708 21433 2742 21467
rect 2776 21433 2810 21467
rect 2844 21433 2878 21467
rect 2912 21433 2946 21467
rect 2980 21433 3014 21467
rect 3048 21433 3082 21467
rect 3116 21433 3150 21467
rect 3184 21433 3218 21467
rect 3252 21433 3286 21467
rect 3320 21433 3354 21467
rect 3388 21433 3422 21467
rect 3456 21433 3574 21467
rect 2352 21365 2386 21433
rect 3540 21365 3574 21433
rect 2450 21331 2466 21365
rect 2500 21331 2516 21365
rect 2642 21331 2658 21365
rect 2692 21331 2708 21365
rect 2834 21331 2850 21365
rect 2884 21331 2900 21365
rect 3026 21331 3042 21365
rect 3076 21331 3092 21365
rect 3218 21331 3234 21365
rect 3268 21331 3284 21365
rect 3410 21331 3426 21365
rect 3460 21331 3476 21365
rect 2352 21297 2386 21331
rect 3540 21297 3574 21305
rect 2352 21229 2386 21263
rect 2352 21161 2386 21195
rect 2352 21093 2386 21127
rect 2352 21025 2386 21059
rect 2466 21266 2500 21287
rect 2466 21198 2500 21202
rect 2466 21092 2500 21096
rect 2466 21007 2500 21028
rect 2562 21266 2596 21287
rect 2562 21198 2596 21202
rect 2562 21092 2596 21096
rect 2562 21007 2596 21028
rect 2658 21266 2692 21287
rect 2658 21198 2692 21202
rect 2658 21092 2692 21096
rect 2658 21007 2692 21028
rect 2754 21266 2788 21287
rect 2754 21198 2788 21202
rect 2754 21092 2788 21096
rect 2754 21007 2788 21028
rect 2850 21266 2884 21287
rect 2850 21198 2884 21202
rect 2850 21092 2884 21096
rect 2850 21007 2884 21028
rect 2946 21266 2980 21287
rect 2946 21198 2980 21202
rect 2946 21092 2980 21096
rect 2946 21007 2980 21028
rect 3042 21266 3076 21287
rect 3042 21198 3076 21202
rect 3042 21092 3076 21096
rect 3042 21007 3076 21028
rect 3138 21266 3172 21287
rect 3138 21198 3172 21202
rect 3138 21092 3172 21096
rect 3138 21007 3172 21028
rect 3234 21266 3268 21287
rect 3234 21198 3268 21202
rect 3234 21092 3268 21096
rect 3234 21007 3268 21028
rect 3330 21266 3364 21287
rect 3330 21198 3364 21202
rect 3330 21092 3364 21096
rect 3330 21007 3364 21028
rect 3426 21266 3460 21287
rect 3426 21198 3460 21202
rect 3426 21092 3460 21096
rect 3426 21007 3460 21028
rect 3540 21229 3574 21233
rect 3540 21123 3574 21127
rect 3540 21051 3574 21059
rect 2352 20923 2386 20991
rect 3540 20923 3574 20991
rect 2352 20889 2470 20923
rect 2504 20889 2538 20923
rect 2572 20889 2606 20923
rect 2640 20889 2674 20923
rect 2708 20889 2742 20923
rect 2776 20889 2810 20923
rect 2844 20889 2878 20923
rect 2912 20889 2946 20923
rect 2980 20889 3014 20923
rect 3048 20889 3082 20923
rect 3116 20889 3150 20923
rect 3184 20889 3218 20923
rect 3252 20889 3286 20923
rect 3320 20889 3354 20923
rect 3388 20889 3422 20923
rect 3456 20889 3574 20923
rect 3873 21433 3991 21467
rect 4025 21433 4059 21467
rect 4093 21433 4127 21467
rect 4161 21433 4195 21467
rect 4229 21433 4263 21467
rect 4297 21433 4331 21467
rect 4365 21433 4399 21467
rect 4433 21433 4467 21467
rect 4501 21433 4535 21467
rect 4569 21433 4603 21467
rect 4637 21433 4671 21467
rect 4705 21433 4739 21467
rect 4773 21433 4807 21467
rect 4841 21433 4875 21467
rect 4909 21433 4943 21467
rect 4977 21433 5095 21467
rect 3873 21365 3907 21433
rect 5061 21365 5095 21433
rect 3971 21331 3987 21365
rect 4021 21331 4037 21365
rect 4163 21331 4179 21365
rect 4213 21331 4229 21365
rect 4355 21331 4371 21365
rect 4405 21331 4421 21365
rect 4547 21331 4563 21365
rect 4597 21331 4613 21365
rect 4739 21331 4755 21365
rect 4789 21331 4805 21365
rect 4931 21331 4947 21365
rect 4981 21331 4997 21365
rect 3873 21297 3907 21331
rect 5061 21297 5095 21305
rect 3873 21229 3907 21263
rect 3873 21161 3907 21195
rect 3873 21093 3907 21127
rect 3873 21025 3907 21059
rect 3987 21266 4021 21287
rect 3987 21198 4021 21202
rect 3987 21092 4021 21096
rect 3987 21007 4021 21028
rect 4083 21266 4117 21287
rect 4083 21198 4117 21202
rect 4083 21092 4117 21096
rect 4083 21007 4117 21028
rect 4179 21266 4213 21287
rect 4179 21198 4213 21202
rect 4179 21092 4213 21096
rect 4179 21007 4213 21028
rect 4275 21266 4309 21287
rect 4275 21198 4309 21202
rect 4275 21092 4309 21096
rect 4275 21007 4309 21028
rect 4371 21266 4405 21287
rect 4371 21198 4405 21202
rect 4371 21092 4405 21096
rect 4371 21007 4405 21028
rect 4467 21266 4501 21287
rect 4467 21198 4501 21202
rect 4467 21092 4501 21096
rect 4467 21007 4501 21028
rect 4563 21266 4597 21287
rect 4563 21198 4597 21202
rect 4563 21092 4597 21096
rect 4563 21007 4597 21028
rect 4659 21266 4693 21287
rect 4659 21198 4693 21202
rect 4659 21092 4693 21096
rect 4659 21007 4693 21028
rect 4755 21266 4789 21287
rect 4755 21198 4789 21202
rect 4755 21092 4789 21096
rect 4755 21007 4789 21028
rect 4851 21266 4885 21287
rect 4851 21198 4885 21202
rect 4851 21092 4885 21096
rect 4851 21007 4885 21028
rect 4947 21266 4981 21287
rect 4947 21198 4981 21202
rect 4947 21092 4981 21096
rect 4947 21007 4981 21028
rect 5061 21229 5095 21233
rect 5061 21123 5095 21127
rect 5274 21100 5303 21134
rect 5337 21100 5395 21134
rect 5429 21100 5487 21134
rect 5521 21100 5550 21134
rect 5061 21051 5095 21059
rect 3873 20923 3907 20991
rect 5061 20923 5095 20991
rect 3873 20889 3991 20923
rect 4025 20889 4059 20923
rect 4093 20889 4127 20923
rect 4161 20889 4195 20923
rect 4229 20889 4263 20923
rect 4297 20889 4331 20923
rect 4365 20889 4399 20923
rect 4433 20889 4467 20923
rect 4501 20889 4535 20923
rect 4569 20889 4603 20923
rect 4637 20889 4671 20923
rect 4705 20889 4739 20923
rect 4773 20889 4807 20923
rect 4841 20889 4875 20923
rect 4909 20889 4943 20923
rect 4977 20889 5095 20923
rect 5340 21058 5406 21066
rect 5340 21024 5356 21058
rect 5390 21024 5406 21058
rect 5340 20990 5406 21024
rect 5340 20956 5356 20990
rect 5390 20956 5406 20990
rect 5340 20922 5406 20956
rect 5340 20888 5356 20922
rect 5390 20888 5406 20922
rect 5340 20870 5406 20888
rect 5440 21058 5482 21100
rect 5474 21024 5482 21058
rect 5440 20990 5482 21024
rect 5474 20956 5482 20990
rect 5440 20922 5482 20956
rect 5474 20888 5482 20922
rect 5440 20872 5482 20888
rect 5340 20820 5386 20870
rect 199 20777 317 20811
rect 351 20777 385 20811
rect 419 20777 453 20811
rect 487 20777 521 20811
rect 555 20777 589 20811
rect 623 20777 657 20811
rect 691 20777 725 20811
rect 759 20777 793 20811
rect 827 20777 861 20811
rect 895 20777 929 20811
rect 963 20777 997 20811
rect 1031 20777 1065 20811
rect 1099 20777 1133 20811
rect 1167 20777 1201 20811
rect 1235 20777 1269 20811
rect 1303 20777 1421 20811
rect 199 20701 233 20777
rect 1387 20706 1421 20777
rect 199 20633 233 20667
rect 199 20565 233 20599
rect 313 20664 347 20703
rect 313 20591 347 20630
rect 409 20664 443 20703
rect 409 20591 443 20630
rect 505 20664 539 20703
rect 505 20591 539 20630
rect 601 20664 635 20703
rect 601 20591 635 20630
rect 697 20664 731 20703
rect 697 20591 731 20630
rect 793 20664 827 20703
rect 793 20591 827 20630
rect 889 20664 923 20703
rect 889 20591 923 20630
rect 985 20664 1019 20703
rect 985 20591 1019 20630
rect 1081 20664 1115 20703
rect 1081 20591 1115 20630
rect 1177 20664 1211 20703
rect 1177 20591 1211 20630
rect 1273 20664 1307 20703
rect 1273 20591 1307 20630
rect 1387 20634 1421 20667
rect 1387 20565 1421 20599
rect 199 20455 233 20531
rect 297 20519 313 20553
rect 347 20519 363 20553
rect 489 20519 505 20553
rect 539 20519 555 20553
rect 681 20519 697 20553
rect 731 20519 747 20553
rect 873 20519 889 20553
rect 923 20519 939 20553
rect 1065 20519 1081 20553
rect 1115 20519 1131 20553
rect 1257 20519 1273 20553
rect 1307 20519 1323 20553
rect 1387 20455 1421 20528
rect 199 20421 317 20455
rect 351 20421 385 20455
rect 419 20421 453 20455
rect 487 20421 521 20455
rect 555 20421 589 20455
rect 623 20421 657 20455
rect 691 20421 725 20455
rect 759 20421 793 20455
rect 827 20421 861 20455
rect 895 20421 929 20455
rect 963 20421 997 20455
rect 1031 20421 1065 20455
rect 1099 20421 1133 20455
rect 1167 20421 1201 20455
rect 1235 20421 1269 20455
rect 1303 20421 1421 20455
rect 2352 20781 2470 20815
rect 2504 20781 2538 20815
rect 2572 20781 2606 20815
rect 2640 20781 2674 20815
rect 2708 20781 2742 20815
rect 2776 20781 2810 20815
rect 2844 20781 2878 20815
rect 2912 20781 2946 20815
rect 2980 20781 3014 20815
rect 3048 20781 3082 20815
rect 3116 20781 3150 20815
rect 3184 20781 3218 20815
rect 3252 20781 3286 20815
rect 3320 20781 3354 20815
rect 3388 20781 3422 20815
rect 3456 20781 3574 20815
rect 2352 20705 2386 20781
rect 3540 20710 3574 20781
rect 3873 20781 3991 20815
rect 4025 20781 4059 20815
rect 4093 20781 4127 20815
rect 4161 20781 4195 20815
rect 4229 20781 4263 20815
rect 4297 20781 4331 20815
rect 4365 20781 4399 20815
rect 4433 20781 4467 20815
rect 4501 20781 4535 20815
rect 4569 20781 4603 20815
rect 4637 20781 4671 20815
rect 4705 20781 4739 20815
rect 4773 20781 4807 20815
rect 4841 20781 4875 20815
rect 4909 20781 4943 20815
rect 4977 20781 5095 20815
rect 3675 20745 3691 20779
rect 3725 20745 3741 20779
rect 2352 20637 2386 20671
rect 2352 20569 2386 20603
rect 2466 20668 2500 20707
rect 2466 20595 2500 20634
rect 2562 20668 2596 20707
rect 2562 20595 2596 20634
rect 2658 20668 2692 20707
rect 2658 20595 2692 20634
rect 2754 20668 2788 20707
rect 2754 20595 2788 20634
rect 2850 20668 2884 20707
rect 2850 20595 2884 20634
rect 2946 20668 2980 20707
rect 2946 20595 2980 20634
rect 3042 20668 3076 20707
rect 3042 20595 3076 20634
rect 3138 20668 3172 20707
rect 3138 20595 3172 20634
rect 3234 20668 3268 20707
rect 3234 20595 3268 20634
rect 3330 20668 3364 20707
rect 3330 20595 3364 20634
rect 3426 20668 3460 20707
rect 3426 20595 3460 20634
rect 3540 20638 3574 20671
rect 3647 20695 3681 20711
rect 3647 20603 3681 20619
rect 3735 20695 3769 20711
rect 3735 20603 3769 20619
rect 3873 20705 3907 20781
rect 5061 20710 5095 20781
rect 3873 20637 3907 20671
rect 3540 20569 3574 20603
rect 2352 20459 2386 20535
rect 2450 20523 2466 20557
rect 2500 20523 2516 20557
rect 2642 20523 2658 20557
rect 2692 20523 2708 20557
rect 2834 20523 2850 20557
rect 2884 20523 2900 20557
rect 3026 20523 3042 20557
rect 3076 20523 3092 20557
rect 3218 20523 3234 20557
rect 3268 20523 3284 20557
rect 3410 20523 3426 20557
rect 3460 20523 3476 20557
rect 3540 20459 3574 20532
rect 2352 20425 2470 20459
rect 2504 20425 2538 20459
rect 2572 20425 2606 20459
rect 2640 20425 2674 20459
rect 2708 20425 2742 20459
rect 2776 20425 2810 20459
rect 2844 20425 2878 20459
rect 2912 20425 2946 20459
rect 2980 20425 3014 20459
rect 3048 20425 3082 20459
rect 3116 20425 3150 20459
rect 3184 20425 3218 20459
rect 3252 20425 3286 20459
rect 3320 20425 3354 20459
rect 3388 20425 3422 20459
rect 3456 20425 3574 20459
rect 3873 20569 3907 20603
rect 3987 20668 4021 20707
rect 3987 20595 4021 20634
rect 4083 20668 4117 20707
rect 4083 20595 4117 20634
rect 4179 20668 4213 20707
rect 4179 20595 4213 20634
rect 4275 20668 4309 20707
rect 4275 20595 4309 20634
rect 4371 20668 4405 20707
rect 4371 20595 4405 20634
rect 4467 20668 4501 20707
rect 4467 20595 4501 20634
rect 4563 20668 4597 20707
rect 4563 20595 4597 20634
rect 4659 20668 4693 20707
rect 4659 20595 4693 20634
rect 4755 20668 4789 20707
rect 4755 20595 4789 20634
rect 4851 20668 4885 20707
rect 4851 20595 4885 20634
rect 4947 20668 4981 20707
rect 4947 20595 4981 20634
rect 5061 20638 5095 20671
rect 5340 20786 5348 20820
rect 5382 20786 5386 20820
rect 5420 20825 5486 20836
rect 5420 20822 5450 20825
rect 5420 20788 5436 20822
rect 5484 20791 5486 20825
rect 5470 20788 5486 20791
rect 5340 20750 5386 20786
rect 5340 20738 5406 20750
rect 5340 20704 5356 20738
rect 5390 20704 5406 20738
rect 5340 20670 5406 20704
rect 5340 20636 5356 20670
rect 5390 20636 5406 20670
rect 5340 20624 5406 20636
rect 5440 20738 5486 20754
rect 5474 20704 5486 20738
rect 5440 20670 5486 20704
rect 5474 20636 5486 20670
rect 5061 20569 5095 20603
rect 5440 20590 5486 20636
rect 3873 20459 3907 20535
rect 3971 20523 3987 20557
rect 4021 20523 4037 20557
rect 4163 20523 4179 20557
rect 4213 20523 4229 20557
rect 4355 20523 4371 20557
rect 4405 20523 4421 20557
rect 4547 20523 4563 20557
rect 4597 20523 4613 20557
rect 4739 20523 4755 20557
rect 4789 20523 4805 20557
rect 4931 20523 4947 20557
rect 4981 20523 4997 20557
rect 5274 20556 5303 20590
rect 5337 20556 5395 20590
rect 5429 20556 5487 20590
rect 5521 20556 5550 20590
rect 5061 20459 5095 20532
rect 3873 20425 3991 20459
rect 4025 20425 4059 20459
rect 4093 20425 4127 20459
rect 4161 20425 4195 20459
rect 4229 20425 4263 20459
rect 4297 20425 4331 20459
rect 4365 20425 4399 20459
rect 4433 20425 4467 20459
rect 4501 20425 4535 20459
rect 4569 20425 4603 20459
rect 4637 20425 4671 20459
rect 4705 20425 4739 20459
rect 4773 20425 4807 20459
rect 4841 20425 4875 20459
rect 4909 20425 4943 20459
rect 4977 20425 5095 20459
rect 199 20142 317 20176
rect 351 20142 385 20176
rect 419 20142 453 20176
rect 487 20142 521 20176
rect 555 20142 589 20176
rect 623 20142 657 20176
rect 691 20142 725 20176
rect 759 20142 793 20176
rect 827 20142 861 20176
rect 895 20142 929 20176
rect 963 20142 997 20176
rect 1031 20142 1065 20176
rect 1099 20142 1133 20176
rect 1167 20142 1201 20176
rect 1235 20142 1269 20176
rect 1303 20142 1421 20176
rect 199 20074 233 20142
rect 1387 20074 1421 20142
rect 297 20040 313 20074
rect 347 20040 363 20074
rect 489 20040 505 20074
rect 539 20040 555 20074
rect 681 20040 697 20074
rect 731 20040 747 20074
rect 873 20040 889 20074
rect 923 20040 939 20074
rect 1065 20040 1081 20074
rect 1115 20040 1131 20074
rect 1257 20040 1273 20074
rect 1307 20040 1323 20074
rect 199 20006 233 20040
rect 1387 20006 1421 20014
rect 199 19938 233 19972
rect 199 19870 233 19904
rect 199 19802 233 19836
rect 199 19734 233 19768
rect 313 19975 347 19996
rect 313 19907 347 19911
rect 313 19801 347 19805
rect 313 19716 347 19737
rect 409 19975 443 19996
rect 409 19907 443 19911
rect 409 19801 443 19805
rect 409 19716 443 19737
rect 505 19975 539 19996
rect 505 19907 539 19911
rect 505 19801 539 19805
rect 505 19716 539 19737
rect 601 19975 635 19996
rect 601 19907 635 19911
rect 601 19801 635 19805
rect 601 19716 635 19737
rect 697 19975 731 19996
rect 697 19907 731 19911
rect 697 19801 731 19805
rect 697 19716 731 19737
rect 793 19975 827 19996
rect 793 19907 827 19911
rect 793 19801 827 19805
rect 793 19716 827 19737
rect 889 19975 923 19996
rect 889 19907 923 19911
rect 889 19801 923 19805
rect 889 19716 923 19737
rect 985 19975 1019 19996
rect 985 19907 1019 19911
rect 985 19801 1019 19805
rect 985 19716 1019 19737
rect 1081 19975 1115 19996
rect 1081 19907 1115 19911
rect 1081 19801 1115 19805
rect 1081 19716 1115 19737
rect 1177 19975 1211 19996
rect 1177 19907 1211 19911
rect 1177 19801 1211 19805
rect 1177 19716 1211 19737
rect 1273 19975 1307 19996
rect 1273 19907 1307 19911
rect 1273 19801 1307 19805
rect 1273 19716 1307 19737
rect 1387 19938 1421 19942
rect 1387 19832 1421 19836
rect 1387 19760 1421 19768
rect 199 19632 233 19700
rect 1387 19632 1421 19700
rect 199 19598 317 19632
rect 351 19598 385 19632
rect 419 19598 453 19632
rect 487 19598 521 19632
rect 555 19598 589 19632
rect 623 19598 657 19632
rect 691 19598 725 19632
rect 759 19598 793 19632
rect 827 19598 861 19632
rect 895 19598 929 19632
rect 963 19598 997 19632
rect 1031 19598 1065 19632
rect 1099 19598 1133 19632
rect 1167 19598 1201 19632
rect 1235 19598 1269 19632
rect 1303 19598 1421 19632
rect 2352 20146 2470 20180
rect 2504 20146 2538 20180
rect 2572 20146 2606 20180
rect 2640 20146 2674 20180
rect 2708 20146 2742 20180
rect 2776 20146 2810 20180
rect 2844 20146 2878 20180
rect 2912 20146 2946 20180
rect 2980 20146 3014 20180
rect 3048 20146 3082 20180
rect 3116 20146 3150 20180
rect 3184 20146 3218 20180
rect 3252 20146 3286 20180
rect 3320 20146 3354 20180
rect 3388 20146 3422 20180
rect 3456 20146 3574 20180
rect 2352 20078 2386 20146
rect 3540 20078 3574 20146
rect 2450 20044 2466 20078
rect 2500 20044 2516 20078
rect 2642 20044 2658 20078
rect 2692 20044 2708 20078
rect 2834 20044 2850 20078
rect 2884 20044 2900 20078
rect 3026 20044 3042 20078
rect 3076 20044 3092 20078
rect 3218 20044 3234 20078
rect 3268 20044 3284 20078
rect 3410 20044 3426 20078
rect 3460 20044 3476 20078
rect 2352 20010 2386 20044
rect 3540 20010 3574 20018
rect 2352 19942 2386 19976
rect 2352 19874 2386 19908
rect 2352 19806 2386 19840
rect 2352 19738 2386 19772
rect 2466 19979 2500 20000
rect 2466 19911 2500 19915
rect 2466 19805 2500 19809
rect 2466 19720 2500 19741
rect 2562 19979 2596 20000
rect 2562 19911 2596 19915
rect 2562 19805 2596 19809
rect 2562 19720 2596 19741
rect 2658 19979 2692 20000
rect 2658 19911 2692 19915
rect 2658 19805 2692 19809
rect 2658 19720 2692 19741
rect 2754 19979 2788 20000
rect 2754 19911 2788 19915
rect 2754 19805 2788 19809
rect 2754 19720 2788 19741
rect 2850 19979 2884 20000
rect 2850 19911 2884 19915
rect 2850 19805 2884 19809
rect 2850 19720 2884 19741
rect 2946 19979 2980 20000
rect 2946 19911 2980 19915
rect 2946 19805 2980 19809
rect 2946 19720 2980 19741
rect 3042 19979 3076 20000
rect 3042 19911 3076 19915
rect 3042 19805 3076 19809
rect 3042 19720 3076 19741
rect 3138 19979 3172 20000
rect 3138 19911 3172 19915
rect 3138 19805 3172 19809
rect 3138 19720 3172 19741
rect 3234 19979 3268 20000
rect 3234 19911 3268 19915
rect 3234 19805 3268 19809
rect 3234 19720 3268 19741
rect 3330 19979 3364 20000
rect 3330 19911 3364 19915
rect 3330 19805 3364 19809
rect 3330 19720 3364 19741
rect 3426 19979 3460 20000
rect 3426 19911 3460 19915
rect 3426 19805 3460 19809
rect 3426 19720 3460 19741
rect 3540 19942 3574 19946
rect 3540 19836 3574 19840
rect 3540 19764 3574 19772
rect 2352 19636 2386 19704
rect 3540 19636 3574 19704
rect 2352 19602 2470 19636
rect 2504 19602 2538 19636
rect 2572 19602 2606 19636
rect 2640 19602 2674 19636
rect 2708 19602 2742 19636
rect 2776 19602 2810 19636
rect 2844 19602 2878 19636
rect 2912 19602 2946 19636
rect 2980 19602 3014 19636
rect 3048 19602 3082 19636
rect 3116 19602 3150 19636
rect 3184 19602 3218 19636
rect 3252 19602 3286 19636
rect 3320 19602 3354 19636
rect 3388 19602 3422 19636
rect 3456 19602 3574 19636
rect 3873 20146 3991 20180
rect 4025 20146 4059 20180
rect 4093 20146 4127 20180
rect 4161 20146 4195 20180
rect 4229 20146 4263 20180
rect 4297 20146 4331 20180
rect 4365 20146 4399 20180
rect 4433 20146 4467 20180
rect 4501 20146 4535 20180
rect 4569 20146 4603 20180
rect 4637 20146 4671 20180
rect 4705 20146 4739 20180
rect 4773 20146 4807 20180
rect 4841 20146 4875 20180
rect 4909 20146 4943 20180
rect 4977 20146 5095 20180
rect 3873 20078 3907 20146
rect 5061 20078 5095 20146
rect 3971 20044 3987 20078
rect 4021 20044 4037 20078
rect 4163 20044 4179 20078
rect 4213 20044 4229 20078
rect 4355 20044 4371 20078
rect 4405 20044 4421 20078
rect 4547 20044 4563 20078
rect 4597 20044 4613 20078
rect 4739 20044 4755 20078
rect 4789 20044 4805 20078
rect 4931 20044 4947 20078
rect 4981 20044 4997 20078
rect 3873 20010 3907 20044
rect 5061 20010 5095 20018
rect 3873 19942 3907 19976
rect 3873 19874 3907 19908
rect 3873 19806 3907 19840
rect 3873 19738 3907 19772
rect 3987 19979 4021 20000
rect 3987 19911 4021 19915
rect 3987 19805 4021 19809
rect 3987 19720 4021 19741
rect 4083 19979 4117 20000
rect 4083 19911 4117 19915
rect 4083 19805 4117 19809
rect 4083 19720 4117 19741
rect 4179 19979 4213 20000
rect 4179 19911 4213 19915
rect 4179 19805 4213 19809
rect 4179 19720 4213 19741
rect 4275 19979 4309 20000
rect 4275 19911 4309 19915
rect 4275 19805 4309 19809
rect 4275 19720 4309 19741
rect 4371 19979 4405 20000
rect 4371 19911 4405 19915
rect 4371 19805 4405 19809
rect 4371 19720 4405 19741
rect 4467 19979 4501 20000
rect 4467 19911 4501 19915
rect 4467 19805 4501 19809
rect 4467 19720 4501 19741
rect 4563 19979 4597 20000
rect 4563 19911 4597 19915
rect 4563 19805 4597 19809
rect 4563 19720 4597 19741
rect 4659 19979 4693 20000
rect 4659 19911 4693 19915
rect 4659 19805 4693 19809
rect 4659 19720 4693 19741
rect 4755 19979 4789 20000
rect 4755 19911 4789 19915
rect 4755 19805 4789 19809
rect 4755 19720 4789 19741
rect 4851 19979 4885 20000
rect 4851 19911 4885 19915
rect 4851 19805 4885 19809
rect 4851 19720 4885 19741
rect 4947 19979 4981 20000
rect 4947 19911 4981 19915
rect 4947 19805 4981 19809
rect 4947 19720 4981 19741
rect 5061 19942 5095 19946
rect 5061 19836 5095 19840
rect 5274 19813 5303 19847
rect 5337 19813 5395 19847
rect 5429 19813 5487 19847
rect 5521 19813 5550 19847
rect 5061 19764 5095 19772
rect 3873 19636 3907 19704
rect 5061 19636 5095 19704
rect 3873 19602 3991 19636
rect 4025 19602 4059 19636
rect 4093 19602 4127 19636
rect 4161 19602 4195 19636
rect 4229 19602 4263 19636
rect 4297 19602 4331 19636
rect 4365 19602 4399 19636
rect 4433 19602 4467 19636
rect 4501 19602 4535 19636
rect 4569 19602 4603 19636
rect 4637 19602 4671 19636
rect 4705 19602 4739 19636
rect 4773 19602 4807 19636
rect 4841 19602 4875 19636
rect 4909 19602 4943 19636
rect 4977 19602 5095 19636
rect 5340 19771 5406 19779
rect 5340 19737 5356 19771
rect 5390 19737 5406 19771
rect 5340 19703 5406 19737
rect 5340 19669 5356 19703
rect 5390 19669 5406 19703
rect 5340 19635 5406 19669
rect 5340 19601 5356 19635
rect 5390 19601 5406 19635
rect 5340 19583 5406 19601
rect 5440 19771 5482 19813
rect 5474 19737 5482 19771
rect 5440 19703 5482 19737
rect 5474 19669 5482 19703
rect 5440 19635 5482 19669
rect 5474 19601 5482 19635
rect 5440 19585 5482 19601
rect 5340 19533 5386 19583
rect 199 19490 317 19524
rect 351 19490 385 19524
rect 419 19490 453 19524
rect 487 19490 521 19524
rect 555 19490 589 19524
rect 623 19490 657 19524
rect 691 19490 725 19524
rect 759 19490 793 19524
rect 827 19490 861 19524
rect 895 19490 929 19524
rect 963 19490 997 19524
rect 1031 19490 1065 19524
rect 1099 19490 1133 19524
rect 1167 19490 1201 19524
rect 1235 19490 1269 19524
rect 1303 19490 1421 19524
rect 199 19414 233 19490
rect 1387 19419 1421 19490
rect 199 19346 233 19380
rect 199 19278 233 19312
rect 313 19377 347 19416
rect 313 19304 347 19343
rect 409 19377 443 19416
rect 409 19304 443 19343
rect 505 19377 539 19416
rect 505 19304 539 19343
rect 601 19377 635 19416
rect 601 19304 635 19343
rect 697 19377 731 19416
rect 697 19304 731 19343
rect 793 19377 827 19416
rect 793 19304 827 19343
rect 889 19377 923 19416
rect 889 19304 923 19343
rect 985 19377 1019 19416
rect 985 19304 1019 19343
rect 1081 19377 1115 19416
rect 1081 19304 1115 19343
rect 1177 19377 1211 19416
rect 1177 19304 1211 19343
rect 1273 19377 1307 19416
rect 1273 19304 1307 19343
rect 1387 19347 1421 19380
rect 1387 19278 1421 19312
rect 199 19168 233 19244
rect 297 19232 313 19266
rect 347 19232 363 19266
rect 489 19232 505 19266
rect 539 19232 555 19266
rect 681 19232 697 19266
rect 731 19232 747 19266
rect 873 19232 889 19266
rect 923 19232 939 19266
rect 1065 19232 1081 19266
rect 1115 19232 1131 19266
rect 1257 19232 1273 19266
rect 1307 19232 1323 19266
rect 1387 19168 1421 19241
rect 199 19134 317 19168
rect 351 19134 385 19168
rect 419 19134 453 19168
rect 487 19134 521 19168
rect 555 19134 589 19168
rect 623 19134 657 19168
rect 691 19134 725 19168
rect 759 19134 793 19168
rect 827 19134 861 19168
rect 895 19134 929 19168
rect 963 19134 997 19168
rect 1031 19134 1065 19168
rect 1099 19134 1133 19168
rect 1167 19134 1201 19168
rect 1235 19134 1269 19168
rect 1303 19134 1421 19168
rect 2352 19494 2470 19528
rect 2504 19494 2538 19528
rect 2572 19494 2606 19528
rect 2640 19494 2674 19528
rect 2708 19494 2742 19528
rect 2776 19494 2810 19528
rect 2844 19494 2878 19528
rect 2912 19494 2946 19528
rect 2980 19494 3014 19528
rect 3048 19494 3082 19528
rect 3116 19494 3150 19528
rect 3184 19494 3218 19528
rect 3252 19494 3286 19528
rect 3320 19494 3354 19528
rect 3388 19494 3422 19528
rect 3456 19494 3574 19528
rect 2352 19418 2386 19494
rect 3540 19423 3574 19494
rect 3873 19494 3991 19528
rect 4025 19494 4059 19528
rect 4093 19494 4127 19528
rect 4161 19494 4195 19528
rect 4229 19494 4263 19528
rect 4297 19494 4331 19528
rect 4365 19494 4399 19528
rect 4433 19494 4467 19528
rect 4501 19494 4535 19528
rect 4569 19494 4603 19528
rect 4637 19494 4671 19528
rect 4705 19494 4739 19528
rect 4773 19494 4807 19528
rect 4841 19494 4875 19528
rect 4909 19494 4943 19528
rect 4977 19494 5095 19528
rect 3675 19458 3691 19492
rect 3725 19458 3741 19492
rect 2352 19350 2386 19384
rect 2352 19282 2386 19316
rect 2466 19381 2500 19420
rect 2466 19308 2500 19347
rect 2562 19381 2596 19420
rect 2562 19308 2596 19347
rect 2658 19381 2692 19420
rect 2658 19308 2692 19347
rect 2754 19381 2788 19420
rect 2754 19308 2788 19347
rect 2850 19381 2884 19420
rect 2850 19308 2884 19347
rect 2946 19381 2980 19420
rect 2946 19308 2980 19347
rect 3042 19381 3076 19420
rect 3042 19308 3076 19347
rect 3138 19381 3172 19420
rect 3138 19308 3172 19347
rect 3234 19381 3268 19420
rect 3234 19308 3268 19347
rect 3330 19381 3364 19420
rect 3330 19308 3364 19347
rect 3426 19381 3460 19420
rect 3426 19308 3460 19347
rect 3540 19351 3574 19384
rect 3647 19408 3681 19424
rect 3647 19316 3681 19332
rect 3735 19408 3769 19424
rect 3735 19316 3769 19332
rect 3873 19418 3907 19494
rect 5061 19423 5095 19494
rect 3873 19350 3907 19384
rect 3540 19282 3574 19316
rect 2352 19172 2386 19248
rect 2450 19236 2466 19270
rect 2500 19236 2516 19270
rect 2642 19236 2658 19270
rect 2692 19236 2708 19270
rect 2834 19236 2850 19270
rect 2884 19236 2900 19270
rect 3026 19236 3042 19270
rect 3076 19236 3092 19270
rect 3218 19236 3234 19270
rect 3268 19236 3284 19270
rect 3410 19236 3426 19270
rect 3460 19236 3476 19270
rect 3540 19172 3574 19245
rect 2352 19138 2470 19172
rect 2504 19138 2538 19172
rect 2572 19138 2606 19172
rect 2640 19138 2674 19172
rect 2708 19138 2742 19172
rect 2776 19138 2810 19172
rect 2844 19138 2878 19172
rect 2912 19138 2946 19172
rect 2980 19138 3014 19172
rect 3048 19138 3082 19172
rect 3116 19138 3150 19172
rect 3184 19138 3218 19172
rect 3252 19138 3286 19172
rect 3320 19138 3354 19172
rect 3388 19138 3422 19172
rect 3456 19138 3574 19172
rect 3873 19282 3907 19316
rect 3987 19381 4021 19420
rect 3987 19308 4021 19347
rect 4083 19381 4117 19420
rect 4083 19308 4117 19347
rect 4179 19381 4213 19420
rect 4179 19308 4213 19347
rect 4275 19381 4309 19420
rect 4275 19308 4309 19347
rect 4371 19381 4405 19420
rect 4371 19308 4405 19347
rect 4467 19381 4501 19420
rect 4467 19308 4501 19347
rect 4563 19381 4597 19420
rect 4563 19308 4597 19347
rect 4659 19381 4693 19420
rect 4659 19308 4693 19347
rect 4755 19381 4789 19420
rect 4755 19308 4789 19347
rect 4851 19381 4885 19420
rect 4851 19308 4885 19347
rect 4947 19381 4981 19420
rect 4947 19308 4981 19347
rect 5061 19351 5095 19384
rect 5340 19499 5348 19533
rect 5382 19499 5386 19533
rect 5420 19538 5486 19549
rect 5420 19535 5450 19538
rect 5420 19501 5436 19535
rect 5484 19504 5486 19538
rect 5470 19501 5486 19504
rect 5340 19463 5386 19499
rect 5340 19451 5406 19463
rect 5340 19417 5356 19451
rect 5390 19417 5406 19451
rect 5340 19383 5406 19417
rect 5340 19349 5356 19383
rect 5390 19349 5406 19383
rect 5340 19337 5406 19349
rect 5440 19451 5486 19467
rect 5474 19417 5486 19451
rect 5440 19383 5486 19417
rect 5474 19349 5486 19383
rect 5061 19282 5095 19316
rect 5440 19303 5486 19349
rect 3873 19172 3907 19248
rect 3971 19236 3987 19270
rect 4021 19236 4037 19270
rect 4163 19236 4179 19270
rect 4213 19236 4229 19270
rect 4355 19236 4371 19270
rect 4405 19236 4421 19270
rect 4547 19236 4563 19270
rect 4597 19236 4613 19270
rect 4739 19236 4755 19270
rect 4789 19236 4805 19270
rect 4931 19236 4947 19270
rect 4981 19236 4997 19270
rect 5274 19269 5303 19303
rect 5337 19269 5395 19303
rect 5429 19269 5487 19303
rect 5521 19269 5550 19303
rect 5061 19172 5095 19245
rect 3873 19138 3991 19172
rect 4025 19138 4059 19172
rect 4093 19138 4127 19172
rect 4161 19138 4195 19172
rect 4229 19138 4263 19172
rect 4297 19138 4331 19172
rect 4365 19138 4399 19172
rect 4433 19138 4467 19172
rect 4501 19138 4535 19172
rect 4569 19138 4603 19172
rect 4637 19138 4671 19172
rect 4705 19138 4739 19172
rect 4773 19138 4807 19172
rect 4841 19138 4875 19172
rect 4909 19138 4943 19172
rect 4977 19138 5095 19172
rect 199 18855 317 18889
rect 351 18855 385 18889
rect 419 18855 453 18889
rect 487 18855 521 18889
rect 555 18855 589 18889
rect 623 18855 657 18889
rect 691 18855 725 18889
rect 759 18855 793 18889
rect 827 18855 861 18889
rect 895 18855 929 18889
rect 963 18855 997 18889
rect 1031 18855 1065 18889
rect 1099 18855 1133 18889
rect 1167 18855 1201 18889
rect 1235 18855 1269 18889
rect 1303 18855 1421 18889
rect 199 18787 233 18855
rect 1387 18787 1421 18855
rect 297 18753 313 18787
rect 347 18753 363 18787
rect 489 18753 505 18787
rect 539 18753 555 18787
rect 681 18753 697 18787
rect 731 18753 747 18787
rect 873 18753 889 18787
rect 923 18753 939 18787
rect 1065 18753 1081 18787
rect 1115 18753 1131 18787
rect 1257 18753 1273 18787
rect 1307 18753 1323 18787
rect 199 18719 233 18753
rect 1387 18719 1421 18727
rect 199 18651 233 18685
rect 199 18583 233 18617
rect 199 18515 233 18549
rect 199 18447 233 18481
rect 313 18688 347 18709
rect 313 18620 347 18624
rect 313 18514 347 18518
rect 313 18429 347 18450
rect 409 18688 443 18709
rect 409 18620 443 18624
rect 409 18514 443 18518
rect 409 18429 443 18450
rect 505 18688 539 18709
rect 505 18620 539 18624
rect 505 18514 539 18518
rect 505 18429 539 18450
rect 601 18688 635 18709
rect 601 18620 635 18624
rect 601 18514 635 18518
rect 601 18429 635 18450
rect 697 18688 731 18709
rect 697 18620 731 18624
rect 697 18514 731 18518
rect 697 18429 731 18450
rect 793 18688 827 18709
rect 793 18620 827 18624
rect 793 18514 827 18518
rect 793 18429 827 18450
rect 889 18688 923 18709
rect 889 18620 923 18624
rect 889 18514 923 18518
rect 889 18429 923 18450
rect 985 18688 1019 18709
rect 985 18620 1019 18624
rect 985 18514 1019 18518
rect 985 18429 1019 18450
rect 1081 18688 1115 18709
rect 1081 18620 1115 18624
rect 1081 18514 1115 18518
rect 1081 18429 1115 18450
rect 1177 18688 1211 18709
rect 1177 18620 1211 18624
rect 1177 18514 1211 18518
rect 1177 18429 1211 18450
rect 1273 18688 1307 18709
rect 1273 18620 1307 18624
rect 1273 18514 1307 18518
rect 1273 18429 1307 18450
rect 1387 18651 1421 18655
rect 1387 18545 1421 18549
rect 1387 18473 1421 18481
rect 199 18345 233 18413
rect 1387 18345 1421 18413
rect 199 18311 317 18345
rect 351 18311 385 18345
rect 419 18311 453 18345
rect 487 18311 521 18345
rect 555 18311 589 18345
rect 623 18311 657 18345
rect 691 18311 725 18345
rect 759 18311 793 18345
rect 827 18311 861 18345
rect 895 18311 929 18345
rect 963 18311 997 18345
rect 1031 18311 1065 18345
rect 1099 18311 1133 18345
rect 1167 18311 1201 18345
rect 1235 18311 1269 18345
rect 1303 18311 1421 18345
rect 2352 18859 2470 18893
rect 2504 18859 2538 18893
rect 2572 18859 2606 18893
rect 2640 18859 2674 18893
rect 2708 18859 2742 18893
rect 2776 18859 2810 18893
rect 2844 18859 2878 18893
rect 2912 18859 2946 18893
rect 2980 18859 3014 18893
rect 3048 18859 3082 18893
rect 3116 18859 3150 18893
rect 3184 18859 3218 18893
rect 3252 18859 3286 18893
rect 3320 18859 3354 18893
rect 3388 18859 3422 18893
rect 3456 18859 3574 18893
rect 2352 18791 2386 18859
rect 3540 18791 3574 18859
rect 2450 18757 2466 18791
rect 2500 18757 2516 18791
rect 2642 18757 2658 18791
rect 2692 18757 2708 18791
rect 2834 18757 2850 18791
rect 2884 18757 2900 18791
rect 3026 18757 3042 18791
rect 3076 18757 3092 18791
rect 3218 18757 3234 18791
rect 3268 18757 3284 18791
rect 3410 18757 3426 18791
rect 3460 18757 3476 18791
rect 2352 18723 2386 18757
rect 3540 18723 3574 18731
rect 2352 18655 2386 18689
rect 2352 18587 2386 18621
rect 2352 18519 2386 18553
rect 2352 18451 2386 18485
rect 2466 18692 2500 18713
rect 2466 18624 2500 18628
rect 2466 18518 2500 18522
rect 2466 18433 2500 18454
rect 2562 18692 2596 18713
rect 2562 18624 2596 18628
rect 2562 18518 2596 18522
rect 2562 18433 2596 18454
rect 2658 18692 2692 18713
rect 2658 18624 2692 18628
rect 2658 18518 2692 18522
rect 2658 18433 2692 18454
rect 2754 18692 2788 18713
rect 2754 18624 2788 18628
rect 2754 18518 2788 18522
rect 2754 18433 2788 18454
rect 2850 18692 2884 18713
rect 2850 18624 2884 18628
rect 2850 18518 2884 18522
rect 2850 18433 2884 18454
rect 2946 18692 2980 18713
rect 2946 18624 2980 18628
rect 2946 18518 2980 18522
rect 2946 18433 2980 18454
rect 3042 18692 3076 18713
rect 3042 18624 3076 18628
rect 3042 18518 3076 18522
rect 3042 18433 3076 18454
rect 3138 18692 3172 18713
rect 3138 18624 3172 18628
rect 3138 18518 3172 18522
rect 3138 18433 3172 18454
rect 3234 18692 3268 18713
rect 3234 18624 3268 18628
rect 3234 18518 3268 18522
rect 3234 18433 3268 18454
rect 3330 18692 3364 18713
rect 3330 18624 3364 18628
rect 3330 18518 3364 18522
rect 3330 18433 3364 18454
rect 3426 18692 3460 18713
rect 3426 18624 3460 18628
rect 3426 18518 3460 18522
rect 3426 18433 3460 18454
rect 3540 18655 3574 18659
rect 3540 18549 3574 18553
rect 3540 18477 3574 18485
rect 2352 18349 2386 18417
rect 3540 18349 3574 18417
rect 2352 18315 2470 18349
rect 2504 18315 2538 18349
rect 2572 18315 2606 18349
rect 2640 18315 2674 18349
rect 2708 18315 2742 18349
rect 2776 18315 2810 18349
rect 2844 18315 2878 18349
rect 2912 18315 2946 18349
rect 2980 18315 3014 18349
rect 3048 18315 3082 18349
rect 3116 18315 3150 18349
rect 3184 18315 3218 18349
rect 3252 18315 3286 18349
rect 3320 18315 3354 18349
rect 3388 18315 3422 18349
rect 3456 18315 3574 18349
rect 3873 18859 3991 18893
rect 4025 18859 4059 18893
rect 4093 18859 4127 18893
rect 4161 18859 4195 18893
rect 4229 18859 4263 18893
rect 4297 18859 4331 18893
rect 4365 18859 4399 18893
rect 4433 18859 4467 18893
rect 4501 18859 4535 18893
rect 4569 18859 4603 18893
rect 4637 18859 4671 18893
rect 4705 18859 4739 18893
rect 4773 18859 4807 18893
rect 4841 18859 4875 18893
rect 4909 18859 4943 18893
rect 4977 18859 5095 18893
rect 3873 18791 3907 18859
rect 5061 18791 5095 18859
rect 3971 18757 3987 18791
rect 4021 18757 4037 18791
rect 4163 18757 4179 18791
rect 4213 18757 4229 18791
rect 4355 18757 4371 18791
rect 4405 18757 4421 18791
rect 4547 18757 4563 18791
rect 4597 18757 4613 18791
rect 4739 18757 4755 18791
rect 4789 18757 4805 18791
rect 4931 18757 4947 18791
rect 4981 18757 4997 18791
rect 3873 18723 3907 18757
rect 5061 18723 5095 18731
rect 3873 18655 3907 18689
rect 3873 18587 3907 18621
rect 3873 18519 3907 18553
rect 3873 18451 3907 18485
rect 3987 18692 4021 18713
rect 3987 18624 4021 18628
rect 3987 18518 4021 18522
rect 3987 18433 4021 18454
rect 4083 18692 4117 18713
rect 4083 18624 4117 18628
rect 4083 18518 4117 18522
rect 4083 18433 4117 18454
rect 4179 18692 4213 18713
rect 4179 18624 4213 18628
rect 4179 18518 4213 18522
rect 4179 18433 4213 18454
rect 4275 18692 4309 18713
rect 4275 18624 4309 18628
rect 4275 18518 4309 18522
rect 4275 18433 4309 18454
rect 4371 18692 4405 18713
rect 4371 18624 4405 18628
rect 4371 18518 4405 18522
rect 4371 18433 4405 18454
rect 4467 18692 4501 18713
rect 4467 18624 4501 18628
rect 4467 18518 4501 18522
rect 4467 18433 4501 18454
rect 4563 18692 4597 18713
rect 4563 18624 4597 18628
rect 4563 18518 4597 18522
rect 4563 18433 4597 18454
rect 4659 18692 4693 18713
rect 4659 18624 4693 18628
rect 4659 18518 4693 18522
rect 4659 18433 4693 18454
rect 4755 18692 4789 18713
rect 4755 18624 4789 18628
rect 4755 18518 4789 18522
rect 4755 18433 4789 18454
rect 4851 18692 4885 18713
rect 4851 18624 4885 18628
rect 4851 18518 4885 18522
rect 4851 18433 4885 18454
rect 4947 18692 4981 18713
rect 4947 18624 4981 18628
rect 4947 18518 4981 18522
rect 4947 18433 4981 18454
rect 5061 18655 5095 18659
rect 5061 18549 5095 18553
rect 5274 18526 5303 18560
rect 5337 18526 5395 18560
rect 5429 18526 5487 18560
rect 5521 18526 5550 18560
rect 5061 18477 5095 18485
rect 3873 18349 3907 18417
rect 5061 18349 5095 18417
rect 3873 18315 3991 18349
rect 4025 18315 4059 18349
rect 4093 18315 4127 18349
rect 4161 18315 4195 18349
rect 4229 18315 4263 18349
rect 4297 18315 4331 18349
rect 4365 18315 4399 18349
rect 4433 18315 4467 18349
rect 4501 18315 4535 18349
rect 4569 18315 4603 18349
rect 4637 18315 4671 18349
rect 4705 18315 4739 18349
rect 4773 18315 4807 18349
rect 4841 18315 4875 18349
rect 4909 18315 4943 18349
rect 4977 18315 5095 18349
rect 5340 18484 5406 18492
rect 5340 18450 5356 18484
rect 5390 18450 5406 18484
rect 5340 18416 5406 18450
rect 5340 18382 5356 18416
rect 5390 18382 5406 18416
rect 5340 18348 5406 18382
rect 5340 18314 5356 18348
rect 5390 18314 5406 18348
rect 5340 18296 5406 18314
rect 5440 18484 5482 18526
rect 5474 18450 5482 18484
rect 5440 18416 5482 18450
rect 5474 18382 5482 18416
rect 5440 18348 5482 18382
rect 5474 18314 5482 18348
rect 5440 18298 5482 18314
rect 5340 18246 5386 18296
rect 199 18203 317 18237
rect 351 18203 385 18237
rect 419 18203 453 18237
rect 487 18203 521 18237
rect 555 18203 589 18237
rect 623 18203 657 18237
rect 691 18203 725 18237
rect 759 18203 793 18237
rect 827 18203 861 18237
rect 895 18203 929 18237
rect 963 18203 997 18237
rect 1031 18203 1065 18237
rect 1099 18203 1133 18237
rect 1167 18203 1201 18237
rect 1235 18203 1269 18237
rect 1303 18203 1421 18237
rect 199 18127 233 18203
rect 1387 18132 1421 18203
rect 199 18059 233 18093
rect 199 17991 233 18025
rect 313 18090 347 18129
rect 313 18017 347 18056
rect 409 18090 443 18129
rect 409 18017 443 18056
rect 505 18090 539 18129
rect 505 18017 539 18056
rect 601 18090 635 18129
rect 601 18017 635 18056
rect 697 18090 731 18129
rect 697 18017 731 18056
rect 793 18090 827 18129
rect 793 18017 827 18056
rect 889 18090 923 18129
rect 889 18017 923 18056
rect 985 18090 1019 18129
rect 985 18017 1019 18056
rect 1081 18090 1115 18129
rect 1081 18017 1115 18056
rect 1177 18090 1211 18129
rect 1177 18017 1211 18056
rect 1273 18090 1307 18129
rect 1273 18017 1307 18056
rect 1387 18060 1421 18093
rect 1387 17991 1421 18025
rect 199 17881 233 17957
rect 297 17945 313 17979
rect 347 17945 363 17979
rect 489 17945 505 17979
rect 539 17945 555 17979
rect 681 17945 697 17979
rect 731 17945 747 17979
rect 873 17945 889 17979
rect 923 17945 939 17979
rect 1065 17945 1081 17979
rect 1115 17945 1131 17979
rect 1257 17945 1273 17979
rect 1307 17945 1323 17979
rect 1387 17881 1421 17954
rect 199 17847 317 17881
rect 351 17847 385 17881
rect 419 17847 453 17881
rect 487 17847 521 17881
rect 555 17847 589 17881
rect 623 17847 657 17881
rect 691 17847 725 17881
rect 759 17847 793 17881
rect 827 17847 861 17881
rect 895 17847 929 17881
rect 963 17847 997 17881
rect 1031 17847 1065 17881
rect 1099 17847 1133 17881
rect 1167 17847 1201 17881
rect 1235 17847 1269 17881
rect 1303 17847 1421 17881
rect 2352 18207 2470 18241
rect 2504 18207 2538 18241
rect 2572 18207 2606 18241
rect 2640 18207 2674 18241
rect 2708 18207 2742 18241
rect 2776 18207 2810 18241
rect 2844 18207 2878 18241
rect 2912 18207 2946 18241
rect 2980 18207 3014 18241
rect 3048 18207 3082 18241
rect 3116 18207 3150 18241
rect 3184 18207 3218 18241
rect 3252 18207 3286 18241
rect 3320 18207 3354 18241
rect 3388 18207 3422 18241
rect 3456 18207 3574 18241
rect 2352 18131 2386 18207
rect 3540 18136 3574 18207
rect 3873 18207 3991 18241
rect 4025 18207 4059 18241
rect 4093 18207 4127 18241
rect 4161 18207 4195 18241
rect 4229 18207 4263 18241
rect 4297 18207 4331 18241
rect 4365 18207 4399 18241
rect 4433 18207 4467 18241
rect 4501 18207 4535 18241
rect 4569 18207 4603 18241
rect 4637 18207 4671 18241
rect 4705 18207 4739 18241
rect 4773 18207 4807 18241
rect 4841 18207 4875 18241
rect 4909 18207 4943 18241
rect 4977 18207 5095 18241
rect 3675 18171 3691 18205
rect 3725 18171 3741 18205
rect 2352 18063 2386 18097
rect 2352 17995 2386 18029
rect 2466 18094 2500 18133
rect 2466 18021 2500 18060
rect 2562 18094 2596 18133
rect 2562 18021 2596 18060
rect 2658 18094 2692 18133
rect 2658 18021 2692 18060
rect 2754 18094 2788 18133
rect 2754 18021 2788 18060
rect 2850 18094 2884 18133
rect 2850 18021 2884 18060
rect 2946 18094 2980 18133
rect 2946 18021 2980 18060
rect 3042 18094 3076 18133
rect 3042 18021 3076 18060
rect 3138 18094 3172 18133
rect 3138 18021 3172 18060
rect 3234 18094 3268 18133
rect 3234 18021 3268 18060
rect 3330 18094 3364 18133
rect 3330 18021 3364 18060
rect 3426 18094 3460 18133
rect 3426 18021 3460 18060
rect 3540 18064 3574 18097
rect 3647 18121 3681 18137
rect 3647 18029 3681 18045
rect 3735 18121 3769 18137
rect 3735 18029 3769 18045
rect 3873 18131 3907 18207
rect 5061 18136 5095 18207
rect 3873 18063 3907 18097
rect 3540 17995 3574 18029
rect 2352 17885 2386 17961
rect 2450 17949 2466 17983
rect 2500 17949 2516 17983
rect 2642 17949 2658 17983
rect 2692 17949 2708 17983
rect 2834 17949 2850 17983
rect 2884 17949 2900 17983
rect 3026 17949 3042 17983
rect 3076 17949 3092 17983
rect 3218 17949 3234 17983
rect 3268 17949 3284 17983
rect 3410 17949 3426 17983
rect 3460 17949 3476 17983
rect 3540 17885 3574 17958
rect 2352 17851 2470 17885
rect 2504 17851 2538 17885
rect 2572 17851 2606 17885
rect 2640 17851 2674 17885
rect 2708 17851 2742 17885
rect 2776 17851 2810 17885
rect 2844 17851 2878 17885
rect 2912 17851 2946 17885
rect 2980 17851 3014 17885
rect 3048 17851 3082 17885
rect 3116 17851 3150 17885
rect 3184 17851 3218 17885
rect 3252 17851 3286 17885
rect 3320 17851 3354 17885
rect 3388 17851 3422 17885
rect 3456 17851 3574 17885
rect 3873 17995 3907 18029
rect 3987 18094 4021 18133
rect 3987 18021 4021 18060
rect 4083 18094 4117 18133
rect 4083 18021 4117 18060
rect 4179 18094 4213 18133
rect 4179 18021 4213 18060
rect 4275 18094 4309 18133
rect 4275 18021 4309 18060
rect 4371 18094 4405 18133
rect 4371 18021 4405 18060
rect 4467 18094 4501 18133
rect 4467 18021 4501 18060
rect 4563 18094 4597 18133
rect 4563 18021 4597 18060
rect 4659 18094 4693 18133
rect 4659 18021 4693 18060
rect 4755 18094 4789 18133
rect 4755 18021 4789 18060
rect 4851 18094 4885 18133
rect 4851 18021 4885 18060
rect 4947 18094 4981 18133
rect 4947 18021 4981 18060
rect 5061 18064 5095 18097
rect 5340 18212 5348 18246
rect 5382 18212 5386 18246
rect 5420 18251 5486 18262
rect 5420 18248 5450 18251
rect 5420 18214 5436 18248
rect 5484 18217 5486 18251
rect 5470 18214 5486 18217
rect 5340 18176 5386 18212
rect 5340 18164 5406 18176
rect 5340 18130 5356 18164
rect 5390 18130 5406 18164
rect 5340 18096 5406 18130
rect 5340 18062 5356 18096
rect 5390 18062 5406 18096
rect 5340 18050 5406 18062
rect 5440 18164 5486 18180
rect 5474 18130 5486 18164
rect 5440 18096 5486 18130
rect 5474 18062 5486 18096
rect 5061 17995 5095 18029
rect 5440 18016 5486 18062
rect 3873 17885 3907 17961
rect 3971 17949 3987 17983
rect 4021 17949 4037 17983
rect 4163 17949 4179 17983
rect 4213 17949 4229 17983
rect 4355 17949 4371 17983
rect 4405 17949 4421 17983
rect 4547 17949 4563 17983
rect 4597 17949 4613 17983
rect 4739 17949 4755 17983
rect 4789 17949 4805 17983
rect 4931 17949 4947 17983
rect 4981 17949 4997 17983
rect 5274 17982 5303 18016
rect 5337 17982 5395 18016
rect 5429 17982 5487 18016
rect 5521 17982 5550 18016
rect 5061 17885 5095 17958
rect 3873 17851 3991 17885
rect 4025 17851 4059 17885
rect 4093 17851 4127 17885
rect 4161 17851 4195 17885
rect 4229 17851 4263 17885
rect 4297 17851 4331 17885
rect 4365 17851 4399 17885
rect 4433 17851 4467 17885
rect 4501 17851 4535 17885
rect 4569 17851 4603 17885
rect 4637 17851 4671 17885
rect 4705 17851 4739 17885
rect 4773 17851 4807 17885
rect 4841 17851 4875 17885
rect 4909 17851 4943 17885
rect 4977 17851 5095 17885
rect 199 17568 317 17602
rect 351 17568 385 17602
rect 419 17568 453 17602
rect 487 17568 521 17602
rect 555 17568 589 17602
rect 623 17568 657 17602
rect 691 17568 725 17602
rect 759 17568 793 17602
rect 827 17568 861 17602
rect 895 17568 929 17602
rect 963 17568 997 17602
rect 1031 17568 1065 17602
rect 1099 17568 1133 17602
rect 1167 17568 1201 17602
rect 1235 17568 1269 17602
rect 1303 17568 1421 17602
rect 199 17500 233 17568
rect 1387 17500 1421 17568
rect 297 17466 313 17500
rect 347 17466 363 17500
rect 489 17466 505 17500
rect 539 17466 555 17500
rect 681 17466 697 17500
rect 731 17466 747 17500
rect 873 17466 889 17500
rect 923 17466 939 17500
rect 1065 17466 1081 17500
rect 1115 17466 1131 17500
rect 1257 17466 1273 17500
rect 1307 17466 1323 17500
rect 199 17432 233 17466
rect 1387 17432 1421 17440
rect 199 17364 233 17398
rect 199 17296 233 17330
rect 199 17228 233 17262
rect 199 17160 233 17194
rect 313 17401 347 17422
rect 313 17333 347 17337
rect 313 17227 347 17231
rect 313 17142 347 17163
rect 409 17401 443 17422
rect 409 17333 443 17337
rect 409 17227 443 17231
rect 409 17142 443 17163
rect 505 17401 539 17422
rect 505 17333 539 17337
rect 505 17227 539 17231
rect 505 17142 539 17163
rect 601 17401 635 17422
rect 601 17333 635 17337
rect 601 17227 635 17231
rect 601 17142 635 17163
rect 697 17401 731 17422
rect 697 17333 731 17337
rect 697 17227 731 17231
rect 697 17142 731 17163
rect 793 17401 827 17422
rect 793 17333 827 17337
rect 793 17227 827 17231
rect 793 17142 827 17163
rect 889 17401 923 17422
rect 889 17333 923 17337
rect 889 17227 923 17231
rect 889 17142 923 17163
rect 985 17401 1019 17422
rect 985 17333 1019 17337
rect 985 17227 1019 17231
rect 985 17142 1019 17163
rect 1081 17401 1115 17422
rect 1081 17333 1115 17337
rect 1081 17227 1115 17231
rect 1081 17142 1115 17163
rect 1177 17401 1211 17422
rect 1177 17333 1211 17337
rect 1177 17227 1211 17231
rect 1177 17142 1211 17163
rect 1273 17401 1307 17422
rect 1273 17333 1307 17337
rect 1273 17227 1307 17231
rect 1273 17142 1307 17163
rect 1387 17364 1421 17368
rect 1387 17258 1421 17262
rect 1387 17186 1421 17194
rect 199 17058 233 17126
rect 1387 17058 1421 17126
rect 199 17024 317 17058
rect 351 17024 385 17058
rect 419 17024 453 17058
rect 487 17024 521 17058
rect 555 17024 589 17058
rect 623 17024 657 17058
rect 691 17024 725 17058
rect 759 17024 793 17058
rect 827 17024 861 17058
rect 895 17024 929 17058
rect 963 17024 997 17058
rect 1031 17024 1065 17058
rect 1099 17024 1133 17058
rect 1167 17024 1201 17058
rect 1235 17024 1269 17058
rect 1303 17024 1421 17058
rect 2352 17572 2470 17606
rect 2504 17572 2538 17606
rect 2572 17572 2606 17606
rect 2640 17572 2674 17606
rect 2708 17572 2742 17606
rect 2776 17572 2810 17606
rect 2844 17572 2878 17606
rect 2912 17572 2946 17606
rect 2980 17572 3014 17606
rect 3048 17572 3082 17606
rect 3116 17572 3150 17606
rect 3184 17572 3218 17606
rect 3252 17572 3286 17606
rect 3320 17572 3354 17606
rect 3388 17572 3422 17606
rect 3456 17572 3574 17606
rect 2352 17504 2386 17572
rect 3540 17504 3574 17572
rect 2450 17470 2466 17504
rect 2500 17470 2516 17504
rect 2642 17470 2658 17504
rect 2692 17470 2708 17504
rect 2834 17470 2850 17504
rect 2884 17470 2900 17504
rect 3026 17470 3042 17504
rect 3076 17470 3092 17504
rect 3218 17470 3234 17504
rect 3268 17470 3284 17504
rect 3410 17470 3426 17504
rect 3460 17470 3476 17504
rect 2352 17436 2386 17470
rect 3540 17436 3574 17444
rect 2352 17368 2386 17402
rect 2352 17300 2386 17334
rect 2352 17232 2386 17266
rect 2352 17164 2386 17198
rect 2466 17405 2500 17426
rect 2466 17337 2500 17341
rect 2466 17231 2500 17235
rect 2466 17146 2500 17167
rect 2562 17405 2596 17426
rect 2562 17337 2596 17341
rect 2562 17231 2596 17235
rect 2562 17146 2596 17167
rect 2658 17405 2692 17426
rect 2658 17337 2692 17341
rect 2658 17231 2692 17235
rect 2658 17146 2692 17167
rect 2754 17405 2788 17426
rect 2754 17337 2788 17341
rect 2754 17231 2788 17235
rect 2754 17146 2788 17167
rect 2850 17405 2884 17426
rect 2850 17337 2884 17341
rect 2850 17231 2884 17235
rect 2850 17146 2884 17167
rect 2946 17405 2980 17426
rect 2946 17337 2980 17341
rect 2946 17231 2980 17235
rect 2946 17146 2980 17167
rect 3042 17405 3076 17426
rect 3042 17337 3076 17341
rect 3042 17231 3076 17235
rect 3042 17146 3076 17167
rect 3138 17405 3172 17426
rect 3138 17337 3172 17341
rect 3138 17231 3172 17235
rect 3138 17146 3172 17167
rect 3234 17405 3268 17426
rect 3234 17337 3268 17341
rect 3234 17231 3268 17235
rect 3234 17146 3268 17167
rect 3330 17405 3364 17426
rect 3330 17337 3364 17341
rect 3330 17231 3364 17235
rect 3330 17146 3364 17167
rect 3426 17405 3460 17426
rect 3426 17337 3460 17341
rect 3426 17231 3460 17235
rect 3426 17146 3460 17167
rect 3540 17368 3574 17372
rect 3540 17262 3574 17266
rect 3540 17190 3574 17198
rect 2352 17062 2386 17130
rect 3540 17062 3574 17130
rect 2352 17028 2470 17062
rect 2504 17028 2538 17062
rect 2572 17028 2606 17062
rect 2640 17028 2674 17062
rect 2708 17028 2742 17062
rect 2776 17028 2810 17062
rect 2844 17028 2878 17062
rect 2912 17028 2946 17062
rect 2980 17028 3014 17062
rect 3048 17028 3082 17062
rect 3116 17028 3150 17062
rect 3184 17028 3218 17062
rect 3252 17028 3286 17062
rect 3320 17028 3354 17062
rect 3388 17028 3422 17062
rect 3456 17028 3574 17062
rect 3873 17572 3991 17606
rect 4025 17572 4059 17606
rect 4093 17572 4127 17606
rect 4161 17572 4195 17606
rect 4229 17572 4263 17606
rect 4297 17572 4331 17606
rect 4365 17572 4399 17606
rect 4433 17572 4467 17606
rect 4501 17572 4535 17606
rect 4569 17572 4603 17606
rect 4637 17572 4671 17606
rect 4705 17572 4739 17606
rect 4773 17572 4807 17606
rect 4841 17572 4875 17606
rect 4909 17572 4943 17606
rect 4977 17572 5095 17606
rect 3873 17504 3907 17572
rect 5061 17504 5095 17572
rect 3971 17470 3987 17504
rect 4021 17470 4037 17504
rect 4163 17470 4179 17504
rect 4213 17470 4229 17504
rect 4355 17470 4371 17504
rect 4405 17470 4421 17504
rect 4547 17470 4563 17504
rect 4597 17470 4613 17504
rect 4739 17470 4755 17504
rect 4789 17470 4805 17504
rect 4931 17470 4947 17504
rect 4981 17470 4997 17504
rect 3873 17436 3907 17470
rect 5061 17436 5095 17444
rect 3873 17368 3907 17402
rect 3873 17300 3907 17334
rect 3873 17232 3907 17266
rect 3873 17164 3907 17198
rect 3987 17405 4021 17426
rect 3987 17337 4021 17341
rect 3987 17231 4021 17235
rect 3987 17146 4021 17167
rect 4083 17405 4117 17426
rect 4083 17337 4117 17341
rect 4083 17231 4117 17235
rect 4083 17146 4117 17167
rect 4179 17405 4213 17426
rect 4179 17337 4213 17341
rect 4179 17231 4213 17235
rect 4179 17146 4213 17167
rect 4275 17405 4309 17426
rect 4275 17337 4309 17341
rect 4275 17231 4309 17235
rect 4275 17146 4309 17167
rect 4371 17405 4405 17426
rect 4371 17337 4405 17341
rect 4371 17231 4405 17235
rect 4371 17146 4405 17167
rect 4467 17405 4501 17426
rect 4467 17337 4501 17341
rect 4467 17231 4501 17235
rect 4467 17146 4501 17167
rect 4563 17405 4597 17426
rect 4563 17337 4597 17341
rect 4563 17231 4597 17235
rect 4563 17146 4597 17167
rect 4659 17405 4693 17426
rect 4659 17337 4693 17341
rect 4659 17231 4693 17235
rect 4659 17146 4693 17167
rect 4755 17405 4789 17426
rect 4755 17337 4789 17341
rect 4755 17231 4789 17235
rect 4755 17146 4789 17167
rect 4851 17405 4885 17426
rect 4851 17337 4885 17341
rect 4851 17231 4885 17235
rect 4851 17146 4885 17167
rect 4947 17405 4981 17426
rect 4947 17337 4981 17341
rect 4947 17231 4981 17235
rect 4947 17146 4981 17167
rect 5061 17368 5095 17372
rect 5061 17262 5095 17266
rect 5274 17239 5303 17273
rect 5337 17239 5395 17273
rect 5429 17239 5487 17273
rect 5521 17239 5550 17273
rect 5061 17190 5095 17198
rect 3873 17062 3907 17130
rect 5061 17062 5095 17130
rect 3873 17028 3991 17062
rect 4025 17028 4059 17062
rect 4093 17028 4127 17062
rect 4161 17028 4195 17062
rect 4229 17028 4263 17062
rect 4297 17028 4331 17062
rect 4365 17028 4399 17062
rect 4433 17028 4467 17062
rect 4501 17028 4535 17062
rect 4569 17028 4603 17062
rect 4637 17028 4671 17062
rect 4705 17028 4739 17062
rect 4773 17028 4807 17062
rect 4841 17028 4875 17062
rect 4909 17028 4943 17062
rect 4977 17028 5095 17062
rect 5340 17197 5406 17205
rect 5340 17163 5356 17197
rect 5390 17163 5406 17197
rect 5340 17129 5406 17163
rect 5340 17095 5356 17129
rect 5390 17095 5406 17129
rect 5340 17061 5406 17095
rect 5340 17027 5356 17061
rect 5390 17027 5406 17061
rect 5340 17009 5406 17027
rect 5440 17197 5482 17239
rect 5474 17163 5482 17197
rect 5440 17129 5482 17163
rect 5474 17095 5482 17129
rect 5440 17061 5482 17095
rect 5474 17027 5482 17061
rect 5440 17011 5482 17027
rect 5340 16959 5386 17009
rect 199 16916 317 16950
rect 351 16916 385 16950
rect 419 16916 453 16950
rect 487 16916 521 16950
rect 555 16916 589 16950
rect 623 16916 657 16950
rect 691 16916 725 16950
rect 759 16916 793 16950
rect 827 16916 861 16950
rect 895 16916 929 16950
rect 963 16916 997 16950
rect 1031 16916 1065 16950
rect 1099 16916 1133 16950
rect 1167 16916 1201 16950
rect 1235 16916 1269 16950
rect 1303 16916 1421 16950
rect 199 16840 233 16916
rect 1387 16845 1421 16916
rect 199 16772 233 16806
rect 199 16704 233 16738
rect 313 16803 347 16842
rect 313 16730 347 16769
rect 409 16803 443 16842
rect 409 16730 443 16769
rect 505 16803 539 16842
rect 505 16730 539 16769
rect 601 16803 635 16842
rect 601 16730 635 16769
rect 697 16803 731 16842
rect 697 16730 731 16769
rect 793 16803 827 16842
rect 793 16730 827 16769
rect 889 16803 923 16842
rect 889 16730 923 16769
rect 985 16803 1019 16842
rect 985 16730 1019 16769
rect 1081 16803 1115 16842
rect 1081 16730 1115 16769
rect 1177 16803 1211 16842
rect 1177 16730 1211 16769
rect 1273 16803 1307 16842
rect 1273 16730 1307 16769
rect 1387 16773 1421 16806
rect 1387 16704 1421 16738
rect 199 16594 233 16670
rect 297 16658 313 16692
rect 347 16658 363 16692
rect 489 16658 505 16692
rect 539 16658 555 16692
rect 681 16658 697 16692
rect 731 16658 747 16692
rect 873 16658 889 16692
rect 923 16658 939 16692
rect 1065 16658 1081 16692
rect 1115 16658 1131 16692
rect 1257 16658 1273 16692
rect 1307 16658 1323 16692
rect 1387 16594 1421 16667
rect 199 16560 317 16594
rect 351 16560 385 16594
rect 419 16560 453 16594
rect 487 16560 521 16594
rect 555 16560 589 16594
rect 623 16560 657 16594
rect 691 16560 725 16594
rect 759 16560 793 16594
rect 827 16560 861 16594
rect 895 16560 929 16594
rect 963 16560 997 16594
rect 1031 16560 1065 16594
rect 1099 16560 1133 16594
rect 1167 16560 1201 16594
rect 1235 16560 1269 16594
rect 1303 16560 1421 16594
rect 2352 16920 2470 16954
rect 2504 16920 2538 16954
rect 2572 16920 2606 16954
rect 2640 16920 2674 16954
rect 2708 16920 2742 16954
rect 2776 16920 2810 16954
rect 2844 16920 2878 16954
rect 2912 16920 2946 16954
rect 2980 16920 3014 16954
rect 3048 16920 3082 16954
rect 3116 16920 3150 16954
rect 3184 16920 3218 16954
rect 3252 16920 3286 16954
rect 3320 16920 3354 16954
rect 3388 16920 3422 16954
rect 3456 16920 3574 16954
rect 2352 16844 2386 16920
rect 3540 16849 3574 16920
rect 3873 16920 3991 16954
rect 4025 16920 4059 16954
rect 4093 16920 4127 16954
rect 4161 16920 4195 16954
rect 4229 16920 4263 16954
rect 4297 16920 4331 16954
rect 4365 16920 4399 16954
rect 4433 16920 4467 16954
rect 4501 16920 4535 16954
rect 4569 16920 4603 16954
rect 4637 16920 4671 16954
rect 4705 16920 4739 16954
rect 4773 16920 4807 16954
rect 4841 16920 4875 16954
rect 4909 16920 4943 16954
rect 4977 16920 5095 16954
rect 3675 16884 3691 16918
rect 3725 16884 3741 16918
rect 2352 16776 2386 16810
rect 2352 16708 2386 16742
rect 2466 16807 2500 16846
rect 2466 16734 2500 16773
rect 2562 16807 2596 16846
rect 2562 16734 2596 16773
rect 2658 16807 2692 16846
rect 2658 16734 2692 16773
rect 2754 16807 2788 16846
rect 2754 16734 2788 16773
rect 2850 16807 2884 16846
rect 2850 16734 2884 16773
rect 2946 16807 2980 16846
rect 2946 16734 2980 16773
rect 3042 16807 3076 16846
rect 3042 16734 3076 16773
rect 3138 16807 3172 16846
rect 3138 16734 3172 16773
rect 3234 16807 3268 16846
rect 3234 16734 3268 16773
rect 3330 16807 3364 16846
rect 3330 16734 3364 16773
rect 3426 16807 3460 16846
rect 3426 16734 3460 16773
rect 3540 16777 3574 16810
rect 3647 16834 3681 16850
rect 3647 16742 3681 16758
rect 3735 16834 3769 16850
rect 3735 16742 3769 16758
rect 3873 16844 3907 16920
rect 5061 16849 5095 16920
rect 3873 16776 3907 16810
rect 3540 16708 3574 16742
rect 2352 16598 2386 16674
rect 2450 16662 2466 16696
rect 2500 16662 2516 16696
rect 2642 16662 2658 16696
rect 2692 16662 2708 16696
rect 2834 16662 2850 16696
rect 2884 16662 2900 16696
rect 3026 16662 3042 16696
rect 3076 16662 3092 16696
rect 3218 16662 3234 16696
rect 3268 16662 3284 16696
rect 3410 16662 3426 16696
rect 3460 16662 3476 16696
rect 3540 16598 3574 16671
rect 2352 16564 2470 16598
rect 2504 16564 2538 16598
rect 2572 16564 2606 16598
rect 2640 16564 2674 16598
rect 2708 16564 2742 16598
rect 2776 16564 2810 16598
rect 2844 16564 2878 16598
rect 2912 16564 2946 16598
rect 2980 16564 3014 16598
rect 3048 16564 3082 16598
rect 3116 16564 3150 16598
rect 3184 16564 3218 16598
rect 3252 16564 3286 16598
rect 3320 16564 3354 16598
rect 3388 16564 3422 16598
rect 3456 16564 3574 16598
rect 3873 16708 3907 16742
rect 3987 16807 4021 16846
rect 3987 16734 4021 16773
rect 4083 16807 4117 16846
rect 4083 16734 4117 16773
rect 4179 16807 4213 16846
rect 4179 16734 4213 16773
rect 4275 16807 4309 16846
rect 4275 16734 4309 16773
rect 4371 16807 4405 16846
rect 4371 16734 4405 16773
rect 4467 16807 4501 16846
rect 4467 16734 4501 16773
rect 4563 16807 4597 16846
rect 4563 16734 4597 16773
rect 4659 16807 4693 16846
rect 4659 16734 4693 16773
rect 4755 16807 4789 16846
rect 4755 16734 4789 16773
rect 4851 16807 4885 16846
rect 4851 16734 4885 16773
rect 4947 16807 4981 16846
rect 4947 16734 4981 16773
rect 5061 16777 5095 16810
rect 5340 16925 5348 16959
rect 5382 16925 5386 16959
rect 5420 16964 5486 16975
rect 5420 16961 5450 16964
rect 5420 16927 5436 16961
rect 5484 16930 5486 16964
rect 5470 16927 5486 16930
rect 5340 16889 5386 16925
rect 5340 16877 5406 16889
rect 5340 16843 5356 16877
rect 5390 16843 5406 16877
rect 5340 16809 5406 16843
rect 5340 16775 5356 16809
rect 5390 16775 5406 16809
rect 5340 16763 5406 16775
rect 5440 16877 5486 16893
rect 5474 16843 5486 16877
rect 5440 16809 5486 16843
rect 5474 16775 5486 16809
rect 5061 16708 5095 16742
rect 5440 16729 5486 16775
rect 3873 16598 3907 16674
rect 3971 16662 3987 16696
rect 4021 16662 4037 16696
rect 4163 16662 4179 16696
rect 4213 16662 4229 16696
rect 4355 16662 4371 16696
rect 4405 16662 4421 16696
rect 4547 16662 4563 16696
rect 4597 16662 4613 16696
rect 4739 16662 4755 16696
rect 4789 16662 4805 16696
rect 4931 16662 4947 16696
rect 4981 16662 4997 16696
rect 5274 16695 5303 16729
rect 5337 16695 5395 16729
rect 5429 16695 5487 16729
rect 5521 16695 5550 16729
rect 5061 16598 5095 16671
rect 3873 16564 3991 16598
rect 4025 16564 4059 16598
rect 4093 16564 4127 16598
rect 4161 16564 4195 16598
rect 4229 16564 4263 16598
rect 4297 16564 4331 16598
rect 4365 16564 4399 16598
rect 4433 16564 4467 16598
rect 4501 16564 4535 16598
rect 4569 16564 4603 16598
rect 4637 16564 4671 16598
rect 4705 16564 4739 16598
rect 4773 16564 4807 16598
rect 4841 16564 4875 16598
rect 4909 16564 4943 16598
rect 4977 16564 5095 16598
rect 199 16281 317 16315
rect 351 16281 385 16315
rect 419 16281 453 16315
rect 487 16281 521 16315
rect 555 16281 589 16315
rect 623 16281 657 16315
rect 691 16281 725 16315
rect 759 16281 793 16315
rect 827 16281 861 16315
rect 895 16281 929 16315
rect 963 16281 997 16315
rect 1031 16281 1065 16315
rect 1099 16281 1133 16315
rect 1167 16281 1201 16315
rect 1235 16281 1269 16315
rect 1303 16281 1421 16315
rect 199 16213 233 16281
rect 1387 16213 1421 16281
rect 297 16179 313 16213
rect 347 16179 363 16213
rect 489 16179 505 16213
rect 539 16179 555 16213
rect 681 16179 697 16213
rect 731 16179 747 16213
rect 873 16179 889 16213
rect 923 16179 939 16213
rect 1065 16179 1081 16213
rect 1115 16179 1131 16213
rect 1257 16179 1273 16213
rect 1307 16179 1323 16213
rect 199 16145 233 16179
rect 1387 16145 1421 16153
rect 199 16077 233 16111
rect 199 16009 233 16043
rect 199 15941 233 15975
rect 199 15873 233 15907
rect 313 16114 347 16135
rect 313 16046 347 16050
rect 313 15940 347 15944
rect 313 15855 347 15876
rect 409 16114 443 16135
rect 409 16046 443 16050
rect 409 15940 443 15944
rect 409 15855 443 15876
rect 505 16114 539 16135
rect 505 16046 539 16050
rect 505 15940 539 15944
rect 505 15855 539 15876
rect 601 16114 635 16135
rect 601 16046 635 16050
rect 601 15940 635 15944
rect 601 15855 635 15876
rect 697 16114 731 16135
rect 697 16046 731 16050
rect 697 15940 731 15944
rect 697 15855 731 15876
rect 793 16114 827 16135
rect 793 16046 827 16050
rect 793 15940 827 15944
rect 793 15855 827 15876
rect 889 16114 923 16135
rect 889 16046 923 16050
rect 889 15940 923 15944
rect 889 15855 923 15876
rect 985 16114 1019 16135
rect 985 16046 1019 16050
rect 985 15940 1019 15944
rect 985 15855 1019 15876
rect 1081 16114 1115 16135
rect 1081 16046 1115 16050
rect 1081 15940 1115 15944
rect 1081 15855 1115 15876
rect 1177 16114 1211 16135
rect 1177 16046 1211 16050
rect 1177 15940 1211 15944
rect 1177 15855 1211 15876
rect 1273 16114 1307 16135
rect 1273 16046 1307 16050
rect 1273 15940 1307 15944
rect 1273 15855 1307 15876
rect 1387 16077 1421 16081
rect 1387 15971 1421 15975
rect 1387 15899 1421 15907
rect 199 15771 233 15839
rect 1387 15771 1421 15839
rect 199 15737 317 15771
rect 351 15737 385 15771
rect 419 15737 453 15771
rect 487 15737 521 15771
rect 555 15737 589 15771
rect 623 15737 657 15771
rect 691 15737 725 15771
rect 759 15737 793 15771
rect 827 15737 861 15771
rect 895 15737 929 15771
rect 963 15737 997 15771
rect 1031 15737 1065 15771
rect 1099 15737 1133 15771
rect 1167 15737 1201 15771
rect 1235 15737 1269 15771
rect 1303 15737 1421 15771
rect 2352 16285 2470 16319
rect 2504 16285 2538 16319
rect 2572 16285 2606 16319
rect 2640 16285 2674 16319
rect 2708 16285 2742 16319
rect 2776 16285 2810 16319
rect 2844 16285 2878 16319
rect 2912 16285 2946 16319
rect 2980 16285 3014 16319
rect 3048 16285 3082 16319
rect 3116 16285 3150 16319
rect 3184 16285 3218 16319
rect 3252 16285 3286 16319
rect 3320 16285 3354 16319
rect 3388 16285 3422 16319
rect 3456 16285 3574 16319
rect 2352 16217 2386 16285
rect 3540 16217 3574 16285
rect 2450 16183 2466 16217
rect 2500 16183 2516 16217
rect 2642 16183 2658 16217
rect 2692 16183 2708 16217
rect 2834 16183 2850 16217
rect 2884 16183 2900 16217
rect 3026 16183 3042 16217
rect 3076 16183 3092 16217
rect 3218 16183 3234 16217
rect 3268 16183 3284 16217
rect 3410 16183 3426 16217
rect 3460 16183 3476 16217
rect 2352 16149 2386 16183
rect 3540 16149 3574 16157
rect 2352 16081 2386 16115
rect 2352 16013 2386 16047
rect 2352 15945 2386 15979
rect 2352 15877 2386 15911
rect 2466 16118 2500 16139
rect 2466 16050 2500 16054
rect 2466 15944 2500 15948
rect 2466 15859 2500 15880
rect 2562 16118 2596 16139
rect 2562 16050 2596 16054
rect 2562 15944 2596 15948
rect 2562 15859 2596 15880
rect 2658 16118 2692 16139
rect 2658 16050 2692 16054
rect 2658 15944 2692 15948
rect 2658 15859 2692 15880
rect 2754 16118 2788 16139
rect 2754 16050 2788 16054
rect 2754 15944 2788 15948
rect 2754 15859 2788 15880
rect 2850 16118 2884 16139
rect 2850 16050 2884 16054
rect 2850 15944 2884 15948
rect 2850 15859 2884 15880
rect 2946 16118 2980 16139
rect 2946 16050 2980 16054
rect 2946 15944 2980 15948
rect 2946 15859 2980 15880
rect 3042 16118 3076 16139
rect 3042 16050 3076 16054
rect 3042 15944 3076 15948
rect 3042 15859 3076 15880
rect 3138 16118 3172 16139
rect 3138 16050 3172 16054
rect 3138 15944 3172 15948
rect 3138 15859 3172 15880
rect 3234 16118 3268 16139
rect 3234 16050 3268 16054
rect 3234 15944 3268 15948
rect 3234 15859 3268 15880
rect 3330 16118 3364 16139
rect 3330 16050 3364 16054
rect 3330 15944 3364 15948
rect 3330 15859 3364 15880
rect 3426 16118 3460 16139
rect 3426 16050 3460 16054
rect 3426 15944 3460 15948
rect 3426 15859 3460 15880
rect 3540 16081 3574 16085
rect 3540 15975 3574 15979
rect 3540 15903 3574 15911
rect 2352 15775 2386 15843
rect 3540 15775 3574 15843
rect 2352 15741 2470 15775
rect 2504 15741 2538 15775
rect 2572 15741 2606 15775
rect 2640 15741 2674 15775
rect 2708 15741 2742 15775
rect 2776 15741 2810 15775
rect 2844 15741 2878 15775
rect 2912 15741 2946 15775
rect 2980 15741 3014 15775
rect 3048 15741 3082 15775
rect 3116 15741 3150 15775
rect 3184 15741 3218 15775
rect 3252 15741 3286 15775
rect 3320 15741 3354 15775
rect 3388 15741 3422 15775
rect 3456 15741 3574 15775
rect 3873 16285 3991 16319
rect 4025 16285 4059 16319
rect 4093 16285 4127 16319
rect 4161 16285 4195 16319
rect 4229 16285 4263 16319
rect 4297 16285 4331 16319
rect 4365 16285 4399 16319
rect 4433 16285 4467 16319
rect 4501 16285 4535 16319
rect 4569 16285 4603 16319
rect 4637 16285 4671 16319
rect 4705 16285 4739 16319
rect 4773 16285 4807 16319
rect 4841 16285 4875 16319
rect 4909 16285 4943 16319
rect 4977 16285 5095 16319
rect 3873 16217 3907 16285
rect 5061 16217 5095 16285
rect 3971 16183 3987 16217
rect 4021 16183 4037 16217
rect 4163 16183 4179 16217
rect 4213 16183 4229 16217
rect 4355 16183 4371 16217
rect 4405 16183 4421 16217
rect 4547 16183 4563 16217
rect 4597 16183 4613 16217
rect 4739 16183 4755 16217
rect 4789 16183 4805 16217
rect 4931 16183 4947 16217
rect 4981 16183 4997 16217
rect 3873 16149 3907 16183
rect 5061 16149 5095 16157
rect 3873 16081 3907 16115
rect 3873 16013 3907 16047
rect 3873 15945 3907 15979
rect 3873 15877 3907 15911
rect 3987 16118 4021 16139
rect 3987 16050 4021 16054
rect 3987 15944 4021 15948
rect 3987 15859 4021 15880
rect 4083 16118 4117 16139
rect 4083 16050 4117 16054
rect 4083 15944 4117 15948
rect 4083 15859 4117 15880
rect 4179 16118 4213 16139
rect 4179 16050 4213 16054
rect 4179 15944 4213 15948
rect 4179 15859 4213 15880
rect 4275 16118 4309 16139
rect 4275 16050 4309 16054
rect 4275 15944 4309 15948
rect 4275 15859 4309 15880
rect 4371 16118 4405 16139
rect 4371 16050 4405 16054
rect 4371 15944 4405 15948
rect 4371 15859 4405 15880
rect 4467 16118 4501 16139
rect 4467 16050 4501 16054
rect 4467 15944 4501 15948
rect 4467 15859 4501 15880
rect 4563 16118 4597 16139
rect 4563 16050 4597 16054
rect 4563 15944 4597 15948
rect 4563 15859 4597 15880
rect 4659 16118 4693 16139
rect 4659 16050 4693 16054
rect 4659 15944 4693 15948
rect 4659 15859 4693 15880
rect 4755 16118 4789 16139
rect 4755 16050 4789 16054
rect 4755 15944 4789 15948
rect 4755 15859 4789 15880
rect 4851 16118 4885 16139
rect 4851 16050 4885 16054
rect 4851 15944 4885 15948
rect 4851 15859 4885 15880
rect 4947 16118 4981 16139
rect 4947 16050 4981 16054
rect 4947 15944 4981 15948
rect 4947 15859 4981 15880
rect 5061 16081 5095 16085
rect 5061 15975 5095 15979
rect 5274 15952 5303 15986
rect 5337 15952 5395 15986
rect 5429 15952 5487 15986
rect 5521 15952 5550 15986
rect 5061 15903 5095 15911
rect 3873 15775 3907 15843
rect 5061 15775 5095 15843
rect 3873 15741 3991 15775
rect 4025 15741 4059 15775
rect 4093 15741 4127 15775
rect 4161 15741 4195 15775
rect 4229 15741 4263 15775
rect 4297 15741 4331 15775
rect 4365 15741 4399 15775
rect 4433 15741 4467 15775
rect 4501 15741 4535 15775
rect 4569 15741 4603 15775
rect 4637 15741 4671 15775
rect 4705 15741 4739 15775
rect 4773 15741 4807 15775
rect 4841 15741 4875 15775
rect 4909 15741 4943 15775
rect 4977 15741 5095 15775
rect 5340 15910 5406 15918
rect 5340 15876 5356 15910
rect 5390 15876 5406 15910
rect 5340 15842 5406 15876
rect 5340 15808 5356 15842
rect 5390 15808 5406 15842
rect 5340 15774 5406 15808
rect 5340 15740 5356 15774
rect 5390 15740 5406 15774
rect 5340 15722 5406 15740
rect 5440 15910 5482 15952
rect 5474 15876 5482 15910
rect 5440 15842 5482 15876
rect 5474 15808 5482 15842
rect 5440 15774 5482 15808
rect 5474 15740 5482 15774
rect 5440 15724 5482 15740
rect 5340 15672 5386 15722
rect 199 15629 317 15663
rect 351 15629 385 15663
rect 419 15629 453 15663
rect 487 15629 521 15663
rect 555 15629 589 15663
rect 623 15629 657 15663
rect 691 15629 725 15663
rect 759 15629 793 15663
rect 827 15629 861 15663
rect 895 15629 929 15663
rect 963 15629 997 15663
rect 1031 15629 1065 15663
rect 1099 15629 1133 15663
rect 1167 15629 1201 15663
rect 1235 15629 1269 15663
rect 1303 15629 1421 15663
rect 199 15553 233 15629
rect 1387 15558 1421 15629
rect 199 15485 233 15519
rect 199 15417 233 15451
rect 313 15516 347 15555
rect 313 15443 347 15482
rect 409 15516 443 15555
rect 409 15443 443 15482
rect 505 15516 539 15555
rect 505 15443 539 15482
rect 601 15516 635 15555
rect 601 15443 635 15482
rect 697 15516 731 15555
rect 697 15443 731 15482
rect 793 15516 827 15555
rect 793 15443 827 15482
rect 889 15516 923 15555
rect 889 15443 923 15482
rect 985 15516 1019 15555
rect 985 15443 1019 15482
rect 1081 15516 1115 15555
rect 1081 15443 1115 15482
rect 1177 15516 1211 15555
rect 1177 15443 1211 15482
rect 1273 15516 1307 15555
rect 1273 15443 1307 15482
rect 1387 15486 1421 15519
rect 1387 15417 1421 15451
rect 199 15307 233 15383
rect 297 15371 313 15405
rect 347 15371 363 15405
rect 489 15371 505 15405
rect 539 15371 555 15405
rect 681 15371 697 15405
rect 731 15371 747 15405
rect 873 15371 889 15405
rect 923 15371 939 15405
rect 1065 15371 1081 15405
rect 1115 15371 1131 15405
rect 1257 15371 1273 15405
rect 1307 15371 1323 15405
rect 1387 15307 1421 15380
rect 199 15273 317 15307
rect 351 15273 385 15307
rect 419 15273 453 15307
rect 487 15273 521 15307
rect 555 15273 589 15307
rect 623 15273 657 15307
rect 691 15273 725 15307
rect 759 15273 793 15307
rect 827 15273 861 15307
rect 895 15273 929 15307
rect 963 15273 997 15307
rect 1031 15273 1065 15307
rect 1099 15273 1133 15307
rect 1167 15273 1201 15307
rect 1235 15273 1269 15307
rect 1303 15273 1421 15307
rect 2352 15633 2470 15667
rect 2504 15633 2538 15667
rect 2572 15633 2606 15667
rect 2640 15633 2674 15667
rect 2708 15633 2742 15667
rect 2776 15633 2810 15667
rect 2844 15633 2878 15667
rect 2912 15633 2946 15667
rect 2980 15633 3014 15667
rect 3048 15633 3082 15667
rect 3116 15633 3150 15667
rect 3184 15633 3218 15667
rect 3252 15633 3286 15667
rect 3320 15633 3354 15667
rect 3388 15633 3422 15667
rect 3456 15633 3574 15667
rect 2352 15557 2386 15633
rect 3540 15562 3574 15633
rect 3873 15633 3991 15667
rect 4025 15633 4059 15667
rect 4093 15633 4127 15667
rect 4161 15633 4195 15667
rect 4229 15633 4263 15667
rect 4297 15633 4331 15667
rect 4365 15633 4399 15667
rect 4433 15633 4467 15667
rect 4501 15633 4535 15667
rect 4569 15633 4603 15667
rect 4637 15633 4671 15667
rect 4705 15633 4739 15667
rect 4773 15633 4807 15667
rect 4841 15633 4875 15667
rect 4909 15633 4943 15667
rect 4977 15633 5095 15667
rect 3675 15597 3691 15631
rect 3725 15597 3741 15631
rect 2352 15489 2386 15523
rect 2352 15421 2386 15455
rect 2466 15520 2500 15559
rect 2466 15447 2500 15486
rect 2562 15520 2596 15559
rect 2562 15447 2596 15486
rect 2658 15520 2692 15559
rect 2658 15447 2692 15486
rect 2754 15520 2788 15559
rect 2754 15447 2788 15486
rect 2850 15520 2884 15559
rect 2850 15447 2884 15486
rect 2946 15520 2980 15559
rect 2946 15447 2980 15486
rect 3042 15520 3076 15559
rect 3042 15447 3076 15486
rect 3138 15520 3172 15559
rect 3138 15447 3172 15486
rect 3234 15520 3268 15559
rect 3234 15447 3268 15486
rect 3330 15520 3364 15559
rect 3330 15447 3364 15486
rect 3426 15520 3460 15559
rect 3426 15447 3460 15486
rect 3540 15490 3574 15523
rect 3647 15547 3681 15563
rect 3647 15455 3681 15471
rect 3735 15547 3769 15563
rect 3735 15455 3769 15471
rect 3873 15557 3907 15633
rect 5061 15562 5095 15633
rect 3873 15489 3907 15523
rect 3540 15421 3574 15455
rect 2352 15311 2386 15387
rect 2450 15375 2466 15409
rect 2500 15375 2516 15409
rect 2642 15375 2658 15409
rect 2692 15375 2708 15409
rect 2834 15375 2850 15409
rect 2884 15375 2900 15409
rect 3026 15375 3042 15409
rect 3076 15375 3092 15409
rect 3218 15375 3234 15409
rect 3268 15375 3284 15409
rect 3410 15375 3426 15409
rect 3460 15375 3476 15409
rect 3540 15311 3574 15384
rect 2352 15277 2470 15311
rect 2504 15277 2538 15311
rect 2572 15277 2606 15311
rect 2640 15277 2674 15311
rect 2708 15277 2742 15311
rect 2776 15277 2810 15311
rect 2844 15277 2878 15311
rect 2912 15277 2946 15311
rect 2980 15277 3014 15311
rect 3048 15277 3082 15311
rect 3116 15277 3150 15311
rect 3184 15277 3218 15311
rect 3252 15277 3286 15311
rect 3320 15277 3354 15311
rect 3388 15277 3422 15311
rect 3456 15277 3574 15311
rect 3873 15421 3907 15455
rect 3987 15520 4021 15559
rect 3987 15447 4021 15486
rect 4083 15520 4117 15559
rect 4083 15447 4117 15486
rect 4179 15520 4213 15559
rect 4179 15447 4213 15486
rect 4275 15520 4309 15559
rect 4275 15447 4309 15486
rect 4371 15520 4405 15559
rect 4371 15447 4405 15486
rect 4467 15520 4501 15559
rect 4467 15447 4501 15486
rect 4563 15520 4597 15559
rect 4563 15447 4597 15486
rect 4659 15520 4693 15559
rect 4659 15447 4693 15486
rect 4755 15520 4789 15559
rect 4755 15447 4789 15486
rect 4851 15520 4885 15559
rect 4851 15447 4885 15486
rect 4947 15520 4981 15559
rect 4947 15447 4981 15486
rect 5061 15490 5095 15523
rect 5340 15638 5348 15672
rect 5382 15638 5386 15672
rect 5420 15677 5486 15688
rect 5420 15674 5450 15677
rect 5420 15640 5436 15674
rect 5484 15643 5486 15677
rect 5470 15640 5486 15643
rect 5340 15602 5386 15638
rect 5340 15590 5406 15602
rect 5340 15556 5356 15590
rect 5390 15556 5406 15590
rect 5340 15522 5406 15556
rect 5340 15488 5356 15522
rect 5390 15488 5406 15522
rect 5340 15476 5406 15488
rect 5440 15590 5486 15606
rect 5474 15556 5486 15590
rect 5440 15522 5486 15556
rect 5474 15488 5486 15522
rect 5061 15421 5095 15455
rect 5440 15442 5486 15488
rect 3873 15311 3907 15387
rect 3971 15375 3987 15409
rect 4021 15375 4037 15409
rect 4163 15375 4179 15409
rect 4213 15375 4229 15409
rect 4355 15375 4371 15409
rect 4405 15375 4421 15409
rect 4547 15375 4563 15409
rect 4597 15375 4613 15409
rect 4739 15375 4755 15409
rect 4789 15375 4805 15409
rect 4931 15375 4947 15409
rect 4981 15375 4997 15409
rect 5274 15408 5303 15442
rect 5337 15408 5395 15442
rect 5429 15408 5487 15442
rect 5521 15408 5550 15442
rect 5061 15311 5095 15384
rect 3873 15277 3991 15311
rect 4025 15277 4059 15311
rect 4093 15277 4127 15311
rect 4161 15277 4195 15311
rect 4229 15277 4263 15311
rect 4297 15277 4331 15311
rect 4365 15277 4399 15311
rect 4433 15277 4467 15311
rect 4501 15277 4535 15311
rect 4569 15277 4603 15311
rect 4637 15277 4671 15311
rect 4705 15277 4739 15311
rect 4773 15277 4807 15311
rect 4841 15277 4875 15311
rect 4909 15277 4943 15311
rect 4977 15277 5095 15311
rect 199 14994 317 15028
rect 351 14994 385 15028
rect 419 14994 453 15028
rect 487 14994 521 15028
rect 555 14994 589 15028
rect 623 14994 657 15028
rect 691 14994 725 15028
rect 759 14994 793 15028
rect 827 14994 861 15028
rect 895 14994 929 15028
rect 963 14994 997 15028
rect 1031 14994 1065 15028
rect 1099 14994 1133 15028
rect 1167 14994 1201 15028
rect 1235 14994 1269 15028
rect 1303 14994 1421 15028
rect 199 14926 233 14994
rect 1387 14926 1421 14994
rect 297 14892 313 14926
rect 347 14892 363 14926
rect 489 14892 505 14926
rect 539 14892 555 14926
rect 681 14892 697 14926
rect 731 14892 747 14926
rect 873 14892 889 14926
rect 923 14892 939 14926
rect 1065 14892 1081 14926
rect 1115 14892 1131 14926
rect 1257 14892 1273 14926
rect 1307 14892 1323 14926
rect 199 14858 233 14892
rect 1387 14858 1421 14866
rect 199 14790 233 14824
rect 199 14722 233 14756
rect 199 14654 233 14688
rect 199 14586 233 14620
rect 313 14827 347 14848
rect 313 14759 347 14763
rect 313 14653 347 14657
rect 313 14568 347 14589
rect 409 14827 443 14848
rect 409 14759 443 14763
rect 409 14653 443 14657
rect 409 14568 443 14589
rect 505 14827 539 14848
rect 505 14759 539 14763
rect 505 14653 539 14657
rect 505 14568 539 14589
rect 601 14827 635 14848
rect 601 14759 635 14763
rect 601 14653 635 14657
rect 601 14568 635 14589
rect 697 14827 731 14848
rect 697 14759 731 14763
rect 697 14653 731 14657
rect 697 14568 731 14589
rect 793 14827 827 14848
rect 793 14759 827 14763
rect 793 14653 827 14657
rect 793 14568 827 14589
rect 889 14827 923 14848
rect 889 14759 923 14763
rect 889 14653 923 14657
rect 889 14568 923 14589
rect 985 14827 1019 14848
rect 985 14759 1019 14763
rect 985 14653 1019 14657
rect 985 14568 1019 14589
rect 1081 14827 1115 14848
rect 1081 14759 1115 14763
rect 1081 14653 1115 14657
rect 1081 14568 1115 14589
rect 1177 14827 1211 14848
rect 1177 14759 1211 14763
rect 1177 14653 1211 14657
rect 1177 14568 1211 14589
rect 1273 14827 1307 14848
rect 1273 14759 1307 14763
rect 1273 14653 1307 14657
rect 1273 14568 1307 14589
rect 1387 14790 1421 14794
rect 1387 14684 1421 14688
rect 1387 14612 1421 14620
rect 199 14484 233 14552
rect 1387 14484 1421 14552
rect 199 14450 317 14484
rect 351 14450 385 14484
rect 419 14450 453 14484
rect 487 14450 521 14484
rect 555 14450 589 14484
rect 623 14450 657 14484
rect 691 14450 725 14484
rect 759 14450 793 14484
rect 827 14450 861 14484
rect 895 14450 929 14484
rect 963 14450 997 14484
rect 1031 14450 1065 14484
rect 1099 14450 1133 14484
rect 1167 14450 1201 14484
rect 1235 14450 1269 14484
rect 1303 14450 1421 14484
rect 2352 14998 2470 15032
rect 2504 14998 2538 15032
rect 2572 14998 2606 15032
rect 2640 14998 2674 15032
rect 2708 14998 2742 15032
rect 2776 14998 2810 15032
rect 2844 14998 2878 15032
rect 2912 14998 2946 15032
rect 2980 14998 3014 15032
rect 3048 14998 3082 15032
rect 3116 14998 3150 15032
rect 3184 14998 3218 15032
rect 3252 14998 3286 15032
rect 3320 14998 3354 15032
rect 3388 14998 3422 15032
rect 3456 14998 3574 15032
rect 2352 14930 2386 14998
rect 3540 14930 3574 14998
rect 2450 14896 2466 14930
rect 2500 14896 2516 14930
rect 2642 14896 2658 14930
rect 2692 14896 2708 14930
rect 2834 14896 2850 14930
rect 2884 14896 2900 14930
rect 3026 14896 3042 14930
rect 3076 14896 3092 14930
rect 3218 14896 3234 14930
rect 3268 14896 3284 14930
rect 3410 14896 3426 14930
rect 3460 14896 3476 14930
rect 2352 14862 2386 14896
rect 3540 14862 3574 14870
rect 2352 14794 2386 14828
rect 2352 14726 2386 14760
rect 2352 14658 2386 14692
rect 2352 14590 2386 14624
rect 2466 14831 2500 14852
rect 2466 14763 2500 14767
rect 2466 14657 2500 14661
rect 2466 14572 2500 14593
rect 2562 14831 2596 14852
rect 2562 14763 2596 14767
rect 2562 14657 2596 14661
rect 2562 14572 2596 14593
rect 2658 14831 2692 14852
rect 2658 14763 2692 14767
rect 2658 14657 2692 14661
rect 2658 14572 2692 14593
rect 2754 14831 2788 14852
rect 2754 14763 2788 14767
rect 2754 14657 2788 14661
rect 2754 14572 2788 14593
rect 2850 14831 2884 14852
rect 2850 14763 2884 14767
rect 2850 14657 2884 14661
rect 2850 14572 2884 14593
rect 2946 14831 2980 14852
rect 2946 14763 2980 14767
rect 2946 14657 2980 14661
rect 2946 14572 2980 14593
rect 3042 14831 3076 14852
rect 3042 14763 3076 14767
rect 3042 14657 3076 14661
rect 3042 14572 3076 14593
rect 3138 14831 3172 14852
rect 3138 14763 3172 14767
rect 3138 14657 3172 14661
rect 3138 14572 3172 14593
rect 3234 14831 3268 14852
rect 3234 14763 3268 14767
rect 3234 14657 3268 14661
rect 3234 14572 3268 14593
rect 3330 14831 3364 14852
rect 3330 14763 3364 14767
rect 3330 14657 3364 14661
rect 3330 14572 3364 14593
rect 3426 14831 3460 14852
rect 3426 14763 3460 14767
rect 3426 14657 3460 14661
rect 3426 14572 3460 14593
rect 3540 14794 3574 14798
rect 3540 14688 3574 14692
rect 3540 14616 3574 14624
rect 2352 14488 2386 14556
rect 3540 14488 3574 14556
rect 2352 14454 2470 14488
rect 2504 14454 2538 14488
rect 2572 14454 2606 14488
rect 2640 14454 2674 14488
rect 2708 14454 2742 14488
rect 2776 14454 2810 14488
rect 2844 14454 2878 14488
rect 2912 14454 2946 14488
rect 2980 14454 3014 14488
rect 3048 14454 3082 14488
rect 3116 14454 3150 14488
rect 3184 14454 3218 14488
rect 3252 14454 3286 14488
rect 3320 14454 3354 14488
rect 3388 14454 3422 14488
rect 3456 14454 3574 14488
rect 3873 14998 3991 15032
rect 4025 14998 4059 15032
rect 4093 14998 4127 15032
rect 4161 14998 4195 15032
rect 4229 14998 4263 15032
rect 4297 14998 4331 15032
rect 4365 14998 4399 15032
rect 4433 14998 4467 15032
rect 4501 14998 4535 15032
rect 4569 14998 4603 15032
rect 4637 14998 4671 15032
rect 4705 14998 4739 15032
rect 4773 14998 4807 15032
rect 4841 14998 4875 15032
rect 4909 14998 4943 15032
rect 4977 14998 5095 15032
rect 3873 14930 3907 14998
rect 5061 14930 5095 14998
rect 3971 14896 3987 14930
rect 4021 14896 4037 14930
rect 4163 14896 4179 14930
rect 4213 14896 4229 14930
rect 4355 14896 4371 14930
rect 4405 14896 4421 14930
rect 4547 14896 4563 14930
rect 4597 14896 4613 14930
rect 4739 14896 4755 14930
rect 4789 14896 4805 14930
rect 4931 14896 4947 14930
rect 4981 14896 4997 14930
rect 3873 14862 3907 14896
rect 5061 14862 5095 14870
rect 3873 14794 3907 14828
rect 3873 14726 3907 14760
rect 3873 14658 3907 14692
rect 3873 14590 3907 14624
rect 3987 14831 4021 14852
rect 3987 14763 4021 14767
rect 3987 14657 4021 14661
rect 3987 14572 4021 14593
rect 4083 14831 4117 14852
rect 4083 14763 4117 14767
rect 4083 14657 4117 14661
rect 4083 14572 4117 14593
rect 4179 14831 4213 14852
rect 4179 14763 4213 14767
rect 4179 14657 4213 14661
rect 4179 14572 4213 14593
rect 4275 14831 4309 14852
rect 4275 14763 4309 14767
rect 4275 14657 4309 14661
rect 4275 14572 4309 14593
rect 4371 14831 4405 14852
rect 4371 14763 4405 14767
rect 4371 14657 4405 14661
rect 4371 14572 4405 14593
rect 4467 14831 4501 14852
rect 4467 14763 4501 14767
rect 4467 14657 4501 14661
rect 4467 14572 4501 14593
rect 4563 14831 4597 14852
rect 4563 14763 4597 14767
rect 4563 14657 4597 14661
rect 4563 14572 4597 14593
rect 4659 14831 4693 14852
rect 4659 14763 4693 14767
rect 4659 14657 4693 14661
rect 4659 14572 4693 14593
rect 4755 14831 4789 14852
rect 4755 14763 4789 14767
rect 4755 14657 4789 14661
rect 4755 14572 4789 14593
rect 4851 14831 4885 14852
rect 4851 14763 4885 14767
rect 4851 14657 4885 14661
rect 4851 14572 4885 14593
rect 4947 14831 4981 14852
rect 4947 14763 4981 14767
rect 4947 14657 4981 14661
rect 4947 14572 4981 14593
rect 5061 14794 5095 14798
rect 5061 14688 5095 14692
rect 5274 14665 5303 14699
rect 5337 14665 5395 14699
rect 5429 14665 5487 14699
rect 5521 14665 5550 14699
rect 5061 14616 5095 14624
rect 3873 14488 3907 14556
rect 5061 14488 5095 14556
rect 3873 14454 3991 14488
rect 4025 14454 4059 14488
rect 4093 14454 4127 14488
rect 4161 14454 4195 14488
rect 4229 14454 4263 14488
rect 4297 14454 4331 14488
rect 4365 14454 4399 14488
rect 4433 14454 4467 14488
rect 4501 14454 4535 14488
rect 4569 14454 4603 14488
rect 4637 14454 4671 14488
rect 4705 14454 4739 14488
rect 4773 14454 4807 14488
rect 4841 14454 4875 14488
rect 4909 14454 4943 14488
rect 4977 14454 5095 14488
rect 5340 14623 5406 14631
rect 5340 14589 5356 14623
rect 5390 14589 5406 14623
rect 5340 14555 5406 14589
rect 5340 14521 5356 14555
rect 5390 14521 5406 14555
rect 5340 14487 5406 14521
rect 5340 14453 5356 14487
rect 5390 14453 5406 14487
rect 5340 14435 5406 14453
rect 5440 14623 5482 14665
rect 5474 14589 5482 14623
rect 5440 14555 5482 14589
rect 5474 14521 5482 14555
rect 5440 14487 5482 14521
rect 5474 14453 5482 14487
rect 5440 14437 5482 14453
rect 5340 14385 5386 14435
rect 199 14342 317 14376
rect 351 14342 385 14376
rect 419 14342 453 14376
rect 487 14342 521 14376
rect 555 14342 589 14376
rect 623 14342 657 14376
rect 691 14342 725 14376
rect 759 14342 793 14376
rect 827 14342 861 14376
rect 895 14342 929 14376
rect 963 14342 997 14376
rect 1031 14342 1065 14376
rect 1099 14342 1133 14376
rect 1167 14342 1201 14376
rect 1235 14342 1269 14376
rect 1303 14342 1421 14376
rect 199 14266 233 14342
rect 1387 14271 1421 14342
rect 199 14198 233 14232
rect 199 14130 233 14164
rect 313 14229 347 14268
rect 313 14156 347 14195
rect 409 14229 443 14268
rect 409 14156 443 14195
rect 505 14229 539 14268
rect 505 14156 539 14195
rect 601 14229 635 14268
rect 601 14156 635 14195
rect 697 14229 731 14268
rect 697 14156 731 14195
rect 793 14229 827 14268
rect 793 14156 827 14195
rect 889 14229 923 14268
rect 889 14156 923 14195
rect 985 14229 1019 14268
rect 985 14156 1019 14195
rect 1081 14229 1115 14268
rect 1081 14156 1115 14195
rect 1177 14229 1211 14268
rect 1177 14156 1211 14195
rect 1273 14229 1307 14268
rect 1273 14156 1307 14195
rect 1387 14199 1421 14232
rect 1387 14130 1421 14164
rect 199 14020 233 14096
rect 297 14084 313 14118
rect 347 14084 363 14118
rect 489 14084 505 14118
rect 539 14084 555 14118
rect 681 14084 697 14118
rect 731 14084 747 14118
rect 873 14084 889 14118
rect 923 14084 939 14118
rect 1065 14084 1081 14118
rect 1115 14084 1131 14118
rect 1257 14084 1273 14118
rect 1307 14084 1323 14118
rect 1387 14020 1421 14093
rect 199 13986 317 14020
rect 351 13986 385 14020
rect 419 13986 453 14020
rect 487 13986 521 14020
rect 555 13986 589 14020
rect 623 13986 657 14020
rect 691 13986 725 14020
rect 759 13986 793 14020
rect 827 13986 861 14020
rect 895 13986 929 14020
rect 963 13986 997 14020
rect 1031 13986 1065 14020
rect 1099 13986 1133 14020
rect 1167 13986 1201 14020
rect 1235 13986 1269 14020
rect 1303 13986 1421 14020
rect 2352 14346 2470 14380
rect 2504 14346 2538 14380
rect 2572 14346 2606 14380
rect 2640 14346 2674 14380
rect 2708 14346 2742 14380
rect 2776 14346 2810 14380
rect 2844 14346 2878 14380
rect 2912 14346 2946 14380
rect 2980 14346 3014 14380
rect 3048 14346 3082 14380
rect 3116 14346 3150 14380
rect 3184 14346 3218 14380
rect 3252 14346 3286 14380
rect 3320 14346 3354 14380
rect 3388 14346 3422 14380
rect 3456 14346 3574 14380
rect 2352 14270 2386 14346
rect 3540 14275 3574 14346
rect 3873 14346 3991 14380
rect 4025 14346 4059 14380
rect 4093 14346 4127 14380
rect 4161 14346 4195 14380
rect 4229 14346 4263 14380
rect 4297 14346 4331 14380
rect 4365 14346 4399 14380
rect 4433 14346 4467 14380
rect 4501 14346 4535 14380
rect 4569 14346 4603 14380
rect 4637 14346 4671 14380
rect 4705 14346 4739 14380
rect 4773 14346 4807 14380
rect 4841 14346 4875 14380
rect 4909 14346 4943 14380
rect 4977 14346 5095 14380
rect 3675 14310 3691 14344
rect 3725 14310 3741 14344
rect 2352 14202 2386 14236
rect 2352 14134 2386 14168
rect 2466 14233 2500 14272
rect 2466 14160 2500 14199
rect 2562 14233 2596 14272
rect 2562 14160 2596 14199
rect 2658 14233 2692 14272
rect 2658 14160 2692 14199
rect 2754 14233 2788 14272
rect 2754 14160 2788 14199
rect 2850 14233 2884 14272
rect 2850 14160 2884 14199
rect 2946 14233 2980 14272
rect 2946 14160 2980 14199
rect 3042 14233 3076 14272
rect 3042 14160 3076 14199
rect 3138 14233 3172 14272
rect 3138 14160 3172 14199
rect 3234 14233 3268 14272
rect 3234 14160 3268 14199
rect 3330 14233 3364 14272
rect 3330 14160 3364 14199
rect 3426 14233 3460 14272
rect 3426 14160 3460 14199
rect 3540 14203 3574 14236
rect 3647 14260 3681 14276
rect 3647 14168 3681 14184
rect 3735 14260 3769 14276
rect 3735 14168 3769 14184
rect 3873 14270 3907 14346
rect 5061 14275 5095 14346
rect 3873 14202 3907 14236
rect 3540 14134 3574 14168
rect 2352 14024 2386 14100
rect 2450 14088 2466 14122
rect 2500 14088 2516 14122
rect 2642 14088 2658 14122
rect 2692 14088 2708 14122
rect 2834 14088 2850 14122
rect 2884 14088 2900 14122
rect 3026 14088 3042 14122
rect 3076 14088 3092 14122
rect 3218 14088 3234 14122
rect 3268 14088 3284 14122
rect 3410 14088 3426 14122
rect 3460 14088 3476 14122
rect 3540 14024 3574 14097
rect 2352 13990 2470 14024
rect 2504 13990 2538 14024
rect 2572 13990 2606 14024
rect 2640 13990 2674 14024
rect 2708 13990 2742 14024
rect 2776 13990 2810 14024
rect 2844 13990 2878 14024
rect 2912 13990 2946 14024
rect 2980 13990 3014 14024
rect 3048 13990 3082 14024
rect 3116 13990 3150 14024
rect 3184 13990 3218 14024
rect 3252 13990 3286 14024
rect 3320 13990 3354 14024
rect 3388 13990 3422 14024
rect 3456 13990 3574 14024
rect 3873 14134 3907 14168
rect 3987 14233 4021 14272
rect 3987 14160 4021 14199
rect 4083 14233 4117 14272
rect 4083 14160 4117 14199
rect 4179 14233 4213 14272
rect 4179 14160 4213 14199
rect 4275 14233 4309 14272
rect 4275 14160 4309 14199
rect 4371 14233 4405 14272
rect 4371 14160 4405 14199
rect 4467 14233 4501 14272
rect 4467 14160 4501 14199
rect 4563 14233 4597 14272
rect 4563 14160 4597 14199
rect 4659 14233 4693 14272
rect 4659 14160 4693 14199
rect 4755 14233 4789 14272
rect 4755 14160 4789 14199
rect 4851 14233 4885 14272
rect 4851 14160 4885 14199
rect 4947 14233 4981 14272
rect 4947 14160 4981 14199
rect 5061 14203 5095 14236
rect 5340 14351 5348 14385
rect 5382 14351 5386 14385
rect 5420 14390 5486 14401
rect 5420 14387 5450 14390
rect 5420 14353 5436 14387
rect 5484 14356 5486 14390
rect 5470 14353 5486 14356
rect 5340 14315 5386 14351
rect 5340 14303 5406 14315
rect 5340 14269 5356 14303
rect 5390 14269 5406 14303
rect 5340 14235 5406 14269
rect 5340 14201 5356 14235
rect 5390 14201 5406 14235
rect 5340 14189 5406 14201
rect 5440 14303 5486 14319
rect 5474 14269 5486 14303
rect 5440 14235 5486 14269
rect 5474 14201 5486 14235
rect 5061 14134 5095 14168
rect 5440 14155 5486 14201
rect 3873 14024 3907 14100
rect 3971 14088 3987 14122
rect 4021 14088 4037 14122
rect 4163 14088 4179 14122
rect 4213 14088 4229 14122
rect 4355 14088 4371 14122
rect 4405 14088 4421 14122
rect 4547 14088 4563 14122
rect 4597 14088 4613 14122
rect 4739 14088 4755 14122
rect 4789 14088 4805 14122
rect 4931 14088 4947 14122
rect 4981 14088 4997 14122
rect 5274 14121 5303 14155
rect 5337 14121 5395 14155
rect 5429 14121 5487 14155
rect 5521 14121 5550 14155
rect 5061 14024 5095 14097
rect 3873 13990 3991 14024
rect 4025 13990 4059 14024
rect 4093 13990 4127 14024
rect 4161 13990 4195 14024
rect 4229 13990 4263 14024
rect 4297 13990 4331 14024
rect 4365 13990 4399 14024
rect 4433 13990 4467 14024
rect 4501 13990 4535 14024
rect 4569 13990 4603 14024
rect 4637 13990 4671 14024
rect 4705 13990 4739 14024
rect 4773 13990 4807 14024
rect 4841 13990 4875 14024
rect 4909 13990 4943 14024
rect 4977 13990 5095 14024
rect 199 13707 317 13741
rect 351 13707 385 13741
rect 419 13707 453 13741
rect 487 13707 521 13741
rect 555 13707 589 13741
rect 623 13707 657 13741
rect 691 13707 725 13741
rect 759 13707 793 13741
rect 827 13707 861 13741
rect 895 13707 929 13741
rect 963 13707 997 13741
rect 1031 13707 1065 13741
rect 1099 13707 1133 13741
rect 1167 13707 1201 13741
rect 1235 13707 1269 13741
rect 1303 13707 1421 13741
rect 199 13639 233 13707
rect 1387 13639 1421 13707
rect 297 13605 313 13639
rect 347 13605 363 13639
rect 489 13605 505 13639
rect 539 13605 555 13639
rect 681 13605 697 13639
rect 731 13605 747 13639
rect 873 13605 889 13639
rect 923 13605 939 13639
rect 1065 13605 1081 13639
rect 1115 13605 1131 13639
rect 1257 13605 1273 13639
rect 1307 13605 1323 13639
rect 199 13571 233 13605
rect 1387 13571 1421 13579
rect 199 13503 233 13537
rect 199 13435 233 13469
rect 199 13367 233 13401
rect 199 13299 233 13333
rect 313 13540 347 13561
rect 313 13472 347 13476
rect 313 13366 347 13370
rect 313 13281 347 13302
rect 409 13540 443 13561
rect 409 13472 443 13476
rect 409 13366 443 13370
rect 409 13281 443 13302
rect 505 13540 539 13561
rect 505 13472 539 13476
rect 505 13366 539 13370
rect 505 13281 539 13302
rect 601 13540 635 13561
rect 601 13472 635 13476
rect 601 13366 635 13370
rect 601 13281 635 13302
rect 697 13540 731 13561
rect 697 13472 731 13476
rect 697 13366 731 13370
rect 697 13281 731 13302
rect 793 13540 827 13561
rect 793 13472 827 13476
rect 793 13366 827 13370
rect 793 13281 827 13302
rect 889 13540 923 13561
rect 889 13472 923 13476
rect 889 13366 923 13370
rect 889 13281 923 13302
rect 985 13540 1019 13561
rect 985 13472 1019 13476
rect 985 13366 1019 13370
rect 985 13281 1019 13302
rect 1081 13540 1115 13561
rect 1081 13472 1115 13476
rect 1081 13366 1115 13370
rect 1081 13281 1115 13302
rect 1177 13540 1211 13561
rect 1177 13472 1211 13476
rect 1177 13366 1211 13370
rect 1177 13281 1211 13302
rect 1273 13540 1307 13561
rect 1273 13472 1307 13476
rect 1273 13366 1307 13370
rect 1273 13281 1307 13302
rect 1387 13503 1421 13507
rect 1387 13397 1421 13401
rect 1387 13325 1421 13333
rect 199 13197 233 13265
rect 1387 13197 1421 13265
rect 199 13163 317 13197
rect 351 13163 385 13197
rect 419 13163 453 13197
rect 487 13163 521 13197
rect 555 13163 589 13197
rect 623 13163 657 13197
rect 691 13163 725 13197
rect 759 13163 793 13197
rect 827 13163 861 13197
rect 895 13163 929 13197
rect 963 13163 997 13197
rect 1031 13163 1065 13197
rect 1099 13163 1133 13197
rect 1167 13163 1201 13197
rect 1235 13163 1269 13197
rect 1303 13163 1421 13197
rect 2352 13711 2470 13745
rect 2504 13711 2538 13745
rect 2572 13711 2606 13745
rect 2640 13711 2674 13745
rect 2708 13711 2742 13745
rect 2776 13711 2810 13745
rect 2844 13711 2878 13745
rect 2912 13711 2946 13745
rect 2980 13711 3014 13745
rect 3048 13711 3082 13745
rect 3116 13711 3150 13745
rect 3184 13711 3218 13745
rect 3252 13711 3286 13745
rect 3320 13711 3354 13745
rect 3388 13711 3422 13745
rect 3456 13711 3574 13745
rect 2352 13643 2386 13711
rect 3540 13643 3574 13711
rect 2450 13609 2466 13643
rect 2500 13609 2516 13643
rect 2642 13609 2658 13643
rect 2692 13609 2708 13643
rect 2834 13609 2850 13643
rect 2884 13609 2900 13643
rect 3026 13609 3042 13643
rect 3076 13609 3092 13643
rect 3218 13609 3234 13643
rect 3268 13609 3284 13643
rect 3410 13609 3426 13643
rect 3460 13609 3476 13643
rect 2352 13575 2386 13609
rect 3540 13575 3574 13583
rect 2352 13507 2386 13541
rect 2352 13439 2386 13473
rect 2352 13371 2386 13405
rect 2352 13303 2386 13337
rect 2466 13544 2500 13565
rect 2466 13476 2500 13480
rect 2466 13370 2500 13374
rect 2466 13285 2500 13306
rect 2562 13544 2596 13565
rect 2562 13476 2596 13480
rect 2562 13370 2596 13374
rect 2562 13285 2596 13306
rect 2658 13544 2692 13565
rect 2658 13476 2692 13480
rect 2658 13370 2692 13374
rect 2658 13285 2692 13306
rect 2754 13544 2788 13565
rect 2754 13476 2788 13480
rect 2754 13370 2788 13374
rect 2754 13285 2788 13306
rect 2850 13544 2884 13565
rect 2850 13476 2884 13480
rect 2850 13370 2884 13374
rect 2850 13285 2884 13306
rect 2946 13544 2980 13565
rect 2946 13476 2980 13480
rect 2946 13370 2980 13374
rect 2946 13285 2980 13306
rect 3042 13544 3076 13565
rect 3042 13476 3076 13480
rect 3042 13370 3076 13374
rect 3042 13285 3076 13306
rect 3138 13544 3172 13565
rect 3138 13476 3172 13480
rect 3138 13370 3172 13374
rect 3138 13285 3172 13306
rect 3234 13544 3268 13565
rect 3234 13476 3268 13480
rect 3234 13370 3268 13374
rect 3234 13285 3268 13306
rect 3330 13544 3364 13565
rect 3330 13476 3364 13480
rect 3330 13370 3364 13374
rect 3330 13285 3364 13306
rect 3426 13544 3460 13565
rect 3426 13476 3460 13480
rect 3426 13370 3460 13374
rect 3426 13285 3460 13306
rect 3540 13507 3574 13511
rect 3540 13401 3574 13405
rect 3540 13329 3574 13337
rect 2352 13201 2386 13269
rect 3540 13201 3574 13269
rect 2352 13167 2470 13201
rect 2504 13167 2538 13201
rect 2572 13167 2606 13201
rect 2640 13167 2674 13201
rect 2708 13167 2742 13201
rect 2776 13167 2810 13201
rect 2844 13167 2878 13201
rect 2912 13167 2946 13201
rect 2980 13167 3014 13201
rect 3048 13167 3082 13201
rect 3116 13167 3150 13201
rect 3184 13167 3218 13201
rect 3252 13167 3286 13201
rect 3320 13167 3354 13201
rect 3388 13167 3422 13201
rect 3456 13167 3574 13201
rect 3873 13711 3991 13745
rect 4025 13711 4059 13745
rect 4093 13711 4127 13745
rect 4161 13711 4195 13745
rect 4229 13711 4263 13745
rect 4297 13711 4331 13745
rect 4365 13711 4399 13745
rect 4433 13711 4467 13745
rect 4501 13711 4535 13745
rect 4569 13711 4603 13745
rect 4637 13711 4671 13745
rect 4705 13711 4739 13745
rect 4773 13711 4807 13745
rect 4841 13711 4875 13745
rect 4909 13711 4943 13745
rect 4977 13711 5095 13745
rect 3873 13643 3907 13711
rect 5061 13643 5095 13711
rect 3971 13609 3987 13643
rect 4021 13609 4037 13643
rect 4163 13609 4179 13643
rect 4213 13609 4229 13643
rect 4355 13609 4371 13643
rect 4405 13609 4421 13643
rect 4547 13609 4563 13643
rect 4597 13609 4613 13643
rect 4739 13609 4755 13643
rect 4789 13609 4805 13643
rect 4931 13609 4947 13643
rect 4981 13609 4997 13643
rect 3873 13575 3907 13609
rect 5061 13575 5095 13583
rect 3873 13507 3907 13541
rect 3873 13439 3907 13473
rect 3873 13371 3907 13405
rect 3873 13303 3907 13337
rect 3987 13544 4021 13565
rect 3987 13476 4021 13480
rect 3987 13370 4021 13374
rect 3987 13285 4021 13306
rect 4083 13544 4117 13565
rect 4083 13476 4117 13480
rect 4083 13370 4117 13374
rect 4083 13285 4117 13306
rect 4179 13544 4213 13565
rect 4179 13476 4213 13480
rect 4179 13370 4213 13374
rect 4179 13285 4213 13306
rect 4275 13544 4309 13565
rect 4275 13476 4309 13480
rect 4275 13370 4309 13374
rect 4275 13285 4309 13306
rect 4371 13544 4405 13565
rect 4371 13476 4405 13480
rect 4371 13370 4405 13374
rect 4371 13285 4405 13306
rect 4467 13544 4501 13565
rect 4467 13476 4501 13480
rect 4467 13370 4501 13374
rect 4467 13285 4501 13306
rect 4563 13544 4597 13565
rect 4563 13476 4597 13480
rect 4563 13370 4597 13374
rect 4563 13285 4597 13306
rect 4659 13544 4693 13565
rect 4659 13476 4693 13480
rect 4659 13370 4693 13374
rect 4659 13285 4693 13306
rect 4755 13544 4789 13565
rect 4755 13476 4789 13480
rect 4755 13370 4789 13374
rect 4755 13285 4789 13306
rect 4851 13544 4885 13565
rect 4851 13476 4885 13480
rect 4851 13370 4885 13374
rect 4851 13285 4885 13306
rect 4947 13544 4981 13565
rect 4947 13476 4981 13480
rect 4947 13370 4981 13374
rect 4947 13285 4981 13306
rect 5061 13507 5095 13511
rect 5061 13401 5095 13405
rect 5274 13378 5303 13412
rect 5337 13378 5395 13412
rect 5429 13378 5487 13412
rect 5521 13378 5550 13412
rect 5061 13329 5095 13337
rect 3873 13201 3907 13269
rect 5061 13201 5095 13269
rect 3873 13167 3991 13201
rect 4025 13167 4059 13201
rect 4093 13167 4127 13201
rect 4161 13167 4195 13201
rect 4229 13167 4263 13201
rect 4297 13167 4331 13201
rect 4365 13167 4399 13201
rect 4433 13167 4467 13201
rect 4501 13167 4535 13201
rect 4569 13167 4603 13201
rect 4637 13167 4671 13201
rect 4705 13167 4739 13201
rect 4773 13167 4807 13201
rect 4841 13167 4875 13201
rect 4909 13167 4943 13201
rect 4977 13167 5095 13201
rect 5340 13336 5406 13344
rect 5340 13302 5356 13336
rect 5390 13302 5406 13336
rect 5340 13268 5406 13302
rect 5340 13234 5356 13268
rect 5390 13234 5406 13268
rect 5340 13200 5406 13234
rect 5340 13166 5356 13200
rect 5390 13166 5406 13200
rect 5340 13148 5406 13166
rect 5440 13336 5482 13378
rect 5474 13302 5482 13336
rect 5440 13268 5482 13302
rect 5474 13234 5482 13268
rect 5440 13200 5482 13234
rect 5474 13166 5482 13200
rect 5440 13150 5482 13166
rect 5340 13098 5386 13148
rect 199 13055 317 13089
rect 351 13055 385 13089
rect 419 13055 453 13089
rect 487 13055 521 13089
rect 555 13055 589 13089
rect 623 13055 657 13089
rect 691 13055 725 13089
rect 759 13055 793 13089
rect 827 13055 861 13089
rect 895 13055 929 13089
rect 963 13055 997 13089
rect 1031 13055 1065 13089
rect 1099 13055 1133 13089
rect 1167 13055 1201 13089
rect 1235 13055 1269 13089
rect 1303 13055 1421 13089
rect 199 12979 233 13055
rect 1387 12984 1421 13055
rect 199 12911 233 12945
rect 199 12843 233 12877
rect 313 12942 347 12981
rect 313 12869 347 12908
rect 409 12942 443 12981
rect 409 12869 443 12908
rect 505 12942 539 12981
rect 505 12869 539 12908
rect 601 12942 635 12981
rect 601 12869 635 12908
rect 697 12942 731 12981
rect 697 12869 731 12908
rect 793 12942 827 12981
rect 793 12869 827 12908
rect 889 12942 923 12981
rect 889 12869 923 12908
rect 985 12942 1019 12981
rect 985 12869 1019 12908
rect 1081 12942 1115 12981
rect 1081 12869 1115 12908
rect 1177 12942 1211 12981
rect 1177 12869 1211 12908
rect 1273 12942 1307 12981
rect 1273 12869 1307 12908
rect 1387 12912 1421 12945
rect 1387 12843 1421 12877
rect 199 12733 233 12809
rect 297 12797 313 12831
rect 347 12797 363 12831
rect 489 12797 505 12831
rect 539 12797 555 12831
rect 681 12797 697 12831
rect 731 12797 747 12831
rect 873 12797 889 12831
rect 923 12797 939 12831
rect 1065 12797 1081 12831
rect 1115 12797 1131 12831
rect 1257 12797 1273 12831
rect 1307 12797 1323 12831
rect 1387 12733 1421 12806
rect 199 12699 317 12733
rect 351 12699 385 12733
rect 419 12699 453 12733
rect 487 12699 521 12733
rect 555 12699 589 12733
rect 623 12699 657 12733
rect 691 12699 725 12733
rect 759 12699 793 12733
rect 827 12699 861 12733
rect 895 12699 929 12733
rect 963 12699 997 12733
rect 1031 12699 1065 12733
rect 1099 12699 1133 12733
rect 1167 12699 1201 12733
rect 1235 12699 1269 12733
rect 1303 12699 1421 12733
rect 2352 13059 2470 13093
rect 2504 13059 2538 13093
rect 2572 13059 2606 13093
rect 2640 13059 2674 13093
rect 2708 13059 2742 13093
rect 2776 13059 2810 13093
rect 2844 13059 2878 13093
rect 2912 13059 2946 13093
rect 2980 13059 3014 13093
rect 3048 13059 3082 13093
rect 3116 13059 3150 13093
rect 3184 13059 3218 13093
rect 3252 13059 3286 13093
rect 3320 13059 3354 13093
rect 3388 13059 3422 13093
rect 3456 13059 3574 13093
rect 2352 12983 2386 13059
rect 3540 12988 3574 13059
rect 3873 13059 3991 13093
rect 4025 13059 4059 13093
rect 4093 13059 4127 13093
rect 4161 13059 4195 13093
rect 4229 13059 4263 13093
rect 4297 13059 4331 13093
rect 4365 13059 4399 13093
rect 4433 13059 4467 13093
rect 4501 13059 4535 13093
rect 4569 13059 4603 13093
rect 4637 13059 4671 13093
rect 4705 13059 4739 13093
rect 4773 13059 4807 13093
rect 4841 13059 4875 13093
rect 4909 13059 4943 13093
rect 4977 13059 5095 13093
rect 3675 13023 3691 13057
rect 3725 13023 3741 13057
rect 2352 12915 2386 12949
rect 2352 12847 2386 12881
rect 2466 12946 2500 12985
rect 2466 12873 2500 12912
rect 2562 12946 2596 12985
rect 2562 12873 2596 12912
rect 2658 12946 2692 12985
rect 2658 12873 2692 12912
rect 2754 12946 2788 12985
rect 2754 12873 2788 12912
rect 2850 12946 2884 12985
rect 2850 12873 2884 12912
rect 2946 12946 2980 12985
rect 2946 12873 2980 12912
rect 3042 12946 3076 12985
rect 3042 12873 3076 12912
rect 3138 12946 3172 12985
rect 3138 12873 3172 12912
rect 3234 12946 3268 12985
rect 3234 12873 3268 12912
rect 3330 12946 3364 12985
rect 3330 12873 3364 12912
rect 3426 12946 3460 12985
rect 3426 12873 3460 12912
rect 3540 12916 3574 12949
rect 3647 12973 3681 12989
rect 3647 12881 3681 12897
rect 3735 12973 3769 12989
rect 3735 12881 3769 12897
rect 3873 12983 3907 13059
rect 5061 12988 5095 13059
rect 3873 12915 3907 12949
rect 3540 12847 3574 12881
rect 2352 12737 2386 12813
rect 2450 12801 2466 12835
rect 2500 12801 2516 12835
rect 2642 12801 2658 12835
rect 2692 12801 2708 12835
rect 2834 12801 2850 12835
rect 2884 12801 2900 12835
rect 3026 12801 3042 12835
rect 3076 12801 3092 12835
rect 3218 12801 3234 12835
rect 3268 12801 3284 12835
rect 3410 12801 3426 12835
rect 3460 12801 3476 12835
rect 3540 12737 3574 12810
rect 2352 12703 2470 12737
rect 2504 12703 2538 12737
rect 2572 12703 2606 12737
rect 2640 12703 2674 12737
rect 2708 12703 2742 12737
rect 2776 12703 2810 12737
rect 2844 12703 2878 12737
rect 2912 12703 2946 12737
rect 2980 12703 3014 12737
rect 3048 12703 3082 12737
rect 3116 12703 3150 12737
rect 3184 12703 3218 12737
rect 3252 12703 3286 12737
rect 3320 12703 3354 12737
rect 3388 12703 3422 12737
rect 3456 12703 3574 12737
rect 3873 12847 3907 12881
rect 3987 12946 4021 12985
rect 3987 12873 4021 12912
rect 4083 12946 4117 12985
rect 4083 12873 4117 12912
rect 4179 12946 4213 12985
rect 4179 12873 4213 12912
rect 4275 12946 4309 12985
rect 4275 12873 4309 12912
rect 4371 12946 4405 12985
rect 4371 12873 4405 12912
rect 4467 12946 4501 12985
rect 4467 12873 4501 12912
rect 4563 12946 4597 12985
rect 4563 12873 4597 12912
rect 4659 12946 4693 12985
rect 4659 12873 4693 12912
rect 4755 12946 4789 12985
rect 4755 12873 4789 12912
rect 4851 12946 4885 12985
rect 4851 12873 4885 12912
rect 4947 12946 4981 12985
rect 4947 12873 4981 12912
rect 5061 12916 5095 12949
rect 5340 13064 5348 13098
rect 5382 13064 5386 13098
rect 5420 13103 5486 13114
rect 5420 13100 5450 13103
rect 5420 13066 5436 13100
rect 5484 13069 5486 13103
rect 5470 13066 5486 13069
rect 5340 13028 5386 13064
rect 5340 13016 5406 13028
rect 5340 12982 5356 13016
rect 5390 12982 5406 13016
rect 5340 12948 5406 12982
rect 5340 12914 5356 12948
rect 5390 12914 5406 12948
rect 5340 12902 5406 12914
rect 5440 13016 5486 13032
rect 5474 12982 5486 13016
rect 5440 12948 5486 12982
rect 5474 12914 5486 12948
rect 5061 12847 5095 12881
rect 5440 12868 5486 12914
rect 3873 12737 3907 12813
rect 3971 12801 3987 12835
rect 4021 12801 4037 12835
rect 4163 12801 4179 12835
rect 4213 12801 4229 12835
rect 4355 12801 4371 12835
rect 4405 12801 4421 12835
rect 4547 12801 4563 12835
rect 4597 12801 4613 12835
rect 4739 12801 4755 12835
rect 4789 12801 4805 12835
rect 4931 12801 4947 12835
rect 4981 12801 4997 12835
rect 5274 12834 5303 12868
rect 5337 12834 5395 12868
rect 5429 12834 5487 12868
rect 5521 12834 5550 12868
rect 5061 12737 5095 12810
rect 3873 12703 3991 12737
rect 4025 12703 4059 12737
rect 4093 12703 4127 12737
rect 4161 12703 4195 12737
rect 4229 12703 4263 12737
rect 4297 12703 4331 12737
rect 4365 12703 4399 12737
rect 4433 12703 4467 12737
rect 4501 12703 4535 12737
rect 4569 12703 4603 12737
rect 4637 12703 4671 12737
rect 4705 12703 4739 12737
rect 4773 12703 4807 12737
rect 4841 12703 4875 12737
rect 4909 12703 4943 12737
rect 4977 12703 5095 12737
rect 199 12420 317 12454
rect 351 12420 385 12454
rect 419 12420 453 12454
rect 487 12420 521 12454
rect 555 12420 589 12454
rect 623 12420 657 12454
rect 691 12420 725 12454
rect 759 12420 793 12454
rect 827 12420 861 12454
rect 895 12420 929 12454
rect 963 12420 997 12454
rect 1031 12420 1065 12454
rect 1099 12420 1133 12454
rect 1167 12420 1201 12454
rect 1235 12420 1269 12454
rect 1303 12420 1421 12454
rect 199 12352 233 12420
rect 1387 12352 1421 12420
rect 297 12318 313 12352
rect 347 12318 363 12352
rect 489 12318 505 12352
rect 539 12318 555 12352
rect 681 12318 697 12352
rect 731 12318 747 12352
rect 873 12318 889 12352
rect 923 12318 939 12352
rect 1065 12318 1081 12352
rect 1115 12318 1131 12352
rect 1257 12318 1273 12352
rect 1307 12318 1323 12352
rect 199 12284 233 12318
rect 1387 12284 1421 12292
rect 199 12216 233 12250
rect 199 12148 233 12182
rect 199 12080 233 12114
rect 199 12012 233 12046
rect 313 12253 347 12274
rect 313 12185 347 12189
rect 313 12079 347 12083
rect 313 11994 347 12015
rect 409 12253 443 12274
rect 409 12185 443 12189
rect 409 12079 443 12083
rect 409 11994 443 12015
rect 505 12253 539 12274
rect 505 12185 539 12189
rect 505 12079 539 12083
rect 505 11994 539 12015
rect 601 12253 635 12274
rect 601 12185 635 12189
rect 601 12079 635 12083
rect 601 11994 635 12015
rect 697 12253 731 12274
rect 697 12185 731 12189
rect 697 12079 731 12083
rect 697 11994 731 12015
rect 793 12253 827 12274
rect 793 12185 827 12189
rect 793 12079 827 12083
rect 793 11994 827 12015
rect 889 12253 923 12274
rect 889 12185 923 12189
rect 889 12079 923 12083
rect 889 11994 923 12015
rect 985 12253 1019 12274
rect 985 12185 1019 12189
rect 985 12079 1019 12083
rect 985 11994 1019 12015
rect 1081 12253 1115 12274
rect 1081 12185 1115 12189
rect 1081 12079 1115 12083
rect 1081 11994 1115 12015
rect 1177 12253 1211 12274
rect 1177 12185 1211 12189
rect 1177 12079 1211 12083
rect 1177 11994 1211 12015
rect 1273 12253 1307 12274
rect 1273 12185 1307 12189
rect 1273 12079 1307 12083
rect 1273 11994 1307 12015
rect 1387 12216 1421 12220
rect 1387 12110 1421 12114
rect 1387 12038 1421 12046
rect 199 11910 233 11978
rect 1387 11910 1421 11978
rect 199 11876 317 11910
rect 351 11876 385 11910
rect 419 11876 453 11910
rect 487 11876 521 11910
rect 555 11876 589 11910
rect 623 11876 657 11910
rect 691 11876 725 11910
rect 759 11876 793 11910
rect 827 11876 861 11910
rect 895 11876 929 11910
rect 963 11876 997 11910
rect 1031 11876 1065 11910
rect 1099 11876 1133 11910
rect 1167 11876 1201 11910
rect 1235 11876 1269 11910
rect 1303 11876 1421 11910
rect 2352 12424 2470 12458
rect 2504 12424 2538 12458
rect 2572 12424 2606 12458
rect 2640 12424 2674 12458
rect 2708 12424 2742 12458
rect 2776 12424 2810 12458
rect 2844 12424 2878 12458
rect 2912 12424 2946 12458
rect 2980 12424 3014 12458
rect 3048 12424 3082 12458
rect 3116 12424 3150 12458
rect 3184 12424 3218 12458
rect 3252 12424 3286 12458
rect 3320 12424 3354 12458
rect 3388 12424 3422 12458
rect 3456 12424 3574 12458
rect 2352 12356 2386 12424
rect 3540 12356 3574 12424
rect 2450 12322 2466 12356
rect 2500 12322 2516 12356
rect 2642 12322 2658 12356
rect 2692 12322 2708 12356
rect 2834 12322 2850 12356
rect 2884 12322 2900 12356
rect 3026 12322 3042 12356
rect 3076 12322 3092 12356
rect 3218 12322 3234 12356
rect 3268 12322 3284 12356
rect 3410 12322 3426 12356
rect 3460 12322 3476 12356
rect 2352 12288 2386 12322
rect 3540 12288 3574 12296
rect 2352 12220 2386 12254
rect 2352 12152 2386 12186
rect 2352 12084 2386 12118
rect 2352 12016 2386 12050
rect 2466 12257 2500 12278
rect 2466 12189 2500 12193
rect 2466 12083 2500 12087
rect 2466 11998 2500 12019
rect 2562 12257 2596 12278
rect 2562 12189 2596 12193
rect 2562 12083 2596 12087
rect 2562 11998 2596 12019
rect 2658 12257 2692 12278
rect 2658 12189 2692 12193
rect 2658 12083 2692 12087
rect 2658 11998 2692 12019
rect 2754 12257 2788 12278
rect 2754 12189 2788 12193
rect 2754 12083 2788 12087
rect 2754 11998 2788 12019
rect 2850 12257 2884 12278
rect 2850 12189 2884 12193
rect 2850 12083 2884 12087
rect 2850 11998 2884 12019
rect 2946 12257 2980 12278
rect 2946 12189 2980 12193
rect 2946 12083 2980 12087
rect 2946 11998 2980 12019
rect 3042 12257 3076 12278
rect 3042 12189 3076 12193
rect 3042 12083 3076 12087
rect 3042 11998 3076 12019
rect 3138 12257 3172 12278
rect 3138 12189 3172 12193
rect 3138 12083 3172 12087
rect 3138 11998 3172 12019
rect 3234 12257 3268 12278
rect 3234 12189 3268 12193
rect 3234 12083 3268 12087
rect 3234 11998 3268 12019
rect 3330 12257 3364 12278
rect 3330 12189 3364 12193
rect 3330 12083 3364 12087
rect 3330 11998 3364 12019
rect 3426 12257 3460 12278
rect 3426 12189 3460 12193
rect 3426 12083 3460 12087
rect 3426 11998 3460 12019
rect 3540 12220 3574 12224
rect 3540 12114 3574 12118
rect 3540 12042 3574 12050
rect 2352 11914 2386 11982
rect 3540 11914 3574 11982
rect 2352 11880 2470 11914
rect 2504 11880 2538 11914
rect 2572 11880 2606 11914
rect 2640 11880 2674 11914
rect 2708 11880 2742 11914
rect 2776 11880 2810 11914
rect 2844 11880 2878 11914
rect 2912 11880 2946 11914
rect 2980 11880 3014 11914
rect 3048 11880 3082 11914
rect 3116 11880 3150 11914
rect 3184 11880 3218 11914
rect 3252 11880 3286 11914
rect 3320 11880 3354 11914
rect 3388 11880 3422 11914
rect 3456 11880 3574 11914
rect 3873 12424 3991 12458
rect 4025 12424 4059 12458
rect 4093 12424 4127 12458
rect 4161 12424 4195 12458
rect 4229 12424 4263 12458
rect 4297 12424 4331 12458
rect 4365 12424 4399 12458
rect 4433 12424 4467 12458
rect 4501 12424 4535 12458
rect 4569 12424 4603 12458
rect 4637 12424 4671 12458
rect 4705 12424 4739 12458
rect 4773 12424 4807 12458
rect 4841 12424 4875 12458
rect 4909 12424 4943 12458
rect 4977 12424 5095 12458
rect 3873 12356 3907 12424
rect 5061 12356 5095 12424
rect 3971 12322 3987 12356
rect 4021 12322 4037 12356
rect 4163 12322 4179 12356
rect 4213 12322 4229 12356
rect 4355 12322 4371 12356
rect 4405 12322 4421 12356
rect 4547 12322 4563 12356
rect 4597 12322 4613 12356
rect 4739 12322 4755 12356
rect 4789 12322 4805 12356
rect 4931 12322 4947 12356
rect 4981 12322 4997 12356
rect 3873 12288 3907 12322
rect 5061 12288 5095 12296
rect 3873 12220 3907 12254
rect 3873 12152 3907 12186
rect 3873 12084 3907 12118
rect 3873 12016 3907 12050
rect 3987 12257 4021 12278
rect 3987 12189 4021 12193
rect 3987 12083 4021 12087
rect 3987 11998 4021 12019
rect 4083 12257 4117 12278
rect 4083 12189 4117 12193
rect 4083 12083 4117 12087
rect 4083 11998 4117 12019
rect 4179 12257 4213 12278
rect 4179 12189 4213 12193
rect 4179 12083 4213 12087
rect 4179 11998 4213 12019
rect 4275 12257 4309 12278
rect 4275 12189 4309 12193
rect 4275 12083 4309 12087
rect 4275 11998 4309 12019
rect 4371 12257 4405 12278
rect 4371 12189 4405 12193
rect 4371 12083 4405 12087
rect 4371 11998 4405 12019
rect 4467 12257 4501 12278
rect 4467 12189 4501 12193
rect 4467 12083 4501 12087
rect 4467 11998 4501 12019
rect 4563 12257 4597 12278
rect 4563 12189 4597 12193
rect 4563 12083 4597 12087
rect 4563 11998 4597 12019
rect 4659 12257 4693 12278
rect 4659 12189 4693 12193
rect 4659 12083 4693 12087
rect 4659 11998 4693 12019
rect 4755 12257 4789 12278
rect 4755 12189 4789 12193
rect 4755 12083 4789 12087
rect 4755 11998 4789 12019
rect 4851 12257 4885 12278
rect 4851 12189 4885 12193
rect 4851 12083 4885 12087
rect 4851 11998 4885 12019
rect 4947 12257 4981 12278
rect 4947 12189 4981 12193
rect 4947 12083 4981 12087
rect 4947 11998 4981 12019
rect 5061 12220 5095 12224
rect 5061 12114 5095 12118
rect 5274 12091 5303 12125
rect 5337 12091 5395 12125
rect 5429 12091 5487 12125
rect 5521 12091 5550 12125
rect 5061 12042 5095 12050
rect 3873 11914 3907 11982
rect 5061 11914 5095 11982
rect 3873 11880 3991 11914
rect 4025 11880 4059 11914
rect 4093 11880 4127 11914
rect 4161 11880 4195 11914
rect 4229 11880 4263 11914
rect 4297 11880 4331 11914
rect 4365 11880 4399 11914
rect 4433 11880 4467 11914
rect 4501 11880 4535 11914
rect 4569 11880 4603 11914
rect 4637 11880 4671 11914
rect 4705 11880 4739 11914
rect 4773 11880 4807 11914
rect 4841 11880 4875 11914
rect 4909 11880 4943 11914
rect 4977 11880 5095 11914
rect 5340 12049 5406 12057
rect 5340 12015 5356 12049
rect 5390 12015 5406 12049
rect 5340 11981 5406 12015
rect 5340 11947 5356 11981
rect 5390 11947 5406 11981
rect 5340 11913 5406 11947
rect 5340 11879 5356 11913
rect 5390 11879 5406 11913
rect 5340 11861 5406 11879
rect 5440 12049 5482 12091
rect 5474 12015 5482 12049
rect 5440 11981 5482 12015
rect 5474 11947 5482 11981
rect 5440 11913 5482 11947
rect 5474 11879 5482 11913
rect 5440 11863 5482 11879
rect 5340 11811 5386 11861
rect 199 11768 317 11802
rect 351 11768 385 11802
rect 419 11768 453 11802
rect 487 11768 521 11802
rect 555 11768 589 11802
rect 623 11768 657 11802
rect 691 11768 725 11802
rect 759 11768 793 11802
rect 827 11768 861 11802
rect 895 11768 929 11802
rect 963 11768 997 11802
rect 1031 11768 1065 11802
rect 1099 11768 1133 11802
rect 1167 11768 1201 11802
rect 1235 11768 1269 11802
rect 1303 11768 1421 11802
rect 199 11692 233 11768
rect 1387 11697 1421 11768
rect 199 11624 233 11658
rect 199 11556 233 11590
rect 313 11655 347 11694
rect 313 11582 347 11621
rect 409 11655 443 11694
rect 409 11582 443 11621
rect 505 11655 539 11694
rect 505 11582 539 11621
rect 601 11655 635 11694
rect 601 11582 635 11621
rect 697 11655 731 11694
rect 697 11582 731 11621
rect 793 11655 827 11694
rect 793 11582 827 11621
rect 889 11655 923 11694
rect 889 11582 923 11621
rect 985 11655 1019 11694
rect 985 11582 1019 11621
rect 1081 11655 1115 11694
rect 1081 11582 1115 11621
rect 1177 11655 1211 11694
rect 1177 11582 1211 11621
rect 1273 11655 1307 11694
rect 1273 11582 1307 11621
rect 1387 11625 1421 11658
rect 1387 11556 1421 11590
rect 199 11446 233 11522
rect 297 11510 313 11544
rect 347 11510 363 11544
rect 489 11510 505 11544
rect 539 11510 555 11544
rect 681 11510 697 11544
rect 731 11510 747 11544
rect 873 11510 889 11544
rect 923 11510 939 11544
rect 1065 11510 1081 11544
rect 1115 11510 1131 11544
rect 1257 11510 1273 11544
rect 1307 11510 1323 11544
rect 1387 11446 1421 11519
rect 199 11412 317 11446
rect 351 11412 385 11446
rect 419 11412 453 11446
rect 487 11412 521 11446
rect 555 11412 589 11446
rect 623 11412 657 11446
rect 691 11412 725 11446
rect 759 11412 793 11446
rect 827 11412 861 11446
rect 895 11412 929 11446
rect 963 11412 997 11446
rect 1031 11412 1065 11446
rect 1099 11412 1133 11446
rect 1167 11412 1201 11446
rect 1235 11412 1269 11446
rect 1303 11412 1421 11446
rect 2352 11772 2470 11806
rect 2504 11772 2538 11806
rect 2572 11772 2606 11806
rect 2640 11772 2674 11806
rect 2708 11772 2742 11806
rect 2776 11772 2810 11806
rect 2844 11772 2878 11806
rect 2912 11772 2946 11806
rect 2980 11772 3014 11806
rect 3048 11772 3082 11806
rect 3116 11772 3150 11806
rect 3184 11772 3218 11806
rect 3252 11772 3286 11806
rect 3320 11772 3354 11806
rect 3388 11772 3422 11806
rect 3456 11772 3574 11806
rect 2352 11696 2386 11772
rect 3540 11701 3574 11772
rect 3873 11772 3991 11806
rect 4025 11772 4059 11806
rect 4093 11772 4127 11806
rect 4161 11772 4195 11806
rect 4229 11772 4263 11806
rect 4297 11772 4331 11806
rect 4365 11772 4399 11806
rect 4433 11772 4467 11806
rect 4501 11772 4535 11806
rect 4569 11772 4603 11806
rect 4637 11772 4671 11806
rect 4705 11772 4739 11806
rect 4773 11772 4807 11806
rect 4841 11772 4875 11806
rect 4909 11772 4943 11806
rect 4977 11772 5095 11806
rect 3675 11736 3691 11770
rect 3725 11736 3741 11770
rect 2352 11628 2386 11662
rect 2352 11560 2386 11594
rect 2466 11659 2500 11698
rect 2466 11586 2500 11625
rect 2562 11659 2596 11698
rect 2562 11586 2596 11625
rect 2658 11659 2692 11698
rect 2658 11586 2692 11625
rect 2754 11659 2788 11698
rect 2754 11586 2788 11625
rect 2850 11659 2884 11698
rect 2850 11586 2884 11625
rect 2946 11659 2980 11698
rect 2946 11586 2980 11625
rect 3042 11659 3076 11698
rect 3042 11586 3076 11625
rect 3138 11659 3172 11698
rect 3138 11586 3172 11625
rect 3234 11659 3268 11698
rect 3234 11586 3268 11625
rect 3330 11659 3364 11698
rect 3330 11586 3364 11625
rect 3426 11659 3460 11698
rect 3426 11586 3460 11625
rect 3540 11629 3574 11662
rect 3647 11686 3681 11702
rect 3647 11594 3681 11610
rect 3735 11686 3769 11702
rect 3735 11594 3769 11610
rect 3873 11696 3907 11772
rect 5061 11701 5095 11772
rect 3873 11628 3907 11662
rect 3540 11560 3574 11594
rect 2352 11450 2386 11526
rect 2450 11514 2466 11548
rect 2500 11514 2516 11548
rect 2642 11514 2658 11548
rect 2692 11514 2708 11548
rect 2834 11514 2850 11548
rect 2884 11514 2900 11548
rect 3026 11514 3042 11548
rect 3076 11514 3092 11548
rect 3218 11514 3234 11548
rect 3268 11514 3284 11548
rect 3410 11514 3426 11548
rect 3460 11514 3476 11548
rect 3540 11450 3574 11523
rect 2352 11416 2470 11450
rect 2504 11416 2538 11450
rect 2572 11416 2606 11450
rect 2640 11416 2674 11450
rect 2708 11416 2742 11450
rect 2776 11416 2810 11450
rect 2844 11416 2878 11450
rect 2912 11416 2946 11450
rect 2980 11416 3014 11450
rect 3048 11416 3082 11450
rect 3116 11416 3150 11450
rect 3184 11416 3218 11450
rect 3252 11416 3286 11450
rect 3320 11416 3354 11450
rect 3388 11416 3422 11450
rect 3456 11416 3574 11450
rect 3873 11560 3907 11594
rect 3987 11659 4021 11698
rect 3987 11586 4021 11625
rect 4083 11659 4117 11698
rect 4083 11586 4117 11625
rect 4179 11659 4213 11698
rect 4179 11586 4213 11625
rect 4275 11659 4309 11698
rect 4275 11586 4309 11625
rect 4371 11659 4405 11698
rect 4371 11586 4405 11625
rect 4467 11659 4501 11698
rect 4467 11586 4501 11625
rect 4563 11659 4597 11698
rect 4563 11586 4597 11625
rect 4659 11659 4693 11698
rect 4659 11586 4693 11625
rect 4755 11659 4789 11698
rect 4755 11586 4789 11625
rect 4851 11659 4885 11698
rect 4851 11586 4885 11625
rect 4947 11659 4981 11698
rect 4947 11586 4981 11625
rect 5061 11629 5095 11662
rect 5340 11777 5348 11811
rect 5382 11777 5386 11811
rect 5420 11816 5486 11827
rect 5420 11813 5450 11816
rect 5420 11779 5436 11813
rect 5484 11782 5486 11816
rect 5470 11779 5486 11782
rect 5340 11741 5386 11777
rect 5340 11729 5406 11741
rect 5340 11695 5356 11729
rect 5390 11695 5406 11729
rect 5340 11661 5406 11695
rect 5340 11627 5356 11661
rect 5390 11627 5406 11661
rect 5340 11615 5406 11627
rect 5440 11729 5486 11745
rect 5474 11695 5486 11729
rect 5440 11661 5486 11695
rect 5474 11627 5486 11661
rect 5061 11560 5095 11594
rect 5440 11581 5486 11627
rect 3873 11450 3907 11526
rect 3971 11514 3987 11548
rect 4021 11514 4037 11548
rect 4163 11514 4179 11548
rect 4213 11514 4229 11548
rect 4355 11514 4371 11548
rect 4405 11514 4421 11548
rect 4547 11514 4563 11548
rect 4597 11514 4613 11548
rect 4739 11514 4755 11548
rect 4789 11514 4805 11548
rect 4931 11514 4947 11548
rect 4981 11514 4997 11548
rect 5274 11547 5303 11581
rect 5337 11547 5395 11581
rect 5429 11547 5487 11581
rect 5521 11547 5550 11581
rect 5061 11450 5095 11523
rect 3873 11416 3991 11450
rect 4025 11416 4059 11450
rect 4093 11416 4127 11450
rect 4161 11416 4195 11450
rect 4229 11416 4263 11450
rect 4297 11416 4331 11450
rect 4365 11416 4399 11450
rect 4433 11416 4467 11450
rect 4501 11416 4535 11450
rect 4569 11416 4603 11450
rect 4637 11416 4671 11450
rect 4705 11416 4739 11450
rect 4773 11416 4807 11450
rect 4841 11416 4875 11450
rect 4909 11416 4943 11450
rect 4977 11416 5095 11450
rect 199 11133 317 11167
rect 351 11133 385 11167
rect 419 11133 453 11167
rect 487 11133 521 11167
rect 555 11133 589 11167
rect 623 11133 657 11167
rect 691 11133 725 11167
rect 759 11133 793 11167
rect 827 11133 861 11167
rect 895 11133 929 11167
rect 963 11133 997 11167
rect 1031 11133 1065 11167
rect 1099 11133 1133 11167
rect 1167 11133 1201 11167
rect 1235 11133 1269 11167
rect 1303 11133 1421 11167
rect 199 11065 233 11133
rect 1387 11065 1421 11133
rect 297 11031 313 11065
rect 347 11031 363 11065
rect 489 11031 505 11065
rect 539 11031 555 11065
rect 681 11031 697 11065
rect 731 11031 747 11065
rect 873 11031 889 11065
rect 923 11031 939 11065
rect 1065 11031 1081 11065
rect 1115 11031 1131 11065
rect 1257 11031 1273 11065
rect 1307 11031 1323 11065
rect 199 10997 233 11031
rect 1387 10997 1421 11005
rect 199 10929 233 10963
rect 199 10861 233 10895
rect 199 10793 233 10827
rect 199 10725 233 10759
rect 313 10966 347 10987
rect 313 10898 347 10902
rect 313 10792 347 10796
rect 313 10707 347 10728
rect 409 10966 443 10987
rect 409 10898 443 10902
rect 409 10792 443 10796
rect 409 10707 443 10728
rect 505 10966 539 10987
rect 505 10898 539 10902
rect 505 10792 539 10796
rect 505 10707 539 10728
rect 601 10966 635 10987
rect 601 10898 635 10902
rect 601 10792 635 10796
rect 601 10707 635 10728
rect 697 10966 731 10987
rect 697 10898 731 10902
rect 697 10792 731 10796
rect 697 10707 731 10728
rect 793 10966 827 10987
rect 793 10898 827 10902
rect 793 10792 827 10796
rect 793 10707 827 10728
rect 889 10966 923 10987
rect 889 10898 923 10902
rect 889 10792 923 10796
rect 889 10707 923 10728
rect 985 10966 1019 10987
rect 985 10898 1019 10902
rect 985 10792 1019 10796
rect 985 10707 1019 10728
rect 1081 10966 1115 10987
rect 1081 10898 1115 10902
rect 1081 10792 1115 10796
rect 1081 10707 1115 10728
rect 1177 10966 1211 10987
rect 1177 10898 1211 10902
rect 1177 10792 1211 10796
rect 1177 10707 1211 10728
rect 1273 10966 1307 10987
rect 1273 10898 1307 10902
rect 1273 10792 1307 10796
rect 1273 10707 1307 10728
rect 1387 10929 1421 10933
rect 1387 10823 1421 10827
rect 1387 10751 1421 10759
rect 199 10623 233 10691
rect 1387 10623 1421 10691
rect 199 10589 317 10623
rect 351 10589 385 10623
rect 419 10589 453 10623
rect 487 10589 521 10623
rect 555 10589 589 10623
rect 623 10589 657 10623
rect 691 10589 725 10623
rect 759 10589 793 10623
rect 827 10589 861 10623
rect 895 10589 929 10623
rect 963 10589 997 10623
rect 1031 10589 1065 10623
rect 1099 10589 1133 10623
rect 1167 10589 1201 10623
rect 1235 10589 1269 10623
rect 1303 10589 1421 10623
rect 2352 11137 2470 11171
rect 2504 11137 2538 11171
rect 2572 11137 2606 11171
rect 2640 11137 2674 11171
rect 2708 11137 2742 11171
rect 2776 11137 2810 11171
rect 2844 11137 2878 11171
rect 2912 11137 2946 11171
rect 2980 11137 3014 11171
rect 3048 11137 3082 11171
rect 3116 11137 3150 11171
rect 3184 11137 3218 11171
rect 3252 11137 3286 11171
rect 3320 11137 3354 11171
rect 3388 11137 3422 11171
rect 3456 11137 3574 11171
rect 2352 11069 2386 11137
rect 3540 11069 3574 11137
rect 2450 11035 2466 11069
rect 2500 11035 2516 11069
rect 2642 11035 2658 11069
rect 2692 11035 2708 11069
rect 2834 11035 2850 11069
rect 2884 11035 2900 11069
rect 3026 11035 3042 11069
rect 3076 11035 3092 11069
rect 3218 11035 3234 11069
rect 3268 11035 3284 11069
rect 3410 11035 3426 11069
rect 3460 11035 3476 11069
rect 2352 11001 2386 11035
rect 3540 11001 3574 11009
rect 2352 10933 2386 10967
rect 2352 10865 2386 10899
rect 2352 10797 2386 10831
rect 2352 10729 2386 10763
rect 2466 10970 2500 10991
rect 2466 10902 2500 10906
rect 2466 10796 2500 10800
rect 2466 10711 2500 10732
rect 2562 10970 2596 10991
rect 2562 10902 2596 10906
rect 2562 10796 2596 10800
rect 2562 10711 2596 10732
rect 2658 10970 2692 10991
rect 2658 10902 2692 10906
rect 2658 10796 2692 10800
rect 2658 10711 2692 10732
rect 2754 10970 2788 10991
rect 2754 10902 2788 10906
rect 2754 10796 2788 10800
rect 2754 10711 2788 10732
rect 2850 10970 2884 10991
rect 2850 10902 2884 10906
rect 2850 10796 2884 10800
rect 2850 10711 2884 10732
rect 2946 10970 2980 10991
rect 2946 10902 2980 10906
rect 2946 10796 2980 10800
rect 2946 10711 2980 10732
rect 3042 10970 3076 10991
rect 3042 10902 3076 10906
rect 3042 10796 3076 10800
rect 3042 10711 3076 10732
rect 3138 10970 3172 10991
rect 3138 10902 3172 10906
rect 3138 10796 3172 10800
rect 3138 10711 3172 10732
rect 3234 10970 3268 10991
rect 3234 10902 3268 10906
rect 3234 10796 3268 10800
rect 3234 10711 3268 10732
rect 3330 10970 3364 10991
rect 3330 10902 3364 10906
rect 3330 10796 3364 10800
rect 3330 10711 3364 10732
rect 3426 10970 3460 10991
rect 3426 10902 3460 10906
rect 3426 10796 3460 10800
rect 3426 10711 3460 10732
rect 3540 10933 3574 10937
rect 3540 10827 3574 10831
rect 3540 10755 3574 10763
rect 2352 10627 2386 10695
rect 3540 10627 3574 10695
rect 2352 10593 2470 10627
rect 2504 10593 2538 10627
rect 2572 10593 2606 10627
rect 2640 10593 2674 10627
rect 2708 10593 2742 10627
rect 2776 10593 2810 10627
rect 2844 10593 2878 10627
rect 2912 10593 2946 10627
rect 2980 10593 3014 10627
rect 3048 10593 3082 10627
rect 3116 10593 3150 10627
rect 3184 10593 3218 10627
rect 3252 10593 3286 10627
rect 3320 10593 3354 10627
rect 3388 10593 3422 10627
rect 3456 10593 3574 10627
rect 3873 11137 3991 11171
rect 4025 11137 4059 11171
rect 4093 11137 4127 11171
rect 4161 11137 4195 11171
rect 4229 11137 4263 11171
rect 4297 11137 4331 11171
rect 4365 11137 4399 11171
rect 4433 11137 4467 11171
rect 4501 11137 4535 11171
rect 4569 11137 4603 11171
rect 4637 11137 4671 11171
rect 4705 11137 4739 11171
rect 4773 11137 4807 11171
rect 4841 11137 4875 11171
rect 4909 11137 4943 11171
rect 4977 11137 5095 11171
rect 3873 11069 3907 11137
rect 5061 11069 5095 11137
rect 3971 11035 3987 11069
rect 4021 11035 4037 11069
rect 4163 11035 4179 11069
rect 4213 11035 4229 11069
rect 4355 11035 4371 11069
rect 4405 11035 4421 11069
rect 4547 11035 4563 11069
rect 4597 11035 4613 11069
rect 4739 11035 4755 11069
rect 4789 11035 4805 11069
rect 4931 11035 4947 11069
rect 4981 11035 4997 11069
rect 3873 11001 3907 11035
rect 5061 11001 5095 11009
rect 3873 10933 3907 10967
rect 3873 10865 3907 10899
rect 3873 10797 3907 10831
rect 3873 10729 3907 10763
rect 3987 10970 4021 10991
rect 3987 10902 4021 10906
rect 3987 10796 4021 10800
rect 3987 10711 4021 10732
rect 4083 10970 4117 10991
rect 4083 10902 4117 10906
rect 4083 10796 4117 10800
rect 4083 10711 4117 10732
rect 4179 10970 4213 10991
rect 4179 10902 4213 10906
rect 4179 10796 4213 10800
rect 4179 10711 4213 10732
rect 4275 10970 4309 10991
rect 4275 10902 4309 10906
rect 4275 10796 4309 10800
rect 4275 10711 4309 10732
rect 4371 10970 4405 10991
rect 4371 10902 4405 10906
rect 4371 10796 4405 10800
rect 4371 10711 4405 10732
rect 4467 10970 4501 10991
rect 4467 10902 4501 10906
rect 4467 10796 4501 10800
rect 4467 10711 4501 10732
rect 4563 10970 4597 10991
rect 4563 10902 4597 10906
rect 4563 10796 4597 10800
rect 4563 10711 4597 10732
rect 4659 10970 4693 10991
rect 4659 10902 4693 10906
rect 4659 10796 4693 10800
rect 4659 10711 4693 10732
rect 4755 10970 4789 10991
rect 4755 10902 4789 10906
rect 4755 10796 4789 10800
rect 4755 10711 4789 10732
rect 4851 10970 4885 10991
rect 4851 10902 4885 10906
rect 4851 10796 4885 10800
rect 4851 10711 4885 10732
rect 4947 10970 4981 10991
rect 4947 10902 4981 10906
rect 4947 10796 4981 10800
rect 4947 10711 4981 10732
rect 5061 10933 5095 10937
rect 5061 10827 5095 10831
rect 5274 10804 5303 10838
rect 5337 10804 5395 10838
rect 5429 10804 5487 10838
rect 5521 10804 5550 10838
rect 5061 10755 5095 10763
rect 3873 10627 3907 10695
rect 5061 10627 5095 10695
rect 3873 10593 3991 10627
rect 4025 10593 4059 10627
rect 4093 10593 4127 10627
rect 4161 10593 4195 10627
rect 4229 10593 4263 10627
rect 4297 10593 4331 10627
rect 4365 10593 4399 10627
rect 4433 10593 4467 10627
rect 4501 10593 4535 10627
rect 4569 10593 4603 10627
rect 4637 10593 4671 10627
rect 4705 10593 4739 10627
rect 4773 10593 4807 10627
rect 4841 10593 4875 10627
rect 4909 10593 4943 10627
rect 4977 10593 5095 10627
rect 5340 10762 5406 10770
rect 5340 10728 5356 10762
rect 5390 10728 5406 10762
rect 5340 10694 5406 10728
rect 5340 10660 5356 10694
rect 5390 10660 5406 10694
rect 5340 10626 5406 10660
rect 5340 10592 5356 10626
rect 5390 10592 5406 10626
rect 5340 10574 5406 10592
rect 5440 10762 5482 10804
rect 5474 10728 5482 10762
rect 5440 10694 5482 10728
rect 5474 10660 5482 10694
rect 5440 10626 5482 10660
rect 5474 10592 5482 10626
rect 5440 10576 5482 10592
rect 5340 10524 5386 10574
rect 199 10481 317 10515
rect 351 10481 385 10515
rect 419 10481 453 10515
rect 487 10481 521 10515
rect 555 10481 589 10515
rect 623 10481 657 10515
rect 691 10481 725 10515
rect 759 10481 793 10515
rect 827 10481 861 10515
rect 895 10481 929 10515
rect 963 10481 997 10515
rect 1031 10481 1065 10515
rect 1099 10481 1133 10515
rect 1167 10481 1201 10515
rect 1235 10481 1269 10515
rect 1303 10481 1421 10515
rect 199 10405 233 10481
rect 1387 10410 1421 10481
rect 199 10337 233 10371
rect 199 10269 233 10303
rect 313 10368 347 10407
rect 313 10295 347 10334
rect 409 10368 443 10407
rect 409 10295 443 10334
rect 505 10368 539 10407
rect 505 10295 539 10334
rect 601 10368 635 10407
rect 601 10295 635 10334
rect 697 10368 731 10407
rect 697 10295 731 10334
rect 793 10368 827 10407
rect 793 10295 827 10334
rect 889 10368 923 10407
rect 889 10295 923 10334
rect 985 10368 1019 10407
rect 985 10295 1019 10334
rect 1081 10368 1115 10407
rect 1081 10295 1115 10334
rect 1177 10368 1211 10407
rect 1177 10295 1211 10334
rect 1273 10368 1307 10407
rect 1273 10295 1307 10334
rect 1387 10338 1421 10371
rect 1387 10269 1421 10303
rect 199 10159 233 10235
rect 297 10223 313 10257
rect 347 10223 363 10257
rect 489 10223 505 10257
rect 539 10223 555 10257
rect 681 10223 697 10257
rect 731 10223 747 10257
rect 873 10223 889 10257
rect 923 10223 939 10257
rect 1065 10223 1081 10257
rect 1115 10223 1131 10257
rect 1257 10223 1273 10257
rect 1307 10223 1323 10257
rect 1387 10159 1421 10232
rect 199 10125 317 10159
rect 351 10125 385 10159
rect 419 10125 453 10159
rect 487 10125 521 10159
rect 555 10125 589 10159
rect 623 10125 657 10159
rect 691 10125 725 10159
rect 759 10125 793 10159
rect 827 10125 861 10159
rect 895 10125 929 10159
rect 963 10125 997 10159
rect 1031 10125 1065 10159
rect 1099 10125 1133 10159
rect 1167 10125 1201 10159
rect 1235 10125 1269 10159
rect 1303 10125 1421 10159
rect 2352 10485 2470 10519
rect 2504 10485 2538 10519
rect 2572 10485 2606 10519
rect 2640 10485 2674 10519
rect 2708 10485 2742 10519
rect 2776 10485 2810 10519
rect 2844 10485 2878 10519
rect 2912 10485 2946 10519
rect 2980 10485 3014 10519
rect 3048 10485 3082 10519
rect 3116 10485 3150 10519
rect 3184 10485 3218 10519
rect 3252 10485 3286 10519
rect 3320 10485 3354 10519
rect 3388 10485 3422 10519
rect 3456 10485 3574 10519
rect 2352 10409 2386 10485
rect 3540 10414 3574 10485
rect 3873 10485 3991 10519
rect 4025 10485 4059 10519
rect 4093 10485 4127 10519
rect 4161 10485 4195 10519
rect 4229 10485 4263 10519
rect 4297 10485 4331 10519
rect 4365 10485 4399 10519
rect 4433 10485 4467 10519
rect 4501 10485 4535 10519
rect 4569 10485 4603 10519
rect 4637 10485 4671 10519
rect 4705 10485 4739 10519
rect 4773 10485 4807 10519
rect 4841 10485 4875 10519
rect 4909 10485 4943 10519
rect 4977 10485 5095 10519
rect 3675 10449 3691 10483
rect 3725 10449 3741 10483
rect 2352 10341 2386 10375
rect 2352 10273 2386 10307
rect 2466 10372 2500 10411
rect 2466 10299 2500 10338
rect 2562 10372 2596 10411
rect 2562 10299 2596 10338
rect 2658 10372 2692 10411
rect 2658 10299 2692 10338
rect 2754 10372 2788 10411
rect 2754 10299 2788 10338
rect 2850 10372 2884 10411
rect 2850 10299 2884 10338
rect 2946 10372 2980 10411
rect 2946 10299 2980 10338
rect 3042 10372 3076 10411
rect 3042 10299 3076 10338
rect 3138 10372 3172 10411
rect 3138 10299 3172 10338
rect 3234 10372 3268 10411
rect 3234 10299 3268 10338
rect 3330 10372 3364 10411
rect 3330 10299 3364 10338
rect 3426 10372 3460 10411
rect 3426 10299 3460 10338
rect 3540 10342 3574 10375
rect 3647 10399 3681 10415
rect 3647 10307 3681 10323
rect 3735 10399 3769 10415
rect 3735 10307 3769 10323
rect 3873 10409 3907 10485
rect 5061 10414 5095 10485
rect 3873 10341 3907 10375
rect 3540 10273 3574 10307
rect 2352 10163 2386 10239
rect 2450 10227 2466 10261
rect 2500 10227 2516 10261
rect 2642 10227 2658 10261
rect 2692 10227 2708 10261
rect 2834 10227 2850 10261
rect 2884 10227 2900 10261
rect 3026 10227 3042 10261
rect 3076 10227 3092 10261
rect 3218 10227 3234 10261
rect 3268 10227 3284 10261
rect 3410 10227 3426 10261
rect 3460 10227 3476 10261
rect 3540 10163 3574 10236
rect 2352 10129 2470 10163
rect 2504 10129 2538 10163
rect 2572 10129 2606 10163
rect 2640 10129 2674 10163
rect 2708 10129 2742 10163
rect 2776 10129 2810 10163
rect 2844 10129 2878 10163
rect 2912 10129 2946 10163
rect 2980 10129 3014 10163
rect 3048 10129 3082 10163
rect 3116 10129 3150 10163
rect 3184 10129 3218 10163
rect 3252 10129 3286 10163
rect 3320 10129 3354 10163
rect 3388 10129 3422 10163
rect 3456 10129 3574 10163
rect 3873 10273 3907 10307
rect 3987 10372 4021 10411
rect 3987 10299 4021 10338
rect 4083 10372 4117 10411
rect 4083 10299 4117 10338
rect 4179 10372 4213 10411
rect 4179 10299 4213 10338
rect 4275 10372 4309 10411
rect 4275 10299 4309 10338
rect 4371 10372 4405 10411
rect 4371 10299 4405 10338
rect 4467 10372 4501 10411
rect 4467 10299 4501 10338
rect 4563 10372 4597 10411
rect 4563 10299 4597 10338
rect 4659 10372 4693 10411
rect 4659 10299 4693 10338
rect 4755 10372 4789 10411
rect 4755 10299 4789 10338
rect 4851 10372 4885 10411
rect 4851 10299 4885 10338
rect 4947 10372 4981 10411
rect 4947 10299 4981 10338
rect 5061 10342 5095 10375
rect 5340 10490 5348 10524
rect 5382 10490 5386 10524
rect 5420 10529 5486 10540
rect 5420 10526 5450 10529
rect 5420 10492 5436 10526
rect 5484 10495 5486 10529
rect 5470 10492 5486 10495
rect 5340 10454 5386 10490
rect 5340 10442 5406 10454
rect 5340 10408 5356 10442
rect 5390 10408 5406 10442
rect 5340 10374 5406 10408
rect 5340 10340 5356 10374
rect 5390 10340 5406 10374
rect 5340 10328 5406 10340
rect 5440 10442 5486 10458
rect 5474 10408 5486 10442
rect 5440 10374 5486 10408
rect 5474 10340 5486 10374
rect 5061 10273 5095 10307
rect 5440 10294 5486 10340
rect 3873 10163 3907 10239
rect 3971 10227 3987 10261
rect 4021 10227 4037 10261
rect 4163 10227 4179 10261
rect 4213 10227 4229 10261
rect 4355 10227 4371 10261
rect 4405 10227 4421 10261
rect 4547 10227 4563 10261
rect 4597 10227 4613 10261
rect 4739 10227 4755 10261
rect 4789 10227 4805 10261
rect 4931 10227 4947 10261
rect 4981 10227 4997 10261
rect 5274 10260 5303 10294
rect 5337 10260 5395 10294
rect 5429 10260 5487 10294
rect 5521 10260 5550 10294
rect 5061 10163 5095 10236
rect 3873 10129 3991 10163
rect 4025 10129 4059 10163
rect 4093 10129 4127 10163
rect 4161 10129 4195 10163
rect 4229 10129 4263 10163
rect 4297 10129 4331 10163
rect 4365 10129 4399 10163
rect 4433 10129 4467 10163
rect 4501 10129 4535 10163
rect 4569 10129 4603 10163
rect 4637 10129 4671 10163
rect 4705 10129 4739 10163
rect 4773 10129 4807 10163
rect 4841 10129 4875 10163
rect 4909 10129 4943 10163
rect 4977 10129 5095 10163
rect 199 9846 317 9880
rect 351 9846 385 9880
rect 419 9846 453 9880
rect 487 9846 521 9880
rect 555 9846 589 9880
rect 623 9846 657 9880
rect 691 9846 725 9880
rect 759 9846 793 9880
rect 827 9846 861 9880
rect 895 9846 929 9880
rect 963 9846 997 9880
rect 1031 9846 1065 9880
rect 1099 9846 1133 9880
rect 1167 9846 1201 9880
rect 1235 9846 1269 9880
rect 1303 9846 1421 9880
rect 199 9778 233 9846
rect 1387 9778 1421 9846
rect 297 9744 313 9778
rect 347 9744 363 9778
rect 489 9744 505 9778
rect 539 9744 555 9778
rect 681 9744 697 9778
rect 731 9744 747 9778
rect 873 9744 889 9778
rect 923 9744 939 9778
rect 1065 9744 1081 9778
rect 1115 9744 1131 9778
rect 1257 9744 1273 9778
rect 1307 9744 1323 9778
rect 199 9710 233 9744
rect 1387 9710 1421 9718
rect 199 9642 233 9676
rect 199 9574 233 9608
rect 199 9506 233 9540
rect 199 9438 233 9472
rect 313 9679 347 9700
rect 313 9611 347 9615
rect 313 9505 347 9509
rect 313 9420 347 9441
rect 409 9679 443 9700
rect 409 9611 443 9615
rect 409 9505 443 9509
rect 409 9420 443 9441
rect 505 9679 539 9700
rect 505 9611 539 9615
rect 505 9505 539 9509
rect 505 9420 539 9441
rect 601 9679 635 9700
rect 601 9611 635 9615
rect 601 9505 635 9509
rect 601 9420 635 9441
rect 697 9679 731 9700
rect 697 9611 731 9615
rect 697 9505 731 9509
rect 697 9420 731 9441
rect 793 9679 827 9700
rect 793 9611 827 9615
rect 793 9505 827 9509
rect 793 9420 827 9441
rect 889 9679 923 9700
rect 889 9611 923 9615
rect 889 9505 923 9509
rect 889 9420 923 9441
rect 985 9679 1019 9700
rect 985 9611 1019 9615
rect 985 9505 1019 9509
rect 985 9420 1019 9441
rect 1081 9679 1115 9700
rect 1081 9611 1115 9615
rect 1081 9505 1115 9509
rect 1081 9420 1115 9441
rect 1177 9679 1211 9700
rect 1177 9611 1211 9615
rect 1177 9505 1211 9509
rect 1177 9420 1211 9441
rect 1273 9679 1307 9700
rect 1273 9611 1307 9615
rect 1273 9505 1307 9509
rect 1273 9420 1307 9441
rect 1387 9642 1421 9646
rect 1387 9536 1421 9540
rect 1387 9464 1421 9472
rect 199 9336 233 9404
rect 1387 9336 1421 9404
rect 199 9302 317 9336
rect 351 9302 385 9336
rect 419 9302 453 9336
rect 487 9302 521 9336
rect 555 9302 589 9336
rect 623 9302 657 9336
rect 691 9302 725 9336
rect 759 9302 793 9336
rect 827 9302 861 9336
rect 895 9302 929 9336
rect 963 9302 997 9336
rect 1031 9302 1065 9336
rect 1099 9302 1133 9336
rect 1167 9302 1201 9336
rect 1235 9302 1269 9336
rect 1303 9302 1421 9336
rect 2352 9850 2470 9884
rect 2504 9850 2538 9884
rect 2572 9850 2606 9884
rect 2640 9850 2674 9884
rect 2708 9850 2742 9884
rect 2776 9850 2810 9884
rect 2844 9850 2878 9884
rect 2912 9850 2946 9884
rect 2980 9850 3014 9884
rect 3048 9850 3082 9884
rect 3116 9850 3150 9884
rect 3184 9850 3218 9884
rect 3252 9850 3286 9884
rect 3320 9850 3354 9884
rect 3388 9850 3422 9884
rect 3456 9850 3574 9884
rect 2352 9782 2386 9850
rect 3540 9782 3574 9850
rect 2450 9748 2466 9782
rect 2500 9748 2516 9782
rect 2642 9748 2658 9782
rect 2692 9748 2708 9782
rect 2834 9748 2850 9782
rect 2884 9748 2900 9782
rect 3026 9748 3042 9782
rect 3076 9748 3092 9782
rect 3218 9748 3234 9782
rect 3268 9748 3284 9782
rect 3410 9748 3426 9782
rect 3460 9748 3476 9782
rect 2352 9714 2386 9748
rect 3540 9714 3574 9722
rect 2352 9646 2386 9680
rect 2352 9578 2386 9612
rect 2352 9510 2386 9544
rect 2352 9442 2386 9476
rect 2466 9683 2500 9704
rect 2466 9615 2500 9619
rect 2466 9509 2500 9513
rect 2466 9424 2500 9445
rect 2562 9683 2596 9704
rect 2562 9615 2596 9619
rect 2562 9509 2596 9513
rect 2562 9424 2596 9445
rect 2658 9683 2692 9704
rect 2658 9615 2692 9619
rect 2658 9509 2692 9513
rect 2658 9424 2692 9445
rect 2754 9683 2788 9704
rect 2754 9615 2788 9619
rect 2754 9509 2788 9513
rect 2754 9424 2788 9445
rect 2850 9683 2884 9704
rect 2850 9615 2884 9619
rect 2850 9509 2884 9513
rect 2850 9424 2884 9445
rect 2946 9683 2980 9704
rect 2946 9615 2980 9619
rect 2946 9509 2980 9513
rect 2946 9424 2980 9445
rect 3042 9683 3076 9704
rect 3042 9615 3076 9619
rect 3042 9509 3076 9513
rect 3042 9424 3076 9445
rect 3138 9683 3172 9704
rect 3138 9615 3172 9619
rect 3138 9509 3172 9513
rect 3138 9424 3172 9445
rect 3234 9683 3268 9704
rect 3234 9615 3268 9619
rect 3234 9509 3268 9513
rect 3234 9424 3268 9445
rect 3330 9683 3364 9704
rect 3330 9615 3364 9619
rect 3330 9509 3364 9513
rect 3330 9424 3364 9445
rect 3426 9683 3460 9704
rect 3426 9615 3460 9619
rect 3426 9509 3460 9513
rect 3426 9424 3460 9445
rect 3540 9646 3574 9650
rect 3540 9540 3574 9544
rect 3540 9468 3574 9476
rect 2352 9340 2386 9408
rect 3540 9340 3574 9408
rect 2352 9306 2470 9340
rect 2504 9306 2538 9340
rect 2572 9306 2606 9340
rect 2640 9306 2674 9340
rect 2708 9306 2742 9340
rect 2776 9306 2810 9340
rect 2844 9306 2878 9340
rect 2912 9306 2946 9340
rect 2980 9306 3014 9340
rect 3048 9306 3082 9340
rect 3116 9306 3150 9340
rect 3184 9306 3218 9340
rect 3252 9306 3286 9340
rect 3320 9306 3354 9340
rect 3388 9306 3422 9340
rect 3456 9306 3574 9340
rect 3873 9850 3991 9884
rect 4025 9850 4059 9884
rect 4093 9850 4127 9884
rect 4161 9850 4195 9884
rect 4229 9850 4263 9884
rect 4297 9850 4331 9884
rect 4365 9850 4399 9884
rect 4433 9850 4467 9884
rect 4501 9850 4535 9884
rect 4569 9850 4603 9884
rect 4637 9850 4671 9884
rect 4705 9850 4739 9884
rect 4773 9850 4807 9884
rect 4841 9850 4875 9884
rect 4909 9850 4943 9884
rect 4977 9850 5095 9884
rect 3873 9782 3907 9850
rect 5061 9782 5095 9850
rect 3971 9748 3987 9782
rect 4021 9748 4037 9782
rect 4163 9748 4179 9782
rect 4213 9748 4229 9782
rect 4355 9748 4371 9782
rect 4405 9748 4421 9782
rect 4547 9748 4563 9782
rect 4597 9748 4613 9782
rect 4739 9748 4755 9782
rect 4789 9748 4805 9782
rect 4931 9748 4947 9782
rect 4981 9748 4997 9782
rect 3873 9714 3907 9748
rect 5061 9714 5095 9722
rect 3873 9646 3907 9680
rect 3873 9578 3907 9612
rect 3873 9510 3907 9544
rect 3873 9442 3907 9476
rect 3987 9683 4021 9704
rect 3987 9615 4021 9619
rect 3987 9509 4021 9513
rect 3987 9424 4021 9445
rect 4083 9683 4117 9704
rect 4083 9615 4117 9619
rect 4083 9509 4117 9513
rect 4083 9424 4117 9445
rect 4179 9683 4213 9704
rect 4179 9615 4213 9619
rect 4179 9509 4213 9513
rect 4179 9424 4213 9445
rect 4275 9683 4309 9704
rect 4275 9615 4309 9619
rect 4275 9509 4309 9513
rect 4275 9424 4309 9445
rect 4371 9683 4405 9704
rect 4371 9615 4405 9619
rect 4371 9509 4405 9513
rect 4371 9424 4405 9445
rect 4467 9683 4501 9704
rect 4467 9615 4501 9619
rect 4467 9509 4501 9513
rect 4467 9424 4501 9445
rect 4563 9683 4597 9704
rect 4563 9615 4597 9619
rect 4563 9509 4597 9513
rect 4563 9424 4597 9445
rect 4659 9683 4693 9704
rect 4659 9615 4693 9619
rect 4659 9509 4693 9513
rect 4659 9424 4693 9445
rect 4755 9683 4789 9704
rect 4755 9615 4789 9619
rect 4755 9509 4789 9513
rect 4755 9424 4789 9445
rect 4851 9683 4885 9704
rect 4851 9615 4885 9619
rect 4851 9509 4885 9513
rect 4851 9424 4885 9445
rect 4947 9683 4981 9704
rect 4947 9615 4981 9619
rect 4947 9509 4981 9513
rect 4947 9424 4981 9445
rect 5061 9646 5095 9650
rect 5061 9540 5095 9544
rect 5274 9517 5303 9551
rect 5337 9517 5395 9551
rect 5429 9517 5487 9551
rect 5521 9517 5550 9551
rect 5061 9468 5095 9476
rect 3873 9340 3907 9408
rect 5061 9340 5095 9408
rect 3873 9306 3991 9340
rect 4025 9306 4059 9340
rect 4093 9306 4127 9340
rect 4161 9306 4195 9340
rect 4229 9306 4263 9340
rect 4297 9306 4331 9340
rect 4365 9306 4399 9340
rect 4433 9306 4467 9340
rect 4501 9306 4535 9340
rect 4569 9306 4603 9340
rect 4637 9306 4671 9340
rect 4705 9306 4739 9340
rect 4773 9306 4807 9340
rect 4841 9306 4875 9340
rect 4909 9306 4943 9340
rect 4977 9306 5095 9340
rect 5340 9475 5406 9483
rect 5340 9441 5356 9475
rect 5390 9441 5406 9475
rect 5340 9407 5406 9441
rect 5340 9373 5356 9407
rect 5390 9373 5406 9407
rect 5340 9339 5406 9373
rect 5340 9305 5356 9339
rect 5390 9305 5406 9339
rect 5340 9287 5406 9305
rect 5440 9475 5482 9517
rect 5474 9441 5482 9475
rect 5440 9407 5482 9441
rect 5474 9373 5482 9407
rect 5440 9339 5482 9373
rect 5474 9305 5482 9339
rect 5440 9289 5482 9305
rect 5340 9237 5386 9287
rect 199 9194 317 9228
rect 351 9194 385 9228
rect 419 9194 453 9228
rect 487 9194 521 9228
rect 555 9194 589 9228
rect 623 9194 657 9228
rect 691 9194 725 9228
rect 759 9194 793 9228
rect 827 9194 861 9228
rect 895 9194 929 9228
rect 963 9194 997 9228
rect 1031 9194 1065 9228
rect 1099 9194 1133 9228
rect 1167 9194 1201 9228
rect 1235 9194 1269 9228
rect 1303 9194 1421 9228
rect 199 9118 233 9194
rect 1387 9123 1421 9194
rect 199 9050 233 9084
rect 199 8982 233 9016
rect 313 9081 347 9120
rect 313 9008 347 9047
rect 409 9081 443 9120
rect 409 9008 443 9047
rect 505 9081 539 9120
rect 505 9008 539 9047
rect 601 9081 635 9120
rect 601 9008 635 9047
rect 697 9081 731 9120
rect 697 9008 731 9047
rect 793 9081 827 9120
rect 793 9008 827 9047
rect 889 9081 923 9120
rect 889 9008 923 9047
rect 985 9081 1019 9120
rect 985 9008 1019 9047
rect 1081 9081 1115 9120
rect 1081 9008 1115 9047
rect 1177 9081 1211 9120
rect 1177 9008 1211 9047
rect 1273 9081 1307 9120
rect 1273 9008 1307 9047
rect 1387 9051 1421 9084
rect 1387 8982 1421 9016
rect 199 8872 233 8948
rect 297 8936 313 8970
rect 347 8936 363 8970
rect 489 8936 505 8970
rect 539 8936 555 8970
rect 681 8936 697 8970
rect 731 8936 747 8970
rect 873 8936 889 8970
rect 923 8936 939 8970
rect 1065 8936 1081 8970
rect 1115 8936 1131 8970
rect 1257 8936 1273 8970
rect 1307 8936 1323 8970
rect 1387 8872 1421 8945
rect 199 8838 317 8872
rect 351 8838 385 8872
rect 419 8838 453 8872
rect 487 8838 521 8872
rect 555 8838 589 8872
rect 623 8838 657 8872
rect 691 8838 725 8872
rect 759 8838 793 8872
rect 827 8838 861 8872
rect 895 8838 929 8872
rect 963 8838 997 8872
rect 1031 8838 1065 8872
rect 1099 8838 1133 8872
rect 1167 8838 1201 8872
rect 1235 8838 1269 8872
rect 1303 8838 1421 8872
rect 2352 9198 2470 9232
rect 2504 9198 2538 9232
rect 2572 9198 2606 9232
rect 2640 9198 2674 9232
rect 2708 9198 2742 9232
rect 2776 9198 2810 9232
rect 2844 9198 2878 9232
rect 2912 9198 2946 9232
rect 2980 9198 3014 9232
rect 3048 9198 3082 9232
rect 3116 9198 3150 9232
rect 3184 9198 3218 9232
rect 3252 9198 3286 9232
rect 3320 9198 3354 9232
rect 3388 9198 3422 9232
rect 3456 9198 3574 9232
rect 2352 9122 2386 9198
rect 3540 9127 3574 9198
rect 3873 9198 3991 9232
rect 4025 9198 4059 9232
rect 4093 9198 4127 9232
rect 4161 9198 4195 9232
rect 4229 9198 4263 9232
rect 4297 9198 4331 9232
rect 4365 9198 4399 9232
rect 4433 9198 4467 9232
rect 4501 9198 4535 9232
rect 4569 9198 4603 9232
rect 4637 9198 4671 9232
rect 4705 9198 4739 9232
rect 4773 9198 4807 9232
rect 4841 9198 4875 9232
rect 4909 9198 4943 9232
rect 4977 9198 5095 9232
rect 3675 9162 3691 9196
rect 3725 9162 3741 9196
rect 2352 9054 2386 9088
rect 2352 8986 2386 9020
rect 2466 9085 2500 9124
rect 2466 9012 2500 9051
rect 2562 9085 2596 9124
rect 2562 9012 2596 9051
rect 2658 9085 2692 9124
rect 2658 9012 2692 9051
rect 2754 9085 2788 9124
rect 2754 9012 2788 9051
rect 2850 9085 2884 9124
rect 2850 9012 2884 9051
rect 2946 9085 2980 9124
rect 2946 9012 2980 9051
rect 3042 9085 3076 9124
rect 3042 9012 3076 9051
rect 3138 9085 3172 9124
rect 3138 9012 3172 9051
rect 3234 9085 3268 9124
rect 3234 9012 3268 9051
rect 3330 9085 3364 9124
rect 3330 9012 3364 9051
rect 3426 9085 3460 9124
rect 3426 9012 3460 9051
rect 3540 9055 3574 9088
rect 3647 9112 3681 9128
rect 3647 9020 3681 9036
rect 3735 9112 3769 9128
rect 3735 9020 3769 9036
rect 3873 9122 3907 9198
rect 5061 9127 5095 9198
rect 3873 9054 3907 9088
rect 3540 8986 3574 9020
rect 2352 8876 2386 8952
rect 2450 8940 2466 8974
rect 2500 8940 2516 8974
rect 2642 8940 2658 8974
rect 2692 8940 2708 8974
rect 2834 8940 2850 8974
rect 2884 8940 2900 8974
rect 3026 8940 3042 8974
rect 3076 8940 3092 8974
rect 3218 8940 3234 8974
rect 3268 8940 3284 8974
rect 3410 8940 3426 8974
rect 3460 8940 3476 8974
rect 3540 8876 3574 8949
rect 2352 8842 2470 8876
rect 2504 8842 2538 8876
rect 2572 8842 2606 8876
rect 2640 8842 2674 8876
rect 2708 8842 2742 8876
rect 2776 8842 2810 8876
rect 2844 8842 2878 8876
rect 2912 8842 2946 8876
rect 2980 8842 3014 8876
rect 3048 8842 3082 8876
rect 3116 8842 3150 8876
rect 3184 8842 3218 8876
rect 3252 8842 3286 8876
rect 3320 8842 3354 8876
rect 3388 8842 3422 8876
rect 3456 8842 3574 8876
rect 3873 8986 3907 9020
rect 3987 9085 4021 9124
rect 3987 9012 4021 9051
rect 4083 9085 4117 9124
rect 4083 9012 4117 9051
rect 4179 9085 4213 9124
rect 4179 9012 4213 9051
rect 4275 9085 4309 9124
rect 4275 9012 4309 9051
rect 4371 9085 4405 9124
rect 4371 9012 4405 9051
rect 4467 9085 4501 9124
rect 4467 9012 4501 9051
rect 4563 9085 4597 9124
rect 4563 9012 4597 9051
rect 4659 9085 4693 9124
rect 4659 9012 4693 9051
rect 4755 9085 4789 9124
rect 4755 9012 4789 9051
rect 4851 9085 4885 9124
rect 4851 9012 4885 9051
rect 4947 9085 4981 9124
rect 4947 9012 4981 9051
rect 5061 9055 5095 9088
rect 5340 9203 5348 9237
rect 5382 9203 5386 9237
rect 5420 9242 5486 9253
rect 5420 9239 5450 9242
rect 5420 9205 5436 9239
rect 5484 9208 5486 9242
rect 5470 9205 5486 9208
rect 5340 9167 5386 9203
rect 5340 9155 5406 9167
rect 5340 9121 5356 9155
rect 5390 9121 5406 9155
rect 5340 9087 5406 9121
rect 5340 9053 5356 9087
rect 5390 9053 5406 9087
rect 5340 9041 5406 9053
rect 5440 9155 5486 9171
rect 5474 9121 5486 9155
rect 5440 9087 5486 9121
rect 5474 9053 5486 9087
rect 5061 8986 5095 9020
rect 5440 9007 5486 9053
rect 3873 8876 3907 8952
rect 3971 8940 3987 8974
rect 4021 8940 4037 8974
rect 4163 8940 4179 8974
rect 4213 8940 4229 8974
rect 4355 8940 4371 8974
rect 4405 8940 4421 8974
rect 4547 8940 4563 8974
rect 4597 8940 4613 8974
rect 4739 8940 4755 8974
rect 4789 8940 4805 8974
rect 4931 8940 4947 8974
rect 4981 8940 4997 8974
rect 5274 8973 5303 9007
rect 5337 8973 5395 9007
rect 5429 8973 5487 9007
rect 5521 8973 5550 9007
rect 5061 8876 5095 8949
rect 3873 8842 3991 8876
rect 4025 8842 4059 8876
rect 4093 8842 4127 8876
rect 4161 8842 4195 8876
rect 4229 8842 4263 8876
rect 4297 8842 4331 8876
rect 4365 8842 4399 8876
rect 4433 8842 4467 8876
rect 4501 8842 4535 8876
rect 4569 8842 4603 8876
rect 4637 8842 4671 8876
rect 4705 8842 4739 8876
rect 4773 8842 4807 8876
rect 4841 8842 4875 8876
rect 4909 8842 4943 8876
rect 4977 8842 5095 8876
rect 199 8559 317 8593
rect 351 8559 385 8593
rect 419 8559 453 8593
rect 487 8559 521 8593
rect 555 8559 589 8593
rect 623 8559 657 8593
rect 691 8559 725 8593
rect 759 8559 793 8593
rect 827 8559 861 8593
rect 895 8559 929 8593
rect 963 8559 997 8593
rect 1031 8559 1065 8593
rect 1099 8559 1133 8593
rect 1167 8559 1201 8593
rect 1235 8559 1269 8593
rect 1303 8559 1421 8593
rect 199 8491 233 8559
rect 1387 8491 1421 8559
rect 297 8457 313 8491
rect 347 8457 363 8491
rect 489 8457 505 8491
rect 539 8457 555 8491
rect 681 8457 697 8491
rect 731 8457 747 8491
rect 873 8457 889 8491
rect 923 8457 939 8491
rect 1065 8457 1081 8491
rect 1115 8457 1131 8491
rect 1257 8457 1273 8491
rect 1307 8457 1323 8491
rect 199 8423 233 8457
rect 1387 8423 1421 8431
rect 199 8355 233 8389
rect 199 8287 233 8321
rect 199 8219 233 8253
rect 199 8151 233 8185
rect 313 8392 347 8413
rect 313 8324 347 8328
rect 313 8218 347 8222
rect 313 8133 347 8154
rect 409 8392 443 8413
rect 409 8324 443 8328
rect 409 8218 443 8222
rect 409 8133 443 8154
rect 505 8392 539 8413
rect 505 8324 539 8328
rect 505 8218 539 8222
rect 505 8133 539 8154
rect 601 8392 635 8413
rect 601 8324 635 8328
rect 601 8218 635 8222
rect 601 8133 635 8154
rect 697 8392 731 8413
rect 697 8324 731 8328
rect 697 8218 731 8222
rect 697 8133 731 8154
rect 793 8392 827 8413
rect 793 8324 827 8328
rect 793 8218 827 8222
rect 793 8133 827 8154
rect 889 8392 923 8413
rect 889 8324 923 8328
rect 889 8218 923 8222
rect 889 8133 923 8154
rect 985 8392 1019 8413
rect 985 8324 1019 8328
rect 985 8218 1019 8222
rect 985 8133 1019 8154
rect 1081 8392 1115 8413
rect 1081 8324 1115 8328
rect 1081 8218 1115 8222
rect 1081 8133 1115 8154
rect 1177 8392 1211 8413
rect 1177 8324 1211 8328
rect 1177 8218 1211 8222
rect 1177 8133 1211 8154
rect 1273 8392 1307 8413
rect 1273 8324 1307 8328
rect 1273 8218 1307 8222
rect 1273 8133 1307 8154
rect 1387 8355 1421 8359
rect 1387 8249 1421 8253
rect 1387 8177 1421 8185
rect 199 8049 233 8117
rect 1387 8049 1421 8117
rect 199 8015 317 8049
rect 351 8015 385 8049
rect 419 8015 453 8049
rect 487 8015 521 8049
rect 555 8015 589 8049
rect 623 8015 657 8049
rect 691 8015 725 8049
rect 759 8015 793 8049
rect 827 8015 861 8049
rect 895 8015 929 8049
rect 963 8015 997 8049
rect 1031 8015 1065 8049
rect 1099 8015 1133 8049
rect 1167 8015 1201 8049
rect 1235 8015 1269 8049
rect 1303 8015 1421 8049
rect 2352 8563 2470 8597
rect 2504 8563 2538 8597
rect 2572 8563 2606 8597
rect 2640 8563 2674 8597
rect 2708 8563 2742 8597
rect 2776 8563 2810 8597
rect 2844 8563 2878 8597
rect 2912 8563 2946 8597
rect 2980 8563 3014 8597
rect 3048 8563 3082 8597
rect 3116 8563 3150 8597
rect 3184 8563 3218 8597
rect 3252 8563 3286 8597
rect 3320 8563 3354 8597
rect 3388 8563 3422 8597
rect 3456 8563 3574 8597
rect 2352 8495 2386 8563
rect 3540 8495 3574 8563
rect 2450 8461 2466 8495
rect 2500 8461 2516 8495
rect 2642 8461 2658 8495
rect 2692 8461 2708 8495
rect 2834 8461 2850 8495
rect 2884 8461 2900 8495
rect 3026 8461 3042 8495
rect 3076 8461 3092 8495
rect 3218 8461 3234 8495
rect 3268 8461 3284 8495
rect 3410 8461 3426 8495
rect 3460 8461 3476 8495
rect 2352 8427 2386 8461
rect 3540 8427 3574 8435
rect 2352 8359 2386 8393
rect 2352 8291 2386 8325
rect 2352 8223 2386 8257
rect 2352 8155 2386 8189
rect 2466 8396 2500 8417
rect 2466 8328 2500 8332
rect 2466 8222 2500 8226
rect 2466 8137 2500 8158
rect 2562 8396 2596 8417
rect 2562 8328 2596 8332
rect 2562 8222 2596 8226
rect 2562 8137 2596 8158
rect 2658 8396 2692 8417
rect 2658 8328 2692 8332
rect 2658 8222 2692 8226
rect 2658 8137 2692 8158
rect 2754 8396 2788 8417
rect 2754 8328 2788 8332
rect 2754 8222 2788 8226
rect 2754 8137 2788 8158
rect 2850 8396 2884 8417
rect 2850 8328 2884 8332
rect 2850 8222 2884 8226
rect 2850 8137 2884 8158
rect 2946 8396 2980 8417
rect 2946 8328 2980 8332
rect 2946 8222 2980 8226
rect 2946 8137 2980 8158
rect 3042 8396 3076 8417
rect 3042 8328 3076 8332
rect 3042 8222 3076 8226
rect 3042 8137 3076 8158
rect 3138 8396 3172 8417
rect 3138 8328 3172 8332
rect 3138 8222 3172 8226
rect 3138 8137 3172 8158
rect 3234 8396 3268 8417
rect 3234 8328 3268 8332
rect 3234 8222 3268 8226
rect 3234 8137 3268 8158
rect 3330 8396 3364 8417
rect 3330 8328 3364 8332
rect 3330 8222 3364 8226
rect 3330 8137 3364 8158
rect 3426 8396 3460 8417
rect 3426 8328 3460 8332
rect 3426 8222 3460 8226
rect 3426 8137 3460 8158
rect 3540 8359 3574 8363
rect 3540 8253 3574 8257
rect 3540 8181 3574 8189
rect 2352 8053 2386 8121
rect 3540 8053 3574 8121
rect 2352 8019 2470 8053
rect 2504 8019 2538 8053
rect 2572 8019 2606 8053
rect 2640 8019 2674 8053
rect 2708 8019 2742 8053
rect 2776 8019 2810 8053
rect 2844 8019 2878 8053
rect 2912 8019 2946 8053
rect 2980 8019 3014 8053
rect 3048 8019 3082 8053
rect 3116 8019 3150 8053
rect 3184 8019 3218 8053
rect 3252 8019 3286 8053
rect 3320 8019 3354 8053
rect 3388 8019 3422 8053
rect 3456 8019 3574 8053
rect 3873 8563 3991 8597
rect 4025 8563 4059 8597
rect 4093 8563 4127 8597
rect 4161 8563 4195 8597
rect 4229 8563 4263 8597
rect 4297 8563 4331 8597
rect 4365 8563 4399 8597
rect 4433 8563 4467 8597
rect 4501 8563 4535 8597
rect 4569 8563 4603 8597
rect 4637 8563 4671 8597
rect 4705 8563 4739 8597
rect 4773 8563 4807 8597
rect 4841 8563 4875 8597
rect 4909 8563 4943 8597
rect 4977 8563 5095 8597
rect 3873 8495 3907 8563
rect 5061 8495 5095 8563
rect 3971 8461 3987 8495
rect 4021 8461 4037 8495
rect 4163 8461 4179 8495
rect 4213 8461 4229 8495
rect 4355 8461 4371 8495
rect 4405 8461 4421 8495
rect 4547 8461 4563 8495
rect 4597 8461 4613 8495
rect 4739 8461 4755 8495
rect 4789 8461 4805 8495
rect 4931 8461 4947 8495
rect 4981 8461 4997 8495
rect 3873 8427 3907 8461
rect 5061 8427 5095 8435
rect 3873 8359 3907 8393
rect 3873 8291 3907 8325
rect 3873 8223 3907 8257
rect 3873 8155 3907 8189
rect 3987 8396 4021 8417
rect 3987 8328 4021 8332
rect 3987 8222 4021 8226
rect 3987 8137 4021 8158
rect 4083 8396 4117 8417
rect 4083 8328 4117 8332
rect 4083 8222 4117 8226
rect 4083 8137 4117 8158
rect 4179 8396 4213 8417
rect 4179 8328 4213 8332
rect 4179 8222 4213 8226
rect 4179 8137 4213 8158
rect 4275 8396 4309 8417
rect 4275 8328 4309 8332
rect 4275 8222 4309 8226
rect 4275 8137 4309 8158
rect 4371 8396 4405 8417
rect 4371 8328 4405 8332
rect 4371 8222 4405 8226
rect 4371 8137 4405 8158
rect 4467 8396 4501 8417
rect 4467 8328 4501 8332
rect 4467 8222 4501 8226
rect 4467 8137 4501 8158
rect 4563 8396 4597 8417
rect 4563 8328 4597 8332
rect 4563 8222 4597 8226
rect 4563 8137 4597 8158
rect 4659 8396 4693 8417
rect 4659 8328 4693 8332
rect 4659 8222 4693 8226
rect 4659 8137 4693 8158
rect 4755 8396 4789 8417
rect 4755 8328 4789 8332
rect 4755 8222 4789 8226
rect 4755 8137 4789 8158
rect 4851 8396 4885 8417
rect 4851 8328 4885 8332
rect 4851 8222 4885 8226
rect 4851 8137 4885 8158
rect 4947 8396 4981 8417
rect 4947 8328 4981 8332
rect 4947 8222 4981 8226
rect 4947 8137 4981 8158
rect 5061 8359 5095 8363
rect 5061 8253 5095 8257
rect 5274 8230 5303 8264
rect 5337 8230 5395 8264
rect 5429 8230 5487 8264
rect 5521 8230 5550 8264
rect 5061 8181 5095 8189
rect 3873 8053 3907 8121
rect 5061 8053 5095 8121
rect 3873 8019 3991 8053
rect 4025 8019 4059 8053
rect 4093 8019 4127 8053
rect 4161 8019 4195 8053
rect 4229 8019 4263 8053
rect 4297 8019 4331 8053
rect 4365 8019 4399 8053
rect 4433 8019 4467 8053
rect 4501 8019 4535 8053
rect 4569 8019 4603 8053
rect 4637 8019 4671 8053
rect 4705 8019 4739 8053
rect 4773 8019 4807 8053
rect 4841 8019 4875 8053
rect 4909 8019 4943 8053
rect 4977 8019 5095 8053
rect 5340 8188 5406 8196
rect 5340 8154 5356 8188
rect 5390 8154 5406 8188
rect 5340 8120 5406 8154
rect 5340 8086 5356 8120
rect 5390 8086 5406 8120
rect 5340 8052 5406 8086
rect 5340 8018 5356 8052
rect 5390 8018 5406 8052
rect 5340 8000 5406 8018
rect 5440 8188 5482 8230
rect 5474 8154 5482 8188
rect 5440 8120 5482 8154
rect 5474 8086 5482 8120
rect 5440 8052 5482 8086
rect 5474 8018 5482 8052
rect 5440 8002 5482 8018
rect 5340 7950 5386 8000
rect 199 7907 317 7941
rect 351 7907 385 7941
rect 419 7907 453 7941
rect 487 7907 521 7941
rect 555 7907 589 7941
rect 623 7907 657 7941
rect 691 7907 725 7941
rect 759 7907 793 7941
rect 827 7907 861 7941
rect 895 7907 929 7941
rect 963 7907 997 7941
rect 1031 7907 1065 7941
rect 1099 7907 1133 7941
rect 1167 7907 1201 7941
rect 1235 7907 1269 7941
rect 1303 7907 1421 7941
rect 199 7831 233 7907
rect 1387 7836 1421 7907
rect 199 7763 233 7797
rect 199 7695 233 7729
rect 313 7794 347 7833
rect 313 7721 347 7760
rect 409 7794 443 7833
rect 409 7721 443 7760
rect 505 7794 539 7833
rect 505 7721 539 7760
rect 601 7794 635 7833
rect 601 7721 635 7760
rect 697 7794 731 7833
rect 697 7721 731 7760
rect 793 7794 827 7833
rect 793 7721 827 7760
rect 889 7794 923 7833
rect 889 7721 923 7760
rect 985 7794 1019 7833
rect 985 7721 1019 7760
rect 1081 7794 1115 7833
rect 1081 7721 1115 7760
rect 1177 7794 1211 7833
rect 1177 7721 1211 7760
rect 1273 7794 1307 7833
rect 1273 7721 1307 7760
rect 1387 7764 1421 7797
rect 1387 7695 1421 7729
rect 199 7585 233 7661
rect 297 7649 313 7683
rect 347 7649 363 7683
rect 489 7649 505 7683
rect 539 7649 555 7683
rect 681 7649 697 7683
rect 731 7649 747 7683
rect 873 7649 889 7683
rect 923 7649 939 7683
rect 1065 7649 1081 7683
rect 1115 7649 1131 7683
rect 1257 7649 1273 7683
rect 1307 7649 1323 7683
rect 1387 7585 1421 7658
rect 199 7551 317 7585
rect 351 7551 385 7585
rect 419 7551 453 7585
rect 487 7551 521 7585
rect 555 7551 589 7585
rect 623 7551 657 7585
rect 691 7551 725 7585
rect 759 7551 793 7585
rect 827 7551 861 7585
rect 895 7551 929 7585
rect 963 7551 997 7585
rect 1031 7551 1065 7585
rect 1099 7551 1133 7585
rect 1167 7551 1201 7585
rect 1235 7551 1269 7585
rect 1303 7551 1421 7585
rect 2352 7911 2470 7945
rect 2504 7911 2538 7945
rect 2572 7911 2606 7945
rect 2640 7911 2674 7945
rect 2708 7911 2742 7945
rect 2776 7911 2810 7945
rect 2844 7911 2878 7945
rect 2912 7911 2946 7945
rect 2980 7911 3014 7945
rect 3048 7911 3082 7945
rect 3116 7911 3150 7945
rect 3184 7911 3218 7945
rect 3252 7911 3286 7945
rect 3320 7911 3354 7945
rect 3388 7911 3422 7945
rect 3456 7911 3574 7945
rect 2352 7835 2386 7911
rect 3540 7840 3574 7911
rect 3873 7911 3991 7945
rect 4025 7911 4059 7945
rect 4093 7911 4127 7945
rect 4161 7911 4195 7945
rect 4229 7911 4263 7945
rect 4297 7911 4331 7945
rect 4365 7911 4399 7945
rect 4433 7911 4467 7945
rect 4501 7911 4535 7945
rect 4569 7911 4603 7945
rect 4637 7911 4671 7945
rect 4705 7911 4739 7945
rect 4773 7911 4807 7945
rect 4841 7911 4875 7945
rect 4909 7911 4943 7945
rect 4977 7911 5095 7945
rect 3675 7875 3691 7909
rect 3725 7875 3741 7909
rect 2352 7767 2386 7801
rect 2352 7699 2386 7733
rect 2466 7798 2500 7837
rect 2466 7725 2500 7764
rect 2562 7798 2596 7837
rect 2562 7725 2596 7764
rect 2658 7798 2692 7837
rect 2658 7725 2692 7764
rect 2754 7798 2788 7837
rect 2754 7725 2788 7764
rect 2850 7798 2884 7837
rect 2850 7725 2884 7764
rect 2946 7798 2980 7837
rect 2946 7725 2980 7764
rect 3042 7798 3076 7837
rect 3042 7725 3076 7764
rect 3138 7798 3172 7837
rect 3138 7725 3172 7764
rect 3234 7798 3268 7837
rect 3234 7725 3268 7764
rect 3330 7798 3364 7837
rect 3330 7725 3364 7764
rect 3426 7798 3460 7837
rect 3426 7725 3460 7764
rect 3540 7768 3574 7801
rect 3647 7825 3681 7841
rect 3647 7733 3681 7749
rect 3735 7825 3769 7841
rect 3735 7733 3769 7749
rect 3873 7835 3907 7911
rect 5061 7840 5095 7911
rect 3873 7767 3907 7801
rect 3540 7699 3574 7733
rect 2352 7589 2386 7665
rect 2450 7653 2466 7687
rect 2500 7653 2516 7687
rect 2642 7653 2658 7687
rect 2692 7653 2708 7687
rect 2834 7653 2850 7687
rect 2884 7653 2900 7687
rect 3026 7653 3042 7687
rect 3076 7653 3092 7687
rect 3218 7653 3234 7687
rect 3268 7653 3284 7687
rect 3410 7653 3426 7687
rect 3460 7653 3476 7687
rect 3540 7589 3574 7662
rect 2352 7555 2470 7589
rect 2504 7555 2538 7589
rect 2572 7555 2606 7589
rect 2640 7555 2674 7589
rect 2708 7555 2742 7589
rect 2776 7555 2810 7589
rect 2844 7555 2878 7589
rect 2912 7555 2946 7589
rect 2980 7555 3014 7589
rect 3048 7555 3082 7589
rect 3116 7555 3150 7589
rect 3184 7555 3218 7589
rect 3252 7555 3286 7589
rect 3320 7555 3354 7589
rect 3388 7555 3422 7589
rect 3456 7555 3574 7589
rect 3873 7699 3907 7733
rect 3987 7798 4021 7837
rect 3987 7725 4021 7764
rect 4083 7798 4117 7837
rect 4083 7725 4117 7764
rect 4179 7798 4213 7837
rect 4179 7725 4213 7764
rect 4275 7798 4309 7837
rect 4275 7725 4309 7764
rect 4371 7798 4405 7837
rect 4371 7725 4405 7764
rect 4467 7798 4501 7837
rect 4467 7725 4501 7764
rect 4563 7798 4597 7837
rect 4563 7725 4597 7764
rect 4659 7798 4693 7837
rect 4659 7725 4693 7764
rect 4755 7798 4789 7837
rect 4755 7725 4789 7764
rect 4851 7798 4885 7837
rect 4851 7725 4885 7764
rect 4947 7798 4981 7837
rect 4947 7725 4981 7764
rect 5061 7768 5095 7801
rect 5340 7916 5348 7950
rect 5382 7916 5386 7950
rect 5420 7955 5486 7966
rect 5420 7952 5450 7955
rect 5420 7918 5436 7952
rect 5484 7921 5486 7955
rect 5470 7918 5486 7921
rect 5340 7880 5386 7916
rect 5340 7868 5406 7880
rect 5340 7834 5356 7868
rect 5390 7834 5406 7868
rect 5340 7800 5406 7834
rect 5340 7766 5356 7800
rect 5390 7766 5406 7800
rect 5340 7754 5406 7766
rect 5440 7868 5486 7884
rect 5474 7834 5486 7868
rect 5440 7800 5486 7834
rect 5474 7766 5486 7800
rect 5061 7699 5095 7733
rect 5440 7720 5486 7766
rect 3873 7589 3907 7665
rect 3971 7653 3987 7687
rect 4021 7653 4037 7687
rect 4163 7653 4179 7687
rect 4213 7653 4229 7687
rect 4355 7653 4371 7687
rect 4405 7653 4421 7687
rect 4547 7653 4563 7687
rect 4597 7653 4613 7687
rect 4739 7653 4755 7687
rect 4789 7653 4805 7687
rect 4931 7653 4947 7687
rect 4981 7653 4997 7687
rect 5274 7686 5303 7720
rect 5337 7686 5395 7720
rect 5429 7686 5487 7720
rect 5521 7686 5550 7720
rect 5061 7589 5095 7662
rect 3873 7555 3991 7589
rect 4025 7555 4059 7589
rect 4093 7555 4127 7589
rect 4161 7555 4195 7589
rect 4229 7555 4263 7589
rect 4297 7555 4331 7589
rect 4365 7555 4399 7589
rect 4433 7555 4467 7589
rect 4501 7555 4535 7589
rect 4569 7555 4603 7589
rect 4637 7555 4671 7589
rect 4705 7555 4739 7589
rect 4773 7555 4807 7589
rect 4841 7555 4875 7589
rect 4909 7555 4943 7589
rect 4977 7555 5095 7589
rect 199 7272 317 7306
rect 351 7272 385 7306
rect 419 7272 453 7306
rect 487 7272 521 7306
rect 555 7272 589 7306
rect 623 7272 657 7306
rect 691 7272 725 7306
rect 759 7272 793 7306
rect 827 7272 861 7306
rect 895 7272 929 7306
rect 963 7272 997 7306
rect 1031 7272 1065 7306
rect 1099 7272 1133 7306
rect 1167 7272 1201 7306
rect 1235 7272 1269 7306
rect 1303 7272 1421 7306
rect 199 7204 233 7272
rect 1387 7204 1421 7272
rect 297 7170 313 7204
rect 347 7170 363 7204
rect 489 7170 505 7204
rect 539 7170 555 7204
rect 681 7170 697 7204
rect 731 7170 747 7204
rect 873 7170 889 7204
rect 923 7170 939 7204
rect 1065 7170 1081 7204
rect 1115 7170 1131 7204
rect 1257 7170 1273 7204
rect 1307 7170 1323 7204
rect 199 7136 233 7170
rect 1387 7136 1421 7144
rect 199 7068 233 7102
rect 199 7000 233 7034
rect 199 6932 233 6966
rect 199 6864 233 6898
rect 313 7105 347 7126
rect 313 7037 347 7041
rect 313 6931 347 6935
rect 313 6846 347 6867
rect 409 7105 443 7126
rect 409 7037 443 7041
rect 409 6931 443 6935
rect 409 6846 443 6867
rect 505 7105 539 7126
rect 505 7037 539 7041
rect 505 6931 539 6935
rect 505 6846 539 6867
rect 601 7105 635 7126
rect 601 7037 635 7041
rect 601 6931 635 6935
rect 601 6846 635 6867
rect 697 7105 731 7126
rect 697 7037 731 7041
rect 697 6931 731 6935
rect 697 6846 731 6867
rect 793 7105 827 7126
rect 793 7037 827 7041
rect 793 6931 827 6935
rect 793 6846 827 6867
rect 889 7105 923 7126
rect 889 7037 923 7041
rect 889 6931 923 6935
rect 889 6846 923 6867
rect 985 7105 1019 7126
rect 985 7037 1019 7041
rect 985 6931 1019 6935
rect 985 6846 1019 6867
rect 1081 7105 1115 7126
rect 1081 7037 1115 7041
rect 1081 6931 1115 6935
rect 1081 6846 1115 6867
rect 1177 7105 1211 7126
rect 1177 7037 1211 7041
rect 1177 6931 1211 6935
rect 1177 6846 1211 6867
rect 1273 7105 1307 7126
rect 1273 7037 1307 7041
rect 1273 6931 1307 6935
rect 1273 6846 1307 6867
rect 1387 7068 1421 7072
rect 1387 6962 1421 6966
rect 1387 6890 1421 6898
rect 199 6762 233 6830
rect 1387 6762 1421 6830
rect 199 6728 317 6762
rect 351 6728 385 6762
rect 419 6728 453 6762
rect 487 6728 521 6762
rect 555 6728 589 6762
rect 623 6728 657 6762
rect 691 6728 725 6762
rect 759 6728 793 6762
rect 827 6728 861 6762
rect 895 6728 929 6762
rect 963 6728 997 6762
rect 1031 6728 1065 6762
rect 1099 6728 1133 6762
rect 1167 6728 1201 6762
rect 1235 6728 1269 6762
rect 1303 6728 1421 6762
rect 2352 7276 2470 7310
rect 2504 7276 2538 7310
rect 2572 7276 2606 7310
rect 2640 7276 2674 7310
rect 2708 7276 2742 7310
rect 2776 7276 2810 7310
rect 2844 7276 2878 7310
rect 2912 7276 2946 7310
rect 2980 7276 3014 7310
rect 3048 7276 3082 7310
rect 3116 7276 3150 7310
rect 3184 7276 3218 7310
rect 3252 7276 3286 7310
rect 3320 7276 3354 7310
rect 3388 7276 3422 7310
rect 3456 7276 3574 7310
rect 2352 7208 2386 7276
rect 3540 7208 3574 7276
rect 2450 7174 2466 7208
rect 2500 7174 2516 7208
rect 2642 7174 2658 7208
rect 2692 7174 2708 7208
rect 2834 7174 2850 7208
rect 2884 7174 2900 7208
rect 3026 7174 3042 7208
rect 3076 7174 3092 7208
rect 3218 7174 3234 7208
rect 3268 7174 3284 7208
rect 3410 7174 3426 7208
rect 3460 7174 3476 7208
rect 2352 7140 2386 7174
rect 3540 7140 3574 7148
rect 2352 7072 2386 7106
rect 2352 7004 2386 7038
rect 2352 6936 2386 6970
rect 2352 6868 2386 6902
rect 2466 7109 2500 7130
rect 2466 7041 2500 7045
rect 2466 6935 2500 6939
rect 2466 6850 2500 6871
rect 2562 7109 2596 7130
rect 2562 7041 2596 7045
rect 2562 6935 2596 6939
rect 2562 6850 2596 6871
rect 2658 7109 2692 7130
rect 2658 7041 2692 7045
rect 2658 6935 2692 6939
rect 2658 6850 2692 6871
rect 2754 7109 2788 7130
rect 2754 7041 2788 7045
rect 2754 6935 2788 6939
rect 2754 6850 2788 6871
rect 2850 7109 2884 7130
rect 2850 7041 2884 7045
rect 2850 6935 2884 6939
rect 2850 6850 2884 6871
rect 2946 7109 2980 7130
rect 2946 7041 2980 7045
rect 2946 6935 2980 6939
rect 2946 6850 2980 6871
rect 3042 7109 3076 7130
rect 3042 7041 3076 7045
rect 3042 6935 3076 6939
rect 3042 6850 3076 6871
rect 3138 7109 3172 7130
rect 3138 7041 3172 7045
rect 3138 6935 3172 6939
rect 3138 6850 3172 6871
rect 3234 7109 3268 7130
rect 3234 7041 3268 7045
rect 3234 6935 3268 6939
rect 3234 6850 3268 6871
rect 3330 7109 3364 7130
rect 3330 7041 3364 7045
rect 3330 6935 3364 6939
rect 3330 6850 3364 6871
rect 3426 7109 3460 7130
rect 3426 7041 3460 7045
rect 3426 6935 3460 6939
rect 3426 6850 3460 6871
rect 3540 7072 3574 7076
rect 3540 6966 3574 6970
rect 3540 6894 3574 6902
rect 2352 6766 2386 6834
rect 3540 6766 3574 6834
rect 2352 6732 2470 6766
rect 2504 6732 2538 6766
rect 2572 6732 2606 6766
rect 2640 6732 2674 6766
rect 2708 6732 2742 6766
rect 2776 6732 2810 6766
rect 2844 6732 2878 6766
rect 2912 6732 2946 6766
rect 2980 6732 3014 6766
rect 3048 6732 3082 6766
rect 3116 6732 3150 6766
rect 3184 6732 3218 6766
rect 3252 6732 3286 6766
rect 3320 6732 3354 6766
rect 3388 6732 3422 6766
rect 3456 6732 3574 6766
rect 3873 7276 3991 7310
rect 4025 7276 4059 7310
rect 4093 7276 4127 7310
rect 4161 7276 4195 7310
rect 4229 7276 4263 7310
rect 4297 7276 4331 7310
rect 4365 7276 4399 7310
rect 4433 7276 4467 7310
rect 4501 7276 4535 7310
rect 4569 7276 4603 7310
rect 4637 7276 4671 7310
rect 4705 7276 4739 7310
rect 4773 7276 4807 7310
rect 4841 7276 4875 7310
rect 4909 7276 4943 7310
rect 4977 7276 5095 7310
rect 3873 7208 3907 7276
rect 5061 7208 5095 7276
rect 3971 7174 3987 7208
rect 4021 7174 4037 7208
rect 4163 7174 4179 7208
rect 4213 7174 4229 7208
rect 4355 7174 4371 7208
rect 4405 7174 4421 7208
rect 4547 7174 4563 7208
rect 4597 7174 4613 7208
rect 4739 7174 4755 7208
rect 4789 7174 4805 7208
rect 4931 7174 4947 7208
rect 4981 7174 4997 7208
rect 3873 7140 3907 7174
rect 5061 7140 5095 7148
rect 3873 7072 3907 7106
rect 3873 7004 3907 7038
rect 3873 6936 3907 6970
rect 3873 6868 3907 6902
rect 3987 7109 4021 7130
rect 3987 7041 4021 7045
rect 3987 6935 4021 6939
rect 3987 6850 4021 6871
rect 4083 7109 4117 7130
rect 4083 7041 4117 7045
rect 4083 6935 4117 6939
rect 4083 6850 4117 6871
rect 4179 7109 4213 7130
rect 4179 7041 4213 7045
rect 4179 6935 4213 6939
rect 4179 6850 4213 6871
rect 4275 7109 4309 7130
rect 4275 7041 4309 7045
rect 4275 6935 4309 6939
rect 4275 6850 4309 6871
rect 4371 7109 4405 7130
rect 4371 7041 4405 7045
rect 4371 6935 4405 6939
rect 4371 6850 4405 6871
rect 4467 7109 4501 7130
rect 4467 7041 4501 7045
rect 4467 6935 4501 6939
rect 4467 6850 4501 6871
rect 4563 7109 4597 7130
rect 4563 7041 4597 7045
rect 4563 6935 4597 6939
rect 4563 6850 4597 6871
rect 4659 7109 4693 7130
rect 4659 7041 4693 7045
rect 4659 6935 4693 6939
rect 4659 6850 4693 6871
rect 4755 7109 4789 7130
rect 4755 7041 4789 7045
rect 4755 6935 4789 6939
rect 4755 6850 4789 6871
rect 4851 7109 4885 7130
rect 4851 7041 4885 7045
rect 4851 6935 4885 6939
rect 4851 6850 4885 6871
rect 4947 7109 4981 7130
rect 4947 7041 4981 7045
rect 4947 6935 4981 6939
rect 4947 6850 4981 6871
rect 5061 7072 5095 7076
rect 5061 6966 5095 6970
rect 5274 6943 5303 6977
rect 5337 6943 5395 6977
rect 5429 6943 5487 6977
rect 5521 6943 5550 6977
rect 5061 6894 5095 6902
rect 3873 6766 3907 6834
rect 5061 6766 5095 6834
rect 3873 6732 3991 6766
rect 4025 6732 4059 6766
rect 4093 6732 4127 6766
rect 4161 6732 4195 6766
rect 4229 6732 4263 6766
rect 4297 6732 4331 6766
rect 4365 6732 4399 6766
rect 4433 6732 4467 6766
rect 4501 6732 4535 6766
rect 4569 6732 4603 6766
rect 4637 6732 4671 6766
rect 4705 6732 4739 6766
rect 4773 6732 4807 6766
rect 4841 6732 4875 6766
rect 4909 6732 4943 6766
rect 4977 6732 5095 6766
rect 5340 6901 5406 6909
rect 5340 6867 5356 6901
rect 5390 6867 5406 6901
rect 5340 6833 5406 6867
rect 5340 6799 5356 6833
rect 5390 6799 5406 6833
rect 5340 6765 5406 6799
rect 5340 6731 5356 6765
rect 5390 6731 5406 6765
rect 5340 6713 5406 6731
rect 5440 6901 5482 6943
rect 5474 6867 5482 6901
rect 5440 6833 5482 6867
rect 5474 6799 5482 6833
rect 5440 6765 5482 6799
rect 5474 6731 5482 6765
rect 5440 6715 5482 6731
rect 5340 6663 5386 6713
rect 199 6620 317 6654
rect 351 6620 385 6654
rect 419 6620 453 6654
rect 487 6620 521 6654
rect 555 6620 589 6654
rect 623 6620 657 6654
rect 691 6620 725 6654
rect 759 6620 793 6654
rect 827 6620 861 6654
rect 895 6620 929 6654
rect 963 6620 997 6654
rect 1031 6620 1065 6654
rect 1099 6620 1133 6654
rect 1167 6620 1201 6654
rect 1235 6620 1269 6654
rect 1303 6620 1421 6654
rect 199 6544 233 6620
rect 1387 6549 1421 6620
rect 199 6476 233 6510
rect 199 6408 233 6442
rect 313 6507 347 6546
rect 313 6434 347 6473
rect 409 6507 443 6546
rect 409 6434 443 6473
rect 505 6507 539 6546
rect 505 6434 539 6473
rect 601 6507 635 6546
rect 601 6434 635 6473
rect 697 6507 731 6546
rect 697 6434 731 6473
rect 793 6507 827 6546
rect 793 6434 827 6473
rect 889 6507 923 6546
rect 889 6434 923 6473
rect 985 6507 1019 6546
rect 985 6434 1019 6473
rect 1081 6507 1115 6546
rect 1081 6434 1115 6473
rect 1177 6507 1211 6546
rect 1177 6434 1211 6473
rect 1273 6507 1307 6546
rect 1273 6434 1307 6473
rect 1387 6477 1421 6510
rect 1387 6408 1421 6442
rect 199 6298 233 6374
rect 297 6362 313 6396
rect 347 6362 363 6396
rect 489 6362 505 6396
rect 539 6362 555 6396
rect 681 6362 697 6396
rect 731 6362 747 6396
rect 873 6362 889 6396
rect 923 6362 939 6396
rect 1065 6362 1081 6396
rect 1115 6362 1131 6396
rect 1257 6362 1273 6396
rect 1307 6362 1323 6396
rect 1387 6298 1421 6371
rect 199 6264 317 6298
rect 351 6264 385 6298
rect 419 6264 453 6298
rect 487 6264 521 6298
rect 555 6264 589 6298
rect 623 6264 657 6298
rect 691 6264 725 6298
rect 759 6264 793 6298
rect 827 6264 861 6298
rect 895 6264 929 6298
rect 963 6264 997 6298
rect 1031 6264 1065 6298
rect 1099 6264 1133 6298
rect 1167 6264 1201 6298
rect 1235 6264 1269 6298
rect 1303 6264 1421 6298
rect 2352 6624 2470 6658
rect 2504 6624 2538 6658
rect 2572 6624 2606 6658
rect 2640 6624 2674 6658
rect 2708 6624 2742 6658
rect 2776 6624 2810 6658
rect 2844 6624 2878 6658
rect 2912 6624 2946 6658
rect 2980 6624 3014 6658
rect 3048 6624 3082 6658
rect 3116 6624 3150 6658
rect 3184 6624 3218 6658
rect 3252 6624 3286 6658
rect 3320 6624 3354 6658
rect 3388 6624 3422 6658
rect 3456 6624 3574 6658
rect 2352 6548 2386 6624
rect 3540 6553 3574 6624
rect 3873 6624 3991 6658
rect 4025 6624 4059 6658
rect 4093 6624 4127 6658
rect 4161 6624 4195 6658
rect 4229 6624 4263 6658
rect 4297 6624 4331 6658
rect 4365 6624 4399 6658
rect 4433 6624 4467 6658
rect 4501 6624 4535 6658
rect 4569 6624 4603 6658
rect 4637 6624 4671 6658
rect 4705 6624 4739 6658
rect 4773 6624 4807 6658
rect 4841 6624 4875 6658
rect 4909 6624 4943 6658
rect 4977 6624 5095 6658
rect 3675 6588 3691 6622
rect 3725 6588 3741 6622
rect 2352 6480 2386 6514
rect 2352 6412 2386 6446
rect 2466 6511 2500 6550
rect 2466 6438 2500 6477
rect 2562 6511 2596 6550
rect 2562 6438 2596 6477
rect 2658 6511 2692 6550
rect 2658 6438 2692 6477
rect 2754 6511 2788 6550
rect 2754 6438 2788 6477
rect 2850 6511 2884 6550
rect 2850 6438 2884 6477
rect 2946 6511 2980 6550
rect 2946 6438 2980 6477
rect 3042 6511 3076 6550
rect 3042 6438 3076 6477
rect 3138 6511 3172 6550
rect 3138 6438 3172 6477
rect 3234 6511 3268 6550
rect 3234 6438 3268 6477
rect 3330 6511 3364 6550
rect 3330 6438 3364 6477
rect 3426 6511 3460 6550
rect 3426 6438 3460 6477
rect 3540 6481 3574 6514
rect 3647 6538 3681 6554
rect 3647 6446 3681 6462
rect 3735 6538 3769 6554
rect 3735 6446 3769 6462
rect 3873 6548 3907 6624
rect 5061 6553 5095 6624
rect 3873 6480 3907 6514
rect 3540 6412 3574 6446
rect 2352 6302 2386 6378
rect 2450 6366 2466 6400
rect 2500 6366 2516 6400
rect 2642 6366 2658 6400
rect 2692 6366 2708 6400
rect 2834 6366 2850 6400
rect 2884 6366 2900 6400
rect 3026 6366 3042 6400
rect 3076 6366 3092 6400
rect 3218 6366 3234 6400
rect 3268 6366 3284 6400
rect 3410 6366 3426 6400
rect 3460 6366 3476 6400
rect 3540 6302 3574 6375
rect 2352 6268 2470 6302
rect 2504 6268 2538 6302
rect 2572 6268 2606 6302
rect 2640 6268 2674 6302
rect 2708 6268 2742 6302
rect 2776 6268 2810 6302
rect 2844 6268 2878 6302
rect 2912 6268 2946 6302
rect 2980 6268 3014 6302
rect 3048 6268 3082 6302
rect 3116 6268 3150 6302
rect 3184 6268 3218 6302
rect 3252 6268 3286 6302
rect 3320 6268 3354 6302
rect 3388 6268 3422 6302
rect 3456 6268 3574 6302
rect 3873 6412 3907 6446
rect 3987 6511 4021 6550
rect 3987 6438 4021 6477
rect 4083 6511 4117 6550
rect 4083 6438 4117 6477
rect 4179 6511 4213 6550
rect 4179 6438 4213 6477
rect 4275 6511 4309 6550
rect 4275 6438 4309 6477
rect 4371 6511 4405 6550
rect 4371 6438 4405 6477
rect 4467 6511 4501 6550
rect 4467 6438 4501 6477
rect 4563 6511 4597 6550
rect 4563 6438 4597 6477
rect 4659 6511 4693 6550
rect 4659 6438 4693 6477
rect 4755 6511 4789 6550
rect 4755 6438 4789 6477
rect 4851 6511 4885 6550
rect 4851 6438 4885 6477
rect 4947 6511 4981 6550
rect 4947 6438 4981 6477
rect 5061 6481 5095 6514
rect 5340 6629 5348 6663
rect 5382 6629 5386 6663
rect 5420 6668 5486 6679
rect 5420 6665 5450 6668
rect 5420 6631 5436 6665
rect 5484 6634 5486 6668
rect 5470 6631 5486 6634
rect 5340 6593 5386 6629
rect 5340 6581 5406 6593
rect 5340 6547 5356 6581
rect 5390 6547 5406 6581
rect 5340 6513 5406 6547
rect 5340 6479 5356 6513
rect 5390 6479 5406 6513
rect 5340 6467 5406 6479
rect 5440 6581 5486 6597
rect 5474 6547 5486 6581
rect 5440 6513 5486 6547
rect 5474 6479 5486 6513
rect 5061 6412 5095 6446
rect 5440 6433 5486 6479
rect 3873 6302 3907 6378
rect 3971 6366 3987 6400
rect 4021 6366 4037 6400
rect 4163 6366 4179 6400
rect 4213 6366 4229 6400
rect 4355 6366 4371 6400
rect 4405 6366 4421 6400
rect 4547 6366 4563 6400
rect 4597 6366 4613 6400
rect 4739 6366 4755 6400
rect 4789 6366 4805 6400
rect 4931 6366 4947 6400
rect 4981 6366 4997 6400
rect 5274 6399 5303 6433
rect 5337 6399 5395 6433
rect 5429 6399 5487 6433
rect 5521 6399 5550 6433
rect 5061 6302 5095 6375
rect 3873 6268 3991 6302
rect 4025 6268 4059 6302
rect 4093 6268 4127 6302
rect 4161 6268 4195 6302
rect 4229 6268 4263 6302
rect 4297 6268 4331 6302
rect 4365 6268 4399 6302
rect 4433 6268 4467 6302
rect 4501 6268 4535 6302
rect 4569 6268 4603 6302
rect 4637 6268 4671 6302
rect 4705 6268 4739 6302
rect 4773 6268 4807 6302
rect 4841 6268 4875 6302
rect 4909 6268 4943 6302
rect 4977 6268 5095 6302
rect 199 5985 317 6019
rect 351 5985 385 6019
rect 419 5985 453 6019
rect 487 5985 521 6019
rect 555 5985 589 6019
rect 623 5985 657 6019
rect 691 5985 725 6019
rect 759 5985 793 6019
rect 827 5985 861 6019
rect 895 5985 929 6019
rect 963 5985 997 6019
rect 1031 5985 1065 6019
rect 1099 5985 1133 6019
rect 1167 5985 1201 6019
rect 1235 5985 1269 6019
rect 1303 5985 1421 6019
rect 199 5917 233 5985
rect 1387 5917 1421 5985
rect 297 5883 313 5917
rect 347 5883 363 5917
rect 489 5883 505 5917
rect 539 5883 555 5917
rect 681 5883 697 5917
rect 731 5883 747 5917
rect 873 5883 889 5917
rect 923 5883 939 5917
rect 1065 5883 1081 5917
rect 1115 5883 1131 5917
rect 1257 5883 1273 5917
rect 1307 5883 1323 5917
rect 199 5849 233 5883
rect 1387 5849 1421 5857
rect 199 5781 233 5815
rect 199 5713 233 5747
rect 199 5645 233 5679
rect 199 5577 233 5611
rect 313 5818 347 5839
rect 313 5750 347 5754
rect 313 5644 347 5648
rect 313 5559 347 5580
rect 409 5818 443 5839
rect 409 5750 443 5754
rect 409 5644 443 5648
rect 409 5559 443 5580
rect 505 5818 539 5839
rect 505 5750 539 5754
rect 505 5644 539 5648
rect 505 5559 539 5580
rect 601 5818 635 5839
rect 601 5750 635 5754
rect 601 5644 635 5648
rect 601 5559 635 5580
rect 697 5818 731 5839
rect 697 5750 731 5754
rect 697 5644 731 5648
rect 697 5559 731 5580
rect 793 5818 827 5839
rect 793 5750 827 5754
rect 793 5644 827 5648
rect 793 5559 827 5580
rect 889 5818 923 5839
rect 889 5750 923 5754
rect 889 5644 923 5648
rect 889 5559 923 5580
rect 985 5818 1019 5839
rect 985 5750 1019 5754
rect 985 5644 1019 5648
rect 985 5559 1019 5580
rect 1081 5818 1115 5839
rect 1081 5750 1115 5754
rect 1081 5644 1115 5648
rect 1081 5559 1115 5580
rect 1177 5818 1211 5839
rect 1177 5750 1211 5754
rect 1177 5644 1211 5648
rect 1177 5559 1211 5580
rect 1273 5818 1307 5839
rect 1273 5750 1307 5754
rect 1273 5644 1307 5648
rect 1273 5559 1307 5580
rect 1387 5781 1421 5785
rect 1387 5675 1421 5679
rect 1387 5603 1421 5611
rect 199 5475 233 5543
rect 1387 5475 1421 5543
rect 199 5441 317 5475
rect 351 5441 385 5475
rect 419 5441 453 5475
rect 487 5441 521 5475
rect 555 5441 589 5475
rect 623 5441 657 5475
rect 691 5441 725 5475
rect 759 5441 793 5475
rect 827 5441 861 5475
rect 895 5441 929 5475
rect 963 5441 997 5475
rect 1031 5441 1065 5475
rect 1099 5441 1133 5475
rect 1167 5441 1201 5475
rect 1235 5441 1269 5475
rect 1303 5441 1421 5475
rect 2352 5989 2470 6023
rect 2504 5989 2538 6023
rect 2572 5989 2606 6023
rect 2640 5989 2674 6023
rect 2708 5989 2742 6023
rect 2776 5989 2810 6023
rect 2844 5989 2878 6023
rect 2912 5989 2946 6023
rect 2980 5989 3014 6023
rect 3048 5989 3082 6023
rect 3116 5989 3150 6023
rect 3184 5989 3218 6023
rect 3252 5989 3286 6023
rect 3320 5989 3354 6023
rect 3388 5989 3422 6023
rect 3456 5989 3574 6023
rect 2352 5921 2386 5989
rect 3540 5921 3574 5989
rect 2450 5887 2466 5921
rect 2500 5887 2516 5921
rect 2642 5887 2658 5921
rect 2692 5887 2708 5921
rect 2834 5887 2850 5921
rect 2884 5887 2900 5921
rect 3026 5887 3042 5921
rect 3076 5887 3092 5921
rect 3218 5887 3234 5921
rect 3268 5887 3284 5921
rect 3410 5887 3426 5921
rect 3460 5887 3476 5921
rect 2352 5853 2386 5887
rect 3540 5853 3574 5861
rect 2352 5785 2386 5819
rect 2352 5717 2386 5751
rect 2352 5649 2386 5683
rect 2352 5581 2386 5615
rect 2466 5822 2500 5843
rect 2466 5754 2500 5758
rect 2466 5648 2500 5652
rect 2466 5563 2500 5584
rect 2562 5822 2596 5843
rect 2562 5754 2596 5758
rect 2562 5648 2596 5652
rect 2562 5563 2596 5584
rect 2658 5822 2692 5843
rect 2658 5754 2692 5758
rect 2658 5648 2692 5652
rect 2658 5563 2692 5584
rect 2754 5822 2788 5843
rect 2754 5754 2788 5758
rect 2754 5648 2788 5652
rect 2754 5563 2788 5584
rect 2850 5822 2884 5843
rect 2850 5754 2884 5758
rect 2850 5648 2884 5652
rect 2850 5563 2884 5584
rect 2946 5822 2980 5843
rect 2946 5754 2980 5758
rect 2946 5648 2980 5652
rect 2946 5563 2980 5584
rect 3042 5822 3076 5843
rect 3042 5754 3076 5758
rect 3042 5648 3076 5652
rect 3042 5563 3076 5584
rect 3138 5822 3172 5843
rect 3138 5754 3172 5758
rect 3138 5648 3172 5652
rect 3138 5563 3172 5584
rect 3234 5822 3268 5843
rect 3234 5754 3268 5758
rect 3234 5648 3268 5652
rect 3234 5563 3268 5584
rect 3330 5822 3364 5843
rect 3330 5754 3364 5758
rect 3330 5648 3364 5652
rect 3330 5563 3364 5584
rect 3426 5822 3460 5843
rect 3426 5754 3460 5758
rect 3426 5648 3460 5652
rect 3426 5563 3460 5584
rect 3540 5785 3574 5789
rect 3540 5679 3574 5683
rect 3540 5607 3574 5615
rect 2352 5479 2386 5547
rect 3540 5479 3574 5547
rect 2352 5445 2470 5479
rect 2504 5445 2538 5479
rect 2572 5445 2606 5479
rect 2640 5445 2674 5479
rect 2708 5445 2742 5479
rect 2776 5445 2810 5479
rect 2844 5445 2878 5479
rect 2912 5445 2946 5479
rect 2980 5445 3014 5479
rect 3048 5445 3082 5479
rect 3116 5445 3150 5479
rect 3184 5445 3218 5479
rect 3252 5445 3286 5479
rect 3320 5445 3354 5479
rect 3388 5445 3422 5479
rect 3456 5445 3574 5479
rect 3873 5989 3991 6023
rect 4025 5989 4059 6023
rect 4093 5989 4127 6023
rect 4161 5989 4195 6023
rect 4229 5989 4263 6023
rect 4297 5989 4331 6023
rect 4365 5989 4399 6023
rect 4433 5989 4467 6023
rect 4501 5989 4535 6023
rect 4569 5989 4603 6023
rect 4637 5989 4671 6023
rect 4705 5989 4739 6023
rect 4773 5989 4807 6023
rect 4841 5989 4875 6023
rect 4909 5989 4943 6023
rect 4977 5989 5095 6023
rect 3873 5921 3907 5989
rect 5061 5921 5095 5989
rect 3971 5887 3987 5921
rect 4021 5887 4037 5921
rect 4163 5887 4179 5921
rect 4213 5887 4229 5921
rect 4355 5887 4371 5921
rect 4405 5887 4421 5921
rect 4547 5887 4563 5921
rect 4597 5887 4613 5921
rect 4739 5887 4755 5921
rect 4789 5887 4805 5921
rect 4931 5887 4947 5921
rect 4981 5887 4997 5921
rect 3873 5853 3907 5887
rect 5061 5853 5095 5861
rect 3873 5785 3907 5819
rect 3873 5717 3907 5751
rect 3873 5649 3907 5683
rect 3873 5581 3907 5615
rect 3987 5822 4021 5843
rect 3987 5754 4021 5758
rect 3987 5648 4021 5652
rect 3987 5563 4021 5584
rect 4083 5822 4117 5843
rect 4083 5754 4117 5758
rect 4083 5648 4117 5652
rect 4083 5563 4117 5584
rect 4179 5822 4213 5843
rect 4179 5754 4213 5758
rect 4179 5648 4213 5652
rect 4179 5563 4213 5584
rect 4275 5822 4309 5843
rect 4275 5754 4309 5758
rect 4275 5648 4309 5652
rect 4275 5563 4309 5584
rect 4371 5822 4405 5843
rect 4371 5754 4405 5758
rect 4371 5648 4405 5652
rect 4371 5563 4405 5584
rect 4467 5822 4501 5843
rect 4467 5754 4501 5758
rect 4467 5648 4501 5652
rect 4467 5563 4501 5584
rect 4563 5822 4597 5843
rect 4563 5754 4597 5758
rect 4563 5648 4597 5652
rect 4563 5563 4597 5584
rect 4659 5822 4693 5843
rect 4659 5754 4693 5758
rect 4659 5648 4693 5652
rect 4659 5563 4693 5584
rect 4755 5822 4789 5843
rect 4755 5754 4789 5758
rect 4755 5648 4789 5652
rect 4755 5563 4789 5584
rect 4851 5822 4885 5843
rect 4851 5754 4885 5758
rect 4851 5648 4885 5652
rect 4851 5563 4885 5584
rect 4947 5822 4981 5843
rect 4947 5754 4981 5758
rect 4947 5648 4981 5652
rect 4947 5563 4981 5584
rect 5061 5785 5095 5789
rect 5061 5679 5095 5683
rect 5274 5656 5303 5690
rect 5337 5656 5395 5690
rect 5429 5656 5487 5690
rect 5521 5656 5550 5690
rect 5061 5607 5095 5615
rect 3873 5479 3907 5547
rect 5061 5479 5095 5547
rect 3873 5445 3991 5479
rect 4025 5445 4059 5479
rect 4093 5445 4127 5479
rect 4161 5445 4195 5479
rect 4229 5445 4263 5479
rect 4297 5445 4331 5479
rect 4365 5445 4399 5479
rect 4433 5445 4467 5479
rect 4501 5445 4535 5479
rect 4569 5445 4603 5479
rect 4637 5445 4671 5479
rect 4705 5445 4739 5479
rect 4773 5445 4807 5479
rect 4841 5445 4875 5479
rect 4909 5445 4943 5479
rect 4977 5445 5095 5479
rect 5340 5614 5406 5622
rect 5340 5580 5356 5614
rect 5390 5580 5406 5614
rect 5340 5546 5406 5580
rect 5340 5512 5356 5546
rect 5390 5512 5406 5546
rect 5340 5478 5406 5512
rect 5340 5444 5356 5478
rect 5390 5444 5406 5478
rect 5340 5426 5406 5444
rect 5440 5614 5482 5656
rect 5474 5580 5482 5614
rect 5440 5546 5482 5580
rect 5474 5512 5482 5546
rect 5440 5478 5482 5512
rect 5474 5444 5482 5478
rect 5440 5428 5482 5444
rect 5340 5376 5386 5426
rect 199 5333 317 5367
rect 351 5333 385 5367
rect 419 5333 453 5367
rect 487 5333 521 5367
rect 555 5333 589 5367
rect 623 5333 657 5367
rect 691 5333 725 5367
rect 759 5333 793 5367
rect 827 5333 861 5367
rect 895 5333 929 5367
rect 963 5333 997 5367
rect 1031 5333 1065 5367
rect 1099 5333 1133 5367
rect 1167 5333 1201 5367
rect 1235 5333 1269 5367
rect 1303 5333 1421 5367
rect 199 5257 233 5333
rect 1387 5262 1421 5333
rect 199 5189 233 5223
rect 199 5121 233 5155
rect 313 5220 347 5259
rect 313 5147 347 5186
rect 409 5220 443 5259
rect 409 5147 443 5186
rect 505 5220 539 5259
rect 505 5147 539 5186
rect 601 5220 635 5259
rect 601 5147 635 5186
rect 697 5220 731 5259
rect 697 5147 731 5186
rect 793 5220 827 5259
rect 793 5147 827 5186
rect 889 5220 923 5259
rect 889 5147 923 5186
rect 985 5220 1019 5259
rect 985 5147 1019 5186
rect 1081 5220 1115 5259
rect 1081 5147 1115 5186
rect 1177 5220 1211 5259
rect 1177 5147 1211 5186
rect 1273 5220 1307 5259
rect 1273 5147 1307 5186
rect 1387 5190 1421 5223
rect 1387 5121 1421 5155
rect 199 5011 233 5087
rect 297 5075 313 5109
rect 347 5075 363 5109
rect 489 5075 505 5109
rect 539 5075 555 5109
rect 681 5075 697 5109
rect 731 5075 747 5109
rect 873 5075 889 5109
rect 923 5075 939 5109
rect 1065 5075 1081 5109
rect 1115 5075 1131 5109
rect 1257 5075 1273 5109
rect 1307 5075 1323 5109
rect 1387 5011 1421 5084
rect 199 4977 317 5011
rect 351 4977 385 5011
rect 419 4977 453 5011
rect 487 4977 521 5011
rect 555 4977 589 5011
rect 623 4977 657 5011
rect 691 4977 725 5011
rect 759 4977 793 5011
rect 827 4977 861 5011
rect 895 4977 929 5011
rect 963 4977 997 5011
rect 1031 4977 1065 5011
rect 1099 4977 1133 5011
rect 1167 4977 1201 5011
rect 1235 4977 1269 5011
rect 1303 4977 1421 5011
rect 2352 5337 2470 5371
rect 2504 5337 2538 5371
rect 2572 5337 2606 5371
rect 2640 5337 2674 5371
rect 2708 5337 2742 5371
rect 2776 5337 2810 5371
rect 2844 5337 2878 5371
rect 2912 5337 2946 5371
rect 2980 5337 3014 5371
rect 3048 5337 3082 5371
rect 3116 5337 3150 5371
rect 3184 5337 3218 5371
rect 3252 5337 3286 5371
rect 3320 5337 3354 5371
rect 3388 5337 3422 5371
rect 3456 5337 3574 5371
rect 2352 5261 2386 5337
rect 3540 5266 3574 5337
rect 3873 5337 3991 5371
rect 4025 5337 4059 5371
rect 4093 5337 4127 5371
rect 4161 5337 4195 5371
rect 4229 5337 4263 5371
rect 4297 5337 4331 5371
rect 4365 5337 4399 5371
rect 4433 5337 4467 5371
rect 4501 5337 4535 5371
rect 4569 5337 4603 5371
rect 4637 5337 4671 5371
rect 4705 5337 4739 5371
rect 4773 5337 4807 5371
rect 4841 5337 4875 5371
rect 4909 5337 4943 5371
rect 4977 5337 5095 5371
rect 3675 5301 3691 5335
rect 3725 5301 3741 5335
rect 2352 5193 2386 5227
rect 2352 5125 2386 5159
rect 2466 5224 2500 5263
rect 2466 5151 2500 5190
rect 2562 5224 2596 5263
rect 2562 5151 2596 5190
rect 2658 5224 2692 5263
rect 2658 5151 2692 5190
rect 2754 5224 2788 5263
rect 2754 5151 2788 5190
rect 2850 5224 2884 5263
rect 2850 5151 2884 5190
rect 2946 5224 2980 5263
rect 2946 5151 2980 5190
rect 3042 5224 3076 5263
rect 3042 5151 3076 5190
rect 3138 5224 3172 5263
rect 3138 5151 3172 5190
rect 3234 5224 3268 5263
rect 3234 5151 3268 5190
rect 3330 5224 3364 5263
rect 3330 5151 3364 5190
rect 3426 5224 3460 5263
rect 3426 5151 3460 5190
rect 3540 5194 3574 5227
rect 3647 5251 3681 5267
rect 3647 5159 3681 5175
rect 3735 5251 3769 5267
rect 3735 5159 3769 5175
rect 3873 5261 3907 5337
rect 5061 5266 5095 5337
rect 3873 5193 3907 5227
rect 3540 5125 3574 5159
rect 2352 5015 2386 5091
rect 2450 5079 2466 5113
rect 2500 5079 2516 5113
rect 2642 5079 2658 5113
rect 2692 5079 2708 5113
rect 2834 5079 2850 5113
rect 2884 5079 2900 5113
rect 3026 5079 3042 5113
rect 3076 5079 3092 5113
rect 3218 5079 3234 5113
rect 3268 5079 3284 5113
rect 3410 5079 3426 5113
rect 3460 5079 3476 5113
rect 3540 5015 3574 5088
rect 2352 4981 2470 5015
rect 2504 4981 2538 5015
rect 2572 4981 2606 5015
rect 2640 4981 2674 5015
rect 2708 4981 2742 5015
rect 2776 4981 2810 5015
rect 2844 4981 2878 5015
rect 2912 4981 2946 5015
rect 2980 4981 3014 5015
rect 3048 4981 3082 5015
rect 3116 4981 3150 5015
rect 3184 4981 3218 5015
rect 3252 4981 3286 5015
rect 3320 4981 3354 5015
rect 3388 4981 3422 5015
rect 3456 4981 3574 5015
rect 3873 5125 3907 5159
rect 3987 5224 4021 5263
rect 3987 5151 4021 5190
rect 4083 5224 4117 5263
rect 4083 5151 4117 5190
rect 4179 5224 4213 5263
rect 4179 5151 4213 5190
rect 4275 5224 4309 5263
rect 4275 5151 4309 5190
rect 4371 5224 4405 5263
rect 4371 5151 4405 5190
rect 4467 5224 4501 5263
rect 4467 5151 4501 5190
rect 4563 5224 4597 5263
rect 4563 5151 4597 5190
rect 4659 5224 4693 5263
rect 4659 5151 4693 5190
rect 4755 5224 4789 5263
rect 4755 5151 4789 5190
rect 4851 5224 4885 5263
rect 4851 5151 4885 5190
rect 4947 5224 4981 5263
rect 4947 5151 4981 5190
rect 5061 5194 5095 5227
rect 5340 5342 5348 5376
rect 5382 5342 5386 5376
rect 5420 5381 5486 5392
rect 5420 5378 5450 5381
rect 5420 5344 5436 5378
rect 5484 5347 5486 5381
rect 5470 5344 5486 5347
rect 5340 5306 5386 5342
rect 5340 5294 5406 5306
rect 5340 5260 5356 5294
rect 5390 5260 5406 5294
rect 5340 5226 5406 5260
rect 5340 5192 5356 5226
rect 5390 5192 5406 5226
rect 5340 5180 5406 5192
rect 5440 5294 5486 5310
rect 5474 5260 5486 5294
rect 5440 5226 5486 5260
rect 5474 5192 5486 5226
rect 5061 5125 5095 5159
rect 5440 5146 5486 5192
rect 3873 5015 3907 5091
rect 3971 5079 3987 5113
rect 4021 5079 4037 5113
rect 4163 5079 4179 5113
rect 4213 5079 4229 5113
rect 4355 5079 4371 5113
rect 4405 5079 4421 5113
rect 4547 5079 4563 5113
rect 4597 5079 4613 5113
rect 4739 5079 4755 5113
rect 4789 5079 4805 5113
rect 4931 5079 4947 5113
rect 4981 5079 4997 5113
rect 5274 5112 5303 5146
rect 5337 5112 5395 5146
rect 5429 5112 5487 5146
rect 5521 5112 5550 5146
rect 5061 5015 5095 5088
rect 3873 4981 3991 5015
rect 4025 4981 4059 5015
rect 4093 4981 4127 5015
rect 4161 4981 4195 5015
rect 4229 4981 4263 5015
rect 4297 4981 4331 5015
rect 4365 4981 4399 5015
rect 4433 4981 4467 5015
rect 4501 4981 4535 5015
rect 4569 4981 4603 5015
rect 4637 4981 4671 5015
rect 4705 4981 4739 5015
rect 4773 4981 4807 5015
rect 4841 4981 4875 5015
rect 4909 4981 4943 5015
rect 4977 4981 5095 5015
rect 199 4698 317 4732
rect 351 4698 385 4732
rect 419 4698 453 4732
rect 487 4698 521 4732
rect 555 4698 589 4732
rect 623 4698 657 4732
rect 691 4698 725 4732
rect 759 4698 793 4732
rect 827 4698 861 4732
rect 895 4698 929 4732
rect 963 4698 997 4732
rect 1031 4698 1065 4732
rect 1099 4698 1133 4732
rect 1167 4698 1201 4732
rect 1235 4698 1269 4732
rect 1303 4698 1421 4732
rect 199 4630 233 4698
rect 1387 4630 1421 4698
rect 297 4596 313 4630
rect 347 4596 363 4630
rect 489 4596 505 4630
rect 539 4596 555 4630
rect 681 4596 697 4630
rect 731 4596 747 4630
rect 873 4596 889 4630
rect 923 4596 939 4630
rect 1065 4596 1081 4630
rect 1115 4596 1131 4630
rect 1257 4596 1273 4630
rect 1307 4596 1323 4630
rect 199 4562 233 4596
rect 1387 4562 1421 4570
rect 199 4494 233 4528
rect 199 4426 233 4460
rect 199 4358 233 4392
rect 199 4290 233 4324
rect 313 4531 347 4552
rect 313 4463 347 4467
rect 313 4357 347 4361
rect 313 4272 347 4293
rect 409 4531 443 4552
rect 409 4463 443 4467
rect 409 4357 443 4361
rect 409 4272 443 4293
rect 505 4531 539 4552
rect 505 4463 539 4467
rect 505 4357 539 4361
rect 505 4272 539 4293
rect 601 4531 635 4552
rect 601 4463 635 4467
rect 601 4357 635 4361
rect 601 4272 635 4293
rect 697 4531 731 4552
rect 697 4463 731 4467
rect 697 4357 731 4361
rect 697 4272 731 4293
rect 793 4531 827 4552
rect 793 4463 827 4467
rect 793 4357 827 4361
rect 793 4272 827 4293
rect 889 4531 923 4552
rect 889 4463 923 4467
rect 889 4357 923 4361
rect 889 4272 923 4293
rect 985 4531 1019 4552
rect 985 4463 1019 4467
rect 985 4357 1019 4361
rect 985 4272 1019 4293
rect 1081 4531 1115 4552
rect 1081 4463 1115 4467
rect 1081 4357 1115 4361
rect 1081 4272 1115 4293
rect 1177 4531 1211 4552
rect 1177 4463 1211 4467
rect 1177 4357 1211 4361
rect 1177 4272 1211 4293
rect 1273 4531 1307 4552
rect 1273 4463 1307 4467
rect 1273 4357 1307 4361
rect 1273 4272 1307 4293
rect 1387 4494 1421 4498
rect 1387 4388 1421 4392
rect 1387 4316 1421 4324
rect 199 4188 233 4256
rect 1387 4188 1421 4256
rect 199 4154 317 4188
rect 351 4154 385 4188
rect 419 4154 453 4188
rect 487 4154 521 4188
rect 555 4154 589 4188
rect 623 4154 657 4188
rect 691 4154 725 4188
rect 759 4154 793 4188
rect 827 4154 861 4188
rect 895 4154 929 4188
rect 963 4154 997 4188
rect 1031 4154 1065 4188
rect 1099 4154 1133 4188
rect 1167 4154 1201 4188
rect 1235 4154 1269 4188
rect 1303 4154 1421 4188
rect 2352 4702 2470 4736
rect 2504 4702 2538 4736
rect 2572 4702 2606 4736
rect 2640 4702 2674 4736
rect 2708 4702 2742 4736
rect 2776 4702 2810 4736
rect 2844 4702 2878 4736
rect 2912 4702 2946 4736
rect 2980 4702 3014 4736
rect 3048 4702 3082 4736
rect 3116 4702 3150 4736
rect 3184 4702 3218 4736
rect 3252 4702 3286 4736
rect 3320 4702 3354 4736
rect 3388 4702 3422 4736
rect 3456 4702 3574 4736
rect 2352 4634 2386 4702
rect 3540 4634 3574 4702
rect 2450 4600 2466 4634
rect 2500 4600 2516 4634
rect 2642 4600 2658 4634
rect 2692 4600 2708 4634
rect 2834 4600 2850 4634
rect 2884 4600 2900 4634
rect 3026 4600 3042 4634
rect 3076 4600 3092 4634
rect 3218 4600 3234 4634
rect 3268 4600 3284 4634
rect 3410 4600 3426 4634
rect 3460 4600 3476 4634
rect 2352 4566 2386 4600
rect 3540 4566 3574 4574
rect 2352 4498 2386 4532
rect 2352 4430 2386 4464
rect 2352 4362 2386 4396
rect 2352 4294 2386 4328
rect 2466 4535 2500 4556
rect 2466 4467 2500 4471
rect 2466 4361 2500 4365
rect 2466 4276 2500 4297
rect 2562 4535 2596 4556
rect 2562 4467 2596 4471
rect 2562 4361 2596 4365
rect 2562 4276 2596 4297
rect 2658 4535 2692 4556
rect 2658 4467 2692 4471
rect 2658 4361 2692 4365
rect 2658 4276 2692 4297
rect 2754 4535 2788 4556
rect 2754 4467 2788 4471
rect 2754 4361 2788 4365
rect 2754 4276 2788 4297
rect 2850 4535 2884 4556
rect 2850 4467 2884 4471
rect 2850 4361 2884 4365
rect 2850 4276 2884 4297
rect 2946 4535 2980 4556
rect 2946 4467 2980 4471
rect 2946 4361 2980 4365
rect 2946 4276 2980 4297
rect 3042 4535 3076 4556
rect 3042 4467 3076 4471
rect 3042 4361 3076 4365
rect 3042 4276 3076 4297
rect 3138 4535 3172 4556
rect 3138 4467 3172 4471
rect 3138 4361 3172 4365
rect 3138 4276 3172 4297
rect 3234 4535 3268 4556
rect 3234 4467 3268 4471
rect 3234 4361 3268 4365
rect 3234 4276 3268 4297
rect 3330 4535 3364 4556
rect 3330 4467 3364 4471
rect 3330 4361 3364 4365
rect 3330 4276 3364 4297
rect 3426 4535 3460 4556
rect 3426 4467 3460 4471
rect 3426 4361 3460 4365
rect 3426 4276 3460 4297
rect 3540 4498 3574 4502
rect 3540 4392 3574 4396
rect 3540 4320 3574 4328
rect 2352 4192 2386 4260
rect 3540 4192 3574 4260
rect 2352 4158 2470 4192
rect 2504 4158 2538 4192
rect 2572 4158 2606 4192
rect 2640 4158 2674 4192
rect 2708 4158 2742 4192
rect 2776 4158 2810 4192
rect 2844 4158 2878 4192
rect 2912 4158 2946 4192
rect 2980 4158 3014 4192
rect 3048 4158 3082 4192
rect 3116 4158 3150 4192
rect 3184 4158 3218 4192
rect 3252 4158 3286 4192
rect 3320 4158 3354 4192
rect 3388 4158 3422 4192
rect 3456 4158 3574 4192
rect 3873 4702 3991 4736
rect 4025 4702 4059 4736
rect 4093 4702 4127 4736
rect 4161 4702 4195 4736
rect 4229 4702 4263 4736
rect 4297 4702 4331 4736
rect 4365 4702 4399 4736
rect 4433 4702 4467 4736
rect 4501 4702 4535 4736
rect 4569 4702 4603 4736
rect 4637 4702 4671 4736
rect 4705 4702 4739 4736
rect 4773 4702 4807 4736
rect 4841 4702 4875 4736
rect 4909 4702 4943 4736
rect 4977 4702 5095 4736
rect 3873 4634 3907 4702
rect 5061 4634 5095 4702
rect 3971 4600 3987 4634
rect 4021 4600 4037 4634
rect 4163 4600 4179 4634
rect 4213 4600 4229 4634
rect 4355 4600 4371 4634
rect 4405 4600 4421 4634
rect 4547 4600 4563 4634
rect 4597 4600 4613 4634
rect 4739 4600 4755 4634
rect 4789 4600 4805 4634
rect 4931 4600 4947 4634
rect 4981 4600 4997 4634
rect 3873 4566 3907 4600
rect 5061 4566 5095 4574
rect 3873 4498 3907 4532
rect 3873 4430 3907 4464
rect 3873 4362 3907 4396
rect 3873 4294 3907 4328
rect 3987 4535 4021 4556
rect 3987 4467 4021 4471
rect 3987 4361 4021 4365
rect 3987 4276 4021 4297
rect 4083 4535 4117 4556
rect 4083 4467 4117 4471
rect 4083 4361 4117 4365
rect 4083 4276 4117 4297
rect 4179 4535 4213 4556
rect 4179 4467 4213 4471
rect 4179 4361 4213 4365
rect 4179 4276 4213 4297
rect 4275 4535 4309 4556
rect 4275 4467 4309 4471
rect 4275 4361 4309 4365
rect 4275 4276 4309 4297
rect 4371 4535 4405 4556
rect 4371 4467 4405 4471
rect 4371 4361 4405 4365
rect 4371 4276 4405 4297
rect 4467 4535 4501 4556
rect 4467 4467 4501 4471
rect 4467 4361 4501 4365
rect 4467 4276 4501 4297
rect 4563 4535 4597 4556
rect 4563 4467 4597 4471
rect 4563 4361 4597 4365
rect 4563 4276 4597 4297
rect 4659 4535 4693 4556
rect 4659 4467 4693 4471
rect 4659 4361 4693 4365
rect 4659 4276 4693 4297
rect 4755 4535 4789 4556
rect 4755 4467 4789 4471
rect 4755 4361 4789 4365
rect 4755 4276 4789 4297
rect 4851 4535 4885 4556
rect 4851 4467 4885 4471
rect 4851 4361 4885 4365
rect 4851 4276 4885 4297
rect 4947 4535 4981 4556
rect 4947 4467 4981 4471
rect 4947 4361 4981 4365
rect 4947 4276 4981 4297
rect 5061 4498 5095 4502
rect 5061 4392 5095 4396
rect 5274 4369 5303 4403
rect 5337 4369 5395 4403
rect 5429 4369 5487 4403
rect 5521 4369 5550 4403
rect 5061 4320 5095 4328
rect 3873 4192 3907 4260
rect 5061 4192 5095 4260
rect 3873 4158 3991 4192
rect 4025 4158 4059 4192
rect 4093 4158 4127 4192
rect 4161 4158 4195 4192
rect 4229 4158 4263 4192
rect 4297 4158 4331 4192
rect 4365 4158 4399 4192
rect 4433 4158 4467 4192
rect 4501 4158 4535 4192
rect 4569 4158 4603 4192
rect 4637 4158 4671 4192
rect 4705 4158 4739 4192
rect 4773 4158 4807 4192
rect 4841 4158 4875 4192
rect 4909 4158 4943 4192
rect 4977 4158 5095 4192
rect 5340 4327 5406 4335
rect 5340 4293 5356 4327
rect 5390 4293 5406 4327
rect 5340 4259 5406 4293
rect 5340 4225 5356 4259
rect 5390 4225 5406 4259
rect 5340 4191 5406 4225
rect 5340 4157 5356 4191
rect 5390 4157 5406 4191
rect 5340 4139 5406 4157
rect 5440 4327 5482 4369
rect 5474 4293 5482 4327
rect 5440 4259 5482 4293
rect 5474 4225 5482 4259
rect 5440 4191 5482 4225
rect 5474 4157 5482 4191
rect 5440 4141 5482 4157
rect 5340 4089 5386 4139
rect 199 4046 317 4080
rect 351 4046 385 4080
rect 419 4046 453 4080
rect 487 4046 521 4080
rect 555 4046 589 4080
rect 623 4046 657 4080
rect 691 4046 725 4080
rect 759 4046 793 4080
rect 827 4046 861 4080
rect 895 4046 929 4080
rect 963 4046 997 4080
rect 1031 4046 1065 4080
rect 1099 4046 1133 4080
rect 1167 4046 1201 4080
rect 1235 4046 1269 4080
rect 1303 4046 1421 4080
rect 199 3970 233 4046
rect 1387 3975 1421 4046
rect 199 3902 233 3936
rect 199 3834 233 3868
rect 313 3933 347 3972
rect 313 3860 347 3899
rect 409 3933 443 3972
rect 409 3860 443 3899
rect 505 3933 539 3972
rect 505 3860 539 3899
rect 601 3933 635 3972
rect 601 3860 635 3899
rect 697 3933 731 3972
rect 697 3860 731 3899
rect 793 3933 827 3972
rect 793 3860 827 3899
rect 889 3933 923 3972
rect 889 3860 923 3899
rect 985 3933 1019 3972
rect 985 3860 1019 3899
rect 1081 3933 1115 3972
rect 1081 3860 1115 3899
rect 1177 3933 1211 3972
rect 1177 3860 1211 3899
rect 1273 3933 1307 3972
rect 1273 3860 1307 3899
rect 1387 3903 1421 3936
rect 1387 3834 1421 3868
rect 199 3724 233 3800
rect 297 3788 313 3822
rect 347 3788 363 3822
rect 489 3788 505 3822
rect 539 3788 555 3822
rect 681 3788 697 3822
rect 731 3788 747 3822
rect 873 3788 889 3822
rect 923 3788 939 3822
rect 1065 3788 1081 3822
rect 1115 3788 1131 3822
rect 1257 3788 1273 3822
rect 1307 3788 1323 3822
rect 1387 3724 1421 3797
rect 199 3690 317 3724
rect 351 3690 385 3724
rect 419 3690 453 3724
rect 487 3690 521 3724
rect 555 3690 589 3724
rect 623 3690 657 3724
rect 691 3690 725 3724
rect 759 3690 793 3724
rect 827 3690 861 3724
rect 895 3690 929 3724
rect 963 3690 997 3724
rect 1031 3690 1065 3724
rect 1099 3690 1133 3724
rect 1167 3690 1201 3724
rect 1235 3690 1269 3724
rect 1303 3690 1421 3724
rect 2352 4050 2470 4084
rect 2504 4050 2538 4084
rect 2572 4050 2606 4084
rect 2640 4050 2674 4084
rect 2708 4050 2742 4084
rect 2776 4050 2810 4084
rect 2844 4050 2878 4084
rect 2912 4050 2946 4084
rect 2980 4050 3014 4084
rect 3048 4050 3082 4084
rect 3116 4050 3150 4084
rect 3184 4050 3218 4084
rect 3252 4050 3286 4084
rect 3320 4050 3354 4084
rect 3388 4050 3422 4084
rect 3456 4050 3574 4084
rect 2352 3974 2386 4050
rect 3540 3979 3574 4050
rect 3873 4050 3991 4084
rect 4025 4050 4059 4084
rect 4093 4050 4127 4084
rect 4161 4050 4195 4084
rect 4229 4050 4263 4084
rect 4297 4050 4331 4084
rect 4365 4050 4399 4084
rect 4433 4050 4467 4084
rect 4501 4050 4535 4084
rect 4569 4050 4603 4084
rect 4637 4050 4671 4084
rect 4705 4050 4739 4084
rect 4773 4050 4807 4084
rect 4841 4050 4875 4084
rect 4909 4050 4943 4084
rect 4977 4050 5095 4084
rect 3675 4014 3691 4048
rect 3725 4014 3741 4048
rect 2352 3906 2386 3940
rect 2352 3838 2386 3872
rect 2466 3937 2500 3976
rect 2466 3864 2500 3903
rect 2562 3937 2596 3976
rect 2562 3864 2596 3903
rect 2658 3937 2692 3976
rect 2658 3864 2692 3903
rect 2754 3937 2788 3976
rect 2754 3864 2788 3903
rect 2850 3937 2884 3976
rect 2850 3864 2884 3903
rect 2946 3937 2980 3976
rect 2946 3864 2980 3903
rect 3042 3937 3076 3976
rect 3042 3864 3076 3903
rect 3138 3937 3172 3976
rect 3138 3864 3172 3903
rect 3234 3937 3268 3976
rect 3234 3864 3268 3903
rect 3330 3937 3364 3976
rect 3330 3864 3364 3903
rect 3426 3937 3460 3976
rect 3426 3864 3460 3903
rect 3540 3907 3574 3940
rect 3647 3964 3681 3980
rect 3647 3872 3681 3888
rect 3735 3964 3769 3980
rect 3735 3872 3769 3888
rect 3873 3974 3907 4050
rect 5061 3979 5095 4050
rect 3873 3906 3907 3940
rect 3540 3838 3574 3872
rect 2352 3728 2386 3804
rect 2450 3792 2466 3826
rect 2500 3792 2516 3826
rect 2642 3792 2658 3826
rect 2692 3792 2708 3826
rect 2834 3792 2850 3826
rect 2884 3792 2900 3826
rect 3026 3792 3042 3826
rect 3076 3792 3092 3826
rect 3218 3792 3234 3826
rect 3268 3792 3284 3826
rect 3410 3792 3426 3826
rect 3460 3792 3476 3826
rect 3540 3728 3574 3801
rect 2352 3694 2470 3728
rect 2504 3694 2538 3728
rect 2572 3694 2606 3728
rect 2640 3694 2674 3728
rect 2708 3694 2742 3728
rect 2776 3694 2810 3728
rect 2844 3694 2878 3728
rect 2912 3694 2946 3728
rect 2980 3694 3014 3728
rect 3048 3694 3082 3728
rect 3116 3694 3150 3728
rect 3184 3694 3218 3728
rect 3252 3694 3286 3728
rect 3320 3694 3354 3728
rect 3388 3694 3422 3728
rect 3456 3694 3574 3728
rect 3873 3838 3907 3872
rect 3987 3937 4021 3976
rect 3987 3864 4021 3903
rect 4083 3937 4117 3976
rect 4083 3864 4117 3903
rect 4179 3937 4213 3976
rect 4179 3864 4213 3903
rect 4275 3937 4309 3976
rect 4275 3864 4309 3903
rect 4371 3937 4405 3976
rect 4371 3864 4405 3903
rect 4467 3937 4501 3976
rect 4467 3864 4501 3903
rect 4563 3937 4597 3976
rect 4563 3864 4597 3903
rect 4659 3937 4693 3976
rect 4659 3864 4693 3903
rect 4755 3937 4789 3976
rect 4755 3864 4789 3903
rect 4851 3937 4885 3976
rect 4851 3864 4885 3903
rect 4947 3937 4981 3976
rect 4947 3864 4981 3903
rect 5061 3907 5095 3940
rect 5340 4055 5348 4089
rect 5382 4055 5386 4089
rect 5420 4094 5486 4105
rect 5420 4091 5450 4094
rect 5420 4057 5436 4091
rect 5484 4060 5486 4094
rect 5470 4057 5486 4060
rect 5340 4019 5386 4055
rect 5340 4007 5406 4019
rect 5340 3973 5356 4007
rect 5390 3973 5406 4007
rect 5340 3939 5406 3973
rect 5340 3905 5356 3939
rect 5390 3905 5406 3939
rect 5340 3893 5406 3905
rect 5440 4007 5486 4023
rect 5474 3973 5486 4007
rect 5440 3939 5486 3973
rect 5474 3905 5486 3939
rect 5061 3838 5095 3872
rect 5440 3859 5486 3905
rect 3873 3728 3907 3804
rect 3971 3792 3987 3826
rect 4021 3792 4037 3826
rect 4163 3792 4179 3826
rect 4213 3792 4229 3826
rect 4355 3792 4371 3826
rect 4405 3792 4421 3826
rect 4547 3792 4563 3826
rect 4597 3792 4613 3826
rect 4739 3792 4755 3826
rect 4789 3792 4805 3826
rect 4931 3792 4947 3826
rect 4981 3792 4997 3826
rect 5274 3825 5303 3859
rect 5337 3825 5395 3859
rect 5429 3825 5487 3859
rect 5521 3825 5550 3859
rect 5061 3728 5095 3801
rect 3873 3694 3991 3728
rect 4025 3694 4059 3728
rect 4093 3694 4127 3728
rect 4161 3694 4195 3728
rect 4229 3694 4263 3728
rect 4297 3694 4331 3728
rect 4365 3694 4399 3728
rect 4433 3694 4467 3728
rect 4501 3694 4535 3728
rect 4569 3694 4603 3728
rect 4637 3694 4671 3728
rect 4705 3694 4739 3728
rect 4773 3694 4807 3728
rect 4841 3694 4875 3728
rect 4909 3694 4943 3728
rect 4977 3694 5095 3728
rect 199 3411 317 3445
rect 351 3411 385 3445
rect 419 3411 453 3445
rect 487 3411 521 3445
rect 555 3411 589 3445
rect 623 3411 657 3445
rect 691 3411 725 3445
rect 759 3411 793 3445
rect 827 3411 861 3445
rect 895 3411 929 3445
rect 963 3411 997 3445
rect 1031 3411 1065 3445
rect 1099 3411 1133 3445
rect 1167 3411 1201 3445
rect 1235 3411 1269 3445
rect 1303 3411 1421 3445
rect 199 3343 233 3411
rect 1387 3343 1421 3411
rect 297 3309 313 3343
rect 347 3309 363 3343
rect 489 3309 505 3343
rect 539 3309 555 3343
rect 681 3309 697 3343
rect 731 3309 747 3343
rect 873 3309 889 3343
rect 923 3309 939 3343
rect 1065 3309 1081 3343
rect 1115 3309 1131 3343
rect 1257 3309 1273 3343
rect 1307 3309 1323 3343
rect 199 3275 233 3309
rect 1387 3275 1421 3283
rect 199 3207 233 3241
rect 199 3139 233 3173
rect 199 3071 233 3105
rect 199 3003 233 3037
rect 313 3244 347 3265
rect 313 3176 347 3180
rect 313 3070 347 3074
rect 313 2985 347 3006
rect 409 3244 443 3265
rect 409 3176 443 3180
rect 409 3070 443 3074
rect 409 2985 443 3006
rect 505 3244 539 3265
rect 505 3176 539 3180
rect 505 3070 539 3074
rect 505 2985 539 3006
rect 601 3244 635 3265
rect 601 3176 635 3180
rect 601 3070 635 3074
rect 601 2985 635 3006
rect 697 3244 731 3265
rect 697 3176 731 3180
rect 697 3070 731 3074
rect 697 2985 731 3006
rect 793 3244 827 3265
rect 793 3176 827 3180
rect 793 3070 827 3074
rect 793 2985 827 3006
rect 889 3244 923 3265
rect 889 3176 923 3180
rect 889 3070 923 3074
rect 889 2985 923 3006
rect 985 3244 1019 3265
rect 985 3176 1019 3180
rect 985 3070 1019 3074
rect 985 2985 1019 3006
rect 1081 3244 1115 3265
rect 1081 3176 1115 3180
rect 1081 3070 1115 3074
rect 1081 2985 1115 3006
rect 1177 3244 1211 3265
rect 1177 3176 1211 3180
rect 1177 3070 1211 3074
rect 1177 2985 1211 3006
rect 1273 3244 1307 3265
rect 1273 3176 1307 3180
rect 1273 3070 1307 3074
rect 1273 2985 1307 3006
rect 1387 3207 1421 3211
rect 1387 3101 1421 3105
rect 1387 3029 1421 3037
rect 199 2901 233 2969
rect 1387 2901 1421 2969
rect 199 2867 317 2901
rect 351 2867 385 2901
rect 419 2867 453 2901
rect 487 2867 521 2901
rect 555 2867 589 2901
rect 623 2867 657 2901
rect 691 2867 725 2901
rect 759 2867 793 2901
rect 827 2867 861 2901
rect 895 2867 929 2901
rect 963 2867 997 2901
rect 1031 2867 1065 2901
rect 1099 2867 1133 2901
rect 1167 2867 1201 2901
rect 1235 2867 1269 2901
rect 1303 2867 1421 2901
rect 2352 3415 2470 3449
rect 2504 3415 2538 3449
rect 2572 3415 2606 3449
rect 2640 3415 2674 3449
rect 2708 3415 2742 3449
rect 2776 3415 2810 3449
rect 2844 3415 2878 3449
rect 2912 3415 2946 3449
rect 2980 3415 3014 3449
rect 3048 3415 3082 3449
rect 3116 3415 3150 3449
rect 3184 3415 3218 3449
rect 3252 3415 3286 3449
rect 3320 3415 3354 3449
rect 3388 3415 3422 3449
rect 3456 3415 3574 3449
rect 2352 3347 2386 3415
rect 3540 3347 3574 3415
rect 2450 3313 2466 3347
rect 2500 3313 2516 3347
rect 2642 3313 2658 3347
rect 2692 3313 2708 3347
rect 2834 3313 2850 3347
rect 2884 3313 2900 3347
rect 3026 3313 3042 3347
rect 3076 3313 3092 3347
rect 3218 3313 3234 3347
rect 3268 3313 3284 3347
rect 3410 3313 3426 3347
rect 3460 3313 3476 3347
rect 2352 3279 2386 3313
rect 3540 3279 3574 3287
rect 2352 3211 2386 3245
rect 2352 3143 2386 3177
rect 2352 3075 2386 3109
rect 2352 3007 2386 3041
rect 2466 3248 2500 3269
rect 2466 3180 2500 3184
rect 2466 3074 2500 3078
rect 2466 2989 2500 3010
rect 2562 3248 2596 3269
rect 2562 3180 2596 3184
rect 2562 3074 2596 3078
rect 2562 2989 2596 3010
rect 2658 3248 2692 3269
rect 2658 3180 2692 3184
rect 2658 3074 2692 3078
rect 2658 2989 2692 3010
rect 2754 3248 2788 3269
rect 2754 3180 2788 3184
rect 2754 3074 2788 3078
rect 2754 2989 2788 3010
rect 2850 3248 2884 3269
rect 2850 3180 2884 3184
rect 2850 3074 2884 3078
rect 2850 2989 2884 3010
rect 2946 3248 2980 3269
rect 2946 3180 2980 3184
rect 2946 3074 2980 3078
rect 2946 2989 2980 3010
rect 3042 3248 3076 3269
rect 3042 3180 3076 3184
rect 3042 3074 3076 3078
rect 3042 2989 3076 3010
rect 3138 3248 3172 3269
rect 3138 3180 3172 3184
rect 3138 3074 3172 3078
rect 3138 2989 3172 3010
rect 3234 3248 3268 3269
rect 3234 3180 3268 3184
rect 3234 3074 3268 3078
rect 3234 2989 3268 3010
rect 3330 3248 3364 3269
rect 3330 3180 3364 3184
rect 3330 3074 3364 3078
rect 3330 2989 3364 3010
rect 3426 3248 3460 3269
rect 3426 3180 3460 3184
rect 3426 3074 3460 3078
rect 3426 2989 3460 3010
rect 3540 3211 3574 3215
rect 3540 3105 3574 3109
rect 3540 3033 3574 3041
rect 2352 2905 2386 2973
rect 3540 2905 3574 2973
rect 2352 2871 2470 2905
rect 2504 2871 2538 2905
rect 2572 2871 2606 2905
rect 2640 2871 2674 2905
rect 2708 2871 2742 2905
rect 2776 2871 2810 2905
rect 2844 2871 2878 2905
rect 2912 2871 2946 2905
rect 2980 2871 3014 2905
rect 3048 2871 3082 2905
rect 3116 2871 3150 2905
rect 3184 2871 3218 2905
rect 3252 2871 3286 2905
rect 3320 2871 3354 2905
rect 3388 2871 3422 2905
rect 3456 2871 3574 2905
rect 3873 3415 3991 3449
rect 4025 3415 4059 3449
rect 4093 3415 4127 3449
rect 4161 3415 4195 3449
rect 4229 3415 4263 3449
rect 4297 3415 4331 3449
rect 4365 3415 4399 3449
rect 4433 3415 4467 3449
rect 4501 3415 4535 3449
rect 4569 3415 4603 3449
rect 4637 3415 4671 3449
rect 4705 3415 4739 3449
rect 4773 3415 4807 3449
rect 4841 3415 4875 3449
rect 4909 3415 4943 3449
rect 4977 3415 5095 3449
rect 3873 3347 3907 3415
rect 5061 3347 5095 3415
rect 3971 3313 3987 3347
rect 4021 3313 4037 3347
rect 4163 3313 4179 3347
rect 4213 3313 4229 3347
rect 4355 3313 4371 3347
rect 4405 3313 4421 3347
rect 4547 3313 4563 3347
rect 4597 3313 4613 3347
rect 4739 3313 4755 3347
rect 4789 3313 4805 3347
rect 4931 3313 4947 3347
rect 4981 3313 4997 3347
rect 3873 3279 3907 3313
rect 5061 3279 5095 3287
rect 3873 3211 3907 3245
rect 3873 3143 3907 3177
rect 3873 3075 3907 3109
rect 3873 3007 3907 3041
rect 3987 3248 4021 3269
rect 3987 3180 4021 3184
rect 3987 3074 4021 3078
rect 3987 2989 4021 3010
rect 4083 3248 4117 3269
rect 4083 3180 4117 3184
rect 4083 3074 4117 3078
rect 4083 2989 4117 3010
rect 4179 3248 4213 3269
rect 4179 3180 4213 3184
rect 4179 3074 4213 3078
rect 4179 2989 4213 3010
rect 4275 3248 4309 3269
rect 4275 3180 4309 3184
rect 4275 3074 4309 3078
rect 4275 2989 4309 3010
rect 4371 3248 4405 3269
rect 4371 3180 4405 3184
rect 4371 3074 4405 3078
rect 4371 2989 4405 3010
rect 4467 3248 4501 3269
rect 4467 3180 4501 3184
rect 4467 3074 4501 3078
rect 4467 2989 4501 3010
rect 4563 3248 4597 3269
rect 4563 3180 4597 3184
rect 4563 3074 4597 3078
rect 4563 2989 4597 3010
rect 4659 3248 4693 3269
rect 4659 3180 4693 3184
rect 4659 3074 4693 3078
rect 4659 2989 4693 3010
rect 4755 3248 4789 3269
rect 4755 3180 4789 3184
rect 4755 3074 4789 3078
rect 4755 2989 4789 3010
rect 4851 3248 4885 3269
rect 4851 3180 4885 3184
rect 4851 3074 4885 3078
rect 4851 2989 4885 3010
rect 4947 3248 4981 3269
rect 4947 3180 4981 3184
rect 4947 3074 4981 3078
rect 4947 2989 4981 3010
rect 5061 3211 5095 3215
rect 5061 3105 5095 3109
rect 5274 3082 5303 3116
rect 5337 3082 5395 3116
rect 5429 3082 5487 3116
rect 5521 3082 5550 3116
rect 5061 3033 5095 3041
rect 3873 2905 3907 2973
rect 5061 2905 5095 2973
rect 3873 2871 3991 2905
rect 4025 2871 4059 2905
rect 4093 2871 4127 2905
rect 4161 2871 4195 2905
rect 4229 2871 4263 2905
rect 4297 2871 4331 2905
rect 4365 2871 4399 2905
rect 4433 2871 4467 2905
rect 4501 2871 4535 2905
rect 4569 2871 4603 2905
rect 4637 2871 4671 2905
rect 4705 2871 4739 2905
rect 4773 2871 4807 2905
rect 4841 2871 4875 2905
rect 4909 2871 4943 2905
rect 4977 2871 5095 2905
rect 5340 3040 5406 3048
rect 5340 3006 5356 3040
rect 5390 3006 5406 3040
rect 5340 2972 5406 3006
rect 5340 2938 5356 2972
rect 5390 2938 5406 2972
rect 5340 2904 5406 2938
rect 5340 2870 5356 2904
rect 5390 2870 5406 2904
rect 5340 2852 5406 2870
rect 5440 3040 5482 3082
rect 5474 3006 5482 3040
rect 5440 2972 5482 3006
rect 5474 2938 5482 2972
rect 5440 2904 5482 2938
rect 5474 2870 5482 2904
rect 5440 2854 5482 2870
rect 5340 2802 5386 2852
rect 199 2759 317 2793
rect 351 2759 385 2793
rect 419 2759 453 2793
rect 487 2759 521 2793
rect 555 2759 589 2793
rect 623 2759 657 2793
rect 691 2759 725 2793
rect 759 2759 793 2793
rect 827 2759 861 2793
rect 895 2759 929 2793
rect 963 2759 997 2793
rect 1031 2759 1065 2793
rect 1099 2759 1133 2793
rect 1167 2759 1201 2793
rect 1235 2759 1269 2793
rect 1303 2759 1421 2793
rect 199 2683 233 2759
rect 1387 2688 1421 2759
rect 199 2615 233 2649
rect 199 2547 233 2581
rect 313 2646 347 2685
rect 313 2573 347 2612
rect 409 2646 443 2685
rect 409 2573 443 2612
rect 505 2646 539 2685
rect 505 2573 539 2612
rect 601 2646 635 2685
rect 601 2573 635 2612
rect 697 2646 731 2685
rect 697 2573 731 2612
rect 793 2646 827 2685
rect 793 2573 827 2612
rect 889 2646 923 2685
rect 889 2573 923 2612
rect 985 2646 1019 2685
rect 985 2573 1019 2612
rect 1081 2646 1115 2685
rect 1081 2573 1115 2612
rect 1177 2646 1211 2685
rect 1177 2573 1211 2612
rect 1273 2646 1307 2685
rect 1273 2573 1307 2612
rect 1387 2616 1421 2649
rect 1387 2547 1421 2581
rect 199 2437 233 2513
rect 297 2501 313 2535
rect 347 2501 363 2535
rect 489 2501 505 2535
rect 539 2501 555 2535
rect 681 2501 697 2535
rect 731 2501 747 2535
rect 873 2501 889 2535
rect 923 2501 939 2535
rect 1065 2501 1081 2535
rect 1115 2501 1131 2535
rect 1257 2501 1273 2535
rect 1307 2501 1323 2535
rect 1387 2437 1421 2510
rect 199 2403 317 2437
rect 351 2403 385 2437
rect 419 2403 453 2437
rect 487 2403 521 2437
rect 555 2403 589 2437
rect 623 2403 657 2437
rect 691 2403 725 2437
rect 759 2403 793 2437
rect 827 2403 861 2437
rect 895 2403 929 2437
rect 963 2403 997 2437
rect 1031 2403 1065 2437
rect 1099 2403 1133 2437
rect 1167 2403 1201 2437
rect 1235 2403 1269 2437
rect 1303 2403 1421 2437
rect 2352 2763 2470 2797
rect 2504 2763 2538 2797
rect 2572 2763 2606 2797
rect 2640 2763 2674 2797
rect 2708 2763 2742 2797
rect 2776 2763 2810 2797
rect 2844 2763 2878 2797
rect 2912 2763 2946 2797
rect 2980 2763 3014 2797
rect 3048 2763 3082 2797
rect 3116 2763 3150 2797
rect 3184 2763 3218 2797
rect 3252 2763 3286 2797
rect 3320 2763 3354 2797
rect 3388 2763 3422 2797
rect 3456 2763 3574 2797
rect 2352 2687 2386 2763
rect 3540 2692 3574 2763
rect 3873 2763 3991 2797
rect 4025 2763 4059 2797
rect 4093 2763 4127 2797
rect 4161 2763 4195 2797
rect 4229 2763 4263 2797
rect 4297 2763 4331 2797
rect 4365 2763 4399 2797
rect 4433 2763 4467 2797
rect 4501 2763 4535 2797
rect 4569 2763 4603 2797
rect 4637 2763 4671 2797
rect 4705 2763 4739 2797
rect 4773 2763 4807 2797
rect 4841 2763 4875 2797
rect 4909 2763 4943 2797
rect 4977 2763 5095 2797
rect 3675 2727 3691 2761
rect 3725 2727 3741 2761
rect 2352 2619 2386 2653
rect 2352 2551 2386 2585
rect 2466 2650 2500 2689
rect 2466 2577 2500 2616
rect 2562 2650 2596 2689
rect 2562 2577 2596 2616
rect 2658 2650 2692 2689
rect 2658 2577 2692 2616
rect 2754 2650 2788 2689
rect 2754 2577 2788 2616
rect 2850 2650 2884 2689
rect 2850 2577 2884 2616
rect 2946 2650 2980 2689
rect 2946 2577 2980 2616
rect 3042 2650 3076 2689
rect 3042 2577 3076 2616
rect 3138 2650 3172 2689
rect 3138 2577 3172 2616
rect 3234 2650 3268 2689
rect 3234 2577 3268 2616
rect 3330 2650 3364 2689
rect 3330 2577 3364 2616
rect 3426 2650 3460 2689
rect 3426 2577 3460 2616
rect 3540 2620 3574 2653
rect 3647 2677 3681 2693
rect 3647 2585 3681 2601
rect 3735 2677 3769 2693
rect 3735 2585 3769 2601
rect 3873 2687 3907 2763
rect 5061 2692 5095 2763
rect 3873 2619 3907 2653
rect 3540 2551 3574 2585
rect 2352 2441 2386 2517
rect 2450 2505 2466 2539
rect 2500 2505 2516 2539
rect 2642 2505 2658 2539
rect 2692 2505 2708 2539
rect 2834 2505 2850 2539
rect 2884 2505 2900 2539
rect 3026 2505 3042 2539
rect 3076 2505 3092 2539
rect 3218 2505 3234 2539
rect 3268 2505 3284 2539
rect 3410 2505 3426 2539
rect 3460 2505 3476 2539
rect 3540 2441 3574 2514
rect 2352 2407 2470 2441
rect 2504 2407 2538 2441
rect 2572 2407 2606 2441
rect 2640 2407 2674 2441
rect 2708 2407 2742 2441
rect 2776 2407 2810 2441
rect 2844 2407 2878 2441
rect 2912 2407 2946 2441
rect 2980 2407 3014 2441
rect 3048 2407 3082 2441
rect 3116 2407 3150 2441
rect 3184 2407 3218 2441
rect 3252 2407 3286 2441
rect 3320 2407 3354 2441
rect 3388 2407 3422 2441
rect 3456 2407 3574 2441
rect 3873 2551 3907 2585
rect 3987 2650 4021 2689
rect 3987 2577 4021 2616
rect 4083 2650 4117 2689
rect 4083 2577 4117 2616
rect 4179 2650 4213 2689
rect 4179 2577 4213 2616
rect 4275 2650 4309 2689
rect 4275 2577 4309 2616
rect 4371 2650 4405 2689
rect 4371 2577 4405 2616
rect 4467 2650 4501 2689
rect 4467 2577 4501 2616
rect 4563 2650 4597 2689
rect 4563 2577 4597 2616
rect 4659 2650 4693 2689
rect 4659 2577 4693 2616
rect 4755 2650 4789 2689
rect 4755 2577 4789 2616
rect 4851 2650 4885 2689
rect 4851 2577 4885 2616
rect 4947 2650 4981 2689
rect 4947 2577 4981 2616
rect 5061 2620 5095 2653
rect 5340 2768 5348 2802
rect 5382 2768 5386 2802
rect 5420 2807 5486 2818
rect 5420 2804 5450 2807
rect 5420 2770 5436 2804
rect 5484 2773 5486 2807
rect 5470 2770 5486 2773
rect 5340 2732 5386 2768
rect 5340 2720 5406 2732
rect 5340 2686 5356 2720
rect 5390 2686 5406 2720
rect 5340 2652 5406 2686
rect 5340 2618 5356 2652
rect 5390 2618 5406 2652
rect 5340 2606 5406 2618
rect 5440 2720 5486 2736
rect 5474 2686 5486 2720
rect 5440 2652 5486 2686
rect 5474 2618 5486 2652
rect 5061 2551 5095 2585
rect 5440 2572 5486 2618
rect 3873 2441 3907 2517
rect 3971 2505 3987 2539
rect 4021 2505 4037 2539
rect 4163 2505 4179 2539
rect 4213 2505 4229 2539
rect 4355 2505 4371 2539
rect 4405 2505 4421 2539
rect 4547 2505 4563 2539
rect 4597 2505 4613 2539
rect 4739 2505 4755 2539
rect 4789 2505 4805 2539
rect 4931 2505 4947 2539
rect 4981 2505 4997 2539
rect 5274 2538 5303 2572
rect 5337 2538 5395 2572
rect 5429 2538 5487 2572
rect 5521 2538 5550 2572
rect 5061 2441 5095 2514
rect 3873 2407 3991 2441
rect 4025 2407 4059 2441
rect 4093 2407 4127 2441
rect 4161 2407 4195 2441
rect 4229 2407 4263 2441
rect 4297 2407 4331 2441
rect 4365 2407 4399 2441
rect 4433 2407 4467 2441
rect 4501 2407 4535 2441
rect 4569 2407 4603 2441
rect 4637 2407 4671 2441
rect 4705 2407 4739 2441
rect 4773 2407 4807 2441
rect 4841 2407 4875 2441
rect 4909 2407 4943 2441
rect 4977 2407 5095 2441
rect 199 2124 317 2158
rect 351 2124 385 2158
rect 419 2124 453 2158
rect 487 2124 521 2158
rect 555 2124 589 2158
rect 623 2124 657 2158
rect 691 2124 725 2158
rect 759 2124 793 2158
rect 827 2124 861 2158
rect 895 2124 929 2158
rect 963 2124 997 2158
rect 1031 2124 1065 2158
rect 1099 2124 1133 2158
rect 1167 2124 1201 2158
rect 1235 2124 1269 2158
rect 1303 2124 1421 2158
rect 199 2056 233 2124
rect 1387 2056 1421 2124
rect 297 2022 313 2056
rect 347 2022 363 2056
rect 489 2022 505 2056
rect 539 2022 555 2056
rect 681 2022 697 2056
rect 731 2022 747 2056
rect 873 2022 889 2056
rect 923 2022 939 2056
rect 1065 2022 1081 2056
rect 1115 2022 1131 2056
rect 1257 2022 1273 2056
rect 1307 2022 1323 2056
rect 199 1988 233 2022
rect 1387 1988 1421 1996
rect 199 1920 233 1954
rect 199 1852 233 1886
rect 199 1784 233 1818
rect 199 1716 233 1750
rect 313 1957 347 1978
rect 313 1889 347 1893
rect 313 1783 347 1787
rect 313 1698 347 1719
rect 409 1957 443 1978
rect 409 1889 443 1893
rect 409 1783 443 1787
rect 409 1698 443 1719
rect 505 1957 539 1978
rect 505 1889 539 1893
rect 505 1783 539 1787
rect 505 1698 539 1719
rect 601 1957 635 1978
rect 601 1889 635 1893
rect 601 1783 635 1787
rect 601 1698 635 1719
rect 697 1957 731 1978
rect 697 1889 731 1893
rect 697 1783 731 1787
rect 697 1698 731 1719
rect 793 1957 827 1978
rect 793 1889 827 1893
rect 793 1783 827 1787
rect 793 1698 827 1719
rect 889 1957 923 1978
rect 889 1889 923 1893
rect 889 1783 923 1787
rect 889 1698 923 1719
rect 985 1957 1019 1978
rect 985 1889 1019 1893
rect 985 1783 1019 1787
rect 985 1698 1019 1719
rect 1081 1957 1115 1978
rect 1081 1889 1115 1893
rect 1081 1783 1115 1787
rect 1081 1698 1115 1719
rect 1177 1957 1211 1978
rect 1177 1889 1211 1893
rect 1177 1783 1211 1787
rect 1177 1698 1211 1719
rect 1273 1957 1307 1978
rect 1273 1889 1307 1893
rect 1273 1783 1307 1787
rect 1273 1698 1307 1719
rect 1387 1920 1421 1924
rect 1387 1814 1421 1818
rect 1387 1742 1421 1750
rect 199 1614 233 1682
rect 1387 1614 1421 1682
rect 199 1580 317 1614
rect 351 1580 385 1614
rect 419 1580 453 1614
rect 487 1580 521 1614
rect 555 1580 589 1614
rect 623 1580 657 1614
rect 691 1580 725 1614
rect 759 1580 793 1614
rect 827 1580 861 1614
rect 895 1580 929 1614
rect 963 1580 997 1614
rect 1031 1580 1065 1614
rect 1099 1580 1133 1614
rect 1167 1580 1201 1614
rect 1235 1580 1269 1614
rect 1303 1580 1421 1614
rect 2352 2128 2470 2162
rect 2504 2128 2538 2162
rect 2572 2128 2606 2162
rect 2640 2128 2674 2162
rect 2708 2128 2742 2162
rect 2776 2128 2810 2162
rect 2844 2128 2878 2162
rect 2912 2128 2946 2162
rect 2980 2128 3014 2162
rect 3048 2128 3082 2162
rect 3116 2128 3150 2162
rect 3184 2128 3218 2162
rect 3252 2128 3286 2162
rect 3320 2128 3354 2162
rect 3388 2128 3422 2162
rect 3456 2128 3574 2162
rect 2352 2060 2386 2128
rect 3540 2060 3574 2128
rect 2450 2026 2466 2060
rect 2500 2026 2516 2060
rect 2642 2026 2658 2060
rect 2692 2026 2708 2060
rect 2834 2026 2850 2060
rect 2884 2026 2900 2060
rect 3026 2026 3042 2060
rect 3076 2026 3092 2060
rect 3218 2026 3234 2060
rect 3268 2026 3284 2060
rect 3410 2026 3426 2060
rect 3460 2026 3476 2060
rect 2352 1992 2386 2026
rect 3540 1992 3574 2000
rect 2352 1924 2386 1958
rect 2352 1856 2386 1890
rect 2352 1788 2386 1822
rect 2352 1720 2386 1754
rect 2466 1961 2500 1982
rect 2466 1893 2500 1897
rect 2466 1787 2500 1791
rect 2466 1702 2500 1723
rect 2562 1961 2596 1982
rect 2562 1893 2596 1897
rect 2562 1787 2596 1791
rect 2562 1702 2596 1723
rect 2658 1961 2692 1982
rect 2658 1893 2692 1897
rect 2658 1787 2692 1791
rect 2658 1702 2692 1723
rect 2754 1961 2788 1982
rect 2754 1893 2788 1897
rect 2754 1787 2788 1791
rect 2754 1702 2788 1723
rect 2850 1961 2884 1982
rect 2850 1893 2884 1897
rect 2850 1787 2884 1791
rect 2850 1702 2884 1723
rect 2946 1961 2980 1982
rect 2946 1893 2980 1897
rect 2946 1787 2980 1791
rect 2946 1702 2980 1723
rect 3042 1961 3076 1982
rect 3042 1893 3076 1897
rect 3042 1787 3076 1791
rect 3042 1702 3076 1723
rect 3138 1961 3172 1982
rect 3138 1893 3172 1897
rect 3138 1787 3172 1791
rect 3138 1702 3172 1723
rect 3234 1961 3268 1982
rect 3234 1893 3268 1897
rect 3234 1787 3268 1791
rect 3234 1702 3268 1723
rect 3330 1961 3364 1982
rect 3330 1893 3364 1897
rect 3330 1787 3364 1791
rect 3330 1702 3364 1723
rect 3426 1961 3460 1982
rect 3426 1893 3460 1897
rect 3426 1787 3460 1791
rect 3426 1702 3460 1723
rect 3540 1924 3574 1928
rect 3540 1818 3574 1822
rect 3540 1746 3574 1754
rect 2352 1618 2386 1686
rect 3540 1618 3574 1686
rect 2352 1584 2470 1618
rect 2504 1584 2538 1618
rect 2572 1584 2606 1618
rect 2640 1584 2674 1618
rect 2708 1584 2742 1618
rect 2776 1584 2810 1618
rect 2844 1584 2878 1618
rect 2912 1584 2946 1618
rect 2980 1584 3014 1618
rect 3048 1584 3082 1618
rect 3116 1584 3150 1618
rect 3184 1584 3218 1618
rect 3252 1584 3286 1618
rect 3320 1584 3354 1618
rect 3388 1584 3422 1618
rect 3456 1584 3574 1618
rect 3873 2128 3991 2162
rect 4025 2128 4059 2162
rect 4093 2128 4127 2162
rect 4161 2128 4195 2162
rect 4229 2128 4263 2162
rect 4297 2128 4331 2162
rect 4365 2128 4399 2162
rect 4433 2128 4467 2162
rect 4501 2128 4535 2162
rect 4569 2128 4603 2162
rect 4637 2128 4671 2162
rect 4705 2128 4739 2162
rect 4773 2128 4807 2162
rect 4841 2128 4875 2162
rect 4909 2128 4943 2162
rect 4977 2128 5095 2162
rect 3873 2060 3907 2128
rect 5061 2060 5095 2128
rect 3971 2026 3987 2060
rect 4021 2026 4037 2060
rect 4163 2026 4179 2060
rect 4213 2026 4229 2060
rect 4355 2026 4371 2060
rect 4405 2026 4421 2060
rect 4547 2026 4563 2060
rect 4597 2026 4613 2060
rect 4739 2026 4755 2060
rect 4789 2026 4805 2060
rect 4931 2026 4947 2060
rect 4981 2026 4997 2060
rect 3873 1992 3907 2026
rect 5061 1992 5095 2000
rect 3873 1924 3907 1958
rect 3873 1856 3907 1890
rect 3873 1788 3907 1822
rect 3873 1720 3907 1754
rect 3987 1961 4021 1982
rect 3987 1893 4021 1897
rect 3987 1787 4021 1791
rect 3987 1702 4021 1723
rect 4083 1961 4117 1982
rect 4083 1893 4117 1897
rect 4083 1787 4117 1791
rect 4083 1702 4117 1723
rect 4179 1961 4213 1982
rect 4179 1893 4213 1897
rect 4179 1787 4213 1791
rect 4179 1702 4213 1723
rect 4275 1961 4309 1982
rect 4275 1893 4309 1897
rect 4275 1787 4309 1791
rect 4275 1702 4309 1723
rect 4371 1961 4405 1982
rect 4371 1893 4405 1897
rect 4371 1787 4405 1791
rect 4371 1702 4405 1723
rect 4467 1961 4501 1982
rect 4467 1893 4501 1897
rect 4467 1787 4501 1791
rect 4467 1702 4501 1723
rect 4563 1961 4597 1982
rect 4563 1893 4597 1897
rect 4563 1787 4597 1791
rect 4563 1702 4597 1723
rect 4659 1961 4693 1982
rect 4659 1893 4693 1897
rect 4659 1787 4693 1791
rect 4659 1702 4693 1723
rect 4755 1961 4789 1982
rect 4755 1893 4789 1897
rect 4755 1787 4789 1791
rect 4755 1702 4789 1723
rect 4851 1961 4885 1982
rect 4851 1893 4885 1897
rect 4851 1787 4885 1791
rect 4851 1702 4885 1723
rect 4947 1961 4981 1982
rect 4947 1893 4981 1897
rect 4947 1787 4981 1791
rect 4947 1702 4981 1723
rect 5061 1924 5095 1928
rect 5061 1818 5095 1822
rect 5274 1795 5303 1829
rect 5337 1795 5395 1829
rect 5429 1795 5487 1829
rect 5521 1795 5550 1829
rect 5061 1746 5095 1754
rect 3873 1618 3907 1686
rect 5061 1618 5095 1686
rect 3873 1584 3991 1618
rect 4025 1584 4059 1618
rect 4093 1584 4127 1618
rect 4161 1584 4195 1618
rect 4229 1584 4263 1618
rect 4297 1584 4331 1618
rect 4365 1584 4399 1618
rect 4433 1584 4467 1618
rect 4501 1584 4535 1618
rect 4569 1584 4603 1618
rect 4637 1584 4671 1618
rect 4705 1584 4739 1618
rect 4773 1584 4807 1618
rect 4841 1584 4875 1618
rect 4909 1584 4943 1618
rect 4977 1584 5095 1618
rect 5340 1753 5406 1761
rect 5340 1719 5356 1753
rect 5390 1719 5406 1753
rect 5340 1685 5406 1719
rect 5340 1651 5356 1685
rect 5390 1651 5406 1685
rect 5340 1617 5406 1651
rect 5340 1583 5356 1617
rect 5390 1583 5406 1617
rect 5340 1565 5406 1583
rect 5440 1753 5482 1795
rect 5474 1719 5482 1753
rect 5440 1685 5482 1719
rect 5474 1651 5482 1685
rect 5440 1617 5482 1651
rect 5474 1583 5482 1617
rect 5440 1567 5482 1583
rect 5340 1515 5386 1565
rect 199 1472 317 1506
rect 351 1472 385 1506
rect 419 1472 453 1506
rect 487 1472 521 1506
rect 555 1472 589 1506
rect 623 1472 657 1506
rect 691 1472 725 1506
rect 759 1472 793 1506
rect 827 1472 861 1506
rect 895 1472 929 1506
rect 963 1472 997 1506
rect 1031 1472 1065 1506
rect 1099 1472 1133 1506
rect 1167 1472 1201 1506
rect 1235 1472 1269 1506
rect 1303 1472 1421 1506
rect 199 1396 233 1472
rect 1387 1401 1421 1472
rect 199 1328 233 1362
rect 199 1260 233 1294
rect 313 1359 347 1398
rect 313 1286 347 1325
rect 409 1359 443 1398
rect 409 1286 443 1325
rect 505 1359 539 1398
rect 505 1286 539 1325
rect 601 1359 635 1398
rect 601 1286 635 1325
rect 697 1359 731 1398
rect 697 1286 731 1325
rect 793 1359 827 1398
rect 793 1286 827 1325
rect 889 1359 923 1398
rect 889 1286 923 1325
rect 985 1359 1019 1398
rect 985 1286 1019 1325
rect 1081 1359 1115 1398
rect 1081 1286 1115 1325
rect 1177 1359 1211 1398
rect 1177 1286 1211 1325
rect 1273 1359 1307 1398
rect 1273 1286 1307 1325
rect 1387 1329 1421 1362
rect 1387 1260 1421 1294
rect 199 1150 233 1226
rect 297 1214 313 1248
rect 347 1214 363 1248
rect 489 1214 505 1248
rect 539 1214 555 1248
rect 681 1214 697 1248
rect 731 1214 747 1248
rect 873 1214 889 1248
rect 923 1214 939 1248
rect 1065 1214 1081 1248
rect 1115 1214 1131 1248
rect 1257 1214 1273 1248
rect 1307 1214 1323 1248
rect 1387 1150 1421 1223
rect 199 1116 317 1150
rect 351 1116 385 1150
rect 419 1116 453 1150
rect 487 1116 521 1150
rect 555 1116 589 1150
rect 623 1116 657 1150
rect 691 1116 725 1150
rect 759 1116 793 1150
rect 827 1116 861 1150
rect 895 1116 929 1150
rect 963 1116 997 1150
rect 1031 1116 1065 1150
rect 1099 1116 1133 1150
rect 1167 1116 1201 1150
rect 1235 1116 1269 1150
rect 1303 1116 1421 1150
rect 2352 1476 2470 1510
rect 2504 1476 2538 1510
rect 2572 1476 2606 1510
rect 2640 1476 2674 1510
rect 2708 1476 2742 1510
rect 2776 1476 2810 1510
rect 2844 1476 2878 1510
rect 2912 1476 2946 1510
rect 2980 1476 3014 1510
rect 3048 1476 3082 1510
rect 3116 1476 3150 1510
rect 3184 1476 3218 1510
rect 3252 1476 3286 1510
rect 3320 1476 3354 1510
rect 3388 1476 3422 1510
rect 3456 1476 3574 1510
rect 2352 1400 2386 1476
rect 3540 1405 3574 1476
rect 3873 1476 3991 1510
rect 4025 1476 4059 1510
rect 4093 1476 4127 1510
rect 4161 1476 4195 1510
rect 4229 1476 4263 1510
rect 4297 1476 4331 1510
rect 4365 1476 4399 1510
rect 4433 1476 4467 1510
rect 4501 1476 4535 1510
rect 4569 1476 4603 1510
rect 4637 1476 4671 1510
rect 4705 1476 4739 1510
rect 4773 1476 4807 1510
rect 4841 1476 4875 1510
rect 4909 1476 4943 1510
rect 4977 1476 5095 1510
rect 3675 1440 3691 1474
rect 3725 1440 3741 1474
rect 2352 1332 2386 1366
rect 2352 1264 2386 1298
rect 2466 1363 2500 1402
rect 2466 1290 2500 1329
rect 2562 1363 2596 1402
rect 2562 1290 2596 1329
rect 2658 1363 2692 1402
rect 2658 1290 2692 1329
rect 2754 1363 2788 1402
rect 2754 1290 2788 1329
rect 2850 1363 2884 1402
rect 2850 1290 2884 1329
rect 2946 1363 2980 1402
rect 2946 1290 2980 1329
rect 3042 1363 3076 1402
rect 3042 1290 3076 1329
rect 3138 1363 3172 1402
rect 3138 1290 3172 1329
rect 3234 1363 3268 1402
rect 3234 1290 3268 1329
rect 3330 1363 3364 1402
rect 3330 1290 3364 1329
rect 3426 1363 3460 1402
rect 3426 1290 3460 1329
rect 3540 1333 3574 1366
rect 3647 1390 3681 1406
rect 3647 1298 3681 1314
rect 3735 1390 3769 1406
rect 3735 1298 3769 1314
rect 3873 1400 3907 1476
rect 5061 1405 5095 1476
rect 3873 1332 3907 1366
rect 3540 1264 3574 1298
rect 2352 1154 2386 1230
rect 2450 1218 2466 1252
rect 2500 1218 2516 1252
rect 2642 1218 2658 1252
rect 2692 1218 2708 1252
rect 2834 1218 2850 1252
rect 2884 1218 2900 1252
rect 3026 1218 3042 1252
rect 3076 1218 3092 1252
rect 3218 1218 3234 1252
rect 3268 1218 3284 1252
rect 3410 1218 3426 1252
rect 3460 1218 3476 1252
rect 3540 1154 3574 1227
rect 2352 1120 2470 1154
rect 2504 1120 2538 1154
rect 2572 1120 2606 1154
rect 2640 1120 2674 1154
rect 2708 1120 2742 1154
rect 2776 1120 2810 1154
rect 2844 1120 2878 1154
rect 2912 1120 2946 1154
rect 2980 1120 3014 1154
rect 3048 1120 3082 1154
rect 3116 1120 3150 1154
rect 3184 1120 3218 1154
rect 3252 1120 3286 1154
rect 3320 1120 3354 1154
rect 3388 1120 3422 1154
rect 3456 1120 3574 1154
rect 3873 1264 3907 1298
rect 3987 1363 4021 1402
rect 3987 1290 4021 1329
rect 4083 1363 4117 1402
rect 4083 1290 4117 1329
rect 4179 1363 4213 1402
rect 4179 1290 4213 1329
rect 4275 1363 4309 1402
rect 4275 1290 4309 1329
rect 4371 1363 4405 1402
rect 4371 1290 4405 1329
rect 4467 1363 4501 1402
rect 4467 1290 4501 1329
rect 4563 1363 4597 1402
rect 4563 1290 4597 1329
rect 4659 1363 4693 1402
rect 4659 1290 4693 1329
rect 4755 1363 4789 1402
rect 4755 1290 4789 1329
rect 4851 1363 4885 1402
rect 4851 1290 4885 1329
rect 4947 1363 4981 1402
rect 4947 1290 4981 1329
rect 5061 1333 5095 1366
rect 5340 1481 5348 1515
rect 5382 1481 5386 1515
rect 5420 1520 5486 1531
rect 5420 1517 5450 1520
rect 5420 1483 5436 1517
rect 5484 1486 5486 1520
rect 5470 1483 5486 1486
rect 5340 1445 5386 1481
rect 5340 1433 5406 1445
rect 5340 1399 5356 1433
rect 5390 1399 5406 1433
rect 5340 1365 5406 1399
rect 5340 1331 5356 1365
rect 5390 1331 5406 1365
rect 5340 1319 5406 1331
rect 5440 1433 5486 1449
rect 5474 1399 5486 1433
rect 5440 1365 5486 1399
rect 5474 1331 5486 1365
rect 5061 1264 5095 1298
rect 5440 1285 5486 1331
rect 3873 1154 3907 1230
rect 3971 1218 3987 1252
rect 4021 1218 4037 1252
rect 4163 1218 4179 1252
rect 4213 1218 4229 1252
rect 4355 1218 4371 1252
rect 4405 1218 4421 1252
rect 4547 1218 4563 1252
rect 4597 1218 4613 1252
rect 4739 1218 4755 1252
rect 4789 1218 4805 1252
rect 4931 1218 4947 1252
rect 4981 1218 4997 1252
rect 5274 1251 5303 1285
rect 5337 1251 5395 1285
rect 5429 1251 5487 1285
rect 5521 1251 5550 1285
rect 5061 1154 5095 1227
rect 3873 1120 3991 1154
rect 4025 1120 4059 1154
rect 4093 1120 4127 1154
rect 4161 1120 4195 1154
rect 4229 1120 4263 1154
rect 4297 1120 4331 1154
rect 4365 1120 4399 1154
rect 4433 1120 4467 1154
rect 4501 1120 4535 1154
rect 4569 1120 4603 1154
rect 4637 1120 4671 1154
rect 4705 1120 4739 1154
rect 4773 1120 4807 1154
rect 4841 1120 4875 1154
rect 4909 1120 4943 1154
rect 4977 1120 5095 1154
<< viali >>
rect 313 41919 347 41953
rect 505 41919 539 41953
rect 697 41919 731 41953
rect 889 41919 923 41953
rect 1081 41919 1115 41953
rect 1273 41919 1307 41953
rect 1387 41919 1421 41927
rect 1387 41893 1421 41919
rect 313 41820 347 41824
rect 313 41790 347 41820
rect 313 41718 347 41752
rect 313 41650 347 41680
rect 313 41646 347 41650
rect 409 41820 443 41824
rect 409 41790 443 41820
rect 409 41718 443 41752
rect 409 41650 443 41680
rect 409 41646 443 41650
rect 505 41820 539 41824
rect 505 41790 539 41820
rect 505 41718 539 41752
rect 505 41650 539 41680
rect 505 41646 539 41650
rect 601 41820 635 41824
rect 601 41790 635 41820
rect 601 41718 635 41752
rect 601 41650 635 41680
rect 601 41646 635 41650
rect 697 41820 731 41824
rect 697 41790 731 41820
rect 697 41718 731 41752
rect 697 41650 731 41680
rect 697 41646 731 41650
rect 793 41820 827 41824
rect 793 41790 827 41820
rect 793 41718 827 41752
rect 793 41650 827 41680
rect 793 41646 827 41650
rect 889 41820 923 41824
rect 889 41790 923 41820
rect 889 41718 923 41752
rect 889 41650 923 41680
rect 889 41646 923 41650
rect 985 41820 1019 41824
rect 985 41790 1019 41820
rect 985 41718 1019 41752
rect 985 41650 1019 41680
rect 985 41646 1019 41650
rect 1081 41820 1115 41824
rect 1081 41790 1115 41820
rect 1081 41718 1115 41752
rect 1081 41650 1115 41680
rect 1081 41646 1115 41650
rect 1177 41820 1211 41824
rect 1177 41790 1211 41820
rect 1177 41718 1211 41752
rect 1177 41650 1211 41680
rect 1177 41646 1211 41650
rect 1273 41820 1307 41824
rect 1273 41790 1307 41820
rect 1273 41718 1307 41752
rect 1273 41650 1307 41680
rect 1273 41646 1307 41650
rect 1387 41851 1421 41855
rect 1387 41821 1421 41851
rect 1387 41749 1421 41783
rect 1387 41681 1421 41711
rect 1387 41677 1421 41681
rect 1387 41613 1421 41639
rect 1387 41605 1421 41613
rect 2466 41923 2500 41957
rect 2658 41923 2692 41957
rect 2850 41923 2884 41957
rect 3042 41923 3076 41957
rect 3234 41923 3268 41957
rect 3426 41923 3460 41957
rect 3540 41923 3574 41931
rect 3540 41897 3574 41923
rect 2466 41824 2500 41828
rect 2466 41794 2500 41824
rect 2466 41722 2500 41756
rect 2466 41654 2500 41684
rect 2466 41650 2500 41654
rect 2562 41824 2596 41828
rect 2562 41794 2596 41824
rect 2562 41722 2596 41756
rect 2562 41654 2596 41684
rect 2562 41650 2596 41654
rect 2658 41824 2692 41828
rect 2658 41794 2692 41824
rect 2658 41722 2692 41756
rect 2658 41654 2692 41684
rect 2658 41650 2692 41654
rect 2754 41824 2788 41828
rect 2754 41794 2788 41824
rect 2754 41722 2788 41756
rect 2754 41654 2788 41684
rect 2754 41650 2788 41654
rect 2850 41824 2884 41828
rect 2850 41794 2884 41824
rect 2850 41722 2884 41756
rect 2850 41654 2884 41684
rect 2850 41650 2884 41654
rect 2946 41824 2980 41828
rect 2946 41794 2980 41824
rect 2946 41722 2980 41756
rect 2946 41654 2980 41684
rect 2946 41650 2980 41654
rect 3042 41824 3076 41828
rect 3042 41794 3076 41824
rect 3042 41722 3076 41756
rect 3042 41654 3076 41684
rect 3042 41650 3076 41654
rect 3138 41824 3172 41828
rect 3138 41794 3172 41824
rect 3138 41722 3172 41756
rect 3138 41654 3172 41684
rect 3138 41650 3172 41654
rect 3234 41824 3268 41828
rect 3234 41794 3268 41824
rect 3234 41722 3268 41756
rect 3234 41654 3268 41684
rect 3234 41650 3268 41654
rect 3330 41824 3364 41828
rect 3330 41794 3364 41824
rect 3330 41722 3364 41756
rect 3330 41654 3364 41684
rect 3330 41650 3364 41654
rect 3426 41824 3460 41828
rect 3426 41794 3460 41824
rect 3426 41722 3460 41756
rect 3426 41654 3460 41684
rect 3426 41650 3460 41654
rect 3540 41855 3574 41859
rect 3540 41825 3574 41855
rect 3540 41753 3574 41787
rect 3540 41685 3574 41715
rect 3540 41681 3574 41685
rect 3540 41617 3574 41643
rect 3540 41609 3574 41617
rect 3987 41923 4021 41957
rect 4179 41923 4213 41957
rect 4371 41923 4405 41957
rect 4563 41923 4597 41957
rect 4755 41923 4789 41957
rect 4947 41923 4981 41957
rect 5061 41923 5095 41931
rect 5061 41897 5095 41923
rect 3987 41824 4021 41828
rect 3987 41794 4021 41824
rect 3987 41722 4021 41756
rect 3987 41654 4021 41684
rect 3987 41650 4021 41654
rect 4083 41824 4117 41828
rect 4083 41794 4117 41824
rect 4083 41722 4117 41756
rect 4083 41654 4117 41684
rect 4083 41650 4117 41654
rect 4179 41824 4213 41828
rect 4179 41794 4213 41824
rect 4179 41722 4213 41756
rect 4179 41654 4213 41684
rect 4179 41650 4213 41654
rect 4275 41824 4309 41828
rect 4275 41794 4309 41824
rect 4275 41722 4309 41756
rect 4275 41654 4309 41684
rect 4275 41650 4309 41654
rect 4371 41824 4405 41828
rect 4371 41794 4405 41824
rect 4371 41722 4405 41756
rect 4371 41654 4405 41684
rect 4371 41650 4405 41654
rect 4467 41824 4501 41828
rect 4467 41794 4501 41824
rect 4467 41722 4501 41756
rect 4467 41654 4501 41684
rect 4467 41650 4501 41654
rect 4563 41824 4597 41828
rect 4563 41794 4597 41824
rect 4563 41722 4597 41756
rect 4563 41654 4597 41684
rect 4563 41650 4597 41654
rect 4659 41824 4693 41828
rect 4659 41794 4693 41824
rect 4659 41722 4693 41756
rect 4659 41654 4693 41684
rect 4659 41650 4693 41654
rect 4755 41824 4789 41828
rect 4755 41794 4789 41824
rect 4755 41722 4789 41756
rect 4755 41654 4789 41684
rect 4755 41650 4789 41654
rect 4851 41824 4885 41828
rect 4851 41794 4885 41824
rect 4851 41722 4885 41756
rect 4851 41654 4885 41684
rect 4851 41650 4885 41654
rect 4947 41824 4981 41828
rect 4947 41794 4981 41824
rect 4947 41722 4981 41756
rect 4947 41654 4981 41684
rect 4947 41650 4981 41654
rect 5061 41855 5095 41859
rect 5061 41825 5095 41855
rect 5061 41753 5095 41787
rect 5061 41685 5095 41715
rect 5303 41692 5337 41726
rect 5395 41692 5429 41726
rect 5487 41692 5521 41726
rect 5061 41681 5095 41685
rect 5061 41617 5095 41643
rect 5061 41609 5095 41617
rect 313 41222 347 41256
rect 409 41222 443 41256
rect 505 41222 539 41256
rect 601 41222 635 41256
rect 697 41222 731 41256
rect 793 41222 827 41256
rect 889 41222 923 41256
rect 985 41222 1019 41256
rect 1081 41222 1115 41256
rect 1177 41222 1211 41256
rect 1273 41222 1307 41256
rect 1387 41293 1421 41298
rect 1387 41264 1421 41293
rect 1387 41225 1421 41226
rect 1387 41192 1421 41225
rect 313 41111 347 41145
rect 505 41111 539 41145
rect 697 41111 731 41145
rect 889 41111 923 41145
rect 1081 41111 1115 41145
rect 1273 41111 1307 41145
rect 1387 41123 1421 41154
rect 1387 41120 1421 41123
rect 3691 41337 3725 41371
rect 2466 41226 2500 41260
rect 2562 41226 2596 41260
rect 2658 41226 2692 41260
rect 2754 41226 2788 41260
rect 2850 41226 2884 41260
rect 2946 41226 2980 41260
rect 3042 41226 3076 41260
rect 3138 41226 3172 41260
rect 3234 41226 3268 41260
rect 3330 41226 3364 41260
rect 3426 41226 3460 41260
rect 3540 41297 3574 41302
rect 3540 41268 3574 41297
rect 3540 41229 3574 41230
rect 3540 41196 3574 41229
rect 3647 41211 3681 41287
rect 3735 41211 3769 41287
rect 2466 41115 2500 41149
rect 2658 41115 2692 41149
rect 2850 41115 2884 41149
rect 3042 41115 3076 41149
rect 3234 41115 3268 41149
rect 3426 41115 3460 41149
rect 3540 41127 3574 41158
rect 3540 41124 3574 41127
rect 3987 41226 4021 41260
rect 4083 41226 4117 41260
rect 4179 41226 4213 41260
rect 4275 41226 4309 41260
rect 4371 41226 4405 41260
rect 4467 41226 4501 41260
rect 4563 41226 4597 41260
rect 4659 41226 4693 41260
rect 4755 41226 4789 41260
rect 4851 41226 4885 41260
rect 4947 41226 4981 41260
rect 5061 41297 5095 41302
rect 5061 41268 5095 41297
rect 5061 41229 5095 41230
rect 5061 41196 5095 41229
rect 5348 41378 5382 41412
rect 5450 41414 5484 41417
rect 5450 41383 5470 41414
rect 5470 41383 5484 41414
rect 3987 41115 4021 41149
rect 4179 41115 4213 41149
rect 4371 41115 4405 41149
rect 4563 41115 4597 41149
rect 4755 41115 4789 41149
rect 4947 41115 4981 41149
rect 5061 41127 5095 41158
rect 5303 41148 5337 41182
rect 5395 41148 5429 41182
rect 5487 41148 5521 41182
rect 5061 41124 5095 41127
rect 313 40632 347 40666
rect 505 40632 539 40666
rect 697 40632 731 40666
rect 889 40632 923 40666
rect 1081 40632 1115 40666
rect 1273 40632 1307 40666
rect 1387 40632 1421 40640
rect 1387 40606 1421 40632
rect 313 40533 347 40537
rect 313 40503 347 40533
rect 313 40431 347 40465
rect 313 40363 347 40393
rect 313 40359 347 40363
rect 409 40533 443 40537
rect 409 40503 443 40533
rect 409 40431 443 40465
rect 409 40363 443 40393
rect 409 40359 443 40363
rect 505 40533 539 40537
rect 505 40503 539 40533
rect 505 40431 539 40465
rect 505 40363 539 40393
rect 505 40359 539 40363
rect 601 40533 635 40537
rect 601 40503 635 40533
rect 601 40431 635 40465
rect 601 40363 635 40393
rect 601 40359 635 40363
rect 697 40533 731 40537
rect 697 40503 731 40533
rect 697 40431 731 40465
rect 697 40363 731 40393
rect 697 40359 731 40363
rect 793 40533 827 40537
rect 793 40503 827 40533
rect 793 40431 827 40465
rect 793 40363 827 40393
rect 793 40359 827 40363
rect 889 40533 923 40537
rect 889 40503 923 40533
rect 889 40431 923 40465
rect 889 40363 923 40393
rect 889 40359 923 40363
rect 985 40533 1019 40537
rect 985 40503 1019 40533
rect 985 40431 1019 40465
rect 985 40363 1019 40393
rect 985 40359 1019 40363
rect 1081 40533 1115 40537
rect 1081 40503 1115 40533
rect 1081 40431 1115 40465
rect 1081 40363 1115 40393
rect 1081 40359 1115 40363
rect 1177 40533 1211 40537
rect 1177 40503 1211 40533
rect 1177 40431 1211 40465
rect 1177 40363 1211 40393
rect 1177 40359 1211 40363
rect 1273 40533 1307 40537
rect 1273 40503 1307 40533
rect 1273 40431 1307 40465
rect 1273 40363 1307 40393
rect 1273 40359 1307 40363
rect 1387 40564 1421 40568
rect 1387 40534 1421 40564
rect 1387 40462 1421 40496
rect 1387 40394 1421 40424
rect 1387 40390 1421 40394
rect 1387 40326 1421 40352
rect 1387 40318 1421 40326
rect 2466 40636 2500 40670
rect 2658 40636 2692 40670
rect 2850 40636 2884 40670
rect 3042 40636 3076 40670
rect 3234 40636 3268 40670
rect 3426 40636 3460 40670
rect 3540 40636 3574 40644
rect 3540 40610 3574 40636
rect 2466 40537 2500 40541
rect 2466 40507 2500 40537
rect 2466 40435 2500 40469
rect 2466 40367 2500 40397
rect 2466 40363 2500 40367
rect 2562 40537 2596 40541
rect 2562 40507 2596 40537
rect 2562 40435 2596 40469
rect 2562 40367 2596 40397
rect 2562 40363 2596 40367
rect 2658 40537 2692 40541
rect 2658 40507 2692 40537
rect 2658 40435 2692 40469
rect 2658 40367 2692 40397
rect 2658 40363 2692 40367
rect 2754 40537 2788 40541
rect 2754 40507 2788 40537
rect 2754 40435 2788 40469
rect 2754 40367 2788 40397
rect 2754 40363 2788 40367
rect 2850 40537 2884 40541
rect 2850 40507 2884 40537
rect 2850 40435 2884 40469
rect 2850 40367 2884 40397
rect 2850 40363 2884 40367
rect 2946 40537 2980 40541
rect 2946 40507 2980 40537
rect 2946 40435 2980 40469
rect 2946 40367 2980 40397
rect 2946 40363 2980 40367
rect 3042 40537 3076 40541
rect 3042 40507 3076 40537
rect 3042 40435 3076 40469
rect 3042 40367 3076 40397
rect 3042 40363 3076 40367
rect 3138 40537 3172 40541
rect 3138 40507 3172 40537
rect 3138 40435 3172 40469
rect 3138 40367 3172 40397
rect 3138 40363 3172 40367
rect 3234 40537 3268 40541
rect 3234 40507 3268 40537
rect 3234 40435 3268 40469
rect 3234 40367 3268 40397
rect 3234 40363 3268 40367
rect 3330 40537 3364 40541
rect 3330 40507 3364 40537
rect 3330 40435 3364 40469
rect 3330 40367 3364 40397
rect 3330 40363 3364 40367
rect 3426 40537 3460 40541
rect 3426 40507 3460 40537
rect 3426 40435 3460 40469
rect 3426 40367 3460 40397
rect 3426 40363 3460 40367
rect 3540 40568 3574 40572
rect 3540 40538 3574 40568
rect 3540 40466 3574 40500
rect 3540 40398 3574 40428
rect 3540 40394 3574 40398
rect 3540 40330 3574 40356
rect 3540 40322 3574 40330
rect 3987 40636 4021 40670
rect 4179 40636 4213 40670
rect 4371 40636 4405 40670
rect 4563 40636 4597 40670
rect 4755 40636 4789 40670
rect 4947 40636 4981 40670
rect 5061 40636 5095 40644
rect 5061 40610 5095 40636
rect 3987 40537 4021 40541
rect 3987 40507 4021 40537
rect 3987 40435 4021 40469
rect 3987 40367 4021 40397
rect 3987 40363 4021 40367
rect 4083 40537 4117 40541
rect 4083 40507 4117 40537
rect 4083 40435 4117 40469
rect 4083 40367 4117 40397
rect 4083 40363 4117 40367
rect 4179 40537 4213 40541
rect 4179 40507 4213 40537
rect 4179 40435 4213 40469
rect 4179 40367 4213 40397
rect 4179 40363 4213 40367
rect 4275 40537 4309 40541
rect 4275 40507 4309 40537
rect 4275 40435 4309 40469
rect 4275 40367 4309 40397
rect 4275 40363 4309 40367
rect 4371 40537 4405 40541
rect 4371 40507 4405 40537
rect 4371 40435 4405 40469
rect 4371 40367 4405 40397
rect 4371 40363 4405 40367
rect 4467 40537 4501 40541
rect 4467 40507 4501 40537
rect 4467 40435 4501 40469
rect 4467 40367 4501 40397
rect 4467 40363 4501 40367
rect 4563 40537 4597 40541
rect 4563 40507 4597 40537
rect 4563 40435 4597 40469
rect 4563 40367 4597 40397
rect 4563 40363 4597 40367
rect 4659 40537 4693 40541
rect 4659 40507 4693 40537
rect 4659 40435 4693 40469
rect 4659 40367 4693 40397
rect 4659 40363 4693 40367
rect 4755 40537 4789 40541
rect 4755 40507 4789 40537
rect 4755 40435 4789 40469
rect 4755 40367 4789 40397
rect 4755 40363 4789 40367
rect 4851 40537 4885 40541
rect 4851 40507 4885 40537
rect 4851 40435 4885 40469
rect 4851 40367 4885 40397
rect 4851 40363 4885 40367
rect 4947 40537 4981 40541
rect 4947 40507 4981 40537
rect 4947 40435 4981 40469
rect 4947 40367 4981 40397
rect 4947 40363 4981 40367
rect 5061 40568 5095 40572
rect 5061 40538 5095 40568
rect 5061 40466 5095 40500
rect 5061 40398 5095 40428
rect 5303 40405 5337 40439
rect 5395 40405 5429 40439
rect 5487 40405 5521 40439
rect 5061 40394 5095 40398
rect 5061 40330 5095 40356
rect 5061 40322 5095 40330
rect 313 39935 347 39969
rect 409 39935 443 39969
rect 505 39935 539 39969
rect 601 39935 635 39969
rect 697 39935 731 39969
rect 793 39935 827 39969
rect 889 39935 923 39969
rect 985 39935 1019 39969
rect 1081 39935 1115 39969
rect 1177 39935 1211 39969
rect 1273 39935 1307 39969
rect 1387 40006 1421 40011
rect 1387 39977 1421 40006
rect 1387 39938 1421 39939
rect 1387 39905 1421 39938
rect 313 39824 347 39858
rect 505 39824 539 39858
rect 697 39824 731 39858
rect 889 39824 923 39858
rect 1081 39824 1115 39858
rect 1273 39824 1307 39858
rect 1387 39836 1421 39867
rect 1387 39833 1421 39836
rect 3691 40050 3725 40084
rect 2466 39939 2500 39973
rect 2562 39939 2596 39973
rect 2658 39939 2692 39973
rect 2754 39939 2788 39973
rect 2850 39939 2884 39973
rect 2946 39939 2980 39973
rect 3042 39939 3076 39973
rect 3138 39939 3172 39973
rect 3234 39939 3268 39973
rect 3330 39939 3364 39973
rect 3426 39939 3460 39973
rect 3540 40010 3574 40015
rect 3540 39981 3574 40010
rect 3540 39942 3574 39943
rect 3540 39909 3574 39942
rect 3647 39924 3681 40000
rect 3735 39924 3769 40000
rect 2466 39828 2500 39862
rect 2658 39828 2692 39862
rect 2850 39828 2884 39862
rect 3042 39828 3076 39862
rect 3234 39828 3268 39862
rect 3426 39828 3460 39862
rect 3540 39840 3574 39871
rect 3540 39837 3574 39840
rect 3987 39939 4021 39973
rect 4083 39939 4117 39973
rect 4179 39939 4213 39973
rect 4275 39939 4309 39973
rect 4371 39939 4405 39973
rect 4467 39939 4501 39973
rect 4563 39939 4597 39973
rect 4659 39939 4693 39973
rect 4755 39939 4789 39973
rect 4851 39939 4885 39973
rect 4947 39939 4981 39973
rect 5061 40010 5095 40015
rect 5061 39981 5095 40010
rect 5061 39942 5095 39943
rect 5061 39909 5095 39942
rect 5348 40091 5382 40125
rect 5450 40127 5484 40130
rect 5450 40096 5470 40127
rect 5470 40096 5484 40127
rect 3987 39828 4021 39862
rect 4179 39828 4213 39862
rect 4371 39828 4405 39862
rect 4563 39828 4597 39862
rect 4755 39828 4789 39862
rect 4947 39828 4981 39862
rect 5061 39840 5095 39871
rect 5303 39861 5337 39895
rect 5395 39861 5429 39895
rect 5487 39861 5521 39895
rect 5061 39837 5095 39840
rect 313 39345 347 39379
rect 505 39345 539 39379
rect 697 39345 731 39379
rect 889 39345 923 39379
rect 1081 39345 1115 39379
rect 1273 39345 1307 39379
rect 1387 39345 1421 39353
rect 1387 39319 1421 39345
rect 313 39246 347 39250
rect 313 39216 347 39246
rect 313 39144 347 39178
rect 313 39076 347 39106
rect 313 39072 347 39076
rect 409 39246 443 39250
rect 409 39216 443 39246
rect 409 39144 443 39178
rect 409 39076 443 39106
rect 409 39072 443 39076
rect 505 39246 539 39250
rect 505 39216 539 39246
rect 505 39144 539 39178
rect 505 39076 539 39106
rect 505 39072 539 39076
rect 601 39246 635 39250
rect 601 39216 635 39246
rect 601 39144 635 39178
rect 601 39076 635 39106
rect 601 39072 635 39076
rect 697 39246 731 39250
rect 697 39216 731 39246
rect 697 39144 731 39178
rect 697 39076 731 39106
rect 697 39072 731 39076
rect 793 39246 827 39250
rect 793 39216 827 39246
rect 793 39144 827 39178
rect 793 39076 827 39106
rect 793 39072 827 39076
rect 889 39246 923 39250
rect 889 39216 923 39246
rect 889 39144 923 39178
rect 889 39076 923 39106
rect 889 39072 923 39076
rect 985 39246 1019 39250
rect 985 39216 1019 39246
rect 985 39144 1019 39178
rect 985 39076 1019 39106
rect 985 39072 1019 39076
rect 1081 39246 1115 39250
rect 1081 39216 1115 39246
rect 1081 39144 1115 39178
rect 1081 39076 1115 39106
rect 1081 39072 1115 39076
rect 1177 39246 1211 39250
rect 1177 39216 1211 39246
rect 1177 39144 1211 39178
rect 1177 39076 1211 39106
rect 1177 39072 1211 39076
rect 1273 39246 1307 39250
rect 1273 39216 1307 39246
rect 1273 39144 1307 39178
rect 1273 39076 1307 39106
rect 1273 39072 1307 39076
rect 1387 39277 1421 39281
rect 1387 39247 1421 39277
rect 1387 39175 1421 39209
rect 1387 39107 1421 39137
rect 1387 39103 1421 39107
rect 1387 39039 1421 39065
rect 1387 39031 1421 39039
rect 2466 39349 2500 39383
rect 2658 39349 2692 39383
rect 2850 39349 2884 39383
rect 3042 39349 3076 39383
rect 3234 39349 3268 39383
rect 3426 39349 3460 39383
rect 3540 39349 3574 39357
rect 3540 39323 3574 39349
rect 2466 39250 2500 39254
rect 2466 39220 2500 39250
rect 2466 39148 2500 39182
rect 2466 39080 2500 39110
rect 2466 39076 2500 39080
rect 2562 39250 2596 39254
rect 2562 39220 2596 39250
rect 2562 39148 2596 39182
rect 2562 39080 2596 39110
rect 2562 39076 2596 39080
rect 2658 39250 2692 39254
rect 2658 39220 2692 39250
rect 2658 39148 2692 39182
rect 2658 39080 2692 39110
rect 2658 39076 2692 39080
rect 2754 39250 2788 39254
rect 2754 39220 2788 39250
rect 2754 39148 2788 39182
rect 2754 39080 2788 39110
rect 2754 39076 2788 39080
rect 2850 39250 2884 39254
rect 2850 39220 2884 39250
rect 2850 39148 2884 39182
rect 2850 39080 2884 39110
rect 2850 39076 2884 39080
rect 2946 39250 2980 39254
rect 2946 39220 2980 39250
rect 2946 39148 2980 39182
rect 2946 39080 2980 39110
rect 2946 39076 2980 39080
rect 3042 39250 3076 39254
rect 3042 39220 3076 39250
rect 3042 39148 3076 39182
rect 3042 39080 3076 39110
rect 3042 39076 3076 39080
rect 3138 39250 3172 39254
rect 3138 39220 3172 39250
rect 3138 39148 3172 39182
rect 3138 39080 3172 39110
rect 3138 39076 3172 39080
rect 3234 39250 3268 39254
rect 3234 39220 3268 39250
rect 3234 39148 3268 39182
rect 3234 39080 3268 39110
rect 3234 39076 3268 39080
rect 3330 39250 3364 39254
rect 3330 39220 3364 39250
rect 3330 39148 3364 39182
rect 3330 39080 3364 39110
rect 3330 39076 3364 39080
rect 3426 39250 3460 39254
rect 3426 39220 3460 39250
rect 3426 39148 3460 39182
rect 3426 39080 3460 39110
rect 3426 39076 3460 39080
rect 3540 39281 3574 39285
rect 3540 39251 3574 39281
rect 3540 39179 3574 39213
rect 3540 39111 3574 39141
rect 3540 39107 3574 39111
rect 3540 39043 3574 39069
rect 3540 39035 3574 39043
rect 3987 39349 4021 39383
rect 4179 39349 4213 39383
rect 4371 39349 4405 39383
rect 4563 39349 4597 39383
rect 4755 39349 4789 39383
rect 4947 39349 4981 39383
rect 5061 39349 5095 39357
rect 5061 39323 5095 39349
rect 3987 39250 4021 39254
rect 3987 39220 4021 39250
rect 3987 39148 4021 39182
rect 3987 39080 4021 39110
rect 3987 39076 4021 39080
rect 4083 39250 4117 39254
rect 4083 39220 4117 39250
rect 4083 39148 4117 39182
rect 4083 39080 4117 39110
rect 4083 39076 4117 39080
rect 4179 39250 4213 39254
rect 4179 39220 4213 39250
rect 4179 39148 4213 39182
rect 4179 39080 4213 39110
rect 4179 39076 4213 39080
rect 4275 39250 4309 39254
rect 4275 39220 4309 39250
rect 4275 39148 4309 39182
rect 4275 39080 4309 39110
rect 4275 39076 4309 39080
rect 4371 39250 4405 39254
rect 4371 39220 4405 39250
rect 4371 39148 4405 39182
rect 4371 39080 4405 39110
rect 4371 39076 4405 39080
rect 4467 39250 4501 39254
rect 4467 39220 4501 39250
rect 4467 39148 4501 39182
rect 4467 39080 4501 39110
rect 4467 39076 4501 39080
rect 4563 39250 4597 39254
rect 4563 39220 4597 39250
rect 4563 39148 4597 39182
rect 4563 39080 4597 39110
rect 4563 39076 4597 39080
rect 4659 39250 4693 39254
rect 4659 39220 4693 39250
rect 4659 39148 4693 39182
rect 4659 39080 4693 39110
rect 4659 39076 4693 39080
rect 4755 39250 4789 39254
rect 4755 39220 4789 39250
rect 4755 39148 4789 39182
rect 4755 39080 4789 39110
rect 4755 39076 4789 39080
rect 4851 39250 4885 39254
rect 4851 39220 4885 39250
rect 4851 39148 4885 39182
rect 4851 39080 4885 39110
rect 4851 39076 4885 39080
rect 4947 39250 4981 39254
rect 4947 39220 4981 39250
rect 4947 39148 4981 39182
rect 4947 39080 4981 39110
rect 4947 39076 4981 39080
rect 5061 39281 5095 39285
rect 5061 39251 5095 39281
rect 5061 39179 5095 39213
rect 5061 39111 5095 39141
rect 5303 39118 5337 39152
rect 5395 39118 5429 39152
rect 5487 39118 5521 39152
rect 5061 39107 5095 39111
rect 5061 39043 5095 39069
rect 5061 39035 5095 39043
rect 313 38648 347 38682
rect 409 38648 443 38682
rect 505 38648 539 38682
rect 601 38648 635 38682
rect 697 38648 731 38682
rect 793 38648 827 38682
rect 889 38648 923 38682
rect 985 38648 1019 38682
rect 1081 38648 1115 38682
rect 1177 38648 1211 38682
rect 1273 38648 1307 38682
rect 1387 38719 1421 38724
rect 1387 38690 1421 38719
rect 1387 38651 1421 38652
rect 1387 38618 1421 38651
rect 313 38537 347 38571
rect 505 38537 539 38571
rect 697 38537 731 38571
rect 889 38537 923 38571
rect 1081 38537 1115 38571
rect 1273 38537 1307 38571
rect 1387 38549 1421 38580
rect 1387 38546 1421 38549
rect 3691 38763 3725 38797
rect 2466 38652 2500 38686
rect 2562 38652 2596 38686
rect 2658 38652 2692 38686
rect 2754 38652 2788 38686
rect 2850 38652 2884 38686
rect 2946 38652 2980 38686
rect 3042 38652 3076 38686
rect 3138 38652 3172 38686
rect 3234 38652 3268 38686
rect 3330 38652 3364 38686
rect 3426 38652 3460 38686
rect 3540 38723 3574 38728
rect 3540 38694 3574 38723
rect 3540 38655 3574 38656
rect 3540 38622 3574 38655
rect 3647 38637 3681 38713
rect 3735 38637 3769 38713
rect 2466 38541 2500 38575
rect 2658 38541 2692 38575
rect 2850 38541 2884 38575
rect 3042 38541 3076 38575
rect 3234 38541 3268 38575
rect 3426 38541 3460 38575
rect 3540 38553 3574 38584
rect 3540 38550 3574 38553
rect 3987 38652 4021 38686
rect 4083 38652 4117 38686
rect 4179 38652 4213 38686
rect 4275 38652 4309 38686
rect 4371 38652 4405 38686
rect 4467 38652 4501 38686
rect 4563 38652 4597 38686
rect 4659 38652 4693 38686
rect 4755 38652 4789 38686
rect 4851 38652 4885 38686
rect 4947 38652 4981 38686
rect 5061 38723 5095 38728
rect 5061 38694 5095 38723
rect 5061 38655 5095 38656
rect 5061 38622 5095 38655
rect 5348 38804 5382 38838
rect 5450 38840 5484 38843
rect 5450 38809 5470 38840
rect 5470 38809 5484 38840
rect 3987 38541 4021 38575
rect 4179 38541 4213 38575
rect 4371 38541 4405 38575
rect 4563 38541 4597 38575
rect 4755 38541 4789 38575
rect 4947 38541 4981 38575
rect 5061 38553 5095 38584
rect 5303 38574 5337 38608
rect 5395 38574 5429 38608
rect 5487 38574 5521 38608
rect 5061 38550 5095 38553
rect 313 38058 347 38092
rect 505 38058 539 38092
rect 697 38058 731 38092
rect 889 38058 923 38092
rect 1081 38058 1115 38092
rect 1273 38058 1307 38092
rect 1387 38058 1421 38066
rect 1387 38032 1421 38058
rect 313 37959 347 37963
rect 313 37929 347 37959
rect 313 37857 347 37891
rect 313 37789 347 37819
rect 313 37785 347 37789
rect 409 37959 443 37963
rect 409 37929 443 37959
rect 409 37857 443 37891
rect 409 37789 443 37819
rect 409 37785 443 37789
rect 505 37959 539 37963
rect 505 37929 539 37959
rect 505 37857 539 37891
rect 505 37789 539 37819
rect 505 37785 539 37789
rect 601 37959 635 37963
rect 601 37929 635 37959
rect 601 37857 635 37891
rect 601 37789 635 37819
rect 601 37785 635 37789
rect 697 37959 731 37963
rect 697 37929 731 37959
rect 697 37857 731 37891
rect 697 37789 731 37819
rect 697 37785 731 37789
rect 793 37959 827 37963
rect 793 37929 827 37959
rect 793 37857 827 37891
rect 793 37789 827 37819
rect 793 37785 827 37789
rect 889 37959 923 37963
rect 889 37929 923 37959
rect 889 37857 923 37891
rect 889 37789 923 37819
rect 889 37785 923 37789
rect 985 37959 1019 37963
rect 985 37929 1019 37959
rect 985 37857 1019 37891
rect 985 37789 1019 37819
rect 985 37785 1019 37789
rect 1081 37959 1115 37963
rect 1081 37929 1115 37959
rect 1081 37857 1115 37891
rect 1081 37789 1115 37819
rect 1081 37785 1115 37789
rect 1177 37959 1211 37963
rect 1177 37929 1211 37959
rect 1177 37857 1211 37891
rect 1177 37789 1211 37819
rect 1177 37785 1211 37789
rect 1273 37959 1307 37963
rect 1273 37929 1307 37959
rect 1273 37857 1307 37891
rect 1273 37789 1307 37819
rect 1273 37785 1307 37789
rect 1387 37990 1421 37994
rect 1387 37960 1421 37990
rect 1387 37888 1421 37922
rect 1387 37820 1421 37850
rect 1387 37816 1421 37820
rect 1387 37752 1421 37778
rect 1387 37744 1421 37752
rect 2466 38062 2500 38096
rect 2658 38062 2692 38096
rect 2850 38062 2884 38096
rect 3042 38062 3076 38096
rect 3234 38062 3268 38096
rect 3426 38062 3460 38096
rect 3540 38062 3574 38070
rect 3540 38036 3574 38062
rect 2466 37963 2500 37967
rect 2466 37933 2500 37963
rect 2466 37861 2500 37895
rect 2466 37793 2500 37823
rect 2466 37789 2500 37793
rect 2562 37963 2596 37967
rect 2562 37933 2596 37963
rect 2562 37861 2596 37895
rect 2562 37793 2596 37823
rect 2562 37789 2596 37793
rect 2658 37963 2692 37967
rect 2658 37933 2692 37963
rect 2658 37861 2692 37895
rect 2658 37793 2692 37823
rect 2658 37789 2692 37793
rect 2754 37963 2788 37967
rect 2754 37933 2788 37963
rect 2754 37861 2788 37895
rect 2754 37793 2788 37823
rect 2754 37789 2788 37793
rect 2850 37963 2884 37967
rect 2850 37933 2884 37963
rect 2850 37861 2884 37895
rect 2850 37793 2884 37823
rect 2850 37789 2884 37793
rect 2946 37963 2980 37967
rect 2946 37933 2980 37963
rect 2946 37861 2980 37895
rect 2946 37793 2980 37823
rect 2946 37789 2980 37793
rect 3042 37963 3076 37967
rect 3042 37933 3076 37963
rect 3042 37861 3076 37895
rect 3042 37793 3076 37823
rect 3042 37789 3076 37793
rect 3138 37963 3172 37967
rect 3138 37933 3172 37963
rect 3138 37861 3172 37895
rect 3138 37793 3172 37823
rect 3138 37789 3172 37793
rect 3234 37963 3268 37967
rect 3234 37933 3268 37963
rect 3234 37861 3268 37895
rect 3234 37793 3268 37823
rect 3234 37789 3268 37793
rect 3330 37963 3364 37967
rect 3330 37933 3364 37963
rect 3330 37861 3364 37895
rect 3330 37793 3364 37823
rect 3330 37789 3364 37793
rect 3426 37963 3460 37967
rect 3426 37933 3460 37963
rect 3426 37861 3460 37895
rect 3426 37793 3460 37823
rect 3426 37789 3460 37793
rect 3540 37994 3574 37998
rect 3540 37964 3574 37994
rect 3540 37892 3574 37926
rect 3540 37824 3574 37854
rect 3540 37820 3574 37824
rect 3540 37756 3574 37782
rect 3540 37748 3574 37756
rect 3987 38062 4021 38096
rect 4179 38062 4213 38096
rect 4371 38062 4405 38096
rect 4563 38062 4597 38096
rect 4755 38062 4789 38096
rect 4947 38062 4981 38096
rect 5061 38062 5095 38070
rect 5061 38036 5095 38062
rect 3987 37963 4021 37967
rect 3987 37933 4021 37963
rect 3987 37861 4021 37895
rect 3987 37793 4021 37823
rect 3987 37789 4021 37793
rect 4083 37963 4117 37967
rect 4083 37933 4117 37963
rect 4083 37861 4117 37895
rect 4083 37793 4117 37823
rect 4083 37789 4117 37793
rect 4179 37963 4213 37967
rect 4179 37933 4213 37963
rect 4179 37861 4213 37895
rect 4179 37793 4213 37823
rect 4179 37789 4213 37793
rect 4275 37963 4309 37967
rect 4275 37933 4309 37963
rect 4275 37861 4309 37895
rect 4275 37793 4309 37823
rect 4275 37789 4309 37793
rect 4371 37963 4405 37967
rect 4371 37933 4405 37963
rect 4371 37861 4405 37895
rect 4371 37793 4405 37823
rect 4371 37789 4405 37793
rect 4467 37963 4501 37967
rect 4467 37933 4501 37963
rect 4467 37861 4501 37895
rect 4467 37793 4501 37823
rect 4467 37789 4501 37793
rect 4563 37963 4597 37967
rect 4563 37933 4597 37963
rect 4563 37861 4597 37895
rect 4563 37793 4597 37823
rect 4563 37789 4597 37793
rect 4659 37963 4693 37967
rect 4659 37933 4693 37963
rect 4659 37861 4693 37895
rect 4659 37793 4693 37823
rect 4659 37789 4693 37793
rect 4755 37963 4789 37967
rect 4755 37933 4789 37963
rect 4755 37861 4789 37895
rect 4755 37793 4789 37823
rect 4755 37789 4789 37793
rect 4851 37963 4885 37967
rect 4851 37933 4885 37963
rect 4851 37861 4885 37895
rect 4851 37793 4885 37823
rect 4851 37789 4885 37793
rect 4947 37963 4981 37967
rect 4947 37933 4981 37963
rect 4947 37861 4981 37895
rect 4947 37793 4981 37823
rect 4947 37789 4981 37793
rect 5061 37994 5095 37998
rect 5061 37964 5095 37994
rect 5061 37892 5095 37926
rect 5061 37824 5095 37854
rect 5303 37831 5337 37865
rect 5395 37831 5429 37865
rect 5487 37831 5521 37865
rect 5061 37820 5095 37824
rect 5061 37756 5095 37782
rect 5061 37748 5095 37756
rect 313 37361 347 37395
rect 409 37361 443 37395
rect 505 37361 539 37395
rect 601 37361 635 37395
rect 697 37361 731 37395
rect 793 37361 827 37395
rect 889 37361 923 37395
rect 985 37361 1019 37395
rect 1081 37361 1115 37395
rect 1177 37361 1211 37395
rect 1273 37361 1307 37395
rect 1387 37432 1421 37437
rect 1387 37403 1421 37432
rect 1387 37364 1421 37365
rect 1387 37331 1421 37364
rect 313 37250 347 37284
rect 505 37250 539 37284
rect 697 37250 731 37284
rect 889 37250 923 37284
rect 1081 37250 1115 37284
rect 1273 37250 1307 37284
rect 1387 37262 1421 37293
rect 1387 37259 1421 37262
rect 3691 37476 3725 37510
rect 2466 37365 2500 37399
rect 2562 37365 2596 37399
rect 2658 37365 2692 37399
rect 2754 37365 2788 37399
rect 2850 37365 2884 37399
rect 2946 37365 2980 37399
rect 3042 37365 3076 37399
rect 3138 37365 3172 37399
rect 3234 37365 3268 37399
rect 3330 37365 3364 37399
rect 3426 37365 3460 37399
rect 3540 37436 3574 37441
rect 3540 37407 3574 37436
rect 3540 37368 3574 37369
rect 3540 37335 3574 37368
rect 3647 37350 3681 37426
rect 3735 37350 3769 37426
rect 2466 37254 2500 37288
rect 2658 37254 2692 37288
rect 2850 37254 2884 37288
rect 3042 37254 3076 37288
rect 3234 37254 3268 37288
rect 3426 37254 3460 37288
rect 3540 37266 3574 37297
rect 3540 37263 3574 37266
rect 3987 37365 4021 37399
rect 4083 37365 4117 37399
rect 4179 37365 4213 37399
rect 4275 37365 4309 37399
rect 4371 37365 4405 37399
rect 4467 37365 4501 37399
rect 4563 37365 4597 37399
rect 4659 37365 4693 37399
rect 4755 37365 4789 37399
rect 4851 37365 4885 37399
rect 4947 37365 4981 37399
rect 5061 37436 5095 37441
rect 5061 37407 5095 37436
rect 5061 37368 5095 37369
rect 5061 37335 5095 37368
rect 5348 37517 5382 37551
rect 5450 37553 5484 37556
rect 5450 37522 5470 37553
rect 5470 37522 5484 37553
rect 3987 37254 4021 37288
rect 4179 37254 4213 37288
rect 4371 37254 4405 37288
rect 4563 37254 4597 37288
rect 4755 37254 4789 37288
rect 4947 37254 4981 37288
rect 5061 37266 5095 37297
rect 5303 37287 5337 37321
rect 5395 37287 5429 37321
rect 5487 37287 5521 37321
rect 5061 37263 5095 37266
rect 313 36771 347 36805
rect 505 36771 539 36805
rect 697 36771 731 36805
rect 889 36771 923 36805
rect 1081 36771 1115 36805
rect 1273 36771 1307 36805
rect 1387 36771 1421 36779
rect 1387 36745 1421 36771
rect 313 36672 347 36676
rect 313 36642 347 36672
rect 313 36570 347 36604
rect 313 36502 347 36532
rect 313 36498 347 36502
rect 409 36672 443 36676
rect 409 36642 443 36672
rect 409 36570 443 36604
rect 409 36502 443 36532
rect 409 36498 443 36502
rect 505 36672 539 36676
rect 505 36642 539 36672
rect 505 36570 539 36604
rect 505 36502 539 36532
rect 505 36498 539 36502
rect 601 36672 635 36676
rect 601 36642 635 36672
rect 601 36570 635 36604
rect 601 36502 635 36532
rect 601 36498 635 36502
rect 697 36672 731 36676
rect 697 36642 731 36672
rect 697 36570 731 36604
rect 697 36502 731 36532
rect 697 36498 731 36502
rect 793 36672 827 36676
rect 793 36642 827 36672
rect 793 36570 827 36604
rect 793 36502 827 36532
rect 793 36498 827 36502
rect 889 36672 923 36676
rect 889 36642 923 36672
rect 889 36570 923 36604
rect 889 36502 923 36532
rect 889 36498 923 36502
rect 985 36672 1019 36676
rect 985 36642 1019 36672
rect 985 36570 1019 36604
rect 985 36502 1019 36532
rect 985 36498 1019 36502
rect 1081 36672 1115 36676
rect 1081 36642 1115 36672
rect 1081 36570 1115 36604
rect 1081 36502 1115 36532
rect 1081 36498 1115 36502
rect 1177 36672 1211 36676
rect 1177 36642 1211 36672
rect 1177 36570 1211 36604
rect 1177 36502 1211 36532
rect 1177 36498 1211 36502
rect 1273 36672 1307 36676
rect 1273 36642 1307 36672
rect 1273 36570 1307 36604
rect 1273 36502 1307 36532
rect 1273 36498 1307 36502
rect 1387 36703 1421 36707
rect 1387 36673 1421 36703
rect 1387 36601 1421 36635
rect 1387 36533 1421 36563
rect 1387 36529 1421 36533
rect 1387 36465 1421 36491
rect 1387 36457 1421 36465
rect 2466 36775 2500 36809
rect 2658 36775 2692 36809
rect 2850 36775 2884 36809
rect 3042 36775 3076 36809
rect 3234 36775 3268 36809
rect 3426 36775 3460 36809
rect 3540 36775 3574 36783
rect 3540 36749 3574 36775
rect 2466 36676 2500 36680
rect 2466 36646 2500 36676
rect 2466 36574 2500 36608
rect 2466 36506 2500 36536
rect 2466 36502 2500 36506
rect 2562 36676 2596 36680
rect 2562 36646 2596 36676
rect 2562 36574 2596 36608
rect 2562 36506 2596 36536
rect 2562 36502 2596 36506
rect 2658 36676 2692 36680
rect 2658 36646 2692 36676
rect 2658 36574 2692 36608
rect 2658 36506 2692 36536
rect 2658 36502 2692 36506
rect 2754 36676 2788 36680
rect 2754 36646 2788 36676
rect 2754 36574 2788 36608
rect 2754 36506 2788 36536
rect 2754 36502 2788 36506
rect 2850 36676 2884 36680
rect 2850 36646 2884 36676
rect 2850 36574 2884 36608
rect 2850 36506 2884 36536
rect 2850 36502 2884 36506
rect 2946 36676 2980 36680
rect 2946 36646 2980 36676
rect 2946 36574 2980 36608
rect 2946 36506 2980 36536
rect 2946 36502 2980 36506
rect 3042 36676 3076 36680
rect 3042 36646 3076 36676
rect 3042 36574 3076 36608
rect 3042 36506 3076 36536
rect 3042 36502 3076 36506
rect 3138 36676 3172 36680
rect 3138 36646 3172 36676
rect 3138 36574 3172 36608
rect 3138 36506 3172 36536
rect 3138 36502 3172 36506
rect 3234 36676 3268 36680
rect 3234 36646 3268 36676
rect 3234 36574 3268 36608
rect 3234 36506 3268 36536
rect 3234 36502 3268 36506
rect 3330 36676 3364 36680
rect 3330 36646 3364 36676
rect 3330 36574 3364 36608
rect 3330 36506 3364 36536
rect 3330 36502 3364 36506
rect 3426 36676 3460 36680
rect 3426 36646 3460 36676
rect 3426 36574 3460 36608
rect 3426 36506 3460 36536
rect 3426 36502 3460 36506
rect 3540 36707 3574 36711
rect 3540 36677 3574 36707
rect 3540 36605 3574 36639
rect 3540 36537 3574 36567
rect 3540 36533 3574 36537
rect 3540 36469 3574 36495
rect 3540 36461 3574 36469
rect 3987 36775 4021 36809
rect 4179 36775 4213 36809
rect 4371 36775 4405 36809
rect 4563 36775 4597 36809
rect 4755 36775 4789 36809
rect 4947 36775 4981 36809
rect 5061 36775 5095 36783
rect 5061 36749 5095 36775
rect 3987 36676 4021 36680
rect 3987 36646 4021 36676
rect 3987 36574 4021 36608
rect 3987 36506 4021 36536
rect 3987 36502 4021 36506
rect 4083 36676 4117 36680
rect 4083 36646 4117 36676
rect 4083 36574 4117 36608
rect 4083 36506 4117 36536
rect 4083 36502 4117 36506
rect 4179 36676 4213 36680
rect 4179 36646 4213 36676
rect 4179 36574 4213 36608
rect 4179 36506 4213 36536
rect 4179 36502 4213 36506
rect 4275 36676 4309 36680
rect 4275 36646 4309 36676
rect 4275 36574 4309 36608
rect 4275 36506 4309 36536
rect 4275 36502 4309 36506
rect 4371 36676 4405 36680
rect 4371 36646 4405 36676
rect 4371 36574 4405 36608
rect 4371 36506 4405 36536
rect 4371 36502 4405 36506
rect 4467 36676 4501 36680
rect 4467 36646 4501 36676
rect 4467 36574 4501 36608
rect 4467 36506 4501 36536
rect 4467 36502 4501 36506
rect 4563 36676 4597 36680
rect 4563 36646 4597 36676
rect 4563 36574 4597 36608
rect 4563 36506 4597 36536
rect 4563 36502 4597 36506
rect 4659 36676 4693 36680
rect 4659 36646 4693 36676
rect 4659 36574 4693 36608
rect 4659 36506 4693 36536
rect 4659 36502 4693 36506
rect 4755 36676 4789 36680
rect 4755 36646 4789 36676
rect 4755 36574 4789 36608
rect 4755 36506 4789 36536
rect 4755 36502 4789 36506
rect 4851 36676 4885 36680
rect 4851 36646 4885 36676
rect 4851 36574 4885 36608
rect 4851 36506 4885 36536
rect 4851 36502 4885 36506
rect 4947 36676 4981 36680
rect 4947 36646 4981 36676
rect 4947 36574 4981 36608
rect 4947 36506 4981 36536
rect 4947 36502 4981 36506
rect 5061 36707 5095 36711
rect 5061 36677 5095 36707
rect 5061 36605 5095 36639
rect 5061 36537 5095 36567
rect 5303 36544 5337 36578
rect 5395 36544 5429 36578
rect 5487 36544 5521 36578
rect 5061 36533 5095 36537
rect 5061 36469 5095 36495
rect 5061 36461 5095 36469
rect 313 36074 347 36108
rect 409 36074 443 36108
rect 505 36074 539 36108
rect 601 36074 635 36108
rect 697 36074 731 36108
rect 793 36074 827 36108
rect 889 36074 923 36108
rect 985 36074 1019 36108
rect 1081 36074 1115 36108
rect 1177 36074 1211 36108
rect 1273 36074 1307 36108
rect 1387 36145 1421 36150
rect 1387 36116 1421 36145
rect 1387 36077 1421 36078
rect 1387 36044 1421 36077
rect 313 35963 347 35997
rect 505 35963 539 35997
rect 697 35963 731 35997
rect 889 35963 923 35997
rect 1081 35963 1115 35997
rect 1273 35963 1307 35997
rect 1387 35975 1421 36006
rect 1387 35972 1421 35975
rect 3691 36189 3725 36223
rect 2466 36078 2500 36112
rect 2562 36078 2596 36112
rect 2658 36078 2692 36112
rect 2754 36078 2788 36112
rect 2850 36078 2884 36112
rect 2946 36078 2980 36112
rect 3042 36078 3076 36112
rect 3138 36078 3172 36112
rect 3234 36078 3268 36112
rect 3330 36078 3364 36112
rect 3426 36078 3460 36112
rect 3540 36149 3574 36154
rect 3540 36120 3574 36149
rect 3540 36081 3574 36082
rect 3540 36048 3574 36081
rect 3647 36063 3681 36139
rect 3735 36063 3769 36139
rect 2466 35967 2500 36001
rect 2658 35967 2692 36001
rect 2850 35967 2884 36001
rect 3042 35967 3076 36001
rect 3234 35967 3268 36001
rect 3426 35967 3460 36001
rect 3540 35979 3574 36010
rect 3540 35976 3574 35979
rect 3987 36078 4021 36112
rect 4083 36078 4117 36112
rect 4179 36078 4213 36112
rect 4275 36078 4309 36112
rect 4371 36078 4405 36112
rect 4467 36078 4501 36112
rect 4563 36078 4597 36112
rect 4659 36078 4693 36112
rect 4755 36078 4789 36112
rect 4851 36078 4885 36112
rect 4947 36078 4981 36112
rect 5061 36149 5095 36154
rect 5061 36120 5095 36149
rect 5061 36081 5095 36082
rect 5061 36048 5095 36081
rect 5348 36230 5382 36264
rect 5450 36266 5484 36269
rect 5450 36235 5470 36266
rect 5470 36235 5484 36266
rect 3987 35967 4021 36001
rect 4179 35967 4213 36001
rect 4371 35967 4405 36001
rect 4563 35967 4597 36001
rect 4755 35967 4789 36001
rect 4947 35967 4981 36001
rect 5061 35979 5095 36010
rect 5303 36000 5337 36034
rect 5395 36000 5429 36034
rect 5487 36000 5521 36034
rect 5061 35976 5095 35979
rect 313 35484 347 35518
rect 505 35484 539 35518
rect 697 35484 731 35518
rect 889 35484 923 35518
rect 1081 35484 1115 35518
rect 1273 35484 1307 35518
rect 1387 35484 1421 35492
rect 1387 35458 1421 35484
rect 313 35385 347 35389
rect 313 35355 347 35385
rect 313 35283 347 35317
rect 313 35215 347 35245
rect 313 35211 347 35215
rect 409 35385 443 35389
rect 409 35355 443 35385
rect 409 35283 443 35317
rect 409 35215 443 35245
rect 409 35211 443 35215
rect 505 35385 539 35389
rect 505 35355 539 35385
rect 505 35283 539 35317
rect 505 35215 539 35245
rect 505 35211 539 35215
rect 601 35385 635 35389
rect 601 35355 635 35385
rect 601 35283 635 35317
rect 601 35215 635 35245
rect 601 35211 635 35215
rect 697 35385 731 35389
rect 697 35355 731 35385
rect 697 35283 731 35317
rect 697 35215 731 35245
rect 697 35211 731 35215
rect 793 35385 827 35389
rect 793 35355 827 35385
rect 793 35283 827 35317
rect 793 35215 827 35245
rect 793 35211 827 35215
rect 889 35385 923 35389
rect 889 35355 923 35385
rect 889 35283 923 35317
rect 889 35215 923 35245
rect 889 35211 923 35215
rect 985 35385 1019 35389
rect 985 35355 1019 35385
rect 985 35283 1019 35317
rect 985 35215 1019 35245
rect 985 35211 1019 35215
rect 1081 35385 1115 35389
rect 1081 35355 1115 35385
rect 1081 35283 1115 35317
rect 1081 35215 1115 35245
rect 1081 35211 1115 35215
rect 1177 35385 1211 35389
rect 1177 35355 1211 35385
rect 1177 35283 1211 35317
rect 1177 35215 1211 35245
rect 1177 35211 1211 35215
rect 1273 35385 1307 35389
rect 1273 35355 1307 35385
rect 1273 35283 1307 35317
rect 1273 35215 1307 35245
rect 1273 35211 1307 35215
rect 1387 35416 1421 35420
rect 1387 35386 1421 35416
rect 1387 35314 1421 35348
rect 1387 35246 1421 35276
rect 1387 35242 1421 35246
rect 1387 35178 1421 35204
rect 1387 35170 1421 35178
rect 2466 35488 2500 35522
rect 2658 35488 2692 35522
rect 2850 35488 2884 35522
rect 3042 35488 3076 35522
rect 3234 35488 3268 35522
rect 3426 35488 3460 35522
rect 3540 35488 3574 35496
rect 3540 35462 3574 35488
rect 2466 35389 2500 35393
rect 2466 35359 2500 35389
rect 2466 35287 2500 35321
rect 2466 35219 2500 35249
rect 2466 35215 2500 35219
rect 2562 35389 2596 35393
rect 2562 35359 2596 35389
rect 2562 35287 2596 35321
rect 2562 35219 2596 35249
rect 2562 35215 2596 35219
rect 2658 35389 2692 35393
rect 2658 35359 2692 35389
rect 2658 35287 2692 35321
rect 2658 35219 2692 35249
rect 2658 35215 2692 35219
rect 2754 35389 2788 35393
rect 2754 35359 2788 35389
rect 2754 35287 2788 35321
rect 2754 35219 2788 35249
rect 2754 35215 2788 35219
rect 2850 35389 2884 35393
rect 2850 35359 2884 35389
rect 2850 35287 2884 35321
rect 2850 35219 2884 35249
rect 2850 35215 2884 35219
rect 2946 35389 2980 35393
rect 2946 35359 2980 35389
rect 2946 35287 2980 35321
rect 2946 35219 2980 35249
rect 2946 35215 2980 35219
rect 3042 35389 3076 35393
rect 3042 35359 3076 35389
rect 3042 35287 3076 35321
rect 3042 35219 3076 35249
rect 3042 35215 3076 35219
rect 3138 35389 3172 35393
rect 3138 35359 3172 35389
rect 3138 35287 3172 35321
rect 3138 35219 3172 35249
rect 3138 35215 3172 35219
rect 3234 35389 3268 35393
rect 3234 35359 3268 35389
rect 3234 35287 3268 35321
rect 3234 35219 3268 35249
rect 3234 35215 3268 35219
rect 3330 35389 3364 35393
rect 3330 35359 3364 35389
rect 3330 35287 3364 35321
rect 3330 35219 3364 35249
rect 3330 35215 3364 35219
rect 3426 35389 3460 35393
rect 3426 35359 3460 35389
rect 3426 35287 3460 35321
rect 3426 35219 3460 35249
rect 3426 35215 3460 35219
rect 3540 35420 3574 35424
rect 3540 35390 3574 35420
rect 3540 35318 3574 35352
rect 3540 35250 3574 35280
rect 3540 35246 3574 35250
rect 3540 35182 3574 35208
rect 3540 35174 3574 35182
rect 3987 35488 4021 35522
rect 4179 35488 4213 35522
rect 4371 35488 4405 35522
rect 4563 35488 4597 35522
rect 4755 35488 4789 35522
rect 4947 35488 4981 35522
rect 5061 35488 5095 35496
rect 5061 35462 5095 35488
rect 3987 35389 4021 35393
rect 3987 35359 4021 35389
rect 3987 35287 4021 35321
rect 3987 35219 4021 35249
rect 3987 35215 4021 35219
rect 4083 35389 4117 35393
rect 4083 35359 4117 35389
rect 4083 35287 4117 35321
rect 4083 35219 4117 35249
rect 4083 35215 4117 35219
rect 4179 35389 4213 35393
rect 4179 35359 4213 35389
rect 4179 35287 4213 35321
rect 4179 35219 4213 35249
rect 4179 35215 4213 35219
rect 4275 35389 4309 35393
rect 4275 35359 4309 35389
rect 4275 35287 4309 35321
rect 4275 35219 4309 35249
rect 4275 35215 4309 35219
rect 4371 35389 4405 35393
rect 4371 35359 4405 35389
rect 4371 35287 4405 35321
rect 4371 35219 4405 35249
rect 4371 35215 4405 35219
rect 4467 35389 4501 35393
rect 4467 35359 4501 35389
rect 4467 35287 4501 35321
rect 4467 35219 4501 35249
rect 4467 35215 4501 35219
rect 4563 35389 4597 35393
rect 4563 35359 4597 35389
rect 4563 35287 4597 35321
rect 4563 35219 4597 35249
rect 4563 35215 4597 35219
rect 4659 35389 4693 35393
rect 4659 35359 4693 35389
rect 4659 35287 4693 35321
rect 4659 35219 4693 35249
rect 4659 35215 4693 35219
rect 4755 35389 4789 35393
rect 4755 35359 4789 35389
rect 4755 35287 4789 35321
rect 4755 35219 4789 35249
rect 4755 35215 4789 35219
rect 4851 35389 4885 35393
rect 4851 35359 4885 35389
rect 4851 35287 4885 35321
rect 4851 35219 4885 35249
rect 4851 35215 4885 35219
rect 4947 35389 4981 35393
rect 4947 35359 4981 35389
rect 4947 35287 4981 35321
rect 4947 35219 4981 35249
rect 4947 35215 4981 35219
rect 5061 35420 5095 35424
rect 5061 35390 5095 35420
rect 5061 35318 5095 35352
rect 5061 35250 5095 35280
rect 5303 35257 5337 35291
rect 5395 35257 5429 35291
rect 5487 35257 5521 35291
rect 5061 35246 5095 35250
rect 5061 35182 5095 35208
rect 5061 35174 5095 35182
rect 313 34787 347 34821
rect 409 34787 443 34821
rect 505 34787 539 34821
rect 601 34787 635 34821
rect 697 34787 731 34821
rect 793 34787 827 34821
rect 889 34787 923 34821
rect 985 34787 1019 34821
rect 1081 34787 1115 34821
rect 1177 34787 1211 34821
rect 1273 34787 1307 34821
rect 1387 34858 1421 34863
rect 1387 34829 1421 34858
rect 1387 34790 1421 34791
rect 1387 34757 1421 34790
rect 313 34676 347 34710
rect 505 34676 539 34710
rect 697 34676 731 34710
rect 889 34676 923 34710
rect 1081 34676 1115 34710
rect 1273 34676 1307 34710
rect 1387 34688 1421 34719
rect 1387 34685 1421 34688
rect 3691 34902 3725 34936
rect 2466 34791 2500 34825
rect 2562 34791 2596 34825
rect 2658 34791 2692 34825
rect 2754 34791 2788 34825
rect 2850 34791 2884 34825
rect 2946 34791 2980 34825
rect 3042 34791 3076 34825
rect 3138 34791 3172 34825
rect 3234 34791 3268 34825
rect 3330 34791 3364 34825
rect 3426 34791 3460 34825
rect 3540 34862 3574 34867
rect 3540 34833 3574 34862
rect 3540 34794 3574 34795
rect 3540 34761 3574 34794
rect 3647 34776 3681 34852
rect 3735 34776 3769 34852
rect 2466 34680 2500 34714
rect 2658 34680 2692 34714
rect 2850 34680 2884 34714
rect 3042 34680 3076 34714
rect 3234 34680 3268 34714
rect 3426 34680 3460 34714
rect 3540 34692 3574 34723
rect 3540 34689 3574 34692
rect 3987 34791 4021 34825
rect 4083 34791 4117 34825
rect 4179 34791 4213 34825
rect 4275 34791 4309 34825
rect 4371 34791 4405 34825
rect 4467 34791 4501 34825
rect 4563 34791 4597 34825
rect 4659 34791 4693 34825
rect 4755 34791 4789 34825
rect 4851 34791 4885 34825
rect 4947 34791 4981 34825
rect 5061 34862 5095 34867
rect 5061 34833 5095 34862
rect 5061 34794 5095 34795
rect 5061 34761 5095 34794
rect 5348 34943 5382 34977
rect 5450 34979 5484 34982
rect 5450 34948 5470 34979
rect 5470 34948 5484 34979
rect 3987 34680 4021 34714
rect 4179 34680 4213 34714
rect 4371 34680 4405 34714
rect 4563 34680 4597 34714
rect 4755 34680 4789 34714
rect 4947 34680 4981 34714
rect 5061 34692 5095 34723
rect 5303 34713 5337 34747
rect 5395 34713 5429 34747
rect 5487 34713 5521 34747
rect 5061 34689 5095 34692
rect 313 34197 347 34231
rect 505 34197 539 34231
rect 697 34197 731 34231
rect 889 34197 923 34231
rect 1081 34197 1115 34231
rect 1273 34197 1307 34231
rect 1387 34197 1421 34205
rect 1387 34171 1421 34197
rect 313 34098 347 34102
rect 313 34068 347 34098
rect 313 33996 347 34030
rect 313 33928 347 33958
rect 313 33924 347 33928
rect 409 34098 443 34102
rect 409 34068 443 34098
rect 409 33996 443 34030
rect 409 33928 443 33958
rect 409 33924 443 33928
rect 505 34098 539 34102
rect 505 34068 539 34098
rect 505 33996 539 34030
rect 505 33928 539 33958
rect 505 33924 539 33928
rect 601 34098 635 34102
rect 601 34068 635 34098
rect 601 33996 635 34030
rect 601 33928 635 33958
rect 601 33924 635 33928
rect 697 34098 731 34102
rect 697 34068 731 34098
rect 697 33996 731 34030
rect 697 33928 731 33958
rect 697 33924 731 33928
rect 793 34098 827 34102
rect 793 34068 827 34098
rect 793 33996 827 34030
rect 793 33928 827 33958
rect 793 33924 827 33928
rect 889 34098 923 34102
rect 889 34068 923 34098
rect 889 33996 923 34030
rect 889 33928 923 33958
rect 889 33924 923 33928
rect 985 34098 1019 34102
rect 985 34068 1019 34098
rect 985 33996 1019 34030
rect 985 33928 1019 33958
rect 985 33924 1019 33928
rect 1081 34098 1115 34102
rect 1081 34068 1115 34098
rect 1081 33996 1115 34030
rect 1081 33928 1115 33958
rect 1081 33924 1115 33928
rect 1177 34098 1211 34102
rect 1177 34068 1211 34098
rect 1177 33996 1211 34030
rect 1177 33928 1211 33958
rect 1177 33924 1211 33928
rect 1273 34098 1307 34102
rect 1273 34068 1307 34098
rect 1273 33996 1307 34030
rect 1273 33928 1307 33958
rect 1273 33924 1307 33928
rect 1387 34129 1421 34133
rect 1387 34099 1421 34129
rect 1387 34027 1421 34061
rect 1387 33959 1421 33989
rect 1387 33955 1421 33959
rect 1387 33891 1421 33917
rect 1387 33883 1421 33891
rect 2466 34201 2500 34235
rect 2658 34201 2692 34235
rect 2850 34201 2884 34235
rect 3042 34201 3076 34235
rect 3234 34201 3268 34235
rect 3426 34201 3460 34235
rect 3540 34201 3574 34209
rect 3540 34175 3574 34201
rect 2466 34102 2500 34106
rect 2466 34072 2500 34102
rect 2466 34000 2500 34034
rect 2466 33932 2500 33962
rect 2466 33928 2500 33932
rect 2562 34102 2596 34106
rect 2562 34072 2596 34102
rect 2562 34000 2596 34034
rect 2562 33932 2596 33962
rect 2562 33928 2596 33932
rect 2658 34102 2692 34106
rect 2658 34072 2692 34102
rect 2658 34000 2692 34034
rect 2658 33932 2692 33962
rect 2658 33928 2692 33932
rect 2754 34102 2788 34106
rect 2754 34072 2788 34102
rect 2754 34000 2788 34034
rect 2754 33932 2788 33962
rect 2754 33928 2788 33932
rect 2850 34102 2884 34106
rect 2850 34072 2884 34102
rect 2850 34000 2884 34034
rect 2850 33932 2884 33962
rect 2850 33928 2884 33932
rect 2946 34102 2980 34106
rect 2946 34072 2980 34102
rect 2946 34000 2980 34034
rect 2946 33932 2980 33962
rect 2946 33928 2980 33932
rect 3042 34102 3076 34106
rect 3042 34072 3076 34102
rect 3042 34000 3076 34034
rect 3042 33932 3076 33962
rect 3042 33928 3076 33932
rect 3138 34102 3172 34106
rect 3138 34072 3172 34102
rect 3138 34000 3172 34034
rect 3138 33932 3172 33962
rect 3138 33928 3172 33932
rect 3234 34102 3268 34106
rect 3234 34072 3268 34102
rect 3234 34000 3268 34034
rect 3234 33932 3268 33962
rect 3234 33928 3268 33932
rect 3330 34102 3364 34106
rect 3330 34072 3364 34102
rect 3330 34000 3364 34034
rect 3330 33932 3364 33962
rect 3330 33928 3364 33932
rect 3426 34102 3460 34106
rect 3426 34072 3460 34102
rect 3426 34000 3460 34034
rect 3426 33932 3460 33962
rect 3426 33928 3460 33932
rect 3540 34133 3574 34137
rect 3540 34103 3574 34133
rect 3540 34031 3574 34065
rect 3540 33963 3574 33993
rect 3540 33959 3574 33963
rect 3540 33895 3574 33921
rect 3540 33887 3574 33895
rect 3987 34201 4021 34235
rect 4179 34201 4213 34235
rect 4371 34201 4405 34235
rect 4563 34201 4597 34235
rect 4755 34201 4789 34235
rect 4947 34201 4981 34235
rect 5061 34201 5095 34209
rect 5061 34175 5095 34201
rect 3987 34102 4021 34106
rect 3987 34072 4021 34102
rect 3987 34000 4021 34034
rect 3987 33932 4021 33962
rect 3987 33928 4021 33932
rect 4083 34102 4117 34106
rect 4083 34072 4117 34102
rect 4083 34000 4117 34034
rect 4083 33932 4117 33962
rect 4083 33928 4117 33932
rect 4179 34102 4213 34106
rect 4179 34072 4213 34102
rect 4179 34000 4213 34034
rect 4179 33932 4213 33962
rect 4179 33928 4213 33932
rect 4275 34102 4309 34106
rect 4275 34072 4309 34102
rect 4275 34000 4309 34034
rect 4275 33932 4309 33962
rect 4275 33928 4309 33932
rect 4371 34102 4405 34106
rect 4371 34072 4405 34102
rect 4371 34000 4405 34034
rect 4371 33932 4405 33962
rect 4371 33928 4405 33932
rect 4467 34102 4501 34106
rect 4467 34072 4501 34102
rect 4467 34000 4501 34034
rect 4467 33932 4501 33962
rect 4467 33928 4501 33932
rect 4563 34102 4597 34106
rect 4563 34072 4597 34102
rect 4563 34000 4597 34034
rect 4563 33932 4597 33962
rect 4563 33928 4597 33932
rect 4659 34102 4693 34106
rect 4659 34072 4693 34102
rect 4659 34000 4693 34034
rect 4659 33932 4693 33962
rect 4659 33928 4693 33932
rect 4755 34102 4789 34106
rect 4755 34072 4789 34102
rect 4755 34000 4789 34034
rect 4755 33932 4789 33962
rect 4755 33928 4789 33932
rect 4851 34102 4885 34106
rect 4851 34072 4885 34102
rect 4851 34000 4885 34034
rect 4851 33932 4885 33962
rect 4851 33928 4885 33932
rect 4947 34102 4981 34106
rect 4947 34072 4981 34102
rect 4947 34000 4981 34034
rect 4947 33932 4981 33962
rect 4947 33928 4981 33932
rect 5061 34133 5095 34137
rect 5061 34103 5095 34133
rect 5061 34031 5095 34065
rect 5061 33963 5095 33993
rect 5303 33970 5337 34004
rect 5395 33970 5429 34004
rect 5487 33970 5521 34004
rect 5061 33959 5095 33963
rect 5061 33895 5095 33921
rect 5061 33887 5095 33895
rect 313 33500 347 33534
rect 409 33500 443 33534
rect 505 33500 539 33534
rect 601 33500 635 33534
rect 697 33500 731 33534
rect 793 33500 827 33534
rect 889 33500 923 33534
rect 985 33500 1019 33534
rect 1081 33500 1115 33534
rect 1177 33500 1211 33534
rect 1273 33500 1307 33534
rect 1387 33571 1421 33576
rect 1387 33542 1421 33571
rect 1387 33503 1421 33504
rect 1387 33470 1421 33503
rect 313 33389 347 33423
rect 505 33389 539 33423
rect 697 33389 731 33423
rect 889 33389 923 33423
rect 1081 33389 1115 33423
rect 1273 33389 1307 33423
rect 1387 33401 1421 33432
rect 1387 33398 1421 33401
rect 3691 33615 3725 33649
rect 2466 33504 2500 33538
rect 2562 33504 2596 33538
rect 2658 33504 2692 33538
rect 2754 33504 2788 33538
rect 2850 33504 2884 33538
rect 2946 33504 2980 33538
rect 3042 33504 3076 33538
rect 3138 33504 3172 33538
rect 3234 33504 3268 33538
rect 3330 33504 3364 33538
rect 3426 33504 3460 33538
rect 3540 33575 3574 33580
rect 3540 33546 3574 33575
rect 3540 33507 3574 33508
rect 3540 33474 3574 33507
rect 3647 33489 3681 33565
rect 3735 33489 3769 33565
rect 2466 33393 2500 33427
rect 2658 33393 2692 33427
rect 2850 33393 2884 33427
rect 3042 33393 3076 33427
rect 3234 33393 3268 33427
rect 3426 33393 3460 33427
rect 3540 33405 3574 33436
rect 3540 33402 3574 33405
rect 3987 33504 4021 33538
rect 4083 33504 4117 33538
rect 4179 33504 4213 33538
rect 4275 33504 4309 33538
rect 4371 33504 4405 33538
rect 4467 33504 4501 33538
rect 4563 33504 4597 33538
rect 4659 33504 4693 33538
rect 4755 33504 4789 33538
rect 4851 33504 4885 33538
rect 4947 33504 4981 33538
rect 5061 33575 5095 33580
rect 5061 33546 5095 33575
rect 5061 33507 5095 33508
rect 5061 33474 5095 33507
rect 5348 33656 5382 33690
rect 5450 33692 5484 33695
rect 5450 33661 5470 33692
rect 5470 33661 5484 33692
rect 3987 33393 4021 33427
rect 4179 33393 4213 33427
rect 4371 33393 4405 33427
rect 4563 33393 4597 33427
rect 4755 33393 4789 33427
rect 4947 33393 4981 33427
rect 5061 33405 5095 33436
rect 5303 33426 5337 33460
rect 5395 33426 5429 33460
rect 5487 33426 5521 33460
rect 5061 33402 5095 33405
rect 313 32910 347 32944
rect 505 32910 539 32944
rect 697 32910 731 32944
rect 889 32910 923 32944
rect 1081 32910 1115 32944
rect 1273 32910 1307 32944
rect 1387 32910 1421 32918
rect 1387 32884 1421 32910
rect 313 32811 347 32815
rect 313 32781 347 32811
rect 313 32709 347 32743
rect 313 32641 347 32671
rect 313 32637 347 32641
rect 409 32811 443 32815
rect 409 32781 443 32811
rect 409 32709 443 32743
rect 409 32641 443 32671
rect 409 32637 443 32641
rect 505 32811 539 32815
rect 505 32781 539 32811
rect 505 32709 539 32743
rect 505 32641 539 32671
rect 505 32637 539 32641
rect 601 32811 635 32815
rect 601 32781 635 32811
rect 601 32709 635 32743
rect 601 32641 635 32671
rect 601 32637 635 32641
rect 697 32811 731 32815
rect 697 32781 731 32811
rect 697 32709 731 32743
rect 697 32641 731 32671
rect 697 32637 731 32641
rect 793 32811 827 32815
rect 793 32781 827 32811
rect 793 32709 827 32743
rect 793 32641 827 32671
rect 793 32637 827 32641
rect 889 32811 923 32815
rect 889 32781 923 32811
rect 889 32709 923 32743
rect 889 32641 923 32671
rect 889 32637 923 32641
rect 985 32811 1019 32815
rect 985 32781 1019 32811
rect 985 32709 1019 32743
rect 985 32641 1019 32671
rect 985 32637 1019 32641
rect 1081 32811 1115 32815
rect 1081 32781 1115 32811
rect 1081 32709 1115 32743
rect 1081 32641 1115 32671
rect 1081 32637 1115 32641
rect 1177 32811 1211 32815
rect 1177 32781 1211 32811
rect 1177 32709 1211 32743
rect 1177 32641 1211 32671
rect 1177 32637 1211 32641
rect 1273 32811 1307 32815
rect 1273 32781 1307 32811
rect 1273 32709 1307 32743
rect 1273 32641 1307 32671
rect 1273 32637 1307 32641
rect 1387 32842 1421 32846
rect 1387 32812 1421 32842
rect 1387 32740 1421 32774
rect 1387 32672 1421 32702
rect 1387 32668 1421 32672
rect 1387 32604 1421 32630
rect 1387 32596 1421 32604
rect 2466 32914 2500 32948
rect 2658 32914 2692 32948
rect 2850 32914 2884 32948
rect 3042 32914 3076 32948
rect 3234 32914 3268 32948
rect 3426 32914 3460 32948
rect 3540 32914 3574 32922
rect 3540 32888 3574 32914
rect 2466 32815 2500 32819
rect 2466 32785 2500 32815
rect 2466 32713 2500 32747
rect 2466 32645 2500 32675
rect 2466 32641 2500 32645
rect 2562 32815 2596 32819
rect 2562 32785 2596 32815
rect 2562 32713 2596 32747
rect 2562 32645 2596 32675
rect 2562 32641 2596 32645
rect 2658 32815 2692 32819
rect 2658 32785 2692 32815
rect 2658 32713 2692 32747
rect 2658 32645 2692 32675
rect 2658 32641 2692 32645
rect 2754 32815 2788 32819
rect 2754 32785 2788 32815
rect 2754 32713 2788 32747
rect 2754 32645 2788 32675
rect 2754 32641 2788 32645
rect 2850 32815 2884 32819
rect 2850 32785 2884 32815
rect 2850 32713 2884 32747
rect 2850 32645 2884 32675
rect 2850 32641 2884 32645
rect 2946 32815 2980 32819
rect 2946 32785 2980 32815
rect 2946 32713 2980 32747
rect 2946 32645 2980 32675
rect 2946 32641 2980 32645
rect 3042 32815 3076 32819
rect 3042 32785 3076 32815
rect 3042 32713 3076 32747
rect 3042 32645 3076 32675
rect 3042 32641 3076 32645
rect 3138 32815 3172 32819
rect 3138 32785 3172 32815
rect 3138 32713 3172 32747
rect 3138 32645 3172 32675
rect 3138 32641 3172 32645
rect 3234 32815 3268 32819
rect 3234 32785 3268 32815
rect 3234 32713 3268 32747
rect 3234 32645 3268 32675
rect 3234 32641 3268 32645
rect 3330 32815 3364 32819
rect 3330 32785 3364 32815
rect 3330 32713 3364 32747
rect 3330 32645 3364 32675
rect 3330 32641 3364 32645
rect 3426 32815 3460 32819
rect 3426 32785 3460 32815
rect 3426 32713 3460 32747
rect 3426 32645 3460 32675
rect 3426 32641 3460 32645
rect 3540 32846 3574 32850
rect 3540 32816 3574 32846
rect 3540 32744 3574 32778
rect 3540 32676 3574 32706
rect 3540 32672 3574 32676
rect 3540 32608 3574 32634
rect 3540 32600 3574 32608
rect 3987 32914 4021 32948
rect 4179 32914 4213 32948
rect 4371 32914 4405 32948
rect 4563 32914 4597 32948
rect 4755 32914 4789 32948
rect 4947 32914 4981 32948
rect 5061 32914 5095 32922
rect 5061 32888 5095 32914
rect 3987 32815 4021 32819
rect 3987 32785 4021 32815
rect 3987 32713 4021 32747
rect 3987 32645 4021 32675
rect 3987 32641 4021 32645
rect 4083 32815 4117 32819
rect 4083 32785 4117 32815
rect 4083 32713 4117 32747
rect 4083 32645 4117 32675
rect 4083 32641 4117 32645
rect 4179 32815 4213 32819
rect 4179 32785 4213 32815
rect 4179 32713 4213 32747
rect 4179 32645 4213 32675
rect 4179 32641 4213 32645
rect 4275 32815 4309 32819
rect 4275 32785 4309 32815
rect 4275 32713 4309 32747
rect 4275 32645 4309 32675
rect 4275 32641 4309 32645
rect 4371 32815 4405 32819
rect 4371 32785 4405 32815
rect 4371 32713 4405 32747
rect 4371 32645 4405 32675
rect 4371 32641 4405 32645
rect 4467 32815 4501 32819
rect 4467 32785 4501 32815
rect 4467 32713 4501 32747
rect 4467 32645 4501 32675
rect 4467 32641 4501 32645
rect 4563 32815 4597 32819
rect 4563 32785 4597 32815
rect 4563 32713 4597 32747
rect 4563 32645 4597 32675
rect 4563 32641 4597 32645
rect 4659 32815 4693 32819
rect 4659 32785 4693 32815
rect 4659 32713 4693 32747
rect 4659 32645 4693 32675
rect 4659 32641 4693 32645
rect 4755 32815 4789 32819
rect 4755 32785 4789 32815
rect 4755 32713 4789 32747
rect 4755 32645 4789 32675
rect 4755 32641 4789 32645
rect 4851 32815 4885 32819
rect 4851 32785 4885 32815
rect 4851 32713 4885 32747
rect 4851 32645 4885 32675
rect 4851 32641 4885 32645
rect 4947 32815 4981 32819
rect 4947 32785 4981 32815
rect 4947 32713 4981 32747
rect 4947 32645 4981 32675
rect 4947 32641 4981 32645
rect 5061 32846 5095 32850
rect 5061 32816 5095 32846
rect 5061 32744 5095 32778
rect 5061 32676 5095 32706
rect 5303 32683 5337 32717
rect 5395 32683 5429 32717
rect 5487 32683 5521 32717
rect 5061 32672 5095 32676
rect 5061 32608 5095 32634
rect 5061 32600 5095 32608
rect 313 32213 347 32247
rect 409 32213 443 32247
rect 505 32213 539 32247
rect 601 32213 635 32247
rect 697 32213 731 32247
rect 793 32213 827 32247
rect 889 32213 923 32247
rect 985 32213 1019 32247
rect 1081 32213 1115 32247
rect 1177 32213 1211 32247
rect 1273 32213 1307 32247
rect 1387 32284 1421 32289
rect 1387 32255 1421 32284
rect 1387 32216 1421 32217
rect 1387 32183 1421 32216
rect 313 32102 347 32136
rect 505 32102 539 32136
rect 697 32102 731 32136
rect 889 32102 923 32136
rect 1081 32102 1115 32136
rect 1273 32102 1307 32136
rect 1387 32114 1421 32145
rect 1387 32111 1421 32114
rect 3691 32328 3725 32362
rect 2466 32217 2500 32251
rect 2562 32217 2596 32251
rect 2658 32217 2692 32251
rect 2754 32217 2788 32251
rect 2850 32217 2884 32251
rect 2946 32217 2980 32251
rect 3042 32217 3076 32251
rect 3138 32217 3172 32251
rect 3234 32217 3268 32251
rect 3330 32217 3364 32251
rect 3426 32217 3460 32251
rect 3540 32288 3574 32293
rect 3540 32259 3574 32288
rect 3540 32220 3574 32221
rect 3540 32187 3574 32220
rect 3647 32202 3681 32278
rect 3735 32202 3769 32278
rect 2466 32106 2500 32140
rect 2658 32106 2692 32140
rect 2850 32106 2884 32140
rect 3042 32106 3076 32140
rect 3234 32106 3268 32140
rect 3426 32106 3460 32140
rect 3540 32118 3574 32149
rect 3540 32115 3574 32118
rect 3987 32217 4021 32251
rect 4083 32217 4117 32251
rect 4179 32217 4213 32251
rect 4275 32217 4309 32251
rect 4371 32217 4405 32251
rect 4467 32217 4501 32251
rect 4563 32217 4597 32251
rect 4659 32217 4693 32251
rect 4755 32217 4789 32251
rect 4851 32217 4885 32251
rect 4947 32217 4981 32251
rect 5061 32288 5095 32293
rect 5061 32259 5095 32288
rect 5061 32220 5095 32221
rect 5061 32187 5095 32220
rect 5348 32369 5382 32403
rect 5450 32405 5484 32408
rect 5450 32374 5470 32405
rect 5470 32374 5484 32405
rect 3987 32106 4021 32140
rect 4179 32106 4213 32140
rect 4371 32106 4405 32140
rect 4563 32106 4597 32140
rect 4755 32106 4789 32140
rect 4947 32106 4981 32140
rect 5061 32118 5095 32149
rect 5303 32139 5337 32173
rect 5395 32139 5429 32173
rect 5487 32139 5521 32173
rect 5061 32115 5095 32118
rect 313 31623 347 31657
rect 505 31623 539 31657
rect 697 31623 731 31657
rect 889 31623 923 31657
rect 1081 31623 1115 31657
rect 1273 31623 1307 31657
rect 1387 31623 1421 31631
rect 1387 31597 1421 31623
rect 313 31524 347 31528
rect 313 31494 347 31524
rect 313 31422 347 31456
rect 313 31354 347 31384
rect 313 31350 347 31354
rect 409 31524 443 31528
rect 409 31494 443 31524
rect 409 31422 443 31456
rect 409 31354 443 31384
rect 409 31350 443 31354
rect 505 31524 539 31528
rect 505 31494 539 31524
rect 505 31422 539 31456
rect 505 31354 539 31384
rect 505 31350 539 31354
rect 601 31524 635 31528
rect 601 31494 635 31524
rect 601 31422 635 31456
rect 601 31354 635 31384
rect 601 31350 635 31354
rect 697 31524 731 31528
rect 697 31494 731 31524
rect 697 31422 731 31456
rect 697 31354 731 31384
rect 697 31350 731 31354
rect 793 31524 827 31528
rect 793 31494 827 31524
rect 793 31422 827 31456
rect 793 31354 827 31384
rect 793 31350 827 31354
rect 889 31524 923 31528
rect 889 31494 923 31524
rect 889 31422 923 31456
rect 889 31354 923 31384
rect 889 31350 923 31354
rect 985 31524 1019 31528
rect 985 31494 1019 31524
rect 985 31422 1019 31456
rect 985 31354 1019 31384
rect 985 31350 1019 31354
rect 1081 31524 1115 31528
rect 1081 31494 1115 31524
rect 1081 31422 1115 31456
rect 1081 31354 1115 31384
rect 1081 31350 1115 31354
rect 1177 31524 1211 31528
rect 1177 31494 1211 31524
rect 1177 31422 1211 31456
rect 1177 31354 1211 31384
rect 1177 31350 1211 31354
rect 1273 31524 1307 31528
rect 1273 31494 1307 31524
rect 1273 31422 1307 31456
rect 1273 31354 1307 31384
rect 1273 31350 1307 31354
rect 1387 31555 1421 31559
rect 1387 31525 1421 31555
rect 1387 31453 1421 31487
rect 1387 31385 1421 31415
rect 1387 31381 1421 31385
rect 1387 31317 1421 31343
rect 1387 31309 1421 31317
rect 2466 31627 2500 31661
rect 2658 31627 2692 31661
rect 2850 31627 2884 31661
rect 3042 31627 3076 31661
rect 3234 31627 3268 31661
rect 3426 31627 3460 31661
rect 3540 31627 3574 31635
rect 3540 31601 3574 31627
rect 2466 31528 2500 31532
rect 2466 31498 2500 31528
rect 2466 31426 2500 31460
rect 2466 31358 2500 31388
rect 2466 31354 2500 31358
rect 2562 31528 2596 31532
rect 2562 31498 2596 31528
rect 2562 31426 2596 31460
rect 2562 31358 2596 31388
rect 2562 31354 2596 31358
rect 2658 31528 2692 31532
rect 2658 31498 2692 31528
rect 2658 31426 2692 31460
rect 2658 31358 2692 31388
rect 2658 31354 2692 31358
rect 2754 31528 2788 31532
rect 2754 31498 2788 31528
rect 2754 31426 2788 31460
rect 2754 31358 2788 31388
rect 2754 31354 2788 31358
rect 2850 31528 2884 31532
rect 2850 31498 2884 31528
rect 2850 31426 2884 31460
rect 2850 31358 2884 31388
rect 2850 31354 2884 31358
rect 2946 31528 2980 31532
rect 2946 31498 2980 31528
rect 2946 31426 2980 31460
rect 2946 31358 2980 31388
rect 2946 31354 2980 31358
rect 3042 31528 3076 31532
rect 3042 31498 3076 31528
rect 3042 31426 3076 31460
rect 3042 31358 3076 31388
rect 3042 31354 3076 31358
rect 3138 31528 3172 31532
rect 3138 31498 3172 31528
rect 3138 31426 3172 31460
rect 3138 31358 3172 31388
rect 3138 31354 3172 31358
rect 3234 31528 3268 31532
rect 3234 31498 3268 31528
rect 3234 31426 3268 31460
rect 3234 31358 3268 31388
rect 3234 31354 3268 31358
rect 3330 31528 3364 31532
rect 3330 31498 3364 31528
rect 3330 31426 3364 31460
rect 3330 31358 3364 31388
rect 3330 31354 3364 31358
rect 3426 31528 3460 31532
rect 3426 31498 3460 31528
rect 3426 31426 3460 31460
rect 3426 31358 3460 31388
rect 3426 31354 3460 31358
rect 3540 31559 3574 31563
rect 3540 31529 3574 31559
rect 3540 31457 3574 31491
rect 3540 31389 3574 31419
rect 3540 31385 3574 31389
rect 3540 31321 3574 31347
rect 3540 31313 3574 31321
rect 3987 31627 4021 31661
rect 4179 31627 4213 31661
rect 4371 31627 4405 31661
rect 4563 31627 4597 31661
rect 4755 31627 4789 31661
rect 4947 31627 4981 31661
rect 5061 31627 5095 31635
rect 5061 31601 5095 31627
rect 3987 31528 4021 31532
rect 3987 31498 4021 31528
rect 3987 31426 4021 31460
rect 3987 31358 4021 31388
rect 3987 31354 4021 31358
rect 4083 31528 4117 31532
rect 4083 31498 4117 31528
rect 4083 31426 4117 31460
rect 4083 31358 4117 31388
rect 4083 31354 4117 31358
rect 4179 31528 4213 31532
rect 4179 31498 4213 31528
rect 4179 31426 4213 31460
rect 4179 31358 4213 31388
rect 4179 31354 4213 31358
rect 4275 31528 4309 31532
rect 4275 31498 4309 31528
rect 4275 31426 4309 31460
rect 4275 31358 4309 31388
rect 4275 31354 4309 31358
rect 4371 31528 4405 31532
rect 4371 31498 4405 31528
rect 4371 31426 4405 31460
rect 4371 31358 4405 31388
rect 4371 31354 4405 31358
rect 4467 31528 4501 31532
rect 4467 31498 4501 31528
rect 4467 31426 4501 31460
rect 4467 31358 4501 31388
rect 4467 31354 4501 31358
rect 4563 31528 4597 31532
rect 4563 31498 4597 31528
rect 4563 31426 4597 31460
rect 4563 31358 4597 31388
rect 4563 31354 4597 31358
rect 4659 31528 4693 31532
rect 4659 31498 4693 31528
rect 4659 31426 4693 31460
rect 4659 31358 4693 31388
rect 4659 31354 4693 31358
rect 4755 31528 4789 31532
rect 4755 31498 4789 31528
rect 4755 31426 4789 31460
rect 4755 31358 4789 31388
rect 4755 31354 4789 31358
rect 4851 31528 4885 31532
rect 4851 31498 4885 31528
rect 4851 31426 4885 31460
rect 4851 31358 4885 31388
rect 4851 31354 4885 31358
rect 4947 31528 4981 31532
rect 4947 31498 4981 31528
rect 4947 31426 4981 31460
rect 4947 31358 4981 31388
rect 4947 31354 4981 31358
rect 5061 31559 5095 31563
rect 5061 31529 5095 31559
rect 5061 31457 5095 31491
rect 5061 31389 5095 31419
rect 5303 31396 5337 31430
rect 5395 31396 5429 31430
rect 5487 31396 5521 31430
rect 5061 31385 5095 31389
rect 5061 31321 5095 31347
rect 5061 31313 5095 31321
rect 313 30926 347 30960
rect 409 30926 443 30960
rect 505 30926 539 30960
rect 601 30926 635 30960
rect 697 30926 731 30960
rect 793 30926 827 30960
rect 889 30926 923 30960
rect 985 30926 1019 30960
rect 1081 30926 1115 30960
rect 1177 30926 1211 30960
rect 1273 30926 1307 30960
rect 1387 30997 1421 31002
rect 1387 30968 1421 30997
rect 1387 30929 1421 30930
rect 1387 30896 1421 30929
rect 313 30815 347 30849
rect 505 30815 539 30849
rect 697 30815 731 30849
rect 889 30815 923 30849
rect 1081 30815 1115 30849
rect 1273 30815 1307 30849
rect 1387 30827 1421 30858
rect 1387 30824 1421 30827
rect 3691 31041 3725 31075
rect 2466 30930 2500 30964
rect 2562 30930 2596 30964
rect 2658 30930 2692 30964
rect 2754 30930 2788 30964
rect 2850 30930 2884 30964
rect 2946 30930 2980 30964
rect 3042 30930 3076 30964
rect 3138 30930 3172 30964
rect 3234 30930 3268 30964
rect 3330 30930 3364 30964
rect 3426 30930 3460 30964
rect 3540 31001 3574 31006
rect 3540 30972 3574 31001
rect 3540 30933 3574 30934
rect 3540 30900 3574 30933
rect 3647 30915 3681 30991
rect 3735 30915 3769 30991
rect 2466 30819 2500 30853
rect 2658 30819 2692 30853
rect 2850 30819 2884 30853
rect 3042 30819 3076 30853
rect 3234 30819 3268 30853
rect 3426 30819 3460 30853
rect 3540 30831 3574 30862
rect 3540 30828 3574 30831
rect 3987 30930 4021 30964
rect 4083 30930 4117 30964
rect 4179 30930 4213 30964
rect 4275 30930 4309 30964
rect 4371 30930 4405 30964
rect 4467 30930 4501 30964
rect 4563 30930 4597 30964
rect 4659 30930 4693 30964
rect 4755 30930 4789 30964
rect 4851 30930 4885 30964
rect 4947 30930 4981 30964
rect 5061 31001 5095 31006
rect 5061 30972 5095 31001
rect 5061 30933 5095 30934
rect 5061 30900 5095 30933
rect 5348 31082 5382 31116
rect 5450 31118 5484 31121
rect 5450 31087 5470 31118
rect 5470 31087 5484 31118
rect 3987 30819 4021 30853
rect 4179 30819 4213 30853
rect 4371 30819 4405 30853
rect 4563 30819 4597 30853
rect 4755 30819 4789 30853
rect 4947 30819 4981 30853
rect 5061 30831 5095 30862
rect 5303 30852 5337 30886
rect 5395 30852 5429 30886
rect 5487 30852 5521 30886
rect 5061 30828 5095 30831
rect 313 30336 347 30370
rect 505 30336 539 30370
rect 697 30336 731 30370
rect 889 30336 923 30370
rect 1081 30336 1115 30370
rect 1273 30336 1307 30370
rect 1387 30336 1421 30344
rect 1387 30310 1421 30336
rect 313 30237 347 30241
rect 313 30207 347 30237
rect 313 30135 347 30169
rect 313 30067 347 30097
rect 313 30063 347 30067
rect 409 30237 443 30241
rect 409 30207 443 30237
rect 409 30135 443 30169
rect 409 30067 443 30097
rect 409 30063 443 30067
rect 505 30237 539 30241
rect 505 30207 539 30237
rect 505 30135 539 30169
rect 505 30067 539 30097
rect 505 30063 539 30067
rect 601 30237 635 30241
rect 601 30207 635 30237
rect 601 30135 635 30169
rect 601 30067 635 30097
rect 601 30063 635 30067
rect 697 30237 731 30241
rect 697 30207 731 30237
rect 697 30135 731 30169
rect 697 30067 731 30097
rect 697 30063 731 30067
rect 793 30237 827 30241
rect 793 30207 827 30237
rect 793 30135 827 30169
rect 793 30067 827 30097
rect 793 30063 827 30067
rect 889 30237 923 30241
rect 889 30207 923 30237
rect 889 30135 923 30169
rect 889 30067 923 30097
rect 889 30063 923 30067
rect 985 30237 1019 30241
rect 985 30207 1019 30237
rect 985 30135 1019 30169
rect 985 30067 1019 30097
rect 985 30063 1019 30067
rect 1081 30237 1115 30241
rect 1081 30207 1115 30237
rect 1081 30135 1115 30169
rect 1081 30067 1115 30097
rect 1081 30063 1115 30067
rect 1177 30237 1211 30241
rect 1177 30207 1211 30237
rect 1177 30135 1211 30169
rect 1177 30067 1211 30097
rect 1177 30063 1211 30067
rect 1273 30237 1307 30241
rect 1273 30207 1307 30237
rect 1273 30135 1307 30169
rect 1273 30067 1307 30097
rect 1273 30063 1307 30067
rect 1387 30268 1421 30272
rect 1387 30238 1421 30268
rect 1387 30166 1421 30200
rect 1387 30098 1421 30128
rect 1387 30094 1421 30098
rect 1387 30030 1421 30056
rect 1387 30022 1421 30030
rect 2466 30340 2500 30374
rect 2658 30340 2692 30374
rect 2850 30340 2884 30374
rect 3042 30340 3076 30374
rect 3234 30340 3268 30374
rect 3426 30340 3460 30374
rect 3540 30340 3574 30348
rect 3540 30314 3574 30340
rect 2466 30241 2500 30245
rect 2466 30211 2500 30241
rect 2466 30139 2500 30173
rect 2466 30071 2500 30101
rect 2466 30067 2500 30071
rect 2562 30241 2596 30245
rect 2562 30211 2596 30241
rect 2562 30139 2596 30173
rect 2562 30071 2596 30101
rect 2562 30067 2596 30071
rect 2658 30241 2692 30245
rect 2658 30211 2692 30241
rect 2658 30139 2692 30173
rect 2658 30071 2692 30101
rect 2658 30067 2692 30071
rect 2754 30241 2788 30245
rect 2754 30211 2788 30241
rect 2754 30139 2788 30173
rect 2754 30071 2788 30101
rect 2754 30067 2788 30071
rect 2850 30241 2884 30245
rect 2850 30211 2884 30241
rect 2850 30139 2884 30173
rect 2850 30071 2884 30101
rect 2850 30067 2884 30071
rect 2946 30241 2980 30245
rect 2946 30211 2980 30241
rect 2946 30139 2980 30173
rect 2946 30071 2980 30101
rect 2946 30067 2980 30071
rect 3042 30241 3076 30245
rect 3042 30211 3076 30241
rect 3042 30139 3076 30173
rect 3042 30071 3076 30101
rect 3042 30067 3076 30071
rect 3138 30241 3172 30245
rect 3138 30211 3172 30241
rect 3138 30139 3172 30173
rect 3138 30071 3172 30101
rect 3138 30067 3172 30071
rect 3234 30241 3268 30245
rect 3234 30211 3268 30241
rect 3234 30139 3268 30173
rect 3234 30071 3268 30101
rect 3234 30067 3268 30071
rect 3330 30241 3364 30245
rect 3330 30211 3364 30241
rect 3330 30139 3364 30173
rect 3330 30071 3364 30101
rect 3330 30067 3364 30071
rect 3426 30241 3460 30245
rect 3426 30211 3460 30241
rect 3426 30139 3460 30173
rect 3426 30071 3460 30101
rect 3426 30067 3460 30071
rect 3540 30272 3574 30276
rect 3540 30242 3574 30272
rect 3540 30170 3574 30204
rect 3540 30102 3574 30132
rect 3540 30098 3574 30102
rect 3540 30034 3574 30060
rect 3540 30026 3574 30034
rect 3987 30340 4021 30374
rect 4179 30340 4213 30374
rect 4371 30340 4405 30374
rect 4563 30340 4597 30374
rect 4755 30340 4789 30374
rect 4947 30340 4981 30374
rect 5061 30340 5095 30348
rect 5061 30314 5095 30340
rect 3987 30241 4021 30245
rect 3987 30211 4021 30241
rect 3987 30139 4021 30173
rect 3987 30071 4021 30101
rect 3987 30067 4021 30071
rect 4083 30241 4117 30245
rect 4083 30211 4117 30241
rect 4083 30139 4117 30173
rect 4083 30071 4117 30101
rect 4083 30067 4117 30071
rect 4179 30241 4213 30245
rect 4179 30211 4213 30241
rect 4179 30139 4213 30173
rect 4179 30071 4213 30101
rect 4179 30067 4213 30071
rect 4275 30241 4309 30245
rect 4275 30211 4309 30241
rect 4275 30139 4309 30173
rect 4275 30071 4309 30101
rect 4275 30067 4309 30071
rect 4371 30241 4405 30245
rect 4371 30211 4405 30241
rect 4371 30139 4405 30173
rect 4371 30071 4405 30101
rect 4371 30067 4405 30071
rect 4467 30241 4501 30245
rect 4467 30211 4501 30241
rect 4467 30139 4501 30173
rect 4467 30071 4501 30101
rect 4467 30067 4501 30071
rect 4563 30241 4597 30245
rect 4563 30211 4597 30241
rect 4563 30139 4597 30173
rect 4563 30071 4597 30101
rect 4563 30067 4597 30071
rect 4659 30241 4693 30245
rect 4659 30211 4693 30241
rect 4659 30139 4693 30173
rect 4659 30071 4693 30101
rect 4659 30067 4693 30071
rect 4755 30241 4789 30245
rect 4755 30211 4789 30241
rect 4755 30139 4789 30173
rect 4755 30071 4789 30101
rect 4755 30067 4789 30071
rect 4851 30241 4885 30245
rect 4851 30211 4885 30241
rect 4851 30139 4885 30173
rect 4851 30071 4885 30101
rect 4851 30067 4885 30071
rect 4947 30241 4981 30245
rect 4947 30211 4981 30241
rect 4947 30139 4981 30173
rect 4947 30071 4981 30101
rect 4947 30067 4981 30071
rect 5061 30272 5095 30276
rect 5061 30242 5095 30272
rect 5061 30170 5095 30204
rect 5061 30102 5095 30132
rect 5303 30109 5337 30143
rect 5395 30109 5429 30143
rect 5487 30109 5521 30143
rect 5061 30098 5095 30102
rect 5061 30034 5095 30060
rect 5061 30026 5095 30034
rect 313 29639 347 29673
rect 409 29639 443 29673
rect 505 29639 539 29673
rect 601 29639 635 29673
rect 697 29639 731 29673
rect 793 29639 827 29673
rect 889 29639 923 29673
rect 985 29639 1019 29673
rect 1081 29639 1115 29673
rect 1177 29639 1211 29673
rect 1273 29639 1307 29673
rect 1387 29710 1421 29715
rect 1387 29681 1421 29710
rect 1387 29642 1421 29643
rect 1387 29609 1421 29642
rect 313 29528 347 29562
rect 505 29528 539 29562
rect 697 29528 731 29562
rect 889 29528 923 29562
rect 1081 29528 1115 29562
rect 1273 29528 1307 29562
rect 1387 29540 1421 29571
rect 1387 29537 1421 29540
rect 3691 29754 3725 29788
rect 2466 29643 2500 29677
rect 2562 29643 2596 29677
rect 2658 29643 2692 29677
rect 2754 29643 2788 29677
rect 2850 29643 2884 29677
rect 2946 29643 2980 29677
rect 3042 29643 3076 29677
rect 3138 29643 3172 29677
rect 3234 29643 3268 29677
rect 3330 29643 3364 29677
rect 3426 29643 3460 29677
rect 3540 29714 3574 29719
rect 3540 29685 3574 29714
rect 3540 29646 3574 29647
rect 3540 29613 3574 29646
rect 3647 29628 3681 29704
rect 3735 29628 3769 29704
rect 2466 29532 2500 29566
rect 2658 29532 2692 29566
rect 2850 29532 2884 29566
rect 3042 29532 3076 29566
rect 3234 29532 3268 29566
rect 3426 29532 3460 29566
rect 3540 29544 3574 29575
rect 3540 29541 3574 29544
rect 3987 29643 4021 29677
rect 4083 29643 4117 29677
rect 4179 29643 4213 29677
rect 4275 29643 4309 29677
rect 4371 29643 4405 29677
rect 4467 29643 4501 29677
rect 4563 29643 4597 29677
rect 4659 29643 4693 29677
rect 4755 29643 4789 29677
rect 4851 29643 4885 29677
rect 4947 29643 4981 29677
rect 5061 29714 5095 29719
rect 5061 29685 5095 29714
rect 5061 29646 5095 29647
rect 5061 29613 5095 29646
rect 5348 29795 5382 29829
rect 5450 29831 5484 29834
rect 5450 29800 5470 29831
rect 5470 29800 5484 29831
rect 3987 29532 4021 29566
rect 4179 29532 4213 29566
rect 4371 29532 4405 29566
rect 4563 29532 4597 29566
rect 4755 29532 4789 29566
rect 4947 29532 4981 29566
rect 5061 29544 5095 29575
rect 5303 29565 5337 29599
rect 5395 29565 5429 29599
rect 5487 29565 5521 29599
rect 5061 29541 5095 29544
rect 313 29049 347 29083
rect 505 29049 539 29083
rect 697 29049 731 29083
rect 889 29049 923 29083
rect 1081 29049 1115 29083
rect 1273 29049 1307 29083
rect 1387 29049 1421 29057
rect 1387 29023 1421 29049
rect 313 28950 347 28954
rect 313 28920 347 28950
rect 313 28848 347 28882
rect 313 28780 347 28810
rect 313 28776 347 28780
rect 409 28950 443 28954
rect 409 28920 443 28950
rect 409 28848 443 28882
rect 409 28780 443 28810
rect 409 28776 443 28780
rect 505 28950 539 28954
rect 505 28920 539 28950
rect 505 28848 539 28882
rect 505 28780 539 28810
rect 505 28776 539 28780
rect 601 28950 635 28954
rect 601 28920 635 28950
rect 601 28848 635 28882
rect 601 28780 635 28810
rect 601 28776 635 28780
rect 697 28950 731 28954
rect 697 28920 731 28950
rect 697 28848 731 28882
rect 697 28780 731 28810
rect 697 28776 731 28780
rect 793 28950 827 28954
rect 793 28920 827 28950
rect 793 28848 827 28882
rect 793 28780 827 28810
rect 793 28776 827 28780
rect 889 28950 923 28954
rect 889 28920 923 28950
rect 889 28848 923 28882
rect 889 28780 923 28810
rect 889 28776 923 28780
rect 985 28950 1019 28954
rect 985 28920 1019 28950
rect 985 28848 1019 28882
rect 985 28780 1019 28810
rect 985 28776 1019 28780
rect 1081 28950 1115 28954
rect 1081 28920 1115 28950
rect 1081 28848 1115 28882
rect 1081 28780 1115 28810
rect 1081 28776 1115 28780
rect 1177 28950 1211 28954
rect 1177 28920 1211 28950
rect 1177 28848 1211 28882
rect 1177 28780 1211 28810
rect 1177 28776 1211 28780
rect 1273 28950 1307 28954
rect 1273 28920 1307 28950
rect 1273 28848 1307 28882
rect 1273 28780 1307 28810
rect 1273 28776 1307 28780
rect 1387 28981 1421 28985
rect 1387 28951 1421 28981
rect 1387 28879 1421 28913
rect 1387 28811 1421 28841
rect 1387 28807 1421 28811
rect 1387 28743 1421 28769
rect 1387 28735 1421 28743
rect 2466 29053 2500 29087
rect 2658 29053 2692 29087
rect 2850 29053 2884 29087
rect 3042 29053 3076 29087
rect 3234 29053 3268 29087
rect 3426 29053 3460 29087
rect 3540 29053 3574 29061
rect 3540 29027 3574 29053
rect 2466 28954 2500 28958
rect 2466 28924 2500 28954
rect 2466 28852 2500 28886
rect 2466 28784 2500 28814
rect 2466 28780 2500 28784
rect 2562 28954 2596 28958
rect 2562 28924 2596 28954
rect 2562 28852 2596 28886
rect 2562 28784 2596 28814
rect 2562 28780 2596 28784
rect 2658 28954 2692 28958
rect 2658 28924 2692 28954
rect 2658 28852 2692 28886
rect 2658 28784 2692 28814
rect 2658 28780 2692 28784
rect 2754 28954 2788 28958
rect 2754 28924 2788 28954
rect 2754 28852 2788 28886
rect 2754 28784 2788 28814
rect 2754 28780 2788 28784
rect 2850 28954 2884 28958
rect 2850 28924 2884 28954
rect 2850 28852 2884 28886
rect 2850 28784 2884 28814
rect 2850 28780 2884 28784
rect 2946 28954 2980 28958
rect 2946 28924 2980 28954
rect 2946 28852 2980 28886
rect 2946 28784 2980 28814
rect 2946 28780 2980 28784
rect 3042 28954 3076 28958
rect 3042 28924 3076 28954
rect 3042 28852 3076 28886
rect 3042 28784 3076 28814
rect 3042 28780 3076 28784
rect 3138 28954 3172 28958
rect 3138 28924 3172 28954
rect 3138 28852 3172 28886
rect 3138 28784 3172 28814
rect 3138 28780 3172 28784
rect 3234 28954 3268 28958
rect 3234 28924 3268 28954
rect 3234 28852 3268 28886
rect 3234 28784 3268 28814
rect 3234 28780 3268 28784
rect 3330 28954 3364 28958
rect 3330 28924 3364 28954
rect 3330 28852 3364 28886
rect 3330 28784 3364 28814
rect 3330 28780 3364 28784
rect 3426 28954 3460 28958
rect 3426 28924 3460 28954
rect 3426 28852 3460 28886
rect 3426 28784 3460 28814
rect 3426 28780 3460 28784
rect 3540 28985 3574 28989
rect 3540 28955 3574 28985
rect 3540 28883 3574 28917
rect 3540 28815 3574 28845
rect 3540 28811 3574 28815
rect 3540 28747 3574 28773
rect 3540 28739 3574 28747
rect 3987 29053 4021 29087
rect 4179 29053 4213 29087
rect 4371 29053 4405 29087
rect 4563 29053 4597 29087
rect 4755 29053 4789 29087
rect 4947 29053 4981 29087
rect 5061 29053 5095 29061
rect 5061 29027 5095 29053
rect 3987 28954 4021 28958
rect 3987 28924 4021 28954
rect 3987 28852 4021 28886
rect 3987 28784 4021 28814
rect 3987 28780 4021 28784
rect 4083 28954 4117 28958
rect 4083 28924 4117 28954
rect 4083 28852 4117 28886
rect 4083 28784 4117 28814
rect 4083 28780 4117 28784
rect 4179 28954 4213 28958
rect 4179 28924 4213 28954
rect 4179 28852 4213 28886
rect 4179 28784 4213 28814
rect 4179 28780 4213 28784
rect 4275 28954 4309 28958
rect 4275 28924 4309 28954
rect 4275 28852 4309 28886
rect 4275 28784 4309 28814
rect 4275 28780 4309 28784
rect 4371 28954 4405 28958
rect 4371 28924 4405 28954
rect 4371 28852 4405 28886
rect 4371 28784 4405 28814
rect 4371 28780 4405 28784
rect 4467 28954 4501 28958
rect 4467 28924 4501 28954
rect 4467 28852 4501 28886
rect 4467 28784 4501 28814
rect 4467 28780 4501 28784
rect 4563 28954 4597 28958
rect 4563 28924 4597 28954
rect 4563 28852 4597 28886
rect 4563 28784 4597 28814
rect 4563 28780 4597 28784
rect 4659 28954 4693 28958
rect 4659 28924 4693 28954
rect 4659 28852 4693 28886
rect 4659 28784 4693 28814
rect 4659 28780 4693 28784
rect 4755 28954 4789 28958
rect 4755 28924 4789 28954
rect 4755 28852 4789 28886
rect 4755 28784 4789 28814
rect 4755 28780 4789 28784
rect 4851 28954 4885 28958
rect 4851 28924 4885 28954
rect 4851 28852 4885 28886
rect 4851 28784 4885 28814
rect 4851 28780 4885 28784
rect 4947 28954 4981 28958
rect 4947 28924 4981 28954
rect 4947 28852 4981 28886
rect 4947 28784 4981 28814
rect 4947 28780 4981 28784
rect 5061 28985 5095 28989
rect 5061 28955 5095 28985
rect 5061 28883 5095 28917
rect 5061 28815 5095 28845
rect 5303 28822 5337 28856
rect 5395 28822 5429 28856
rect 5487 28822 5521 28856
rect 5061 28811 5095 28815
rect 5061 28747 5095 28773
rect 5061 28739 5095 28747
rect 313 28352 347 28386
rect 409 28352 443 28386
rect 505 28352 539 28386
rect 601 28352 635 28386
rect 697 28352 731 28386
rect 793 28352 827 28386
rect 889 28352 923 28386
rect 985 28352 1019 28386
rect 1081 28352 1115 28386
rect 1177 28352 1211 28386
rect 1273 28352 1307 28386
rect 1387 28423 1421 28428
rect 1387 28394 1421 28423
rect 1387 28355 1421 28356
rect 1387 28322 1421 28355
rect 313 28241 347 28275
rect 505 28241 539 28275
rect 697 28241 731 28275
rect 889 28241 923 28275
rect 1081 28241 1115 28275
rect 1273 28241 1307 28275
rect 1387 28253 1421 28284
rect 1387 28250 1421 28253
rect 3691 28467 3725 28501
rect 2466 28356 2500 28390
rect 2562 28356 2596 28390
rect 2658 28356 2692 28390
rect 2754 28356 2788 28390
rect 2850 28356 2884 28390
rect 2946 28356 2980 28390
rect 3042 28356 3076 28390
rect 3138 28356 3172 28390
rect 3234 28356 3268 28390
rect 3330 28356 3364 28390
rect 3426 28356 3460 28390
rect 3540 28427 3574 28432
rect 3540 28398 3574 28427
rect 3540 28359 3574 28360
rect 3540 28326 3574 28359
rect 3647 28341 3681 28417
rect 3735 28341 3769 28417
rect 2466 28245 2500 28279
rect 2658 28245 2692 28279
rect 2850 28245 2884 28279
rect 3042 28245 3076 28279
rect 3234 28245 3268 28279
rect 3426 28245 3460 28279
rect 3540 28257 3574 28288
rect 3540 28254 3574 28257
rect 3987 28356 4021 28390
rect 4083 28356 4117 28390
rect 4179 28356 4213 28390
rect 4275 28356 4309 28390
rect 4371 28356 4405 28390
rect 4467 28356 4501 28390
rect 4563 28356 4597 28390
rect 4659 28356 4693 28390
rect 4755 28356 4789 28390
rect 4851 28356 4885 28390
rect 4947 28356 4981 28390
rect 5061 28427 5095 28432
rect 5061 28398 5095 28427
rect 5061 28359 5095 28360
rect 5061 28326 5095 28359
rect 5348 28508 5382 28542
rect 5450 28544 5484 28547
rect 5450 28513 5470 28544
rect 5470 28513 5484 28544
rect 3987 28245 4021 28279
rect 4179 28245 4213 28279
rect 4371 28245 4405 28279
rect 4563 28245 4597 28279
rect 4755 28245 4789 28279
rect 4947 28245 4981 28279
rect 5061 28257 5095 28288
rect 5303 28278 5337 28312
rect 5395 28278 5429 28312
rect 5487 28278 5521 28312
rect 5061 28254 5095 28257
rect 313 27762 347 27796
rect 505 27762 539 27796
rect 697 27762 731 27796
rect 889 27762 923 27796
rect 1081 27762 1115 27796
rect 1273 27762 1307 27796
rect 1387 27762 1421 27770
rect 1387 27736 1421 27762
rect 313 27663 347 27667
rect 313 27633 347 27663
rect 313 27561 347 27595
rect 313 27493 347 27523
rect 313 27489 347 27493
rect 409 27663 443 27667
rect 409 27633 443 27663
rect 409 27561 443 27595
rect 409 27493 443 27523
rect 409 27489 443 27493
rect 505 27663 539 27667
rect 505 27633 539 27663
rect 505 27561 539 27595
rect 505 27493 539 27523
rect 505 27489 539 27493
rect 601 27663 635 27667
rect 601 27633 635 27663
rect 601 27561 635 27595
rect 601 27493 635 27523
rect 601 27489 635 27493
rect 697 27663 731 27667
rect 697 27633 731 27663
rect 697 27561 731 27595
rect 697 27493 731 27523
rect 697 27489 731 27493
rect 793 27663 827 27667
rect 793 27633 827 27663
rect 793 27561 827 27595
rect 793 27493 827 27523
rect 793 27489 827 27493
rect 889 27663 923 27667
rect 889 27633 923 27663
rect 889 27561 923 27595
rect 889 27493 923 27523
rect 889 27489 923 27493
rect 985 27663 1019 27667
rect 985 27633 1019 27663
rect 985 27561 1019 27595
rect 985 27493 1019 27523
rect 985 27489 1019 27493
rect 1081 27663 1115 27667
rect 1081 27633 1115 27663
rect 1081 27561 1115 27595
rect 1081 27493 1115 27523
rect 1081 27489 1115 27493
rect 1177 27663 1211 27667
rect 1177 27633 1211 27663
rect 1177 27561 1211 27595
rect 1177 27493 1211 27523
rect 1177 27489 1211 27493
rect 1273 27663 1307 27667
rect 1273 27633 1307 27663
rect 1273 27561 1307 27595
rect 1273 27493 1307 27523
rect 1273 27489 1307 27493
rect 1387 27694 1421 27698
rect 1387 27664 1421 27694
rect 1387 27592 1421 27626
rect 1387 27524 1421 27554
rect 1387 27520 1421 27524
rect 1387 27456 1421 27482
rect 1387 27448 1421 27456
rect 2466 27766 2500 27800
rect 2658 27766 2692 27800
rect 2850 27766 2884 27800
rect 3042 27766 3076 27800
rect 3234 27766 3268 27800
rect 3426 27766 3460 27800
rect 3540 27766 3574 27774
rect 3540 27740 3574 27766
rect 2466 27667 2500 27671
rect 2466 27637 2500 27667
rect 2466 27565 2500 27599
rect 2466 27497 2500 27527
rect 2466 27493 2500 27497
rect 2562 27667 2596 27671
rect 2562 27637 2596 27667
rect 2562 27565 2596 27599
rect 2562 27497 2596 27527
rect 2562 27493 2596 27497
rect 2658 27667 2692 27671
rect 2658 27637 2692 27667
rect 2658 27565 2692 27599
rect 2658 27497 2692 27527
rect 2658 27493 2692 27497
rect 2754 27667 2788 27671
rect 2754 27637 2788 27667
rect 2754 27565 2788 27599
rect 2754 27497 2788 27527
rect 2754 27493 2788 27497
rect 2850 27667 2884 27671
rect 2850 27637 2884 27667
rect 2850 27565 2884 27599
rect 2850 27497 2884 27527
rect 2850 27493 2884 27497
rect 2946 27667 2980 27671
rect 2946 27637 2980 27667
rect 2946 27565 2980 27599
rect 2946 27497 2980 27527
rect 2946 27493 2980 27497
rect 3042 27667 3076 27671
rect 3042 27637 3076 27667
rect 3042 27565 3076 27599
rect 3042 27497 3076 27527
rect 3042 27493 3076 27497
rect 3138 27667 3172 27671
rect 3138 27637 3172 27667
rect 3138 27565 3172 27599
rect 3138 27497 3172 27527
rect 3138 27493 3172 27497
rect 3234 27667 3268 27671
rect 3234 27637 3268 27667
rect 3234 27565 3268 27599
rect 3234 27497 3268 27527
rect 3234 27493 3268 27497
rect 3330 27667 3364 27671
rect 3330 27637 3364 27667
rect 3330 27565 3364 27599
rect 3330 27497 3364 27527
rect 3330 27493 3364 27497
rect 3426 27667 3460 27671
rect 3426 27637 3460 27667
rect 3426 27565 3460 27599
rect 3426 27497 3460 27527
rect 3426 27493 3460 27497
rect 3540 27698 3574 27702
rect 3540 27668 3574 27698
rect 3540 27596 3574 27630
rect 3540 27528 3574 27558
rect 3540 27524 3574 27528
rect 3540 27460 3574 27486
rect 3540 27452 3574 27460
rect 3987 27766 4021 27800
rect 4179 27766 4213 27800
rect 4371 27766 4405 27800
rect 4563 27766 4597 27800
rect 4755 27766 4789 27800
rect 4947 27766 4981 27800
rect 5061 27766 5095 27774
rect 5061 27740 5095 27766
rect 3987 27667 4021 27671
rect 3987 27637 4021 27667
rect 3987 27565 4021 27599
rect 3987 27497 4021 27527
rect 3987 27493 4021 27497
rect 4083 27667 4117 27671
rect 4083 27637 4117 27667
rect 4083 27565 4117 27599
rect 4083 27497 4117 27527
rect 4083 27493 4117 27497
rect 4179 27667 4213 27671
rect 4179 27637 4213 27667
rect 4179 27565 4213 27599
rect 4179 27497 4213 27527
rect 4179 27493 4213 27497
rect 4275 27667 4309 27671
rect 4275 27637 4309 27667
rect 4275 27565 4309 27599
rect 4275 27497 4309 27527
rect 4275 27493 4309 27497
rect 4371 27667 4405 27671
rect 4371 27637 4405 27667
rect 4371 27565 4405 27599
rect 4371 27497 4405 27527
rect 4371 27493 4405 27497
rect 4467 27667 4501 27671
rect 4467 27637 4501 27667
rect 4467 27565 4501 27599
rect 4467 27497 4501 27527
rect 4467 27493 4501 27497
rect 4563 27667 4597 27671
rect 4563 27637 4597 27667
rect 4563 27565 4597 27599
rect 4563 27497 4597 27527
rect 4563 27493 4597 27497
rect 4659 27667 4693 27671
rect 4659 27637 4693 27667
rect 4659 27565 4693 27599
rect 4659 27497 4693 27527
rect 4659 27493 4693 27497
rect 4755 27667 4789 27671
rect 4755 27637 4789 27667
rect 4755 27565 4789 27599
rect 4755 27497 4789 27527
rect 4755 27493 4789 27497
rect 4851 27667 4885 27671
rect 4851 27637 4885 27667
rect 4851 27565 4885 27599
rect 4851 27497 4885 27527
rect 4851 27493 4885 27497
rect 4947 27667 4981 27671
rect 4947 27637 4981 27667
rect 4947 27565 4981 27599
rect 4947 27497 4981 27527
rect 4947 27493 4981 27497
rect 5061 27698 5095 27702
rect 5061 27668 5095 27698
rect 5061 27596 5095 27630
rect 5061 27528 5095 27558
rect 5303 27535 5337 27569
rect 5395 27535 5429 27569
rect 5487 27535 5521 27569
rect 5061 27524 5095 27528
rect 5061 27460 5095 27486
rect 5061 27452 5095 27460
rect 313 27065 347 27099
rect 409 27065 443 27099
rect 505 27065 539 27099
rect 601 27065 635 27099
rect 697 27065 731 27099
rect 793 27065 827 27099
rect 889 27065 923 27099
rect 985 27065 1019 27099
rect 1081 27065 1115 27099
rect 1177 27065 1211 27099
rect 1273 27065 1307 27099
rect 1387 27136 1421 27141
rect 1387 27107 1421 27136
rect 1387 27068 1421 27069
rect 1387 27035 1421 27068
rect 313 26954 347 26988
rect 505 26954 539 26988
rect 697 26954 731 26988
rect 889 26954 923 26988
rect 1081 26954 1115 26988
rect 1273 26954 1307 26988
rect 1387 26966 1421 26997
rect 1387 26963 1421 26966
rect 3691 27180 3725 27214
rect 2466 27069 2500 27103
rect 2562 27069 2596 27103
rect 2658 27069 2692 27103
rect 2754 27069 2788 27103
rect 2850 27069 2884 27103
rect 2946 27069 2980 27103
rect 3042 27069 3076 27103
rect 3138 27069 3172 27103
rect 3234 27069 3268 27103
rect 3330 27069 3364 27103
rect 3426 27069 3460 27103
rect 3540 27140 3574 27145
rect 3540 27111 3574 27140
rect 3540 27072 3574 27073
rect 3540 27039 3574 27072
rect 3647 27054 3681 27130
rect 3735 27054 3769 27130
rect 2466 26958 2500 26992
rect 2658 26958 2692 26992
rect 2850 26958 2884 26992
rect 3042 26958 3076 26992
rect 3234 26958 3268 26992
rect 3426 26958 3460 26992
rect 3540 26970 3574 27001
rect 3540 26967 3574 26970
rect 3987 27069 4021 27103
rect 4083 27069 4117 27103
rect 4179 27069 4213 27103
rect 4275 27069 4309 27103
rect 4371 27069 4405 27103
rect 4467 27069 4501 27103
rect 4563 27069 4597 27103
rect 4659 27069 4693 27103
rect 4755 27069 4789 27103
rect 4851 27069 4885 27103
rect 4947 27069 4981 27103
rect 5061 27140 5095 27145
rect 5061 27111 5095 27140
rect 5061 27072 5095 27073
rect 5061 27039 5095 27072
rect 5348 27221 5382 27255
rect 5450 27257 5484 27260
rect 5450 27226 5470 27257
rect 5470 27226 5484 27257
rect 3987 26958 4021 26992
rect 4179 26958 4213 26992
rect 4371 26958 4405 26992
rect 4563 26958 4597 26992
rect 4755 26958 4789 26992
rect 4947 26958 4981 26992
rect 5061 26970 5095 27001
rect 5303 26991 5337 27025
rect 5395 26991 5429 27025
rect 5487 26991 5521 27025
rect 5061 26967 5095 26970
rect 313 26475 347 26509
rect 505 26475 539 26509
rect 697 26475 731 26509
rect 889 26475 923 26509
rect 1081 26475 1115 26509
rect 1273 26475 1307 26509
rect 1387 26475 1421 26483
rect 1387 26449 1421 26475
rect 313 26376 347 26380
rect 313 26346 347 26376
rect 313 26274 347 26308
rect 313 26206 347 26236
rect 313 26202 347 26206
rect 409 26376 443 26380
rect 409 26346 443 26376
rect 409 26274 443 26308
rect 409 26206 443 26236
rect 409 26202 443 26206
rect 505 26376 539 26380
rect 505 26346 539 26376
rect 505 26274 539 26308
rect 505 26206 539 26236
rect 505 26202 539 26206
rect 601 26376 635 26380
rect 601 26346 635 26376
rect 601 26274 635 26308
rect 601 26206 635 26236
rect 601 26202 635 26206
rect 697 26376 731 26380
rect 697 26346 731 26376
rect 697 26274 731 26308
rect 697 26206 731 26236
rect 697 26202 731 26206
rect 793 26376 827 26380
rect 793 26346 827 26376
rect 793 26274 827 26308
rect 793 26206 827 26236
rect 793 26202 827 26206
rect 889 26376 923 26380
rect 889 26346 923 26376
rect 889 26274 923 26308
rect 889 26206 923 26236
rect 889 26202 923 26206
rect 985 26376 1019 26380
rect 985 26346 1019 26376
rect 985 26274 1019 26308
rect 985 26206 1019 26236
rect 985 26202 1019 26206
rect 1081 26376 1115 26380
rect 1081 26346 1115 26376
rect 1081 26274 1115 26308
rect 1081 26206 1115 26236
rect 1081 26202 1115 26206
rect 1177 26376 1211 26380
rect 1177 26346 1211 26376
rect 1177 26274 1211 26308
rect 1177 26206 1211 26236
rect 1177 26202 1211 26206
rect 1273 26376 1307 26380
rect 1273 26346 1307 26376
rect 1273 26274 1307 26308
rect 1273 26206 1307 26236
rect 1273 26202 1307 26206
rect 1387 26407 1421 26411
rect 1387 26377 1421 26407
rect 1387 26305 1421 26339
rect 1387 26237 1421 26267
rect 1387 26233 1421 26237
rect 1387 26169 1421 26195
rect 1387 26161 1421 26169
rect 2466 26479 2500 26513
rect 2658 26479 2692 26513
rect 2850 26479 2884 26513
rect 3042 26479 3076 26513
rect 3234 26479 3268 26513
rect 3426 26479 3460 26513
rect 3540 26479 3574 26487
rect 3540 26453 3574 26479
rect 2466 26380 2500 26384
rect 2466 26350 2500 26380
rect 2466 26278 2500 26312
rect 2466 26210 2500 26240
rect 2466 26206 2500 26210
rect 2562 26380 2596 26384
rect 2562 26350 2596 26380
rect 2562 26278 2596 26312
rect 2562 26210 2596 26240
rect 2562 26206 2596 26210
rect 2658 26380 2692 26384
rect 2658 26350 2692 26380
rect 2658 26278 2692 26312
rect 2658 26210 2692 26240
rect 2658 26206 2692 26210
rect 2754 26380 2788 26384
rect 2754 26350 2788 26380
rect 2754 26278 2788 26312
rect 2754 26210 2788 26240
rect 2754 26206 2788 26210
rect 2850 26380 2884 26384
rect 2850 26350 2884 26380
rect 2850 26278 2884 26312
rect 2850 26210 2884 26240
rect 2850 26206 2884 26210
rect 2946 26380 2980 26384
rect 2946 26350 2980 26380
rect 2946 26278 2980 26312
rect 2946 26210 2980 26240
rect 2946 26206 2980 26210
rect 3042 26380 3076 26384
rect 3042 26350 3076 26380
rect 3042 26278 3076 26312
rect 3042 26210 3076 26240
rect 3042 26206 3076 26210
rect 3138 26380 3172 26384
rect 3138 26350 3172 26380
rect 3138 26278 3172 26312
rect 3138 26210 3172 26240
rect 3138 26206 3172 26210
rect 3234 26380 3268 26384
rect 3234 26350 3268 26380
rect 3234 26278 3268 26312
rect 3234 26210 3268 26240
rect 3234 26206 3268 26210
rect 3330 26380 3364 26384
rect 3330 26350 3364 26380
rect 3330 26278 3364 26312
rect 3330 26210 3364 26240
rect 3330 26206 3364 26210
rect 3426 26380 3460 26384
rect 3426 26350 3460 26380
rect 3426 26278 3460 26312
rect 3426 26210 3460 26240
rect 3426 26206 3460 26210
rect 3540 26411 3574 26415
rect 3540 26381 3574 26411
rect 3540 26309 3574 26343
rect 3540 26241 3574 26271
rect 3540 26237 3574 26241
rect 3540 26173 3574 26199
rect 3540 26165 3574 26173
rect 3987 26479 4021 26513
rect 4179 26479 4213 26513
rect 4371 26479 4405 26513
rect 4563 26479 4597 26513
rect 4755 26479 4789 26513
rect 4947 26479 4981 26513
rect 5061 26479 5095 26487
rect 5061 26453 5095 26479
rect 3987 26380 4021 26384
rect 3987 26350 4021 26380
rect 3987 26278 4021 26312
rect 3987 26210 4021 26240
rect 3987 26206 4021 26210
rect 4083 26380 4117 26384
rect 4083 26350 4117 26380
rect 4083 26278 4117 26312
rect 4083 26210 4117 26240
rect 4083 26206 4117 26210
rect 4179 26380 4213 26384
rect 4179 26350 4213 26380
rect 4179 26278 4213 26312
rect 4179 26210 4213 26240
rect 4179 26206 4213 26210
rect 4275 26380 4309 26384
rect 4275 26350 4309 26380
rect 4275 26278 4309 26312
rect 4275 26210 4309 26240
rect 4275 26206 4309 26210
rect 4371 26380 4405 26384
rect 4371 26350 4405 26380
rect 4371 26278 4405 26312
rect 4371 26210 4405 26240
rect 4371 26206 4405 26210
rect 4467 26380 4501 26384
rect 4467 26350 4501 26380
rect 4467 26278 4501 26312
rect 4467 26210 4501 26240
rect 4467 26206 4501 26210
rect 4563 26380 4597 26384
rect 4563 26350 4597 26380
rect 4563 26278 4597 26312
rect 4563 26210 4597 26240
rect 4563 26206 4597 26210
rect 4659 26380 4693 26384
rect 4659 26350 4693 26380
rect 4659 26278 4693 26312
rect 4659 26210 4693 26240
rect 4659 26206 4693 26210
rect 4755 26380 4789 26384
rect 4755 26350 4789 26380
rect 4755 26278 4789 26312
rect 4755 26210 4789 26240
rect 4755 26206 4789 26210
rect 4851 26380 4885 26384
rect 4851 26350 4885 26380
rect 4851 26278 4885 26312
rect 4851 26210 4885 26240
rect 4851 26206 4885 26210
rect 4947 26380 4981 26384
rect 4947 26350 4981 26380
rect 4947 26278 4981 26312
rect 4947 26210 4981 26240
rect 4947 26206 4981 26210
rect 5061 26411 5095 26415
rect 5061 26381 5095 26411
rect 5061 26309 5095 26343
rect 5061 26241 5095 26271
rect 5303 26248 5337 26282
rect 5395 26248 5429 26282
rect 5487 26248 5521 26282
rect 5061 26237 5095 26241
rect 5061 26173 5095 26199
rect 5061 26165 5095 26173
rect 313 25778 347 25812
rect 409 25778 443 25812
rect 505 25778 539 25812
rect 601 25778 635 25812
rect 697 25778 731 25812
rect 793 25778 827 25812
rect 889 25778 923 25812
rect 985 25778 1019 25812
rect 1081 25778 1115 25812
rect 1177 25778 1211 25812
rect 1273 25778 1307 25812
rect 1387 25849 1421 25854
rect 1387 25820 1421 25849
rect 1387 25781 1421 25782
rect 1387 25748 1421 25781
rect 313 25667 347 25701
rect 505 25667 539 25701
rect 697 25667 731 25701
rect 889 25667 923 25701
rect 1081 25667 1115 25701
rect 1273 25667 1307 25701
rect 1387 25679 1421 25710
rect 1387 25676 1421 25679
rect 3691 25893 3725 25927
rect 2466 25782 2500 25816
rect 2562 25782 2596 25816
rect 2658 25782 2692 25816
rect 2754 25782 2788 25816
rect 2850 25782 2884 25816
rect 2946 25782 2980 25816
rect 3042 25782 3076 25816
rect 3138 25782 3172 25816
rect 3234 25782 3268 25816
rect 3330 25782 3364 25816
rect 3426 25782 3460 25816
rect 3540 25853 3574 25858
rect 3540 25824 3574 25853
rect 3540 25785 3574 25786
rect 3540 25752 3574 25785
rect 3647 25767 3681 25843
rect 3735 25767 3769 25843
rect 2466 25671 2500 25705
rect 2658 25671 2692 25705
rect 2850 25671 2884 25705
rect 3042 25671 3076 25705
rect 3234 25671 3268 25705
rect 3426 25671 3460 25705
rect 3540 25683 3574 25714
rect 3540 25680 3574 25683
rect 3987 25782 4021 25816
rect 4083 25782 4117 25816
rect 4179 25782 4213 25816
rect 4275 25782 4309 25816
rect 4371 25782 4405 25816
rect 4467 25782 4501 25816
rect 4563 25782 4597 25816
rect 4659 25782 4693 25816
rect 4755 25782 4789 25816
rect 4851 25782 4885 25816
rect 4947 25782 4981 25816
rect 5061 25853 5095 25858
rect 5061 25824 5095 25853
rect 5061 25785 5095 25786
rect 5061 25752 5095 25785
rect 5348 25934 5382 25968
rect 5450 25970 5484 25973
rect 5450 25939 5470 25970
rect 5470 25939 5484 25970
rect 3987 25671 4021 25705
rect 4179 25671 4213 25705
rect 4371 25671 4405 25705
rect 4563 25671 4597 25705
rect 4755 25671 4789 25705
rect 4947 25671 4981 25705
rect 5061 25683 5095 25714
rect 5303 25704 5337 25738
rect 5395 25704 5429 25738
rect 5487 25704 5521 25738
rect 5061 25680 5095 25683
rect 313 25188 347 25222
rect 505 25188 539 25222
rect 697 25188 731 25222
rect 889 25188 923 25222
rect 1081 25188 1115 25222
rect 1273 25188 1307 25222
rect 1387 25188 1421 25196
rect 1387 25162 1421 25188
rect 313 25089 347 25093
rect 313 25059 347 25089
rect 313 24987 347 25021
rect 313 24919 347 24949
rect 313 24915 347 24919
rect 409 25089 443 25093
rect 409 25059 443 25089
rect 409 24987 443 25021
rect 409 24919 443 24949
rect 409 24915 443 24919
rect 505 25089 539 25093
rect 505 25059 539 25089
rect 505 24987 539 25021
rect 505 24919 539 24949
rect 505 24915 539 24919
rect 601 25089 635 25093
rect 601 25059 635 25089
rect 601 24987 635 25021
rect 601 24919 635 24949
rect 601 24915 635 24919
rect 697 25089 731 25093
rect 697 25059 731 25089
rect 697 24987 731 25021
rect 697 24919 731 24949
rect 697 24915 731 24919
rect 793 25089 827 25093
rect 793 25059 827 25089
rect 793 24987 827 25021
rect 793 24919 827 24949
rect 793 24915 827 24919
rect 889 25089 923 25093
rect 889 25059 923 25089
rect 889 24987 923 25021
rect 889 24919 923 24949
rect 889 24915 923 24919
rect 985 25089 1019 25093
rect 985 25059 1019 25089
rect 985 24987 1019 25021
rect 985 24919 1019 24949
rect 985 24915 1019 24919
rect 1081 25089 1115 25093
rect 1081 25059 1115 25089
rect 1081 24987 1115 25021
rect 1081 24919 1115 24949
rect 1081 24915 1115 24919
rect 1177 25089 1211 25093
rect 1177 25059 1211 25089
rect 1177 24987 1211 25021
rect 1177 24919 1211 24949
rect 1177 24915 1211 24919
rect 1273 25089 1307 25093
rect 1273 25059 1307 25089
rect 1273 24987 1307 25021
rect 1273 24919 1307 24949
rect 1273 24915 1307 24919
rect 1387 25120 1421 25124
rect 1387 25090 1421 25120
rect 1387 25018 1421 25052
rect 1387 24950 1421 24980
rect 1387 24946 1421 24950
rect 1387 24882 1421 24908
rect 1387 24874 1421 24882
rect 2466 25192 2500 25226
rect 2658 25192 2692 25226
rect 2850 25192 2884 25226
rect 3042 25192 3076 25226
rect 3234 25192 3268 25226
rect 3426 25192 3460 25226
rect 3540 25192 3574 25200
rect 3540 25166 3574 25192
rect 2466 25093 2500 25097
rect 2466 25063 2500 25093
rect 2466 24991 2500 25025
rect 2466 24923 2500 24953
rect 2466 24919 2500 24923
rect 2562 25093 2596 25097
rect 2562 25063 2596 25093
rect 2562 24991 2596 25025
rect 2562 24923 2596 24953
rect 2562 24919 2596 24923
rect 2658 25093 2692 25097
rect 2658 25063 2692 25093
rect 2658 24991 2692 25025
rect 2658 24923 2692 24953
rect 2658 24919 2692 24923
rect 2754 25093 2788 25097
rect 2754 25063 2788 25093
rect 2754 24991 2788 25025
rect 2754 24923 2788 24953
rect 2754 24919 2788 24923
rect 2850 25093 2884 25097
rect 2850 25063 2884 25093
rect 2850 24991 2884 25025
rect 2850 24923 2884 24953
rect 2850 24919 2884 24923
rect 2946 25093 2980 25097
rect 2946 25063 2980 25093
rect 2946 24991 2980 25025
rect 2946 24923 2980 24953
rect 2946 24919 2980 24923
rect 3042 25093 3076 25097
rect 3042 25063 3076 25093
rect 3042 24991 3076 25025
rect 3042 24923 3076 24953
rect 3042 24919 3076 24923
rect 3138 25093 3172 25097
rect 3138 25063 3172 25093
rect 3138 24991 3172 25025
rect 3138 24923 3172 24953
rect 3138 24919 3172 24923
rect 3234 25093 3268 25097
rect 3234 25063 3268 25093
rect 3234 24991 3268 25025
rect 3234 24923 3268 24953
rect 3234 24919 3268 24923
rect 3330 25093 3364 25097
rect 3330 25063 3364 25093
rect 3330 24991 3364 25025
rect 3330 24923 3364 24953
rect 3330 24919 3364 24923
rect 3426 25093 3460 25097
rect 3426 25063 3460 25093
rect 3426 24991 3460 25025
rect 3426 24923 3460 24953
rect 3426 24919 3460 24923
rect 3540 25124 3574 25128
rect 3540 25094 3574 25124
rect 3540 25022 3574 25056
rect 3540 24954 3574 24984
rect 3540 24950 3574 24954
rect 3540 24886 3574 24912
rect 3540 24878 3574 24886
rect 3987 25192 4021 25226
rect 4179 25192 4213 25226
rect 4371 25192 4405 25226
rect 4563 25192 4597 25226
rect 4755 25192 4789 25226
rect 4947 25192 4981 25226
rect 5061 25192 5095 25200
rect 5061 25166 5095 25192
rect 3987 25093 4021 25097
rect 3987 25063 4021 25093
rect 3987 24991 4021 25025
rect 3987 24923 4021 24953
rect 3987 24919 4021 24923
rect 4083 25093 4117 25097
rect 4083 25063 4117 25093
rect 4083 24991 4117 25025
rect 4083 24923 4117 24953
rect 4083 24919 4117 24923
rect 4179 25093 4213 25097
rect 4179 25063 4213 25093
rect 4179 24991 4213 25025
rect 4179 24923 4213 24953
rect 4179 24919 4213 24923
rect 4275 25093 4309 25097
rect 4275 25063 4309 25093
rect 4275 24991 4309 25025
rect 4275 24923 4309 24953
rect 4275 24919 4309 24923
rect 4371 25093 4405 25097
rect 4371 25063 4405 25093
rect 4371 24991 4405 25025
rect 4371 24923 4405 24953
rect 4371 24919 4405 24923
rect 4467 25093 4501 25097
rect 4467 25063 4501 25093
rect 4467 24991 4501 25025
rect 4467 24923 4501 24953
rect 4467 24919 4501 24923
rect 4563 25093 4597 25097
rect 4563 25063 4597 25093
rect 4563 24991 4597 25025
rect 4563 24923 4597 24953
rect 4563 24919 4597 24923
rect 4659 25093 4693 25097
rect 4659 25063 4693 25093
rect 4659 24991 4693 25025
rect 4659 24923 4693 24953
rect 4659 24919 4693 24923
rect 4755 25093 4789 25097
rect 4755 25063 4789 25093
rect 4755 24991 4789 25025
rect 4755 24923 4789 24953
rect 4755 24919 4789 24923
rect 4851 25093 4885 25097
rect 4851 25063 4885 25093
rect 4851 24991 4885 25025
rect 4851 24923 4885 24953
rect 4851 24919 4885 24923
rect 4947 25093 4981 25097
rect 4947 25063 4981 25093
rect 4947 24991 4981 25025
rect 4947 24923 4981 24953
rect 4947 24919 4981 24923
rect 5061 25124 5095 25128
rect 5061 25094 5095 25124
rect 5061 25022 5095 25056
rect 5061 24954 5095 24984
rect 5303 24961 5337 24995
rect 5395 24961 5429 24995
rect 5487 24961 5521 24995
rect 5061 24950 5095 24954
rect 5061 24886 5095 24912
rect 5061 24878 5095 24886
rect 313 24491 347 24525
rect 409 24491 443 24525
rect 505 24491 539 24525
rect 601 24491 635 24525
rect 697 24491 731 24525
rect 793 24491 827 24525
rect 889 24491 923 24525
rect 985 24491 1019 24525
rect 1081 24491 1115 24525
rect 1177 24491 1211 24525
rect 1273 24491 1307 24525
rect 1387 24562 1421 24567
rect 1387 24533 1421 24562
rect 1387 24494 1421 24495
rect 1387 24461 1421 24494
rect 313 24380 347 24414
rect 505 24380 539 24414
rect 697 24380 731 24414
rect 889 24380 923 24414
rect 1081 24380 1115 24414
rect 1273 24380 1307 24414
rect 1387 24392 1421 24423
rect 1387 24389 1421 24392
rect 3691 24606 3725 24640
rect 2466 24495 2500 24529
rect 2562 24495 2596 24529
rect 2658 24495 2692 24529
rect 2754 24495 2788 24529
rect 2850 24495 2884 24529
rect 2946 24495 2980 24529
rect 3042 24495 3076 24529
rect 3138 24495 3172 24529
rect 3234 24495 3268 24529
rect 3330 24495 3364 24529
rect 3426 24495 3460 24529
rect 3540 24566 3574 24571
rect 3540 24537 3574 24566
rect 3540 24498 3574 24499
rect 3540 24465 3574 24498
rect 3647 24480 3681 24556
rect 3735 24480 3769 24556
rect 2466 24384 2500 24418
rect 2658 24384 2692 24418
rect 2850 24384 2884 24418
rect 3042 24384 3076 24418
rect 3234 24384 3268 24418
rect 3426 24384 3460 24418
rect 3540 24396 3574 24427
rect 3540 24393 3574 24396
rect 3987 24495 4021 24529
rect 4083 24495 4117 24529
rect 4179 24495 4213 24529
rect 4275 24495 4309 24529
rect 4371 24495 4405 24529
rect 4467 24495 4501 24529
rect 4563 24495 4597 24529
rect 4659 24495 4693 24529
rect 4755 24495 4789 24529
rect 4851 24495 4885 24529
rect 4947 24495 4981 24529
rect 5061 24566 5095 24571
rect 5061 24537 5095 24566
rect 5061 24498 5095 24499
rect 5061 24465 5095 24498
rect 5348 24647 5382 24681
rect 5450 24683 5484 24686
rect 5450 24652 5470 24683
rect 5470 24652 5484 24683
rect 3987 24384 4021 24418
rect 4179 24384 4213 24418
rect 4371 24384 4405 24418
rect 4563 24384 4597 24418
rect 4755 24384 4789 24418
rect 4947 24384 4981 24418
rect 5061 24396 5095 24427
rect 5303 24417 5337 24451
rect 5395 24417 5429 24451
rect 5487 24417 5521 24451
rect 5061 24393 5095 24396
rect 313 23901 347 23935
rect 505 23901 539 23935
rect 697 23901 731 23935
rect 889 23901 923 23935
rect 1081 23901 1115 23935
rect 1273 23901 1307 23935
rect 1387 23901 1421 23909
rect 1387 23875 1421 23901
rect 313 23802 347 23806
rect 313 23772 347 23802
rect 313 23700 347 23734
rect 313 23632 347 23662
rect 313 23628 347 23632
rect 409 23802 443 23806
rect 409 23772 443 23802
rect 409 23700 443 23734
rect 409 23632 443 23662
rect 409 23628 443 23632
rect 505 23802 539 23806
rect 505 23772 539 23802
rect 505 23700 539 23734
rect 505 23632 539 23662
rect 505 23628 539 23632
rect 601 23802 635 23806
rect 601 23772 635 23802
rect 601 23700 635 23734
rect 601 23632 635 23662
rect 601 23628 635 23632
rect 697 23802 731 23806
rect 697 23772 731 23802
rect 697 23700 731 23734
rect 697 23632 731 23662
rect 697 23628 731 23632
rect 793 23802 827 23806
rect 793 23772 827 23802
rect 793 23700 827 23734
rect 793 23632 827 23662
rect 793 23628 827 23632
rect 889 23802 923 23806
rect 889 23772 923 23802
rect 889 23700 923 23734
rect 889 23632 923 23662
rect 889 23628 923 23632
rect 985 23802 1019 23806
rect 985 23772 1019 23802
rect 985 23700 1019 23734
rect 985 23632 1019 23662
rect 985 23628 1019 23632
rect 1081 23802 1115 23806
rect 1081 23772 1115 23802
rect 1081 23700 1115 23734
rect 1081 23632 1115 23662
rect 1081 23628 1115 23632
rect 1177 23802 1211 23806
rect 1177 23772 1211 23802
rect 1177 23700 1211 23734
rect 1177 23632 1211 23662
rect 1177 23628 1211 23632
rect 1273 23802 1307 23806
rect 1273 23772 1307 23802
rect 1273 23700 1307 23734
rect 1273 23632 1307 23662
rect 1273 23628 1307 23632
rect 1387 23833 1421 23837
rect 1387 23803 1421 23833
rect 1387 23731 1421 23765
rect 1387 23663 1421 23693
rect 1387 23659 1421 23663
rect 1387 23595 1421 23621
rect 1387 23587 1421 23595
rect 2466 23905 2500 23939
rect 2658 23905 2692 23939
rect 2850 23905 2884 23939
rect 3042 23905 3076 23939
rect 3234 23905 3268 23939
rect 3426 23905 3460 23939
rect 3540 23905 3574 23913
rect 3540 23879 3574 23905
rect 2466 23806 2500 23810
rect 2466 23776 2500 23806
rect 2466 23704 2500 23738
rect 2466 23636 2500 23666
rect 2466 23632 2500 23636
rect 2562 23806 2596 23810
rect 2562 23776 2596 23806
rect 2562 23704 2596 23738
rect 2562 23636 2596 23666
rect 2562 23632 2596 23636
rect 2658 23806 2692 23810
rect 2658 23776 2692 23806
rect 2658 23704 2692 23738
rect 2658 23636 2692 23666
rect 2658 23632 2692 23636
rect 2754 23806 2788 23810
rect 2754 23776 2788 23806
rect 2754 23704 2788 23738
rect 2754 23636 2788 23666
rect 2754 23632 2788 23636
rect 2850 23806 2884 23810
rect 2850 23776 2884 23806
rect 2850 23704 2884 23738
rect 2850 23636 2884 23666
rect 2850 23632 2884 23636
rect 2946 23806 2980 23810
rect 2946 23776 2980 23806
rect 2946 23704 2980 23738
rect 2946 23636 2980 23666
rect 2946 23632 2980 23636
rect 3042 23806 3076 23810
rect 3042 23776 3076 23806
rect 3042 23704 3076 23738
rect 3042 23636 3076 23666
rect 3042 23632 3076 23636
rect 3138 23806 3172 23810
rect 3138 23776 3172 23806
rect 3138 23704 3172 23738
rect 3138 23636 3172 23666
rect 3138 23632 3172 23636
rect 3234 23806 3268 23810
rect 3234 23776 3268 23806
rect 3234 23704 3268 23738
rect 3234 23636 3268 23666
rect 3234 23632 3268 23636
rect 3330 23806 3364 23810
rect 3330 23776 3364 23806
rect 3330 23704 3364 23738
rect 3330 23636 3364 23666
rect 3330 23632 3364 23636
rect 3426 23806 3460 23810
rect 3426 23776 3460 23806
rect 3426 23704 3460 23738
rect 3426 23636 3460 23666
rect 3426 23632 3460 23636
rect 3540 23837 3574 23841
rect 3540 23807 3574 23837
rect 3540 23735 3574 23769
rect 3540 23667 3574 23697
rect 3540 23663 3574 23667
rect 3540 23599 3574 23625
rect 3540 23591 3574 23599
rect 3987 23905 4021 23939
rect 4179 23905 4213 23939
rect 4371 23905 4405 23939
rect 4563 23905 4597 23939
rect 4755 23905 4789 23939
rect 4947 23905 4981 23939
rect 5061 23905 5095 23913
rect 5061 23879 5095 23905
rect 3987 23806 4021 23810
rect 3987 23776 4021 23806
rect 3987 23704 4021 23738
rect 3987 23636 4021 23666
rect 3987 23632 4021 23636
rect 4083 23806 4117 23810
rect 4083 23776 4117 23806
rect 4083 23704 4117 23738
rect 4083 23636 4117 23666
rect 4083 23632 4117 23636
rect 4179 23806 4213 23810
rect 4179 23776 4213 23806
rect 4179 23704 4213 23738
rect 4179 23636 4213 23666
rect 4179 23632 4213 23636
rect 4275 23806 4309 23810
rect 4275 23776 4309 23806
rect 4275 23704 4309 23738
rect 4275 23636 4309 23666
rect 4275 23632 4309 23636
rect 4371 23806 4405 23810
rect 4371 23776 4405 23806
rect 4371 23704 4405 23738
rect 4371 23636 4405 23666
rect 4371 23632 4405 23636
rect 4467 23806 4501 23810
rect 4467 23776 4501 23806
rect 4467 23704 4501 23738
rect 4467 23636 4501 23666
rect 4467 23632 4501 23636
rect 4563 23806 4597 23810
rect 4563 23776 4597 23806
rect 4563 23704 4597 23738
rect 4563 23636 4597 23666
rect 4563 23632 4597 23636
rect 4659 23806 4693 23810
rect 4659 23776 4693 23806
rect 4659 23704 4693 23738
rect 4659 23636 4693 23666
rect 4659 23632 4693 23636
rect 4755 23806 4789 23810
rect 4755 23776 4789 23806
rect 4755 23704 4789 23738
rect 4755 23636 4789 23666
rect 4755 23632 4789 23636
rect 4851 23806 4885 23810
rect 4851 23776 4885 23806
rect 4851 23704 4885 23738
rect 4851 23636 4885 23666
rect 4851 23632 4885 23636
rect 4947 23806 4981 23810
rect 4947 23776 4981 23806
rect 4947 23704 4981 23738
rect 4947 23636 4981 23666
rect 4947 23632 4981 23636
rect 5061 23837 5095 23841
rect 5061 23807 5095 23837
rect 5061 23735 5095 23769
rect 5061 23667 5095 23697
rect 5303 23674 5337 23708
rect 5395 23674 5429 23708
rect 5487 23674 5521 23708
rect 5061 23663 5095 23667
rect 5061 23599 5095 23625
rect 5061 23591 5095 23599
rect 313 23204 347 23238
rect 409 23204 443 23238
rect 505 23204 539 23238
rect 601 23204 635 23238
rect 697 23204 731 23238
rect 793 23204 827 23238
rect 889 23204 923 23238
rect 985 23204 1019 23238
rect 1081 23204 1115 23238
rect 1177 23204 1211 23238
rect 1273 23204 1307 23238
rect 1387 23275 1421 23280
rect 1387 23246 1421 23275
rect 1387 23207 1421 23208
rect 1387 23174 1421 23207
rect 313 23093 347 23127
rect 505 23093 539 23127
rect 697 23093 731 23127
rect 889 23093 923 23127
rect 1081 23093 1115 23127
rect 1273 23093 1307 23127
rect 1387 23105 1421 23136
rect 1387 23102 1421 23105
rect 3691 23319 3725 23353
rect 2466 23208 2500 23242
rect 2562 23208 2596 23242
rect 2658 23208 2692 23242
rect 2754 23208 2788 23242
rect 2850 23208 2884 23242
rect 2946 23208 2980 23242
rect 3042 23208 3076 23242
rect 3138 23208 3172 23242
rect 3234 23208 3268 23242
rect 3330 23208 3364 23242
rect 3426 23208 3460 23242
rect 3540 23279 3574 23284
rect 3540 23250 3574 23279
rect 3540 23211 3574 23212
rect 3540 23178 3574 23211
rect 3647 23193 3681 23269
rect 3735 23193 3769 23269
rect 2466 23097 2500 23131
rect 2658 23097 2692 23131
rect 2850 23097 2884 23131
rect 3042 23097 3076 23131
rect 3234 23097 3268 23131
rect 3426 23097 3460 23131
rect 3540 23109 3574 23140
rect 3540 23106 3574 23109
rect 3987 23208 4021 23242
rect 4083 23208 4117 23242
rect 4179 23208 4213 23242
rect 4275 23208 4309 23242
rect 4371 23208 4405 23242
rect 4467 23208 4501 23242
rect 4563 23208 4597 23242
rect 4659 23208 4693 23242
rect 4755 23208 4789 23242
rect 4851 23208 4885 23242
rect 4947 23208 4981 23242
rect 5061 23279 5095 23284
rect 5061 23250 5095 23279
rect 5061 23211 5095 23212
rect 5061 23178 5095 23211
rect 5348 23360 5382 23394
rect 5450 23396 5484 23399
rect 5450 23365 5470 23396
rect 5470 23365 5484 23396
rect 3987 23097 4021 23131
rect 4179 23097 4213 23131
rect 4371 23097 4405 23131
rect 4563 23097 4597 23131
rect 4755 23097 4789 23131
rect 4947 23097 4981 23131
rect 5061 23109 5095 23140
rect 5303 23130 5337 23164
rect 5395 23130 5429 23164
rect 5487 23130 5521 23164
rect 5061 23106 5095 23109
rect 313 22614 347 22648
rect 505 22614 539 22648
rect 697 22614 731 22648
rect 889 22614 923 22648
rect 1081 22614 1115 22648
rect 1273 22614 1307 22648
rect 1387 22614 1421 22622
rect 1387 22588 1421 22614
rect 313 22515 347 22519
rect 313 22485 347 22515
rect 313 22413 347 22447
rect 313 22345 347 22375
rect 313 22341 347 22345
rect 409 22515 443 22519
rect 409 22485 443 22515
rect 409 22413 443 22447
rect 409 22345 443 22375
rect 409 22341 443 22345
rect 505 22515 539 22519
rect 505 22485 539 22515
rect 505 22413 539 22447
rect 505 22345 539 22375
rect 505 22341 539 22345
rect 601 22515 635 22519
rect 601 22485 635 22515
rect 601 22413 635 22447
rect 601 22345 635 22375
rect 601 22341 635 22345
rect 697 22515 731 22519
rect 697 22485 731 22515
rect 697 22413 731 22447
rect 697 22345 731 22375
rect 697 22341 731 22345
rect 793 22515 827 22519
rect 793 22485 827 22515
rect 793 22413 827 22447
rect 793 22345 827 22375
rect 793 22341 827 22345
rect 889 22515 923 22519
rect 889 22485 923 22515
rect 889 22413 923 22447
rect 889 22345 923 22375
rect 889 22341 923 22345
rect 985 22515 1019 22519
rect 985 22485 1019 22515
rect 985 22413 1019 22447
rect 985 22345 1019 22375
rect 985 22341 1019 22345
rect 1081 22515 1115 22519
rect 1081 22485 1115 22515
rect 1081 22413 1115 22447
rect 1081 22345 1115 22375
rect 1081 22341 1115 22345
rect 1177 22515 1211 22519
rect 1177 22485 1211 22515
rect 1177 22413 1211 22447
rect 1177 22345 1211 22375
rect 1177 22341 1211 22345
rect 1273 22515 1307 22519
rect 1273 22485 1307 22515
rect 1273 22413 1307 22447
rect 1273 22345 1307 22375
rect 1273 22341 1307 22345
rect 1387 22546 1421 22550
rect 1387 22516 1421 22546
rect 1387 22444 1421 22478
rect 1387 22376 1421 22406
rect 1387 22372 1421 22376
rect 1387 22308 1421 22334
rect 1387 22300 1421 22308
rect 2466 22618 2500 22652
rect 2658 22618 2692 22652
rect 2850 22618 2884 22652
rect 3042 22618 3076 22652
rect 3234 22618 3268 22652
rect 3426 22618 3460 22652
rect 3540 22618 3574 22626
rect 3540 22592 3574 22618
rect 2466 22519 2500 22523
rect 2466 22489 2500 22519
rect 2466 22417 2500 22451
rect 2466 22349 2500 22379
rect 2466 22345 2500 22349
rect 2562 22519 2596 22523
rect 2562 22489 2596 22519
rect 2562 22417 2596 22451
rect 2562 22349 2596 22379
rect 2562 22345 2596 22349
rect 2658 22519 2692 22523
rect 2658 22489 2692 22519
rect 2658 22417 2692 22451
rect 2658 22349 2692 22379
rect 2658 22345 2692 22349
rect 2754 22519 2788 22523
rect 2754 22489 2788 22519
rect 2754 22417 2788 22451
rect 2754 22349 2788 22379
rect 2754 22345 2788 22349
rect 2850 22519 2884 22523
rect 2850 22489 2884 22519
rect 2850 22417 2884 22451
rect 2850 22349 2884 22379
rect 2850 22345 2884 22349
rect 2946 22519 2980 22523
rect 2946 22489 2980 22519
rect 2946 22417 2980 22451
rect 2946 22349 2980 22379
rect 2946 22345 2980 22349
rect 3042 22519 3076 22523
rect 3042 22489 3076 22519
rect 3042 22417 3076 22451
rect 3042 22349 3076 22379
rect 3042 22345 3076 22349
rect 3138 22519 3172 22523
rect 3138 22489 3172 22519
rect 3138 22417 3172 22451
rect 3138 22349 3172 22379
rect 3138 22345 3172 22349
rect 3234 22519 3268 22523
rect 3234 22489 3268 22519
rect 3234 22417 3268 22451
rect 3234 22349 3268 22379
rect 3234 22345 3268 22349
rect 3330 22519 3364 22523
rect 3330 22489 3364 22519
rect 3330 22417 3364 22451
rect 3330 22349 3364 22379
rect 3330 22345 3364 22349
rect 3426 22519 3460 22523
rect 3426 22489 3460 22519
rect 3426 22417 3460 22451
rect 3426 22349 3460 22379
rect 3426 22345 3460 22349
rect 3540 22550 3574 22554
rect 3540 22520 3574 22550
rect 3540 22448 3574 22482
rect 3540 22380 3574 22410
rect 3540 22376 3574 22380
rect 3540 22312 3574 22338
rect 3540 22304 3574 22312
rect 3987 22618 4021 22652
rect 4179 22618 4213 22652
rect 4371 22618 4405 22652
rect 4563 22618 4597 22652
rect 4755 22618 4789 22652
rect 4947 22618 4981 22652
rect 5061 22618 5095 22626
rect 5061 22592 5095 22618
rect 3987 22519 4021 22523
rect 3987 22489 4021 22519
rect 3987 22417 4021 22451
rect 3987 22349 4021 22379
rect 3987 22345 4021 22349
rect 4083 22519 4117 22523
rect 4083 22489 4117 22519
rect 4083 22417 4117 22451
rect 4083 22349 4117 22379
rect 4083 22345 4117 22349
rect 4179 22519 4213 22523
rect 4179 22489 4213 22519
rect 4179 22417 4213 22451
rect 4179 22349 4213 22379
rect 4179 22345 4213 22349
rect 4275 22519 4309 22523
rect 4275 22489 4309 22519
rect 4275 22417 4309 22451
rect 4275 22349 4309 22379
rect 4275 22345 4309 22349
rect 4371 22519 4405 22523
rect 4371 22489 4405 22519
rect 4371 22417 4405 22451
rect 4371 22349 4405 22379
rect 4371 22345 4405 22349
rect 4467 22519 4501 22523
rect 4467 22489 4501 22519
rect 4467 22417 4501 22451
rect 4467 22349 4501 22379
rect 4467 22345 4501 22349
rect 4563 22519 4597 22523
rect 4563 22489 4597 22519
rect 4563 22417 4597 22451
rect 4563 22349 4597 22379
rect 4563 22345 4597 22349
rect 4659 22519 4693 22523
rect 4659 22489 4693 22519
rect 4659 22417 4693 22451
rect 4659 22349 4693 22379
rect 4659 22345 4693 22349
rect 4755 22519 4789 22523
rect 4755 22489 4789 22519
rect 4755 22417 4789 22451
rect 4755 22349 4789 22379
rect 4755 22345 4789 22349
rect 4851 22519 4885 22523
rect 4851 22489 4885 22519
rect 4851 22417 4885 22451
rect 4851 22349 4885 22379
rect 4851 22345 4885 22349
rect 4947 22519 4981 22523
rect 4947 22489 4981 22519
rect 4947 22417 4981 22451
rect 4947 22349 4981 22379
rect 4947 22345 4981 22349
rect 5061 22550 5095 22554
rect 5061 22520 5095 22550
rect 5061 22448 5095 22482
rect 5061 22380 5095 22410
rect 5303 22387 5337 22421
rect 5395 22387 5429 22421
rect 5487 22387 5521 22421
rect 5061 22376 5095 22380
rect 5061 22312 5095 22338
rect 5061 22304 5095 22312
rect 313 21917 347 21951
rect 409 21917 443 21951
rect 505 21917 539 21951
rect 601 21917 635 21951
rect 697 21917 731 21951
rect 793 21917 827 21951
rect 889 21917 923 21951
rect 985 21917 1019 21951
rect 1081 21917 1115 21951
rect 1177 21917 1211 21951
rect 1273 21917 1307 21951
rect 1387 21988 1421 21993
rect 1387 21959 1421 21988
rect 1387 21920 1421 21921
rect 1387 21887 1421 21920
rect 313 21806 347 21840
rect 505 21806 539 21840
rect 697 21806 731 21840
rect 889 21806 923 21840
rect 1081 21806 1115 21840
rect 1273 21806 1307 21840
rect 1387 21818 1421 21849
rect 1387 21815 1421 21818
rect 3691 22032 3725 22066
rect 2466 21921 2500 21955
rect 2562 21921 2596 21955
rect 2658 21921 2692 21955
rect 2754 21921 2788 21955
rect 2850 21921 2884 21955
rect 2946 21921 2980 21955
rect 3042 21921 3076 21955
rect 3138 21921 3172 21955
rect 3234 21921 3268 21955
rect 3330 21921 3364 21955
rect 3426 21921 3460 21955
rect 3540 21992 3574 21997
rect 3540 21963 3574 21992
rect 3540 21924 3574 21925
rect 3540 21891 3574 21924
rect 3647 21906 3681 21982
rect 3735 21906 3769 21982
rect 2466 21810 2500 21844
rect 2658 21810 2692 21844
rect 2850 21810 2884 21844
rect 3042 21810 3076 21844
rect 3234 21810 3268 21844
rect 3426 21810 3460 21844
rect 3540 21822 3574 21853
rect 3540 21819 3574 21822
rect 3987 21921 4021 21955
rect 4083 21921 4117 21955
rect 4179 21921 4213 21955
rect 4275 21921 4309 21955
rect 4371 21921 4405 21955
rect 4467 21921 4501 21955
rect 4563 21921 4597 21955
rect 4659 21921 4693 21955
rect 4755 21921 4789 21955
rect 4851 21921 4885 21955
rect 4947 21921 4981 21955
rect 5061 21992 5095 21997
rect 5061 21963 5095 21992
rect 5061 21924 5095 21925
rect 5061 21891 5095 21924
rect 5348 22073 5382 22107
rect 5450 22109 5484 22112
rect 5450 22078 5470 22109
rect 5470 22078 5484 22109
rect 3987 21810 4021 21844
rect 4179 21810 4213 21844
rect 4371 21810 4405 21844
rect 4563 21810 4597 21844
rect 4755 21810 4789 21844
rect 4947 21810 4981 21844
rect 5061 21822 5095 21853
rect 5303 21843 5337 21877
rect 5395 21843 5429 21877
rect 5487 21843 5521 21877
rect 5061 21819 5095 21822
rect 313 21327 347 21361
rect 505 21327 539 21361
rect 697 21327 731 21361
rect 889 21327 923 21361
rect 1081 21327 1115 21361
rect 1273 21327 1307 21361
rect 1387 21327 1421 21335
rect 1387 21301 1421 21327
rect 313 21228 347 21232
rect 313 21198 347 21228
rect 313 21126 347 21160
rect 313 21058 347 21088
rect 313 21054 347 21058
rect 409 21228 443 21232
rect 409 21198 443 21228
rect 409 21126 443 21160
rect 409 21058 443 21088
rect 409 21054 443 21058
rect 505 21228 539 21232
rect 505 21198 539 21228
rect 505 21126 539 21160
rect 505 21058 539 21088
rect 505 21054 539 21058
rect 601 21228 635 21232
rect 601 21198 635 21228
rect 601 21126 635 21160
rect 601 21058 635 21088
rect 601 21054 635 21058
rect 697 21228 731 21232
rect 697 21198 731 21228
rect 697 21126 731 21160
rect 697 21058 731 21088
rect 697 21054 731 21058
rect 793 21228 827 21232
rect 793 21198 827 21228
rect 793 21126 827 21160
rect 793 21058 827 21088
rect 793 21054 827 21058
rect 889 21228 923 21232
rect 889 21198 923 21228
rect 889 21126 923 21160
rect 889 21058 923 21088
rect 889 21054 923 21058
rect 985 21228 1019 21232
rect 985 21198 1019 21228
rect 985 21126 1019 21160
rect 985 21058 1019 21088
rect 985 21054 1019 21058
rect 1081 21228 1115 21232
rect 1081 21198 1115 21228
rect 1081 21126 1115 21160
rect 1081 21058 1115 21088
rect 1081 21054 1115 21058
rect 1177 21228 1211 21232
rect 1177 21198 1211 21228
rect 1177 21126 1211 21160
rect 1177 21058 1211 21088
rect 1177 21054 1211 21058
rect 1273 21228 1307 21232
rect 1273 21198 1307 21228
rect 1273 21126 1307 21160
rect 1273 21058 1307 21088
rect 1273 21054 1307 21058
rect 1387 21259 1421 21263
rect 1387 21229 1421 21259
rect 1387 21157 1421 21191
rect 1387 21089 1421 21119
rect 1387 21085 1421 21089
rect 1387 21021 1421 21047
rect 1387 21013 1421 21021
rect 2466 21331 2500 21365
rect 2658 21331 2692 21365
rect 2850 21331 2884 21365
rect 3042 21331 3076 21365
rect 3234 21331 3268 21365
rect 3426 21331 3460 21365
rect 3540 21331 3574 21339
rect 3540 21305 3574 21331
rect 2466 21232 2500 21236
rect 2466 21202 2500 21232
rect 2466 21130 2500 21164
rect 2466 21062 2500 21092
rect 2466 21058 2500 21062
rect 2562 21232 2596 21236
rect 2562 21202 2596 21232
rect 2562 21130 2596 21164
rect 2562 21062 2596 21092
rect 2562 21058 2596 21062
rect 2658 21232 2692 21236
rect 2658 21202 2692 21232
rect 2658 21130 2692 21164
rect 2658 21062 2692 21092
rect 2658 21058 2692 21062
rect 2754 21232 2788 21236
rect 2754 21202 2788 21232
rect 2754 21130 2788 21164
rect 2754 21062 2788 21092
rect 2754 21058 2788 21062
rect 2850 21232 2884 21236
rect 2850 21202 2884 21232
rect 2850 21130 2884 21164
rect 2850 21062 2884 21092
rect 2850 21058 2884 21062
rect 2946 21232 2980 21236
rect 2946 21202 2980 21232
rect 2946 21130 2980 21164
rect 2946 21062 2980 21092
rect 2946 21058 2980 21062
rect 3042 21232 3076 21236
rect 3042 21202 3076 21232
rect 3042 21130 3076 21164
rect 3042 21062 3076 21092
rect 3042 21058 3076 21062
rect 3138 21232 3172 21236
rect 3138 21202 3172 21232
rect 3138 21130 3172 21164
rect 3138 21062 3172 21092
rect 3138 21058 3172 21062
rect 3234 21232 3268 21236
rect 3234 21202 3268 21232
rect 3234 21130 3268 21164
rect 3234 21062 3268 21092
rect 3234 21058 3268 21062
rect 3330 21232 3364 21236
rect 3330 21202 3364 21232
rect 3330 21130 3364 21164
rect 3330 21062 3364 21092
rect 3330 21058 3364 21062
rect 3426 21232 3460 21236
rect 3426 21202 3460 21232
rect 3426 21130 3460 21164
rect 3426 21062 3460 21092
rect 3426 21058 3460 21062
rect 3540 21263 3574 21267
rect 3540 21233 3574 21263
rect 3540 21161 3574 21195
rect 3540 21093 3574 21123
rect 3540 21089 3574 21093
rect 3540 21025 3574 21051
rect 3540 21017 3574 21025
rect 3987 21331 4021 21365
rect 4179 21331 4213 21365
rect 4371 21331 4405 21365
rect 4563 21331 4597 21365
rect 4755 21331 4789 21365
rect 4947 21331 4981 21365
rect 5061 21331 5095 21339
rect 5061 21305 5095 21331
rect 3987 21232 4021 21236
rect 3987 21202 4021 21232
rect 3987 21130 4021 21164
rect 3987 21062 4021 21092
rect 3987 21058 4021 21062
rect 4083 21232 4117 21236
rect 4083 21202 4117 21232
rect 4083 21130 4117 21164
rect 4083 21062 4117 21092
rect 4083 21058 4117 21062
rect 4179 21232 4213 21236
rect 4179 21202 4213 21232
rect 4179 21130 4213 21164
rect 4179 21062 4213 21092
rect 4179 21058 4213 21062
rect 4275 21232 4309 21236
rect 4275 21202 4309 21232
rect 4275 21130 4309 21164
rect 4275 21062 4309 21092
rect 4275 21058 4309 21062
rect 4371 21232 4405 21236
rect 4371 21202 4405 21232
rect 4371 21130 4405 21164
rect 4371 21062 4405 21092
rect 4371 21058 4405 21062
rect 4467 21232 4501 21236
rect 4467 21202 4501 21232
rect 4467 21130 4501 21164
rect 4467 21062 4501 21092
rect 4467 21058 4501 21062
rect 4563 21232 4597 21236
rect 4563 21202 4597 21232
rect 4563 21130 4597 21164
rect 4563 21062 4597 21092
rect 4563 21058 4597 21062
rect 4659 21232 4693 21236
rect 4659 21202 4693 21232
rect 4659 21130 4693 21164
rect 4659 21062 4693 21092
rect 4659 21058 4693 21062
rect 4755 21232 4789 21236
rect 4755 21202 4789 21232
rect 4755 21130 4789 21164
rect 4755 21062 4789 21092
rect 4755 21058 4789 21062
rect 4851 21232 4885 21236
rect 4851 21202 4885 21232
rect 4851 21130 4885 21164
rect 4851 21062 4885 21092
rect 4851 21058 4885 21062
rect 4947 21232 4981 21236
rect 4947 21202 4981 21232
rect 4947 21130 4981 21164
rect 4947 21062 4981 21092
rect 4947 21058 4981 21062
rect 5061 21263 5095 21267
rect 5061 21233 5095 21263
rect 5061 21161 5095 21195
rect 5061 21093 5095 21123
rect 5303 21100 5337 21134
rect 5395 21100 5429 21134
rect 5487 21100 5521 21134
rect 5061 21089 5095 21093
rect 5061 21025 5095 21051
rect 5061 21017 5095 21025
rect 313 20630 347 20664
rect 409 20630 443 20664
rect 505 20630 539 20664
rect 601 20630 635 20664
rect 697 20630 731 20664
rect 793 20630 827 20664
rect 889 20630 923 20664
rect 985 20630 1019 20664
rect 1081 20630 1115 20664
rect 1177 20630 1211 20664
rect 1273 20630 1307 20664
rect 1387 20701 1421 20706
rect 1387 20672 1421 20701
rect 1387 20633 1421 20634
rect 1387 20600 1421 20633
rect 313 20519 347 20553
rect 505 20519 539 20553
rect 697 20519 731 20553
rect 889 20519 923 20553
rect 1081 20519 1115 20553
rect 1273 20519 1307 20553
rect 1387 20531 1421 20562
rect 1387 20528 1421 20531
rect 3691 20745 3725 20779
rect 2466 20634 2500 20668
rect 2562 20634 2596 20668
rect 2658 20634 2692 20668
rect 2754 20634 2788 20668
rect 2850 20634 2884 20668
rect 2946 20634 2980 20668
rect 3042 20634 3076 20668
rect 3138 20634 3172 20668
rect 3234 20634 3268 20668
rect 3330 20634 3364 20668
rect 3426 20634 3460 20668
rect 3540 20705 3574 20710
rect 3540 20676 3574 20705
rect 3540 20637 3574 20638
rect 3540 20604 3574 20637
rect 3647 20619 3681 20695
rect 3735 20619 3769 20695
rect 2466 20523 2500 20557
rect 2658 20523 2692 20557
rect 2850 20523 2884 20557
rect 3042 20523 3076 20557
rect 3234 20523 3268 20557
rect 3426 20523 3460 20557
rect 3540 20535 3574 20566
rect 3540 20532 3574 20535
rect 3987 20634 4021 20668
rect 4083 20634 4117 20668
rect 4179 20634 4213 20668
rect 4275 20634 4309 20668
rect 4371 20634 4405 20668
rect 4467 20634 4501 20668
rect 4563 20634 4597 20668
rect 4659 20634 4693 20668
rect 4755 20634 4789 20668
rect 4851 20634 4885 20668
rect 4947 20634 4981 20668
rect 5061 20705 5095 20710
rect 5061 20676 5095 20705
rect 5061 20637 5095 20638
rect 5061 20604 5095 20637
rect 5348 20786 5382 20820
rect 5450 20822 5484 20825
rect 5450 20791 5470 20822
rect 5470 20791 5484 20822
rect 3987 20523 4021 20557
rect 4179 20523 4213 20557
rect 4371 20523 4405 20557
rect 4563 20523 4597 20557
rect 4755 20523 4789 20557
rect 4947 20523 4981 20557
rect 5061 20535 5095 20566
rect 5303 20556 5337 20590
rect 5395 20556 5429 20590
rect 5487 20556 5521 20590
rect 5061 20532 5095 20535
rect 313 20040 347 20074
rect 505 20040 539 20074
rect 697 20040 731 20074
rect 889 20040 923 20074
rect 1081 20040 1115 20074
rect 1273 20040 1307 20074
rect 1387 20040 1421 20048
rect 1387 20014 1421 20040
rect 313 19941 347 19945
rect 313 19911 347 19941
rect 313 19839 347 19873
rect 313 19771 347 19801
rect 313 19767 347 19771
rect 409 19941 443 19945
rect 409 19911 443 19941
rect 409 19839 443 19873
rect 409 19771 443 19801
rect 409 19767 443 19771
rect 505 19941 539 19945
rect 505 19911 539 19941
rect 505 19839 539 19873
rect 505 19771 539 19801
rect 505 19767 539 19771
rect 601 19941 635 19945
rect 601 19911 635 19941
rect 601 19839 635 19873
rect 601 19771 635 19801
rect 601 19767 635 19771
rect 697 19941 731 19945
rect 697 19911 731 19941
rect 697 19839 731 19873
rect 697 19771 731 19801
rect 697 19767 731 19771
rect 793 19941 827 19945
rect 793 19911 827 19941
rect 793 19839 827 19873
rect 793 19771 827 19801
rect 793 19767 827 19771
rect 889 19941 923 19945
rect 889 19911 923 19941
rect 889 19839 923 19873
rect 889 19771 923 19801
rect 889 19767 923 19771
rect 985 19941 1019 19945
rect 985 19911 1019 19941
rect 985 19839 1019 19873
rect 985 19771 1019 19801
rect 985 19767 1019 19771
rect 1081 19941 1115 19945
rect 1081 19911 1115 19941
rect 1081 19839 1115 19873
rect 1081 19771 1115 19801
rect 1081 19767 1115 19771
rect 1177 19941 1211 19945
rect 1177 19911 1211 19941
rect 1177 19839 1211 19873
rect 1177 19771 1211 19801
rect 1177 19767 1211 19771
rect 1273 19941 1307 19945
rect 1273 19911 1307 19941
rect 1273 19839 1307 19873
rect 1273 19771 1307 19801
rect 1273 19767 1307 19771
rect 1387 19972 1421 19976
rect 1387 19942 1421 19972
rect 1387 19870 1421 19904
rect 1387 19802 1421 19832
rect 1387 19798 1421 19802
rect 1387 19734 1421 19760
rect 1387 19726 1421 19734
rect 2466 20044 2500 20078
rect 2658 20044 2692 20078
rect 2850 20044 2884 20078
rect 3042 20044 3076 20078
rect 3234 20044 3268 20078
rect 3426 20044 3460 20078
rect 3540 20044 3574 20052
rect 3540 20018 3574 20044
rect 2466 19945 2500 19949
rect 2466 19915 2500 19945
rect 2466 19843 2500 19877
rect 2466 19775 2500 19805
rect 2466 19771 2500 19775
rect 2562 19945 2596 19949
rect 2562 19915 2596 19945
rect 2562 19843 2596 19877
rect 2562 19775 2596 19805
rect 2562 19771 2596 19775
rect 2658 19945 2692 19949
rect 2658 19915 2692 19945
rect 2658 19843 2692 19877
rect 2658 19775 2692 19805
rect 2658 19771 2692 19775
rect 2754 19945 2788 19949
rect 2754 19915 2788 19945
rect 2754 19843 2788 19877
rect 2754 19775 2788 19805
rect 2754 19771 2788 19775
rect 2850 19945 2884 19949
rect 2850 19915 2884 19945
rect 2850 19843 2884 19877
rect 2850 19775 2884 19805
rect 2850 19771 2884 19775
rect 2946 19945 2980 19949
rect 2946 19915 2980 19945
rect 2946 19843 2980 19877
rect 2946 19775 2980 19805
rect 2946 19771 2980 19775
rect 3042 19945 3076 19949
rect 3042 19915 3076 19945
rect 3042 19843 3076 19877
rect 3042 19775 3076 19805
rect 3042 19771 3076 19775
rect 3138 19945 3172 19949
rect 3138 19915 3172 19945
rect 3138 19843 3172 19877
rect 3138 19775 3172 19805
rect 3138 19771 3172 19775
rect 3234 19945 3268 19949
rect 3234 19915 3268 19945
rect 3234 19843 3268 19877
rect 3234 19775 3268 19805
rect 3234 19771 3268 19775
rect 3330 19945 3364 19949
rect 3330 19915 3364 19945
rect 3330 19843 3364 19877
rect 3330 19775 3364 19805
rect 3330 19771 3364 19775
rect 3426 19945 3460 19949
rect 3426 19915 3460 19945
rect 3426 19843 3460 19877
rect 3426 19775 3460 19805
rect 3426 19771 3460 19775
rect 3540 19976 3574 19980
rect 3540 19946 3574 19976
rect 3540 19874 3574 19908
rect 3540 19806 3574 19836
rect 3540 19802 3574 19806
rect 3540 19738 3574 19764
rect 3540 19730 3574 19738
rect 3987 20044 4021 20078
rect 4179 20044 4213 20078
rect 4371 20044 4405 20078
rect 4563 20044 4597 20078
rect 4755 20044 4789 20078
rect 4947 20044 4981 20078
rect 5061 20044 5095 20052
rect 5061 20018 5095 20044
rect 3987 19945 4021 19949
rect 3987 19915 4021 19945
rect 3987 19843 4021 19877
rect 3987 19775 4021 19805
rect 3987 19771 4021 19775
rect 4083 19945 4117 19949
rect 4083 19915 4117 19945
rect 4083 19843 4117 19877
rect 4083 19775 4117 19805
rect 4083 19771 4117 19775
rect 4179 19945 4213 19949
rect 4179 19915 4213 19945
rect 4179 19843 4213 19877
rect 4179 19775 4213 19805
rect 4179 19771 4213 19775
rect 4275 19945 4309 19949
rect 4275 19915 4309 19945
rect 4275 19843 4309 19877
rect 4275 19775 4309 19805
rect 4275 19771 4309 19775
rect 4371 19945 4405 19949
rect 4371 19915 4405 19945
rect 4371 19843 4405 19877
rect 4371 19775 4405 19805
rect 4371 19771 4405 19775
rect 4467 19945 4501 19949
rect 4467 19915 4501 19945
rect 4467 19843 4501 19877
rect 4467 19775 4501 19805
rect 4467 19771 4501 19775
rect 4563 19945 4597 19949
rect 4563 19915 4597 19945
rect 4563 19843 4597 19877
rect 4563 19775 4597 19805
rect 4563 19771 4597 19775
rect 4659 19945 4693 19949
rect 4659 19915 4693 19945
rect 4659 19843 4693 19877
rect 4659 19775 4693 19805
rect 4659 19771 4693 19775
rect 4755 19945 4789 19949
rect 4755 19915 4789 19945
rect 4755 19843 4789 19877
rect 4755 19775 4789 19805
rect 4755 19771 4789 19775
rect 4851 19945 4885 19949
rect 4851 19915 4885 19945
rect 4851 19843 4885 19877
rect 4851 19775 4885 19805
rect 4851 19771 4885 19775
rect 4947 19945 4981 19949
rect 4947 19915 4981 19945
rect 4947 19843 4981 19877
rect 4947 19775 4981 19805
rect 4947 19771 4981 19775
rect 5061 19976 5095 19980
rect 5061 19946 5095 19976
rect 5061 19874 5095 19908
rect 5061 19806 5095 19836
rect 5303 19813 5337 19847
rect 5395 19813 5429 19847
rect 5487 19813 5521 19847
rect 5061 19802 5095 19806
rect 5061 19738 5095 19764
rect 5061 19730 5095 19738
rect 313 19343 347 19377
rect 409 19343 443 19377
rect 505 19343 539 19377
rect 601 19343 635 19377
rect 697 19343 731 19377
rect 793 19343 827 19377
rect 889 19343 923 19377
rect 985 19343 1019 19377
rect 1081 19343 1115 19377
rect 1177 19343 1211 19377
rect 1273 19343 1307 19377
rect 1387 19414 1421 19419
rect 1387 19385 1421 19414
rect 1387 19346 1421 19347
rect 1387 19313 1421 19346
rect 313 19232 347 19266
rect 505 19232 539 19266
rect 697 19232 731 19266
rect 889 19232 923 19266
rect 1081 19232 1115 19266
rect 1273 19232 1307 19266
rect 1387 19244 1421 19275
rect 1387 19241 1421 19244
rect 3691 19458 3725 19492
rect 2466 19347 2500 19381
rect 2562 19347 2596 19381
rect 2658 19347 2692 19381
rect 2754 19347 2788 19381
rect 2850 19347 2884 19381
rect 2946 19347 2980 19381
rect 3042 19347 3076 19381
rect 3138 19347 3172 19381
rect 3234 19347 3268 19381
rect 3330 19347 3364 19381
rect 3426 19347 3460 19381
rect 3540 19418 3574 19423
rect 3540 19389 3574 19418
rect 3540 19350 3574 19351
rect 3540 19317 3574 19350
rect 3647 19332 3681 19408
rect 3735 19332 3769 19408
rect 2466 19236 2500 19270
rect 2658 19236 2692 19270
rect 2850 19236 2884 19270
rect 3042 19236 3076 19270
rect 3234 19236 3268 19270
rect 3426 19236 3460 19270
rect 3540 19248 3574 19279
rect 3540 19245 3574 19248
rect 3987 19347 4021 19381
rect 4083 19347 4117 19381
rect 4179 19347 4213 19381
rect 4275 19347 4309 19381
rect 4371 19347 4405 19381
rect 4467 19347 4501 19381
rect 4563 19347 4597 19381
rect 4659 19347 4693 19381
rect 4755 19347 4789 19381
rect 4851 19347 4885 19381
rect 4947 19347 4981 19381
rect 5061 19418 5095 19423
rect 5061 19389 5095 19418
rect 5061 19350 5095 19351
rect 5061 19317 5095 19350
rect 5348 19499 5382 19533
rect 5450 19535 5484 19538
rect 5450 19504 5470 19535
rect 5470 19504 5484 19535
rect 3987 19236 4021 19270
rect 4179 19236 4213 19270
rect 4371 19236 4405 19270
rect 4563 19236 4597 19270
rect 4755 19236 4789 19270
rect 4947 19236 4981 19270
rect 5061 19248 5095 19279
rect 5303 19269 5337 19303
rect 5395 19269 5429 19303
rect 5487 19269 5521 19303
rect 5061 19245 5095 19248
rect 313 18753 347 18787
rect 505 18753 539 18787
rect 697 18753 731 18787
rect 889 18753 923 18787
rect 1081 18753 1115 18787
rect 1273 18753 1307 18787
rect 1387 18753 1421 18761
rect 1387 18727 1421 18753
rect 313 18654 347 18658
rect 313 18624 347 18654
rect 313 18552 347 18586
rect 313 18484 347 18514
rect 313 18480 347 18484
rect 409 18654 443 18658
rect 409 18624 443 18654
rect 409 18552 443 18586
rect 409 18484 443 18514
rect 409 18480 443 18484
rect 505 18654 539 18658
rect 505 18624 539 18654
rect 505 18552 539 18586
rect 505 18484 539 18514
rect 505 18480 539 18484
rect 601 18654 635 18658
rect 601 18624 635 18654
rect 601 18552 635 18586
rect 601 18484 635 18514
rect 601 18480 635 18484
rect 697 18654 731 18658
rect 697 18624 731 18654
rect 697 18552 731 18586
rect 697 18484 731 18514
rect 697 18480 731 18484
rect 793 18654 827 18658
rect 793 18624 827 18654
rect 793 18552 827 18586
rect 793 18484 827 18514
rect 793 18480 827 18484
rect 889 18654 923 18658
rect 889 18624 923 18654
rect 889 18552 923 18586
rect 889 18484 923 18514
rect 889 18480 923 18484
rect 985 18654 1019 18658
rect 985 18624 1019 18654
rect 985 18552 1019 18586
rect 985 18484 1019 18514
rect 985 18480 1019 18484
rect 1081 18654 1115 18658
rect 1081 18624 1115 18654
rect 1081 18552 1115 18586
rect 1081 18484 1115 18514
rect 1081 18480 1115 18484
rect 1177 18654 1211 18658
rect 1177 18624 1211 18654
rect 1177 18552 1211 18586
rect 1177 18484 1211 18514
rect 1177 18480 1211 18484
rect 1273 18654 1307 18658
rect 1273 18624 1307 18654
rect 1273 18552 1307 18586
rect 1273 18484 1307 18514
rect 1273 18480 1307 18484
rect 1387 18685 1421 18689
rect 1387 18655 1421 18685
rect 1387 18583 1421 18617
rect 1387 18515 1421 18545
rect 1387 18511 1421 18515
rect 1387 18447 1421 18473
rect 1387 18439 1421 18447
rect 2466 18757 2500 18791
rect 2658 18757 2692 18791
rect 2850 18757 2884 18791
rect 3042 18757 3076 18791
rect 3234 18757 3268 18791
rect 3426 18757 3460 18791
rect 3540 18757 3574 18765
rect 3540 18731 3574 18757
rect 2466 18658 2500 18662
rect 2466 18628 2500 18658
rect 2466 18556 2500 18590
rect 2466 18488 2500 18518
rect 2466 18484 2500 18488
rect 2562 18658 2596 18662
rect 2562 18628 2596 18658
rect 2562 18556 2596 18590
rect 2562 18488 2596 18518
rect 2562 18484 2596 18488
rect 2658 18658 2692 18662
rect 2658 18628 2692 18658
rect 2658 18556 2692 18590
rect 2658 18488 2692 18518
rect 2658 18484 2692 18488
rect 2754 18658 2788 18662
rect 2754 18628 2788 18658
rect 2754 18556 2788 18590
rect 2754 18488 2788 18518
rect 2754 18484 2788 18488
rect 2850 18658 2884 18662
rect 2850 18628 2884 18658
rect 2850 18556 2884 18590
rect 2850 18488 2884 18518
rect 2850 18484 2884 18488
rect 2946 18658 2980 18662
rect 2946 18628 2980 18658
rect 2946 18556 2980 18590
rect 2946 18488 2980 18518
rect 2946 18484 2980 18488
rect 3042 18658 3076 18662
rect 3042 18628 3076 18658
rect 3042 18556 3076 18590
rect 3042 18488 3076 18518
rect 3042 18484 3076 18488
rect 3138 18658 3172 18662
rect 3138 18628 3172 18658
rect 3138 18556 3172 18590
rect 3138 18488 3172 18518
rect 3138 18484 3172 18488
rect 3234 18658 3268 18662
rect 3234 18628 3268 18658
rect 3234 18556 3268 18590
rect 3234 18488 3268 18518
rect 3234 18484 3268 18488
rect 3330 18658 3364 18662
rect 3330 18628 3364 18658
rect 3330 18556 3364 18590
rect 3330 18488 3364 18518
rect 3330 18484 3364 18488
rect 3426 18658 3460 18662
rect 3426 18628 3460 18658
rect 3426 18556 3460 18590
rect 3426 18488 3460 18518
rect 3426 18484 3460 18488
rect 3540 18689 3574 18693
rect 3540 18659 3574 18689
rect 3540 18587 3574 18621
rect 3540 18519 3574 18549
rect 3540 18515 3574 18519
rect 3540 18451 3574 18477
rect 3540 18443 3574 18451
rect 3987 18757 4021 18791
rect 4179 18757 4213 18791
rect 4371 18757 4405 18791
rect 4563 18757 4597 18791
rect 4755 18757 4789 18791
rect 4947 18757 4981 18791
rect 5061 18757 5095 18765
rect 5061 18731 5095 18757
rect 3987 18658 4021 18662
rect 3987 18628 4021 18658
rect 3987 18556 4021 18590
rect 3987 18488 4021 18518
rect 3987 18484 4021 18488
rect 4083 18658 4117 18662
rect 4083 18628 4117 18658
rect 4083 18556 4117 18590
rect 4083 18488 4117 18518
rect 4083 18484 4117 18488
rect 4179 18658 4213 18662
rect 4179 18628 4213 18658
rect 4179 18556 4213 18590
rect 4179 18488 4213 18518
rect 4179 18484 4213 18488
rect 4275 18658 4309 18662
rect 4275 18628 4309 18658
rect 4275 18556 4309 18590
rect 4275 18488 4309 18518
rect 4275 18484 4309 18488
rect 4371 18658 4405 18662
rect 4371 18628 4405 18658
rect 4371 18556 4405 18590
rect 4371 18488 4405 18518
rect 4371 18484 4405 18488
rect 4467 18658 4501 18662
rect 4467 18628 4501 18658
rect 4467 18556 4501 18590
rect 4467 18488 4501 18518
rect 4467 18484 4501 18488
rect 4563 18658 4597 18662
rect 4563 18628 4597 18658
rect 4563 18556 4597 18590
rect 4563 18488 4597 18518
rect 4563 18484 4597 18488
rect 4659 18658 4693 18662
rect 4659 18628 4693 18658
rect 4659 18556 4693 18590
rect 4659 18488 4693 18518
rect 4659 18484 4693 18488
rect 4755 18658 4789 18662
rect 4755 18628 4789 18658
rect 4755 18556 4789 18590
rect 4755 18488 4789 18518
rect 4755 18484 4789 18488
rect 4851 18658 4885 18662
rect 4851 18628 4885 18658
rect 4851 18556 4885 18590
rect 4851 18488 4885 18518
rect 4851 18484 4885 18488
rect 4947 18658 4981 18662
rect 4947 18628 4981 18658
rect 4947 18556 4981 18590
rect 4947 18488 4981 18518
rect 4947 18484 4981 18488
rect 5061 18689 5095 18693
rect 5061 18659 5095 18689
rect 5061 18587 5095 18621
rect 5061 18519 5095 18549
rect 5303 18526 5337 18560
rect 5395 18526 5429 18560
rect 5487 18526 5521 18560
rect 5061 18515 5095 18519
rect 5061 18451 5095 18477
rect 5061 18443 5095 18451
rect 313 18056 347 18090
rect 409 18056 443 18090
rect 505 18056 539 18090
rect 601 18056 635 18090
rect 697 18056 731 18090
rect 793 18056 827 18090
rect 889 18056 923 18090
rect 985 18056 1019 18090
rect 1081 18056 1115 18090
rect 1177 18056 1211 18090
rect 1273 18056 1307 18090
rect 1387 18127 1421 18132
rect 1387 18098 1421 18127
rect 1387 18059 1421 18060
rect 1387 18026 1421 18059
rect 313 17945 347 17979
rect 505 17945 539 17979
rect 697 17945 731 17979
rect 889 17945 923 17979
rect 1081 17945 1115 17979
rect 1273 17945 1307 17979
rect 1387 17957 1421 17988
rect 1387 17954 1421 17957
rect 3691 18171 3725 18205
rect 2466 18060 2500 18094
rect 2562 18060 2596 18094
rect 2658 18060 2692 18094
rect 2754 18060 2788 18094
rect 2850 18060 2884 18094
rect 2946 18060 2980 18094
rect 3042 18060 3076 18094
rect 3138 18060 3172 18094
rect 3234 18060 3268 18094
rect 3330 18060 3364 18094
rect 3426 18060 3460 18094
rect 3540 18131 3574 18136
rect 3540 18102 3574 18131
rect 3540 18063 3574 18064
rect 3540 18030 3574 18063
rect 3647 18045 3681 18121
rect 3735 18045 3769 18121
rect 2466 17949 2500 17983
rect 2658 17949 2692 17983
rect 2850 17949 2884 17983
rect 3042 17949 3076 17983
rect 3234 17949 3268 17983
rect 3426 17949 3460 17983
rect 3540 17961 3574 17992
rect 3540 17958 3574 17961
rect 3987 18060 4021 18094
rect 4083 18060 4117 18094
rect 4179 18060 4213 18094
rect 4275 18060 4309 18094
rect 4371 18060 4405 18094
rect 4467 18060 4501 18094
rect 4563 18060 4597 18094
rect 4659 18060 4693 18094
rect 4755 18060 4789 18094
rect 4851 18060 4885 18094
rect 4947 18060 4981 18094
rect 5061 18131 5095 18136
rect 5061 18102 5095 18131
rect 5061 18063 5095 18064
rect 5061 18030 5095 18063
rect 5348 18212 5382 18246
rect 5450 18248 5484 18251
rect 5450 18217 5470 18248
rect 5470 18217 5484 18248
rect 3987 17949 4021 17983
rect 4179 17949 4213 17983
rect 4371 17949 4405 17983
rect 4563 17949 4597 17983
rect 4755 17949 4789 17983
rect 4947 17949 4981 17983
rect 5061 17961 5095 17992
rect 5303 17982 5337 18016
rect 5395 17982 5429 18016
rect 5487 17982 5521 18016
rect 5061 17958 5095 17961
rect 313 17466 347 17500
rect 505 17466 539 17500
rect 697 17466 731 17500
rect 889 17466 923 17500
rect 1081 17466 1115 17500
rect 1273 17466 1307 17500
rect 1387 17466 1421 17474
rect 1387 17440 1421 17466
rect 313 17367 347 17371
rect 313 17337 347 17367
rect 313 17265 347 17299
rect 313 17197 347 17227
rect 313 17193 347 17197
rect 409 17367 443 17371
rect 409 17337 443 17367
rect 409 17265 443 17299
rect 409 17197 443 17227
rect 409 17193 443 17197
rect 505 17367 539 17371
rect 505 17337 539 17367
rect 505 17265 539 17299
rect 505 17197 539 17227
rect 505 17193 539 17197
rect 601 17367 635 17371
rect 601 17337 635 17367
rect 601 17265 635 17299
rect 601 17197 635 17227
rect 601 17193 635 17197
rect 697 17367 731 17371
rect 697 17337 731 17367
rect 697 17265 731 17299
rect 697 17197 731 17227
rect 697 17193 731 17197
rect 793 17367 827 17371
rect 793 17337 827 17367
rect 793 17265 827 17299
rect 793 17197 827 17227
rect 793 17193 827 17197
rect 889 17367 923 17371
rect 889 17337 923 17367
rect 889 17265 923 17299
rect 889 17197 923 17227
rect 889 17193 923 17197
rect 985 17367 1019 17371
rect 985 17337 1019 17367
rect 985 17265 1019 17299
rect 985 17197 1019 17227
rect 985 17193 1019 17197
rect 1081 17367 1115 17371
rect 1081 17337 1115 17367
rect 1081 17265 1115 17299
rect 1081 17197 1115 17227
rect 1081 17193 1115 17197
rect 1177 17367 1211 17371
rect 1177 17337 1211 17367
rect 1177 17265 1211 17299
rect 1177 17197 1211 17227
rect 1177 17193 1211 17197
rect 1273 17367 1307 17371
rect 1273 17337 1307 17367
rect 1273 17265 1307 17299
rect 1273 17197 1307 17227
rect 1273 17193 1307 17197
rect 1387 17398 1421 17402
rect 1387 17368 1421 17398
rect 1387 17296 1421 17330
rect 1387 17228 1421 17258
rect 1387 17224 1421 17228
rect 1387 17160 1421 17186
rect 1387 17152 1421 17160
rect 2466 17470 2500 17504
rect 2658 17470 2692 17504
rect 2850 17470 2884 17504
rect 3042 17470 3076 17504
rect 3234 17470 3268 17504
rect 3426 17470 3460 17504
rect 3540 17470 3574 17478
rect 3540 17444 3574 17470
rect 2466 17371 2500 17375
rect 2466 17341 2500 17371
rect 2466 17269 2500 17303
rect 2466 17201 2500 17231
rect 2466 17197 2500 17201
rect 2562 17371 2596 17375
rect 2562 17341 2596 17371
rect 2562 17269 2596 17303
rect 2562 17201 2596 17231
rect 2562 17197 2596 17201
rect 2658 17371 2692 17375
rect 2658 17341 2692 17371
rect 2658 17269 2692 17303
rect 2658 17201 2692 17231
rect 2658 17197 2692 17201
rect 2754 17371 2788 17375
rect 2754 17341 2788 17371
rect 2754 17269 2788 17303
rect 2754 17201 2788 17231
rect 2754 17197 2788 17201
rect 2850 17371 2884 17375
rect 2850 17341 2884 17371
rect 2850 17269 2884 17303
rect 2850 17201 2884 17231
rect 2850 17197 2884 17201
rect 2946 17371 2980 17375
rect 2946 17341 2980 17371
rect 2946 17269 2980 17303
rect 2946 17201 2980 17231
rect 2946 17197 2980 17201
rect 3042 17371 3076 17375
rect 3042 17341 3076 17371
rect 3042 17269 3076 17303
rect 3042 17201 3076 17231
rect 3042 17197 3076 17201
rect 3138 17371 3172 17375
rect 3138 17341 3172 17371
rect 3138 17269 3172 17303
rect 3138 17201 3172 17231
rect 3138 17197 3172 17201
rect 3234 17371 3268 17375
rect 3234 17341 3268 17371
rect 3234 17269 3268 17303
rect 3234 17201 3268 17231
rect 3234 17197 3268 17201
rect 3330 17371 3364 17375
rect 3330 17341 3364 17371
rect 3330 17269 3364 17303
rect 3330 17201 3364 17231
rect 3330 17197 3364 17201
rect 3426 17371 3460 17375
rect 3426 17341 3460 17371
rect 3426 17269 3460 17303
rect 3426 17201 3460 17231
rect 3426 17197 3460 17201
rect 3540 17402 3574 17406
rect 3540 17372 3574 17402
rect 3540 17300 3574 17334
rect 3540 17232 3574 17262
rect 3540 17228 3574 17232
rect 3540 17164 3574 17190
rect 3540 17156 3574 17164
rect 3987 17470 4021 17504
rect 4179 17470 4213 17504
rect 4371 17470 4405 17504
rect 4563 17470 4597 17504
rect 4755 17470 4789 17504
rect 4947 17470 4981 17504
rect 5061 17470 5095 17478
rect 5061 17444 5095 17470
rect 3987 17371 4021 17375
rect 3987 17341 4021 17371
rect 3987 17269 4021 17303
rect 3987 17201 4021 17231
rect 3987 17197 4021 17201
rect 4083 17371 4117 17375
rect 4083 17341 4117 17371
rect 4083 17269 4117 17303
rect 4083 17201 4117 17231
rect 4083 17197 4117 17201
rect 4179 17371 4213 17375
rect 4179 17341 4213 17371
rect 4179 17269 4213 17303
rect 4179 17201 4213 17231
rect 4179 17197 4213 17201
rect 4275 17371 4309 17375
rect 4275 17341 4309 17371
rect 4275 17269 4309 17303
rect 4275 17201 4309 17231
rect 4275 17197 4309 17201
rect 4371 17371 4405 17375
rect 4371 17341 4405 17371
rect 4371 17269 4405 17303
rect 4371 17201 4405 17231
rect 4371 17197 4405 17201
rect 4467 17371 4501 17375
rect 4467 17341 4501 17371
rect 4467 17269 4501 17303
rect 4467 17201 4501 17231
rect 4467 17197 4501 17201
rect 4563 17371 4597 17375
rect 4563 17341 4597 17371
rect 4563 17269 4597 17303
rect 4563 17201 4597 17231
rect 4563 17197 4597 17201
rect 4659 17371 4693 17375
rect 4659 17341 4693 17371
rect 4659 17269 4693 17303
rect 4659 17201 4693 17231
rect 4659 17197 4693 17201
rect 4755 17371 4789 17375
rect 4755 17341 4789 17371
rect 4755 17269 4789 17303
rect 4755 17201 4789 17231
rect 4755 17197 4789 17201
rect 4851 17371 4885 17375
rect 4851 17341 4885 17371
rect 4851 17269 4885 17303
rect 4851 17201 4885 17231
rect 4851 17197 4885 17201
rect 4947 17371 4981 17375
rect 4947 17341 4981 17371
rect 4947 17269 4981 17303
rect 4947 17201 4981 17231
rect 4947 17197 4981 17201
rect 5061 17402 5095 17406
rect 5061 17372 5095 17402
rect 5061 17300 5095 17334
rect 5061 17232 5095 17262
rect 5303 17239 5337 17273
rect 5395 17239 5429 17273
rect 5487 17239 5521 17273
rect 5061 17228 5095 17232
rect 5061 17164 5095 17190
rect 5061 17156 5095 17164
rect 313 16769 347 16803
rect 409 16769 443 16803
rect 505 16769 539 16803
rect 601 16769 635 16803
rect 697 16769 731 16803
rect 793 16769 827 16803
rect 889 16769 923 16803
rect 985 16769 1019 16803
rect 1081 16769 1115 16803
rect 1177 16769 1211 16803
rect 1273 16769 1307 16803
rect 1387 16840 1421 16845
rect 1387 16811 1421 16840
rect 1387 16772 1421 16773
rect 1387 16739 1421 16772
rect 313 16658 347 16692
rect 505 16658 539 16692
rect 697 16658 731 16692
rect 889 16658 923 16692
rect 1081 16658 1115 16692
rect 1273 16658 1307 16692
rect 1387 16670 1421 16701
rect 1387 16667 1421 16670
rect 3691 16884 3725 16918
rect 2466 16773 2500 16807
rect 2562 16773 2596 16807
rect 2658 16773 2692 16807
rect 2754 16773 2788 16807
rect 2850 16773 2884 16807
rect 2946 16773 2980 16807
rect 3042 16773 3076 16807
rect 3138 16773 3172 16807
rect 3234 16773 3268 16807
rect 3330 16773 3364 16807
rect 3426 16773 3460 16807
rect 3540 16844 3574 16849
rect 3540 16815 3574 16844
rect 3540 16776 3574 16777
rect 3540 16743 3574 16776
rect 3647 16758 3681 16834
rect 3735 16758 3769 16834
rect 2466 16662 2500 16696
rect 2658 16662 2692 16696
rect 2850 16662 2884 16696
rect 3042 16662 3076 16696
rect 3234 16662 3268 16696
rect 3426 16662 3460 16696
rect 3540 16674 3574 16705
rect 3540 16671 3574 16674
rect 3987 16773 4021 16807
rect 4083 16773 4117 16807
rect 4179 16773 4213 16807
rect 4275 16773 4309 16807
rect 4371 16773 4405 16807
rect 4467 16773 4501 16807
rect 4563 16773 4597 16807
rect 4659 16773 4693 16807
rect 4755 16773 4789 16807
rect 4851 16773 4885 16807
rect 4947 16773 4981 16807
rect 5061 16844 5095 16849
rect 5061 16815 5095 16844
rect 5061 16776 5095 16777
rect 5061 16743 5095 16776
rect 5348 16925 5382 16959
rect 5450 16961 5484 16964
rect 5450 16930 5470 16961
rect 5470 16930 5484 16961
rect 3987 16662 4021 16696
rect 4179 16662 4213 16696
rect 4371 16662 4405 16696
rect 4563 16662 4597 16696
rect 4755 16662 4789 16696
rect 4947 16662 4981 16696
rect 5061 16674 5095 16705
rect 5303 16695 5337 16729
rect 5395 16695 5429 16729
rect 5487 16695 5521 16729
rect 5061 16671 5095 16674
rect 313 16179 347 16213
rect 505 16179 539 16213
rect 697 16179 731 16213
rect 889 16179 923 16213
rect 1081 16179 1115 16213
rect 1273 16179 1307 16213
rect 1387 16179 1421 16187
rect 1387 16153 1421 16179
rect 313 16080 347 16084
rect 313 16050 347 16080
rect 313 15978 347 16012
rect 313 15910 347 15940
rect 313 15906 347 15910
rect 409 16080 443 16084
rect 409 16050 443 16080
rect 409 15978 443 16012
rect 409 15910 443 15940
rect 409 15906 443 15910
rect 505 16080 539 16084
rect 505 16050 539 16080
rect 505 15978 539 16012
rect 505 15910 539 15940
rect 505 15906 539 15910
rect 601 16080 635 16084
rect 601 16050 635 16080
rect 601 15978 635 16012
rect 601 15910 635 15940
rect 601 15906 635 15910
rect 697 16080 731 16084
rect 697 16050 731 16080
rect 697 15978 731 16012
rect 697 15910 731 15940
rect 697 15906 731 15910
rect 793 16080 827 16084
rect 793 16050 827 16080
rect 793 15978 827 16012
rect 793 15910 827 15940
rect 793 15906 827 15910
rect 889 16080 923 16084
rect 889 16050 923 16080
rect 889 15978 923 16012
rect 889 15910 923 15940
rect 889 15906 923 15910
rect 985 16080 1019 16084
rect 985 16050 1019 16080
rect 985 15978 1019 16012
rect 985 15910 1019 15940
rect 985 15906 1019 15910
rect 1081 16080 1115 16084
rect 1081 16050 1115 16080
rect 1081 15978 1115 16012
rect 1081 15910 1115 15940
rect 1081 15906 1115 15910
rect 1177 16080 1211 16084
rect 1177 16050 1211 16080
rect 1177 15978 1211 16012
rect 1177 15910 1211 15940
rect 1177 15906 1211 15910
rect 1273 16080 1307 16084
rect 1273 16050 1307 16080
rect 1273 15978 1307 16012
rect 1273 15910 1307 15940
rect 1273 15906 1307 15910
rect 1387 16111 1421 16115
rect 1387 16081 1421 16111
rect 1387 16009 1421 16043
rect 1387 15941 1421 15971
rect 1387 15937 1421 15941
rect 1387 15873 1421 15899
rect 1387 15865 1421 15873
rect 2466 16183 2500 16217
rect 2658 16183 2692 16217
rect 2850 16183 2884 16217
rect 3042 16183 3076 16217
rect 3234 16183 3268 16217
rect 3426 16183 3460 16217
rect 3540 16183 3574 16191
rect 3540 16157 3574 16183
rect 2466 16084 2500 16088
rect 2466 16054 2500 16084
rect 2466 15982 2500 16016
rect 2466 15914 2500 15944
rect 2466 15910 2500 15914
rect 2562 16084 2596 16088
rect 2562 16054 2596 16084
rect 2562 15982 2596 16016
rect 2562 15914 2596 15944
rect 2562 15910 2596 15914
rect 2658 16084 2692 16088
rect 2658 16054 2692 16084
rect 2658 15982 2692 16016
rect 2658 15914 2692 15944
rect 2658 15910 2692 15914
rect 2754 16084 2788 16088
rect 2754 16054 2788 16084
rect 2754 15982 2788 16016
rect 2754 15914 2788 15944
rect 2754 15910 2788 15914
rect 2850 16084 2884 16088
rect 2850 16054 2884 16084
rect 2850 15982 2884 16016
rect 2850 15914 2884 15944
rect 2850 15910 2884 15914
rect 2946 16084 2980 16088
rect 2946 16054 2980 16084
rect 2946 15982 2980 16016
rect 2946 15914 2980 15944
rect 2946 15910 2980 15914
rect 3042 16084 3076 16088
rect 3042 16054 3076 16084
rect 3042 15982 3076 16016
rect 3042 15914 3076 15944
rect 3042 15910 3076 15914
rect 3138 16084 3172 16088
rect 3138 16054 3172 16084
rect 3138 15982 3172 16016
rect 3138 15914 3172 15944
rect 3138 15910 3172 15914
rect 3234 16084 3268 16088
rect 3234 16054 3268 16084
rect 3234 15982 3268 16016
rect 3234 15914 3268 15944
rect 3234 15910 3268 15914
rect 3330 16084 3364 16088
rect 3330 16054 3364 16084
rect 3330 15982 3364 16016
rect 3330 15914 3364 15944
rect 3330 15910 3364 15914
rect 3426 16084 3460 16088
rect 3426 16054 3460 16084
rect 3426 15982 3460 16016
rect 3426 15914 3460 15944
rect 3426 15910 3460 15914
rect 3540 16115 3574 16119
rect 3540 16085 3574 16115
rect 3540 16013 3574 16047
rect 3540 15945 3574 15975
rect 3540 15941 3574 15945
rect 3540 15877 3574 15903
rect 3540 15869 3574 15877
rect 3987 16183 4021 16217
rect 4179 16183 4213 16217
rect 4371 16183 4405 16217
rect 4563 16183 4597 16217
rect 4755 16183 4789 16217
rect 4947 16183 4981 16217
rect 5061 16183 5095 16191
rect 5061 16157 5095 16183
rect 3987 16084 4021 16088
rect 3987 16054 4021 16084
rect 3987 15982 4021 16016
rect 3987 15914 4021 15944
rect 3987 15910 4021 15914
rect 4083 16084 4117 16088
rect 4083 16054 4117 16084
rect 4083 15982 4117 16016
rect 4083 15914 4117 15944
rect 4083 15910 4117 15914
rect 4179 16084 4213 16088
rect 4179 16054 4213 16084
rect 4179 15982 4213 16016
rect 4179 15914 4213 15944
rect 4179 15910 4213 15914
rect 4275 16084 4309 16088
rect 4275 16054 4309 16084
rect 4275 15982 4309 16016
rect 4275 15914 4309 15944
rect 4275 15910 4309 15914
rect 4371 16084 4405 16088
rect 4371 16054 4405 16084
rect 4371 15982 4405 16016
rect 4371 15914 4405 15944
rect 4371 15910 4405 15914
rect 4467 16084 4501 16088
rect 4467 16054 4501 16084
rect 4467 15982 4501 16016
rect 4467 15914 4501 15944
rect 4467 15910 4501 15914
rect 4563 16084 4597 16088
rect 4563 16054 4597 16084
rect 4563 15982 4597 16016
rect 4563 15914 4597 15944
rect 4563 15910 4597 15914
rect 4659 16084 4693 16088
rect 4659 16054 4693 16084
rect 4659 15982 4693 16016
rect 4659 15914 4693 15944
rect 4659 15910 4693 15914
rect 4755 16084 4789 16088
rect 4755 16054 4789 16084
rect 4755 15982 4789 16016
rect 4755 15914 4789 15944
rect 4755 15910 4789 15914
rect 4851 16084 4885 16088
rect 4851 16054 4885 16084
rect 4851 15982 4885 16016
rect 4851 15914 4885 15944
rect 4851 15910 4885 15914
rect 4947 16084 4981 16088
rect 4947 16054 4981 16084
rect 4947 15982 4981 16016
rect 4947 15914 4981 15944
rect 4947 15910 4981 15914
rect 5061 16115 5095 16119
rect 5061 16085 5095 16115
rect 5061 16013 5095 16047
rect 5061 15945 5095 15975
rect 5303 15952 5337 15986
rect 5395 15952 5429 15986
rect 5487 15952 5521 15986
rect 5061 15941 5095 15945
rect 5061 15877 5095 15903
rect 5061 15869 5095 15877
rect 313 15482 347 15516
rect 409 15482 443 15516
rect 505 15482 539 15516
rect 601 15482 635 15516
rect 697 15482 731 15516
rect 793 15482 827 15516
rect 889 15482 923 15516
rect 985 15482 1019 15516
rect 1081 15482 1115 15516
rect 1177 15482 1211 15516
rect 1273 15482 1307 15516
rect 1387 15553 1421 15558
rect 1387 15524 1421 15553
rect 1387 15485 1421 15486
rect 1387 15452 1421 15485
rect 313 15371 347 15405
rect 505 15371 539 15405
rect 697 15371 731 15405
rect 889 15371 923 15405
rect 1081 15371 1115 15405
rect 1273 15371 1307 15405
rect 1387 15383 1421 15414
rect 1387 15380 1421 15383
rect 3691 15597 3725 15631
rect 2466 15486 2500 15520
rect 2562 15486 2596 15520
rect 2658 15486 2692 15520
rect 2754 15486 2788 15520
rect 2850 15486 2884 15520
rect 2946 15486 2980 15520
rect 3042 15486 3076 15520
rect 3138 15486 3172 15520
rect 3234 15486 3268 15520
rect 3330 15486 3364 15520
rect 3426 15486 3460 15520
rect 3540 15557 3574 15562
rect 3540 15528 3574 15557
rect 3540 15489 3574 15490
rect 3540 15456 3574 15489
rect 3647 15471 3681 15547
rect 3735 15471 3769 15547
rect 2466 15375 2500 15409
rect 2658 15375 2692 15409
rect 2850 15375 2884 15409
rect 3042 15375 3076 15409
rect 3234 15375 3268 15409
rect 3426 15375 3460 15409
rect 3540 15387 3574 15418
rect 3540 15384 3574 15387
rect 3987 15486 4021 15520
rect 4083 15486 4117 15520
rect 4179 15486 4213 15520
rect 4275 15486 4309 15520
rect 4371 15486 4405 15520
rect 4467 15486 4501 15520
rect 4563 15486 4597 15520
rect 4659 15486 4693 15520
rect 4755 15486 4789 15520
rect 4851 15486 4885 15520
rect 4947 15486 4981 15520
rect 5061 15557 5095 15562
rect 5061 15528 5095 15557
rect 5061 15489 5095 15490
rect 5061 15456 5095 15489
rect 5348 15638 5382 15672
rect 5450 15674 5484 15677
rect 5450 15643 5470 15674
rect 5470 15643 5484 15674
rect 3987 15375 4021 15409
rect 4179 15375 4213 15409
rect 4371 15375 4405 15409
rect 4563 15375 4597 15409
rect 4755 15375 4789 15409
rect 4947 15375 4981 15409
rect 5061 15387 5095 15418
rect 5303 15408 5337 15442
rect 5395 15408 5429 15442
rect 5487 15408 5521 15442
rect 5061 15384 5095 15387
rect 313 14892 347 14926
rect 505 14892 539 14926
rect 697 14892 731 14926
rect 889 14892 923 14926
rect 1081 14892 1115 14926
rect 1273 14892 1307 14926
rect 1387 14892 1421 14900
rect 1387 14866 1421 14892
rect 313 14793 347 14797
rect 313 14763 347 14793
rect 313 14691 347 14725
rect 313 14623 347 14653
rect 313 14619 347 14623
rect 409 14793 443 14797
rect 409 14763 443 14793
rect 409 14691 443 14725
rect 409 14623 443 14653
rect 409 14619 443 14623
rect 505 14793 539 14797
rect 505 14763 539 14793
rect 505 14691 539 14725
rect 505 14623 539 14653
rect 505 14619 539 14623
rect 601 14793 635 14797
rect 601 14763 635 14793
rect 601 14691 635 14725
rect 601 14623 635 14653
rect 601 14619 635 14623
rect 697 14793 731 14797
rect 697 14763 731 14793
rect 697 14691 731 14725
rect 697 14623 731 14653
rect 697 14619 731 14623
rect 793 14793 827 14797
rect 793 14763 827 14793
rect 793 14691 827 14725
rect 793 14623 827 14653
rect 793 14619 827 14623
rect 889 14793 923 14797
rect 889 14763 923 14793
rect 889 14691 923 14725
rect 889 14623 923 14653
rect 889 14619 923 14623
rect 985 14793 1019 14797
rect 985 14763 1019 14793
rect 985 14691 1019 14725
rect 985 14623 1019 14653
rect 985 14619 1019 14623
rect 1081 14793 1115 14797
rect 1081 14763 1115 14793
rect 1081 14691 1115 14725
rect 1081 14623 1115 14653
rect 1081 14619 1115 14623
rect 1177 14793 1211 14797
rect 1177 14763 1211 14793
rect 1177 14691 1211 14725
rect 1177 14623 1211 14653
rect 1177 14619 1211 14623
rect 1273 14793 1307 14797
rect 1273 14763 1307 14793
rect 1273 14691 1307 14725
rect 1273 14623 1307 14653
rect 1273 14619 1307 14623
rect 1387 14824 1421 14828
rect 1387 14794 1421 14824
rect 1387 14722 1421 14756
rect 1387 14654 1421 14684
rect 1387 14650 1421 14654
rect 1387 14586 1421 14612
rect 1387 14578 1421 14586
rect 2466 14896 2500 14930
rect 2658 14896 2692 14930
rect 2850 14896 2884 14930
rect 3042 14896 3076 14930
rect 3234 14896 3268 14930
rect 3426 14896 3460 14930
rect 3540 14896 3574 14904
rect 3540 14870 3574 14896
rect 2466 14797 2500 14801
rect 2466 14767 2500 14797
rect 2466 14695 2500 14729
rect 2466 14627 2500 14657
rect 2466 14623 2500 14627
rect 2562 14797 2596 14801
rect 2562 14767 2596 14797
rect 2562 14695 2596 14729
rect 2562 14627 2596 14657
rect 2562 14623 2596 14627
rect 2658 14797 2692 14801
rect 2658 14767 2692 14797
rect 2658 14695 2692 14729
rect 2658 14627 2692 14657
rect 2658 14623 2692 14627
rect 2754 14797 2788 14801
rect 2754 14767 2788 14797
rect 2754 14695 2788 14729
rect 2754 14627 2788 14657
rect 2754 14623 2788 14627
rect 2850 14797 2884 14801
rect 2850 14767 2884 14797
rect 2850 14695 2884 14729
rect 2850 14627 2884 14657
rect 2850 14623 2884 14627
rect 2946 14797 2980 14801
rect 2946 14767 2980 14797
rect 2946 14695 2980 14729
rect 2946 14627 2980 14657
rect 2946 14623 2980 14627
rect 3042 14797 3076 14801
rect 3042 14767 3076 14797
rect 3042 14695 3076 14729
rect 3042 14627 3076 14657
rect 3042 14623 3076 14627
rect 3138 14797 3172 14801
rect 3138 14767 3172 14797
rect 3138 14695 3172 14729
rect 3138 14627 3172 14657
rect 3138 14623 3172 14627
rect 3234 14797 3268 14801
rect 3234 14767 3268 14797
rect 3234 14695 3268 14729
rect 3234 14627 3268 14657
rect 3234 14623 3268 14627
rect 3330 14797 3364 14801
rect 3330 14767 3364 14797
rect 3330 14695 3364 14729
rect 3330 14627 3364 14657
rect 3330 14623 3364 14627
rect 3426 14797 3460 14801
rect 3426 14767 3460 14797
rect 3426 14695 3460 14729
rect 3426 14627 3460 14657
rect 3426 14623 3460 14627
rect 3540 14828 3574 14832
rect 3540 14798 3574 14828
rect 3540 14726 3574 14760
rect 3540 14658 3574 14688
rect 3540 14654 3574 14658
rect 3540 14590 3574 14616
rect 3540 14582 3574 14590
rect 3987 14896 4021 14930
rect 4179 14896 4213 14930
rect 4371 14896 4405 14930
rect 4563 14896 4597 14930
rect 4755 14896 4789 14930
rect 4947 14896 4981 14930
rect 5061 14896 5095 14904
rect 5061 14870 5095 14896
rect 3987 14797 4021 14801
rect 3987 14767 4021 14797
rect 3987 14695 4021 14729
rect 3987 14627 4021 14657
rect 3987 14623 4021 14627
rect 4083 14797 4117 14801
rect 4083 14767 4117 14797
rect 4083 14695 4117 14729
rect 4083 14627 4117 14657
rect 4083 14623 4117 14627
rect 4179 14797 4213 14801
rect 4179 14767 4213 14797
rect 4179 14695 4213 14729
rect 4179 14627 4213 14657
rect 4179 14623 4213 14627
rect 4275 14797 4309 14801
rect 4275 14767 4309 14797
rect 4275 14695 4309 14729
rect 4275 14627 4309 14657
rect 4275 14623 4309 14627
rect 4371 14797 4405 14801
rect 4371 14767 4405 14797
rect 4371 14695 4405 14729
rect 4371 14627 4405 14657
rect 4371 14623 4405 14627
rect 4467 14797 4501 14801
rect 4467 14767 4501 14797
rect 4467 14695 4501 14729
rect 4467 14627 4501 14657
rect 4467 14623 4501 14627
rect 4563 14797 4597 14801
rect 4563 14767 4597 14797
rect 4563 14695 4597 14729
rect 4563 14627 4597 14657
rect 4563 14623 4597 14627
rect 4659 14797 4693 14801
rect 4659 14767 4693 14797
rect 4659 14695 4693 14729
rect 4659 14627 4693 14657
rect 4659 14623 4693 14627
rect 4755 14797 4789 14801
rect 4755 14767 4789 14797
rect 4755 14695 4789 14729
rect 4755 14627 4789 14657
rect 4755 14623 4789 14627
rect 4851 14797 4885 14801
rect 4851 14767 4885 14797
rect 4851 14695 4885 14729
rect 4851 14627 4885 14657
rect 4851 14623 4885 14627
rect 4947 14797 4981 14801
rect 4947 14767 4981 14797
rect 4947 14695 4981 14729
rect 4947 14627 4981 14657
rect 4947 14623 4981 14627
rect 5061 14828 5095 14832
rect 5061 14798 5095 14828
rect 5061 14726 5095 14760
rect 5061 14658 5095 14688
rect 5303 14665 5337 14699
rect 5395 14665 5429 14699
rect 5487 14665 5521 14699
rect 5061 14654 5095 14658
rect 5061 14590 5095 14616
rect 5061 14582 5095 14590
rect 313 14195 347 14229
rect 409 14195 443 14229
rect 505 14195 539 14229
rect 601 14195 635 14229
rect 697 14195 731 14229
rect 793 14195 827 14229
rect 889 14195 923 14229
rect 985 14195 1019 14229
rect 1081 14195 1115 14229
rect 1177 14195 1211 14229
rect 1273 14195 1307 14229
rect 1387 14266 1421 14271
rect 1387 14237 1421 14266
rect 1387 14198 1421 14199
rect 1387 14165 1421 14198
rect 313 14084 347 14118
rect 505 14084 539 14118
rect 697 14084 731 14118
rect 889 14084 923 14118
rect 1081 14084 1115 14118
rect 1273 14084 1307 14118
rect 1387 14096 1421 14127
rect 1387 14093 1421 14096
rect 3691 14310 3725 14344
rect 2466 14199 2500 14233
rect 2562 14199 2596 14233
rect 2658 14199 2692 14233
rect 2754 14199 2788 14233
rect 2850 14199 2884 14233
rect 2946 14199 2980 14233
rect 3042 14199 3076 14233
rect 3138 14199 3172 14233
rect 3234 14199 3268 14233
rect 3330 14199 3364 14233
rect 3426 14199 3460 14233
rect 3540 14270 3574 14275
rect 3540 14241 3574 14270
rect 3540 14202 3574 14203
rect 3540 14169 3574 14202
rect 3647 14184 3681 14260
rect 3735 14184 3769 14260
rect 2466 14088 2500 14122
rect 2658 14088 2692 14122
rect 2850 14088 2884 14122
rect 3042 14088 3076 14122
rect 3234 14088 3268 14122
rect 3426 14088 3460 14122
rect 3540 14100 3574 14131
rect 3540 14097 3574 14100
rect 3987 14199 4021 14233
rect 4083 14199 4117 14233
rect 4179 14199 4213 14233
rect 4275 14199 4309 14233
rect 4371 14199 4405 14233
rect 4467 14199 4501 14233
rect 4563 14199 4597 14233
rect 4659 14199 4693 14233
rect 4755 14199 4789 14233
rect 4851 14199 4885 14233
rect 4947 14199 4981 14233
rect 5061 14270 5095 14275
rect 5061 14241 5095 14270
rect 5061 14202 5095 14203
rect 5061 14169 5095 14202
rect 5348 14351 5382 14385
rect 5450 14387 5484 14390
rect 5450 14356 5470 14387
rect 5470 14356 5484 14387
rect 3987 14088 4021 14122
rect 4179 14088 4213 14122
rect 4371 14088 4405 14122
rect 4563 14088 4597 14122
rect 4755 14088 4789 14122
rect 4947 14088 4981 14122
rect 5061 14100 5095 14131
rect 5303 14121 5337 14155
rect 5395 14121 5429 14155
rect 5487 14121 5521 14155
rect 5061 14097 5095 14100
rect 313 13605 347 13639
rect 505 13605 539 13639
rect 697 13605 731 13639
rect 889 13605 923 13639
rect 1081 13605 1115 13639
rect 1273 13605 1307 13639
rect 1387 13605 1421 13613
rect 1387 13579 1421 13605
rect 313 13506 347 13510
rect 313 13476 347 13506
rect 313 13404 347 13438
rect 313 13336 347 13366
rect 313 13332 347 13336
rect 409 13506 443 13510
rect 409 13476 443 13506
rect 409 13404 443 13438
rect 409 13336 443 13366
rect 409 13332 443 13336
rect 505 13506 539 13510
rect 505 13476 539 13506
rect 505 13404 539 13438
rect 505 13336 539 13366
rect 505 13332 539 13336
rect 601 13506 635 13510
rect 601 13476 635 13506
rect 601 13404 635 13438
rect 601 13336 635 13366
rect 601 13332 635 13336
rect 697 13506 731 13510
rect 697 13476 731 13506
rect 697 13404 731 13438
rect 697 13336 731 13366
rect 697 13332 731 13336
rect 793 13506 827 13510
rect 793 13476 827 13506
rect 793 13404 827 13438
rect 793 13336 827 13366
rect 793 13332 827 13336
rect 889 13506 923 13510
rect 889 13476 923 13506
rect 889 13404 923 13438
rect 889 13336 923 13366
rect 889 13332 923 13336
rect 985 13506 1019 13510
rect 985 13476 1019 13506
rect 985 13404 1019 13438
rect 985 13336 1019 13366
rect 985 13332 1019 13336
rect 1081 13506 1115 13510
rect 1081 13476 1115 13506
rect 1081 13404 1115 13438
rect 1081 13336 1115 13366
rect 1081 13332 1115 13336
rect 1177 13506 1211 13510
rect 1177 13476 1211 13506
rect 1177 13404 1211 13438
rect 1177 13336 1211 13366
rect 1177 13332 1211 13336
rect 1273 13506 1307 13510
rect 1273 13476 1307 13506
rect 1273 13404 1307 13438
rect 1273 13336 1307 13366
rect 1273 13332 1307 13336
rect 1387 13537 1421 13541
rect 1387 13507 1421 13537
rect 1387 13435 1421 13469
rect 1387 13367 1421 13397
rect 1387 13363 1421 13367
rect 1387 13299 1421 13325
rect 1387 13291 1421 13299
rect 2466 13609 2500 13643
rect 2658 13609 2692 13643
rect 2850 13609 2884 13643
rect 3042 13609 3076 13643
rect 3234 13609 3268 13643
rect 3426 13609 3460 13643
rect 3540 13609 3574 13617
rect 3540 13583 3574 13609
rect 2466 13510 2500 13514
rect 2466 13480 2500 13510
rect 2466 13408 2500 13442
rect 2466 13340 2500 13370
rect 2466 13336 2500 13340
rect 2562 13510 2596 13514
rect 2562 13480 2596 13510
rect 2562 13408 2596 13442
rect 2562 13340 2596 13370
rect 2562 13336 2596 13340
rect 2658 13510 2692 13514
rect 2658 13480 2692 13510
rect 2658 13408 2692 13442
rect 2658 13340 2692 13370
rect 2658 13336 2692 13340
rect 2754 13510 2788 13514
rect 2754 13480 2788 13510
rect 2754 13408 2788 13442
rect 2754 13340 2788 13370
rect 2754 13336 2788 13340
rect 2850 13510 2884 13514
rect 2850 13480 2884 13510
rect 2850 13408 2884 13442
rect 2850 13340 2884 13370
rect 2850 13336 2884 13340
rect 2946 13510 2980 13514
rect 2946 13480 2980 13510
rect 2946 13408 2980 13442
rect 2946 13340 2980 13370
rect 2946 13336 2980 13340
rect 3042 13510 3076 13514
rect 3042 13480 3076 13510
rect 3042 13408 3076 13442
rect 3042 13340 3076 13370
rect 3042 13336 3076 13340
rect 3138 13510 3172 13514
rect 3138 13480 3172 13510
rect 3138 13408 3172 13442
rect 3138 13340 3172 13370
rect 3138 13336 3172 13340
rect 3234 13510 3268 13514
rect 3234 13480 3268 13510
rect 3234 13408 3268 13442
rect 3234 13340 3268 13370
rect 3234 13336 3268 13340
rect 3330 13510 3364 13514
rect 3330 13480 3364 13510
rect 3330 13408 3364 13442
rect 3330 13340 3364 13370
rect 3330 13336 3364 13340
rect 3426 13510 3460 13514
rect 3426 13480 3460 13510
rect 3426 13408 3460 13442
rect 3426 13340 3460 13370
rect 3426 13336 3460 13340
rect 3540 13541 3574 13545
rect 3540 13511 3574 13541
rect 3540 13439 3574 13473
rect 3540 13371 3574 13401
rect 3540 13367 3574 13371
rect 3540 13303 3574 13329
rect 3540 13295 3574 13303
rect 3987 13609 4021 13643
rect 4179 13609 4213 13643
rect 4371 13609 4405 13643
rect 4563 13609 4597 13643
rect 4755 13609 4789 13643
rect 4947 13609 4981 13643
rect 5061 13609 5095 13617
rect 5061 13583 5095 13609
rect 3987 13510 4021 13514
rect 3987 13480 4021 13510
rect 3987 13408 4021 13442
rect 3987 13340 4021 13370
rect 3987 13336 4021 13340
rect 4083 13510 4117 13514
rect 4083 13480 4117 13510
rect 4083 13408 4117 13442
rect 4083 13340 4117 13370
rect 4083 13336 4117 13340
rect 4179 13510 4213 13514
rect 4179 13480 4213 13510
rect 4179 13408 4213 13442
rect 4179 13340 4213 13370
rect 4179 13336 4213 13340
rect 4275 13510 4309 13514
rect 4275 13480 4309 13510
rect 4275 13408 4309 13442
rect 4275 13340 4309 13370
rect 4275 13336 4309 13340
rect 4371 13510 4405 13514
rect 4371 13480 4405 13510
rect 4371 13408 4405 13442
rect 4371 13340 4405 13370
rect 4371 13336 4405 13340
rect 4467 13510 4501 13514
rect 4467 13480 4501 13510
rect 4467 13408 4501 13442
rect 4467 13340 4501 13370
rect 4467 13336 4501 13340
rect 4563 13510 4597 13514
rect 4563 13480 4597 13510
rect 4563 13408 4597 13442
rect 4563 13340 4597 13370
rect 4563 13336 4597 13340
rect 4659 13510 4693 13514
rect 4659 13480 4693 13510
rect 4659 13408 4693 13442
rect 4659 13340 4693 13370
rect 4659 13336 4693 13340
rect 4755 13510 4789 13514
rect 4755 13480 4789 13510
rect 4755 13408 4789 13442
rect 4755 13340 4789 13370
rect 4755 13336 4789 13340
rect 4851 13510 4885 13514
rect 4851 13480 4885 13510
rect 4851 13408 4885 13442
rect 4851 13340 4885 13370
rect 4851 13336 4885 13340
rect 4947 13510 4981 13514
rect 4947 13480 4981 13510
rect 4947 13408 4981 13442
rect 4947 13340 4981 13370
rect 4947 13336 4981 13340
rect 5061 13541 5095 13545
rect 5061 13511 5095 13541
rect 5061 13439 5095 13473
rect 5061 13371 5095 13401
rect 5303 13378 5337 13412
rect 5395 13378 5429 13412
rect 5487 13378 5521 13412
rect 5061 13367 5095 13371
rect 5061 13303 5095 13329
rect 5061 13295 5095 13303
rect 313 12908 347 12942
rect 409 12908 443 12942
rect 505 12908 539 12942
rect 601 12908 635 12942
rect 697 12908 731 12942
rect 793 12908 827 12942
rect 889 12908 923 12942
rect 985 12908 1019 12942
rect 1081 12908 1115 12942
rect 1177 12908 1211 12942
rect 1273 12908 1307 12942
rect 1387 12979 1421 12984
rect 1387 12950 1421 12979
rect 1387 12911 1421 12912
rect 1387 12878 1421 12911
rect 313 12797 347 12831
rect 505 12797 539 12831
rect 697 12797 731 12831
rect 889 12797 923 12831
rect 1081 12797 1115 12831
rect 1273 12797 1307 12831
rect 1387 12809 1421 12840
rect 1387 12806 1421 12809
rect 3691 13023 3725 13057
rect 2466 12912 2500 12946
rect 2562 12912 2596 12946
rect 2658 12912 2692 12946
rect 2754 12912 2788 12946
rect 2850 12912 2884 12946
rect 2946 12912 2980 12946
rect 3042 12912 3076 12946
rect 3138 12912 3172 12946
rect 3234 12912 3268 12946
rect 3330 12912 3364 12946
rect 3426 12912 3460 12946
rect 3540 12983 3574 12988
rect 3540 12954 3574 12983
rect 3540 12915 3574 12916
rect 3540 12882 3574 12915
rect 3647 12897 3681 12973
rect 3735 12897 3769 12973
rect 2466 12801 2500 12835
rect 2658 12801 2692 12835
rect 2850 12801 2884 12835
rect 3042 12801 3076 12835
rect 3234 12801 3268 12835
rect 3426 12801 3460 12835
rect 3540 12813 3574 12844
rect 3540 12810 3574 12813
rect 3987 12912 4021 12946
rect 4083 12912 4117 12946
rect 4179 12912 4213 12946
rect 4275 12912 4309 12946
rect 4371 12912 4405 12946
rect 4467 12912 4501 12946
rect 4563 12912 4597 12946
rect 4659 12912 4693 12946
rect 4755 12912 4789 12946
rect 4851 12912 4885 12946
rect 4947 12912 4981 12946
rect 5061 12983 5095 12988
rect 5061 12954 5095 12983
rect 5061 12915 5095 12916
rect 5061 12882 5095 12915
rect 5348 13064 5382 13098
rect 5450 13100 5484 13103
rect 5450 13069 5470 13100
rect 5470 13069 5484 13100
rect 3987 12801 4021 12835
rect 4179 12801 4213 12835
rect 4371 12801 4405 12835
rect 4563 12801 4597 12835
rect 4755 12801 4789 12835
rect 4947 12801 4981 12835
rect 5061 12813 5095 12844
rect 5303 12834 5337 12868
rect 5395 12834 5429 12868
rect 5487 12834 5521 12868
rect 5061 12810 5095 12813
rect 313 12318 347 12352
rect 505 12318 539 12352
rect 697 12318 731 12352
rect 889 12318 923 12352
rect 1081 12318 1115 12352
rect 1273 12318 1307 12352
rect 1387 12318 1421 12326
rect 1387 12292 1421 12318
rect 313 12219 347 12223
rect 313 12189 347 12219
rect 313 12117 347 12151
rect 313 12049 347 12079
rect 313 12045 347 12049
rect 409 12219 443 12223
rect 409 12189 443 12219
rect 409 12117 443 12151
rect 409 12049 443 12079
rect 409 12045 443 12049
rect 505 12219 539 12223
rect 505 12189 539 12219
rect 505 12117 539 12151
rect 505 12049 539 12079
rect 505 12045 539 12049
rect 601 12219 635 12223
rect 601 12189 635 12219
rect 601 12117 635 12151
rect 601 12049 635 12079
rect 601 12045 635 12049
rect 697 12219 731 12223
rect 697 12189 731 12219
rect 697 12117 731 12151
rect 697 12049 731 12079
rect 697 12045 731 12049
rect 793 12219 827 12223
rect 793 12189 827 12219
rect 793 12117 827 12151
rect 793 12049 827 12079
rect 793 12045 827 12049
rect 889 12219 923 12223
rect 889 12189 923 12219
rect 889 12117 923 12151
rect 889 12049 923 12079
rect 889 12045 923 12049
rect 985 12219 1019 12223
rect 985 12189 1019 12219
rect 985 12117 1019 12151
rect 985 12049 1019 12079
rect 985 12045 1019 12049
rect 1081 12219 1115 12223
rect 1081 12189 1115 12219
rect 1081 12117 1115 12151
rect 1081 12049 1115 12079
rect 1081 12045 1115 12049
rect 1177 12219 1211 12223
rect 1177 12189 1211 12219
rect 1177 12117 1211 12151
rect 1177 12049 1211 12079
rect 1177 12045 1211 12049
rect 1273 12219 1307 12223
rect 1273 12189 1307 12219
rect 1273 12117 1307 12151
rect 1273 12049 1307 12079
rect 1273 12045 1307 12049
rect 1387 12250 1421 12254
rect 1387 12220 1421 12250
rect 1387 12148 1421 12182
rect 1387 12080 1421 12110
rect 1387 12076 1421 12080
rect 1387 12012 1421 12038
rect 1387 12004 1421 12012
rect 2466 12322 2500 12356
rect 2658 12322 2692 12356
rect 2850 12322 2884 12356
rect 3042 12322 3076 12356
rect 3234 12322 3268 12356
rect 3426 12322 3460 12356
rect 3540 12322 3574 12330
rect 3540 12296 3574 12322
rect 2466 12223 2500 12227
rect 2466 12193 2500 12223
rect 2466 12121 2500 12155
rect 2466 12053 2500 12083
rect 2466 12049 2500 12053
rect 2562 12223 2596 12227
rect 2562 12193 2596 12223
rect 2562 12121 2596 12155
rect 2562 12053 2596 12083
rect 2562 12049 2596 12053
rect 2658 12223 2692 12227
rect 2658 12193 2692 12223
rect 2658 12121 2692 12155
rect 2658 12053 2692 12083
rect 2658 12049 2692 12053
rect 2754 12223 2788 12227
rect 2754 12193 2788 12223
rect 2754 12121 2788 12155
rect 2754 12053 2788 12083
rect 2754 12049 2788 12053
rect 2850 12223 2884 12227
rect 2850 12193 2884 12223
rect 2850 12121 2884 12155
rect 2850 12053 2884 12083
rect 2850 12049 2884 12053
rect 2946 12223 2980 12227
rect 2946 12193 2980 12223
rect 2946 12121 2980 12155
rect 2946 12053 2980 12083
rect 2946 12049 2980 12053
rect 3042 12223 3076 12227
rect 3042 12193 3076 12223
rect 3042 12121 3076 12155
rect 3042 12053 3076 12083
rect 3042 12049 3076 12053
rect 3138 12223 3172 12227
rect 3138 12193 3172 12223
rect 3138 12121 3172 12155
rect 3138 12053 3172 12083
rect 3138 12049 3172 12053
rect 3234 12223 3268 12227
rect 3234 12193 3268 12223
rect 3234 12121 3268 12155
rect 3234 12053 3268 12083
rect 3234 12049 3268 12053
rect 3330 12223 3364 12227
rect 3330 12193 3364 12223
rect 3330 12121 3364 12155
rect 3330 12053 3364 12083
rect 3330 12049 3364 12053
rect 3426 12223 3460 12227
rect 3426 12193 3460 12223
rect 3426 12121 3460 12155
rect 3426 12053 3460 12083
rect 3426 12049 3460 12053
rect 3540 12254 3574 12258
rect 3540 12224 3574 12254
rect 3540 12152 3574 12186
rect 3540 12084 3574 12114
rect 3540 12080 3574 12084
rect 3540 12016 3574 12042
rect 3540 12008 3574 12016
rect 3987 12322 4021 12356
rect 4179 12322 4213 12356
rect 4371 12322 4405 12356
rect 4563 12322 4597 12356
rect 4755 12322 4789 12356
rect 4947 12322 4981 12356
rect 5061 12322 5095 12330
rect 5061 12296 5095 12322
rect 3987 12223 4021 12227
rect 3987 12193 4021 12223
rect 3987 12121 4021 12155
rect 3987 12053 4021 12083
rect 3987 12049 4021 12053
rect 4083 12223 4117 12227
rect 4083 12193 4117 12223
rect 4083 12121 4117 12155
rect 4083 12053 4117 12083
rect 4083 12049 4117 12053
rect 4179 12223 4213 12227
rect 4179 12193 4213 12223
rect 4179 12121 4213 12155
rect 4179 12053 4213 12083
rect 4179 12049 4213 12053
rect 4275 12223 4309 12227
rect 4275 12193 4309 12223
rect 4275 12121 4309 12155
rect 4275 12053 4309 12083
rect 4275 12049 4309 12053
rect 4371 12223 4405 12227
rect 4371 12193 4405 12223
rect 4371 12121 4405 12155
rect 4371 12053 4405 12083
rect 4371 12049 4405 12053
rect 4467 12223 4501 12227
rect 4467 12193 4501 12223
rect 4467 12121 4501 12155
rect 4467 12053 4501 12083
rect 4467 12049 4501 12053
rect 4563 12223 4597 12227
rect 4563 12193 4597 12223
rect 4563 12121 4597 12155
rect 4563 12053 4597 12083
rect 4563 12049 4597 12053
rect 4659 12223 4693 12227
rect 4659 12193 4693 12223
rect 4659 12121 4693 12155
rect 4659 12053 4693 12083
rect 4659 12049 4693 12053
rect 4755 12223 4789 12227
rect 4755 12193 4789 12223
rect 4755 12121 4789 12155
rect 4755 12053 4789 12083
rect 4755 12049 4789 12053
rect 4851 12223 4885 12227
rect 4851 12193 4885 12223
rect 4851 12121 4885 12155
rect 4851 12053 4885 12083
rect 4851 12049 4885 12053
rect 4947 12223 4981 12227
rect 4947 12193 4981 12223
rect 4947 12121 4981 12155
rect 4947 12053 4981 12083
rect 4947 12049 4981 12053
rect 5061 12254 5095 12258
rect 5061 12224 5095 12254
rect 5061 12152 5095 12186
rect 5061 12084 5095 12114
rect 5303 12091 5337 12125
rect 5395 12091 5429 12125
rect 5487 12091 5521 12125
rect 5061 12080 5095 12084
rect 5061 12016 5095 12042
rect 5061 12008 5095 12016
rect 313 11621 347 11655
rect 409 11621 443 11655
rect 505 11621 539 11655
rect 601 11621 635 11655
rect 697 11621 731 11655
rect 793 11621 827 11655
rect 889 11621 923 11655
rect 985 11621 1019 11655
rect 1081 11621 1115 11655
rect 1177 11621 1211 11655
rect 1273 11621 1307 11655
rect 1387 11692 1421 11697
rect 1387 11663 1421 11692
rect 1387 11624 1421 11625
rect 1387 11591 1421 11624
rect 313 11510 347 11544
rect 505 11510 539 11544
rect 697 11510 731 11544
rect 889 11510 923 11544
rect 1081 11510 1115 11544
rect 1273 11510 1307 11544
rect 1387 11522 1421 11553
rect 1387 11519 1421 11522
rect 3691 11736 3725 11770
rect 2466 11625 2500 11659
rect 2562 11625 2596 11659
rect 2658 11625 2692 11659
rect 2754 11625 2788 11659
rect 2850 11625 2884 11659
rect 2946 11625 2980 11659
rect 3042 11625 3076 11659
rect 3138 11625 3172 11659
rect 3234 11625 3268 11659
rect 3330 11625 3364 11659
rect 3426 11625 3460 11659
rect 3540 11696 3574 11701
rect 3540 11667 3574 11696
rect 3540 11628 3574 11629
rect 3540 11595 3574 11628
rect 3647 11610 3681 11686
rect 3735 11610 3769 11686
rect 2466 11514 2500 11548
rect 2658 11514 2692 11548
rect 2850 11514 2884 11548
rect 3042 11514 3076 11548
rect 3234 11514 3268 11548
rect 3426 11514 3460 11548
rect 3540 11526 3574 11557
rect 3540 11523 3574 11526
rect 3987 11625 4021 11659
rect 4083 11625 4117 11659
rect 4179 11625 4213 11659
rect 4275 11625 4309 11659
rect 4371 11625 4405 11659
rect 4467 11625 4501 11659
rect 4563 11625 4597 11659
rect 4659 11625 4693 11659
rect 4755 11625 4789 11659
rect 4851 11625 4885 11659
rect 4947 11625 4981 11659
rect 5061 11696 5095 11701
rect 5061 11667 5095 11696
rect 5061 11628 5095 11629
rect 5061 11595 5095 11628
rect 5348 11777 5382 11811
rect 5450 11813 5484 11816
rect 5450 11782 5470 11813
rect 5470 11782 5484 11813
rect 3987 11514 4021 11548
rect 4179 11514 4213 11548
rect 4371 11514 4405 11548
rect 4563 11514 4597 11548
rect 4755 11514 4789 11548
rect 4947 11514 4981 11548
rect 5061 11526 5095 11557
rect 5303 11547 5337 11581
rect 5395 11547 5429 11581
rect 5487 11547 5521 11581
rect 5061 11523 5095 11526
rect 313 11031 347 11065
rect 505 11031 539 11065
rect 697 11031 731 11065
rect 889 11031 923 11065
rect 1081 11031 1115 11065
rect 1273 11031 1307 11065
rect 1387 11031 1421 11039
rect 1387 11005 1421 11031
rect 313 10932 347 10936
rect 313 10902 347 10932
rect 313 10830 347 10864
rect 313 10762 347 10792
rect 313 10758 347 10762
rect 409 10932 443 10936
rect 409 10902 443 10932
rect 409 10830 443 10864
rect 409 10762 443 10792
rect 409 10758 443 10762
rect 505 10932 539 10936
rect 505 10902 539 10932
rect 505 10830 539 10864
rect 505 10762 539 10792
rect 505 10758 539 10762
rect 601 10932 635 10936
rect 601 10902 635 10932
rect 601 10830 635 10864
rect 601 10762 635 10792
rect 601 10758 635 10762
rect 697 10932 731 10936
rect 697 10902 731 10932
rect 697 10830 731 10864
rect 697 10762 731 10792
rect 697 10758 731 10762
rect 793 10932 827 10936
rect 793 10902 827 10932
rect 793 10830 827 10864
rect 793 10762 827 10792
rect 793 10758 827 10762
rect 889 10932 923 10936
rect 889 10902 923 10932
rect 889 10830 923 10864
rect 889 10762 923 10792
rect 889 10758 923 10762
rect 985 10932 1019 10936
rect 985 10902 1019 10932
rect 985 10830 1019 10864
rect 985 10762 1019 10792
rect 985 10758 1019 10762
rect 1081 10932 1115 10936
rect 1081 10902 1115 10932
rect 1081 10830 1115 10864
rect 1081 10762 1115 10792
rect 1081 10758 1115 10762
rect 1177 10932 1211 10936
rect 1177 10902 1211 10932
rect 1177 10830 1211 10864
rect 1177 10762 1211 10792
rect 1177 10758 1211 10762
rect 1273 10932 1307 10936
rect 1273 10902 1307 10932
rect 1273 10830 1307 10864
rect 1273 10762 1307 10792
rect 1273 10758 1307 10762
rect 1387 10963 1421 10967
rect 1387 10933 1421 10963
rect 1387 10861 1421 10895
rect 1387 10793 1421 10823
rect 1387 10789 1421 10793
rect 1387 10725 1421 10751
rect 1387 10717 1421 10725
rect 2466 11035 2500 11069
rect 2658 11035 2692 11069
rect 2850 11035 2884 11069
rect 3042 11035 3076 11069
rect 3234 11035 3268 11069
rect 3426 11035 3460 11069
rect 3540 11035 3574 11043
rect 3540 11009 3574 11035
rect 2466 10936 2500 10940
rect 2466 10906 2500 10936
rect 2466 10834 2500 10868
rect 2466 10766 2500 10796
rect 2466 10762 2500 10766
rect 2562 10936 2596 10940
rect 2562 10906 2596 10936
rect 2562 10834 2596 10868
rect 2562 10766 2596 10796
rect 2562 10762 2596 10766
rect 2658 10936 2692 10940
rect 2658 10906 2692 10936
rect 2658 10834 2692 10868
rect 2658 10766 2692 10796
rect 2658 10762 2692 10766
rect 2754 10936 2788 10940
rect 2754 10906 2788 10936
rect 2754 10834 2788 10868
rect 2754 10766 2788 10796
rect 2754 10762 2788 10766
rect 2850 10936 2884 10940
rect 2850 10906 2884 10936
rect 2850 10834 2884 10868
rect 2850 10766 2884 10796
rect 2850 10762 2884 10766
rect 2946 10936 2980 10940
rect 2946 10906 2980 10936
rect 2946 10834 2980 10868
rect 2946 10766 2980 10796
rect 2946 10762 2980 10766
rect 3042 10936 3076 10940
rect 3042 10906 3076 10936
rect 3042 10834 3076 10868
rect 3042 10766 3076 10796
rect 3042 10762 3076 10766
rect 3138 10936 3172 10940
rect 3138 10906 3172 10936
rect 3138 10834 3172 10868
rect 3138 10766 3172 10796
rect 3138 10762 3172 10766
rect 3234 10936 3268 10940
rect 3234 10906 3268 10936
rect 3234 10834 3268 10868
rect 3234 10766 3268 10796
rect 3234 10762 3268 10766
rect 3330 10936 3364 10940
rect 3330 10906 3364 10936
rect 3330 10834 3364 10868
rect 3330 10766 3364 10796
rect 3330 10762 3364 10766
rect 3426 10936 3460 10940
rect 3426 10906 3460 10936
rect 3426 10834 3460 10868
rect 3426 10766 3460 10796
rect 3426 10762 3460 10766
rect 3540 10967 3574 10971
rect 3540 10937 3574 10967
rect 3540 10865 3574 10899
rect 3540 10797 3574 10827
rect 3540 10793 3574 10797
rect 3540 10729 3574 10755
rect 3540 10721 3574 10729
rect 3987 11035 4021 11069
rect 4179 11035 4213 11069
rect 4371 11035 4405 11069
rect 4563 11035 4597 11069
rect 4755 11035 4789 11069
rect 4947 11035 4981 11069
rect 5061 11035 5095 11043
rect 5061 11009 5095 11035
rect 3987 10936 4021 10940
rect 3987 10906 4021 10936
rect 3987 10834 4021 10868
rect 3987 10766 4021 10796
rect 3987 10762 4021 10766
rect 4083 10936 4117 10940
rect 4083 10906 4117 10936
rect 4083 10834 4117 10868
rect 4083 10766 4117 10796
rect 4083 10762 4117 10766
rect 4179 10936 4213 10940
rect 4179 10906 4213 10936
rect 4179 10834 4213 10868
rect 4179 10766 4213 10796
rect 4179 10762 4213 10766
rect 4275 10936 4309 10940
rect 4275 10906 4309 10936
rect 4275 10834 4309 10868
rect 4275 10766 4309 10796
rect 4275 10762 4309 10766
rect 4371 10936 4405 10940
rect 4371 10906 4405 10936
rect 4371 10834 4405 10868
rect 4371 10766 4405 10796
rect 4371 10762 4405 10766
rect 4467 10936 4501 10940
rect 4467 10906 4501 10936
rect 4467 10834 4501 10868
rect 4467 10766 4501 10796
rect 4467 10762 4501 10766
rect 4563 10936 4597 10940
rect 4563 10906 4597 10936
rect 4563 10834 4597 10868
rect 4563 10766 4597 10796
rect 4563 10762 4597 10766
rect 4659 10936 4693 10940
rect 4659 10906 4693 10936
rect 4659 10834 4693 10868
rect 4659 10766 4693 10796
rect 4659 10762 4693 10766
rect 4755 10936 4789 10940
rect 4755 10906 4789 10936
rect 4755 10834 4789 10868
rect 4755 10766 4789 10796
rect 4755 10762 4789 10766
rect 4851 10936 4885 10940
rect 4851 10906 4885 10936
rect 4851 10834 4885 10868
rect 4851 10766 4885 10796
rect 4851 10762 4885 10766
rect 4947 10936 4981 10940
rect 4947 10906 4981 10936
rect 4947 10834 4981 10868
rect 4947 10766 4981 10796
rect 4947 10762 4981 10766
rect 5061 10967 5095 10971
rect 5061 10937 5095 10967
rect 5061 10865 5095 10899
rect 5061 10797 5095 10827
rect 5303 10804 5337 10838
rect 5395 10804 5429 10838
rect 5487 10804 5521 10838
rect 5061 10793 5095 10797
rect 5061 10729 5095 10755
rect 5061 10721 5095 10729
rect 313 10334 347 10368
rect 409 10334 443 10368
rect 505 10334 539 10368
rect 601 10334 635 10368
rect 697 10334 731 10368
rect 793 10334 827 10368
rect 889 10334 923 10368
rect 985 10334 1019 10368
rect 1081 10334 1115 10368
rect 1177 10334 1211 10368
rect 1273 10334 1307 10368
rect 1387 10405 1421 10410
rect 1387 10376 1421 10405
rect 1387 10337 1421 10338
rect 1387 10304 1421 10337
rect 313 10223 347 10257
rect 505 10223 539 10257
rect 697 10223 731 10257
rect 889 10223 923 10257
rect 1081 10223 1115 10257
rect 1273 10223 1307 10257
rect 1387 10235 1421 10266
rect 1387 10232 1421 10235
rect 3691 10449 3725 10483
rect 2466 10338 2500 10372
rect 2562 10338 2596 10372
rect 2658 10338 2692 10372
rect 2754 10338 2788 10372
rect 2850 10338 2884 10372
rect 2946 10338 2980 10372
rect 3042 10338 3076 10372
rect 3138 10338 3172 10372
rect 3234 10338 3268 10372
rect 3330 10338 3364 10372
rect 3426 10338 3460 10372
rect 3540 10409 3574 10414
rect 3540 10380 3574 10409
rect 3540 10341 3574 10342
rect 3540 10308 3574 10341
rect 3647 10323 3681 10399
rect 3735 10323 3769 10399
rect 2466 10227 2500 10261
rect 2658 10227 2692 10261
rect 2850 10227 2884 10261
rect 3042 10227 3076 10261
rect 3234 10227 3268 10261
rect 3426 10227 3460 10261
rect 3540 10239 3574 10270
rect 3540 10236 3574 10239
rect 3987 10338 4021 10372
rect 4083 10338 4117 10372
rect 4179 10338 4213 10372
rect 4275 10338 4309 10372
rect 4371 10338 4405 10372
rect 4467 10338 4501 10372
rect 4563 10338 4597 10372
rect 4659 10338 4693 10372
rect 4755 10338 4789 10372
rect 4851 10338 4885 10372
rect 4947 10338 4981 10372
rect 5061 10409 5095 10414
rect 5061 10380 5095 10409
rect 5061 10341 5095 10342
rect 5061 10308 5095 10341
rect 5348 10490 5382 10524
rect 5450 10526 5484 10529
rect 5450 10495 5470 10526
rect 5470 10495 5484 10526
rect 3987 10227 4021 10261
rect 4179 10227 4213 10261
rect 4371 10227 4405 10261
rect 4563 10227 4597 10261
rect 4755 10227 4789 10261
rect 4947 10227 4981 10261
rect 5061 10239 5095 10270
rect 5303 10260 5337 10294
rect 5395 10260 5429 10294
rect 5487 10260 5521 10294
rect 5061 10236 5095 10239
rect 313 9744 347 9778
rect 505 9744 539 9778
rect 697 9744 731 9778
rect 889 9744 923 9778
rect 1081 9744 1115 9778
rect 1273 9744 1307 9778
rect 1387 9744 1421 9752
rect 1387 9718 1421 9744
rect 313 9645 347 9649
rect 313 9615 347 9645
rect 313 9543 347 9577
rect 313 9475 347 9505
rect 313 9471 347 9475
rect 409 9645 443 9649
rect 409 9615 443 9645
rect 409 9543 443 9577
rect 409 9475 443 9505
rect 409 9471 443 9475
rect 505 9645 539 9649
rect 505 9615 539 9645
rect 505 9543 539 9577
rect 505 9475 539 9505
rect 505 9471 539 9475
rect 601 9645 635 9649
rect 601 9615 635 9645
rect 601 9543 635 9577
rect 601 9475 635 9505
rect 601 9471 635 9475
rect 697 9645 731 9649
rect 697 9615 731 9645
rect 697 9543 731 9577
rect 697 9475 731 9505
rect 697 9471 731 9475
rect 793 9645 827 9649
rect 793 9615 827 9645
rect 793 9543 827 9577
rect 793 9475 827 9505
rect 793 9471 827 9475
rect 889 9645 923 9649
rect 889 9615 923 9645
rect 889 9543 923 9577
rect 889 9475 923 9505
rect 889 9471 923 9475
rect 985 9645 1019 9649
rect 985 9615 1019 9645
rect 985 9543 1019 9577
rect 985 9475 1019 9505
rect 985 9471 1019 9475
rect 1081 9645 1115 9649
rect 1081 9615 1115 9645
rect 1081 9543 1115 9577
rect 1081 9475 1115 9505
rect 1081 9471 1115 9475
rect 1177 9645 1211 9649
rect 1177 9615 1211 9645
rect 1177 9543 1211 9577
rect 1177 9475 1211 9505
rect 1177 9471 1211 9475
rect 1273 9645 1307 9649
rect 1273 9615 1307 9645
rect 1273 9543 1307 9577
rect 1273 9475 1307 9505
rect 1273 9471 1307 9475
rect 1387 9676 1421 9680
rect 1387 9646 1421 9676
rect 1387 9574 1421 9608
rect 1387 9506 1421 9536
rect 1387 9502 1421 9506
rect 1387 9438 1421 9464
rect 1387 9430 1421 9438
rect 2466 9748 2500 9782
rect 2658 9748 2692 9782
rect 2850 9748 2884 9782
rect 3042 9748 3076 9782
rect 3234 9748 3268 9782
rect 3426 9748 3460 9782
rect 3540 9748 3574 9756
rect 3540 9722 3574 9748
rect 2466 9649 2500 9653
rect 2466 9619 2500 9649
rect 2466 9547 2500 9581
rect 2466 9479 2500 9509
rect 2466 9475 2500 9479
rect 2562 9649 2596 9653
rect 2562 9619 2596 9649
rect 2562 9547 2596 9581
rect 2562 9479 2596 9509
rect 2562 9475 2596 9479
rect 2658 9649 2692 9653
rect 2658 9619 2692 9649
rect 2658 9547 2692 9581
rect 2658 9479 2692 9509
rect 2658 9475 2692 9479
rect 2754 9649 2788 9653
rect 2754 9619 2788 9649
rect 2754 9547 2788 9581
rect 2754 9479 2788 9509
rect 2754 9475 2788 9479
rect 2850 9649 2884 9653
rect 2850 9619 2884 9649
rect 2850 9547 2884 9581
rect 2850 9479 2884 9509
rect 2850 9475 2884 9479
rect 2946 9649 2980 9653
rect 2946 9619 2980 9649
rect 2946 9547 2980 9581
rect 2946 9479 2980 9509
rect 2946 9475 2980 9479
rect 3042 9649 3076 9653
rect 3042 9619 3076 9649
rect 3042 9547 3076 9581
rect 3042 9479 3076 9509
rect 3042 9475 3076 9479
rect 3138 9649 3172 9653
rect 3138 9619 3172 9649
rect 3138 9547 3172 9581
rect 3138 9479 3172 9509
rect 3138 9475 3172 9479
rect 3234 9649 3268 9653
rect 3234 9619 3268 9649
rect 3234 9547 3268 9581
rect 3234 9479 3268 9509
rect 3234 9475 3268 9479
rect 3330 9649 3364 9653
rect 3330 9619 3364 9649
rect 3330 9547 3364 9581
rect 3330 9479 3364 9509
rect 3330 9475 3364 9479
rect 3426 9649 3460 9653
rect 3426 9619 3460 9649
rect 3426 9547 3460 9581
rect 3426 9479 3460 9509
rect 3426 9475 3460 9479
rect 3540 9680 3574 9684
rect 3540 9650 3574 9680
rect 3540 9578 3574 9612
rect 3540 9510 3574 9540
rect 3540 9506 3574 9510
rect 3540 9442 3574 9468
rect 3540 9434 3574 9442
rect 3987 9748 4021 9782
rect 4179 9748 4213 9782
rect 4371 9748 4405 9782
rect 4563 9748 4597 9782
rect 4755 9748 4789 9782
rect 4947 9748 4981 9782
rect 5061 9748 5095 9756
rect 5061 9722 5095 9748
rect 3987 9649 4021 9653
rect 3987 9619 4021 9649
rect 3987 9547 4021 9581
rect 3987 9479 4021 9509
rect 3987 9475 4021 9479
rect 4083 9649 4117 9653
rect 4083 9619 4117 9649
rect 4083 9547 4117 9581
rect 4083 9479 4117 9509
rect 4083 9475 4117 9479
rect 4179 9649 4213 9653
rect 4179 9619 4213 9649
rect 4179 9547 4213 9581
rect 4179 9479 4213 9509
rect 4179 9475 4213 9479
rect 4275 9649 4309 9653
rect 4275 9619 4309 9649
rect 4275 9547 4309 9581
rect 4275 9479 4309 9509
rect 4275 9475 4309 9479
rect 4371 9649 4405 9653
rect 4371 9619 4405 9649
rect 4371 9547 4405 9581
rect 4371 9479 4405 9509
rect 4371 9475 4405 9479
rect 4467 9649 4501 9653
rect 4467 9619 4501 9649
rect 4467 9547 4501 9581
rect 4467 9479 4501 9509
rect 4467 9475 4501 9479
rect 4563 9649 4597 9653
rect 4563 9619 4597 9649
rect 4563 9547 4597 9581
rect 4563 9479 4597 9509
rect 4563 9475 4597 9479
rect 4659 9649 4693 9653
rect 4659 9619 4693 9649
rect 4659 9547 4693 9581
rect 4659 9479 4693 9509
rect 4659 9475 4693 9479
rect 4755 9649 4789 9653
rect 4755 9619 4789 9649
rect 4755 9547 4789 9581
rect 4755 9479 4789 9509
rect 4755 9475 4789 9479
rect 4851 9649 4885 9653
rect 4851 9619 4885 9649
rect 4851 9547 4885 9581
rect 4851 9479 4885 9509
rect 4851 9475 4885 9479
rect 4947 9649 4981 9653
rect 4947 9619 4981 9649
rect 4947 9547 4981 9581
rect 4947 9479 4981 9509
rect 4947 9475 4981 9479
rect 5061 9680 5095 9684
rect 5061 9650 5095 9680
rect 5061 9578 5095 9612
rect 5061 9510 5095 9540
rect 5303 9517 5337 9551
rect 5395 9517 5429 9551
rect 5487 9517 5521 9551
rect 5061 9506 5095 9510
rect 5061 9442 5095 9468
rect 5061 9434 5095 9442
rect 313 9047 347 9081
rect 409 9047 443 9081
rect 505 9047 539 9081
rect 601 9047 635 9081
rect 697 9047 731 9081
rect 793 9047 827 9081
rect 889 9047 923 9081
rect 985 9047 1019 9081
rect 1081 9047 1115 9081
rect 1177 9047 1211 9081
rect 1273 9047 1307 9081
rect 1387 9118 1421 9123
rect 1387 9089 1421 9118
rect 1387 9050 1421 9051
rect 1387 9017 1421 9050
rect 313 8936 347 8970
rect 505 8936 539 8970
rect 697 8936 731 8970
rect 889 8936 923 8970
rect 1081 8936 1115 8970
rect 1273 8936 1307 8970
rect 1387 8948 1421 8979
rect 1387 8945 1421 8948
rect 3691 9162 3725 9196
rect 2466 9051 2500 9085
rect 2562 9051 2596 9085
rect 2658 9051 2692 9085
rect 2754 9051 2788 9085
rect 2850 9051 2884 9085
rect 2946 9051 2980 9085
rect 3042 9051 3076 9085
rect 3138 9051 3172 9085
rect 3234 9051 3268 9085
rect 3330 9051 3364 9085
rect 3426 9051 3460 9085
rect 3540 9122 3574 9127
rect 3540 9093 3574 9122
rect 3540 9054 3574 9055
rect 3540 9021 3574 9054
rect 3647 9036 3681 9112
rect 3735 9036 3769 9112
rect 2466 8940 2500 8974
rect 2658 8940 2692 8974
rect 2850 8940 2884 8974
rect 3042 8940 3076 8974
rect 3234 8940 3268 8974
rect 3426 8940 3460 8974
rect 3540 8952 3574 8983
rect 3540 8949 3574 8952
rect 3987 9051 4021 9085
rect 4083 9051 4117 9085
rect 4179 9051 4213 9085
rect 4275 9051 4309 9085
rect 4371 9051 4405 9085
rect 4467 9051 4501 9085
rect 4563 9051 4597 9085
rect 4659 9051 4693 9085
rect 4755 9051 4789 9085
rect 4851 9051 4885 9085
rect 4947 9051 4981 9085
rect 5061 9122 5095 9127
rect 5061 9093 5095 9122
rect 5061 9054 5095 9055
rect 5061 9021 5095 9054
rect 5348 9203 5382 9237
rect 5450 9239 5484 9242
rect 5450 9208 5470 9239
rect 5470 9208 5484 9239
rect 3987 8940 4021 8974
rect 4179 8940 4213 8974
rect 4371 8940 4405 8974
rect 4563 8940 4597 8974
rect 4755 8940 4789 8974
rect 4947 8940 4981 8974
rect 5061 8952 5095 8983
rect 5303 8973 5337 9007
rect 5395 8973 5429 9007
rect 5487 8973 5521 9007
rect 5061 8949 5095 8952
rect 313 8457 347 8491
rect 505 8457 539 8491
rect 697 8457 731 8491
rect 889 8457 923 8491
rect 1081 8457 1115 8491
rect 1273 8457 1307 8491
rect 1387 8457 1421 8465
rect 1387 8431 1421 8457
rect 313 8358 347 8362
rect 313 8328 347 8358
rect 313 8256 347 8290
rect 313 8188 347 8218
rect 313 8184 347 8188
rect 409 8358 443 8362
rect 409 8328 443 8358
rect 409 8256 443 8290
rect 409 8188 443 8218
rect 409 8184 443 8188
rect 505 8358 539 8362
rect 505 8328 539 8358
rect 505 8256 539 8290
rect 505 8188 539 8218
rect 505 8184 539 8188
rect 601 8358 635 8362
rect 601 8328 635 8358
rect 601 8256 635 8290
rect 601 8188 635 8218
rect 601 8184 635 8188
rect 697 8358 731 8362
rect 697 8328 731 8358
rect 697 8256 731 8290
rect 697 8188 731 8218
rect 697 8184 731 8188
rect 793 8358 827 8362
rect 793 8328 827 8358
rect 793 8256 827 8290
rect 793 8188 827 8218
rect 793 8184 827 8188
rect 889 8358 923 8362
rect 889 8328 923 8358
rect 889 8256 923 8290
rect 889 8188 923 8218
rect 889 8184 923 8188
rect 985 8358 1019 8362
rect 985 8328 1019 8358
rect 985 8256 1019 8290
rect 985 8188 1019 8218
rect 985 8184 1019 8188
rect 1081 8358 1115 8362
rect 1081 8328 1115 8358
rect 1081 8256 1115 8290
rect 1081 8188 1115 8218
rect 1081 8184 1115 8188
rect 1177 8358 1211 8362
rect 1177 8328 1211 8358
rect 1177 8256 1211 8290
rect 1177 8188 1211 8218
rect 1177 8184 1211 8188
rect 1273 8358 1307 8362
rect 1273 8328 1307 8358
rect 1273 8256 1307 8290
rect 1273 8188 1307 8218
rect 1273 8184 1307 8188
rect 1387 8389 1421 8393
rect 1387 8359 1421 8389
rect 1387 8287 1421 8321
rect 1387 8219 1421 8249
rect 1387 8215 1421 8219
rect 1387 8151 1421 8177
rect 1387 8143 1421 8151
rect 2466 8461 2500 8495
rect 2658 8461 2692 8495
rect 2850 8461 2884 8495
rect 3042 8461 3076 8495
rect 3234 8461 3268 8495
rect 3426 8461 3460 8495
rect 3540 8461 3574 8469
rect 3540 8435 3574 8461
rect 2466 8362 2500 8366
rect 2466 8332 2500 8362
rect 2466 8260 2500 8294
rect 2466 8192 2500 8222
rect 2466 8188 2500 8192
rect 2562 8362 2596 8366
rect 2562 8332 2596 8362
rect 2562 8260 2596 8294
rect 2562 8192 2596 8222
rect 2562 8188 2596 8192
rect 2658 8362 2692 8366
rect 2658 8332 2692 8362
rect 2658 8260 2692 8294
rect 2658 8192 2692 8222
rect 2658 8188 2692 8192
rect 2754 8362 2788 8366
rect 2754 8332 2788 8362
rect 2754 8260 2788 8294
rect 2754 8192 2788 8222
rect 2754 8188 2788 8192
rect 2850 8362 2884 8366
rect 2850 8332 2884 8362
rect 2850 8260 2884 8294
rect 2850 8192 2884 8222
rect 2850 8188 2884 8192
rect 2946 8362 2980 8366
rect 2946 8332 2980 8362
rect 2946 8260 2980 8294
rect 2946 8192 2980 8222
rect 2946 8188 2980 8192
rect 3042 8362 3076 8366
rect 3042 8332 3076 8362
rect 3042 8260 3076 8294
rect 3042 8192 3076 8222
rect 3042 8188 3076 8192
rect 3138 8362 3172 8366
rect 3138 8332 3172 8362
rect 3138 8260 3172 8294
rect 3138 8192 3172 8222
rect 3138 8188 3172 8192
rect 3234 8362 3268 8366
rect 3234 8332 3268 8362
rect 3234 8260 3268 8294
rect 3234 8192 3268 8222
rect 3234 8188 3268 8192
rect 3330 8362 3364 8366
rect 3330 8332 3364 8362
rect 3330 8260 3364 8294
rect 3330 8192 3364 8222
rect 3330 8188 3364 8192
rect 3426 8362 3460 8366
rect 3426 8332 3460 8362
rect 3426 8260 3460 8294
rect 3426 8192 3460 8222
rect 3426 8188 3460 8192
rect 3540 8393 3574 8397
rect 3540 8363 3574 8393
rect 3540 8291 3574 8325
rect 3540 8223 3574 8253
rect 3540 8219 3574 8223
rect 3540 8155 3574 8181
rect 3540 8147 3574 8155
rect 3987 8461 4021 8495
rect 4179 8461 4213 8495
rect 4371 8461 4405 8495
rect 4563 8461 4597 8495
rect 4755 8461 4789 8495
rect 4947 8461 4981 8495
rect 5061 8461 5095 8469
rect 5061 8435 5095 8461
rect 3987 8362 4021 8366
rect 3987 8332 4021 8362
rect 3987 8260 4021 8294
rect 3987 8192 4021 8222
rect 3987 8188 4021 8192
rect 4083 8362 4117 8366
rect 4083 8332 4117 8362
rect 4083 8260 4117 8294
rect 4083 8192 4117 8222
rect 4083 8188 4117 8192
rect 4179 8362 4213 8366
rect 4179 8332 4213 8362
rect 4179 8260 4213 8294
rect 4179 8192 4213 8222
rect 4179 8188 4213 8192
rect 4275 8362 4309 8366
rect 4275 8332 4309 8362
rect 4275 8260 4309 8294
rect 4275 8192 4309 8222
rect 4275 8188 4309 8192
rect 4371 8362 4405 8366
rect 4371 8332 4405 8362
rect 4371 8260 4405 8294
rect 4371 8192 4405 8222
rect 4371 8188 4405 8192
rect 4467 8362 4501 8366
rect 4467 8332 4501 8362
rect 4467 8260 4501 8294
rect 4467 8192 4501 8222
rect 4467 8188 4501 8192
rect 4563 8362 4597 8366
rect 4563 8332 4597 8362
rect 4563 8260 4597 8294
rect 4563 8192 4597 8222
rect 4563 8188 4597 8192
rect 4659 8362 4693 8366
rect 4659 8332 4693 8362
rect 4659 8260 4693 8294
rect 4659 8192 4693 8222
rect 4659 8188 4693 8192
rect 4755 8362 4789 8366
rect 4755 8332 4789 8362
rect 4755 8260 4789 8294
rect 4755 8192 4789 8222
rect 4755 8188 4789 8192
rect 4851 8362 4885 8366
rect 4851 8332 4885 8362
rect 4851 8260 4885 8294
rect 4851 8192 4885 8222
rect 4851 8188 4885 8192
rect 4947 8362 4981 8366
rect 4947 8332 4981 8362
rect 4947 8260 4981 8294
rect 4947 8192 4981 8222
rect 4947 8188 4981 8192
rect 5061 8393 5095 8397
rect 5061 8363 5095 8393
rect 5061 8291 5095 8325
rect 5061 8223 5095 8253
rect 5303 8230 5337 8264
rect 5395 8230 5429 8264
rect 5487 8230 5521 8264
rect 5061 8219 5095 8223
rect 5061 8155 5095 8181
rect 5061 8147 5095 8155
rect 313 7760 347 7794
rect 409 7760 443 7794
rect 505 7760 539 7794
rect 601 7760 635 7794
rect 697 7760 731 7794
rect 793 7760 827 7794
rect 889 7760 923 7794
rect 985 7760 1019 7794
rect 1081 7760 1115 7794
rect 1177 7760 1211 7794
rect 1273 7760 1307 7794
rect 1387 7831 1421 7836
rect 1387 7802 1421 7831
rect 1387 7763 1421 7764
rect 1387 7730 1421 7763
rect 313 7649 347 7683
rect 505 7649 539 7683
rect 697 7649 731 7683
rect 889 7649 923 7683
rect 1081 7649 1115 7683
rect 1273 7649 1307 7683
rect 1387 7661 1421 7692
rect 1387 7658 1421 7661
rect 3691 7875 3725 7909
rect 2466 7764 2500 7798
rect 2562 7764 2596 7798
rect 2658 7764 2692 7798
rect 2754 7764 2788 7798
rect 2850 7764 2884 7798
rect 2946 7764 2980 7798
rect 3042 7764 3076 7798
rect 3138 7764 3172 7798
rect 3234 7764 3268 7798
rect 3330 7764 3364 7798
rect 3426 7764 3460 7798
rect 3540 7835 3574 7840
rect 3540 7806 3574 7835
rect 3540 7767 3574 7768
rect 3540 7734 3574 7767
rect 3647 7749 3681 7825
rect 3735 7749 3769 7825
rect 2466 7653 2500 7687
rect 2658 7653 2692 7687
rect 2850 7653 2884 7687
rect 3042 7653 3076 7687
rect 3234 7653 3268 7687
rect 3426 7653 3460 7687
rect 3540 7665 3574 7696
rect 3540 7662 3574 7665
rect 3987 7764 4021 7798
rect 4083 7764 4117 7798
rect 4179 7764 4213 7798
rect 4275 7764 4309 7798
rect 4371 7764 4405 7798
rect 4467 7764 4501 7798
rect 4563 7764 4597 7798
rect 4659 7764 4693 7798
rect 4755 7764 4789 7798
rect 4851 7764 4885 7798
rect 4947 7764 4981 7798
rect 5061 7835 5095 7840
rect 5061 7806 5095 7835
rect 5061 7767 5095 7768
rect 5061 7734 5095 7767
rect 5348 7916 5382 7950
rect 5450 7952 5484 7955
rect 5450 7921 5470 7952
rect 5470 7921 5484 7952
rect 3987 7653 4021 7687
rect 4179 7653 4213 7687
rect 4371 7653 4405 7687
rect 4563 7653 4597 7687
rect 4755 7653 4789 7687
rect 4947 7653 4981 7687
rect 5061 7665 5095 7696
rect 5303 7686 5337 7720
rect 5395 7686 5429 7720
rect 5487 7686 5521 7720
rect 5061 7662 5095 7665
rect 313 7170 347 7204
rect 505 7170 539 7204
rect 697 7170 731 7204
rect 889 7170 923 7204
rect 1081 7170 1115 7204
rect 1273 7170 1307 7204
rect 1387 7170 1421 7178
rect 1387 7144 1421 7170
rect 313 7071 347 7075
rect 313 7041 347 7071
rect 313 6969 347 7003
rect 313 6901 347 6931
rect 313 6897 347 6901
rect 409 7071 443 7075
rect 409 7041 443 7071
rect 409 6969 443 7003
rect 409 6901 443 6931
rect 409 6897 443 6901
rect 505 7071 539 7075
rect 505 7041 539 7071
rect 505 6969 539 7003
rect 505 6901 539 6931
rect 505 6897 539 6901
rect 601 7071 635 7075
rect 601 7041 635 7071
rect 601 6969 635 7003
rect 601 6901 635 6931
rect 601 6897 635 6901
rect 697 7071 731 7075
rect 697 7041 731 7071
rect 697 6969 731 7003
rect 697 6901 731 6931
rect 697 6897 731 6901
rect 793 7071 827 7075
rect 793 7041 827 7071
rect 793 6969 827 7003
rect 793 6901 827 6931
rect 793 6897 827 6901
rect 889 7071 923 7075
rect 889 7041 923 7071
rect 889 6969 923 7003
rect 889 6901 923 6931
rect 889 6897 923 6901
rect 985 7071 1019 7075
rect 985 7041 1019 7071
rect 985 6969 1019 7003
rect 985 6901 1019 6931
rect 985 6897 1019 6901
rect 1081 7071 1115 7075
rect 1081 7041 1115 7071
rect 1081 6969 1115 7003
rect 1081 6901 1115 6931
rect 1081 6897 1115 6901
rect 1177 7071 1211 7075
rect 1177 7041 1211 7071
rect 1177 6969 1211 7003
rect 1177 6901 1211 6931
rect 1177 6897 1211 6901
rect 1273 7071 1307 7075
rect 1273 7041 1307 7071
rect 1273 6969 1307 7003
rect 1273 6901 1307 6931
rect 1273 6897 1307 6901
rect 1387 7102 1421 7106
rect 1387 7072 1421 7102
rect 1387 7000 1421 7034
rect 1387 6932 1421 6962
rect 1387 6928 1421 6932
rect 1387 6864 1421 6890
rect 1387 6856 1421 6864
rect 2466 7174 2500 7208
rect 2658 7174 2692 7208
rect 2850 7174 2884 7208
rect 3042 7174 3076 7208
rect 3234 7174 3268 7208
rect 3426 7174 3460 7208
rect 3540 7174 3574 7182
rect 3540 7148 3574 7174
rect 2466 7075 2500 7079
rect 2466 7045 2500 7075
rect 2466 6973 2500 7007
rect 2466 6905 2500 6935
rect 2466 6901 2500 6905
rect 2562 7075 2596 7079
rect 2562 7045 2596 7075
rect 2562 6973 2596 7007
rect 2562 6905 2596 6935
rect 2562 6901 2596 6905
rect 2658 7075 2692 7079
rect 2658 7045 2692 7075
rect 2658 6973 2692 7007
rect 2658 6905 2692 6935
rect 2658 6901 2692 6905
rect 2754 7075 2788 7079
rect 2754 7045 2788 7075
rect 2754 6973 2788 7007
rect 2754 6905 2788 6935
rect 2754 6901 2788 6905
rect 2850 7075 2884 7079
rect 2850 7045 2884 7075
rect 2850 6973 2884 7007
rect 2850 6905 2884 6935
rect 2850 6901 2884 6905
rect 2946 7075 2980 7079
rect 2946 7045 2980 7075
rect 2946 6973 2980 7007
rect 2946 6905 2980 6935
rect 2946 6901 2980 6905
rect 3042 7075 3076 7079
rect 3042 7045 3076 7075
rect 3042 6973 3076 7007
rect 3042 6905 3076 6935
rect 3042 6901 3076 6905
rect 3138 7075 3172 7079
rect 3138 7045 3172 7075
rect 3138 6973 3172 7007
rect 3138 6905 3172 6935
rect 3138 6901 3172 6905
rect 3234 7075 3268 7079
rect 3234 7045 3268 7075
rect 3234 6973 3268 7007
rect 3234 6905 3268 6935
rect 3234 6901 3268 6905
rect 3330 7075 3364 7079
rect 3330 7045 3364 7075
rect 3330 6973 3364 7007
rect 3330 6905 3364 6935
rect 3330 6901 3364 6905
rect 3426 7075 3460 7079
rect 3426 7045 3460 7075
rect 3426 6973 3460 7007
rect 3426 6905 3460 6935
rect 3426 6901 3460 6905
rect 3540 7106 3574 7110
rect 3540 7076 3574 7106
rect 3540 7004 3574 7038
rect 3540 6936 3574 6966
rect 3540 6932 3574 6936
rect 3540 6868 3574 6894
rect 3540 6860 3574 6868
rect 3987 7174 4021 7208
rect 4179 7174 4213 7208
rect 4371 7174 4405 7208
rect 4563 7174 4597 7208
rect 4755 7174 4789 7208
rect 4947 7174 4981 7208
rect 5061 7174 5095 7182
rect 5061 7148 5095 7174
rect 3987 7075 4021 7079
rect 3987 7045 4021 7075
rect 3987 6973 4021 7007
rect 3987 6905 4021 6935
rect 3987 6901 4021 6905
rect 4083 7075 4117 7079
rect 4083 7045 4117 7075
rect 4083 6973 4117 7007
rect 4083 6905 4117 6935
rect 4083 6901 4117 6905
rect 4179 7075 4213 7079
rect 4179 7045 4213 7075
rect 4179 6973 4213 7007
rect 4179 6905 4213 6935
rect 4179 6901 4213 6905
rect 4275 7075 4309 7079
rect 4275 7045 4309 7075
rect 4275 6973 4309 7007
rect 4275 6905 4309 6935
rect 4275 6901 4309 6905
rect 4371 7075 4405 7079
rect 4371 7045 4405 7075
rect 4371 6973 4405 7007
rect 4371 6905 4405 6935
rect 4371 6901 4405 6905
rect 4467 7075 4501 7079
rect 4467 7045 4501 7075
rect 4467 6973 4501 7007
rect 4467 6905 4501 6935
rect 4467 6901 4501 6905
rect 4563 7075 4597 7079
rect 4563 7045 4597 7075
rect 4563 6973 4597 7007
rect 4563 6905 4597 6935
rect 4563 6901 4597 6905
rect 4659 7075 4693 7079
rect 4659 7045 4693 7075
rect 4659 6973 4693 7007
rect 4659 6905 4693 6935
rect 4659 6901 4693 6905
rect 4755 7075 4789 7079
rect 4755 7045 4789 7075
rect 4755 6973 4789 7007
rect 4755 6905 4789 6935
rect 4755 6901 4789 6905
rect 4851 7075 4885 7079
rect 4851 7045 4885 7075
rect 4851 6973 4885 7007
rect 4851 6905 4885 6935
rect 4851 6901 4885 6905
rect 4947 7075 4981 7079
rect 4947 7045 4981 7075
rect 4947 6973 4981 7007
rect 4947 6905 4981 6935
rect 4947 6901 4981 6905
rect 5061 7106 5095 7110
rect 5061 7076 5095 7106
rect 5061 7004 5095 7038
rect 5061 6936 5095 6966
rect 5303 6943 5337 6977
rect 5395 6943 5429 6977
rect 5487 6943 5521 6977
rect 5061 6932 5095 6936
rect 5061 6868 5095 6894
rect 5061 6860 5095 6868
rect 313 6473 347 6507
rect 409 6473 443 6507
rect 505 6473 539 6507
rect 601 6473 635 6507
rect 697 6473 731 6507
rect 793 6473 827 6507
rect 889 6473 923 6507
rect 985 6473 1019 6507
rect 1081 6473 1115 6507
rect 1177 6473 1211 6507
rect 1273 6473 1307 6507
rect 1387 6544 1421 6549
rect 1387 6515 1421 6544
rect 1387 6476 1421 6477
rect 1387 6443 1421 6476
rect 313 6362 347 6396
rect 505 6362 539 6396
rect 697 6362 731 6396
rect 889 6362 923 6396
rect 1081 6362 1115 6396
rect 1273 6362 1307 6396
rect 1387 6374 1421 6405
rect 1387 6371 1421 6374
rect 3691 6588 3725 6622
rect 2466 6477 2500 6511
rect 2562 6477 2596 6511
rect 2658 6477 2692 6511
rect 2754 6477 2788 6511
rect 2850 6477 2884 6511
rect 2946 6477 2980 6511
rect 3042 6477 3076 6511
rect 3138 6477 3172 6511
rect 3234 6477 3268 6511
rect 3330 6477 3364 6511
rect 3426 6477 3460 6511
rect 3540 6548 3574 6553
rect 3540 6519 3574 6548
rect 3540 6480 3574 6481
rect 3540 6447 3574 6480
rect 3647 6462 3681 6538
rect 3735 6462 3769 6538
rect 2466 6366 2500 6400
rect 2658 6366 2692 6400
rect 2850 6366 2884 6400
rect 3042 6366 3076 6400
rect 3234 6366 3268 6400
rect 3426 6366 3460 6400
rect 3540 6378 3574 6409
rect 3540 6375 3574 6378
rect 3987 6477 4021 6511
rect 4083 6477 4117 6511
rect 4179 6477 4213 6511
rect 4275 6477 4309 6511
rect 4371 6477 4405 6511
rect 4467 6477 4501 6511
rect 4563 6477 4597 6511
rect 4659 6477 4693 6511
rect 4755 6477 4789 6511
rect 4851 6477 4885 6511
rect 4947 6477 4981 6511
rect 5061 6548 5095 6553
rect 5061 6519 5095 6548
rect 5061 6480 5095 6481
rect 5061 6447 5095 6480
rect 5348 6629 5382 6663
rect 5450 6665 5484 6668
rect 5450 6634 5470 6665
rect 5470 6634 5484 6665
rect 3987 6366 4021 6400
rect 4179 6366 4213 6400
rect 4371 6366 4405 6400
rect 4563 6366 4597 6400
rect 4755 6366 4789 6400
rect 4947 6366 4981 6400
rect 5061 6378 5095 6409
rect 5303 6399 5337 6433
rect 5395 6399 5429 6433
rect 5487 6399 5521 6433
rect 5061 6375 5095 6378
rect 313 5883 347 5917
rect 505 5883 539 5917
rect 697 5883 731 5917
rect 889 5883 923 5917
rect 1081 5883 1115 5917
rect 1273 5883 1307 5917
rect 1387 5883 1421 5891
rect 1387 5857 1421 5883
rect 313 5784 347 5788
rect 313 5754 347 5784
rect 313 5682 347 5716
rect 313 5614 347 5644
rect 313 5610 347 5614
rect 409 5784 443 5788
rect 409 5754 443 5784
rect 409 5682 443 5716
rect 409 5614 443 5644
rect 409 5610 443 5614
rect 505 5784 539 5788
rect 505 5754 539 5784
rect 505 5682 539 5716
rect 505 5614 539 5644
rect 505 5610 539 5614
rect 601 5784 635 5788
rect 601 5754 635 5784
rect 601 5682 635 5716
rect 601 5614 635 5644
rect 601 5610 635 5614
rect 697 5784 731 5788
rect 697 5754 731 5784
rect 697 5682 731 5716
rect 697 5614 731 5644
rect 697 5610 731 5614
rect 793 5784 827 5788
rect 793 5754 827 5784
rect 793 5682 827 5716
rect 793 5614 827 5644
rect 793 5610 827 5614
rect 889 5784 923 5788
rect 889 5754 923 5784
rect 889 5682 923 5716
rect 889 5614 923 5644
rect 889 5610 923 5614
rect 985 5784 1019 5788
rect 985 5754 1019 5784
rect 985 5682 1019 5716
rect 985 5614 1019 5644
rect 985 5610 1019 5614
rect 1081 5784 1115 5788
rect 1081 5754 1115 5784
rect 1081 5682 1115 5716
rect 1081 5614 1115 5644
rect 1081 5610 1115 5614
rect 1177 5784 1211 5788
rect 1177 5754 1211 5784
rect 1177 5682 1211 5716
rect 1177 5614 1211 5644
rect 1177 5610 1211 5614
rect 1273 5784 1307 5788
rect 1273 5754 1307 5784
rect 1273 5682 1307 5716
rect 1273 5614 1307 5644
rect 1273 5610 1307 5614
rect 1387 5815 1421 5819
rect 1387 5785 1421 5815
rect 1387 5713 1421 5747
rect 1387 5645 1421 5675
rect 1387 5641 1421 5645
rect 1387 5577 1421 5603
rect 1387 5569 1421 5577
rect 2466 5887 2500 5921
rect 2658 5887 2692 5921
rect 2850 5887 2884 5921
rect 3042 5887 3076 5921
rect 3234 5887 3268 5921
rect 3426 5887 3460 5921
rect 3540 5887 3574 5895
rect 3540 5861 3574 5887
rect 2466 5788 2500 5792
rect 2466 5758 2500 5788
rect 2466 5686 2500 5720
rect 2466 5618 2500 5648
rect 2466 5614 2500 5618
rect 2562 5788 2596 5792
rect 2562 5758 2596 5788
rect 2562 5686 2596 5720
rect 2562 5618 2596 5648
rect 2562 5614 2596 5618
rect 2658 5788 2692 5792
rect 2658 5758 2692 5788
rect 2658 5686 2692 5720
rect 2658 5618 2692 5648
rect 2658 5614 2692 5618
rect 2754 5788 2788 5792
rect 2754 5758 2788 5788
rect 2754 5686 2788 5720
rect 2754 5618 2788 5648
rect 2754 5614 2788 5618
rect 2850 5788 2884 5792
rect 2850 5758 2884 5788
rect 2850 5686 2884 5720
rect 2850 5618 2884 5648
rect 2850 5614 2884 5618
rect 2946 5788 2980 5792
rect 2946 5758 2980 5788
rect 2946 5686 2980 5720
rect 2946 5618 2980 5648
rect 2946 5614 2980 5618
rect 3042 5788 3076 5792
rect 3042 5758 3076 5788
rect 3042 5686 3076 5720
rect 3042 5618 3076 5648
rect 3042 5614 3076 5618
rect 3138 5788 3172 5792
rect 3138 5758 3172 5788
rect 3138 5686 3172 5720
rect 3138 5618 3172 5648
rect 3138 5614 3172 5618
rect 3234 5788 3268 5792
rect 3234 5758 3268 5788
rect 3234 5686 3268 5720
rect 3234 5618 3268 5648
rect 3234 5614 3268 5618
rect 3330 5788 3364 5792
rect 3330 5758 3364 5788
rect 3330 5686 3364 5720
rect 3330 5618 3364 5648
rect 3330 5614 3364 5618
rect 3426 5788 3460 5792
rect 3426 5758 3460 5788
rect 3426 5686 3460 5720
rect 3426 5618 3460 5648
rect 3426 5614 3460 5618
rect 3540 5819 3574 5823
rect 3540 5789 3574 5819
rect 3540 5717 3574 5751
rect 3540 5649 3574 5679
rect 3540 5645 3574 5649
rect 3540 5581 3574 5607
rect 3540 5573 3574 5581
rect 3987 5887 4021 5921
rect 4179 5887 4213 5921
rect 4371 5887 4405 5921
rect 4563 5887 4597 5921
rect 4755 5887 4789 5921
rect 4947 5887 4981 5921
rect 5061 5887 5095 5895
rect 5061 5861 5095 5887
rect 3987 5788 4021 5792
rect 3987 5758 4021 5788
rect 3987 5686 4021 5720
rect 3987 5618 4021 5648
rect 3987 5614 4021 5618
rect 4083 5788 4117 5792
rect 4083 5758 4117 5788
rect 4083 5686 4117 5720
rect 4083 5618 4117 5648
rect 4083 5614 4117 5618
rect 4179 5788 4213 5792
rect 4179 5758 4213 5788
rect 4179 5686 4213 5720
rect 4179 5618 4213 5648
rect 4179 5614 4213 5618
rect 4275 5788 4309 5792
rect 4275 5758 4309 5788
rect 4275 5686 4309 5720
rect 4275 5618 4309 5648
rect 4275 5614 4309 5618
rect 4371 5788 4405 5792
rect 4371 5758 4405 5788
rect 4371 5686 4405 5720
rect 4371 5618 4405 5648
rect 4371 5614 4405 5618
rect 4467 5788 4501 5792
rect 4467 5758 4501 5788
rect 4467 5686 4501 5720
rect 4467 5618 4501 5648
rect 4467 5614 4501 5618
rect 4563 5788 4597 5792
rect 4563 5758 4597 5788
rect 4563 5686 4597 5720
rect 4563 5618 4597 5648
rect 4563 5614 4597 5618
rect 4659 5788 4693 5792
rect 4659 5758 4693 5788
rect 4659 5686 4693 5720
rect 4659 5618 4693 5648
rect 4659 5614 4693 5618
rect 4755 5788 4789 5792
rect 4755 5758 4789 5788
rect 4755 5686 4789 5720
rect 4755 5618 4789 5648
rect 4755 5614 4789 5618
rect 4851 5788 4885 5792
rect 4851 5758 4885 5788
rect 4851 5686 4885 5720
rect 4851 5618 4885 5648
rect 4851 5614 4885 5618
rect 4947 5788 4981 5792
rect 4947 5758 4981 5788
rect 4947 5686 4981 5720
rect 4947 5618 4981 5648
rect 4947 5614 4981 5618
rect 5061 5819 5095 5823
rect 5061 5789 5095 5819
rect 5061 5717 5095 5751
rect 5061 5649 5095 5679
rect 5303 5656 5337 5690
rect 5395 5656 5429 5690
rect 5487 5656 5521 5690
rect 5061 5645 5095 5649
rect 5061 5581 5095 5607
rect 5061 5573 5095 5581
rect 313 5186 347 5220
rect 409 5186 443 5220
rect 505 5186 539 5220
rect 601 5186 635 5220
rect 697 5186 731 5220
rect 793 5186 827 5220
rect 889 5186 923 5220
rect 985 5186 1019 5220
rect 1081 5186 1115 5220
rect 1177 5186 1211 5220
rect 1273 5186 1307 5220
rect 1387 5257 1421 5262
rect 1387 5228 1421 5257
rect 1387 5189 1421 5190
rect 1387 5156 1421 5189
rect 313 5075 347 5109
rect 505 5075 539 5109
rect 697 5075 731 5109
rect 889 5075 923 5109
rect 1081 5075 1115 5109
rect 1273 5075 1307 5109
rect 1387 5087 1421 5118
rect 1387 5084 1421 5087
rect 3691 5301 3725 5335
rect 2466 5190 2500 5224
rect 2562 5190 2596 5224
rect 2658 5190 2692 5224
rect 2754 5190 2788 5224
rect 2850 5190 2884 5224
rect 2946 5190 2980 5224
rect 3042 5190 3076 5224
rect 3138 5190 3172 5224
rect 3234 5190 3268 5224
rect 3330 5190 3364 5224
rect 3426 5190 3460 5224
rect 3540 5261 3574 5266
rect 3540 5232 3574 5261
rect 3540 5193 3574 5194
rect 3540 5160 3574 5193
rect 3647 5175 3681 5251
rect 3735 5175 3769 5251
rect 2466 5079 2500 5113
rect 2658 5079 2692 5113
rect 2850 5079 2884 5113
rect 3042 5079 3076 5113
rect 3234 5079 3268 5113
rect 3426 5079 3460 5113
rect 3540 5091 3574 5122
rect 3540 5088 3574 5091
rect 3987 5190 4021 5224
rect 4083 5190 4117 5224
rect 4179 5190 4213 5224
rect 4275 5190 4309 5224
rect 4371 5190 4405 5224
rect 4467 5190 4501 5224
rect 4563 5190 4597 5224
rect 4659 5190 4693 5224
rect 4755 5190 4789 5224
rect 4851 5190 4885 5224
rect 4947 5190 4981 5224
rect 5061 5261 5095 5266
rect 5061 5232 5095 5261
rect 5061 5193 5095 5194
rect 5061 5160 5095 5193
rect 5348 5342 5382 5376
rect 5450 5378 5484 5381
rect 5450 5347 5470 5378
rect 5470 5347 5484 5378
rect 3987 5079 4021 5113
rect 4179 5079 4213 5113
rect 4371 5079 4405 5113
rect 4563 5079 4597 5113
rect 4755 5079 4789 5113
rect 4947 5079 4981 5113
rect 5061 5091 5095 5122
rect 5303 5112 5337 5146
rect 5395 5112 5429 5146
rect 5487 5112 5521 5146
rect 5061 5088 5095 5091
rect 313 4596 347 4630
rect 505 4596 539 4630
rect 697 4596 731 4630
rect 889 4596 923 4630
rect 1081 4596 1115 4630
rect 1273 4596 1307 4630
rect 1387 4596 1421 4604
rect 1387 4570 1421 4596
rect 313 4497 347 4501
rect 313 4467 347 4497
rect 313 4395 347 4429
rect 313 4327 347 4357
rect 313 4323 347 4327
rect 409 4497 443 4501
rect 409 4467 443 4497
rect 409 4395 443 4429
rect 409 4327 443 4357
rect 409 4323 443 4327
rect 505 4497 539 4501
rect 505 4467 539 4497
rect 505 4395 539 4429
rect 505 4327 539 4357
rect 505 4323 539 4327
rect 601 4497 635 4501
rect 601 4467 635 4497
rect 601 4395 635 4429
rect 601 4327 635 4357
rect 601 4323 635 4327
rect 697 4497 731 4501
rect 697 4467 731 4497
rect 697 4395 731 4429
rect 697 4327 731 4357
rect 697 4323 731 4327
rect 793 4497 827 4501
rect 793 4467 827 4497
rect 793 4395 827 4429
rect 793 4327 827 4357
rect 793 4323 827 4327
rect 889 4497 923 4501
rect 889 4467 923 4497
rect 889 4395 923 4429
rect 889 4327 923 4357
rect 889 4323 923 4327
rect 985 4497 1019 4501
rect 985 4467 1019 4497
rect 985 4395 1019 4429
rect 985 4327 1019 4357
rect 985 4323 1019 4327
rect 1081 4497 1115 4501
rect 1081 4467 1115 4497
rect 1081 4395 1115 4429
rect 1081 4327 1115 4357
rect 1081 4323 1115 4327
rect 1177 4497 1211 4501
rect 1177 4467 1211 4497
rect 1177 4395 1211 4429
rect 1177 4327 1211 4357
rect 1177 4323 1211 4327
rect 1273 4497 1307 4501
rect 1273 4467 1307 4497
rect 1273 4395 1307 4429
rect 1273 4327 1307 4357
rect 1273 4323 1307 4327
rect 1387 4528 1421 4532
rect 1387 4498 1421 4528
rect 1387 4426 1421 4460
rect 1387 4358 1421 4388
rect 1387 4354 1421 4358
rect 1387 4290 1421 4316
rect 1387 4282 1421 4290
rect 2466 4600 2500 4634
rect 2658 4600 2692 4634
rect 2850 4600 2884 4634
rect 3042 4600 3076 4634
rect 3234 4600 3268 4634
rect 3426 4600 3460 4634
rect 3540 4600 3574 4608
rect 3540 4574 3574 4600
rect 2466 4501 2500 4505
rect 2466 4471 2500 4501
rect 2466 4399 2500 4433
rect 2466 4331 2500 4361
rect 2466 4327 2500 4331
rect 2562 4501 2596 4505
rect 2562 4471 2596 4501
rect 2562 4399 2596 4433
rect 2562 4331 2596 4361
rect 2562 4327 2596 4331
rect 2658 4501 2692 4505
rect 2658 4471 2692 4501
rect 2658 4399 2692 4433
rect 2658 4331 2692 4361
rect 2658 4327 2692 4331
rect 2754 4501 2788 4505
rect 2754 4471 2788 4501
rect 2754 4399 2788 4433
rect 2754 4331 2788 4361
rect 2754 4327 2788 4331
rect 2850 4501 2884 4505
rect 2850 4471 2884 4501
rect 2850 4399 2884 4433
rect 2850 4331 2884 4361
rect 2850 4327 2884 4331
rect 2946 4501 2980 4505
rect 2946 4471 2980 4501
rect 2946 4399 2980 4433
rect 2946 4331 2980 4361
rect 2946 4327 2980 4331
rect 3042 4501 3076 4505
rect 3042 4471 3076 4501
rect 3042 4399 3076 4433
rect 3042 4331 3076 4361
rect 3042 4327 3076 4331
rect 3138 4501 3172 4505
rect 3138 4471 3172 4501
rect 3138 4399 3172 4433
rect 3138 4331 3172 4361
rect 3138 4327 3172 4331
rect 3234 4501 3268 4505
rect 3234 4471 3268 4501
rect 3234 4399 3268 4433
rect 3234 4331 3268 4361
rect 3234 4327 3268 4331
rect 3330 4501 3364 4505
rect 3330 4471 3364 4501
rect 3330 4399 3364 4433
rect 3330 4331 3364 4361
rect 3330 4327 3364 4331
rect 3426 4501 3460 4505
rect 3426 4471 3460 4501
rect 3426 4399 3460 4433
rect 3426 4331 3460 4361
rect 3426 4327 3460 4331
rect 3540 4532 3574 4536
rect 3540 4502 3574 4532
rect 3540 4430 3574 4464
rect 3540 4362 3574 4392
rect 3540 4358 3574 4362
rect 3540 4294 3574 4320
rect 3540 4286 3574 4294
rect 3987 4600 4021 4634
rect 4179 4600 4213 4634
rect 4371 4600 4405 4634
rect 4563 4600 4597 4634
rect 4755 4600 4789 4634
rect 4947 4600 4981 4634
rect 5061 4600 5095 4608
rect 5061 4574 5095 4600
rect 3987 4501 4021 4505
rect 3987 4471 4021 4501
rect 3987 4399 4021 4433
rect 3987 4331 4021 4361
rect 3987 4327 4021 4331
rect 4083 4501 4117 4505
rect 4083 4471 4117 4501
rect 4083 4399 4117 4433
rect 4083 4331 4117 4361
rect 4083 4327 4117 4331
rect 4179 4501 4213 4505
rect 4179 4471 4213 4501
rect 4179 4399 4213 4433
rect 4179 4331 4213 4361
rect 4179 4327 4213 4331
rect 4275 4501 4309 4505
rect 4275 4471 4309 4501
rect 4275 4399 4309 4433
rect 4275 4331 4309 4361
rect 4275 4327 4309 4331
rect 4371 4501 4405 4505
rect 4371 4471 4405 4501
rect 4371 4399 4405 4433
rect 4371 4331 4405 4361
rect 4371 4327 4405 4331
rect 4467 4501 4501 4505
rect 4467 4471 4501 4501
rect 4467 4399 4501 4433
rect 4467 4331 4501 4361
rect 4467 4327 4501 4331
rect 4563 4501 4597 4505
rect 4563 4471 4597 4501
rect 4563 4399 4597 4433
rect 4563 4331 4597 4361
rect 4563 4327 4597 4331
rect 4659 4501 4693 4505
rect 4659 4471 4693 4501
rect 4659 4399 4693 4433
rect 4659 4331 4693 4361
rect 4659 4327 4693 4331
rect 4755 4501 4789 4505
rect 4755 4471 4789 4501
rect 4755 4399 4789 4433
rect 4755 4331 4789 4361
rect 4755 4327 4789 4331
rect 4851 4501 4885 4505
rect 4851 4471 4885 4501
rect 4851 4399 4885 4433
rect 4851 4331 4885 4361
rect 4851 4327 4885 4331
rect 4947 4501 4981 4505
rect 4947 4471 4981 4501
rect 4947 4399 4981 4433
rect 4947 4331 4981 4361
rect 4947 4327 4981 4331
rect 5061 4532 5095 4536
rect 5061 4502 5095 4532
rect 5061 4430 5095 4464
rect 5061 4362 5095 4392
rect 5303 4369 5337 4403
rect 5395 4369 5429 4403
rect 5487 4369 5521 4403
rect 5061 4358 5095 4362
rect 5061 4294 5095 4320
rect 5061 4286 5095 4294
rect 313 3899 347 3933
rect 409 3899 443 3933
rect 505 3899 539 3933
rect 601 3899 635 3933
rect 697 3899 731 3933
rect 793 3899 827 3933
rect 889 3899 923 3933
rect 985 3899 1019 3933
rect 1081 3899 1115 3933
rect 1177 3899 1211 3933
rect 1273 3899 1307 3933
rect 1387 3970 1421 3975
rect 1387 3941 1421 3970
rect 1387 3902 1421 3903
rect 1387 3869 1421 3902
rect 313 3788 347 3822
rect 505 3788 539 3822
rect 697 3788 731 3822
rect 889 3788 923 3822
rect 1081 3788 1115 3822
rect 1273 3788 1307 3822
rect 1387 3800 1421 3831
rect 1387 3797 1421 3800
rect 3691 4014 3725 4048
rect 2466 3903 2500 3937
rect 2562 3903 2596 3937
rect 2658 3903 2692 3937
rect 2754 3903 2788 3937
rect 2850 3903 2884 3937
rect 2946 3903 2980 3937
rect 3042 3903 3076 3937
rect 3138 3903 3172 3937
rect 3234 3903 3268 3937
rect 3330 3903 3364 3937
rect 3426 3903 3460 3937
rect 3540 3974 3574 3979
rect 3540 3945 3574 3974
rect 3540 3906 3574 3907
rect 3540 3873 3574 3906
rect 3647 3888 3681 3964
rect 3735 3888 3769 3964
rect 2466 3792 2500 3826
rect 2658 3792 2692 3826
rect 2850 3792 2884 3826
rect 3042 3792 3076 3826
rect 3234 3792 3268 3826
rect 3426 3792 3460 3826
rect 3540 3804 3574 3835
rect 3540 3801 3574 3804
rect 3987 3903 4021 3937
rect 4083 3903 4117 3937
rect 4179 3903 4213 3937
rect 4275 3903 4309 3937
rect 4371 3903 4405 3937
rect 4467 3903 4501 3937
rect 4563 3903 4597 3937
rect 4659 3903 4693 3937
rect 4755 3903 4789 3937
rect 4851 3903 4885 3937
rect 4947 3903 4981 3937
rect 5061 3974 5095 3979
rect 5061 3945 5095 3974
rect 5061 3906 5095 3907
rect 5061 3873 5095 3906
rect 5348 4055 5382 4089
rect 5450 4091 5484 4094
rect 5450 4060 5470 4091
rect 5470 4060 5484 4091
rect 3987 3792 4021 3826
rect 4179 3792 4213 3826
rect 4371 3792 4405 3826
rect 4563 3792 4597 3826
rect 4755 3792 4789 3826
rect 4947 3792 4981 3826
rect 5061 3804 5095 3835
rect 5303 3825 5337 3859
rect 5395 3825 5429 3859
rect 5487 3825 5521 3859
rect 5061 3801 5095 3804
rect 313 3309 347 3343
rect 505 3309 539 3343
rect 697 3309 731 3343
rect 889 3309 923 3343
rect 1081 3309 1115 3343
rect 1273 3309 1307 3343
rect 1387 3309 1421 3317
rect 1387 3283 1421 3309
rect 313 3210 347 3214
rect 313 3180 347 3210
rect 313 3108 347 3142
rect 313 3040 347 3070
rect 313 3036 347 3040
rect 409 3210 443 3214
rect 409 3180 443 3210
rect 409 3108 443 3142
rect 409 3040 443 3070
rect 409 3036 443 3040
rect 505 3210 539 3214
rect 505 3180 539 3210
rect 505 3108 539 3142
rect 505 3040 539 3070
rect 505 3036 539 3040
rect 601 3210 635 3214
rect 601 3180 635 3210
rect 601 3108 635 3142
rect 601 3040 635 3070
rect 601 3036 635 3040
rect 697 3210 731 3214
rect 697 3180 731 3210
rect 697 3108 731 3142
rect 697 3040 731 3070
rect 697 3036 731 3040
rect 793 3210 827 3214
rect 793 3180 827 3210
rect 793 3108 827 3142
rect 793 3040 827 3070
rect 793 3036 827 3040
rect 889 3210 923 3214
rect 889 3180 923 3210
rect 889 3108 923 3142
rect 889 3040 923 3070
rect 889 3036 923 3040
rect 985 3210 1019 3214
rect 985 3180 1019 3210
rect 985 3108 1019 3142
rect 985 3040 1019 3070
rect 985 3036 1019 3040
rect 1081 3210 1115 3214
rect 1081 3180 1115 3210
rect 1081 3108 1115 3142
rect 1081 3040 1115 3070
rect 1081 3036 1115 3040
rect 1177 3210 1211 3214
rect 1177 3180 1211 3210
rect 1177 3108 1211 3142
rect 1177 3040 1211 3070
rect 1177 3036 1211 3040
rect 1273 3210 1307 3214
rect 1273 3180 1307 3210
rect 1273 3108 1307 3142
rect 1273 3040 1307 3070
rect 1273 3036 1307 3040
rect 1387 3241 1421 3245
rect 1387 3211 1421 3241
rect 1387 3139 1421 3173
rect 1387 3071 1421 3101
rect 1387 3067 1421 3071
rect 1387 3003 1421 3029
rect 1387 2995 1421 3003
rect 2466 3313 2500 3347
rect 2658 3313 2692 3347
rect 2850 3313 2884 3347
rect 3042 3313 3076 3347
rect 3234 3313 3268 3347
rect 3426 3313 3460 3347
rect 3540 3313 3574 3321
rect 3540 3287 3574 3313
rect 2466 3214 2500 3218
rect 2466 3184 2500 3214
rect 2466 3112 2500 3146
rect 2466 3044 2500 3074
rect 2466 3040 2500 3044
rect 2562 3214 2596 3218
rect 2562 3184 2596 3214
rect 2562 3112 2596 3146
rect 2562 3044 2596 3074
rect 2562 3040 2596 3044
rect 2658 3214 2692 3218
rect 2658 3184 2692 3214
rect 2658 3112 2692 3146
rect 2658 3044 2692 3074
rect 2658 3040 2692 3044
rect 2754 3214 2788 3218
rect 2754 3184 2788 3214
rect 2754 3112 2788 3146
rect 2754 3044 2788 3074
rect 2754 3040 2788 3044
rect 2850 3214 2884 3218
rect 2850 3184 2884 3214
rect 2850 3112 2884 3146
rect 2850 3044 2884 3074
rect 2850 3040 2884 3044
rect 2946 3214 2980 3218
rect 2946 3184 2980 3214
rect 2946 3112 2980 3146
rect 2946 3044 2980 3074
rect 2946 3040 2980 3044
rect 3042 3214 3076 3218
rect 3042 3184 3076 3214
rect 3042 3112 3076 3146
rect 3042 3044 3076 3074
rect 3042 3040 3076 3044
rect 3138 3214 3172 3218
rect 3138 3184 3172 3214
rect 3138 3112 3172 3146
rect 3138 3044 3172 3074
rect 3138 3040 3172 3044
rect 3234 3214 3268 3218
rect 3234 3184 3268 3214
rect 3234 3112 3268 3146
rect 3234 3044 3268 3074
rect 3234 3040 3268 3044
rect 3330 3214 3364 3218
rect 3330 3184 3364 3214
rect 3330 3112 3364 3146
rect 3330 3044 3364 3074
rect 3330 3040 3364 3044
rect 3426 3214 3460 3218
rect 3426 3184 3460 3214
rect 3426 3112 3460 3146
rect 3426 3044 3460 3074
rect 3426 3040 3460 3044
rect 3540 3245 3574 3249
rect 3540 3215 3574 3245
rect 3540 3143 3574 3177
rect 3540 3075 3574 3105
rect 3540 3071 3574 3075
rect 3540 3007 3574 3033
rect 3540 2999 3574 3007
rect 3987 3313 4021 3347
rect 4179 3313 4213 3347
rect 4371 3313 4405 3347
rect 4563 3313 4597 3347
rect 4755 3313 4789 3347
rect 4947 3313 4981 3347
rect 5061 3313 5095 3321
rect 5061 3287 5095 3313
rect 3987 3214 4021 3218
rect 3987 3184 4021 3214
rect 3987 3112 4021 3146
rect 3987 3044 4021 3074
rect 3987 3040 4021 3044
rect 4083 3214 4117 3218
rect 4083 3184 4117 3214
rect 4083 3112 4117 3146
rect 4083 3044 4117 3074
rect 4083 3040 4117 3044
rect 4179 3214 4213 3218
rect 4179 3184 4213 3214
rect 4179 3112 4213 3146
rect 4179 3044 4213 3074
rect 4179 3040 4213 3044
rect 4275 3214 4309 3218
rect 4275 3184 4309 3214
rect 4275 3112 4309 3146
rect 4275 3044 4309 3074
rect 4275 3040 4309 3044
rect 4371 3214 4405 3218
rect 4371 3184 4405 3214
rect 4371 3112 4405 3146
rect 4371 3044 4405 3074
rect 4371 3040 4405 3044
rect 4467 3214 4501 3218
rect 4467 3184 4501 3214
rect 4467 3112 4501 3146
rect 4467 3044 4501 3074
rect 4467 3040 4501 3044
rect 4563 3214 4597 3218
rect 4563 3184 4597 3214
rect 4563 3112 4597 3146
rect 4563 3044 4597 3074
rect 4563 3040 4597 3044
rect 4659 3214 4693 3218
rect 4659 3184 4693 3214
rect 4659 3112 4693 3146
rect 4659 3044 4693 3074
rect 4659 3040 4693 3044
rect 4755 3214 4789 3218
rect 4755 3184 4789 3214
rect 4755 3112 4789 3146
rect 4755 3044 4789 3074
rect 4755 3040 4789 3044
rect 4851 3214 4885 3218
rect 4851 3184 4885 3214
rect 4851 3112 4885 3146
rect 4851 3044 4885 3074
rect 4851 3040 4885 3044
rect 4947 3214 4981 3218
rect 4947 3184 4981 3214
rect 4947 3112 4981 3146
rect 4947 3044 4981 3074
rect 4947 3040 4981 3044
rect 5061 3245 5095 3249
rect 5061 3215 5095 3245
rect 5061 3143 5095 3177
rect 5061 3075 5095 3105
rect 5303 3082 5337 3116
rect 5395 3082 5429 3116
rect 5487 3082 5521 3116
rect 5061 3071 5095 3075
rect 5061 3007 5095 3033
rect 5061 2999 5095 3007
rect 313 2612 347 2646
rect 409 2612 443 2646
rect 505 2612 539 2646
rect 601 2612 635 2646
rect 697 2612 731 2646
rect 793 2612 827 2646
rect 889 2612 923 2646
rect 985 2612 1019 2646
rect 1081 2612 1115 2646
rect 1177 2612 1211 2646
rect 1273 2612 1307 2646
rect 1387 2683 1421 2688
rect 1387 2654 1421 2683
rect 1387 2615 1421 2616
rect 1387 2582 1421 2615
rect 313 2501 347 2535
rect 505 2501 539 2535
rect 697 2501 731 2535
rect 889 2501 923 2535
rect 1081 2501 1115 2535
rect 1273 2501 1307 2535
rect 1387 2513 1421 2544
rect 1387 2510 1421 2513
rect 3691 2727 3725 2761
rect 2466 2616 2500 2650
rect 2562 2616 2596 2650
rect 2658 2616 2692 2650
rect 2754 2616 2788 2650
rect 2850 2616 2884 2650
rect 2946 2616 2980 2650
rect 3042 2616 3076 2650
rect 3138 2616 3172 2650
rect 3234 2616 3268 2650
rect 3330 2616 3364 2650
rect 3426 2616 3460 2650
rect 3540 2687 3574 2692
rect 3540 2658 3574 2687
rect 3540 2619 3574 2620
rect 3540 2586 3574 2619
rect 3647 2601 3681 2677
rect 3735 2601 3769 2677
rect 2466 2505 2500 2539
rect 2658 2505 2692 2539
rect 2850 2505 2884 2539
rect 3042 2505 3076 2539
rect 3234 2505 3268 2539
rect 3426 2505 3460 2539
rect 3540 2517 3574 2548
rect 3540 2514 3574 2517
rect 3987 2616 4021 2650
rect 4083 2616 4117 2650
rect 4179 2616 4213 2650
rect 4275 2616 4309 2650
rect 4371 2616 4405 2650
rect 4467 2616 4501 2650
rect 4563 2616 4597 2650
rect 4659 2616 4693 2650
rect 4755 2616 4789 2650
rect 4851 2616 4885 2650
rect 4947 2616 4981 2650
rect 5061 2687 5095 2692
rect 5061 2658 5095 2687
rect 5061 2619 5095 2620
rect 5061 2586 5095 2619
rect 5348 2768 5382 2802
rect 5450 2804 5484 2807
rect 5450 2773 5470 2804
rect 5470 2773 5484 2804
rect 3987 2505 4021 2539
rect 4179 2505 4213 2539
rect 4371 2505 4405 2539
rect 4563 2505 4597 2539
rect 4755 2505 4789 2539
rect 4947 2505 4981 2539
rect 5061 2517 5095 2548
rect 5303 2538 5337 2572
rect 5395 2538 5429 2572
rect 5487 2538 5521 2572
rect 5061 2514 5095 2517
rect 313 2022 347 2056
rect 505 2022 539 2056
rect 697 2022 731 2056
rect 889 2022 923 2056
rect 1081 2022 1115 2056
rect 1273 2022 1307 2056
rect 1387 2022 1421 2030
rect 1387 1996 1421 2022
rect 313 1923 347 1927
rect 313 1893 347 1923
rect 313 1821 347 1855
rect 313 1753 347 1783
rect 313 1749 347 1753
rect 409 1923 443 1927
rect 409 1893 443 1923
rect 409 1821 443 1855
rect 409 1753 443 1783
rect 409 1749 443 1753
rect 505 1923 539 1927
rect 505 1893 539 1923
rect 505 1821 539 1855
rect 505 1753 539 1783
rect 505 1749 539 1753
rect 601 1923 635 1927
rect 601 1893 635 1923
rect 601 1821 635 1855
rect 601 1753 635 1783
rect 601 1749 635 1753
rect 697 1923 731 1927
rect 697 1893 731 1923
rect 697 1821 731 1855
rect 697 1753 731 1783
rect 697 1749 731 1753
rect 793 1923 827 1927
rect 793 1893 827 1923
rect 793 1821 827 1855
rect 793 1753 827 1783
rect 793 1749 827 1753
rect 889 1923 923 1927
rect 889 1893 923 1923
rect 889 1821 923 1855
rect 889 1753 923 1783
rect 889 1749 923 1753
rect 985 1923 1019 1927
rect 985 1893 1019 1923
rect 985 1821 1019 1855
rect 985 1753 1019 1783
rect 985 1749 1019 1753
rect 1081 1923 1115 1927
rect 1081 1893 1115 1923
rect 1081 1821 1115 1855
rect 1081 1753 1115 1783
rect 1081 1749 1115 1753
rect 1177 1923 1211 1927
rect 1177 1893 1211 1923
rect 1177 1821 1211 1855
rect 1177 1753 1211 1783
rect 1177 1749 1211 1753
rect 1273 1923 1307 1927
rect 1273 1893 1307 1923
rect 1273 1821 1307 1855
rect 1273 1753 1307 1783
rect 1273 1749 1307 1753
rect 1387 1954 1421 1958
rect 1387 1924 1421 1954
rect 1387 1852 1421 1886
rect 1387 1784 1421 1814
rect 1387 1780 1421 1784
rect 1387 1716 1421 1742
rect 1387 1708 1421 1716
rect 2466 2026 2500 2060
rect 2658 2026 2692 2060
rect 2850 2026 2884 2060
rect 3042 2026 3076 2060
rect 3234 2026 3268 2060
rect 3426 2026 3460 2060
rect 3540 2026 3574 2034
rect 3540 2000 3574 2026
rect 2466 1927 2500 1931
rect 2466 1897 2500 1927
rect 2466 1825 2500 1859
rect 2466 1757 2500 1787
rect 2466 1753 2500 1757
rect 2562 1927 2596 1931
rect 2562 1897 2596 1927
rect 2562 1825 2596 1859
rect 2562 1757 2596 1787
rect 2562 1753 2596 1757
rect 2658 1927 2692 1931
rect 2658 1897 2692 1927
rect 2658 1825 2692 1859
rect 2658 1757 2692 1787
rect 2658 1753 2692 1757
rect 2754 1927 2788 1931
rect 2754 1897 2788 1927
rect 2754 1825 2788 1859
rect 2754 1757 2788 1787
rect 2754 1753 2788 1757
rect 2850 1927 2884 1931
rect 2850 1897 2884 1927
rect 2850 1825 2884 1859
rect 2850 1757 2884 1787
rect 2850 1753 2884 1757
rect 2946 1927 2980 1931
rect 2946 1897 2980 1927
rect 2946 1825 2980 1859
rect 2946 1757 2980 1787
rect 2946 1753 2980 1757
rect 3042 1927 3076 1931
rect 3042 1897 3076 1927
rect 3042 1825 3076 1859
rect 3042 1757 3076 1787
rect 3042 1753 3076 1757
rect 3138 1927 3172 1931
rect 3138 1897 3172 1927
rect 3138 1825 3172 1859
rect 3138 1757 3172 1787
rect 3138 1753 3172 1757
rect 3234 1927 3268 1931
rect 3234 1897 3268 1927
rect 3234 1825 3268 1859
rect 3234 1757 3268 1787
rect 3234 1753 3268 1757
rect 3330 1927 3364 1931
rect 3330 1897 3364 1927
rect 3330 1825 3364 1859
rect 3330 1757 3364 1787
rect 3330 1753 3364 1757
rect 3426 1927 3460 1931
rect 3426 1897 3460 1927
rect 3426 1825 3460 1859
rect 3426 1757 3460 1787
rect 3426 1753 3460 1757
rect 3540 1958 3574 1962
rect 3540 1928 3574 1958
rect 3540 1856 3574 1890
rect 3540 1788 3574 1818
rect 3540 1784 3574 1788
rect 3540 1720 3574 1746
rect 3540 1712 3574 1720
rect 3987 2026 4021 2060
rect 4179 2026 4213 2060
rect 4371 2026 4405 2060
rect 4563 2026 4597 2060
rect 4755 2026 4789 2060
rect 4947 2026 4981 2060
rect 5061 2026 5095 2034
rect 5061 2000 5095 2026
rect 3987 1927 4021 1931
rect 3987 1897 4021 1927
rect 3987 1825 4021 1859
rect 3987 1757 4021 1787
rect 3987 1753 4021 1757
rect 4083 1927 4117 1931
rect 4083 1897 4117 1927
rect 4083 1825 4117 1859
rect 4083 1757 4117 1787
rect 4083 1753 4117 1757
rect 4179 1927 4213 1931
rect 4179 1897 4213 1927
rect 4179 1825 4213 1859
rect 4179 1757 4213 1787
rect 4179 1753 4213 1757
rect 4275 1927 4309 1931
rect 4275 1897 4309 1927
rect 4275 1825 4309 1859
rect 4275 1757 4309 1787
rect 4275 1753 4309 1757
rect 4371 1927 4405 1931
rect 4371 1897 4405 1927
rect 4371 1825 4405 1859
rect 4371 1757 4405 1787
rect 4371 1753 4405 1757
rect 4467 1927 4501 1931
rect 4467 1897 4501 1927
rect 4467 1825 4501 1859
rect 4467 1757 4501 1787
rect 4467 1753 4501 1757
rect 4563 1927 4597 1931
rect 4563 1897 4597 1927
rect 4563 1825 4597 1859
rect 4563 1757 4597 1787
rect 4563 1753 4597 1757
rect 4659 1927 4693 1931
rect 4659 1897 4693 1927
rect 4659 1825 4693 1859
rect 4659 1757 4693 1787
rect 4659 1753 4693 1757
rect 4755 1927 4789 1931
rect 4755 1897 4789 1927
rect 4755 1825 4789 1859
rect 4755 1757 4789 1787
rect 4755 1753 4789 1757
rect 4851 1927 4885 1931
rect 4851 1897 4885 1927
rect 4851 1825 4885 1859
rect 4851 1757 4885 1787
rect 4851 1753 4885 1757
rect 4947 1927 4981 1931
rect 4947 1897 4981 1927
rect 4947 1825 4981 1859
rect 4947 1757 4981 1787
rect 4947 1753 4981 1757
rect 5061 1958 5095 1962
rect 5061 1928 5095 1958
rect 5061 1856 5095 1890
rect 5061 1788 5095 1818
rect 5303 1795 5337 1829
rect 5395 1795 5429 1829
rect 5487 1795 5521 1829
rect 5061 1784 5095 1788
rect 5061 1720 5095 1746
rect 5061 1712 5095 1720
rect 313 1325 347 1359
rect 409 1325 443 1359
rect 505 1325 539 1359
rect 601 1325 635 1359
rect 697 1325 731 1359
rect 793 1325 827 1359
rect 889 1325 923 1359
rect 985 1325 1019 1359
rect 1081 1325 1115 1359
rect 1177 1325 1211 1359
rect 1273 1325 1307 1359
rect 1387 1396 1421 1401
rect 1387 1367 1421 1396
rect 1387 1328 1421 1329
rect 1387 1295 1421 1328
rect 313 1214 347 1248
rect 505 1214 539 1248
rect 697 1214 731 1248
rect 889 1214 923 1248
rect 1081 1214 1115 1248
rect 1273 1214 1307 1248
rect 1387 1226 1421 1257
rect 1387 1223 1421 1226
rect 3691 1440 3725 1474
rect 2466 1329 2500 1363
rect 2562 1329 2596 1363
rect 2658 1329 2692 1363
rect 2754 1329 2788 1363
rect 2850 1329 2884 1363
rect 2946 1329 2980 1363
rect 3042 1329 3076 1363
rect 3138 1329 3172 1363
rect 3234 1329 3268 1363
rect 3330 1329 3364 1363
rect 3426 1329 3460 1363
rect 3540 1400 3574 1405
rect 3540 1371 3574 1400
rect 3540 1332 3574 1333
rect 3540 1299 3574 1332
rect 3647 1314 3681 1390
rect 3735 1314 3769 1390
rect 2466 1218 2500 1252
rect 2658 1218 2692 1252
rect 2850 1218 2884 1252
rect 3042 1218 3076 1252
rect 3234 1218 3268 1252
rect 3426 1218 3460 1252
rect 3540 1230 3574 1261
rect 3540 1227 3574 1230
rect 3987 1329 4021 1363
rect 4083 1329 4117 1363
rect 4179 1329 4213 1363
rect 4275 1329 4309 1363
rect 4371 1329 4405 1363
rect 4467 1329 4501 1363
rect 4563 1329 4597 1363
rect 4659 1329 4693 1363
rect 4755 1329 4789 1363
rect 4851 1329 4885 1363
rect 4947 1329 4981 1363
rect 5061 1400 5095 1405
rect 5061 1371 5095 1400
rect 5061 1332 5095 1333
rect 5061 1299 5095 1332
rect 5348 1481 5382 1515
rect 5450 1517 5484 1520
rect 5450 1486 5470 1517
rect 5470 1486 5484 1517
rect 3987 1218 4021 1252
rect 4179 1218 4213 1252
rect 4371 1218 4405 1252
rect 4563 1218 4597 1252
rect 4755 1218 4789 1252
rect 4947 1218 4981 1252
rect 5061 1230 5095 1261
rect 5303 1251 5337 1285
rect 5395 1251 5429 1285
rect 5487 1251 5521 1285
rect 5061 1227 5095 1230
<< metal1 >>
rect 129 42021 1211 42055
rect 129 41458 163 42021
rect 294 41911 304 41963
rect 356 41911 366 41963
rect 409 41871 443 42021
rect 487 41911 497 41963
rect 549 41911 559 41963
rect 601 41871 635 42021
rect 678 41911 688 41963
rect 740 41911 750 41963
rect 793 41871 827 42021
rect 870 41911 880 41963
rect 932 41911 942 41963
rect 985 41871 1019 42021
rect 1062 41911 1072 41963
rect 1124 41911 1134 41963
rect 1177 41871 1211 42021
rect 1254 41911 1264 41963
rect 1316 41911 1326 41963
rect 1381 41927 1427 42091
rect 2282 42025 3364 42059
rect 1381 41893 1387 41927
rect 1421 41893 1427 41927
rect 1512 41904 1522 41964
rect 1578 41904 1792 41964
rect 1852 41904 1862 41964
rect 307 41824 353 41871
rect 307 41790 313 41824
rect 347 41790 353 41824
rect 307 41752 353 41790
rect 307 41718 313 41752
rect 347 41718 353 41752
rect 307 41680 353 41718
rect 307 41646 313 41680
rect 347 41646 353 41680
rect 307 41599 353 41646
rect 403 41824 449 41871
rect 403 41790 409 41824
rect 443 41790 449 41824
rect 403 41752 449 41790
rect 403 41718 409 41752
rect 443 41718 449 41752
rect 403 41680 449 41718
rect 403 41646 409 41680
rect 443 41646 449 41680
rect 403 41599 449 41646
rect 499 41824 545 41871
rect 499 41790 505 41824
rect 539 41790 545 41824
rect 499 41752 545 41790
rect 499 41718 505 41752
rect 539 41718 545 41752
rect 499 41680 545 41718
rect 499 41646 505 41680
rect 539 41646 545 41680
rect 499 41599 545 41646
rect 595 41824 641 41871
rect 595 41790 601 41824
rect 635 41790 641 41824
rect 595 41752 641 41790
rect 595 41718 601 41752
rect 635 41718 641 41752
rect 595 41680 641 41718
rect 595 41646 601 41680
rect 635 41646 641 41680
rect 595 41599 641 41646
rect 691 41824 737 41871
rect 691 41790 697 41824
rect 731 41790 737 41824
rect 691 41752 737 41790
rect 691 41718 697 41752
rect 731 41718 737 41752
rect 691 41680 737 41718
rect 691 41646 697 41680
rect 731 41646 737 41680
rect 691 41599 737 41646
rect 787 41824 833 41871
rect 787 41790 793 41824
rect 827 41790 833 41824
rect 787 41752 833 41790
rect 787 41718 793 41752
rect 827 41718 833 41752
rect 787 41680 833 41718
rect 787 41646 793 41680
rect 827 41646 833 41680
rect 787 41599 833 41646
rect 883 41824 929 41871
rect 883 41790 889 41824
rect 923 41790 929 41824
rect 883 41752 929 41790
rect 883 41718 889 41752
rect 923 41718 929 41752
rect 883 41680 929 41718
rect 883 41646 889 41680
rect 923 41646 929 41680
rect 883 41599 929 41646
rect 979 41824 1025 41871
rect 979 41790 985 41824
rect 1019 41790 1025 41824
rect 979 41752 1025 41790
rect 979 41718 985 41752
rect 1019 41718 1025 41752
rect 979 41680 1025 41718
rect 979 41646 985 41680
rect 1019 41646 1025 41680
rect 979 41599 1025 41646
rect 1075 41824 1121 41871
rect 1075 41790 1081 41824
rect 1115 41790 1121 41824
rect 1075 41752 1121 41790
rect 1075 41718 1081 41752
rect 1115 41718 1121 41752
rect 1075 41680 1121 41718
rect 1075 41646 1081 41680
rect 1115 41646 1121 41680
rect 1075 41599 1121 41646
rect 1171 41824 1217 41871
rect 1171 41790 1177 41824
rect 1211 41790 1217 41824
rect 1171 41752 1217 41790
rect 1171 41718 1177 41752
rect 1211 41718 1217 41752
rect 1171 41680 1217 41718
rect 1171 41646 1177 41680
rect 1211 41646 1217 41680
rect 1171 41599 1217 41646
rect 1267 41824 1313 41871
rect 1267 41790 1273 41824
rect 1307 41790 1313 41824
rect 1267 41752 1313 41790
rect 1267 41718 1273 41752
rect 1307 41718 1313 41752
rect 1267 41680 1313 41718
rect 1267 41646 1273 41680
rect 1307 41646 1313 41680
rect 1267 41599 1313 41646
rect 1381 41855 1427 41893
rect 1381 41821 1387 41855
rect 1421 41821 1427 41855
rect 1381 41783 1427 41821
rect 1381 41749 1387 41783
rect 1421 41749 1427 41783
rect 1381 41711 1427 41749
rect 1381 41677 1387 41711
rect 1421 41677 1427 41711
rect 1381 41667 1427 41677
rect 1381 41665 2160 41667
rect 1381 41639 2056 41665
rect 1381 41614 1387 41639
rect 1380 41605 1387 41614
rect 1421 41605 2056 41639
rect 0 41424 163 41458
rect 129 41047 163 41424
rect 313 41458 347 41599
rect 505 41458 539 41599
rect 697 41458 731 41599
rect 889 41458 923 41599
rect 1081 41458 1115 41599
rect 1273 41458 1307 41599
rect 1380 41557 2056 41605
rect 2190 41557 2200 41665
rect 1380 41555 2160 41557
rect 2282 41462 2316 42025
rect 2447 41915 2457 41967
rect 2509 41915 2519 41967
rect 2562 41875 2596 42025
rect 2640 41915 2650 41967
rect 2702 41915 2712 41967
rect 2754 41875 2788 42025
rect 2831 41915 2841 41967
rect 2893 41915 2903 41967
rect 2946 41875 2980 42025
rect 3023 41915 3033 41967
rect 3085 41915 3095 41967
rect 3138 41875 3172 42025
rect 3215 41915 3225 41967
rect 3277 41915 3287 41967
rect 3330 41875 3364 42025
rect 3407 41915 3417 41967
rect 3469 41915 3479 41967
rect 3534 41931 3580 42139
rect 3534 41897 3540 41931
rect 3574 41897 3580 41931
rect 2460 41828 2506 41875
rect 2460 41794 2466 41828
rect 2500 41794 2506 41828
rect 2460 41756 2506 41794
rect 2460 41722 2466 41756
rect 2500 41722 2506 41756
rect 2460 41684 2506 41722
rect 2460 41650 2466 41684
rect 2500 41650 2506 41684
rect 2460 41603 2506 41650
rect 2556 41828 2602 41875
rect 2556 41794 2562 41828
rect 2596 41794 2602 41828
rect 2556 41756 2602 41794
rect 2556 41722 2562 41756
rect 2596 41722 2602 41756
rect 2556 41684 2602 41722
rect 2556 41650 2562 41684
rect 2596 41650 2602 41684
rect 2556 41603 2602 41650
rect 2652 41828 2698 41875
rect 2652 41794 2658 41828
rect 2692 41794 2698 41828
rect 2652 41756 2698 41794
rect 2652 41722 2658 41756
rect 2692 41722 2698 41756
rect 2652 41684 2698 41722
rect 2652 41650 2658 41684
rect 2692 41650 2698 41684
rect 2652 41603 2698 41650
rect 2748 41828 2794 41875
rect 2748 41794 2754 41828
rect 2788 41794 2794 41828
rect 2748 41756 2794 41794
rect 2748 41722 2754 41756
rect 2788 41722 2794 41756
rect 2748 41684 2794 41722
rect 2748 41650 2754 41684
rect 2788 41650 2794 41684
rect 2748 41603 2794 41650
rect 2844 41828 2890 41875
rect 2844 41794 2850 41828
rect 2884 41794 2890 41828
rect 2844 41756 2890 41794
rect 2844 41722 2850 41756
rect 2884 41722 2890 41756
rect 2844 41684 2890 41722
rect 2844 41650 2850 41684
rect 2884 41650 2890 41684
rect 2844 41603 2890 41650
rect 2940 41828 2986 41875
rect 2940 41794 2946 41828
rect 2980 41794 2986 41828
rect 2940 41756 2986 41794
rect 2940 41722 2946 41756
rect 2980 41722 2986 41756
rect 2940 41684 2986 41722
rect 2940 41650 2946 41684
rect 2980 41650 2986 41684
rect 2940 41603 2986 41650
rect 3036 41828 3082 41875
rect 3036 41794 3042 41828
rect 3076 41794 3082 41828
rect 3036 41756 3082 41794
rect 3036 41722 3042 41756
rect 3076 41722 3082 41756
rect 3036 41684 3082 41722
rect 3036 41650 3042 41684
rect 3076 41650 3082 41684
rect 3036 41603 3082 41650
rect 3132 41828 3178 41875
rect 3132 41794 3138 41828
rect 3172 41794 3178 41828
rect 3132 41756 3178 41794
rect 3132 41722 3138 41756
rect 3172 41722 3178 41756
rect 3132 41684 3178 41722
rect 3132 41650 3138 41684
rect 3172 41650 3178 41684
rect 3132 41603 3178 41650
rect 3228 41828 3274 41875
rect 3228 41794 3234 41828
rect 3268 41794 3274 41828
rect 3228 41756 3274 41794
rect 3228 41722 3234 41756
rect 3268 41722 3274 41756
rect 3228 41684 3274 41722
rect 3228 41650 3234 41684
rect 3268 41650 3274 41684
rect 3228 41603 3274 41650
rect 3324 41828 3370 41875
rect 3324 41794 3330 41828
rect 3364 41794 3370 41828
rect 3324 41756 3370 41794
rect 3324 41722 3330 41756
rect 3364 41722 3370 41756
rect 3324 41684 3370 41722
rect 3324 41650 3330 41684
rect 3364 41650 3370 41684
rect 3324 41603 3370 41650
rect 3420 41828 3466 41875
rect 3420 41794 3426 41828
rect 3460 41794 3466 41828
rect 3420 41756 3466 41794
rect 3420 41722 3426 41756
rect 3460 41722 3466 41756
rect 3420 41684 3466 41722
rect 3420 41650 3426 41684
rect 3460 41650 3466 41684
rect 3420 41603 3466 41650
rect 3534 41859 3580 41897
rect 3534 41825 3540 41859
rect 3574 41825 3580 41859
rect 3534 41787 3580 41825
rect 3534 41753 3540 41787
rect 3574 41753 3580 41787
rect 3534 41715 3580 41753
rect 3534 41681 3540 41715
rect 3574 41681 3580 41715
rect 3534 41643 3580 41681
rect 3534 41609 3540 41643
rect 3574 41609 3580 41643
rect 2101 41458 2316 41462
rect 313 41428 2316 41458
rect 313 41424 2141 41428
rect 313 41291 347 41424
rect 505 41291 539 41424
rect 697 41291 731 41424
rect 889 41291 923 41424
rect 1081 41291 1115 41424
rect 1273 41291 1307 41424
rect 1381 41298 1608 41321
rect 307 41256 353 41291
rect 307 41222 313 41256
rect 347 41222 353 41256
rect 307 41187 353 41222
rect 403 41256 449 41291
rect 403 41222 409 41256
rect 443 41222 449 41256
rect 403 41187 449 41222
rect 499 41256 545 41291
rect 499 41222 505 41256
rect 539 41222 545 41256
rect 499 41187 545 41222
rect 595 41256 641 41291
rect 595 41222 601 41256
rect 635 41222 641 41256
rect 595 41187 641 41222
rect 691 41256 737 41291
rect 691 41222 697 41256
rect 731 41222 737 41256
rect 691 41187 737 41222
rect 787 41256 833 41291
rect 787 41222 793 41256
rect 827 41222 833 41256
rect 787 41187 833 41222
rect 883 41256 929 41291
rect 883 41222 889 41256
rect 923 41222 929 41256
rect 883 41187 929 41222
rect 979 41256 1025 41291
rect 979 41222 985 41256
rect 1019 41222 1025 41256
rect 979 41187 1025 41222
rect 1075 41256 1121 41291
rect 1075 41222 1081 41256
rect 1115 41222 1121 41256
rect 1075 41187 1121 41222
rect 1171 41256 1217 41291
rect 1171 41222 1177 41256
rect 1211 41222 1217 41256
rect 1171 41187 1217 41222
rect 1267 41256 1313 41291
rect 1267 41222 1273 41256
rect 1307 41222 1313 41256
rect 1267 41187 1313 41222
rect 1381 41264 1387 41298
rect 1421 41264 1608 41298
rect 1381 41226 1608 41264
rect 1381 41192 1387 41226
rect 1421 41201 1608 41226
rect 1421 41192 1427 41201
rect 1560 41199 1608 41201
rect 1598 41197 1608 41199
rect 1720 41197 1730 41321
rect 297 41156 363 41159
rect 294 41104 304 41156
rect 356 41104 366 41156
rect 297 41099 363 41104
rect 409 41047 443 41187
rect 489 41156 555 41159
rect 485 41104 495 41156
rect 547 41104 557 41156
rect 489 41099 555 41104
rect 601 41047 635 41187
rect 681 41156 747 41159
rect 677 41104 687 41156
rect 739 41104 749 41156
rect 681 41099 747 41104
rect 793 41047 827 41187
rect 873 41156 939 41159
rect 869 41104 879 41156
rect 931 41104 941 41156
rect 873 41099 939 41104
rect 985 41047 1019 41187
rect 1065 41155 1131 41159
rect 1062 41103 1072 41155
rect 1124 41103 1134 41155
rect 1065 41099 1131 41103
rect 1177 41047 1211 41187
rect 1257 41155 1323 41159
rect 1254 41103 1264 41155
rect 1316 41103 1326 41155
rect 1381 41154 1427 41192
rect 1920 41159 1930 41161
rect 1381 41120 1387 41154
rect 1421 41120 1427 41154
rect 1257 41099 1323 41103
rect 129 41013 1211 41047
rect 1381 40977 1427 41120
rect 1458 41103 1468 41159
rect 1524 41105 1930 41159
rect 1986 41105 1996 41161
rect 1524 41103 1986 41105
rect 2282 41051 2316 41428
rect 2466 41462 2500 41603
rect 2658 41462 2692 41603
rect 2850 41462 2884 41603
rect 3042 41462 3076 41603
rect 3234 41462 3268 41603
rect 3426 41462 3460 41603
rect 3534 41565 3580 41609
rect 3803 42025 4885 42059
rect 3803 41462 3837 42025
rect 3968 41915 3978 41967
rect 4030 41915 4040 41967
rect 4083 41875 4117 42025
rect 4161 41915 4171 41967
rect 4223 41915 4233 41967
rect 4275 41875 4309 42025
rect 4352 41915 4362 41967
rect 4414 41915 4424 41967
rect 4467 41875 4501 42025
rect 4544 41915 4554 41967
rect 4606 41915 4616 41967
rect 4659 41875 4693 42025
rect 4736 41915 4746 41967
rect 4798 41915 4808 41967
rect 4851 41875 4885 42025
rect 4928 41915 4938 41967
rect 4990 41915 5000 41967
rect 5055 41931 5101 42136
rect 5055 41897 5061 41931
rect 5095 41897 5101 41931
rect 3981 41828 4027 41875
rect 3981 41794 3987 41828
rect 4021 41794 4027 41828
rect 3981 41756 4027 41794
rect 3981 41722 3987 41756
rect 4021 41722 4027 41756
rect 3981 41684 4027 41722
rect 3981 41650 3987 41684
rect 4021 41650 4027 41684
rect 3981 41603 4027 41650
rect 4077 41828 4123 41875
rect 4077 41794 4083 41828
rect 4117 41794 4123 41828
rect 4077 41756 4123 41794
rect 4077 41722 4083 41756
rect 4117 41722 4123 41756
rect 4077 41684 4123 41722
rect 4077 41650 4083 41684
rect 4117 41650 4123 41684
rect 4077 41603 4123 41650
rect 4173 41828 4219 41875
rect 4173 41794 4179 41828
rect 4213 41794 4219 41828
rect 4173 41756 4219 41794
rect 4173 41722 4179 41756
rect 4213 41722 4219 41756
rect 4173 41684 4219 41722
rect 4173 41650 4179 41684
rect 4213 41650 4219 41684
rect 4173 41603 4219 41650
rect 4269 41828 4315 41875
rect 4269 41794 4275 41828
rect 4309 41794 4315 41828
rect 4269 41756 4315 41794
rect 4269 41722 4275 41756
rect 4309 41722 4315 41756
rect 4269 41684 4315 41722
rect 4269 41650 4275 41684
rect 4309 41650 4315 41684
rect 4269 41603 4315 41650
rect 4365 41828 4411 41875
rect 4365 41794 4371 41828
rect 4405 41794 4411 41828
rect 4365 41756 4411 41794
rect 4365 41722 4371 41756
rect 4405 41722 4411 41756
rect 4365 41684 4411 41722
rect 4365 41650 4371 41684
rect 4405 41650 4411 41684
rect 4365 41603 4411 41650
rect 4461 41828 4507 41875
rect 4461 41794 4467 41828
rect 4501 41794 4507 41828
rect 4461 41756 4507 41794
rect 4461 41722 4467 41756
rect 4501 41722 4507 41756
rect 4461 41684 4507 41722
rect 4461 41650 4467 41684
rect 4501 41650 4507 41684
rect 4461 41603 4507 41650
rect 4557 41828 4603 41875
rect 4557 41794 4563 41828
rect 4597 41794 4603 41828
rect 4557 41756 4603 41794
rect 4557 41722 4563 41756
rect 4597 41722 4603 41756
rect 4557 41684 4603 41722
rect 4557 41650 4563 41684
rect 4597 41650 4603 41684
rect 4557 41603 4603 41650
rect 4653 41828 4699 41875
rect 4653 41794 4659 41828
rect 4693 41794 4699 41828
rect 4653 41756 4699 41794
rect 4653 41722 4659 41756
rect 4693 41722 4699 41756
rect 4653 41684 4699 41722
rect 4653 41650 4659 41684
rect 4693 41650 4699 41684
rect 4653 41603 4699 41650
rect 4749 41828 4795 41875
rect 4749 41794 4755 41828
rect 4789 41794 4795 41828
rect 4749 41756 4795 41794
rect 4749 41722 4755 41756
rect 4789 41722 4795 41756
rect 4749 41684 4795 41722
rect 4749 41650 4755 41684
rect 4789 41650 4795 41684
rect 4749 41603 4795 41650
rect 4845 41828 4891 41875
rect 4845 41794 4851 41828
rect 4885 41794 4891 41828
rect 4845 41756 4891 41794
rect 4845 41722 4851 41756
rect 4885 41722 4891 41756
rect 4845 41684 4891 41722
rect 4845 41650 4851 41684
rect 4885 41650 4891 41684
rect 4845 41603 4891 41650
rect 4941 41828 4987 41875
rect 4941 41794 4947 41828
rect 4981 41794 4987 41828
rect 4941 41756 4987 41794
rect 4941 41722 4947 41756
rect 4981 41722 4987 41756
rect 4941 41684 4987 41722
rect 4941 41650 4947 41684
rect 4981 41650 4987 41684
rect 4941 41603 4987 41650
rect 5055 41859 5101 41897
rect 5055 41825 5061 41859
rect 5095 41825 5101 41859
rect 5055 41787 5101 41825
rect 5055 41753 5061 41787
rect 5095 41756 5101 41787
rect 5274 41756 5550 41757
rect 5095 41753 5550 41756
rect 5055 41726 5550 41753
rect 5055 41715 5303 41726
rect 5055 41681 5061 41715
rect 5095 41692 5303 41715
rect 5337 41692 5395 41726
rect 5429 41692 5487 41726
rect 5521 41692 5550 41726
rect 5095 41681 5550 41692
rect 5055 41661 5550 41681
rect 5055 41643 5101 41661
rect 5055 41609 5061 41643
rect 5095 41609 5101 41643
rect 2466 41428 3837 41462
rect 2466 41295 2500 41428
rect 2658 41295 2692 41428
rect 2850 41295 2884 41428
rect 3042 41295 3076 41428
rect 3234 41295 3268 41428
rect 3426 41295 3460 41428
rect 3671 41338 3681 41390
rect 3733 41338 3743 41390
rect 3679 41337 3691 41338
rect 3725 41337 3737 41338
rect 3679 41331 3737 41337
rect 3534 41302 3580 41325
rect 2460 41260 2506 41295
rect 2460 41226 2466 41260
rect 2500 41226 2506 41260
rect 2460 41191 2506 41226
rect 2556 41260 2602 41295
rect 2556 41226 2562 41260
rect 2596 41226 2602 41260
rect 2556 41191 2602 41226
rect 2652 41260 2698 41295
rect 2652 41226 2658 41260
rect 2692 41226 2698 41260
rect 2652 41191 2698 41226
rect 2748 41260 2794 41295
rect 2748 41226 2754 41260
rect 2788 41226 2794 41260
rect 2748 41191 2794 41226
rect 2844 41260 2890 41295
rect 2844 41226 2850 41260
rect 2884 41226 2890 41260
rect 2844 41191 2890 41226
rect 2940 41260 2986 41295
rect 2940 41226 2946 41260
rect 2980 41226 2986 41260
rect 2940 41191 2986 41226
rect 3036 41260 3082 41295
rect 3036 41226 3042 41260
rect 3076 41226 3082 41260
rect 3036 41191 3082 41226
rect 3132 41260 3178 41295
rect 3132 41226 3138 41260
rect 3172 41226 3178 41260
rect 3132 41191 3178 41226
rect 3228 41260 3274 41295
rect 3228 41226 3234 41260
rect 3268 41226 3274 41260
rect 3228 41191 3274 41226
rect 3324 41260 3370 41295
rect 3324 41226 3330 41260
rect 3364 41226 3370 41260
rect 3324 41191 3370 41226
rect 3420 41260 3466 41295
rect 3420 41226 3426 41260
rect 3460 41226 3466 41260
rect 3420 41191 3466 41226
rect 3534 41268 3540 41302
rect 3574 41300 3580 41302
rect 3803 41300 3837 41428
rect 3574 41299 3680 41300
rect 3734 41299 3837 41300
rect 3574 41287 3687 41299
rect 3574 41268 3647 41287
rect 3534 41230 3647 41268
rect 3534 41196 3540 41230
rect 3574 41211 3647 41230
rect 3681 41211 3687 41287
rect 3574 41200 3687 41211
rect 3574 41196 3580 41200
rect 3641 41199 3687 41200
rect 3729 41287 3837 41299
rect 3987 41462 4021 41603
rect 4179 41462 4213 41603
rect 4371 41462 4405 41603
rect 4563 41462 4597 41603
rect 4755 41462 4789 41603
rect 4947 41462 4981 41603
rect 5055 41565 5101 41609
rect 5177 41482 5882 41516
rect 5177 41462 5211 41482
rect 3987 41428 5211 41462
rect 3987 41295 4021 41428
rect 4179 41295 4213 41428
rect 4371 41295 4405 41428
rect 4563 41295 4597 41428
rect 4755 41295 4789 41428
rect 4947 41295 4981 41428
rect 5438 41424 5512 41425
rect 5326 41422 5400 41423
rect 5326 41370 5337 41422
rect 5389 41370 5400 41422
rect 5438 41372 5449 41424
rect 5501 41372 5512 41424
rect 5438 41371 5512 41372
rect 5683 41380 5882 41482
rect 5326 41369 5400 41370
rect 5055 41302 5101 41325
rect 3729 41211 3735 41287
rect 3769 41211 3837 41287
rect 3729 41200 3837 41211
rect 3729 41199 3775 41200
rect 2450 41160 2516 41163
rect 2447 41108 2457 41160
rect 2509 41108 2519 41160
rect 2450 41103 2516 41108
rect 2562 41051 2596 41191
rect 2642 41160 2708 41163
rect 2638 41108 2648 41160
rect 2700 41108 2710 41160
rect 2642 41103 2708 41108
rect 2754 41051 2788 41191
rect 2834 41160 2900 41163
rect 2830 41108 2840 41160
rect 2892 41108 2902 41160
rect 2834 41103 2900 41108
rect 2946 41051 2980 41191
rect 3026 41160 3092 41163
rect 3022 41108 3032 41160
rect 3084 41108 3094 41160
rect 3026 41103 3092 41108
rect 3138 41051 3172 41191
rect 3218 41159 3284 41163
rect 3215 41107 3225 41159
rect 3277 41107 3287 41159
rect 3218 41103 3284 41107
rect 3330 41051 3364 41191
rect 3410 41159 3476 41163
rect 3407 41107 3417 41159
rect 3469 41107 3479 41159
rect 3534 41158 3580 41196
rect 3534 41124 3540 41158
rect 3574 41124 3580 41158
rect 3410 41103 3476 41107
rect 2282 41017 3364 41051
rect 3534 40941 3580 41124
rect 3803 41051 3837 41200
rect 3981 41260 4027 41295
rect 3981 41226 3987 41260
rect 4021 41226 4027 41260
rect 3981 41191 4027 41226
rect 4077 41260 4123 41295
rect 4077 41226 4083 41260
rect 4117 41226 4123 41260
rect 4077 41191 4123 41226
rect 4173 41260 4219 41295
rect 4173 41226 4179 41260
rect 4213 41226 4219 41260
rect 4173 41191 4219 41226
rect 4269 41260 4315 41295
rect 4269 41226 4275 41260
rect 4309 41226 4315 41260
rect 4269 41191 4315 41226
rect 4365 41260 4411 41295
rect 4365 41226 4371 41260
rect 4405 41226 4411 41260
rect 4365 41191 4411 41226
rect 4461 41260 4507 41295
rect 4461 41226 4467 41260
rect 4501 41226 4507 41260
rect 4461 41191 4507 41226
rect 4557 41260 4603 41295
rect 4557 41226 4563 41260
rect 4597 41226 4603 41260
rect 4557 41191 4603 41226
rect 4653 41260 4699 41295
rect 4653 41226 4659 41260
rect 4693 41226 4699 41260
rect 4653 41191 4699 41226
rect 4749 41260 4795 41295
rect 4749 41226 4755 41260
rect 4789 41226 4795 41260
rect 4749 41191 4795 41226
rect 4845 41260 4891 41295
rect 4845 41226 4851 41260
rect 4885 41226 4891 41260
rect 4845 41191 4891 41226
rect 4941 41260 4987 41295
rect 4941 41226 4947 41260
rect 4981 41226 4987 41260
rect 4941 41191 4987 41226
rect 5055 41268 5061 41302
rect 5095 41268 5101 41302
rect 5055 41230 5101 41268
rect 5055 41196 5061 41230
rect 5095 41213 5101 41230
rect 5095 41196 5550 41213
rect 3971 41160 4037 41163
rect 3968 41108 3978 41160
rect 4030 41108 4040 41160
rect 3971 41103 4037 41108
rect 4083 41051 4117 41191
rect 4163 41160 4229 41163
rect 4159 41108 4169 41160
rect 4221 41108 4231 41160
rect 4163 41103 4229 41108
rect 4275 41051 4309 41191
rect 4355 41160 4421 41163
rect 4351 41108 4361 41160
rect 4413 41108 4423 41160
rect 4355 41103 4421 41108
rect 4467 41051 4501 41191
rect 4547 41160 4613 41163
rect 4543 41108 4553 41160
rect 4605 41108 4615 41160
rect 4547 41103 4613 41108
rect 4659 41051 4693 41191
rect 4739 41159 4805 41163
rect 4736 41107 4746 41159
rect 4798 41107 4808 41159
rect 4739 41103 4805 41107
rect 4851 41051 4885 41191
rect 5055 41182 5550 41196
rect 4931 41159 4997 41163
rect 4928 41107 4938 41159
rect 4990 41107 5000 41159
rect 5055 41158 5303 41182
rect 5055 41124 5061 41158
rect 5095 41148 5303 41158
rect 5337 41148 5395 41182
rect 5429 41148 5487 41182
rect 5521 41148 5550 41182
rect 5095 41124 5550 41148
rect 5055 41117 5550 41124
rect 4931 41103 4997 41107
rect 3803 41017 4885 41051
rect 5055 40942 5101 41117
rect 129 40734 1211 40768
rect 129 40171 163 40734
rect 294 40624 304 40676
rect 356 40624 366 40676
rect 409 40584 443 40734
rect 487 40624 497 40676
rect 549 40624 559 40676
rect 601 40584 635 40734
rect 678 40624 688 40676
rect 740 40624 750 40676
rect 793 40584 827 40734
rect 870 40624 880 40676
rect 932 40624 942 40676
rect 985 40584 1019 40734
rect 1062 40624 1072 40676
rect 1124 40624 1134 40676
rect 1177 40584 1211 40734
rect 1254 40624 1264 40676
rect 1316 40624 1326 40676
rect 1381 40640 1427 40804
rect 2282 40738 3364 40772
rect 1381 40606 1387 40640
rect 1421 40606 1427 40640
rect 1512 40617 1522 40677
rect 1578 40617 1792 40677
rect 1852 40617 1862 40677
rect 307 40537 353 40584
rect 307 40503 313 40537
rect 347 40503 353 40537
rect 307 40465 353 40503
rect 307 40431 313 40465
rect 347 40431 353 40465
rect 307 40393 353 40431
rect 307 40359 313 40393
rect 347 40359 353 40393
rect 307 40312 353 40359
rect 403 40537 449 40584
rect 403 40503 409 40537
rect 443 40503 449 40537
rect 403 40465 449 40503
rect 403 40431 409 40465
rect 443 40431 449 40465
rect 403 40393 449 40431
rect 403 40359 409 40393
rect 443 40359 449 40393
rect 403 40312 449 40359
rect 499 40537 545 40584
rect 499 40503 505 40537
rect 539 40503 545 40537
rect 499 40465 545 40503
rect 499 40431 505 40465
rect 539 40431 545 40465
rect 499 40393 545 40431
rect 499 40359 505 40393
rect 539 40359 545 40393
rect 499 40312 545 40359
rect 595 40537 641 40584
rect 595 40503 601 40537
rect 635 40503 641 40537
rect 595 40465 641 40503
rect 595 40431 601 40465
rect 635 40431 641 40465
rect 595 40393 641 40431
rect 595 40359 601 40393
rect 635 40359 641 40393
rect 595 40312 641 40359
rect 691 40537 737 40584
rect 691 40503 697 40537
rect 731 40503 737 40537
rect 691 40465 737 40503
rect 691 40431 697 40465
rect 731 40431 737 40465
rect 691 40393 737 40431
rect 691 40359 697 40393
rect 731 40359 737 40393
rect 691 40312 737 40359
rect 787 40537 833 40584
rect 787 40503 793 40537
rect 827 40503 833 40537
rect 787 40465 833 40503
rect 787 40431 793 40465
rect 827 40431 833 40465
rect 787 40393 833 40431
rect 787 40359 793 40393
rect 827 40359 833 40393
rect 787 40312 833 40359
rect 883 40537 929 40584
rect 883 40503 889 40537
rect 923 40503 929 40537
rect 883 40465 929 40503
rect 883 40431 889 40465
rect 923 40431 929 40465
rect 883 40393 929 40431
rect 883 40359 889 40393
rect 923 40359 929 40393
rect 883 40312 929 40359
rect 979 40537 1025 40584
rect 979 40503 985 40537
rect 1019 40503 1025 40537
rect 979 40465 1025 40503
rect 979 40431 985 40465
rect 1019 40431 1025 40465
rect 979 40393 1025 40431
rect 979 40359 985 40393
rect 1019 40359 1025 40393
rect 979 40312 1025 40359
rect 1075 40537 1121 40584
rect 1075 40503 1081 40537
rect 1115 40503 1121 40537
rect 1075 40465 1121 40503
rect 1075 40431 1081 40465
rect 1115 40431 1121 40465
rect 1075 40393 1121 40431
rect 1075 40359 1081 40393
rect 1115 40359 1121 40393
rect 1075 40312 1121 40359
rect 1171 40537 1217 40584
rect 1171 40503 1177 40537
rect 1211 40503 1217 40537
rect 1171 40465 1217 40503
rect 1171 40431 1177 40465
rect 1211 40431 1217 40465
rect 1171 40393 1217 40431
rect 1171 40359 1177 40393
rect 1211 40359 1217 40393
rect 1171 40312 1217 40359
rect 1267 40537 1313 40584
rect 1267 40503 1273 40537
rect 1307 40503 1313 40537
rect 1267 40465 1313 40503
rect 1267 40431 1273 40465
rect 1307 40431 1313 40465
rect 1267 40393 1313 40431
rect 1267 40359 1273 40393
rect 1307 40359 1313 40393
rect 1267 40312 1313 40359
rect 1381 40568 1427 40606
rect 1381 40534 1387 40568
rect 1421 40534 1427 40568
rect 1381 40496 1427 40534
rect 1381 40462 1387 40496
rect 1421 40462 1427 40496
rect 1381 40424 1427 40462
rect 1381 40390 1387 40424
rect 1421 40390 1427 40424
rect 1381 40380 1427 40390
rect 1381 40378 2160 40380
rect 1381 40352 2056 40378
rect 1381 40327 1387 40352
rect 1380 40318 1387 40327
rect 1421 40318 2056 40352
rect 0 40137 163 40171
rect 129 39760 163 40137
rect 313 40171 347 40312
rect 505 40171 539 40312
rect 697 40171 731 40312
rect 889 40171 923 40312
rect 1081 40171 1115 40312
rect 1273 40171 1307 40312
rect 1380 40270 2056 40318
rect 2190 40270 2200 40378
rect 1380 40268 2160 40270
rect 2282 40175 2316 40738
rect 2447 40628 2457 40680
rect 2509 40628 2519 40680
rect 2562 40588 2596 40738
rect 2640 40628 2650 40680
rect 2702 40628 2712 40680
rect 2754 40588 2788 40738
rect 2831 40628 2841 40680
rect 2893 40628 2903 40680
rect 2946 40588 2980 40738
rect 3023 40628 3033 40680
rect 3085 40628 3095 40680
rect 3138 40588 3172 40738
rect 3215 40628 3225 40680
rect 3277 40628 3287 40680
rect 3330 40588 3364 40738
rect 3407 40628 3417 40680
rect 3469 40628 3479 40680
rect 3534 40644 3580 40852
rect 3534 40610 3540 40644
rect 3574 40610 3580 40644
rect 2460 40541 2506 40588
rect 2460 40507 2466 40541
rect 2500 40507 2506 40541
rect 2460 40469 2506 40507
rect 2460 40435 2466 40469
rect 2500 40435 2506 40469
rect 2460 40397 2506 40435
rect 2460 40363 2466 40397
rect 2500 40363 2506 40397
rect 2460 40316 2506 40363
rect 2556 40541 2602 40588
rect 2556 40507 2562 40541
rect 2596 40507 2602 40541
rect 2556 40469 2602 40507
rect 2556 40435 2562 40469
rect 2596 40435 2602 40469
rect 2556 40397 2602 40435
rect 2556 40363 2562 40397
rect 2596 40363 2602 40397
rect 2556 40316 2602 40363
rect 2652 40541 2698 40588
rect 2652 40507 2658 40541
rect 2692 40507 2698 40541
rect 2652 40469 2698 40507
rect 2652 40435 2658 40469
rect 2692 40435 2698 40469
rect 2652 40397 2698 40435
rect 2652 40363 2658 40397
rect 2692 40363 2698 40397
rect 2652 40316 2698 40363
rect 2748 40541 2794 40588
rect 2748 40507 2754 40541
rect 2788 40507 2794 40541
rect 2748 40469 2794 40507
rect 2748 40435 2754 40469
rect 2788 40435 2794 40469
rect 2748 40397 2794 40435
rect 2748 40363 2754 40397
rect 2788 40363 2794 40397
rect 2748 40316 2794 40363
rect 2844 40541 2890 40588
rect 2844 40507 2850 40541
rect 2884 40507 2890 40541
rect 2844 40469 2890 40507
rect 2844 40435 2850 40469
rect 2884 40435 2890 40469
rect 2844 40397 2890 40435
rect 2844 40363 2850 40397
rect 2884 40363 2890 40397
rect 2844 40316 2890 40363
rect 2940 40541 2986 40588
rect 2940 40507 2946 40541
rect 2980 40507 2986 40541
rect 2940 40469 2986 40507
rect 2940 40435 2946 40469
rect 2980 40435 2986 40469
rect 2940 40397 2986 40435
rect 2940 40363 2946 40397
rect 2980 40363 2986 40397
rect 2940 40316 2986 40363
rect 3036 40541 3082 40588
rect 3036 40507 3042 40541
rect 3076 40507 3082 40541
rect 3036 40469 3082 40507
rect 3036 40435 3042 40469
rect 3076 40435 3082 40469
rect 3036 40397 3082 40435
rect 3036 40363 3042 40397
rect 3076 40363 3082 40397
rect 3036 40316 3082 40363
rect 3132 40541 3178 40588
rect 3132 40507 3138 40541
rect 3172 40507 3178 40541
rect 3132 40469 3178 40507
rect 3132 40435 3138 40469
rect 3172 40435 3178 40469
rect 3132 40397 3178 40435
rect 3132 40363 3138 40397
rect 3172 40363 3178 40397
rect 3132 40316 3178 40363
rect 3228 40541 3274 40588
rect 3228 40507 3234 40541
rect 3268 40507 3274 40541
rect 3228 40469 3274 40507
rect 3228 40435 3234 40469
rect 3268 40435 3274 40469
rect 3228 40397 3274 40435
rect 3228 40363 3234 40397
rect 3268 40363 3274 40397
rect 3228 40316 3274 40363
rect 3324 40541 3370 40588
rect 3324 40507 3330 40541
rect 3364 40507 3370 40541
rect 3324 40469 3370 40507
rect 3324 40435 3330 40469
rect 3364 40435 3370 40469
rect 3324 40397 3370 40435
rect 3324 40363 3330 40397
rect 3364 40363 3370 40397
rect 3324 40316 3370 40363
rect 3420 40541 3466 40588
rect 3420 40507 3426 40541
rect 3460 40507 3466 40541
rect 3420 40469 3466 40507
rect 3420 40435 3426 40469
rect 3460 40435 3466 40469
rect 3420 40397 3466 40435
rect 3420 40363 3426 40397
rect 3460 40363 3466 40397
rect 3420 40316 3466 40363
rect 3534 40572 3580 40610
rect 3534 40538 3540 40572
rect 3574 40538 3580 40572
rect 3534 40500 3580 40538
rect 3534 40466 3540 40500
rect 3574 40466 3580 40500
rect 3534 40428 3580 40466
rect 3534 40394 3540 40428
rect 3574 40394 3580 40428
rect 3534 40356 3580 40394
rect 3534 40322 3540 40356
rect 3574 40322 3580 40356
rect 2101 40171 2316 40175
rect 313 40141 2316 40171
rect 313 40137 2141 40141
rect 313 40004 347 40137
rect 505 40004 539 40137
rect 697 40004 731 40137
rect 889 40004 923 40137
rect 1081 40004 1115 40137
rect 1273 40004 1307 40137
rect 1381 40011 1608 40034
rect 307 39969 353 40004
rect 307 39935 313 39969
rect 347 39935 353 39969
rect 307 39900 353 39935
rect 403 39969 449 40004
rect 403 39935 409 39969
rect 443 39935 449 39969
rect 403 39900 449 39935
rect 499 39969 545 40004
rect 499 39935 505 39969
rect 539 39935 545 39969
rect 499 39900 545 39935
rect 595 39969 641 40004
rect 595 39935 601 39969
rect 635 39935 641 39969
rect 595 39900 641 39935
rect 691 39969 737 40004
rect 691 39935 697 39969
rect 731 39935 737 39969
rect 691 39900 737 39935
rect 787 39969 833 40004
rect 787 39935 793 39969
rect 827 39935 833 39969
rect 787 39900 833 39935
rect 883 39969 929 40004
rect 883 39935 889 39969
rect 923 39935 929 39969
rect 883 39900 929 39935
rect 979 39969 1025 40004
rect 979 39935 985 39969
rect 1019 39935 1025 39969
rect 979 39900 1025 39935
rect 1075 39969 1121 40004
rect 1075 39935 1081 39969
rect 1115 39935 1121 39969
rect 1075 39900 1121 39935
rect 1171 39969 1217 40004
rect 1171 39935 1177 39969
rect 1211 39935 1217 39969
rect 1171 39900 1217 39935
rect 1267 39969 1313 40004
rect 1267 39935 1273 39969
rect 1307 39935 1313 39969
rect 1267 39900 1313 39935
rect 1381 39977 1387 40011
rect 1421 39977 1608 40011
rect 1381 39939 1608 39977
rect 1381 39905 1387 39939
rect 1421 39914 1608 39939
rect 1421 39905 1427 39914
rect 1560 39912 1608 39914
rect 1598 39910 1608 39912
rect 1720 39910 1730 40034
rect 297 39869 363 39872
rect 294 39817 304 39869
rect 356 39817 366 39869
rect 297 39812 363 39817
rect 409 39760 443 39900
rect 489 39869 555 39872
rect 485 39817 495 39869
rect 547 39817 557 39869
rect 489 39812 555 39817
rect 601 39760 635 39900
rect 681 39869 747 39872
rect 677 39817 687 39869
rect 739 39817 749 39869
rect 681 39812 747 39817
rect 793 39760 827 39900
rect 873 39869 939 39872
rect 869 39817 879 39869
rect 931 39817 941 39869
rect 873 39812 939 39817
rect 985 39760 1019 39900
rect 1065 39868 1131 39872
rect 1062 39816 1072 39868
rect 1124 39816 1134 39868
rect 1065 39812 1131 39816
rect 1177 39760 1211 39900
rect 1257 39868 1323 39872
rect 1254 39816 1264 39868
rect 1316 39816 1326 39868
rect 1381 39867 1427 39905
rect 1920 39872 1930 39874
rect 1381 39833 1387 39867
rect 1421 39833 1427 39867
rect 1257 39812 1323 39816
rect 129 39726 1211 39760
rect 1381 39690 1427 39833
rect 1458 39816 1468 39872
rect 1524 39818 1930 39872
rect 1986 39818 1996 39874
rect 1524 39816 1986 39818
rect 2282 39764 2316 40141
rect 2466 40175 2500 40316
rect 2658 40175 2692 40316
rect 2850 40175 2884 40316
rect 3042 40175 3076 40316
rect 3234 40175 3268 40316
rect 3426 40175 3460 40316
rect 3534 40278 3580 40322
rect 3803 40738 4885 40772
rect 3803 40175 3837 40738
rect 3968 40628 3978 40680
rect 4030 40628 4040 40680
rect 4083 40588 4117 40738
rect 4161 40628 4171 40680
rect 4223 40628 4233 40680
rect 4275 40588 4309 40738
rect 4352 40628 4362 40680
rect 4414 40628 4424 40680
rect 4467 40588 4501 40738
rect 4544 40628 4554 40680
rect 4606 40628 4616 40680
rect 4659 40588 4693 40738
rect 4736 40628 4746 40680
rect 4798 40628 4808 40680
rect 4851 40588 4885 40738
rect 4928 40628 4938 40680
rect 4990 40628 5000 40680
rect 5055 40644 5101 40849
rect 5055 40610 5061 40644
rect 5095 40610 5101 40644
rect 3981 40541 4027 40588
rect 3981 40507 3987 40541
rect 4021 40507 4027 40541
rect 3981 40469 4027 40507
rect 3981 40435 3987 40469
rect 4021 40435 4027 40469
rect 3981 40397 4027 40435
rect 3981 40363 3987 40397
rect 4021 40363 4027 40397
rect 3981 40316 4027 40363
rect 4077 40541 4123 40588
rect 4077 40507 4083 40541
rect 4117 40507 4123 40541
rect 4077 40469 4123 40507
rect 4077 40435 4083 40469
rect 4117 40435 4123 40469
rect 4077 40397 4123 40435
rect 4077 40363 4083 40397
rect 4117 40363 4123 40397
rect 4077 40316 4123 40363
rect 4173 40541 4219 40588
rect 4173 40507 4179 40541
rect 4213 40507 4219 40541
rect 4173 40469 4219 40507
rect 4173 40435 4179 40469
rect 4213 40435 4219 40469
rect 4173 40397 4219 40435
rect 4173 40363 4179 40397
rect 4213 40363 4219 40397
rect 4173 40316 4219 40363
rect 4269 40541 4315 40588
rect 4269 40507 4275 40541
rect 4309 40507 4315 40541
rect 4269 40469 4315 40507
rect 4269 40435 4275 40469
rect 4309 40435 4315 40469
rect 4269 40397 4315 40435
rect 4269 40363 4275 40397
rect 4309 40363 4315 40397
rect 4269 40316 4315 40363
rect 4365 40541 4411 40588
rect 4365 40507 4371 40541
rect 4405 40507 4411 40541
rect 4365 40469 4411 40507
rect 4365 40435 4371 40469
rect 4405 40435 4411 40469
rect 4365 40397 4411 40435
rect 4365 40363 4371 40397
rect 4405 40363 4411 40397
rect 4365 40316 4411 40363
rect 4461 40541 4507 40588
rect 4461 40507 4467 40541
rect 4501 40507 4507 40541
rect 4461 40469 4507 40507
rect 4461 40435 4467 40469
rect 4501 40435 4507 40469
rect 4461 40397 4507 40435
rect 4461 40363 4467 40397
rect 4501 40363 4507 40397
rect 4461 40316 4507 40363
rect 4557 40541 4603 40588
rect 4557 40507 4563 40541
rect 4597 40507 4603 40541
rect 4557 40469 4603 40507
rect 4557 40435 4563 40469
rect 4597 40435 4603 40469
rect 4557 40397 4603 40435
rect 4557 40363 4563 40397
rect 4597 40363 4603 40397
rect 4557 40316 4603 40363
rect 4653 40541 4699 40588
rect 4653 40507 4659 40541
rect 4693 40507 4699 40541
rect 4653 40469 4699 40507
rect 4653 40435 4659 40469
rect 4693 40435 4699 40469
rect 4653 40397 4699 40435
rect 4653 40363 4659 40397
rect 4693 40363 4699 40397
rect 4653 40316 4699 40363
rect 4749 40541 4795 40588
rect 4749 40507 4755 40541
rect 4789 40507 4795 40541
rect 4749 40469 4795 40507
rect 4749 40435 4755 40469
rect 4789 40435 4795 40469
rect 4749 40397 4795 40435
rect 4749 40363 4755 40397
rect 4789 40363 4795 40397
rect 4749 40316 4795 40363
rect 4845 40541 4891 40588
rect 4845 40507 4851 40541
rect 4885 40507 4891 40541
rect 4845 40469 4891 40507
rect 4845 40435 4851 40469
rect 4885 40435 4891 40469
rect 4845 40397 4891 40435
rect 4845 40363 4851 40397
rect 4885 40363 4891 40397
rect 4845 40316 4891 40363
rect 4941 40541 4987 40588
rect 4941 40507 4947 40541
rect 4981 40507 4987 40541
rect 4941 40469 4987 40507
rect 4941 40435 4947 40469
rect 4981 40435 4987 40469
rect 4941 40397 4987 40435
rect 4941 40363 4947 40397
rect 4981 40363 4987 40397
rect 4941 40316 4987 40363
rect 5055 40572 5101 40610
rect 5055 40538 5061 40572
rect 5095 40538 5101 40572
rect 5055 40500 5101 40538
rect 5055 40466 5061 40500
rect 5095 40469 5101 40500
rect 5274 40469 5550 40470
rect 5095 40466 5550 40469
rect 5055 40439 5550 40466
rect 5055 40428 5303 40439
rect 5055 40394 5061 40428
rect 5095 40405 5303 40428
rect 5337 40405 5395 40439
rect 5429 40405 5487 40439
rect 5521 40405 5550 40439
rect 5095 40394 5550 40405
rect 5055 40374 5550 40394
rect 5055 40356 5101 40374
rect 5055 40322 5061 40356
rect 5095 40322 5101 40356
rect 2466 40141 3837 40175
rect 2466 40008 2500 40141
rect 2658 40008 2692 40141
rect 2850 40008 2884 40141
rect 3042 40008 3076 40141
rect 3234 40008 3268 40141
rect 3426 40008 3460 40141
rect 3671 40051 3681 40103
rect 3733 40051 3743 40103
rect 3679 40050 3691 40051
rect 3725 40050 3737 40051
rect 3679 40044 3737 40050
rect 3534 40015 3580 40038
rect 2460 39973 2506 40008
rect 2460 39939 2466 39973
rect 2500 39939 2506 39973
rect 2460 39904 2506 39939
rect 2556 39973 2602 40008
rect 2556 39939 2562 39973
rect 2596 39939 2602 39973
rect 2556 39904 2602 39939
rect 2652 39973 2698 40008
rect 2652 39939 2658 39973
rect 2692 39939 2698 39973
rect 2652 39904 2698 39939
rect 2748 39973 2794 40008
rect 2748 39939 2754 39973
rect 2788 39939 2794 39973
rect 2748 39904 2794 39939
rect 2844 39973 2890 40008
rect 2844 39939 2850 39973
rect 2884 39939 2890 39973
rect 2844 39904 2890 39939
rect 2940 39973 2986 40008
rect 2940 39939 2946 39973
rect 2980 39939 2986 39973
rect 2940 39904 2986 39939
rect 3036 39973 3082 40008
rect 3036 39939 3042 39973
rect 3076 39939 3082 39973
rect 3036 39904 3082 39939
rect 3132 39973 3178 40008
rect 3132 39939 3138 39973
rect 3172 39939 3178 39973
rect 3132 39904 3178 39939
rect 3228 39973 3274 40008
rect 3228 39939 3234 39973
rect 3268 39939 3274 39973
rect 3228 39904 3274 39939
rect 3324 39973 3370 40008
rect 3324 39939 3330 39973
rect 3364 39939 3370 39973
rect 3324 39904 3370 39939
rect 3420 39973 3466 40008
rect 3420 39939 3426 39973
rect 3460 39939 3466 39973
rect 3420 39904 3466 39939
rect 3534 39981 3540 40015
rect 3574 40013 3580 40015
rect 3803 40013 3837 40141
rect 3574 40012 3680 40013
rect 3734 40012 3837 40013
rect 3574 40000 3687 40012
rect 3574 39981 3647 40000
rect 3534 39943 3647 39981
rect 3534 39909 3540 39943
rect 3574 39924 3647 39943
rect 3681 39924 3687 40000
rect 3574 39913 3687 39924
rect 3574 39909 3580 39913
rect 3641 39912 3687 39913
rect 3729 40000 3837 40012
rect 3987 40175 4021 40316
rect 4179 40175 4213 40316
rect 4371 40175 4405 40316
rect 4563 40175 4597 40316
rect 4755 40175 4789 40316
rect 4947 40175 4981 40316
rect 5055 40278 5101 40322
rect 5683 40229 5743 41380
rect 5177 40195 5743 40229
rect 5177 40175 5211 40195
rect 3987 40141 5211 40175
rect 3987 40008 4021 40141
rect 4179 40008 4213 40141
rect 4371 40008 4405 40141
rect 4563 40008 4597 40141
rect 4755 40008 4789 40141
rect 4947 40008 4981 40141
rect 5438 40137 5512 40138
rect 5326 40135 5400 40136
rect 5326 40083 5337 40135
rect 5389 40083 5400 40135
rect 5438 40085 5449 40137
rect 5501 40085 5512 40137
rect 5438 40084 5512 40085
rect 5326 40082 5400 40083
rect 5055 40015 5101 40038
rect 3729 39924 3735 40000
rect 3769 39924 3837 40000
rect 3729 39913 3837 39924
rect 3729 39912 3775 39913
rect 2450 39873 2516 39876
rect 2447 39821 2457 39873
rect 2509 39821 2519 39873
rect 2450 39816 2516 39821
rect 2562 39764 2596 39904
rect 2642 39873 2708 39876
rect 2638 39821 2648 39873
rect 2700 39821 2710 39873
rect 2642 39816 2708 39821
rect 2754 39764 2788 39904
rect 2834 39873 2900 39876
rect 2830 39821 2840 39873
rect 2892 39821 2902 39873
rect 2834 39816 2900 39821
rect 2946 39764 2980 39904
rect 3026 39873 3092 39876
rect 3022 39821 3032 39873
rect 3084 39821 3094 39873
rect 3026 39816 3092 39821
rect 3138 39764 3172 39904
rect 3218 39872 3284 39876
rect 3215 39820 3225 39872
rect 3277 39820 3287 39872
rect 3218 39816 3284 39820
rect 3330 39764 3364 39904
rect 3410 39872 3476 39876
rect 3407 39820 3417 39872
rect 3469 39820 3479 39872
rect 3534 39871 3580 39909
rect 3534 39837 3540 39871
rect 3574 39837 3580 39871
rect 3410 39816 3476 39820
rect 2282 39730 3364 39764
rect 3534 39654 3580 39837
rect 3803 39764 3837 39913
rect 3981 39973 4027 40008
rect 3981 39939 3987 39973
rect 4021 39939 4027 39973
rect 3981 39904 4027 39939
rect 4077 39973 4123 40008
rect 4077 39939 4083 39973
rect 4117 39939 4123 39973
rect 4077 39904 4123 39939
rect 4173 39973 4219 40008
rect 4173 39939 4179 39973
rect 4213 39939 4219 39973
rect 4173 39904 4219 39939
rect 4269 39973 4315 40008
rect 4269 39939 4275 39973
rect 4309 39939 4315 39973
rect 4269 39904 4315 39939
rect 4365 39973 4411 40008
rect 4365 39939 4371 39973
rect 4405 39939 4411 39973
rect 4365 39904 4411 39939
rect 4461 39973 4507 40008
rect 4461 39939 4467 39973
rect 4501 39939 4507 39973
rect 4461 39904 4507 39939
rect 4557 39973 4603 40008
rect 4557 39939 4563 39973
rect 4597 39939 4603 39973
rect 4557 39904 4603 39939
rect 4653 39973 4699 40008
rect 4653 39939 4659 39973
rect 4693 39939 4699 39973
rect 4653 39904 4699 39939
rect 4749 39973 4795 40008
rect 4749 39939 4755 39973
rect 4789 39939 4795 39973
rect 4749 39904 4795 39939
rect 4845 39973 4891 40008
rect 4845 39939 4851 39973
rect 4885 39939 4891 39973
rect 4845 39904 4891 39939
rect 4941 39973 4987 40008
rect 4941 39939 4947 39973
rect 4981 39939 4987 39973
rect 4941 39904 4987 39939
rect 5055 39981 5061 40015
rect 5095 39981 5101 40015
rect 5055 39943 5101 39981
rect 5055 39909 5061 39943
rect 5095 39926 5101 39943
rect 5095 39909 5550 39926
rect 3971 39873 4037 39876
rect 3968 39821 3978 39873
rect 4030 39821 4040 39873
rect 3971 39816 4037 39821
rect 4083 39764 4117 39904
rect 4163 39873 4229 39876
rect 4159 39821 4169 39873
rect 4221 39821 4231 39873
rect 4163 39816 4229 39821
rect 4275 39764 4309 39904
rect 4355 39873 4421 39876
rect 4351 39821 4361 39873
rect 4413 39821 4423 39873
rect 4355 39816 4421 39821
rect 4467 39764 4501 39904
rect 4547 39873 4613 39876
rect 4543 39821 4553 39873
rect 4605 39821 4615 39873
rect 4547 39816 4613 39821
rect 4659 39764 4693 39904
rect 4739 39872 4805 39876
rect 4736 39820 4746 39872
rect 4798 39820 4808 39872
rect 4739 39816 4805 39820
rect 4851 39764 4885 39904
rect 5055 39895 5550 39909
rect 4931 39872 4997 39876
rect 4928 39820 4938 39872
rect 4990 39820 5000 39872
rect 5055 39871 5303 39895
rect 5055 39837 5061 39871
rect 5095 39861 5303 39871
rect 5337 39861 5395 39895
rect 5429 39861 5487 39895
rect 5521 39861 5550 39895
rect 5095 39837 5550 39861
rect 5055 39830 5550 39837
rect 4931 39816 4997 39820
rect 3803 39730 4885 39764
rect 5055 39655 5101 39830
rect 129 39447 1211 39481
rect 129 38884 163 39447
rect 294 39337 304 39389
rect 356 39337 366 39389
rect 409 39297 443 39447
rect 487 39337 497 39389
rect 549 39337 559 39389
rect 601 39297 635 39447
rect 678 39337 688 39389
rect 740 39337 750 39389
rect 793 39297 827 39447
rect 870 39337 880 39389
rect 932 39337 942 39389
rect 985 39297 1019 39447
rect 1062 39337 1072 39389
rect 1124 39337 1134 39389
rect 1177 39297 1211 39447
rect 1254 39337 1264 39389
rect 1316 39337 1326 39389
rect 1381 39353 1427 39517
rect 2282 39451 3364 39485
rect 1381 39319 1387 39353
rect 1421 39319 1427 39353
rect 1512 39330 1522 39390
rect 1578 39330 1792 39390
rect 1852 39330 1862 39390
rect 307 39250 353 39297
rect 307 39216 313 39250
rect 347 39216 353 39250
rect 307 39178 353 39216
rect 307 39144 313 39178
rect 347 39144 353 39178
rect 307 39106 353 39144
rect 307 39072 313 39106
rect 347 39072 353 39106
rect 307 39025 353 39072
rect 403 39250 449 39297
rect 403 39216 409 39250
rect 443 39216 449 39250
rect 403 39178 449 39216
rect 403 39144 409 39178
rect 443 39144 449 39178
rect 403 39106 449 39144
rect 403 39072 409 39106
rect 443 39072 449 39106
rect 403 39025 449 39072
rect 499 39250 545 39297
rect 499 39216 505 39250
rect 539 39216 545 39250
rect 499 39178 545 39216
rect 499 39144 505 39178
rect 539 39144 545 39178
rect 499 39106 545 39144
rect 499 39072 505 39106
rect 539 39072 545 39106
rect 499 39025 545 39072
rect 595 39250 641 39297
rect 595 39216 601 39250
rect 635 39216 641 39250
rect 595 39178 641 39216
rect 595 39144 601 39178
rect 635 39144 641 39178
rect 595 39106 641 39144
rect 595 39072 601 39106
rect 635 39072 641 39106
rect 595 39025 641 39072
rect 691 39250 737 39297
rect 691 39216 697 39250
rect 731 39216 737 39250
rect 691 39178 737 39216
rect 691 39144 697 39178
rect 731 39144 737 39178
rect 691 39106 737 39144
rect 691 39072 697 39106
rect 731 39072 737 39106
rect 691 39025 737 39072
rect 787 39250 833 39297
rect 787 39216 793 39250
rect 827 39216 833 39250
rect 787 39178 833 39216
rect 787 39144 793 39178
rect 827 39144 833 39178
rect 787 39106 833 39144
rect 787 39072 793 39106
rect 827 39072 833 39106
rect 787 39025 833 39072
rect 883 39250 929 39297
rect 883 39216 889 39250
rect 923 39216 929 39250
rect 883 39178 929 39216
rect 883 39144 889 39178
rect 923 39144 929 39178
rect 883 39106 929 39144
rect 883 39072 889 39106
rect 923 39072 929 39106
rect 883 39025 929 39072
rect 979 39250 1025 39297
rect 979 39216 985 39250
rect 1019 39216 1025 39250
rect 979 39178 1025 39216
rect 979 39144 985 39178
rect 1019 39144 1025 39178
rect 979 39106 1025 39144
rect 979 39072 985 39106
rect 1019 39072 1025 39106
rect 979 39025 1025 39072
rect 1075 39250 1121 39297
rect 1075 39216 1081 39250
rect 1115 39216 1121 39250
rect 1075 39178 1121 39216
rect 1075 39144 1081 39178
rect 1115 39144 1121 39178
rect 1075 39106 1121 39144
rect 1075 39072 1081 39106
rect 1115 39072 1121 39106
rect 1075 39025 1121 39072
rect 1171 39250 1217 39297
rect 1171 39216 1177 39250
rect 1211 39216 1217 39250
rect 1171 39178 1217 39216
rect 1171 39144 1177 39178
rect 1211 39144 1217 39178
rect 1171 39106 1217 39144
rect 1171 39072 1177 39106
rect 1211 39072 1217 39106
rect 1171 39025 1217 39072
rect 1267 39250 1313 39297
rect 1267 39216 1273 39250
rect 1307 39216 1313 39250
rect 1267 39178 1313 39216
rect 1267 39144 1273 39178
rect 1307 39144 1313 39178
rect 1267 39106 1313 39144
rect 1267 39072 1273 39106
rect 1307 39072 1313 39106
rect 1267 39025 1313 39072
rect 1381 39281 1427 39319
rect 1381 39247 1387 39281
rect 1421 39247 1427 39281
rect 1381 39209 1427 39247
rect 1381 39175 1387 39209
rect 1421 39175 1427 39209
rect 1381 39137 1427 39175
rect 1381 39103 1387 39137
rect 1421 39103 1427 39137
rect 1381 39093 1427 39103
rect 1381 39091 2160 39093
rect 1381 39065 2056 39091
rect 1381 39040 1387 39065
rect 1380 39031 1387 39040
rect 1421 39031 2056 39065
rect 0 38850 163 38884
rect 129 38473 163 38850
rect 313 38884 347 39025
rect 505 38884 539 39025
rect 697 38884 731 39025
rect 889 38884 923 39025
rect 1081 38884 1115 39025
rect 1273 38884 1307 39025
rect 1380 38983 2056 39031
rect 2190 38983 2200 39091
rect 1380 38981 2160 38983
rect 2282 38888 2316 39451
rect 2447 39341 2457 39393
rect 2509 39341 2519 39393
rect 2562 39301 2596 39451
rect 2640 39341 2650 39393
rect 2702 39341 2712 39393
rect 2754 39301 2788 39451
rect 2831 39341 2841 39393
rect 2893 39341 2903 39393
rect 2946 39301 2980 39451
rect 3023 39341 3033 39393
rect 3085 39341 3095 39393
rect 3138 39301 3172 39451
rect 3215 39341 3225 39393
rect 3277 39341 3287 39393
rect 3330 39301 3364 39451
rect 3407 39341 3417 39393
rect 3469 39341 3479 39393
rect 3534 39357 3580 39565
rect 3534 39323 3540 39357
rect 3574 39323 3580 39357
rect 2460 39254 2506 39301
rect 2460 39220 2466 39254
rect 2500 39220 2506 39254
rect 2460 39182 2506 39220
rect 2460 39148 2466 39182
rect 2500 39148 2506 39182
rect 2460 39110 2506 39148
rect 2460 39076 2466 39110
rect 2500 39076 2506 39110
rect 2460 39029 2506 39076
rect 2556 39254 2602 39301
rect 2556 39220 2562 39254
rect 2596 39220 2602 39254
rect 2556 39182 2602 39220
rect 2556 39148 2562 39182
rect 2596 39148 2602 39182
rect 2556 39110 2602 39148
rect 2556 39076 2562 39110
rect 2596 39076 2602 39110
rect 2556 39029 2602 39076
rect 2652 39254 2698 39301
rect 2652 39220 2658 39254
rect 2692 39220 2698 39254
rect 2652 39182 2698 39220
rect 2652 39148 2658 39182
rect 2692 39148 2698 39182
rect 2652 39110 2698 39148
rect 2652 39076 2658 39110
rect 2692 39076 2698 39110
rect 2652 39029 2698 39076
rect 2748 39254 2794 39301
rect 2748 39220 2754 39254
rect 2788 39220 2794 39254
rect 2748 39182 2794 39220
rect 2748 39148 2754 39182
rect 2788 39148 2794 39182
rect 2748 39110 2794 39148
rect 2748 39076 2754 39110
rect 2788 39076 2794 39110
rect 2748 39029 2794 39076
rect 2844 39254 2890 39301
rect 2844 39220 2850 39254
rect 2884 39220 2890 39254
rect 2844 39182 2890 39220
rect 2844 39148 2850 39182
rect 2884 39148 2890 39182
rect 2844 39110 2890 39148
rect 2844 39076 2850 39110
rect 2884 39076 2890 39110
rect 2844 39029 2890 39076
rect 2940 39254 2986 39301
rect 2940 39220 2946 39254
rect 2980 39220 2986 39254
rect 2940 39182 2986 39220
rect 2940 39148 2946 39182
rect 2980 39148 2986 39182
rect 2940 39110 2986 39148
rect 2940 39076 2946 39110
rect 2980 39076 2986 39110
rect 2940 39029 2986 39076
rect 3036 39254 3082 39301
rect 3036 39220 3042 39254
rect 3076 39220 3082 39254
rect 3036 39182 3082 39220
rect 3036 39148 3042 39182
rect 3076 39148 3082 39182
rect 3036 39110 3082 39148
rect 3036 39076 3042 39110
rect 3076 39076 3082 39110
rect 3036 39029 3082 39076
rect 3132 39254 3178 39301
rect 3132 39220 3138 39254
rect 3172 39220 3178 39254
rect 3132 39182 3178 39220
rect 3132 39148 3138 39182
rect 3172 39148 3178 39182
rect 3132 39110 3178 39148
rect 3132 39076 3138 39110
rect 3172 39076 3178 39110
rect 3132 39029 3178 39076
rect 3228 39254 3274 39301
rect 3228 39220 3234 39254
rect 3268 39220 3274 39254
rect 3228 39182 3274 39220
rect 3228 39148 3234 39182
rect 3268 39148 3274 39182
rect 3228 39110 3274 39148
rect 3228 39076 3234 39110
rect 3268 39076 3274 39110
rect 3228 39029 3274 39076
rect 3324 39254 3370 39301
rect 3324 39220 3330 39254
rect 3364 39220 3370 39254
rect 3324 39182 3370 39220
rect 3324 39148 3330 39182
rect 3364 39148 3370 39182
rect 3324 39110 3370 39148
rect 3324 39076 3330 39110
rect 3364 39076 3370 39110
rect 3324 39029 3370 39076
rect 3420 39254 3466 39301
rect 3420 39220 3426 39254
rect 3460 39220 3466 39254
rect 3420 39182 3466 39220
rect 3420 39148 3426 39182
rect 3460 39148 3466 39182
rect 3420 39110 3466 39148
rect 3420 39076 3426 39110
rect 3460 39076 3466 39110
rect 3420 39029 3466 39076
rect 3534 39285 3580 39323
rect 3534 39251 3540 39285
rect 3574 39251 3580 39285
rect 3534 39213 3580 39251
rect 3534 39179 3540 39213
rect 3574 39179 3580 39213
rect 3534 39141 3580 39179
rect 3534 39107 3540 39141
rect 3574 39107 3580 39141
rect 3534 39069 3580 39107
rect 3534 39035 3540 39069
rect 3574 39035 3580 39069
rect 2101 38884 2316 38888
rect 313 38854 2316 38884
rect 313 38850 2141 38854
rect 313 38717 347 38850
rect 505 38717 539 38850
rect 697 38717 731 38850
rect 889 38717 923 38850
rect 1081 38717 1115 38850
rect 1273 38717 1307 38850
rect 1381 38724 1608 38747
rect 307 38682 353 38717
rect 307 38648 313 38682
rect 347 38648 353 38682
rect 307 38613 353 38648
rect 403 38682 449 38717
rect 403 38648 409 38682
rect 443 38648 449 38682
rect 403 38613 449 38648
rect 499 38682 545 38717
rect 499 38648 505 38682
rect 539 38648 545 38682
rect 499 38613 545 38648
rect 595 38682 641 38717
rect 595 38648 601 38682
rect 635 38648 641 38682
rect 595 38613 641 38648
rect 691 38682 737 38717
rect 691 38648 697 38682
rect 731 38648 737 38682
rect 691 38613 737 38648
rect 787 38682 833 38717
rect 787 38648 793 38682
rect 827 38648 833 38682
rect 787 38613 833 38648
rect 883 38682 929 38717
rect 883 38648 889 38682
rect 923 38648 929 38682
rect 883 38613 929 38648
rect 979 38682 1025 38717
rect 979 38648 985 38682
rect 1019 38648 1025 38682
rect 979 38613 1025 38648
rect 1075 38682 1121 38717
rect 1075 38648 1081 38682
rect 1115 38648 1121 38682
rect 1075 38613 1121 38648
rect 1171 38682 1217 38717
rect 1171 38648 1177 38682
rect 1211 38648 1217 38682
rect 1171 38613 1217 38648
rect 1267 38682 1313 38717
rect 1267 38648 1273 38682
rect 1307 38648 1313 38682
rect 1267 38613 1313 38648
rect 1381 38690 1387 38724
rect 1421 38690 1608 38724
rect 1381 38652 1608 38690
rect 1381 38618 1387 38652
rect 1421 38627 1608 38652
rect 1421 38618 1427 38627
rect 1560 38625 1608 38627
rect 1598 38623 1608 38625
rect 1720 38623 1730 38747
rect 297 38582 363 38585
rect 294 38530 304 38582
rect 356 38530 366 38582
rect 297 38525 363 38530
rect 409 38473 443 38613
rect 489 38582 555 38585
rect 485 38530 495 38582
rect 547 38530 557 38582
rect 489 38525 555 38530
rect 601 38473 635 38613
rect 681 38582 747 38585
rect 677 38530 687 38582
rect 739 38530 749 38582
rect 681 38525 747 38530
rect 793 38473 827 38613
rect 873 38582 939 38585
rect 869 38530 879 38582
rect 931 38530 941 38582
rect 873 38525 939 38530
rect 985 38473 1019 38613
rect 1065 38581 1131 38585
rect 1062 38529 1072 38581
rect 1124 38529 1134 38581
rect 1065 38525 1131 38529
rect 1177 38473 1211 38613
rect 1257 38581 1323 38585
rect 1254 38529 1264 38581
rect 1316 38529 1326 38581
rect 1381 38580 1427 38618
rect 1920 38585 1930 38587
rect 1381 38546 1387 38580
rect 1421 38546 1427 38580
rect 1257 38525 1323 38529
rect 129 38439 1211 38473
rect 1381 38403 1427 38546
rect 1458 38529 1468 38585
rect 1524 38531 1930 38585
rect 1986 38531 1996 38587
rect 1524 38529 1986 38531
rect 2282 38477 2316 38854
rect 2466 38888 2500 39029
rect 2658 38888 2692 39029
rect 2850 38888 2884 39029
rect 3042 38888 3076 39029
rect 3234 38888 3268 39029
rect 3426 38888 3460 39029
rect 3534 38991 3580 39035
rect 3803 39451 4885 39485
rect 3803 38888 3837 39451
rect 3968 39341 3978 39393
rect 4030 39341 4040 39393
rect 4083 39301 4117 39451
rect 4161 39341 4171 39393
rect 4223 39341 4233 39393
rect 4275 39301 4309 39451
rect 4352 39341 4362 39393
rect 4414 39341 4424 39393
rect 4467 39301 4501 39451
rect 4544 39341 4554 39393
rect 4606 39341 4616 39393
rect 4659 39301 4693 39451
rect 4736 39341 4746 39393
rect 4798 39341 4808 39393
rect 4851 39301 4885 39451
rect 4928 39341 4938 39393
rect 4990 39341 5000 39393
rect 5055 39357 5101 39562
rect 5055 39323 5061 39357
rect 5095 39323 5101 39357
rect 3981 39254 4027 39301
rect 3981 39220 3987 39254
rect 4021 39220 4027 39254
rect 3981 39182 4027 39220
rect 3981 39148 3987 39182
rect 4021 39148 4027 39182
rect 3981 39110 4027 39148
rect 3981 39076 3987 39110
rect 4021 39076 4027 39110
rect 3981 39029 4027 39076
rect 4077 39254 4123 39301
rect 4077 39220 4083 39254
rect 4117 39220 4123 39254
rect 4077 39182 4123 39220
rect 4077 39148 4083 39182
rect 4117 39148 4123 39182
rect 4077 39110 4123 39148
rect 4077 39076 4083 39110
rect 4117 39076 4123 39110
rect 4077 39029 4123 39076
rect 4173 39254 4219 39301
rect 4173 39220 4179 39254
rect 4213 39220 4219 39254
rect 4173 39182 4219 39220
rect 4173 39148 4179 39182
rect 4213 39148 4219 39182
rect 4173 39110 4219 39148
rect 4173 39076 4179 39110
rect 4213 39076 4219 39110
rect 4173 39029 4219 39076
rect 4269 39254 4315 39301
rect 4269 39220 4275 39254
rect 4309 39220 4315 39254
rect 4269 39182 4315 39220
rect 4269 39148 4275 39182
rect 4309 39148 4315 39182
rect 4269 39110 4315 39148
rect 4269 39076 4275 39110
rect 4309 39076 4315 39110
rect 4269 39029 4315 39076
rect 4365 39254 4411 39301
rect 4365 39220 4371 39254
rect 4405 39220 4411 39254
rect 4365 39182 4411 39220
rect 4365 39148 4371 39182
rect 4405 39148 4411 39182
rect 4365 39110 4411 39148
rect 4365 39076 4371 39110
rect 4405 39076 4411 39110
rect 4365 39029 4411 39076
rect 4461 39254 4507 39301
rect 4461 39220 4467 39254
rect 4501 39220 4507 39254
rect 4461 39182 4507 39220
rect 4461 39148 4467 39182
rect 4501 39148 4507 39182
rect 4461 39110 4507 39148
rect 4461 39076 4467 39110
rect 4501 39076 4507 39110
rect 4461 39029 4507 39076
rect 4557 39254 4603 39301
rect 4557 39220 4563 39254
rect 4597 39220 4603 39254
rect 4557 39182 4603 39220
rect 4557 39148 4563 39182
rect 4597 39148 4603 39182
rect 4557 39110 4603 39148
rect 4557 39076 4563 39110
rect 4597 39076 4603 39110
rect 4557 39029 4603 39076
rect 4653 39254 4699 39301
rect 4653 39220 4659 39254
rect 4693 39220 4699 39254
rect 4653 39182 4699 39220
rect 4653 39148 4659 39182
rect 4693 39148 4699 39182
rect 4653 39110 4699 39148
rect 4653 39076 4659 39110
rect 4693 39076 4699 39110
rect 4653 39029 4699 39076
rect 4749 39254 4795 39301
rect 4749 39220 4755 39254
rect 4789 39220 4795 39254
rect 4749 39182 4795 39220
rect 4749 39148 4755 39182
rect 4789 39148 4795 39182
rect 4749 39110 4795 39148
rect 4749 39076 4755 39110
rect 4789 39076 4795 39110
rect 4749 39029 4795 39076
rect 4845 39254 4891 39301
rect 4845 39220 4851 39254
rect 4885 39220 4891 39254
rect 4845 39182 4891 39220
rect 4845 39148 4851 39182
rect 4885 39148 4891 39182
rect 4845 39110 4891 39148
rect 4845 39076 4851 39110
rect 4885 39076 4891 39110
rect 4845 39029 4891 39076
rect 4941 39254 4987 39301
rect 4941 39220 4947 39254
rect 4981 39220 4987 39254
rect 4941 39182 4987 39220
rect 4941 39148 4947 39182
rect 4981 39148 4987 39182
rect 4941 39110 4987 39148
rect 4941 39076 4947 39110
rect 4981 39076 4987 39110
rect 4941 39029 4987 39076
rect 5055 39285 5101 39323
rect 5055 39251 5061 39285
rect 5095 39251 5101 39285
rect 5055 39213 5101 39251
rect 5055 39179 5061 39213
rect 5095 39182 5101 39213
rect 5274 39182 5550 39183
rect 5095 39179 5550 39182
rect 5055 39152 5550 39179
rect 5055 39141 5303 39152
rect 5055 39107 5061 39141
rect 5095 39118 5303 39141
rect 5337 39118 5395 39152
rect 5429 39118 5487 39152
rect 5521 39118 5550 39152
rect 5095 39107 5550 39118
rect 5055 39087 5550 39107
rect 5055 39069 5101 39087
rect 5055 39035 5061 39069
rect 5095 39035 5101 39069
rect 2466 38854 3837 38888
rect 2466 38721 2500 38854
rect 2658 38721 2692 38854
rect 2850 38721 2884 38854
rect 3042 38721 3076 38854
rect 3234 38721 3268 38854
rect 3426 38721 3460 38854
rect 3671 38764 3681 38816
rect 3733 38764 3743 38816
rect 3679 38763 3691 38764
rect 3725 38763 3737 38764
rect 3679 38757 3737 38763
rect 3534 38728 3580 38751
rect 2460 38686 2506 38721
rect 2460 38652 2466 38686
rect 2500 38652 2506 38686
rect 2460 38617 2506 38652
rect 2556 38686 2602 38721
rect 2556 38652 2562 38686
rect 2596 38652 2602 38686
rect 2556 38617 2602 38652
rect 2652 38686 2698 38721
rect 2652 38652 2658 38686
rect 2692 38652 2698 38686
rect 2652 38617 2698 38652
rect 2748 38686 2794 38721
rect 2748 38652 2754 38686
rect 2788 38652 2794 38686
rect 2748 38617 2794 38652
rect 2844 38686 2890 38721
rect 2844 38652 2850 38686
rect 2884 38652 2890 38686
rect 2844 38617 2890 38652
rect 2940 38686 2986 38721
rect 2940 38652 2946 38686
rect 2980 38652 2986 38686
rect 2940 38617 2986 38652
rect 3036 38686 3082 38721
rect 3036 38652 3042 38686
rect 3076 38652 3082 38686
rect 3036 38617 3082 38652
rect 3132 38686 3178 38721
rect 3132 38652 3138 38686
rect 3172 38652 3178 38686
rect 3132 38617 3178 38652
rect 3228 38686 3274 38721
rect 3228 38652 3234 38686
rect 3268 38652 3274 38686
rect 3228 38617 3274 38652
rect 3324 38686 3370 38721
rect 3324 38652 3330 38686
rect 3364 38652 3370 38686
rect 3324 38617 3370 38652
rect 3420 38686 3466 38721
rect 3420 38652 3426 38686
rect 3460 38652 3466 38686
rect 3420 38617 3466 38652
rect 3534 38694 3540 38728
rect 3574 38726 3580 38728
rect 3803 38726 3837 38854
rect 3574 38725 3680 38726
rect 3734 38725 3837 38726
rect 3574 38713 3687 38725
rect 3574 38694 3647 38713
rect 3534 38656 3647 38694
rect 3534 38622 3540 38656
rect 3574 38637 3647 38656
rect 3681 38637 3687 38713
rect 3574 38626 3687 38637
rect 3574 38622 3580 38626
rect 3641 38625 3687 38626
rect 3729 38713 3837 38725
rect 3987 38888 4021 39029
rect 4179 38888 4213 39029
rect 4371 38888 4405 39029
rect 4563 38888 4597 39029
rect 4755 38888 4789 39029
rect 4947 38888 4981 39029
rect 5055 38991 5101 39035
rect 5683 38942 5743 40195
rect 5177 38908 5743 38942
rect 5177 38888 5211 38908
rect 3987 38854 5211 38888
rect 3987 38721 4021 38854
rect 4179 38721 4213 38854
rect 4371 38721 4405 38854
rect 4563 38721 4597 38854
rect 4755 38721 4789 38854
rect 4947 38721 4981 38854
rect 5438 38850 5512 38851
rect 5326 38848 5400 38849
rect 5326 38796 5337 38848
rect 5389 38796 5400 38848
rect 5438 38798 5449 38850
rect 5501 38798 5512 38850
rect 5438 38797 5512 38798
rect 5326 38795 5400 38796
rect 5055 38728 5101 38751
rect 3729 38637 3735 38713
rect 3769 38637 3837 38713
rect 3729 38626 3837 38637
rect 3729 38625 3775 38626
rect 2450 38586 2516 38589
rect 2447 38534 2457 38586
rect 2509 38534 2519 38586
rect 2450 38529 2516 38534
rect 2562 38477 2596 38617
rect 2642 38586 2708 38589
rect 2638 38534 2648 38586
rect 2700 38534 2710 38586
rect 2642 38529 2708 38534
rect 2754 38477 2788 38617
rect 2834 38586 2900 38589
rect 2830 38534 2840 38586
rect 2892 38534 2902 38586
rect 2834 38529 2900 38534
rect 2946 38477 2980 38617
rect 3026 38586 3092 38589
rect 3022 38534 3032 38586
rect 3084 38534 3094 38586
rect 3026 38529 3092 38534
rect 3138 38477 3172 38617
rect 3218 38585 3284 38589
rect 3215 38533 3225 38585
rect 3277 38533 3287 38585
rect 3218 38529 3284 38533
rect 3330 38477 3364 38617
rect 3410 38585 3476 38589
rect 3407 38533 3417 38585
rect 3469 38533 3479 38585
rect 3534 38584 3580 38622
rect 3534 38550 3540 38584
rect 3574 38550 3580 38584
rect 3410 38529 3476 38533
rect 2282 38443 3364 38477
rect 3534 38367 3580 38550
rect 3803 38477 3837 38626
rect 3981 38686 4027 38721
rect 3981 38652 3987 38686
rect 4021 38652 4027 38686
rect 3981 38617 4027 38652
rect 4077 38686 4123 38721
rect 4077 38652 4083 38686
rect 4117 38652 4123 38686
rect 4077 38617 4123 38652
rect 4173 38686 4219 38721
rect 4173 38652 4179 38686
rect 4213 38652 4219 38686
rect 4173 38617 4219 38652
rect 4269 38686 4315 38721
rect 4269 38652 4275 38686
rect 4309 38652 4315 38686
rect 4269 38617 4315 38652
rect 4365 38686 4411 38721
rect 4365 38652 4371 38686
rect 4405 38652 4411 38686
rect 4365 38617 4411 38652
rect 4461 38686 4507 38721
rect 4461 38652 4467 38686
rect 4501 38652 4507 38686
rect 4461 38617 4507 38652
rect 4557 38686 4603 38721
rect 4557 38652 4563 38686
rect 4597 38652 4603 38686
rect 4557 38617 4603 38652
rect 4653 38686 4699 38721
rect 4653 38652 4659 38686
rect 4693 38652 4699 38686
rect 4653 38617 4699 38652
rect 4749 38686 4795 38721
rect 4749 38652 4755 38686
rect 4789 38652 4795 38686
rect 4749 38617 4795 38652
rect 4845 38686 4891 38721
rect 4845 38652 4851 38686
rect 4885 38652 4891 38686
rect 4845 38617 4891 38652
rect 4941 38686 4987 38721
rect 4941 38652 4947 38686
rect 4981 38652 4987 38686
rect 4941 38617 4987 38652
rect 5055 38694 5061 38728
rect 5095 38694 5101 38728
rect 5055 38656 5101 38694
rect 5055 38622 5061 38656
rect 5095 38639 5101 38656
rect 5095 38622 5550 38639
rect 3971 38586 4037 38589
rect 3968 38534 3978 38586
rect 4030 38534 4040 38586
rect 3971 38529 4037 38534
rect 4083 38477 4117 38617
rect 4163 38586 4229 38589
rect 4159 38534 4169 38586
rect 4221 38534 4231 38586
rect 4163 38529 4229 38534
rect 4275 38477 4309 38617
rect 4355 38586 4421 38589
rect 4351 38534 4361 38586
rect 4413 38534 4423 38586
rect 4355 38529 4421 38534
rect 4467 38477 4501 38617
rect 4547 38586 4613 38589
rect 4543 38534 4553 38586
rect 4605 38534 4615 38586
rect 4547 38529 4613 38534
rect 4659 38477 4693 38617
rect 4739 38585 4805 38589
rect 4736 38533 4746 38585
rect 4798 38533 4808 38585
rect 4739 38529 4805 38533
rect 4851 38477 4885 38617
rect 5055 38608 5550 38622
rect 4931 38585 4997 38589
rect 4928 38533 4938 38585
rect 4990 38533 5000 38585
rect 5055 38584 5303 38608
rect 5055 38550 5061 38584
rect 5095 38574 5303 38584
rect 5337 38574 5395 38608
rect 5429 38574 5487 38608
rect 5521 38574 5550 38608
rect 5095 38550 5550 38574
rect 5055 38543 5550 38550
rect 4931 38529 4997 38533
rect 3803 38443 4885 38477
rect 5055 38368 5101 38543
rect 129 38160 1211 38194
rect 129 37597 163 38160
rect 294 38050 304 38102
rect 356 38050 366 38102
rect 409 38010 443 38160
rect 487 38050 497 38102
rect 549 38050 559 38102
rect 601 38010 635 38160
rect 678 38050 688 38102
rect 740 38050 750 38102
rect 793 38010 827 38160
rect 870 38050 880 38102
rect 932 38050 942 38102
rect 985 38010 1019 38160
rect 1062 38050 1072 38102
rect 1124 38050 1134 38102
rect 1177 38010 1211 38160
rect 1254 38050 1264 38102
rect 1316 38050 1326 38102
rect 1381 38066 1427 38230
rect 2282 38164 3364 38198
rect 1381 38032 1387 38066
rect 1421 38032 1427 38066
rect 1512 38043 1522 38103
rect 1578 38043 1792 38103
rect 1852 38043 1862 38103
rect 307 37963 353 38010
rect 307 37929 313 37963
rect 347 37929 353 37963
rect 307 37891 353 37929
rect 307 37857 313 37891
rect 347 37857 353 37891
rect 307 37819 353 37857
rect 307 37785 313 37819
rect 347 37785 353 37819
rect 307 37738 353 37785
rect 403 37963 449 38010
rect 403 37929 409 37963
rect 443 37929 449 37963
rect 403 37891 449 37929
rect 403 37857 409 37891
rect 443 37857 449 37891
rect 403 37819 449 37857
rect 403 37785 409 37819
rect 443 37785 449 37819
rect 403 37738 449 37785
rect 499 37963 545 38010
rect 499 37929 505 37963
rect 539 37929 545 37963
rect 499 37891 545 37929
rect 499 37857 505 37891
rect 539 37857 545 37891
rect 499 37819 545 37857
rect 499 37785 505 37819
rect 539 37785 545 37819
rect 499 37738 545 37785
rect 595 37963 641 38010
rect 595 37929 601 37963
rect 635 37929 641 37963
rect 595 37891 641 37929
rect 595 37857 601 37891
rect 635 37857 641 37891
rect 595 37819 641 37857
rect 595 37785 601 37819
rect 635 37785 641 37819
rect 595 37738 641 37785
rect 691 37963 737 38010
rect 691 37929 697 37963
rect 731 37929 737 37963
rect 691 37891 737 37929
rect 691 37857 697 37891
rect 731 37857 737 37891
rect 691 37819 737 37857
rect 691 37785 697 37819
rect 731 37785 737 37819
rect 691 37738 737 37785
rect 787 37963 833 38010
rect 787 37929 793 37963
rect 827 37929 833 37963
rect 787 37891 833 37929
rect 787 37857 793 37891
rect 827 37857 833 37891
rect 787 37819 833 37857
rect 787 37785 793 37819
rect 827 37785 833 37819
rect 787 37738 833 37785
rect 883 37963 929 38010
rect 883 37929 889 37963
rect 923 37929 929 37963
rect 883 37891 929 37929
rect 883 37857 889 37891
rect 923 37857 929 37891
rect 883 37819 929 37857
rect 883 37785 889 37819
rect 923 37785 929 37819
rect 883 37738 929 37785
rect 979 37963 1025 38010
rect 979 37929 985 37963
rect 1019 37929 1025 37963
rect 979 37891 1025 37929
rect 979 37857 985 37891
rect 1019 37857 1025 37891
rect 979 37819 1025 37857
rect 979 37785 985 37819
rect 1019 37785 1025 37819
rect 979 37738 1025 37785
rect 1075 37963 1121 38010
rect 1075 37929 1081 37963
rect 1115 37929 1121 37963
rect 1075 37891 1121 37929
rect 1075 37857 1081 37891
rect 1115 37857 1121 37891
rect 1075 37819 1121 37857
rect 1075 37785 1081 37819
rect 1115 37785 1121 37819
rect 1075 37738 1121 37785
rect 1171 37963 1217 38010
rect 1171 37929 1177 37963
rect 1211 37929 1217 37963
rect 1171 37891 1217 37929
rect 1171 37857 1177 37891
rect 1211 37857 1217 37891
rect 1171 37819 1217 37857
rect 1171 37785 1177 37819
rect 1211 37785 1217 37819
rect 1171 37738 1217 37785
rect 1267 37963 1313 38010
rect 1267 37929 1273 37963
rect 1307 37929 1313 37963
rect 1267 37891 1313 37929
rect 1267 37857 1273 37891
rect 1307 37857 1313 37891
rect 1267 37819 1313 37857
rect 1267 37785 1273 37819
rect 1307 37785 1313 37819
rect 1267 37738 1313 37785
rect 1381 37994 1427 38032
rect 1381 37960 1387 37994
rect 1421 37960 1427 37994
rect 1381 37922 1427 37960
rect 1381 37888 1387 37922
rect 1421 37888 1427 37922
rect 1381 37850 1427 37888
rect 1381 37816 1387 37850
rect 1421 37816 1427 37850
rect 1381 37806 1427 37816
rect 1381 37804 2160 37806
rect 1381 37778 2056 37804
rect 1381 37753 1387 37778
rect 1380 37744 1387 37753
rect 1421 37744 2056 37778
rect 0 37563 163 37597
rect 129 37186 163 37563
rect 313 37597 347 37738
rect 505 37597 539 37738
rect 697 37597 731 37738
rect 889 37597 923 37738
rect 1081 37597 1115 37738
rect 1273 37597 1307 37738
rect 1380 37696 2056 37744
rect 2190 37696 2200 37804
rect 1380 37694 2160 37696
rect 2282 37601 2316 38164
rect 2447 38054 2457 38106
rect 2509 38054 2519 38106
rect 2562 38014 2596 38164
rect 2640 38054 2650 38106
rect 2702 38054 2712 38106
rect 2754 38014 2788 38164
rect 2831 38054 2841 38106
rect 2893 38054 2903 38106
rect 2946 38014 2980 38164
rect 3023 38054 3033 38106
rect 3085 38054 3095 38106
rect 3138 38014 3172 38164
rect 3215 38054 3225 38106
rect 3277 38054 3287 38106
rect 3330 38014 3364 38164
rect 3407 38054 3417 38106
rect 3469 38054 3479 38106
rect 3534 38070 3580 38278
rect 3534 38036 3540 38070
rect 3574 38036 3580 38070
rect 2460 37967 2506 38014
rect 2460 37933 2466 37967
rect 2500 37933 2506 37967
rect 2460 37895 2506 37933
rect 2460 37861 2466 37895
rect 2500 37861 2506 37895
rect 2460 37823 2506 37861
rect 2460 37789 2466 37823
rect 2500 37789 2506 37823
rect 2460 37742 2506 37789
rect 2556 37967 2602 38014
rect 2556 37933 2562 37967
rect 2596 37933 2602 37967
rect 2556 37895 2602 37933
rect 2556 37861 2562 37895
rect 2596 37861 2602 37895
rect 2556 37823 2602 37861
rect 2556 37789 2562 37823
rect 2596 37789 2602 37823
rect 2556 37742 2602 37789
rect 2652 37967 2698 38014
rect 2652 37933 2658 37967
rect 2692 37933 2698 37967
rect 2652 37895 2698 37933
rect 2652 37861 2658 37895
rect 2692 37861 2698 37895
rect 2652 37823 2698 37861
rect 2652 37789 2658 37823
rect 2692 37789 2698 37823
rect 2652 37742 2698 37789
rect 2748 37967 2794 38014
rect 2748 37933 2754 37967
rect 2788 37933 2794 37967
rect 2748 37895 2794 37933
rect 2748 37861 2754 37895
rect 2788 37861 2794 37895
rect 2748 37823 2794 37861
rect 2748 37789 2754 37823
rect 2788 37789 2794 37823
rect 2748 37742 2794 37789
rect 2844 37967 2890 38014
rect 2844 37933 2850 37967
rect 2884 37933 2890 37967
rect 2844 37895 2890 37933
rect 2844 37861 2850 37895
rect 2884 37861 2890 37895
rect 2844 37823 2890 37861
rect 2844 37789 2850 37823
rect 2884 37789 2890 37823
rect 2844 37742 2890 37789
rect 2940 37967 2986 38014
rect 2940 37933 2946 37967
rect 2980 37933 2986 37967
rect 2940 37895 2986 37933
rect 2940 37861 2946 37895
rect 2980 37861 2986 37895
rect 2940 37823 2986 37861
rect 2940 37789 2946 37823
rect 2980 37789 2986 37823
rect 2940 37742 2986 37789
rect 3036 37967 3082 38014
rect 3036 37933 3042 37967
rect 3076 37933 3082 37967
rect 3036 37895 3082 37933
rect 3036 37861 3042 37895
rect 3076 37861 3082 37895
rect 3036 37823 3082 37861
rect 3036 37789 3042 37823
rect 3076 37789 3082 37823
rect 3036 37742 3082 37789
rect 3132 37967 3178 38014
rect 3132 37933 3138 37967
rect 3172 37933 3178 37967
rect 3132 37895 3178 37933
rect 3132 37861 3138 37895
rect 3172 37861 3178 37895
rect 3132 37823 3178 37861
rect 3132 37789 3138 37823
rect 3172 37789 3178 37823
rect 3132 37742 3178 37789
rect 3228 37967 3274 38014
rect 3228 37933 3234 37967
rect 3268 37933 3274 37967
rect 3228 37895 3274 37933
rect 3228 37861 3234 37895
rect 3268 37861 3274 37895
rect 3228 37823 3274 37861
rect 3228 37789 3234 37823
rect 3268 37789 3274 37823
rect 3228 37742 3274 37789
rect 3324 37967 3370 38014
rect 3324 37933 3330 37967
rect 3364 37933 3370 37967
rect 3324 37895 3370 37933
rect 3324 37861 3330 37895
rect 3364 37861 3370 37895
rect 3324 37823 3370 37861
rect 3324 37789 3330 37823
rect 3364 37789 3370 37823
rect 3324 37742 3370 37789
rect 3420 37967 3466 38014
rect 3420 37933 3426 37967
rect 3460 37933 3466 37967
rect 3420 37895 3466 37933
rect 3420 37861 3426 37895
rect 3460 37861 3466 37895
rect 3420 37823 3466 37861
rect 3420 37789 3426 37823
rect 3460 37789 3466 37823
rect 3420 37742 3466 37789
rect 3534 37998 3580 38036
rect 3534 37964 3540 37998
rect 3574 37964 3580 37998
rect 3534 37926 3580 37964
rect 3534 37892 3540 37926
rect 3574 37892 3580 37926
rect 3534 37854 3580 37892
rect 3534 37820 3540 37854
rect 3574 37820 3580 37854
rect 3534 37782 3580 37820
rect 3534 37748 3540 37782
rect 3574 37748 3580 37782
rect 2101 37597 2316 37601
rect 313 37567 2316 37597
rect 313 37563 2141 37567
rect 313 37430 347 37563
rect 505 37430 539 37563
rect 697 37430 731 37563
rect 889 37430 923 37563
rect 1081 37430 1115 37563
rect 1273 37430 1307 37563
rect 1381 37437 1608 37460
rect 307 37395 353 37430
rect 307 37361 313 37395
rect 347 37361 353 37395
rect 307 37326 353 37361
rect 403 37395 449 37430
rect 403 37361 409 37395
rect 443 37361 449 37395
rect 403 37326 449 37361
rect 499 37395 545 37430
rect 499 37361 505 37395
rect 539 37361 545 37395
rect 499 37326 545 37361
rect 595 37395 641 37430
rect 595 37361 601 37395
rect 635 37361 641 37395
rect 595 37326 641 37361
rect 691 37395 737 37430
rect 691 37361 697 37395
rect 731 37361 737 37395
rect 691 37326 737 37361
rect 787 37395 833 37430
rect 787 37361 793 37395
rect 827 37361 833 37395
rect 787 37326 833 37361
rect 883 37395 929 37430
rect 883 37361 889 37395
rect 923 37361 929 37395
rect 883 37326 929 37361
rect 979 37395 1025 37430
rect 979 37361 985 37395
rect 1019 37361 1025 37395
rect 979 37326 1025 37361
rect 1075 37395 1121 37430
rect 1075 37361 1081 37395
rect 1115 37361 1121 37395
rect 1075 37326 1121 37361
rect 1171 37395 1217 37430
rect 1171 37361 1177 37395
rect 1211 37361 1217 37395
rect 1171 37326 1217 37361
rect 1267 37395 1313 37430
rect 1267 37361 1273 37395
rect 1307 37361 1313 37395
rect 1267 37326 1313 37361
rect 1381 37403 1387 37437
rect 1421 37403 1608 37437
rect 1381 37365 1608 37403
rect 1381 37331 1387 37365
rect 1421 37340 1608 37365
rect 1421 37331 1427 37340
rect 1560 37338 1608 37340
rect 1598 37336 1608 37338
rect 1720 37336 1730 37460
rect 297 37295 363 37298
rect 294 37243 304 37295
rect 356 37243 366 37295
rect 297 37238 363 37243
rect 409 37186 443 37326
rect 489 37295 555 37298
rect 485 37243 495 37295
rect 547 37243 557 37295
rect 489 37238 555 37243
rect 601 37186 635 37326
rect 681 37295 747 37298
rect 677 37243 687 37295
rect 739 37243 749 37295
rect 681 37238 747 37243
rect 793 37186 827 37326
rect 873 37295 939 37298
rect 869 37243 879 37295
rect 931 37243 941 37295
rect 873 37238 939 37243
rect 985 37186 1019 37326
rect 1065 37294 1131 37298
rect 1062 37242 1072 37294
rect 1124 37242 1134 37294
rect 1065 37238 1131 37242
rect 1177 37186 1211 37326
rect 1257 37294 1323 37298
rect 1254 37242 1264 37294
rect 1316 37242 1326 37294
rect 1381 37293 1427 37331
rect 1920 37298 1930 37300
rect 1381 37259 1387 37293
rect 1421 37259 1427 37293
rect 1257 37238 1323 37242
rect 129 37152 1211 37186
rect 1381 37116 1427 37259
rect 1458 37242 1468 37298
rect 1524 37244 1930 37298
rect 1986 37244 1996 37300
rect 1524 37242 1986 37244
rect 2282 37190 2316 37567
rect 2466 37601 2500 37742
rect 2658 37601 2692 37742
rect 2850 37601 2884 37742
rect 3042 37601 3076 37742
rect 3234 37601 3268 37742
rect 3426 37601 3460 37742
rect 3534 37704 3580 37748
rect 3803 38164 4885 38198
rect 3803 37601 3837 38164
rect 3968 38054 3978 38106
rect 4030 38054 4040 38106
rect 4083 38014 4117 38164
rect 4161 38054 4171 38106
rect 4223 38054 4233 38106
rect 4275 38014 4309 38164
rect 4352 38054 4362 38106
rect 4414 38054 4424 38106
rect 4467 38014 4501 38164
rect 4544 38054 4554 38106
rect 4606 38054 4616 38106
rect 4659 38014 4693 38164
rect 4736 38054 4746 38106
rect 4798 38054 4808 38106
rect 4851 38014 4885 38164
rect 4928 38054 4938 38106
rect 4990 38054 5000 38106
rect 5055 38070 5101 38275
rect 5055 38036 5061 38070
rect 5095 38036 5101 38070
rect 3981 37967 4027 38014
rect 3981 37933 3987 37967
rect 4021 37933 4027 37967
rect 3981 37895 4027 37933
rect 3981 37861 3987 37895
rect 4021 37861 4027 37895
rect 3981 37823 4027 37861
rect 3981 37789 3987 37823
rect 4021 37789 4027 37823
rect 3981 37742 4027 37789
rect 4077 37967 4123 38014
rect 4077 37933 4083 37967
rect 4117 37933 4123 37967
rect 4077 37895 4123 37933
rect 4077 37861 4083 37895
rect 4117 37861 4123 37895
rect 4077 37823 4123 37861
rect 4077 37789 4083 37823
rect 4117 37789 4123 37823
rect 4077 37742 4123 37789
rect 4173 37967 4219 38014
rect 4173 37933 4179 37967
rect 4213 37933 4219 37967
rect 4173 37895 4219 37933
rect 4173 37861 4179 37895
rect 4213 37861 4219 37895
rect 4173 37823 4219 37861
rect 4173 37789 4179 37823
rect 4213 37789 4219 37823
rect 4173 37742 4219 37789
rect 4269 37967 4315 38014
rect 4269 37933 4275 37967
rect 4309 37933 4315 37967
rect 4269 37895 4315 37933
rect 4269 37861 4275 37895
rect 4309 37861 4315 37895
rect 4269 37823 4315 37861
rect 4269 37789 4275 37823
rect 4309 37789 4315 37823
rect 4269 37742 4315 37789
rect 4365 37967 4411 38014
rect 4365 37933 4371 37967
rect 4405 37933 4411 37967
rect 4365 37895 4411 37933
rect 4365 37861 4371 37895
rect 4405 37861 4411 37895
rect 4365 37823 4411 37861
rect 4365 37789 4371 37823
rect 4405 37789 4411 37823
rect 4365 37742 4411 37789
rect 4461 37967 4507 38014
rect 4461 37933 4467 37967
rect 4501 37933 4507 37967
rect 4461 37895 4507 37933
rect 4461 37861 4467 37895
rect 4501 37861 4507 37895
rect 4461 37823 4507 37861
rect 4461 37789 4467 37823
rect 4501 37789 4507 37823
rect 4461 37742 4507 37789
rect 4557 37967 4603 38014
rect 4557 37933 4563 37967
rect 4597 37933 4603 37967
rect 4557 37895 4603 37933
rect 4557 37861 4563 37895
rect 4597 37861 4603 37895
rect 4557 37823 4603 37861
rect 4557 37789 4563 37823
rect 4597 37789 4603 37823
rect 4557 37742 4603 37789
rect 4653 37967 4699 38014
rect 4653 37933 4659 37967
rect 4693 37933 4699 37967
rect 4653 37895 4699 37933
rect 4653 37861 4659 37895
rect 4693 37861 4699 37895
rect 4653 37823 4699 37861
rect 4653 37789 4659 37823
rect 4693 37789 4699 37823
rect 4653 37742 4699 37789
rect 4749 37967 4795 38014
rect 4749 37933 4755 37967
rect 4789 37933 4795 37967
rect 4749 37895 4795 37933
rect 4749 37861 4755 37895
rect 4789 37861 4795 37895
rect 4749 37823 4795 37861
rect 4749 37789 4755 37823
rect 4789 37789 4795 37823
rect 4749 37742 4795 37789
rect 4845 37967 4891 38014
rect 4845 37933 4851 37967
rect 4885 37933 4891 37967
rect 4845 37895 4891 37933
rect 4845 37861 4851 37895
rect 4885 37861 4891 37895
rect 4845 37823 4891 37861
rect 4845 37789 4851 37823
rect 4885 37789 4891 37823
rect 4845 37742 4891 37789
rect 4941 37967 4987 38014
rect 4941 37933 4947 37967
rect 4981 37933 4987 37967
rect 4941 37895 4987 37933
rect 4941 37861 4947 37895
rect 4981 37861 4987 37895
rect 4941 37823 4987 37861
rect 4941 37789 4947 37823
rect 4981 37789 4987 37823
rect 4941 37742 4987 37789
rect 5055 37998 5101 38036
rect 5055 37964 5061 37998
rect 5095 37964 5101 37998
rect 5055 37926 5101 37964
rect 5055 37892 5061 37926
rect 5095 37895 5101 37926
rect 5274 37895 5550 37896
rect 5095 37892 5550 37895
rect 5055 37865 5550 37892
rect 5055 37854 5303 37865
rect 5055 37820 5061 37854
rect 5095 37831 5303 37854
rect 5337 37831 5395 37865
rect 5429 37831 5487 37865
rect 5521 37831 5550 37865
rect 5095 37820 5550 37831
rect 5055 37800 5550 37820
rect 5055 37782 5101 37800
rect 5055 37748 5061 37782
rect 5095 37748 5101 37782
rect 2466 37567 3837 37601
rect 2466 37434 2500 37567
rect 2658 37434 2692 37567
rect 2850 37434 2884 37567
rect 3042 37434 3076 37567
rect 3234 37434 3268 37567
rect 3426 37434 3460 37567
rect 3671 37477 3681 37529
rect 3733 37477 3743 37529
rect 3679 37476 3691 37477
rect 3725 37476 3737 37477
rect 3679 37470 3737 37476
rect 3534 37441 3580 37464
rect 2460 37399 2506 37434
rect 2460 37365 2466 37399
rect 2500 37365 2506 37399
rect 2460 37330 2506 37365
rect 2556 37399 2602 37434
rect 2556 37365 2562 37399
rect 2596 37365 2602 37399
rect 2556 37330 2602 37365
rect 2652 37399 2698 37434
rect 2652 37365 2658 37399
rect 2692 37365 2698 37399
rect 2652 37330 2698 37365
rect 2748 37399 2794 37434
rect 2748 37365 2754 37399
rect 2788 37365 2794 37399
rect 2748 37330 2794 37365
rect 2844 37399 2890 37434
rect 2844 37365 2850 37399
rect 2884 37365 2890 37399
rect 2844 37330 2890 37365
rect 2940 37399 2986 37434
rect 2940 37365 2946 37399
rect 2980 37365 2986 37399
rect 2940 37330 2986 37365
rect 3036 37399 3082 37434
rect 3036 37365 3042 37399
rect 3076 37365 3082 37399
rect 3036 37330 3082 37365
rect 3132 37399 3178 37434
rect 3132 37365 3138 37399
rect 3172 37365 3178 37399
rect 3132 37330 3178 37365
rect 3228 37399 3274 37434
rect 3228 37365 3234 37399
rect 3268 37365 3274 37399
rect 3228 37330 3274 37365
rect 3324 37399 3370 37434
rect 3324 37365 3330 37399
rect 3364 37365 3370 37399
rect 3324 37330 3370 37365
rect 3420 37399 3466 37434
rect 3420 37365 3426 37399
rect 3460 37365 3466 37399
rect 3420 37330 3466 37365
rect 3534 37407 3540 37441
rect 3574 37439 3580 37441
rect 3803 37439 3837 37567
rect 3574 37438 3680 37439
rect 3734 37438 3837 37439
rect 3574 37426 3687 37438
rect 3574 37407 3647 37426
rect 3534 37369 3647 37407
rect 3534 37335 3540 37369
rect 3574 37350 3647 37369
rect 3681 37350 3687 37426
rect 3574 37339 3687 37350
rect 3574 37335 3580 37339
rect 3641 37338 3687 37339
rect 3729 37426 3837 37438
rect 3987 37601 4021 37742
rect 4179 37601 4213 37742
rect 4371 37601 4405 37742
rect 4563 37601 4597 37742
rect 4755 37601 4789 37742
rect 4947 37601 4981 37742
rect 5055 37704 5101 37748
rect 5683 37655 5743 38908
rect 5177 37621 5743 37655
rect 5177 37601 5211 37621
rect 3987 37567 5211 37601
rect 3987 37434 4021 37567
rect 4179 37434 4213 37567
rect 4371 37434 4405 37567
rect 4563 37434 4597 37567
rect 4755 37434 4789 37567
rect 4947 37434 4981 37567
rect 5438 37563 5512 37564
rect 5326 37561 5400 37562
rect 5326 37509 5337 37561
rect 5389 37509 5400 37561
rect 5438 37511 5449 37563
rect 5501 37511 5512 37563
rect 5438 37510 5512 37511
rect 5326 37508 5400 37509
rect 5055 37441 5101 37464
rect 3729 37350 3735 37426
rect 3769 37350 3837 37426
rect 3729 37339 3837 37350
rect 3729 37338 3775 37339
rect 2450 37299 2516 37302
rect 2447 37247 2457 37299
rect 2509 37247 2519 37299
rect 2450 37242 2516 37247
rect 2562 37190 2596 37330
rect 2642 37299 2708 37302
rect 2638 37247 2648 37299
rect 2700 37247 2710 37299
rect 2642 37242 2708 37247
rect 2754 37190 2788 37330
rect 2834 37299 2900 37302
rect 2830 37247 2840 37299
rect 2892 37247 2902 37299
rect 2834 37242 2900 37247
rect 2946 37190 2980 37330
rect 3026 37299 3092 37302
rect 3022 37247 3032 37299
rect 3084 37247 3094 37299
rect 3026 37242 3092 37247
rect 3138 37190 3172 37330
rect 3218 37298 3284 37302
rect 3215 37246 3225 37298
rect 3277 37246 3287 37298
rect 3218 37242 3284 37246
rect 3330 37190 3364 37330
rect 3410 37298 3476 37302
rect 3407 37246 3417 37298
rect 3469 37246 3479 37298
rect 3534 37297 3580 37335
rect 3534 37263 3540 37297
rect 3574 37263 3580 37297
rect 3410 37242 3476 37246
rect 2282 37156 3364 37190
rect 3534 37080 3580 37263
rect 3803 37190 3837 37339
rect 3981 37399 4027 37434
rect 3981 37365 3987 37399
rect 4021 37365 4027 37399
rect 3981 37330 4027 37365
rect 4077 37399 4123 37434
rect 4077 37365 4083 37399
rect 4117 37365 4123 37399
rect 4077 37330 4123 37365
rect 4173 37399 4219 37434
rect 4173 37365 4179 37399
rect 4213 37365 4219 37399
rect 4173 37330 4219 37365
rect 4269 37399 4315 37434
rect 4269 37365 4275 37399
rect 4309 37365 4315 37399
rect 4269 37330 4315 37365
rect 4365 37399 4411 37434
rect 4365 37365 4371 37399
rect 4405 37365 4411 37399
rect 4365 37330 4411 37365
rect 4461 37399 4507 37434
rect 4461 37365 4467 37399
rect 4501 37365 4507 37399
rect 4461 37330 4507 37365
rect 4557 37399 4603 37434
rect 4557 37365 4563 37399
rect 4597 37365 4603 37399
rect 4557 37330 4603 37365
rect 4653 37399 4699 37434
rect 4653 37365 4659 37399
rect 4693 37365 4699 37399
rect 4653 37330 4699 37365
rect 4749 37399 4795 37434
rect 4749 37365 4755 37399
rect 4789 37365 4795 37399
rect 4749 37330 4795 37365
rect 4845 37399 4891 37434
rect 4845 37365 4851 37399
rect 4885 37365 4891 37399
rect 4845 37330 4891 37365
rect 4941 37399 4987 37434
rect 4941 37365 4947 37399
rect 4981 37365 4987 37399
rect 4941 37330 4987 37365
rect 5055 37407 5061 37441
rect 5095 37407 5101 37441
rect 5055 37369 5101 37407
rect 5055 37335 5061 37369
rect 5095 37352 5101 37369
rect 5095 37335 5550 37352
rect 3971 37299 4037 37302
rect 3968 37247 3978 37299
rect 4030 37247 4040 37299
rect 3971 37242 4037 37247
rect 4083 37190 4117 37330
rect 4163 37299 4229 37302
rect 4159 37247 4169 37299
rect 4221 37247 4231 37299
rect 4163 37242 4229 37247
rect 4275 37190 4309 37330
rect 4355 37299 4421 37302
rect 4351 37247 4361 37299
rect 4413 37247 4423 37299
rect 4355 37242 4421 37247
rect 4467 37190 4501 37330
rect 4547 37299 4613 37302
rect 4543 37247 4553 37299
rect 4605 37247 4615 37299
rect 4547 37242 4613 37247
rect 4659 37190 4693 37330
rect 4739 37298 4805 37302
rect 4736 37246 4746 37298
rect 4798 37246 4808 37298
rect 4739 37242 4805 37246
rect 4851 37190 4885 37330
rect 5055 37321 5550 37335
rect 4931 37298 4997 37302
rect 4928 37246 4938 37298
rect 4990 37246 5000 37298
rect 5055 37297 5303 37321
rect 5055 37263 5061 37297
rect 5095 37287 5303 37297
rect 5337 37287 5395 37321
rect 5429 37287 5487 37321
rect 5521 37287 5550 37321
rect 5095 37263 5550 37287
rect 5055 37256 5550 37263
rect 4931 37242 4997 37246
rect 3803 37156 4885 37190
rect 5055 37081 5101 37256
rect 129 36873 1211 36907
rect 129 36310 163 36873
rect 294 36763 304 36815
rect 356 36763 366 36815
rect 409 36723 443 36873
rect 487 36763 497 36815
rect 549 36763 559 36815
rect 601 36723 635 36873
rect 678 36763 688 36815
rect 740 36763 750 36815
rect 793 36723 827 36873
rect 870 36763 880 36815
rect 932 36763 942 36815
rect 985 36723 1019 36873
rect 1062 36763 1072 36815
rect 1124 36763 1134 36815
rect 1177 36723 1211 36873
rect 1254 36763 1264 36815
rect 1316 36763 1326 36815
rect 1381 36779 1427 36943
rect 2282 36877 3364 36911
rect 1381 36745 1387 36779
rect 1421 36745 1427 36779
rect 1512 36756 1522 36816
rect 1578 36756 1792 36816
rect 1852 36756 1862 36816
rect 307 36676 353 36723
rect 307 36642 313 36676
rect 347 36642 353 36676
rect 307 36604 353 36642
rect 307 36570 313 36604
rect 347 36570 353 36604
rect 307 36532 353 36570
rect 307 36498 313 36532
rect 347 36498 353 36532
rect 307 36451 353 36498
rect 403 36676 449 36723
rect 403 36642 409 36676
rect 443 36642 449 36676
rect 403 36604 449 36642
rect 403 36570 409 36604
rect 443 36570 449 36604
rect 403 36532 449 36570
rect 403 36498 409 36532
rect 443 36498 449 36532
rect 403 36451 449 36498
rect 499 36676 545 36723
rect 499 36642 505 36676
rect 539 36642 545 36676
rect 499 36604 545 36642
rect 499 36570 505 36604
rect 539 36570 545 36604
rect 499 36532 545 36570
rect 499 36498 505 36532
rect 539 36498 545 36532
rect 499 36451 545 36498
rect 595 36676 641 36723
rect 595 36642 601 36676
rect 635 36642 641 36676
rect 595 36604 641 36642
rect 595 36570 601 36604
rect 635 36570 641 36604
rect 595 36532 641 36570
rect 595 36498 601 36532
rect 635 36498 641 36532
rect 595 36451 641 36498
rect 691 36676 737 36723
rect 691 36642 697 36676
rect 731 36642 737 36676
rect 691 36604 737 36642
rect 691 36570 697 36604
rect 731 36570 737 36604
rect 691 36532 737 36570
rect 691 36498 697 36532
rect 731 36498 737 36532
rect 691 36451 737 36498
rect 787 36676 833 36723
rect 787 36642 793 36676
rect 827 36642 833 36676
rect 787 36604 833 36642
rect 787 36570 793 36604
rect 827 36570 833 36604
rect 787 36532 833 36570
rect 787 36498 793 36532
rect 827 36498 833 36532
rect 787 36451 833 36498
rect 883 36676 929 36723
rect 883 36642 889 36676
rect 923 36642 929 36676
rect 883 36604 929 36642
rect 883 36570 889 36604
rect 923 36570 929 36604
rect 883 36532 929 36570
rect 883 36498 889 36532
rect 923 36498 929 36532
rect 883 36451 929 36498
rect 979 36676 1025 36723
rect 979 36642 985 36676
rect 1019 36642 1025 36676
rect 979 36604 1025 36642
rect 979 36570 985 36604
rect 1019 36570 1025 36604
rect 979 36532 1025 36570
rect 979 36498 985 36532
rect 1019 36498 1025 36532
rect 979 36451 1025 36498
rect 1075 36676 1121 36723
rect 1075 36642 1081 36676
rect 1115 36642 1121 36676
rect 1075 36604 1121 36642
rect 1075 36570 1081 36604
rect 1115 36570 1121 36604
rect 1075 36532 1121 36570
rect 1075 36498 1081 36532
rect 1115 36498 1121 36532
rect 1075 36451 1121 36498
rect 1171 36676 1217 36723
rect 1171 36642 1177 36676
rect 1211 36642 1217 36676
rect 1171 36604 1217 36642
rect 1171 36570 1177 36604
rect 1211 36570 1217 36604
rect 1171 36532 1217 36570
rect 1171 36498 1177 36532
rect 1211 36498 1217 36532
rect 1171 36451 1217 36498
rect 1267 36676 1313 36723
rect 1267 36642 1273 36676
rect 1307 36642 1313 36676
rect 1267 36604 1313 36642
rect 1267 36570 1273 36604
rect 1307 36570 1313 36604
rect 1267 36532 1313 36570
rect 1267 36498 1273 36532
rect 1307 36498 1313 36532
rect 1267 36451 1313 36498
rect 1381 36707 1427 36745
rect 1381 36673 1387 36707
rect 1421 36673 1427 36707
rect 1381 36635 1427 36673
rect 1381 36601 1387 36635
rect 1421 36601 1427 36635
rect 1381 36563 1427 36601
rect 1381 36529 1387 36563
rect 1421 36529 1427 36563
rect 1381 36519 1427 36529
rect 1381 36517 2160 36519
rect 1381 36491 2056 36517
rect 1381 36466 1387 36491
rect 1380 36457 1387 36466
rect 1421 36457 2056 36491
rect 0 36276 163 36310
rect 129 35899 163 36276
rect 313 36310 347 36451
rect 505 36310 539 36451
rect 697 36310 731 36451
rect 889 36310 923 36451
rect 1081 36310 1115 36451
rect 1273 36310 1307 36451
rect 1380 36409 2056 36457
rect 2190 36409 2200 36517
rect 1380 36407 2160 36409
rect 2282 36314 2316 36877
rect 2447 36767 2457 36819
rect 2509 36767 2519 36819
rect 2562 36727 2596 36877
rect 2640 36767 2650 36819
rect 2702 36767 2712 36819
rect 2754 36727 2788 36877
rect 2831 36767 2841 36819
rect 2893 36767 2903 36819
rect 2946 36727 2980 36877
rect 3023 36767 3033 36819
rect 3085 36767 3095 36819
rect 3138 36727 3172 36877
rect 3215 36767 3225 36819
rect 3277 36767 3287 36819
rect 3330 36727 3364 36877
rect 3407 36767 3417 36819
rect 3469 36767 3479 36819
rect 3534 36783 3580 36991
rect 3534 36749 3540 36783
rect 3574 36749 3580 36783
rect 2460 36680 2506 36727
rect 2460 36646 2466 36680
rect 2500 36646 2506 36680
rect 2460 36608 2506 36646
rect 2460 36574 2466 36608
rect 2500 36574 2506 36608
rect 2460 36536 2506 36574
rect 2460 36502 2466 36536
rect 2500 36502 2506 36536
rect 2460 36455 2506 36502
rect 2556 36680 2602 36727
rect 2556 36646 2562 36680
rect 2596 36646 2602 36680
rect 2556 36608 2602 36646
rect 2556 36574 2562 36608
rect 2596 36574 2602 36608
rect 2556 36536 2602 36574
rect 2556 36502 2562 36536
rect 2596 36502 2602 36536
rect 2556 36455 2602 36502
rect 2652 36680 2698 36727
rect 2652 36646 2658 36680
rect 2692 36646 2698 36680
rect 2652 36608 2698 36646
rect 2652 36574 2658 36608
rect 2692 36574 2698 36608
rect 2652 36536 2698 36574
rect 2652 36502 2658 36536
rect 2692 36502 2698 36536
rect 2652 36455 2698 36502
rect 2748 36680 2794 36727
rect 2748 36646 2754 36680
rect 2788 36646 2794 36680
rect 2748 36608 2794 36646
rect 2748 36574 2754 36608
rect 2788 36574 2794 36608
rect 2748 36536 2794 36574
rect 2748 36502 2754 36536
rect 2788 36502 2794 36536
rect 2748 36455 2794 36502
rect 2844 36680 2890 36727
rect 2844 36646 2850 36680
rect 2884 36646 2890 36680
rect 2844 36608 2890 36646
rect 2844 36574 2850 36608
rect 2884 36574 2890 36608
rect 2844 36536 2890 36574
rect 2844 36502 2850 36536
rect 2884 36502 2890 36536
rect 2844 36455 2890 36502
rect 2940 36680 2986 36727
rect 2940 36646 2946 36680
rect 2980 36646 2986 36680
rect 2940 36608 2986 36646
rect 2940 36574 2946 36608
rect 2980 36574 2986 36608
rect 2940 36536 2986 36574
rect 2940 36502 2946 36536
rect 2980 36502 2986 36536
rect 2940 36455 2986 36502
rect 3036 36680 3082 36727
rect 3036 36646 3042 36680
rect 3076 36646 3082 36680
rect 3036 36608 3082 36646
rect 3036 36574 3042 36608
rect 3076 36574 3082 36608
rect 3036 36536 3082 36574
rect 3036 36502 3042 36536
rect 3076 36502 3082 36536
rect 3036 36455 3082 36502
rect 3132 36680 3178 36727
rect 3132 36646 3138 36680
rect 3172 36646 3178 36680
rect 3132 36608 3178 36646
rect 3132 36574 3138 36608
rect 3172 36574 3178 36608
rect 3132 36536 3178 36574
rect 3132 36502 3138 36536
rect 3172 36502 3178 36536
rect 3132 36455 3178 36502
rect 3228 36680 3274 36727
rect 3228 36646 3234 36680
rect 3268 36646 3274 36680
rect 3228 36608 3274 36646
rect 3228 36574 3234 36608
rect 3268 36574 3274 36608
rect 3228 36536 3274 36574
rect 3228 36502 3234 36536
rect 3268 36502 3274 36536
rect 3228 36455 3274 36502
rect 3324 36680 3370 36727
rect 3324 36646 3330 36680
rect 3364 36646 3370 36680
rect 3324 36608 3370 36646
rect 3324 36574 3330 36608
rect 3364 36574 3370 36608
rect 3324 36536 3370 36574
rect 3324 36502 3330 36536
rect 3364 36502 3370 36536
rect 3324 36455 3370 36502
rect 3420 36680 3466 36727
rect 3420 36646 3426 36680
rect 3460 36646 3466 36680
rect 3420 36608 3466 36646
rect 3420 36574 3426 36608
rect 3460 36574 3466 36608
rect 3420 36536 3466 36574
rect 3420 36502 3426 36536
rect 3460 36502 3466 36536
rect 3420 36455 3466 36502
rect 3534 36711 3580 36749
rect 3534 36677 3540 36711
rect 3574 36677 3580 36711
rect 3534 36639 3580 36677
rect 3534 36605 3540 36639
rect 3574 36605 3580 36639
rect 3534 36567 3580 36605
rect 3534 36533 3540 36567
rect 3574 36533 3580 36567
rect 3534 36495 3580 36533
rect 3534 36461 3540 36495
rect 3574 36461 3580 36495
rect 2101 36310 2316 36314
rect 313 36280 2316 36310
rect 313 36276 2141 36280
rect 313 36143 347 36276
rect 505 36143 539 36276
rect 697 36143 731 36276
rect 889 36143 923 36276
rect 1081 36143 1115 36276
rect 1273 36143 1307 36276
rect 1381 36150 1608 36173
rect 307 36108 353 36143
rect 307 36074 313 36108
rect 347 36074 353 36108
rect 307 36039 353 36074
rect 403 36108 449 36143
rect 403 36074 409 36108
rect 443 36074 449 36108
rect 403 36039 449 36074
rect 499 36108 545 36143
rect 499 36074 505 36108
rect 539 36074 545 36108
rect 499 36039 545 36074
rect 595 36108 641 36143
rect 595 36074 601 36108
rect 635 36074 641 36108
rect 595 36039 641 36074
rect 691 36108 737 36143
rect 691 36074 697 36108
rect 731 36074 737 36108
rect 691 36039 737 36074
rect 787 36108 833 36143
rect 787 36074 793 36108
rect 827 36074 833 36108
rect 787 36039 833 36074
rect 883 36108 929 36143
rect 883 36074 889 36108
rect 923 36074 929 36108
rect 883 36039 929 36074
rect 979 36108 1025 36143
rect 979 36074 985 36108
rect 1019 36074 1025 36108
rect 979 36039 1025 36074
rect 1075 36108 1121 36143
rect 1075 36074 1081 36108
rect 1115 36074 1121 36108
rect 1075 36039 1121 36074
rect 1171 36108 1217 36143
rect 1171 36074 1177 36108
rect 1211 36074 1217 36108
rect 1171 36039 1217 36074
rect 1267 36108 1313 36143
rect 1267 36074 1273 36108
rect 1307 36074 1313 36108
rect 1267 36039 1313 36074
rect 1381 36116 1387 36150
rect 1421 36116 1608 36150
rect 1381 36078 1608 36116
rect 1381 36044 1387 36078
rect 1421 36053 1608 36078
rect 1421 36044 1427 36053
rect 1560 36051 1608 36053
rect 1598 36049 1608 36051
rect 1720 36049 1730 36173
rect 297 36008 363 36011
rect 294 35956 304 36008
rect 356 35956 366 36008
rect 297 35951 363 35956
rect 409 35899 443 36039
rect 489 36008 555 36011
rect 485 35956 495 36008
rect 547 35956 557 36008
rect 489 35951 555 35956
rect 601 35899 635 36039
rect 681 36008 747 36011
rect 677 35956 687 36008
rect 739 35956 749 36008
rect 681 35951 747 35956
rect 793 35899 827 36039
rect 873 36008 939 36011
rect 869 35956 879 36008
rect 931 35956 941 36008
rect 873 35951 939 35956
rect 985 35899 1019 36039
rect 1065 36007 1131 36011
rect 1062 35955 1072 36007
rect 1124 35955 1134 36007
rect 1065 35951 1131 35955
rect 1177 35899 1211 36039
rect 1257 36007 1323 36011
rect 1254 35955 1264 36007
rect 1316 35955 1326 36007
rect 1381 36006 1427 36044
rect 1920 36011 1930 36013
rect 1381 35972 1387 36006
rect 1421 35972 1427 36006
rect 1257 35951 1323 35955
rect 129 35865 1211 35899
rect 1381 35829 1427 35972
rect 1458 35955 1468 36011
rect 1524 35957 1930 36011
rect 1986 35957 1996 36013
rect 1524 35955 1986 35957
rect 2282 35903 2316 36280
rect 2466 36314 2500 36455
rect 2658 36314 2692 36455
rect 2850 36314 2884 36455
rect 3042 36314 3076 36455
rect 3234 36314 3268 36455
rect 3426 36314 3460 36455
rect 3534 36417 3580 36461
rect 3803 36877 4885 36911
rect 3803 36314 3837 36877
rect 3968 36767 3978 36819
rect 4030 36767 4040 36819
rect 4083 36727 4117 36877
rect 4161 36767 4171 36819
rect 4223 36767 4233 36819
rect 4275 36727 4309 36877
rect 4352 36767 4362 36819
rect 4414 36767 4424 36819
rect 4467 36727 4501 36877
rect 4544 36767 4554 36819
rect 4606 36767 4616 36819
rect 4659 36727 4693 36877
rect 4736 36767 4746 36819
rect 4798 36767 4808 36819
rect 4851 36727 4885 36877
rect 4928 36767 4938 36819
rect 4990 36767 5000 36819
rect 5055 36783 5101 36988
rect 5055 36749 5061 36783
rect 5095 36749 5101 36783
rect 3981 36680 4027 36727
rect 3981 36646 3987 36680
rect 4021 36646 4027 36680
rect 3981 36608 4027 36646
rect 3981 36574 3987 36608
rect 4021 36574 4027 36608
rect 3981 36536 4027 36574
rect 3981 36502 3987 36536
rect 4021 36502 4027 36536
rect 3981 36455 4027 36502
rect 4077 36680 4123 36727
rect 4077 36646 4083 36680
rect 4117 36646 4123 36680
rect 4077 36608 4123 36646
rect 4077 36574 4083 36608
rect 4117 36574 4123 36608
rect 4077 36536 4123 36574
rect 4077 36502 4083 36536
rect 4117 36502 4123 36536
rect 4077 36455 4123 36502
rect 4173 36680 4219 36727
rect 4173 36646 4179 36680
rect 4213 36646 4219 36680
rect 4173 36608 4219 36646
rect 4173 36574 4179 36608
rect 4213 36574 4219 36608
rect 4173 36536 4219 36574
rect 4173 36502 4179 36536
rect 4213 36502 4219 36536
rect 4173 36455 4219 36502
rect 4269 36680 4315 36727
rect 4269 36646 4275 36680
rect 4309 36646 4315 36680
rect 4269 36608 4315 36646
rect 4269 36574 4275 36608
rect 4309 36574 4315 36608
rect 4269 36536 4315 36574
rect 4269 36502 4275 36536
rect 4309 36502 4315 36536
rect 4269 36455 4315 36502
rect 4365 36680 4411 36727
rect 4365 36646 4371 36680
rect 4405 36646 4411 36680
rect 4365 36608 4411 36646
rect 4365 36574 4371 36608
rect 4405 36574 4411 36608
rect 4365 36536 4411 36574
rect 4365 36502 4371 36536
rect 4405 36502 4411 36536
rect 4365 36455 4411 36502
rect 4461 36680 4507 36727
rect 4461 36646 4467 36680
rect 4501 36646 4507 36680
rect 4461 36608 4507 36646
rect 4461 36574 4467 36608
rect 4501 36574 4507 36608
rect 4461 36536 4507 36574
rect 4461 36502 4467 36536
rect 4501 36502 4507 36536
rect 4461 36455 4507 36502
rect 4557 36680 4603 36727
rect 4557 36646 4563 36680
rect 4597 36646 4603 36680
rect 4557 36608 4603 36646
rect 4557 36574 4563 36608
rect 4597 36574 4603 36608
rect 4557 36536 4603 36574
rect 4557 36502 4563 36536
rect 4597 36502 4603 36536
rect 4557 36455 4603 36502
rect 4653 36680 4699 36727
rect 4653 36646 4659 36680
rect 4693 36646 4699 36680
rect 4653 36608 4699 36646
rect 4653 36574 4659 36608
rect 4693 36574 4699 36608
rect 4653 36536 4699 36574
rect 4653 36502 4659 36536
rect 4693 36502 4699 36536
rect 4653 36455 4699 36502
rect 4749 36680 4795 36727
rect 4749 36646 4755 36680
rect 4789 36646 4795 36680
rect 4749 36608 4795 36646
rect 4749 36574 4755 36608
rect 4789 36574 4795 36608
rect 4749 36536 4795 36574
rect 4749 36502 4755 36536
rect 4789 36502 4795 36536
rect 4749 36455 4795 36502
rect 4845 36680 4891 36727
rect 4845 36646 4851 36680
rect 4885 36646 4891 36680
rect 4845 36608 4891 36646
rect 4845 36574 4851 36608
rect 4885 36574 4891 36608
rect 4845 36536 4891 36574
rect 4845 36502 4851 36536
rect 4885 36502 4891 36536
rect 4845 36455 4891 36502
rect 4941 36680 4987 36727
rect 4941 36646 4947 36680
rect 4981 36646 4987 36680
rect 4941 36608 4987 36646
rect 4941 36574 4947 36608
rect 4981 36574 4987 36608
rect 4941 36536 4987 36574
rect 4941 36502 4947 36536
rect 4981 36502 4987 36536
rect 4941 36455 4987 36502
rect 5055 36711 5101 36749
rect 5055 36677 5061 36711
rect 5095 36677 5101 36711
rect 5055 36639 5101 36677
rect 5055 36605 5061 36639
rect 5095 36608 5101 36639
rect 5274 36608 5550 36609
rect 5095 36605 5550 36608
rect 5055 36578 5550 36605
rect 5055 36567 5303 36578
rect 5055 36533 5061 36567
rect 5095 36544 5303 36567
rect 5337 36544 5395 36578
rect 5429 36544 5487 36578
rect 5521 36544 5550 36578
rect 5095 36533 5550 36544
rect 5055 36513 5550 36533
rect 5055 36495 5101 36513
rect 5055 36461 5061 36495
rect 5095 36461 5101 36495
rect 2466 36280 3837 36314
rect 2466 36147 2500 36280
rect 2658 36147 2692 36280
rect 2850 36147 2884 36280
rect 3042 36147 3076 36280
rect 3234 36147 3268 36280
rect 3426 36147 3460 36280
rect 3671 36190 3681 36242
rect 3733 36190 3743 36242
rect 3679 36189 3691 36190
rect 3725 36189 3737 36190
rect 3679 36183 3737 36189
rect 3534 36154 3580 36177
rect 2460 36112 2506 36147
rect 2460 36078 2466 36112
rect 2500 36078 2506 36112
rect 2460 36043 2506 36078
rect 2556 36112 2602 36147
rect 2556 36078 2562 36112
rect 2596 36078 2602 36112
rect 2556 36043 2602 36078
rect 2652 36112 2698 36147
rect 2652 36078 2658 36112
rect 2692 36078 2698 36112
rect 2652 36043 2698 36078
rect 2748 36112 2794 36147
rect 2748 36078 2754 36112
rect 2788 36078 2794 36112
rect 2748 36043 2794 36078
rect 2844 36112 2890 36147
rect 2844 36078 2850 36112
rect 2884 36078 2890 36112
rect 2844 36043 2890 36078
rect 2940 36112 2986 36147
rect 2940 36078 2946 36112
rect 2980 36078 2986 36112
rect 2940 36043 2986 36078
rect 3036 36112 3082 36147
rect 3036 36078 3042 36112
rect 3076 36078 3082 36112
rect 3036 36043 3082 36078
rect 3132 36112 3178 36147
rect 3132 36078 3138 36112
rect 3172 36078 3178 36112
rect 3132 36043 3178 36078
rect 3228 36112 3274 36147
rect 3228 36078 3234 36112
rect 3268 36078 3274 36112
rect 3228 36043 3274 36078
rect 3324 36112 3370 36147
rect 3324 36078 3330 36112
rect 3364 36078 3370 36112
rect 3324 36043 3370 36078
rect 3420 36112 3466 36147
rect 3420 36078 3426 36112
rect 3460 36078 3466 36112
rect 3420 36043 3466 36078
rect 3534 36120 3540 36154
rect 3574 36152 3580 36154
rect 3803 36152 3837 36280
rect 3574 36151 3680 36152
rect 3734 36151 3837 36152
rect 3574 36139 3687 36151
rect 3574 36120 3647 36139
rect 3534 36082 3647 36120
rect 3534 36048 3540 36082
rect 3574 36063 3647 36082
rect 3681 36063 3687 36139
rect 3574 36052 3687 36063
rect 3574 36048 3580 36052
rect 3641 36051 3687 36052
rect 3729 36139 3837 36151
rect 3987 36314 4021 36455
rect 4179 36314 4213 36455
rect 4371 36314 4405 36455
rect 4563 36314 4597 36455
rect 4755 36314 4789 36455
rect 4947 36314 4981 36455
rect 5055 36417 5101 36461
rect 5683 36368 5743 37621
rect 5177 36334 5743 36368
rect 5177 36314 5211 36334
rect 3987 36280 5211 36314
rect 3987 36147 4021 36280
rect 4179 36147 4213 36280
rect 4371 36147 4405 36280
rect 4563 36147 4597 36280
rect 4755 36147 4789 36280
rect 4947 36147 4981 36280
rect 5438 36276 5512 36277
rect 5326 36274 5400 36275
rect 5326 36222 5337 36274
rect 5389 36222 5400 36274
rect 5438 36224 5449 36276
rect 5501 36224 5512 36276
rect 5438 36223 5512 36224
rect 5326 36221 5400 36222
rect 5055 36154 5101 36177
rect 3729 36063 3735 36139
rect 3769 36063 3837 36139
rect 3729 36052 3837 36063
rect 3729 36051 3775 36052
rect 2450 36012 2516 36015
rect 2447 35960 2457 36012
rect 2509 35960 2519 36012
rect 2450 35955 2516 35960
rect 2562 35903 2596 36043
rect 2642 36012 2708 36015
rect 2638 35960 2648 36012
rect 2700 35960 2710 36012
rect 2642 35955 2708 35960
rect 2754 35903 2788 36043
rect 2834 36012 2900 36015
rect 2830 35960 2840 36012
rect 2892 35960 2902 36012
rect 2834 35955 2900 35960
rect 2946 35903 2980 36043
rect 3026 36012 3092 36015
rect 3022 35960 3032 36012
rect 3084 35960 3094 36012
rect 3026 35955 3092 35960
rect 3138 35903 3172 36043
rect 3218 36011 3284 36015
rect 3215 35959 3225 36011
rect 3277 35959 3287 36011
rect 3218 35955 3284 35959
rect 3330 35903 3364 36043
rect 3410 36011 3476 36015
rect 3407 35959 3417 36011
rect 3469 35959 3479 36011
rect 3534 36010 3580 36048
rect 3534 35976 3540 36010
rect 3574 35976 3580 36010
rect 3410 35955 3476 35959
rect 2282 35869 3364 35903
rect 3534 35793 3580 35976
rect 3803 35903 3837 36052
rect 3981 36112 4027 36147
rect 3981 36078 3987 36112
rect 4021 36078 4027 36112
rect 3981 36043 4027 36078
rect 4077 36112 4123 36147
rect 4077 36078 4083 36112
rect 4117 36078 4123 36112
rect 4077 36043 4123 36078
rect 4173 36112 4219 36147
rect 4173 36078 4179 36112
rect 4213 36078 4219 36112
rect 4173 36043 4219 36078
rect 4269 36112 4315 36147
rect 4269 36078 4275 36112
rect 4309 36078 4315 36112
rect 4269 36043 4315 36078
rect 4365 36112 4411 36147
rect 4365 36078 4371 36112
rect 4405 36078 4411 36112
rect 4365 36043 4411 36078
rect 4461 36112 4507 36147
rect 4461 36078 4467 36112
rect 4501 36078 4507 36112
rect 4461 36043 4507 36078
rect 4557 36112 4603 36147
rect 4557 36078 4563 36112
rect 4597 36078 4603 36112
rect 4557 36043 4603 36078
rect 4653 36112 4699 36147
rect 4653 36078 4659 36112
rect 4693 36078 4699 36112
rect 4653 36043 4699 36078
rect 4749 36112 4795 36147
rect 4749 36078 4755 36112
rect 4789 36078 4795 36112
rect 4749 36043 4795 36078
rect 4845 36112 4891 36147
rect 4845 36078 4851 36112
rect 4885 36078 4891 36112
rect 4845 36043 4891 36078
rect 4941 36112 4987 36147
rect 4941 36078 4947 36112
rect 4981 36078 4987 36112
rect 4941 36043 4987 36078
rect 5055 36120 5061 36154
rect 5095 36120 5101 36154
rect 5055 36082 5101 36120
rect 5055 36048 5061 36082
rect 5095 36065 5101 36082
rect 5095 36048 5550 36065
rect 3971 36012 4037 36015
rect 3968 35960 3978 36012
rect 4030 35960 4040 36012
rect 3971 35955 4037 35960
rect 4083 35903 4117 36043
rect 4163 36012 4229 36015
rect 4159 35960 4169 36012
rect 4221 35960 4231 36012
rect 4163 35955 4229 35960
rect 4275 35903 4309 36043
rect 4355 36012 4421 36015
rect 4351 35960 4361 36012
rect 4413 35960 4423 36012
rect 4355 35955 4421 35960
rect 4467 35903 4501 36043
rect 4547 36012 4613 36015
rect 4543 35960 4553 36012
rect 4605 35960 4615 36012
rect 4547 35955 4613 35960
rect 4659 35903 4693 36043
rect 4739 36011 4805 36015
rect 4736 35959 4746 36011
rect 4798 35959 4808 36011
rect 4739 35955 4805 35959
rect 4851 35903 4885 36043
rect 5055 36034 5550 36048
rect 4931 36011 4997 36015
rect 4928 35959 4938 36011
rect 4990 35959 5000 36011
rect 5055 36010 5303 36034
rect 5055 35976 5061 36010
rect 5095 36000 5303 36010
rect 5337 36000 5395 36034
rect 5429 36000 5487 36034
rect 5521 36000 5550 36034
rect 5095 35976 5550 36000
rect 5055 35969 5550 35976
rect 4931 35955 4997 35959
rect 3803 35869 4885 35903
rect 5055 35794 5101 35969
rect 129 35586 1211 35620
rect 129 35023 163 35586
rect 294 35476 304 35528
rect 356 35476 366 35528
rect 409 35436 443 35586
rect 487 35476 497 35528
rect 549 35476 559 35528
rect 601 35436 635 35586
rect 678 35476 688 35528
rect 740 35476 750 35528
rect 793 35436 827 35586
rect 870 35476 880 35528
rect 932 35476 942 35528
rect 985 35436 1019 35586
rect 1062 35476 1072 35528
rect 1124 35476 1134 35528
rect 1177 35436 1211 35586
rect 1254 35476 1264 35528
rect 1316 35476 1326 35528
rect 1381 35492 1427 35656
rect 2282 35590 3364 35624
rect 1381 35458 1387 35492
rect 1421 35458 1427 35492
rect 1512 35469 1522 35529
rect 1578 35469 1792 35529
rect 1852 35469 1862 35529
rect 307 35389 353 35436
rect 307 35355 313 35389
rect 347 35355 353 35389
rect 307 35317 353 35355
rect 307 35283 313 35317
rect 347 35283 353 35317
rect 307 35245 353 35283
rect 307 35211 313 35245
rect 347 35211 353 35245
rect 307 35164 353 35211
rect 403 35389 449 35436
rect 403 35355 409 35389
rect 443 35355 449 35389
rect 403 35317 449 35355
rect 403 35283 409 35317
rect 443 35283 449 35317
rect 403 35245 449 35283
rect 403 35211 409 35245
rect 443 35211 449 35245
rect 403 35164 449 35211
rect 499 35389 545 35436
rect 499 35355 505 35389
rect 539 35355 545 35389
rect 499 35317 545 35355
rect 499 35283 505 35317
rect 539 35283 545 35317
rect 499 35245 545 35283
rect 499 35211 505 35245
rect 539 35211 545 35245
rect 499 35164 545 35211
rect 595 35389 641 35436
rect 595 35355 601 35389
rect 635 35355 641 35389
rect 595 35317 641 35355
rect 595 35283 601 35317
rect 635 35283 641 35317
rect 595 35245 641 35283
rect 595 35211 601 35245
rect 635 35211 641 35245
rect 595 35164 641 35211
rect 691 35389 737 35436
rect 691 35355 697 35389
rect 731 35355 737 35389
rect 691 35317 737 35355
rect 691 35283 697 35317
rect 731 35283 737 35317
rect 691 35245 737 35283
rect 691 35211 697 35245
rect 731 35211 737 35245
rect 691 35164 737 35211
rect 787 35389 833 35436
rect 787 35355 793 35389
rect 827 35355 833 35389
rect 787 35317 833 35355
rect 787 35283 793 35317
rect 827 35283 833 35317
rect 787 35245 833 35283
rect 787 35211 793 35245
rect 827 35211 833 35245
rect 787 35164 833 35211
rect 883 35389 929 35436
rect 883 35355 889 35389
rect 923 35355 929 35389
rect 883 35317 929 35355
rect 883 35283 889 35317
rect 923 35283 929 35317
rect 883 35245 929 35283
rect 883 35211 889 35245
rect 923 35211 929 35245
rect 883 35164 929 35211
rect 979 35389 1025 35436
rect 979 35355 985 35389
rect 1019 35355 1025 35389
rect 979 35317 1025 35355
rect 979 35283 985 35317
rect 1019 35283 1025 35317
rect 979 35245 1025 35283
rect 979 35211 985 35245
rect 1019 35211 1025 35245
rect 979 35164 1025 35211
rect 1075 35389 1121 35436
rect 1075 35355 1081 35389
rect 1115 35355 1121 35389
rect 1075 35317 1121 35355
rect 1075 35283 1081 35317
rect 1115 35283 1121 35317
rect 1075 35245 1121 35283
rect 1075 35211 1081 35245
rect 1115 35211 1121 35245
rect 1075 35164 1121 35211
rect 1171 35389 1217 35436
rect 1171 35355 1177 35389
rect 1211 35355 1217 35389
rect 1171 35317 1217 35355
rect 1171 35283 1177 35317
rect 1211 35283 1217 35317
rect 1171 35245 1217 35283
rect 1171 35211 1177 35245
rect 1211 35211 1217 35245
rect 1171 35164 1217 35211
rect 1267 35389 1313 35436
rect 1267 35355 1273 35389
rect 1307 35355 1313 35389
rect 1267 35317 1313 35355
rect 1267 35283 1273 35317
rect 1307 35283 1313 35317
rect 1267 35245 1313 35283
rect 1267 35211 1273 35245
rect 1307 35211 1313 35245
rect 1267 35164 1313 35211
rect 1381 35420 1427 35458
rect 1381 35386 1387 35420
rect 1421 35386 1427 35420
rect 1381 35348 1427 35386
rect 1381 35314 1387 35348
rect 1421 35314 1427 35348
rect 1381 35276 1427 35314
rect 1381 35242 1387 35276
rect 1421 35242 1427 35276
rect 1381 35232 1427 35242
rect 1381 35230 2160 35232
rect 1381 35204 2056 35230
rect 1381 35179 1387 35204
rect 1380 35170 1387 35179
rect 1421 35170 2056 35204
rect 0 34989 163 35023
rect 129 34612 163 34989
rect 313 35023 347 35164
rect 505 35023 539 35164
rect 697 35023 731 35164
rect 889 35023 923 35164
rect 1081 35023 1115 35164
rect 1273 35023 1307 35164
rect 1380 35122 2056 35170
rect 2190 35122 2200 35230
rect 1380 35120 2160 35122
rect 2282 35027 2316 35590
rect 2447 35480 2457 35532
rect 2509 35480 2519 35532
rect 2562 35440 2596 35590
rect 2640 35480 2650 35532
rect 2702 35480 2712 35532
rect 2754 35440 2788 35590
rect 2831 35480 2841 35532
rect 2893 35480 2903 35532
rect 2946 35440 2980 35590
rect 3023 35480 3033 35532
rect 3085 35480 3095 35532
rect 3138 35440 3172 35590
rect 3215 35480 3225 35532
rect 3277 35480 3287 35532
rect 3330 35440 3364 35590
rect 3407 35480 3417 35532
rect 3469 35480 3479 35532
rect 3534 35496 3580 35704
rect 3534 35462 3540 35496
rect 3574 35462 3580 35496
rect 2460 35393 2506 35440
rect 2460 35359 2466 35393
rect 2500 35359 2506 35393
rect 2460 35321 2506 35359
rect 2460 35287 2466 35321
rect 2500 35287 2506 35321
rect 2460 35249 2506 35287
rect 2460 35215 2466 35249
rect 2500 35215 2506 35249
rect 2460 35168 2506 35215
rect 2556 35393 2602 35440
rect 2556 35359 2562 35393
rect 2596 35359 2602 35393
rect 2556 35321 2602 35359
rect 2556 35287 2562 35321
rect 2596 35287 2602 35321
rect 2556 35249 2602 35287
rect 2556 35215 2562 35249
rect 2596 35215 2602 35249
rect 2556 35168 2602 35215
rect 2652 35393 2698 35440
rect 2652 35359 2658 35393
rect 2692 35359 2698 35393
rect 2652 35321 2698 35359
rect 2652 35287 2658 35321
rect 2692 35287 2698 35321
rect 2652 35249 2698 35287
rect 2652 35215 2658 35249
rect 2692 35215 2698 35249
rect 2652 35168 2698 35215
rect 2748 35393 2794 35440
rect 2748 35359 2754 35393
rect 2788 35359 2794 35393
rect 2748 35321 2794 35359
rect 2748 35287 2754 35321
rect 2788 35287 2794 35321
rect 2748 35249 2794 35287
rect 2748 35215 2754 35249
rect 2788 35215 2794 35249
rect 2748 35168 2794 35215
rect 2844 35393 2890 35440
rect 2844 35359 2850 35393
rect 2884 35359 2890 35393
rect 2844 35321 2890 35359
rect 2844 35287 2850 35321
rect 2884 35287 2890 35321
rect 2844 35249 2890 35287
rect 2844 35215 2850 35249
rect 2884 35215 2890 35249
rect 2844 35168 2890 35215
rect 2940 35393 2986 35440
rect 2940 35359 2946 35393
rect 2980 35359 2986 35393
rect 2940 35321 2986 35359
rect 2940 35287 2946 35321
rect 2980 35287 2986 35321
rect 2940 35249 2986 35287
rect 2940 35215 2946 35249
rect 2980 35215 2986 35249
rect 2940 35168 2986 35215
rect 3036 35393 3082 35440
rect 3036 35359 3042 35393
rect 3076 35359 3082 35393
rect 3036 35321 3082 35359
rect 3036 35287 3042 35321
rect 3076 35287 3082 35321
rect 3036 35249 3082 35287
rect 3036 35215 3042 35249
rect 3076 35215 3082 35249
rect 3036 35168 3082 35215
rect 3132 35393 3178 35440
rect 3132 35359 3138 35393
rect 3172 35359 3178 35393
rect 3132 35321 3178 35359
rect 3132 35287 3138 35321
rect 3172 35287 3178 35321
rect 3132 35249 3178 35287
rect 3132 35215 3138 35249
rect 3172 35215 3178 35249
rect 3132 35168 3178 35215
rect 3228 35393 3274 35440
rect 3228 35359 3234 35393
rect 3268 35359 3274 35393
rect 3228 35321 3274 35359
rect 3228 35287 3234 35321
rect 3268 35287 3274 35321
rect 3228 35249 3274 35287
rect 3228 35215 3234 35249
rect 3268 35215 3274 35249
rect 3228 35168 3274 35215
rect 3324 35393 3370 35440
rect 3324 35359 3330 35393
rect 3364 35359 3370 35393
rect 3324 35321 3370 35359
rect 3324 35287 3330 35321
rect 3364 35287 3370 35321
rect 3324 35249 3370 35287
rect 3324 35215 3330 35249
rect 3364 35215 3370 35249
rect 3324 35168 3370 35215
rect 3420 35393 3466 35440
rect 3420 35359 3426 35393
rect 3460 35359 3466 35393
rect 3420 35321 3466 35359
rect 3420 35287 3426 35321
rect 3460 35287 3466 35321
rect 3420 35249 3466 35287
rect 3420 35215 3426 35249
rect 3460 35215 3466 35249
rect 3420 35168 3466 35215
rect 3534 35424 3580 35462
rect 3534 35390 3540 35424
rect 3574 35390 3580 35424
rect 3534 35352 3580 35390
rect 3534 35318 3540 35352
rect 3574 35318 3580 35352
rect 3534 35280 3580 35318
rect 3534 35246 3540 35280
rect 3574 35246 3580 35280
rect 3534 35208 3580 35246
rect 3534 35174 3540 35208
rect 3574 35174 3580 35208
rect 2101 35023 2316 35027
rect 313 34993 2316 35023
rect 313 34989 2141 34993
rect 313 34856 347 34989
rect 505 34856 539 34989
rect 697 34856 731 34989
rect 889 34856 923 34989
rect 1081 34856 1115 34989
rect 1273 34856 1307 34989
rect 1381 34863 1608 34886
rect 307 34821 353 34856
rect 307 34787 313 34821
rect 347 34787 353 34821
rect 307 34752 353 34787
rect 403 34821 449 34856
rect 403 34787 409 34821
rect 443 34787 449 34821
rect 403 34752 449 34787
rect 499 34821 545 34856
rect 499 34787 505 34821
rect 539 34787 545 34821
rect 499 34752 545 34787
rect 595 34821 641 34856
rect 595 34787 601 34821
rect 635 34787 641 34821
rect 595 34752 641 34787
rect 691 34821 737 34856
rect 691 34787 697 34821
rect 731 34787 737 34821
rect 691 34752 737 34787
rect 787 34821 833 34856
rect 787 34787 793 34821
rect 827 34787 833 34821
rect 787 34752 833 34787
rect 883 34821 929 34856
rect 883 34787 889 34821
rect 923 34787 929 34821
rect 883 34752 929 34787
rect 979 34821 1025 34856
rect 979 34787 985 34821
rect 1019 34787 1025 34821
rect 979 34752 1025 34787
rect 1075 34821 1121 34856
rect 1075 34787 1081 34821
rect 1115 34787 1121 34821
rect 1075 34752 1121 34787
rect 1171 34821 1217 34856
rect 1171 34787 1177 34821
rect 1211 34787 1217 34821
rect 1171 34752 1217 34787
rect 1267 34821 1313 34856
rect 1267 34787 1273 34821
rect 1307 34787 1313 34821
rect 1267 34752 1313 34787
rect 1381 34829 1387 34863
rect 1421 34829 1608 34863
rect 1381 34791 1608 34829
rect 1381 34757 1387 34791
rect 1421 34766 1608 34791
rect 1421 34757 1427 34766
rect 1560 34764 1608 34766
rect 1598 34762 1608 34764
rect 1720 34762 1730 34886
rect 297 34721 363 34724
rect 294 34669 304 34721
rect 356 34669 366 34721
rect 297 34664 363 34669
rect 409 34612 443 34752
rect 489 34721 555 34724
rect 485 34669 495 34721
rect 547 34669 557 34721
rect 489 34664 555 34669
rect 601 34612 635 34752
rect 681 34721 747 34724
rect 677 34669 687 34721
rect 739 34669 749 34721
rect 681 34664 747 34669
rect 793 34612 827 34752
rect 873 34721 939 34724
rect 869 34669 879 34721
rect 931 34669 941 34721
rect 873 34664 939 34669
rect 985 34612 1019 34752
rect 1065 34720 1131 34724
rect 1062 34668 1072 34720
rect 1124 34668 1134 34720
rect 1065 34664 1131 34668
rect 1177 34612 1211 34752
rect 1257 34720 1323 34724
rect 1254 34668 1264 34720
rect 1316 34668 1326 34720
rect 1381 34719 1427 34757
rect 1920 34724 1930 34726
rect 1381 34685 1387 34719
rect 1421 34685 1427 34719
rect 1257 34664 1323 34668
rect 129 34578 1211 34612
rect 1381 34542 1427 34685
rect 1458 34668 1468 34724
rect 1524 34670 1930 34724
rect 1986 34670 1996 34726
rect 1524 34668 1986 34670
rect 2282 34616 2316 34993
rect 2466 35027 2500 35168
rect 2658 35027 2692 35168
rect 2850 35027 2884 35168
rect 3042 35027 3076 35168
rect 3234 35027 3268 35168
rect 3426 35027 3460 35168
rect 3534 35130 3580 35174
rect 3803 35590 4885 35624
rect 3803 35027 3837 35590
rect 3968 35480 3978 35532
rect 4030 35480 4040 35532
rect 4083 35440 4117 35590
rect 4161 35480 4171 35532
rect 4223 35480 4233 35532
rect 4275 35440 4309 35590
rect 4352 35480 4362 35532
rect 4414 35480 4424 35532
rect 4467 35440 4501 35590
rect 4544 35480 4554 35532
rect 4606 35480 4616 35532
rect 4659 35440 4693 35590
rect 4736 35480 4746 35532
rect 4798 35480 4808 35532
rect 4851 35440 4885 35590
rect 4928 35480 4938 35532
rect 4990 35480 5000 35532
rect 5055 35496 5101 35701
rect 5055 35462 5061 35496
rect 5095 35462 5101 35496
rect 3981 35393 4027 35440
rect 3981 35359 3987 35393
rect 4021 35359 4027 35393
rect 3981 35321 4027 35359
rect 3981 35287 3987 35321
rect 4021 35287 4027 35321
rect 3981 35249 4027 35287
rect 3981 35215 3987 35249
rect 4021 35215 4027 35249
rect 3981 35168 4027 35215
rect 4077 35393 4123 35440
rect 4077 35359 4083 35393
rect 4117 35359 4123 35393
rect 4077 35321 4123 35359
rect 4077 35287 4083 35321
rect 4117 35287 4123 35321
rect 4077 35249 4123 35287
rect 4077 35215 4083 35249
rect 4117 35215 4123 35249
rect 4077 35168 4123 35215
rect 4173 35393 4219 35440
rect 4173 35359 4179 35393
rect 4213 35359 4219 35393
rect 4173 35321 4219 35359
rect 4173 35287 4179 35321
rect 4213 35287 4219 35321
rect 4173 35249 4219 35287
rect 4173 35215 4179 35249
rect 4213 35215 4219 35249
rect 4173 35168 4219 35215
rect 4269 35393 4315 35440
rect 4269 35359 4275 35393
rect 4309 35359 4315 35393
rect 4269 35321 4315 35359
rect 4269 35287 4275 35321
rect 4309 35287 4315 35321
rect 4269 35249 4315 35287
rect 4269 35215 4275 35249
rect 4309 35215 4315 35249
rect 4269 35168 4315 35215
rect 4365 35393 4411 35440
rect 4365 35359 4371 35393
rect 4405 35359 4411 35393
rect 4365 35321 4411 35359
rect 4365 35287 4371 35321
rect 4405 35287 4411 35321
rect 4365 35249 4411 35287
rect 4365 35215 4371 35249
rect 4405 35215 4411 35249
rect 4365 35168 4411 35215
rect 4461 35393 4507 35440
rect 4461 35359 4467 35393
rect 4501 35359 4507 35393
rect 4461 35321 4507 35359
rect 4461 35287 4467 35321
rect 4501 35287 4507 35321
rect 4461 35249 4507 35287
rect 4461 35215 4467 35249
rect 4501 35215 4507 35249
rect 4461 35168 4507 35215
rect 4557 35393 4603 35440
rect 4557 35359 4563 35393
rect 4597 35359 4603 35393
rect 4557 35321 4603 35359
rect 4557 35287 4563 35321
rect 4597 35287 4603 35321
rect 4557 35249 4603 35287
rect 4557 35215 4563 35249
rect 4597 35215 4603 35249
rect 4557 35168 4603 35215
rect 4653 35393 4699 35440
rect 4653 35359 4659 35393
rect 4693 35359 4699 35393
rect 4653 35321 4699 35359
rect 4653 35287 4659 35321
rect 4693 35287 4699 35321
rect 4653 35249 4699 35287
rect 4653 35215 4659 35249
rect 4693 35215 4699 35249
rect 4653 35168 4699 35215
rect 4749 35393 4795 35440
rect 4749 35359 4755 35393
rect 4789 35359 4795 35393
rect 4749 35321 4795 35359
rect 4749 35287 4755 35321
rect 4789 35287 4795 35321
rect 4749 35249 4795 35287
rect 4749 35215 4755 35249
rect 4789 35215 4795 35249
rect 4749 35168 4795 35215
rect 4845 35393 4891 35440
rect 4845 35359 4851 35393
rect 4885 35359 4891 35393
rect 4845 35321 4891 35359
rect 4845 35287 4851 35321
rect 4885 35287 4891 35321
rect 4845 35249 4891 35287
rect 4845 35215 4851 35249
rect 4885 35215 4891 35249
rect 4845 35168 4891 35215
rect 4941 35393 4987 35440
rect 4941 35359 4947 35393
rect 4981 35359 4987 35393
rect 4941 35321 4987 35359
rect 4941 35287 4947 35321
rect 4981 35287 4987 35321
rect 4941 35249 4987 35287
rect 4941 35215 4947 35249
rect 4981 35215 4987 35249
rect 4941 35168 4987 35215
rect 5055 35424 5101 35462
rect 5055 35390 5061 35424
rect 5095 35390 5101 35424
rect 5055 35352 5101 35390
rect 5055 35318 5061 35352
rect 5095 35321 5101 35352
rect 5274 35321 5550 35322
rect 5095 35318 5550 35321
rect 5055 35291 5550 35318
rect 5055 35280 5303 35291
rect 5055 35246 5061 35280
rect 5095 35257 5303 35280
rect 5337 35257 5395 35291
rect 5429 35257 5487 35291
rect 5521 35257 5550 35291
rect 5095 35246 5550 35257
rect 5055 35226 5550 35246
rect 5055 35208 5101 35226
rect 5055 35174 5061 35208
rect 5095 35174 5101 35208
rect 2466 34993 3837 35027
rect 2466 34860 2500 34993
rect 2658 34860 2692 34993
rect 2850 34860 2884 34993
rect 3042 34860 3076 34993
rect 3234 34860 3268 34993
rect 3426 34860 3460 34993
rect 3671 34903 3681 34955
rect 3733 34903 3743 34955
rect 3679 34902 3691 34903
rect 3725 34902 3737 34903
rect 3679 34896 3737 34902
rect 3534 34867 3580 34890
rect 2460 34825 2506 34860
rect 2460 34791 2466 34825
rect 2500 34791 2506 34825
rect 2460 34756 2506 34791
rect 2556 34825 2602 34860
rect 2556 34791 2562 34825
rect 2596 34791 2602 34825
rect 2556 34756 2602 34791
rect 2652 34825 2698 34860
rect 2652 34791 2658 34825
rect 2692 34791 2698 34825
rect 2652 34756 2698 34791
rect 2748 34825 2794 34860
rect 2748 34791 2754 34825
rect 2788 34791 2794 34825
rect 2748 34756 2794 34791
rect 2844 34825 2890 34860
rect 2844 34791 2850 34825
rect 2884 34791 2890 34825
rect 2844 34756 2890 34791
rect 2940 34825 2986 34860
rect 2940 34791 2946 34825
rect 2980 34791 2986 34825
rect 2940 34756 2986 34791
rect 3036 34825 3082 34860
rect 3036 34791 3042 34825
rect 3076 34791 3082 34825
rect 3036 34756 3082 34791
rect 3132 34825 3178 34860
rect 3132 34791 3138 34825
rect 3172 34791 3178 34825
rect 3132 34756 3178 34791
rect 3228 34825 3274 34860
rect 3228 34791 3234 34825
rect 3268 34791 3274 34825
rect 3228 34756 3274 34791
rect 3324 34825 3370 34860
rect 3324 34791 3330 34825
rect 3364 34791 3370 34825
rect 3324 34756 3370 34791
rect 3420 34825 3466 34860
rect 3420 34791 3426 34825
rect 3460 34791 3466 34825
rect 3420 34756 3466 34791
rect 3534 34833 3540 34867
rect 3574 34865 3580 34867
rect 3803 34865 3837 34993
rect 3574 34864 3680 34865
rect 3734 34864 3837 34865
rect 3574 34852 3687 34864
rect 3574 34833 3647 34852
rect 3534 34795 3647 34833
rect 3534 34761 3540 34795
rect 3574 34776 3647 34795
rect 3681 34776 3687 34852
rect 3574 34765 3687 34776
rect 3574 34761 3580 34765
rect 3641 34764 3687 34765
rect 3729 34852 3837 34864
rect 3987 35027 4021 35168
rect 4179 35027 4213 35168
rect 4371 35027 4405 35168
rect 4563 35027 4597 35168
rect 4755 35027 4789 35168
rect 4947 35027 4981 35168
rect 5055 35130 5101 35174
rect 5683 35081 5743 36334
rect 5177 35047 5743 35081
rect 5177 35027 5211 35047
rect 3987 34993 5211 35027
rect 3987 34860 4021 34993
rect 4179 34860 4213 34993
rect 4371 34860 4405 34993
rect 4563 34860 4597 34993
rect 4755 34860 4789 34993
rect 4947 34860 4981 34993
rect 5438 34989 5512 34990
rect 5326 34987 5400 34988
rect 5326 34935 5337 34987
rect 5389 34935 5400 34987
rect 5438 34937 5449 34989
rect 5501 34937 5512 34989
rect 5438 34936 5512 34937
rect 5326 34934 5400 34935
rect 5055 34867 5101 34890
rect 3729 34776 3735 34852
rect 3769 34776 3837 34852
rect 3729 34765 3837 34776
rect 3729 34764 3775 34765
rect 2450 34725 2516 34728
rect 2447 34673 2457 34725
rect 2509 34673 2519 34725
rect 2450 34668 2516 34673
rect 2562 34616 2596 34756
rect 2642 34725 2708 34728
rect 2638 34673 2648 34725
rect 2700 34673 2710 34725
rect 2642 34668 2708 34673
rect 2754 34616 2788 34756
rect 2834 34725 2900 34728
rect 2830 34673 2840 34725
rect 2892 34673 2902 34725
rect 2834 34668 2900 34673
rect 2946 34616 2980 34756
rect 3026 34725 3092 34728
rect 3022 34673 3032 34725
rect 3084 34673 3094 34725
rect 3026 34668 3092 34673
rect 3138 34616 3172 34756
rect 3218 34724 3284 34728
rect 3215 34672 3225 34724
rect 3277 34672 3287 34724
rect 3218 34668 3284 34672
rect 3330 34616 3364 34756
rect 3410 34724 3476 34728
rect 3407 34672 3417 34724
rect 3469 34672 3479 34724
rect 3534 34723 3580 34761
rect 3534 34689 3540 34723
rect 3574 34689 3580 34723
rect 3410 34668 3476 34672
rect 2282 34582 3364 34616
rect 3534 34506 3580 34689
rect 3803 34616 3837 34765
rect 3981 34825 4027 34860
rect 3981 34791 3987 34825
rect 4021 34791 4027 34825
rect 3981 34756 4027 34791
rect 4077 34825 4123 34860
rect 4077 34791 4083 34825
rect 4117 34791 4123 34825
rect 4077 34756 4123 34791
rect 4173 34825 4219 34860
rect 4173 34791 4179 34825
rect 4213 34791 4219 34825
rect 4173 34756 4219 34791
rect 4269 34825 4315 34860
rect 4269 34791 4275 34825
rect 4309 34791 4315 34825
rect 4269 34756 4315 34791
rect 4365 34825 4411 34860
rect 4365 34791 4371 34825
rect 4405 34791 4411 34825
rect 4365 34756 4411 34791
rect 4461 34825 4507 34860
rect 4461 34791 4467 34825
rect 4501 34791 4507 34825
rect 4461 34756 4507 34791
rect 4557 34825 4603 34860
rect 4557 34791 4563 34825
rect 4597 34791 4603 34825
rect 4557 34756 4603 34791
rect 4653 34825 4699 34860
rect 4653 34791 4659 34825
rect 4693 34791 4699 34825
rect 4653 34756 4699 34791
rect 4749 34825 4795 34860
rect 4749 34791 4755 34825
rect 4789 34791 4795 34825
rect 4749 34756 4795 34791
rect 4845 34825 4891 34860
rect 4845 34791 4851 34825
rect 4885 34791 4891 34825
rect 4845 34756 4891 34791
rect 4941 34825 4987 34860
rect 4941 34791 4947 34825
rect 4981 34791 4987 34825
rect 4941 34756 4987 34791
rect 5055 34833 5061 34867
rect 5095 34833 5101 34867
rect 5055 34795 5101 34833
rect 5055 34761 5061 34795
rect 5095 34778 5101 34795
rect 5095 34761 5550 34778
rect 3971 34725 4037 34728
rect 3968 34673 3978 34725
rect 4030 34673 4040 34725
rect 3971 34668 4037 34673
rect 4083 34616 4117 34756
rect 4163 34725 4229 34728
rect 4159 34673 4169 34725
rect 4221 34673 4231 34725
rect 4163 34668 4229 34673
rect 4275 34616 4309 34756
rect 4355 34725 4421 34728
rect 4351 34673 4361 34725
rect 4413 34673 4423 34725
rect 4355 34668 4421 34673
rect 4467 34616 4501 34756
rect 4547 34725 4613 34728
rect 4543 34673 4553 34725
rect 4605 34673 4615 34725
rect 4547 34668 4613 34673
rect 4659 34616 4693 34756
rect 4739 34724 4805 34728
rect 4736 34672 4746 34724
rect 4798 34672 4808 34724
rect 4739 34668 4805 34672
rect 4851 34616 4885 34756
rect 5055 34747 5550 34761
rect 4931 34724 4997 34728
rect 4928 34672 4938 34724
rect 4990 34672 5000 34724
rect 5055 34723 5303 34747
rect 5055 34689 5061 34723
rect 5095 34713 5303 34723
rect 5337 34713 5395 34747
rect 5429 34713 5487 34747
rect 5521 34713 5550 34747
rect 5095 34689 5550 34713
rect 5055 34682 5550 34689
rect 4931 34668 4997 34672
rect 3803 34582 4885 34616
rect 5055 34507 5101 34682
rect 129 34299 1211 34333
rect 129 33736 163 34299
rect 294 34189 304 34241
rect 356 34189 366 34241
rect 409 34149 443 34299
rect 487 34189 497 34241
rect 549 34189 559 34241
rect 601 34149 635 34299
rect 678 34189 688 34241
rect 740 34189 750 34241
rect 793 34149 827 34299
rect 870 34189 880 34241
rect 932 34189 942 34241
rect 985 34149 1019 34299
rect 1062 34189 1072 34241
rect 1124 34189 1134 34241
rect 1177 34149 1211 34299
rect 1254 34189 1264 34241
rect 1316 34189 1326 34241
rect 1381 34205 1427 34369
rect 2282 34303 3364 34337
rect 1381 34171 1387 34205
rect 1421 34171 1427 34205
rect 1512 34182 1522 34242
rect 1578 34182 1792 34242
rect 1852 34182 1862 34242
rect 307 34102 353 34149
rect 307 34068 313 34102
rect 347 34068 353 34102
rect 307 34030 353 34068
rect 307 33996 313 34030
rect 347 33996 353 34030
rect 307 33958 353 33996
rect 307 33924 313 33958
rect 347 33924 353 33958
rect 307 33877 353 33924
rect 403 34102 449 34149
rect 403 34068 409 34102
rect 443 34068 449 34102
rect 403 34030 449 34068
rect 403 33996 409 34030
rect 443 33996 449 34030
rect 403 33958 449 33996
rect 403 33924 409 33958
rect 443 33924 449 33958
rect 403 33877 449 33924
rect 499 34102 545 34149
rect 499 34068 505 34102
rect 539 34068 545 34102
rect 499 34030 545 34068
rect 499 33996 505 34030
rect 539 33996 545 34030
rect 499 33958 545 33996
rect 499 33924 505 33958
rect 539 33924 545 33958
rect 499 33877 545 33924
rect 595 34102 641 34149
rect 595 34068 601 34102
rect 635 34068 641 34102
rect 595 34030 641 34068
rect 595 33996 601 34030
rect 635 33996 641 34030
rect 595 33958 641 33996
rect 595 33924 601 33958
rect 635 33924 641 33958
rect 595 33877 641 33924
rect 691 34102 737 34149
rect 691 34068 697 34102
rect 731 34068 737 34102
rect 691 34030 737 34068
rect 691 33996 697 34030
rect 731 33996 737 34030
rect 691 33958 737 33996
rect 691 33924 697 33958
rect 731 33924 737 33958
rect 691 33877 737 33924
rect 787 34102 833 34149
rect 787 34068 793 34102
rect 827 34068 833 34102
rect 787 34030 833 34068
rect 787 33996 793 34030
rect 827 33996 833 34030
rect 787 33958 833 33996
rect 787 33924 793 33958
rect 827 33924 833 33958
rect 787 33877 833 33924
rect 883 34102 929 34149
rect 883 34068 889 34102
rect 923 34068 929 34102
rect 883 34030 929 34068
rect 883 33996 889 34030
rect 923 33996 929 34030
rect 883 33958 929 33996
rect 883 33924 889 33958
rect 923 33924 929 33958
rect 883 33877 929 33924
rect 979 34102 1025 34149
rect 979 34068 985 34102
rect 1019 34068 1025 34102
rect 979 34030 1025 34068
rect 979 33996 985 34030
rect 1019 33996 1025 34030
rect 979 33958 1025 33996
rect 979 33924 985 33958
rect 1019 33924 1025 33958
rect 979 33877 1025 33924
rect 1075 34102 1121 34149
rect 1075 34068 1081 34102
rect 1115 34068 1121 34102
rect 1075 34030 1121 34068
rect 1075 33996 1081 34030
rect 1115 33996 1121 34030
rect 1075 33958 1121 33996
rect 1075 33924 1081 33958
rect 1115 33924 1121 33958
rect 1075 33877 1121 33924
rect 1171 34102 1217 34149
rect 1171 34068 1177 34102
rect 1211 34068 1217 34102
rect 1171 34030 1217 34068
rect 1171 33996 1177 34030
rect 1211 33996 1217 34030
rect 1171 33958 1217 33996
rect 1171 33924 1177 33958
rect 1211 33924 1217 33958
rect 1171 33877 1217 33924
rect 1267 34102 1313 34149
rect 1267 34068 1273 34102
rect 1307 34068 1313 34102
rect 1267 34030 1313 34068
rect 1267 33996 1273 34030
rect 1307 33996 1313 34030
rect 1267 33958 1313 33996
rect 1267 33924 1273 33958
rect 1307 33924 1313 33958
rect 1267 33877 1313 33924
rect 1381 34133 1427 34171
rect 1381 34099 1387 34133
rect 1421 34099 1427 34133
rect 1381 34061 1427 34099
rect 1381 34027 1387 34061
rect 1421 34027 1427 34061
rect 1381 33989 1427 34027
rect 1381 33955 1387 33989
rect 1421 33955 1427 33989
rect 1381 33945 1427 33955
rect 1381 33943 2160 33945
rect 1381 33917 2056 33943
rect 1381 33892 1387 33917
rect 1380 33883 1387 33892
rect 1421 33883 2056 33917
rect 0 33702 163 33736
rect 129 33325 163 33702
rect 313 33736 347 33877
rect 505 33736 539 33877
rect 697 33736 731 33877
rect 889 33736 923 33877
rect 1081 33736 1115 33877
rect 1273 33736 1307 33877
rect 1380 33835 2056 33883
rect 2190 33835 2200 33943
rect 1380 33833 2160 33835
rect 2282 33740 2316 34303
rect 2447 34193 2457 34245
rect 2509 34193 2519 34245
rect 2562 34153 2596 34303
rect 2640 34193 2650 34245
rect 2702 34193 2712 34245
rect 2754 34153 2788 34303
rect 2831 34193 2841 34245
rect 2893 34193 2903 34245
rect 2946 34153 2980 34303
rect 3023 34193 3033 34245
rect 3085 34193 3095 34245
rect 3138 34153 3172 34303
rect 3215 34193 3225 34245
rect 3277 34193 3287 34245
rect 3330 34153 3364 34303
rect 3407 34193 3417 34245
rect 3469 34193 3479 34245
rect 3534 34209 3580 34417
rect 3534 34175 3540 34209
rect 3574 34175 3580 34209
rect 2460 34106 2506 34153
rect 2460 34072 2466 34106
rect 2500 34072 2506 34106
rect 2460 34034 2506 34072
rect 2460 34000 2466 34034
rect 2500 34000 2506 34034
rect 2460 33962 2506 34000
rect 2460 33928 2466 33962
rect 2500 33928 2506 33962
rect 2460 33881 2506 33928
rect 2556 34106 2602 34153
rect 2556 34072 2562 34106
rect 2596 34072 2602 34106
rect 2556 34034 2602 34072
rect 2556 34000 2562 34034
rect 2596 34000 2602 34034
rect 2556 33962 2602 34000
rect 2556 33928 2562 33962
rect 2596 33928 2602 33962
rect 2556 33881 2602 33928
rect 2652 34106 2698 34153
rect 2652 34072 2658 34106
rect 2692 34072 2698 34106
rect 2652 34034 2698 34072
rect 2652 34000 2658 34034
rect 2692 34000 2698 34034
rect 2652 33962 2698 34000
rect 2652 33928 2658 33962
rect 2692 33928 2698 33962
rect 2652 33881 2698 33928
rect 2748 34106 2794 34153
rect 2748 34072 2754 34106
rect 2788 34072 2794 34106
rect 2748 34034 2794 34072
rect 2748 34000 2754 34034
rect 2788 34000 2794 34034
rect 2748 33962 2794 34000
rect 2748 33928 2754 33962
rect 2788 33928 2794 33962
rect 2748 33881 2794 33928
rect 2844 34106 2890 34153
rect 2844 34072 2850 34106
rect 2884 34072 2890 34106
rect 2844 34034 2890 34072
rect 2844 34000 2850 34034
rect 2884 34000 2890 34034
rect 2844 33962 2890 34000
rect 2844 33928 2850 33962
rect 2884 33928 2890 33962
rect 2844 33881 2890 33928
rect 2940 34106 2986 34153
rect 2940 34072 2946 34106
rect 2980 34072 2986 34106
rect 2940 34034 2986 34072
rect 2940 34000 2946 34034
rect 2980 34000 2986 34034
rect 2940 33962 2986 34000
rect 2940 33928 2946 33962
rect 2980 33928 2986 33962
rect 2940 33881 2986 33928
rect 3036 34106 3082 34153
rect 3036 34072 3042 34106
rect 3076 34072 3082 34106
rect 3036 34034 3082 34072
rect 3036 34000 3042 34034
rect 3076 34000 3082 34034
rect 3036 33962 3082 34000
rect 3036 33928 3042 33962
rect 3076 33928 3082 33962
rect 3036 33881 3082 33928
rect 3132 34106 3178 34153
rect 3132 34072 3138 34106
rect 3172 34072 3178 34106
rect 3132 34034 3178 34072
rect 3132 34000 3138 34034
rect 3172 34000 3178 34034
rect 3132 33962 3178 34000
rect 3132 33928 3138 33962
rect 3172 33928 3178 33962
rect 3132 33881 3178 33928
rect 3228 34106 3274 34153
rect 3228 34072 3234 34106
rect 3268 34072 3274 34106
rect 3228 34034 3274 34072
rect 3228 34000 3234 34034
rect 3268 34000 3274 34034
rect 3228 33962 3274 34000
rect 3228 33928 3234 33962
rect 3268 33928 3274 33962
rect 3228 33881 3274 33928
rect 3324 34106 3370 34153
rect 3324 34072 3330 34106
rect 3364 34072 3370 34106
rect 3324 34034 3370 34072
rect 3324 34000 3330 34034
rect 3364 34000 3370 34034
rect 3324 33962 3370 34000
rect 3324 33928 3330 33962
rect 3364 33928 3370 33962
rect 3324 33881 3370 33928
rect 3420 34106 3466 34153
rect 3420 34072 3426 34106
rect 3460 34072 3466 34106
rect 3420 34034 3466 34072
rect 3420 34000 3426 34034
rect 3460 34000 3466 34034
rect 3420 33962 3466 34000
rect 3420 33928 3426 33962
rect 3460 33928 3466 33962
rect 3420 33881 3466 33928
rect 3534 34137 3580 34175
rect 3534 34103 3540 34137
rect 3574 34103 3580 34137
rect 3534 34065 3580 34103
rect 3534 34031 3540 34065
rect 3574 34031 3580 34065
rect 3534 33993 3580 34031
rect 3534 33959 3540 33993
rect 3574 33959 3580 33993
rect 3534 33921 3580 33959
rect 3534 33887 3540 33921
rect 3574 33887 3580 33921
rect 2101 33736 2316 33740
rect 313 33706 2316 33736
rect 313 33702 2141 33706
rect 313 33569 347 33702
rect 505 33569 539 33702
rect 697 33569 731 33702
rect 889 33569 923 33702
rect 1081 33569 1115 33702
rect 1273 33569 1307 33702
rect 1381 33576 1608 33599
rect 307 33534 353 33569
rect 307 33500 313 33534
rect 347 33500 353 33534
rect 307 33465 353 33500
rect 403 33534 449 33569
rect 403 33500 409 33534
rect 443 33500 449 33534
rect 403 33465 449 33500
rect 499 33534 545 33569
rect 499 33500 505 33534
rect 539 33500 545 33534
rect 499 33465 545 33500
rect 595 33534 641 33569
rect 595 33500 601 33534
rect 635 33500 641 33534
rect 595 33465 641 33500
rect 691 33534 737 33569
rect 691 33500 697 33534
rect 731 33500 737 33534
rect 691 33465 737 33500
rect 787 33534 833 33569
rect 787 33500 793 33534
rect 827 33500 833 33534
rect 787 33465 833 33500
rect 883 33534 929 33569
rect 883 33500 889 33534
rect 923 33500 929 33534
rect 883 33465 929 33500
rect 979 33534 1025 33569
rect 979 33500 985 33534
rect 1019 33500 1025 33534
rect 979 33465 1025 33500
rect 1075 33534 1121 33569
rect 1075 33500 1081 33534
rect 1115 33500 1121 33534
rect 1075 33465 1121 33500
rect 1171 33534 1217 33569
rect 1171 33500 1177 33534
rect 1211 33500 1217 33534
rect 1171 33465 1217 33500
rect 1267 33534 1313 33569
rect 1267 33500 1273 33534
rect 1307 33500 1313 33534
rect 1267 33465 1313 33500
rect 1381 33542 1387 33576
rect 1421 33542 1608 33576
rect 1381 33504 1608 33542
rect 1381 33470 1387 33504
rect 1421 33479 1608 33504
rect 1421 33470 1427 33479
rect 1560 33477 1608 33479
rect 1598 33475 1608 33477
rect 1720 33475 1730 33599
rect 297 33434 363 33437
rect 294 33382 304 33434
rect 356 33382 366 33434
rect 297 33377 363 33382
rect 409 33325 443 33465
rect 489 33434 555 33437
rect 485 33382 495 33434
rect 547 33382 557 33434
rect 489 33377 555 33382
rect 601 33325 635 33465
rect 681 33434 747 33437
rect 677 33382 687 33434
rect 739 33382 749 33434
rect 681 33377 747 33382
rect 793 33325 827 33465
rect 873 33434 939 33437
rect 869 33382 879 33434
rect 931 33382 941 33434
rect 873 33377 939 33382
rect 985 33325 1019 33465
rect 1065 33433 1131 33437
rect 1062 33381 1072 33433
rect 1124 33381 1134 33433
rect 1065 33377 1131 33381
rect 1177 33325 1211 33465
rect 1257 33433 1323 33437
rect 1254 33381 1264 33433
rect 1316 33381 1326 33433
rect 1381 33432 1427 33470
rect 1920 33437 1930 33439
rect 1381 33398 1387 33432
rect 1421 33398 1427 33432
rect 1257 33377 1323 33381
rect 129 33291 1211 33325
rect 1381 33255 1427 33398
rect 1458 33381 1468 33437
rect 1524 33383 1930 33437
rect 1986 33383 1996 33439
rect 1524 33381 1986 33383
rect 2282 33329 2316 33706
rect 2466 33740 2500 33881
rect 2658 33740 2692 33881
rect 2850 33740 2884 33881
rect 3042 33740 3076 33881
rect 3234 33740 3268 33881
rect 3426 33740 3460 33881
rect 3534 33843 3580 33887
rect 3803 34303 4885 34337
rect 3803 33740 3837 34303
rect 3968 34193 3978 34245
rect 4030 34193 4040 34245
rect 4083 34153 4117 34303
rect 4161 34193 4171 34245
rect 4223 34193 4233 34245
rect 4275 34153 4309 34303
rect 4352 34193 4362 34245
rect 4414 34193 4424 34245
rect 4467 34153 4501 34303
rect 4544 34193 4554 34245
rect 4606 34193 4616 34245
rect 4659 34153 4693 34303
rect 4736 34193 4746 34245
rect 4798 34193 4808 34245
rect 4851 34153 4885 34303
rect 4928 34193 4938 34245
rect 4990 34193 5000 34245
rect 5055 34209 5101 34414
rect 5055 34175 5061 34209
rect 5095 34175 5101 34209
rect 3981 34106 4027 34153
rect 3981 34072 3987 34106
rect 4021 34072 4027 34106
rect 3981 34034 4027 34072
rect 3981 34000 3987 34034
rect 4021 34000 4027 34034
rect 3981 33962 4027 34000
rect 3981 33928 3987 33962
rect 4021 33928 4027 33962
rect 3981 33881 4027 33928
rect 4077 34106 4123 34153
rect 4077 34072 4083 34106
rect 4117 34072 4123 34106
rect 4077 34034 4123 34072
rect 4077 34000 4083 34034
rect 4117 34000 4123 34034
rect 4077 33962 4123 34000
rect 4077 33928 4083 33962
rect 4117 33928 4123 33962
rect 4077 33881 4123 33928
rect 4173 34106 4219 34153
rect 4173 34072 4179 34106
rect 4213 34072 4219 34106
rect 4173 34034 4219 34072
rect 4173 34000 4179 34034
rect 4213 34000 4219 34034
rect 4173 33962 4219 34000
rect 4173 33928 4179 33962
rect 4213 33928 4219 33962
rect 4173 33881 4219 33928
rect 4269 34106 4315 34153
rect 4269 34072 4275 34106
rect 4309 34072 4315 34106
rect 4269 34034 4315 34072
rect 4269 34000 4275 34034
rect 4309 34000 4315 34034
rect 4269 33962 4315 34000
rect 4269 33928 4275 33962
rect 4309 33928 4315 33962
rect 4269 33881 4315 33928
rect 4365 34106 4411 34153
rect 4365 34072 4371 34106
rect 4405 34072 4411 34106
rect 4365 34034 4411 34072
rect 4365 34000 4371 34034
rect 4405 34000 4411 34034
rect 4365 33962 4411 34000
rect 4365 33928 4371 33962
rect 4405 33928 4411 33962
rect 4365 33881 4411 33928
rect 4461 34106 4507 34153
rect 4461 34072 4467 34106
rect 4501 34072 4507 34106
rect 4461 34034 4507 34072
rect 4461 34000 4467 34034
rect 4501 34000 4507 34034
rect 4461 33962 4507 34000
rect 4461 33928 4467 33962
rect 4501 33928 4507 33962
rect 4461 33881 4507 33928
rect 4557 34106 4603 34153
rect 4557 34072 4563 34106
rect 4597 34072 4603 34106
rect 4557 34034 4603 34072
rect 4557 34000 4563 34034
rect 4597 34000 4603 34034
rect 4557 33962 4603 34000
rect 4557 33928 4563 33962
rect 4597 33928 4603 33962
rect 4557 33881 4603 33928
rect 4653 34106 4699 34153
rect 4653 34072 4659 34106
rect 4693 34072 4699 34106
rect 4653 34034 4699 34072
rect 4653 34000 4659 34034
rect 4693 34000 4699 34034
rect 4653 33962 4699 34000
rect 4653 33928 4659 33962
rect 4693 33928 4699 33962
rect 4653 33881 4699 33928
rect 4749 34106 4795 34153
rect 4749 34072 4755 34106
rect 4789 34072 4795 34106
rect 4749 34034 4795 34072
rect 4749 34000 4755 34034
rect 4789 34000 4795 34034
rect 4749 33962 4795 34000
rect 4749 33928 4755 33962
rect 4789 33928 4795 33962
rect 4749 33881 4795 33928
rect 4845 34106 4891 34153
rect 4845 34072 4851 34106
rect 4885 34072 4891 34106
rect 4845 34034 4891 34072
rect 4845 34000 4851 34034
rect 4885 34000 4891 34034
rect 4845 33962 4891 34000
rect 4845 33928 4851 33962
rect 4885 33928 4891 33962
rect 4845 33881 4891 33928
rect 4941 34106 4987 34153
rect 4941 34072 4947 34106
rect 4981 34072 4987 34106
rect 4941 34034 4987 34072
rect 4941 34000 4947 34034
rect 4981 34000 4987 34034
rect 4941 33962 4987 34000
rect 4941 33928 4947 33962
rect 4981 33928 4987 33962
rect 4941 33881 4987 33928
rect 5055 34137 5101 34175
rect 5055 34103 5061 34137
rect 5095 34103 5101 34137
rect 5055 34065 5101 34103
rect 5055 34031 5061 34065
rect 5095 34034 5101 34065
rect 5274 34034 5550 34035
rect 5095 34031 5550 34034
rect 5055 34004 5550 34031
rect 5055 33993 5303 34004
rect 5055 33959 5061 33993
rect 5095 33970 5303 33993
rect 5337 33970 5395 34004
rect 5429 33970 5487 34004
rect 5521 33970 5550 34004
rect 5095 33959 5550 33970
rect 5055 33939 5550 33959
rect 5055 33921 5101 33939
rect 5055 33887 5061 33921
rect 5095 33887 5101 33921
rect 2466 33706 3837 33740
rect 2466 33573 2500 33706
rect 2658 33573 2692 33706
rect 2850 33573 2884 33706
rect 3042 33573 3076 33706
rect 3234 33573 3268 33706
rect 3426 33573 3460 33706
rect 3671 33616 3681 33668
rect 3733 33616 3743 33668
rect 3679 33615 3691 33616
rect 3725 33615 3737 33616
rect 3679 33609 3737 33615
rect 3534 33580 3580 33603
rect 2460 33538 2506 33573
rect 2460 33504 2466 33538
rect 2500 33504 2506 33538
rect 2460 33469 2506 33504
rect 2556 33538 2602 33573
rect 2556 33504 2562 33538
rect 2596 33504 2602 33538
rect 2556 33469 2602 33504
rect 2652 33538 2698 33573
rect 2652 33504 2658 33538
rect 2692 33504 2698 33538
rect 2652 33469 2698 33504
rect 2748 33538 2794 33573
rect 2748 33504 2754 33538
rect 2788 33504 2794 33538
rect 2748 33469 2794 33504
rect 2844 33538 2890 33573
rect 2844 33504 2850 33538
rect 2884 33504 2890 33538
rect 2844 33469 2890 33504
rect 2940 33538 2986 33573
rect 2940 33504 2946 33538
rect 2980 33504 2986 33538
rect 2940 33469 2986 33504
rect 3036 33538 3082 33573
rect 3036 33504 3042 33538
rect 3076 33504 3082 33538
rect 3036 33469 3082 33504
rect 3132 33538 3178 33573
rect 3132 33504 3138 33538
rect 3172 33504 3178 33538
rect 3132 33469 3178 33504
rect 3228 33538 3274 33573
rect 3228 33504 3234 33538
rect 3268 33504 3274 33538
rect 3228 33469 3274 33504
rect 3324 33538 3370 33573
rect 3324 33504 3330 33538
rect 3364 33504 3370 33538
rect 3324 33469 3370 33504
rect 3420 33538 3466 33573
rect 3420 33504 3426 33538
rect 3460 33504 3466 33538
rect 3420 33469 3466 33504
rect 3534 33546 3540 33580
rect 3574 33578 3580 33580
rect 3803 33578 3837 33706
rect 3574 33577 3680 33578
rect 3734 33577 3837 33578
rect 3574 33565 3687 33577
rect 3574 33546 3647 33565
rect 3534 33508 3647 33546
rect 3534 33474 3540 33508
rect 3574 33489 3647 33508
rect 3681 33489 3687 33565
rect 3574 33478 3687 33489
rect 3574 33474 3580 33478
rect 3641 33477 3687 33478
rect 3729 33565 3837 33577
rect 3987 33740 4021 33881
rect 4179 33740 4213 33881
rect 4371 33740 4405 33881
rect 4563 33740 4597 33881
rect 4755 33740 4789 33881
rect 4947 33740 4981 33881
rect 5055 33843 5101 33887
rect 5683 33794 5743 35047
rect 5177 33760 5743 33794
rect 5177 33740 5211 33760
rect 3987 33706 5211 33740
rect 3987 33573 4021 33706
rect 4179 33573 4213 33706
rect 4371 33573 4405 33706
rect 4563 33573 4597 33706
rect 4755 33573 4789 33706
rect 4947 33573 4981 33706
rect 5438 33702 5512 33703
rect 5326 33700 5400 33701
rect 5326 33648 5337 33700
rect 5389 33648 5400 33700
rect 5438 33650 5449 33702
rect 5501 33650 5512 33702
rect 5438 33649 5512 33650
rect 5326 33647 5400 33648
rect 5055 33580 5101 33603
rect 3729 33489 3735 33565
rect 3769 33489 3837 33565
rect 3729 33478 3837 33489
rect 3729 33477 3775 33478
rect 2450 33438 2516 33441
rect 2447 33386 2457 33438
rect 2509 33386 2519 33438
rect 2450 33381 2516 33386
rect 2562 33329 2596 33469
rect 2642 33438 2708 33441
rect 2638 33386 2648 33438
rect 2700 33386 2710 33438
rect 2642 33381 2708 33386
rect 2754 33329 2788 33469
rect 2834 33438 2900 33441
rect 2830 33386 2840 33438
rect 2892 33386 2902 33438
rect 2834 33381 2900 33386
rect 2946 33329 2980 33469
rect 3026 33438 3092 33441
rect 3022 33386 3032 33438
rect 3084 33386 3094 33438
rect 3026 33381 3092 33386
rect 3138 33329 3172 33469
rect 3218 33437 3284 33441
rect 3215 33385 3225 33437
rect 3277 33385 3287 33437
rect 3218 33381 3284 33385
rect 3330 33329 3364 33469
rect 3410 33437 3476 33441
rect 3407 33385 3417 33437
rect 3469 33385 3479 33437
rect 3534 33436 3580 33474
rect 3534 33402 3540 33436
rect 3574 33402 3580 33436
rect 3410 33381 3476 33385
rect 2282 33295 3364 33329
rect 3534 33219 3580 33402
rect 3803 33329 3837 33478
rect 3981 33538 4027 33573
rect 3981 33504 3987 33538
rect 4021 33504 4027 33538
rect 3981 33469 4027 33504
rect 4077 33538 4123 33573
rect 4077 33504 4083 33538
rect 4117 33504 4123 33538
rect 4077 33469 4123 33504
rect 4173 33538 4219 33573
rect 4173 33504 4179 33538
rect 4213 33504 4219 33538
rect 4173 33469 4219 33504
rect 4269 33538 4315 33573
rect 4269 33504 4275 33538
rect 4309 33504 4315 33538
rect 4269 33469 4315 33504
rect 4365 33538 4411 33573
rect 4365 33504 4371 33538
rect 4405 33504 4411 33538
rect 4365 33469 4411 33504
rect 4461 33538 4507 33573
rect 4461 33504 4467 33538
rect 4501 33504 4507 33538
rect 4461 33469 4507 33504
rect 4557 33538 4603 33573
rect 4557 33504 4563 33538
rect 4597 33504 4603 33538
rect 4557 33469 4603 33504
rect 4653 33538 4699 33573
rect 4653 33504 4659 33538
rect 4693 33504 4699 33538
rect 4653 33469 4699 33504
rect 4749 33538 4795 33573
rect 4749 33504 4755 33538
rect 4789 33504 4795 33538
rect 4749 33469 4795 33504
rect 4845 33538 4891 33573
rect 4845 33504 4851 33538
rect 4885 33504 4891 33538
rect 4845 33469 4891 33504
rect 4941 33538 4987 33573
rect 4941 33504 4947 33538
rect 4981 33504 4987 33538
rect 4941 33469 4987 33504
rect 5055 33546 5061 33580
rect 5095 33546 5101 33580
rect 5055 33508 5101 33546
rect 5055 33474 5061 33508
rect 5095 33491 5101 33508
rect 5095 33474 5550 33491
rect 3971 33438 4037 33441
rect 3968 33386 3978 33438
rect 4030 33386 4040 33438
rect 3971 33381 4037 33386
rect 4083 33329 4117 33469
rect 4163 33438 4229 33441
rect 4159 33386 4169 33438
rect 4221 33386 4231 33438
rect 4163 33381 4229 33386
rect 4275 33329 4309 33469
rect 4355 33438 4421 33441
rect 4351 33386 4361 33438
rect 4413 33386 4423 33438
rect 4355 33381 4421 33386
rect 4467 33329 4501 33469
rect 4547 33438 4613 33441
rect 4543 33386 4553 33438
rect 4605 33386 4615 33438
rect 4547 33381 4613 33386
rect 4659 33329 4693 33469
rect 4739 33437 4805 33441
rect 4736 33385 4746 33437
rect 4798 33385 4808 33437
rect 4739 33381 4805 33385
rect 4851 33329 4885 33469
rect 5055 33460 5550 33474
rect 4931 33437 4997 33441
rect 4928 33385 4938 33437
rect 4990 33385 5000 33437
rect 5055 33436 5303 33460
rect 5055 33402 5061 33436
rect 5095 33426 5303 33436
rect 5337 33426 5395 33460
rect 5429 33426 5487 33460
rect 5521 33426 5550 33460
rect 5095 33402 5550 33426
rect 5055 33395 5550 33402
rect 4931 33381 4997 33385
rect 3803 33295 4885 33329
rect 5055 33220 5101 33395
rect 129 33012 1211 33046
rect 129 32449 163 33012
rect 294 32902 304 32954
rect 356 32902 366 32954
rect 409 32862 443 33012
rect 487 32902 497 32954
rect 549 32902 559 32954
rect 601 32862 635 33012
rect 678 32902 688 32954
rect 740 32902 750 32954
rect 793 32862 827 33012
rect 870 32902 880 32954
rect 932 32902 942 32954
rect 985 32862 1019 33012
rect 1062 32902 1072 32954
rect 1124 32902 1134 32954
rect 1177 32862 1211 33012
rect 1254 32902 1264 32954
rect 1316 32902 1326 32954
rect 1381 32918 1427 33082
rect 2282 33016 3364 33050
rect 1381 32884 1387 32918
rect 1421 32884 1427 32918
rect 1512 32895 1522 32955
rect 1578 32895 1792 32955
rect 1852 32895 1862 32955
rect 307 32815 353 32862
rect 307 32781 313 32815
rect 347 32781 353 32815
rect 307 32743 353 32781
rect 307 32709 313 32743
rect 347 32709 353 32743
rect 307 32671 353 32709
rect 307 32637 313 32671
rect 347 32637 353 32671
rect 307 32590 353 32637
rect 403 32815 449 32862
rect 403 32781 409 32815
rect 443 32781 449 32815
rect 403 32743 449 32781
rect 403 32709 409 32743
rect 443 32709 449 32743
rect 403 32671 449 32709
rect 403 32637 409 32671
rect 443 32637 449 32671
rect 403 32590 449 32637
rect 499 32815 545 32862
rect 499 32781 505 32815
rect 539 32781 545 32815
rect 499 32743 545 32781
rect 499 32709 505 32743
rect 539 32709 545 32743
rect 499 32671 545 32709
rect 499 32637 505 32671
rect 539 32637 545 32671
rect 499 32590 545 32637
rect 595 32815 641 32862
rect 595 32781 601 32815
rect 635 32781 641 32815
rect 595 32743 641 32781
rect 595 32709 601 32743
rect 635 32709 641 32743
rect 595 32671 641 32709
rect 595 32637 601 32671
rect 635 32637 641 32671
rect 595 32590 641 32637
rect 691 32815 737 32862
rect 691 32781 697 32815
rect 731 32781 737 32815
rect 691 32743 737 32781
rect 691 32709 697 32743
rect 731 32709 737 32743
rect 691 32671 737 32709
rect 691 32637 697 32671
rect 731 32637 737 32671
rect 691 32590 737 32637
rect 787 32815 833 32862
rect 787 32781 793 32815
rect 827 32781 833 32815
rect 787 32743 833 32781
rect 787 32709 793 32743
rect 827 32709 833 32743
rect 787 32671 833 32709
rect 787 32637 793 32671
rect 827 32637 833 32671
rect 787 32590 833 32637
rect 883 32815 929 32862
rect 883 32781 889 32815
rect 923 32781 929 32815
rect 883 32743 929 32781
rect 883 32709 889 32743
rect 923 32709 929 32743
rect 883 32671 929 32709
rect 883 32637 889 32671
rect 923 32637 929 32671
rect 883 32590 929 32637
rect 979 32815 1025 32862
rect 979 32781 985 32815
rect 1019 32781 1025 32815
rect 979 32743 1025 32781
rect 979 32709 985 32743
rect 1019 32709 1025 32743
rect 979 32671 1025 32709
rect 979 32637 985 32671
rect 1019 32637 1025 32671
rect 979 32590 1025 32637
rect 1075 32815 1121 32862
rect 1075 32781 1081 32815
rect 1115 32781 1121 32815
rect 1075 32743 1121 32781
rect 1075 32709 1081 32743
rect 1115 32709 1121 32743
rect 1075 32671 1121 32709
rect 1075 32637 1081 32671
rect 1115 32637 1121 32671
rect 1075 32590 1121 32637
rect 1171 32815 1217 32862
rect 1171 32781 1177 32815
rect 1211 32781 1217 32815
rect 1171 32743 1217 32781
rect 1171 32709 1177 32743
rect 1211 32709 1217 32743
rect 1171 32671 1217 32709
rect 1171 32637 1177 32671
rect 1211 32637 1217 32671
rect 1171 32590 1217 32637
rect 1267 32815 1313 32862
rect 1267 32781 1273 32815
rect 1307 32781 1313 32815
rect 1267 32743 1313 32781
rect 1267 32709 1273 32743
rect 1307 32709 1313 32743
rect 1267 32671 1313 32709
rect 1267 32637 1273 32671
rect 1307 32637 1313 32671
rect 1267 32590 1313 32637
rect 1381 32846 1427 32884
rect 1381 32812 1387 32846
rect 1421 32812 1427 32846
rect 1381 32774 1427 32812
rect 1381 32740 1387 32774
rect 1421 32740 1427 32774
rect 1381 32702 1427 32740
rect 1381 32668 1387 32702
rect 1421 32668 1427 32702
rect 1381 32658 1427 32668
rect 1381 32656 2160 32658
rect 1381 32630 2056 32656
rect 1381 32605 1387 32630
rect 1380 32596 1387 32605
rect 1421 32596 2056 32630
rect 0 32415 163 32449
rect 129 32038 163 32415
rect 313 32449 347 32590
rect 505 32449 539 32590
rect 697 32449 731 32590
rect 889 32449 923 32590
rect 1081 32449 1115 32590
rect 1273 32449 1307 32590
rect 1380 32548 2056 32596
rect 2190 32548 2200 32656
rect 1380 32546 2160 32548
rect 2282 32453 2316 33016
rect 2447 32906 2457 32958
rect 2509 32906 2519 32958
rect 2562 32866 2596 33016
rect 2640 32906 2650 32958
rect 2702 32906 2712 32958
rect 2754 32866 2788 33016
rect 2831 32906 2841 32958
rect 2893 32906 2903 32958
rect 2946 32866 2980 33016
rect 3023 32906 3033 32958
rect 3085 32906 3095 32958
rect 3138 32866 3172 33016
rect 3215 32906 3225 32958
rect 3277 32906 3287 32958
rect 3330 32866 3364 33016
rect 3407 32906 3417 32958
rect 3469 32906 3479 32958
rect 3534 32922 3580 33130
rect 3534 32888 3540 32922
rect 3574 32888 3580 32922
rect 2460 32819 2506 32866
rect 2460 32785 2466 32819
rect 2500 32785 2506 32819
rect 2460 32747 2506 32785
rect 2460 32713 2466 32747
rect 2500 32713 2506 32747
rect 2460 32675 2506 32713
rect 2460 32641 2466 32675
rect 2500 32641 2506 32675
rect 2460 32594 2506 32641
rect 2556 32819 2602 32866
rect 2556 32785 2562 32819
rect 2596 32785 2602 32819
rect 2556 32747 2602 32785
rect 2556 32713 2562 32747
rect 2596 32713 2602 32747
rect 2556 32675 2602 32713
rect 2556 32641 2562 32675
rect 2596 32641 2602 32675
rect 2556 32594 2602 32641
rect 2652 32819 2698 32866
rect 2652 32785 2658 32819
rect 2692 32785 2698 32819
rect 2652 32747 2698 32785
rect 2652 32713 2658 32747
rect 2692 32713 2698 32747
rect 2652 32675 2698 32713
rect 2652 32641 2658 32675
rect 2692 32641 2698 32675
rect 2652 32594 2698 32641
rect 2748 32819 2794 32866
rect 2748 32785 2754 32819
rect 2788 32785 2794 32819
rect 2748 32747 2794 32785
rect 2748 32713 2754 32747
rect 2788 32713 2794 32747
rect 2748 32675 2794 32713
rect 2748 32641 2754 32675
rect 2788 32641 2794 32675
rect 2748 32594 2794 32641
rect 2844 32819 2890 32866
rect 2844 32785 2850 32819
rect 2884 32785 2890 32819
rect 2844 32747 2890 32785
rect 2844 32713 2850 32747
rect 2884 32713 2890 32747
rect 2844 32675 2890 32713
rect 2844 32641 2850 32675
rect 2884 32641 2890 32675
rect 2844 32594 2890 32641
rect 2940 32819 2986 32866
rect 2940 32785 2946 32819
rect 2980 32785 2986 32819
rect 2940 32747 2986 32785
rect 2940 32713 2946 32747
rect 2980 32713 2986 32747
rect 2940 32675 2986 32713
rect 2940 32641 2946 32675
rect 2980 32641 2986 32675
rect 2940 32594 2986 32641
rect 3036 32819 3082 32866
rect 3036 32785 3042 32819
rect 3076 32785 3082 32819
rect 3036 32747 3082 32785
rect 3036 32713 3042 32747
rect 3076 32713 3082 32747
rect 3036 32675 3082 32713
rect 3036 32641 3042 32675
rect 3076 32641 3082 32675
rect 3036 32594 3082 32641
rect 3132 32819 3178 32866
rect 3132 32785 3138 32819
rect 3172 32785 3178 32819
rect 3132 32747 3178 32785
rect 3132 32713 3138 32747
rect 3172 32713 3178 32747
rect 3132 32675 3178 32713
rect 3132 32641 3138 32675
rect 3172 32641 3178 32675
rect 3132 32594 3178 32641
rect 3228 32819 3274 32866
rect 3228 32785 3234 32819
rect 3268 32785 3274 32819
rect 3228 32747 3274 32785
rect 3228 32713 3234 32747
rect 3268 32713 3274 32747
rect 3228 32675 3274 32713
rect 3228 32641 3234 32675
rect 3268 32641 3274 32675
rect 3228 32594 3274 32641
rect 3324 32819 3370 32866
rect 3324 32785 3330 32819
rect 3364 32785 3370 32819
rect 3324 32747 3370 32785
rect 3324 32713 3330 32747
rect 3364 32713 3370 32747
rect 3324 32675 3370 32713
rect 3324 32641 3330 32675
rect 3364 32641 3370 32675
rect 3324 32594 3370 32641
rect 3420 32819 3466 32866
rect 3420 32785 3426 32819
rect 3460 32785 3466 32819
rect 3420 32747 3466 32785
rect 3420 32713 3426 32747
rect 3460 32713 3466 32747
rect 3420 32675 3466 32713
rect 3420 32641 3426 32675
rect 3460 32641 3466 32675
rect 3420 32594 3466 32641
rect 3534 32850 3580 32888
rect 3534 32816 3540 32850
rect 3574 32816 3580 32850
rect 3534 32778 3580 32816
rect 3534 32744 3540 32778
rect 3574 32744 3580 32778
rect 3534 32706 3580 32744
rect 3534 32672 3540 32706
rect 3574 32672 3580 32706
rect 3534 32634 3580 32672
rect 3534 32600 3540 32634
rect 3574 32600 3580 32634
rect 2101 32449 2316 32453
rect 313 32419 2316 32449
rect 313 32415 2141 32419
rect 313 32282 347 32415
rect 505 32282 539 32415
rect 697 32282 731 32415
rect 889 32282 923 32415
rect 1081 32282 1115 32415
rect 1273 32282 1307 32415
rect 1381 32289 1608 32312
rect 307 32247 353 32282
rect 307 32213 313 32247
rect 347 32213 353 32247
rect 307 32178 353 32213
rect 403 32247 449 32282
rect 403 32213 409 32247
rect 443 32213 449 32247
rect 403 32178 449 32213
rect 499 32247 545 32282
rect 499 32213 505 32247
rect 539 32213 545 32247
rect 499 32178 545 32213
rect 595 32247 641 32282
rect 595 32213 601 32247
rect 635 32213 641 32247
rect 595 32178 641 32213
rect 691 32247 737 32282
rect 691 32213 697 32247
rect 731 32213 737 32247
rect 691 32178 737 32213
rect 787 32247 833 32282
rect 787 32213 793 32247
rect 827 32213 833 32247
rect 787 32178 833 32213
rect 883 32247 929 32282
rect 883 32213 889 32247
rect 923 32213 929 32247
rect 883 32178 929 32213
rect 979 32247 1025 32282
rect 979 32213 985 32247
rect 1019 32213 1025 32247
rect 979 32178 1025 32213
rect 1075 32247 1121 32282
rect 1075 32213 1081 32247
rect 1115 32213 1121 32247
rect 1075 32178 1121 32213
rect 1171 32247 1217 32282
rect 1171 32213 1177 32247
rect 1211 32213 1217 32247
rect 1171 32178 1217 32213
rect 1267 32247 1313 32282
rect 1267 32213 1273 32247
rect 1307 32213 1313 32247
rect 1267 32178 1313 32213
rect 1381 32255 1387 32289
rect 1421 32255 1608 32289
rect 1381 32217 1608 32255
rect 1381 32183 1387 32217
rect 1421 32192 1608 32217
rect 1421 32183 1427 32192
rect 1560 32190 1608 32192
rect 1598 32188 1608 32190
rect 1720 32188 1730 32312
rect 297 32147 363 32150
rect 294 32095 304 32147
rect 356 32095 366 32147
rect 297 32090 363 32095
rect 409 32038 443 32178
rect 489 32147 555 32150
rect 485 32095 495 32147
rect 547 32095 557 32147
rect 489 32090 555 32095
rect 601 32038 635 32178
rect 681 32147 747 32150
rect 677 32095 687 32147
rect 739 32095 749 32147
rect 681 32090 747 32095
rect 793 32038 827 32178
rect 873 32147 939 32150
rect 869 32095 879 32147
rect 931 32095 941 32147
rect 873 32090 939 32095
rect 985 32038 1019 32178
rect 1065 32146 1131 32150
rect 1062 32094 1072 32146
rect 1124 32094 1134 32146
rect 1065 32090 1131 32094
rect 1177 32038 1211 32178
rect 1257 32146 1323 32150
rect 1254 32094 1264 32146
rect 1316 32094 1326 32146
rect 1381 32145 1427 32183
rect 1920 32150 1930 32152
rect 1381 32111 1387 32145
rect 1421 32111 1427 32145
rect 1257 32090 1323 32094
rect 129 32004 1211 32038
rect 1381 31968 1427 32111
rect 1458 32094 1468 32150
rect 1524 32096 1930 32150
rect 1986 32096 1996 32152
rect 1524 32094 1986 32096
rect 2282 32042 2316 32419
rect 2466 32453 2500 32594
rect 2658 32453 2692 32594
rect 2850 32453 2884 32594
rect 3042 32453 3076 32594
rect 3234 32453 3268 32594
rect 3426 32453 3460 32594
rect 3534 32556 3580 32600
rect 3803 33016 4885 33050
rect 3803 32453 3837 33016
rect 3968 32906 3978 32958
rect 4030 32906 4040 32958
rect 4083 32866 4117 33016
rect 4161 32906 4171 32958
rect 4223 32906 4233 32958
rect 4275 32866 4309 33016
rect 4352 32906 4362 32958
rect 4414 32906 4424 32958
rect 4467 32866 4501 33016
rect 4544 32906 4554 32958
rect 4606 32906 4616 32958
rect 4659 32866 4693 33016
rect 4736 32906 4746 32958
rect 4798 32906 4808 32958
rect 4851 32866 4885 33016
rect 4928 32906 4938 32958
rect 4990 32906 5000 32958
rect 5055 32922 5101 33127
rect 5055 32888 5061 32922
rect 5095 32888 5101 32922
rect 3981 32819 4027 32866
rect 3981 32785 3987 32819
rect 4021 32785 4027 32819
rect 3981 32747 4027 32785
rect 3981 32713 3987 32747
rect 4021 32713 4027 32747
rect 3981 32675 4027 32713
rect 3981 32641 3987 32675
rect 4021 32641 4027 32675
rect 3981 32594 4027 32641
rect 4077 32819 4123 32866
rect 4077 32785 4083 32819
rect 4117 32785 4123 32819
rect 4077 32747 4123 32785
rect 4077 32713 4083 32747
rect 4117 32713 4123 32747
rect 4077 32675 4123 32713
rect 4077 32641 4083 32675
rect 4117 32641 4123 32675
rect 4077 32594 4123 32641
rect 4173 32819 4219 32866
rect 4173 32785 4179 32819
rect 4213 32785 4219 32819
rect 4173 32747 4219 32785
rect 4173 32713 4179 32747
rect 4213 32713 4219 32747
rect 4173 32675 4219 32713
rect 4173 32641 4179 32675
rect 4213 32641 4219 32675
rect 4173 32594 4219 32641
rect 4269 32819 4315 32866
rect 4269 32785 4275 32819
rect 4309 32785 4315 32819
rect 4269 32747 4315 32785
rect 4269 32713 4275 32747
rect 4309 32713 4315 32747
rect 4269 32675 4315 32713
rect 4269 32641 4275 32675
rect 4309 32641 4315 32675
rect 4269 32594 4315 32641
rect 4365 32819 4411 32866
rect 4365 32785 4371 32819
rect 4405 32785 4411 32819
rect 4365 32747 4411 32785
rect 4365 32713 4371 32747
rect 4405 32713 4411 32747
rect 4365 32675 4411 32713
rect 4365 32641 4371 32675
rect 4405 32641 4411 32675
rect 4365 32594 4411 32641
rect 4461 32819 4507 32866
rect 4461 32785 4467 32819
rect 4501 32785 4507 32819
rect 4461 32747 4507 32785
rect 4461 32713 4467 32747
rect 4501 32713 4507 32747
rect 4461 32675 4507 32713
rect 4461 32641 4467 32675
rect 4501 32641 4507 32675
rect 4461 32594 4507 32641
rect 4557 32819 4603 32866
rect 4557 32785 4563 32819
rect 4597 32785 4603 32819
rect 4557 32747 4603 32785
rect 4557 32713 4563 32747
rect 4597 32713 4603 32747
rect 4557 32675 4603 32713
rect 4557 32641 4563 32675
rect 4597 32641 4603 32675
rect 4557 32594 4603 32641
rect 4653 32819 4699 32866
rect 4653 32785 4659 32819
rect 4693 32785 4699 32819
rect 4653 32747 4699 32785
rect 4653 32713 4659 32747
rect 4693 32713 4699 32747
rect 4653 32675 4699 32713
rect 4653 32641 4659 32675
rect 4693 32641 4699 32675
rect 4653 32594 4699 32641
rect 4749 32819 4795 32866
rect 4749 32785 4755 32819
rect 4789 32785 4795 32819
rect 4749 32747 4795 32785
rect 4749 32713 4755 32747
rect 4789 32713 4795 32747
rect 4749 32675 4795 32713
rect 4749 32641 4755 32675
rect 4789 32641 4795 32675
rect 4749 32594 4795 32641
rect 4845 32819 4891 32866
rect 4845 32785 4851 32819
rect 4885 32785 4891 32819
rect 4845 32747 4891 32785
rect 4845 32713 4851 32747
rect 4885 32713 4891 32747
rect 4845 32675 4891 32713
rect 4845 32641 4851 32675
rect 4885 32641 4891 32675
rect 4845 32594 4891 32641
rect 4941 32819 4987 32866
rect 4941 32785 4947 32819
rect 4981 32785 4987 32819
rect 4941 32747 4987 32785
rect 4941 32713 4947 32747
rect 4981 32713 4987 32747
rect 4941 32675 4987 32713
rect 4941 32641 4947 32675
rect 4981 32641 4987 32675
rect 4941 32594 4987 32641
rect 5055 32850 5101 32888
rect 5055 32816 5061 32850
rect 5095 32816 5101 32850
rect 5055 32778 5101 32816
rect 5055 32744 5061 32778
rect 5095 32747 5101 32778
rect 5274 32747 5550 32748
rect 5095 32744 5550 32747
rect 5055 32717 5550 32744
rect 5055 32706 5303 32717
rect 5055 32672 5061 32706
rect 5095 32683 5303 32706
rect 5337 32683 5395 32717
rect 5429 32683 5487 32717
rect 5521 32683 5550 32717
rect 5095 32672 5550 32683
rect 5055 32652 5550 32672
rect 5055 32634 5101 32652
rect 5055 32600 5061 32634
rect 5095 32600 5101 32634
rect 2466 32419 3837 32453
rect 2466 32286 2500 32419
rect 2658 32286 2692 32419
rect 2850 32286 2884 32419
rect 3042 32286 3076 32419
rect 3234 32286 3268 32419
rect 3426 32286 3460 32419
rect 3671 32329 3681 32381
rect 3733 32329 3743 32381
rect 3679 32328 3691 32329
rect 3725 32328 3737 32329
rect 3679 32322 3737 32328
rect 3534 32293 3580 32316
rect 2460 32251 2506 32286
rect 2460 32217 2466 32251
rect 2500 32217 2506 32251
rect 2460 32182 2506 32217
rect 2556 32251 2602 32286
rect 2556 32217 2562 32251
rect 2596 32217 2602 32251
rect 2556 32182 2602 32217
rect 2652 32251 2698 32286
rect 2652 32217 2658 32251
rect 2692 32217 2698 32251
rect 2652 32182 2698 32217
rect 2748 32251 2794 32286
rect 2748 32217 2754 32251
rect 2788 32217 2794 32251
rect 2748 32182 2794 32217
rect 2844 32251 2890 32286
rect 2844 32217 2850 32251
rect 2884 32217 2890 32251
rect 2844 32182 2890 32217
rect 2940 32251 2986 32286
rect 2940 32217 2946 32251
rect 2980 32217 2986 32251
rect 2940 32182 2986 32217
rect 3036 32251 3082 32286
rect 3036 32217 3042 32251
rect 3076 32217 3082 32251
rect 3036 32182 3082 32217
rect 3132 32251 3178 32286
rect 3132 32217 3138 32251
rect 3172 32217 3178 32251
rect 3132 32182 3178 32217
rect 3228 32251 3274 32286
rect 3228 32217 3234 32251
rect 3268 32217 3274 32251
rect 3228 32182 3274 32217
rect 3324 32251 3370 32286
rect 3324 32217 3330 32251
rect 3364 32217 3370 32251
rect 3324 32182 3370 32217
rect 3420 32251 3466 32286
rect 3420 32217 3426 32251
rect 3460 32217 3466 32251
rect 3420 32182 3466 32217
rect 3534 32259 3540 32293
rect 3574 32291 3580 32293
rect 3803 32291 3837 32419
rect 3574 32290 3680 32291
rect 3734 32290 3837 32291
rect 3574 32278 3687 32290
rect 3574 32259 3647 32278
rect 3534 32221 3647 32259
rect 3534 32187 3540 32221
rect 3574 32202 3647 32221
rect 3681 32202 3687 32278
rect 3574 32191 3687 32202
rect 3574 32187 3580 32191
rect 3641 32190 3687 32191
rect 3729 32278 3837 32290
rect 3987 32453 4021 32594
rect 4179 32453 4213 32594
rect 4371 32453 4405 32594
rect 4563 32453 4597 32594
rect 4755 32453 4789 32594
rect 4947 32453 4981 32594
rect 5055 32556 5101 32600
rect 5683 32507 5743 33760
rect 5177 32473 5743 32507
rect 5177 32453 5211 32473
rect 3987 32419 5211 32453
rect 3987 32286 4021 32419
rect 4179 32286 4213 32419
rect 4371 32286 4405 32419
rect 4563 32286 4597 32419
rect 4755 32286 4789 32419
rect 4947 32286 4981 32419
rect 5438 32415 5512 32416
rect 5326 32413 5400 32414
rect 5326 32361 5337 32413
rect 5389 32361 5400 32413
rect 5438 32363 5449 32415
rect 5501 32363 5512 32415
rect 5438 32362 5512 32363
rect 5326 32360 5400 32361
rect 5055 32293 5101 32316
rect 3729 32202 3735 32278
rect 3769 32202 3837 32278
rect 3729 32191 3837 32202
rect 3729 32190 3775 32191
rect 2450 32151 2516 32154
rect 2447 32099 2457 32151
rect 2509 32099 2519 32151
rect 2450 32094 2516 32099
rect 2562 32042 2596 32182
rect 2642 32151 2708 32154
rect 2638 32099 2648 32151
rect 2700 32099 2710 32151
rect 2642 32094 2708 32099
rect 2754 32042 2788 32182
rect 2834 32151 2900 32154
rect 2830 32099 2840 32151
rect 2892 32099 2902 32151
rect 2834 32094 2900 32099
rect 2946 32042 2980 32182
rect 3026 32151 3092 32154
rect 3022 32099 3032 32151
rect 3084 32099 3094 32151
rect 3026 32094 3092 32099
rect 3138 32042 3172 32182
rect 3218 32150 3284 32154
rect 3215 32098 3225 32150
rect 3277 32098 3287 32150
rect 3218 32094 3284 32098
rect 3330 32042 3364 32182
rect 3410 32150 3476 32154
rect 3407 32098 3417 32150
rect 3469 32098 3479 32150
rect 3534 32149 3580 32187
rect 3534 32115 3540 32149
rect 3574 32115 3580 32149
rect 3410 32094 3476 32098
rect 2282 32008 3364 32042
rect 3534 31932 3580 32115
rect 3803 32042 3837 32191
rect 3981 32251 4027 32286
rect 3981 32217 3987 32251
rect 4021 32217 4027 32251
rect 3981 32182 4027 32217
rect 4077 32251 4123 32286
rect 4077 32217 4083 32251
rect 4117 32217 4123 32251
rect 4077 32182 4123 32217
rect 4173 32251 4219 32286
rect 4173 32217 4179 32251
rect 4213 32217 4219 32251
rect 4173 32182 4219 32217
rect 4269 32251 4315 32286
rect 4269 32217 4275 32251
rect 4309 32217 4315 32251
rect 4269 32182 4315 32217
rect 4365 32251 4411 32286
rect 4365 32217 4371 32251
rect 4405 32217 4411 32251
rect 4365 32182 4411 32217
rect 4461 32251 4507 32286
rect 4461 32217 4467 32251
rect 4501 32217 4507 32251
rect 4461 32182 4507 32217
rect 4557 32251 4603 32286
rect 4557 32217 4563 32251
rect 4597 32217 4603 32251
rect 4557 32182 4603 32217
rect 4653 32251 4699 32286
rect 4653 32217 4659 32251
rect 4693 32217 4699 32251
rect 4653 32182 4699 32217
rect 4749 32251 4795 32286
rect 4749 32217 4755 32251
rect 4789 32217 4795 32251
rect 4749 32182 4795 32217
rect 4845 32251 4891 32286
rect 4845 32217 4851 32251
rect 4885 32217 4891 32251
rect 4845 32182 4891 32217
rect 4941 32251 4987 32286
rect 4941 32217 4947 32251
rect 4981 32217 4987 32251
rect 4941 32182 4987 32217
rect 5055 32259 5061 32293
rect 5095 32259 5101 32293
rect 5055 32221 5101 32259
rect 5055 32187 5061 32221
rect 5095 32204 5101 32221
rect 5095 32187 5550 32204
rect 3971 32151 4037 32154
rect 3968 32099 3978 32151
rect 4030 32099 4040 32151
rect 3971 32094 4037 32099
rect 4083 32042 4117 32182
rect 4163 32151 4229 32154
rect 4159 32099 4169 32151
rect 4221 32099 4231 32151
rect 4163 32094 4229 32099
rect 4275 32042 4309 32182
rect 4355 32151 4421 32154
rect 4351 32099 4361 32151
rect 4413 32099 4423 32151
rect 4355 32094 4421 32099
rect 4467 32042 4501 32182
rect 4547 32151 4613 32154
rect 4543 32099 4553 32151
rect 4605 32099 4615 32151
rect 4547 32094 4613 32099
rect 4659 32042 4693 32182
rect 4739 32150 4805 32154
rect 4736 32098 4746 32150
rect 4798 32098 4808 32150
rect 4739 32094 4805 32098
rect 4851 32042 4885 32182
rect 5055 32173 5550 32187
rect 4931 32150 4997 32154
rect 4928 32098 4938 32150
rect 4990 32098 5000 32150
rect 5055 32149 5303 32173
rect 5055 32115 5061 32149
rect 5095 32139 5303 32149
rect 5337 32139 5395 32173
rect 5429 32139 5487 32173
rect 5521 32139 5550 32173
rect 5095 32115 5550 32139
rect 5055 32108 5550 32115
rect 4931 32094 4997 32098
rect 3803 32008 4885 32042
rect 5055 31933 5101 32108
rect 129 31725 1211 31759
rect 129 31162 163 31725
rect 294 31615 304 31667
rect 356 31615 366 31667
rect 409 31575 443 31725
rect 487 31615 497 31667
rect 549 31615 559 31667
rect 601 31575 635 31725
rect 678 31615 688 31667
rect 740 31615 750 31667
rect 793 31575 827 31725
rect 870 31615 880 31667
rect 932 31615 942 31667
rect 985 31575 1019 31725
rect 1062 31615 1072 31667
rect 1124 31615 1134 31667
rect 1177 31575 1211 31725
rect 1254 31615 1264 31667
rect 1316 31615 1326 31667
rect 1381 31631 1427 31795
rect 2282 31729 3364 31763
rect 1381 31597 1387 31631
rect 1421 31597 1427 31631
rect 1512 31608 1522 31668
rect 1578 31608 1792 31668
rect 1852 31608 1862 31668
rect 307 31528 353 31575
rect 307 31494 313 31528
rect 347 31494 353 31528
rect 307 31456 353 31494
rect 307 31422 313 31456
rect 347 31422 353 31456
rect 307 31384 353 31422
rect 307 31350 313 31384
rect 347 31350 353 31384
rect 307 31303 353 31350
rect 403 31528 449 31575
rect 403 31494 409 31528
rect 443 31494 449 31528
rect 403 31456 449 31494
rect 403 31422 409 31456
rect 443 31422 449 31456
rect 403 31384 449 31422
rect 403 31350 409 31384
rect 443 31350 449 31384
rect 403 31303 449 31350
rect 499 31528 545 31575
rect 499 31494 505 31528
rect 539 31494 545 31528
rect 499 31456 545 31494
rect 499 31422 505 31456
rect 539 31422 545 31456
rect 499 31384 545 31422
rect 499 31350 505 31384
rect 539 31350 545 31384
rect 499 31303 545 31350
rect 595 31528 641 31575
rect 595 31494 601 31528
rect 635 31494 641 31528
rect 595 31456 641 31494
rect 595 31422 601 31456
rect 635 31422 641 31456
rect 595 31384 641 31422
rect 595 31350 601 31384
rect 635 31350 641 31384
rect 595 31303 641 31350
rect 691 31528 737 31575
rect 691 31494 697 31528
rect 731 31494 737 31528
rect 691 31456 737 31494
rect 691 31422 697 31456
rect 731 31422 737 31456
rect 691 31384 737 31422
rect 691 31350 697 31384
rect 731 31350 737 31384
rect 691 31303 737 31350
rect 787 31528 833 31575
rect 787 31494 793 31528
rect 827 31494 833 31528
rect 787 31456 833 31494
rect 787 31422 793 31456
rect 827 31422 833 31456
rect 787 31384 833 31422
rect 787 31350 793 31384
rect 827 31350 833 31384
rect 787 31303 833 31350
rect 883 31528 929 31575
rect 883 31494 889 31528
rect 923 31494 929 31528
rect 883 31456 929 31494
rect 883 31422 889 31456
rect 923 31422 929 31456
rect 883 31384 929 31422
rect 883 31350 889 31384
rect 923 31350 929 31384
rect 883 31303 929 31350
rect 979 31528 1025 31575
rect 979 31494 985 31528
rect 1019 31494 1025 31528
rect 979 31456 1025 31494
rect 979 31422 985 31456
rect 1019 31422 1025 31456
rect 979 31384 1025 31422
rect 979 31350 985 31384
rect 1019 31350 1025 31384
rect 979 31303 1025 31350
rect 1075 31528 1121 31575
rect 1075 31494 1081 31528
rect 1115 31494 1121 31528
rect 1075 31456 1121 31494
rect 1075 31422 1081 31456
rect 1115 31422 1121 31456
rect 1075 31384 1121 31422
rect 1075 31350 1081 31384
rect 1115 31350 1121 31384
rect 1075 31303 1121 31350
rect 1171 31528 1217 31575
rect 1171 31494 1177 31528
rect 1211 31494 1217 31528
rect 1171 31456 1217 31494
rect 1171 31422 1177 31456
rect 1211 31422 1217 31456
rect 1171 31384 1217 31422
rect 1171 31350 1177 31384
rect 1211 31350 1217 31384
rect 1171 31303 1217 31350
rect 1267 31528 1313 31575
rect 1267 31494 1273 31528
rect 1307 31494 1313 31528
rect 1267 31456 1313 31494
rect 1267 31422 1273 31456
rect 1307 31422 1313 31456
rect 1267 31384 1313 31422
rect 1267 31350 1273 31384
rect 1307 31350 1313 31384
rect 1267 31303 1313 31350
rect 1381 31559 1427 31597
rect 1381 31525 1387 31559
rect 1421 31525 1427 31559
rect 1381 31487 1427 31525
rect 1381 31453 1387 31487
rect 1421 31453 1427 31487
rect 1381 31415 1427 31453
rect 1381 31381 1387 31415
rect 1421 31381 1427 31415
rect 1381 31371 1427 31381
rect 1381 31369 2160 31371
rect 1381 31343 2056 31369
rect 1381 31318 1387 31343
rect 1380 31309 1387 31318
rect 1421 31309 2056 31343
rect 0 31128 163 31162
rect 129 30751 163 31128
rect 313 31162 347 31303
rect 505 31162 539 31303
rect 697 31162 731 31303
rect 889 31162 923 31303
rect 1081 31162 1115 31303
rect 1273 31162 1307 31303
rect 1380 31261 2056 31309
rect 2190 31261 2200 31369
rect 1380 31259 2160 31261
rect 2282 31166 2316 31729
rect 2447 31619 2457 31671
rect 2509 31619 2519 31671
rect 2562 31579 2596 31729
rect 2640 31619 2650 31671
rect 2702 31619 2712 31671
rect 2754 31579 2788 31729
rect 2831 31619 2841 31671
rect 2893 31619 2903 31671
rect 2946 31579 2980 31729
rect 3023 31619 3033 31671
rect 3085 31619 3095 31671
rect 3138 31579 3172 31729
rect 3215 31619 3225 31671
rect 3277 31619 3287 31671
rect 3330 31579 3364 31729
rect 3407 31619 3417 31671
rect 3469 31619 3479 31671
rect 3534 31635 3580 31843
rect 3534 31601 3540 31635
rect 3574 31601 3580 31635
rect 2460 31532 2506 31579
rect 2460 31498 2466 31532
rect 2500 31498 2506 31532
rect 2460 31460 2506 31498
rect 2460 31426 2466 31460
rect 2500 31426 2506 31460
rect 2460 31388 2506 31426
rect 2460 31354 2466 31388
rect 2500 31354 2506 31388
rect 2460 31307 2506 31354
rect 2556 31532 2602 31579
rect 2556 31498 2562 31532
rect 2596 31498 2602 31532
rect 2556 31460 2602 31498
rect 2556 31426 2562 31460
rect 2596 31426 2602 31460
rect 2556 31388 2602 31426
rect 2556 31354 2562 31388
rect 2596 31354 2602 31388
rect 2556 31307 2602 31354
rect 2652 31532 2698 31579
rect 2652 31498 2658 31532
rect 2692 31498 2698 31532
rect 2652 31460 2698 31498
rect 2652 31426 2658 31460
rect 2692 31426 2698 31460
rect 2652 31388 2698 31426
rect 2652 31354 2658 31388
rect 2692 31354 2698 31388
rect 2652 31307 2698 31354
rect 2748 31532 2794 31579
rect 2748 31498 2754 31532
rect 2788 31498 2794 31532
rect 2748 31460 2794 31498
rect 2748 31426 2754 31460
rect 2788 31426 2794 31460
rect 2748 31388 2794 31426
rect 2748 31354 2754 31388
rect 2788 31354 2794 31388
rect 2748 31307 2794 31354
rect 2844 31532 2890 31579
rect 2844 31498 2850 31532
rect 2884 31498 2890 31532
rect 2844 31460 2890 31498
rect 2844 31426 2850 31460
rect 2884 31426 2890 31460
rect 2844 31388 2890 31426
rect 2844 31354 2850 31388
rect 2884 31354 2890 31388
rect 2844 31307 2890 31354
rect 2940 31532 2986 31579
rect 2940 31498 2946 31532
rect 2980 31498 2986 31532
rect 2940 31460 2986 31498
rect 2940 31426 2946 31460
rect 2980 31426 2986 31460
rect 2940 31388 2986 31426
rect 2940 31354 2946 31388
rect 2980 31354 2986 31388
rect 2940 31307 2986 31354
rect 3036 31532 3082 31579
rect 3036 31498 3042 31532
rect 3076 31498 3082 31532
rect 3036 31460 3082 31498
rect 3036 31426 3042 31460
rect 3076 31426 3082 31460
rect 3036 31388 3082 31426
rect 3036 31354 3042 31388
rect 3076 31354 3082 31388
rect 3036 31307 3082 31354
rect 3132 31532 3178 31579
rect 3132 31498 3138 31532
rect 3172 31498 3178 31532
rect 3132 31460 3178 31498
rect 3132 31426 3138 31460
rect 3172 31426 3178 31460
rect 3132 31388 3178 31426
rect 3132 31354 3138 31388
rect 3172 31354 3178 31388
rect 3132 31307 3178 31354
rect 3228 31532 3274 31579
rect 3228 31498 3234 31532
rect 3268 31498 3274 31532
rect 3228 31460 3274 31498
rect 3228 31426 3234 31460
rect 3268 31426 3274 31460
rect 3228 31388 3274 31426
rect 3228 31354 3234 31388
rect 3268 31354 3274 31388
rect 3228 31307 3274 31354
rect 3324 31532 3370 31579
rect 3324 31498 3330 31532
rect 3364 31498 3370 31532
rect 3324 31460 3370 31498
rect 3324 31426 3330 31460
rect 3364 31426 3370 31460
rect 3324 31388 3370 31426
rect 3324 31354 3330 31388
rect 3364 31354 3370 31388
rect 3324 31307 3370 31354
rect 3420 31532 3466 31579
rect 3420 31498 3426 31532
rect 3460 31498 3466 31532
rect 3420 31460 3466 31498
rect 3420 31426 3426 31460
rect 3460 31426 3466 31460
rect 3420 31388 3466 31426
rect 3420 31354 3426 31388
rect 3460 31354 3466 31388
rect 3420 31307 3466 31354
rect 3534 31563 3580 31601
rect 3534 31529 3540 31563
rect 3574 31529 3580 31563
rect 3534 31491 3580 31529
rect 3534 31457 3540 31491
rect 3574 31457 3580 31491
rect 3534 31419 3580 31457
rect 3534 31385 3540 31419
rect 3574 31385 3580 31419
rect 3534 31347 3580 31385
rect 3534 31313 3540 31347
rect 3574 31313 3580 31347
rect 2101 31162 2316 31166
rect 313 31132 2316 31162
rect 313 31128 2141 31132
rect 313 30995 347 31128
rect 505 30995 539 31128
rect 697 30995 731 31128
rect 889 30995 923 31128
rect 1081 30995 1115 31128
rect 1273 30995 1307 31128
rect 1381 31002 1608 31025
rect 307 30960 353 30995
rect 307 30926 313 30960
rect 347 30926 353 30960
rect 307 30891 353 30926
rect 403 30960 449 30995
rect 403 30926 409 30960
rect 443 30926 449 30960
rect 403 30891 449 30926
rect 499 30960 545 30995
rect 499 30926 505 30960
rect 539 30926 545 30960
rect 499 30891 545 30926
rect 595 30960 641 30995
rect 595 30926 601 30960
rect 635 30926 641 30960
rect 595 30891 641 30926
rect 691 30960 737 30995
rect 691 30926 697 30960
rect 731 30926 737 30960
rect 691 30891 737 30926
rect 787 30960 833 30995
rect 787 30926 793 30960
rect 827 30926 833 30960
rect 787 30891 833 30926
rect 883 30960 929 30995
rect 883 30926 889 30960
rect 923 30926 929 30960
rect 883 30891 929 30926
rect 979 30960 1025 30995
rect 979 30926 985 30960
rect 1019 30926 1025 30960
rect 979 30891 1025 30926
rect 1075 30960 1121 30995
rect 1075 30926 1081 30960
rect 1115 30926 1121 30960
rect 1075 30891 1121 30926
rect 1171 30960 1217 30995
rect 1171 30926 1177 30960
rect 1211 30926 1217 30960
rect 1171 30891 1217 30926
rect 1267 30960 1313 30995
rect 1267 30926 1273 30960
rect 1307 30926 1313 30960
rect 1267 30891 1313 30926
rect 1381 30968 1387 31002
rect 1421 30968 1608 31002
rect 1381 30930 1608 30968
rect 1381 30896 1387 30930
rect 1421 30905 1608 30930
rect 1421 30896 1427 30905
rect 1560 30903 1608 30905
rect 1598 30901 1608 30903
rect 1720 30901 1730 31025
rect 297 30860 363 30863
rect 294 30808 304 30860
rect 356 30808 366 30860
rect 297 30803 363 30808
rect 409 30751 443 30891
rect 489 30860 555 30863
rect 485 30808 495 30860
rect 547 30808 557 30860
rect 489 30803 555 30808
rect 601 30751 635 30891
rect 681 30860 747 30863
rect 677 30808 687 30860
rect 739 30808 749 30860
rect 681 30803 747 30808
rect 793 30751 827 30891
rect 873 30860 939 30863
rect 869 30808 879 30860
rect 931 30808 941 30860
rect 873 30803 939 30808
rect 985 30751 1019 30891
rect 1065 30859 1131 30863
rect 1062 30807 1072 30859
rect 1124 30807 1134 30859
rect 1065 30803 1131 30807
rect 1177 30751 1211 30891
rect 1257 30859 1323 30863
rect 1254 30807 1264 30859
rect 1316 30807 1326 30859
rect 1381 30858 1427 30896
rect 1920 30863 1930 30865
rect 1381 30824 1387 30858
rect 1421 30824 1427 30858
rect 1257 30803 1323 30807
rect 129 30717 1211 30751
rect 1381 30681 1427 30824
rect 1458 30807 1468 30863
rect 1524 30809 1930 30863
rect 1986 30809 1996 30865
rect 1524 30807 1986 30809
rect 2282 30755 2316 31132
rect 2466 31166 2500 31307
rect 2658 31166 2692 31307
rect 2850 31166 2884 31307
rect 3042 31166 3076 31307
rect 3234 31166 3268 31307
rect 3426 31166 3460 31307
rect 3534 31269 3580 31313
rect 3803 31729 4885 31763
rect 3803 31166 3837 31729
rect 3968 31619 3978 31671
rect 4030 31619 4040 31671
rect 4083 31579 4117 31729
rect 4161 31619 4171 31671
rect 4223 31619 4233 31671
rect 4275 31579 4309 31729
rect 4352 31619 4362 31671
rect 4414 31619 4424 31671
rect 4467 31579 4501 31729
rect 4544 31619 4554 31671
rect 4606 31619 4616 31671
rect 4659 31579 4693 31729
rect 4736 31619 4746 31671
rect 4798 31619 4808 31671
rect 4851 31579 4885 31729
rect 4928 31619 4938 31671
rect 4990 31619 5000 31671
rect 5055 31635 5101 31840
rect 5055 31601 5061 31635
rect 5095 31601 5101 31635
rect 3981 31532 4027 31579
rect 3981 31498 3987 31532
rect 4021 31498 4027 31532
rect 3981 31460 4027 31498
rect 3981 31426 3987 31460
rect 4021 31426 4027 31460
rect 3981 31388 4027 31426
rect 3981 31354 3987 31388
rect 4021 31354 4027 31388
rect 3981 31307 4027 31354
rect 4077 31532 4123 31579
rect 4077 31498 4083 31532
rect 4117 31498 4123 31532
rect 4077 31460 4123 31498
rect 4077 31426 4083 31460
rect 4117 31426 4123 31460
rect 4077 31388 4123 31426
rect 4077 31354 4083 31388
rect 4117 31354 4123 31388
rect 4077 31307 4123 31354
rect 4173 31532 4219 31579
rect 4173 31498 4179 31532
rect 4213 31498 4219 31532
rect 4173 31460 4219 31498
rect 4173 31426 4179 31460
rect 4213 31426 4219 31460
rect 4173 31388 4219 31426
rect 4173 31354 4179 31388
rect 4213 31354 4219 31388
rect 4173 31307 4219 31354
rect 4269 31532 4315 31579
rect 4269 31498 4275 31532
rect 4309 31498 4315 31532
rect 4269 31460 4315 31498
rect 4269 31426 4275 31460
rect 4309 31426 4315 31460
rect 4269 31388 4315 31426
rect 4269 31354 4275 31388
rect 4309 31354 4315 31388
rect 4269 31307 4315 31354
rect 4365 31532 4411 31579
rect 4365 31498 4371 31532
rect 4405 31498 4411 31532
rect 4365 31460 4411 31498
rect 4365 31426 4371 31460
rect 4405 31426 4411 31460
rect 4365 31388 4411 31426
rect 4365 31354 4371 31388
rect 4405 31354 4411 31388
rect 4365 31307 4411 31354
rect 4461 31532 4507 31579
rect 4461 31498 4467 31532
rect 4501 31498 4507 31532
rect 4461 31460 4507 31498
rect 4461 31426 4467 31460
rect 4501 31426 4507 31460
rect 4461 31388 4507 31426
rect 4461 31354 4467 31388
rect 4501 31354 4507 31388
rect 4461 31307 4507 31354
rect 4557 31532 4603 31579
rect 4557 31498 4563 31532
rect 4597 31498 4603 31532
rect 4557 31460 4603 31498
rect 4557 31426 4563 31460
rect 4597 31426 4603 31460
rect 4557 31388 4603 31426
rect 4557 31354 4563 31388
rect 4597 31354 4603 31388
rect 4557 31307 4603 31354
rect 4653 31532 4699 31579
rect 4653 31498 4659 31532
rect 4693 31498 4699 31532
rect 4653 31460 4699 31498
rect 4653 31426 4659 31460
rect 4693 31426 4699 31460
rect 4653 31388 4699 31426
rect 4653 31354 4659 31388
rect 4693 31354 4699 31388
rect 4653 31307 4699 31354
rect 4749 31532 4795 31579
rect 4749 31498 4755 31532
rect 4789 31498 4795 31532
rect 4749 31460 4795 31498
rect 4749 31426 4755 31460
rect 4789 31426 4795 31460
rect 4749 31388 4795 31426
rect 4749 31354 4755 31388
rect 4789 31354 4795 31388
rect 4749 31307 4795 31354
rect 4845 31532 4891 31579
rect 4845 31498 4851 31532
rect 4885 31498 4891 31532
rect 4845 31460 4891 31498
rect 4845 31426 4851 31460
rect 4885 31426 4891 31460
rect 4845 31388 4891 31426
rect 4845 31354 4851 31388
rect 4885 31354 4891 31388
rect 4845 31307 4891 31354
rect 4941 31532 4987 31579
rect 4941 31498 4947 31532
rect 4981 31498 4987 31532
rect 4941 31460 4987 31498
rect 4941 31426 4947 31460
rect 4981 31426 4987 31460
rect 4941 31388 4987 31426
rect 4941 31354 4947 31388
rect 4981 31354 4987 31388
rect 4941 31307 4987 31354
rect 5055 31563 5101 31601
rect 5055 31529 5061 31563
rect 5095 31529 5101 31563
rect 5055 31491 5101 31529
rect 5055 31457 5061 31491
rect 5095 31460 5101 31491
rect 5274 31460 5550 31461
rect 5095 31457 5550 31460
rect 5055 31430 5550 31457
rect 5055 31419 5303 31430
rect 5055 31385 5061 31419
rect 5095 31396 5303 31419
rect 5337 31396 5395 31430
rect 5429 31396 5487 31430
rect 5521 31396 5550 31430
rect 5095 31385 5550 31396
rect 5055 31365 5550 31385
rect 5055 31347 5101 31365
rect 5055 31313 5061 31347
rect 5095 31313 5101 31347
rect 2466 31132 3837 31166
rect 2466 30999 2500 31132
rect 2658 30999 2692 31132
rect 2850 30999 2884 31132
rect 3042 30999 3076 31132
rect 3234 30999 3268 31132
rect 3426 30999 3460 31132
rect 3671 31042 3681 31094
rect 3733 31042 3743 31094
rect 3679 31041 3691 31042
rect 3725 31041 3737 31042
rect 3679 31035 3737 31041
rect 3534 31006 3580 31029
rect 2460 30964 2506 30999
rect 2460 30930 2466 30964
rect 2500 30930 2506 30964
rect 2460 30895 2506 30930
rect 2556 30964 2602 30999
rect 2556 30930 2562 30964
rect 2596 30930 2602 30964
rect 2556 30895 2602 30930
rect 2652 30964 2698 30999
rect 2652 30930 2658 30964
rect 2692 30930 2698 30964
rect 2652 30895 2698 30930
rect 2748 30964 2794 30999
rect 2748 30930 2754 30964
rect 2788 30930 2794 30964
rect 2748 30895 2794 30930
rect 2844 30964 2890 30999
rect 2844 30930 2850 30964
rect 2884 30930 2890 30964
rect 2844 30895 2890 30930
rect 2940 30964 2986 30999
rect 2940 30930 2946 30964
rect 2980 30930 2986 30964
rect 2940 30895 2986 30930
rect 3036 30964 3082 30999
rect 3036 30930 3042 30964
rect 3076 30930 3082 30964
rect 3036 30895 3082 30930
rect 3132 30964 3178 30999
rect 3132 30930 3138 30964
rect 3172 30930 3178 30964
rect 3132 30895 3178 30930
rect 3228 30964 3274 30999
rect 3228 30930 3234 30964
rect 3268 30930 3274 30964
rect 3228 30895 3274 30930
rect 3324 30964 3370 30999
rect 3324 30930 3330 30964
rect 3364 30930 3370 30964
rect 3324 30895 3370 30930
rect 3420 30964 3466 30999
rect 3420 30930 3426 30964
rect 3460 30930 3466 30964
rect 3420 30895 3466 30930
rect 3534 30972 3540 31006
rect 3574 31004 3580 31006
rect 3803 31004 3837 31132
rect 3574 31003 3680 31004
rect 3734 31003 3837 31004
rect 3574 30991 3687 31003
rect 3574 30972 3647 30991
rect 3534 30934 3647 30972
rect 3534 30900 3540 30934
rect 3574 30915 3647 30934
rect 3681 30915 3687 30991
rect 3574 30904 3687 30915
rect 3574 30900 3580 30904
rect 3641 30903 3687 30904
rect 3729 30991 3837 31003
rect 3987 31166 4021 31307
rect 4179 31166 4213 31307
rect 4371 31166 4405 31307
rect 4563 31166 4597 31307
rect 4755 31166 4789 31307
rect 4947 31166 4981 31307
rect 5055 31269 5101 31313
rect 5683 31220 5743 32473
rect 5177 31186 5743 31220
rect 5177 31166 5211 31186
rect 3987 31132 5211 31166
rect 3987 30999 4021 31132
rect 4179 30999 4213 31132
rect 4371 30999 4405 31132
rect 4563 30999 4597 31132
rect 4755 30999 4789 31132
rect 4947 30999 4981 31132
rect 5438 31128 5512 31129
rect 5326 31126 5400 31127
rect 5326 31074 5337 31126
rect 5389 31074 5400 31126
rect 5438 31076 5449 31128
rect 5501 31076 5512 31128
rect 5438 31075 5512 31076
rect 5326 31073 5400 31074
rect 5055 31006 5101 31029
rect 3729 30915 3735 30991
rect 3769 30915 3837 30991
rect 3729 30904 3837 30915
rect 3729 30903 3775 30904
rect 2450 30864 2516 30867
rect 2447 30812 2457 30864
rect 2509 30812 2519 30864
rect 2450 30807 2516 30812
rect 2562 30755 2596 30895
rect 2642 30864 2708 30867
rect 2638 30812 2648 30864
rect 2700 30812 2710 30864
rect 2642 30807 2708 30812
rect 2754 30755 2788 30895
rect 2834 30864 2900 30867
rect 2830 30812 2840 30864
rect 2892 30812 2902 30864
rect 2834 30807 2900 30812
rect 2946 30755 2980 30895
rect 3026 30864 3092 30867
rect 3022 30812 3032 30864
rect 3084 30812 3094 30864
rect 3026 30807 3092 30812
rect 3138 30755 3172 30895
rect 3218 30863 3284 30867
rect 3215 30811 3225 30863
rect 3277 30811 3287 30863
rect 3218 30807 3284 30811
rect 3330 30755 3364 30895
rect 3410 30863 3476 30867
rect 3407 30811 3417 30863
rect 3469 30811 3479 30863
rect 3534 30862 3580 30900
rect 3534 30828 3540 30862
rect 3574 30828 3580 30862
rect 3410 30807 3476 30811
rect 2282 30721 3364 30755
rect 3534 30645 3580 30828
rect 3803 30755 3837 30904
rect 3981 30964 4027 30999
rect 3981 30930 3987 30964
rect 4021 30930 4027 30964
rect 3981 30895 4027 30930
rect 4077 30964 4123 30999
rect 4077 30930 4083 30964
rect 4117 30930 4123 30964
rect 4077 30895 4123 30930
rect 4173 30964 4219 30999
rect 4173 30930 4179 30964
rect 4213 30930 4219 30964
rect 4173 30895 4219 30930
rect 4269 30964 4315 30999
rect 4269 30930 4275 30964
rect 4309 30930 4315 30964
rect 4269 30895 4315 30930
rect 4365 30964 4411 30999
rect 4365 30930 4371 30964
rect 4405 30930 4411 30964
rect 4365 30895 4411 30930
rect 4461 30964 4507 30999
rect 4461 30930 4467 30964
rect 4501 30930 4507 30964
rect 4461 30895 4507 30930
rect 4557 30964 4603 30999
rect 4557 30930 4563 30964
rect 4597 30930 4603 30964
rect 4557 30895 4603 30930
rect 4653 30964 4699 30999
rect 4653 30930 4659 30964
rect 4693 30930 4699 30964
rect 4653 30895 4699 30930
rect 4749 30964 4795 30999
rect 4749 30930 4755 30964
rect 4789 30930 4795 30964
rect 4749 30895 4795 30930
rect 4845 30964 4891 30999
rect 4845 30930 4851 30964
rect 4885 30930 4891 30964
rect 4845 30895 4891 30930
rect 4941 30964 4987 30999
rect 4941 30930 4947 30964
rect 4981 30930 4987 30964
rect 4941 30895 4987 30930
rect 5055 30972 5061 31006
rect 5095 30972 5101 31006
rect 5055 30934 5101 30972
rect 5055 30900 5061 30934
rect 5095 30917 5101 30934
rect 5095 30900 5550 30917
rect 3971 30864 4037 30867
rect 3968 30812 3978 30864
rect 4030 30812 4040 30864
rect 3971 30807 4037 30812
rect 4083 30755 4117 30895
rect 4163 30864 4229 30867
rect 4159 30812 4169 30864
rect 4221 30812 4231 30864
rect 4163 30807 4229 30812
rect 4275 30755 4309 30895
rect 4355 30864 4421 30867
rect 4351 30812 4361 30864
rect 4413 30812 4423 30864
rect 4355 30807 4421 30812
rect 4467 30755 4501 30895
rect 4547 30864 4613 30867
rect 4543 30812 4553 30864
rect 4605 30812 4615 30864
rect 4547 30807 4613 30812
rect 4659 30755 4693 30895
rect 4739 30863 4805 30867
rect 4736 30811 4746 30863
rect 4798 30811 4808 30863
rect 4739 30807 4805 30811
rect 4851 30755 4885 30895
rect 5055 30886 5550 30900
rect 4931 30863 4997 30867
rect 4928 30811 4938 30863
rect 4990 30811 5000 30863
rect 5055 30862 5303 30886
rect 5055 30828 5061 30862
rect 5095 30852 5303 30862
rect 5337 30852 5395 30886
rect 5429 30852 5487 30886
rect 5521 30852 5550 30886
rect 5095 30828 5550 30852
rect 5055 30821 5550 30828
rect 4931 30807 4997 30811
rect 3803 30721 4885 30755
rect 5055 30646 5101 30821
rect 129 30438 1211 30472
rect 129 29875 163 30438
rect 294 30328 304 30380
rect 356 30328 366 30380
rect 409 30288 443 30438
rect 487 30328 497 30380
rect 549 30328 559 30380
rect 601 30288 635 30438
rect 678 30328 688 30380
rect 740 30328 750 30380
rect 793 30288 827 30438
rect 870 30328 880 30380
rect 932 30328 942 30380
rect 985 30288 1019 30438
rect 1062 30328 1072 30380
rect 1124 30328 1134 30380
rect 1177 30288 1211 30438
rect 1254 30328 1264 30380
rect 1316 30328 1326 30380
rect 1381 30344 1427 30508
rect 2282 30442 3364 30476
rect 1381 30310 1387 30344
rect 1421 30310 1427 30344
rect 1512 30321 1522 30381
rect 1578 30321 1792 30381
rect 1852 30321 1862 30381
rect 307 30241 353 30288
rect 307 30207 313 30241
rect 347 30207 353 30241
rect 307 30169 353 30207
rect 307 30135 313 30169
rect 347 30135 353 30169
rect 307 30097 353 30135
rect 307 30063 313 30097
rect 347 30063 353 30097
rect 307 30016 353 30063
rect 403 30241 449 30288
rect 403 30207 409 30241
rect 443 30207 449 30241
rect 403 30169 449 30207
rect 403 30135 409 30169
rect 443 30135 449 30169
rect 403 30097 449 30135
rect 403 30063 409 30097
rect 443 30063 449 30097
rect 403 30016 449 30063
rect 499 30241 545 30288
rect 499 30207 505 30241
rect 539 30207 545 30241
rect 499 30169 545 30207
rect 499 30135 505 30169
rect 539 30135 545 30169
rect 499 30097 545 30135
rect 499 30063 505 30097
rect 539 30063 545 30097
rect 499 30016 545 30063
rect 595 30241 641 30288
rect 595 30207 601 30241
rect 635 30207 641 30241
rect 595 30169 641 30207
rect 595 30135 601 30169
rect 635 30135 641 30169
rect 595 30097 641 30135
rect 595 30063 601 30097
rect 635 30063 641 30097
rect 595 30016 641 30063
rect 691 30241 737 30288
rect 691 30207 697 30241
rect 731 30207 737 30241
rect 691 30169 737 30207
rect 691 30135 697 30169
rect 731 30135 737 30169
rect 691 30097 737 30135
rect 691 30063 697 30097
rect 731 30063 737 30097
rect 691 30016 737 30063
rect 787 30241 833 30288
rect 787 30207 793 30241
rect 827 30207 833 30241
rect 787 30169 833 30207
rect 787 30135 793 30169
rect 827 30135 833 30169
rect 787 30097 833 30135
rect 787 30063 793 30097
rect 827 30063 833 30097
rect 787 30016 833 30063
rect 883 30241 929 30288
rect 883 30207 889 30241
rect 923 30207 929 30241
rect 883 30169 929 30207
rect 883 30135 889 30169
rect 923 30135 929 30169
rect 883 30097 929 30135
rect 883 30063 889 30097
rect 923 30063 929 30097
rect 883 30016 929 30063
rect 979 30241 1025 30288
rect 979 30207 985 30241
rect 1019 30207 1025 30241
rect 979 30169 1025 30207
rect 979 30135 985 30169
rect 1019 30135 1025 30169
rect 979 30097 1025 30135
rect 979 30063 985 30097
rect 1019 30063 1025 30097
rect 979 30016 1025 30063
rect 1075 30241 1121 30288
rect 1075 30207 1081 30241
rect 1115 30207 1121 30241
rect 1075 30169 1121 30207
rect 1075 30135 1081 30169
rect 1115 30135 1121 30169
rect 1075 30097 1121 30135
rect 1075 30063 1081 30097
rect 1115 30063 1121 30097
rect 1075 30016 1121 30063
rect 1171 30241 1217 30288
rect 1171 30207 1177 30241
rect 1211 30207 1217 30241
rect 1171 30169 1217 30207
rect 1171 30135 1177 30169
rect 1211 30135 1217 30169
rect 1171 30097 1217 30135
rect 1171 30063 1177 30097
rect 1211 30063 1217 30097
rect 1171 30016 1217 30063
rect 1267 30241 1313 30288
rect 1267 30207 1273 30241
rect 1307 30207 1313 30241
rect 1267 30169 1313 30207
rect 1267 30135 1273 30169
rect 1307 30135 1313 30169
rect 1267 30097 1313 30135
rect 1267 30063 1273 30097
rect 1307 30063 1313 30097
rect 1267 30016 1313 30063
rect 1381 30272 1427 30310
rect 1381 30238 1387 30272
rect 1421 30238 1427 30272
rect 1381 30200 1427 30238
rect 1381 30166 1387 30200
rect 1421 30166 1427 30200
rect 1381 30128 1427 30166
rect 1381 30094 1387 30128
rect 1421 30094 1427 30128
rect 1381 30084 1427 30094
rect 1381 30082 2160 30084
rect 1381 30056 2056 30082
rect 1381 30031 1387 30056
rect 1380 30022 1387 30031
rect 1421 30022 2056 30056
rect 0 29841 163 29875
rect 129 29464 163 29841
rect 313 29875 347 30016
rect 505 29875 539 30016
rect 697 29875 731 30016
rect 889 29875 923 30016
rect 1081 29875 1115 30016
rect 1273 29875 1307 30016
rect 1380 29974 2056 30022
rect 2190 29974 2200 30082
rect 1380 29972 2160 29974
rect 2282 29879 2316 30442
rect 2447 30332 2457 30384
rect 2509 30332 2519 30384
rect 2562 30292 2596 30442
rect 2640 30332 2650 30384
rect 2702 30332 2712 30384
rect 2754 30292 2788 30442
rect 2831 30332 2841 30384
rect 2893 30332 2903 30384
rect 2946 30292 2980 30442
rect 3023 30332 3033 30384
rect 3085 30332 3095 30384
rect 3138 30292 3172 30442
rect 3215 30332 3225 30384
rect 3277 30332 3287 30384
rect 3330 30292 3364 30442
rect 3407 30332 3417 30384
rect 3469 30332 3479 30384
rect 3534 30348 3580 30556
rect 3534 30314 3540 30348
rect 3574 30314 3580 30348
rect 2460 30245 2506 30292
rect 2460 30211 2466 30245
rect 2500 30211 2506 30245
rect 2460 30173 2506 30211
rect 2460 30139 2466 30173
rect 2500 30139 2506 30173
rect 2460 30101 2506 30139
rect 2460 30067 2466 30101
rect 2500 30067 2506 30101
rect 2460 30020 2506 30067
rect 2556 30245 2602 30292
rect 2556 30211 2562 30245
rect 2596 30211 2602 30245
rect 2556 30173 2602 30211
rect 2556 30139 2562 30173
rect 2596 30139 2602 30173
rect 2556 30101 2602 30139
rect 2556 30067 2562 30101
rect 2596 30067 2602 30101
rect 2556 30020 2602 30067
rect 2652 30245 2698 30292
rect 2652 30211 2658 30245
rect 2692 30211 2698 30245
rect 2652 30173 2698 30211
rect 2652 30139 2658 30173
rect 2692 30139 2698 30173
rect 2652 30101 2698 30139
rect 2652 30067 2658 30101
rect 2692 30067 2698 30101
rect 2652 30020 2698 30067
rect 2748 30245 2794 30292
rect 2748 30211 2754 30245
rect 2788 30211 2794 30245
rect 2748 30173 2794 30211
rect 2748 30139 2754 30173
rect 2788 30139 2794 30173
rect 2748 30101 2794 30139
rect 2748 30067 2754 30101
rect 2788 30067 2794 30101
rect 2748 30020 2794 30067
rect 2844 30245 2890 30292
rect 2844 30211 2850 30245
rect 2884 30211 2890 30245
rect 2844 30173 2890 30211
rect 2844 30139 2850 30173
rect 2884 30139 2890 30173
rect 2844 30101 2890 30139
rect 2844 30067 2850 30101
rect 2884 30067 2890 30101
rect 2844 30020 2890 30067
rect 2940 30245 2986 30292
rect 2940 30211 2946 30245
rect 2980 30211 2986 30245
rect 2940 30173 2986 30211
rect 2940 30139 2946 30173
rect 2980 30139 2986 30173
rect 2940 30101 2986 30139
rect 2940 30067 2946 30101
rect 2980 30067 2986 30101
rect 2940 30020 2986 30067
rect 3036 30245 3082 30292
rect 3036 30211 3042 30245
rect 3076 30211 3082 30245
rect 3036 30173 3082 30211
rect 3036 30139 3042 30173
rect 3076 30139 3082 30173
rect 3036 30101 3082 30139
rect 3036 30067 3042 30101
rect 3076 30067 3082 30101
rect 3036 30020 3082 30067
rect 3132 30245 3178 30292
rect 3132 30211 3138 30245
rect 3172 30211 3178 30245
rect 3132 30173 3178 30211
rect 3132 30139 3138 30173
rect 3172 30139 3178 30173
rect 3132 30101 3178 30139
rect 3132 30067 3138 30101
rect 3172 30067 3178 30101
rect 3132 30020 3178 30067
rect 3228 30245 3274 30292
rect 3228 30211 3234 30245
rect 3268 30211 3274 30245
rect 3228 30173 3274 30211
rect 3228 30139 3234 30173
rect 3268 30139 3274 30173
rect 3228 30101 3274 30139
rect 3228 30067 3234 30101
rect 3268 30067 3274 30101
rect 3228 30020 3274 30067
rect 3324 30245 3370 30292
rect 3324 30211 3330 30245
rect 3364 30211 3370 30245
rect 3324 30173 3370 30211
rect 3324 30139 3330 30173
rect 3364 30139 3370 30173
rect 3324 30101 3370 30139
rect 3324 30067 3330 30101
rect 3364 30067 3370 30101
rect 3324 30020 3370 30067
rect 3420 30245 3466 30292
rect 3420 30211 3426 30245
rect 3460 30211 3466 30245
rect 3420 30173 3466 30211
rect 3420 30139 3426 30173
rect 3460 30139 3466 30173
rect 3420 30101 3466 30139
rect 3420 30067 3426 30101
rect 3460 30067 3466 30101
rect 3420 30020 3466 30067
rect 3534 30276 3580 30314
rect 3534 30242 3540 30276
rect 3574 30242 3580 30276
rect 3534 30204 3580 30242
rect 3534 30170 3540 30204
rect 3574 30170 3580 30204
rect 3534 30132 3580 30170
rect 3534 30098 3540 30132
rect 3574 30098 3580 30132
rect 3534 30060 3580 30098
rect 3534 30026 3540 30060
rect 3574 30026 3580 30060
rect 2101 29875 2316 29879
rect 313 29845 2316 29875
rect 313 29841 2141 29845
rect 313 29708 347 29841
rect 505 29708 539 29841
rect 697 29708 731 29841
rect 889 29708 923 29841
rect 1081 29708 1115 29841
rect 1273 29708 1307 29841
rect 1381 29715 1608 29738
rect 307 29673 353 29708
rect 307 29639 313 29673
rect 347 29639 353 29673
rect 307 29604 353 29639
rect 403 29673 449 29708
rect 403 29639 409 29673
rect 443 29639 449 29673
rect 403 29604 449 29639
rect 499 29673 545 29708
rect 499 29639 505 29673
rect 539 29639 545 29673
rect 499 29604 545 29639
rect 595 29673 641 29708
rect 595 29639 601 29673
rect 635 29639 641 29673
rect 595 29604 641 29639
rect 691 29673 737 29708
rect 691 29639 697 29673
rect 731 29639 737 29673
rect 691 29604 737 29639
rect 787 29673 833 29708
rect 787 29639 793 29673
rect 827 29639 833 29673
rect 787 29604 833 29639
rect 883 29673 929 29708
rect 883 29639 889 29673
rect 923 29639 929 29673
rect 883 29604 929 29639
rect 979 29673 1025 29708
rect 979 29639 985 29673
rect 1019 29639 1025 29673
rect 979 29604 1025 29639
rect 1075 29673 1121 29708
rect 1075 29639 1081 29673
rect 1115 29639 1121 29673
rect 1075 29604 1121 29639
rect 1171 29673 1217 29708
rect 1171 29639 1177 29673
rect 1211 29639 1217 29673
rect 1171 29604 1217 29639
rect 1267 29673 1313 29708
rect 1267 29639 1273 29673
rect 1307 29639 1313 29673
rect 1267 29604 1313 29639
rect 1381 29681 1387 29715
rect 1421 29681 1608 29715
rect 1381 29643 1608 29681
rect 1381 29609 1387 29643
rect 1421 29618 1608 29643
rect 1421 29609 1427 29618
rect 1560 29616 1608 29618
rect 1598 29614 1608 29616
rect 1720 29614 1730 29738
rect 297 29573 363 29576
rect 294 29521 304 29573
rect 356 29521 366 29573
rect 297 29516 363 29521
rect 409 29464 443 29604
rect 489 29573 555 29576
rect 485 29521 495 29573
rect 547 29521 557 29573
rect 489 29516 555 29521
rect 601 29464 635 29604
rect 681 29573 747 29576
rect 677 29521 687 29573
rect 739 29521 749 29573
rect 681 29516 747 29521
rect 793 29464 827 29604
rect 873 29573 939 29576
rect 869 29521 879 29573
rect 931 29521 941 29573
rect 873 29516 939 29521
rect 985 29464 1019 29604
rect 1065 29572 1131 29576
rect 1062 29520 1072 29572
rect 1124 29520 1134 29572
rect 1065 29516 1131 29520
rect 1177 29464 1211 29604
rect 1257 29572 1323 29576
rect 1254 29520 1264 29572
rect 1316 29520 1326 29572
rect 1381 29571 1427 29609
rect 1920 29576 1930 29578
rect 1381 29537 1387 29571
rect 1421 29537 1427 29571
rect 1257 29516 1323 29520
rect 129 29430 1211 29464
rect 1381 29394 1427 29537
rect 1458 29520 1468 29576
rect 1524 29522 1930 29576
rect 1986 29522 1996 29578
rect 1524 29520 1986 29522
rect 2282 29468 2316 29845
rect 2466 29879 2500 30020
rect 2658 29879 2692 30020
rect 2850 29879 2884 30020
rect 3042 29879 3076 30020
rect 3234 29879 3268 30020
rect 3426 29879 3460 30020
rect 3534 29982 3580 30026
rect 3803 30442 4885 30476
rect 3803 29879 3837 30442
rect 3968 30332 3978 30384
rect 4030 30332 4040 30384
rect 4083 30292 4117 30442
rect 4161 30332 4171 30384
rect 4223 30332 4233 30384
rect 4275 30292 4309 30442
rect 4352 30332 4362 30384
rect 4414 30332 4424 30384
rect 4467 30292 4501 30442
rect 4544 30332 4554 30384
rect 4606 30332 4616 30384
rect 4659 30292 4693 30442
rect 4736 30332 4746 30384
rect 4798 30332 4808 30384
rect 4851 30292 4885 30442
rect 4928 30332 4938 30384
rect 4990 30332 5000 30384
rect 5055 30348 5101 30553
rect 5055 30314 5061 30348
rect 5095 30314 5101 30348
rect 3981 30245 4027 30292
rect 3981 30211 3987 30245
rect 4021 30211 4027 30245
rect 3981 30173 4027 30211
rect 3981 30139 3987 30173
rect 4021 30139 4027 30173
rect 3981 30101 4027 30139
rect 3981 30067 3987 30101
rect 4021 30067 4027 30101
rect 3981 30020 4027 30067
rect 4077 30245 4123 30292
rect 4077 30211 4083 30245
rect 4117 30211 4123 30245
rect 4077 30173 4123 30211
rect 4077 30139 4083 30173
rect 4117 30139 4123 30173
rect 4077 30101 4123 30139
rect 4077 30067 4083 30101
rect 4117 30067 4123 30101
rect 4077 30020 4123 30067
rect 4173 30245 4219 30292
rect 4173 30211 4179 30245
rect 4213 30211 4219 30245
rect 4173 30173 4219 30211
rect 4173 30139 4179 30173
rect 4213 30139 4219 30173
rect 4173 30101 4219 30139
rect 4173 30067 4179 30101
rect 4213 30067 4219 30101
rect 4173 30020 4219 30067
rect 4269 30245 4315 30292
rect 4269 30211 4275 30245
rect 4309 30211 4315 30245
rect 4269 30173 4315 30211
rect 4269 30139 4275 30173
rect 4309 30139 4315 30173
rect 4269 30101 4315 30139
rect 4269 30067 4275 30101
rect 4309 30067 4315 30101
rect 4269 30020 4315 30067
rect 4365 30245 4411 30292
rect 4365 30211 4371 30245
rect 4405 30211 4411 30245
rect 4365 30173 4411 30211
rect 4365 30139 4371 30173
rect 4405 30139 4411 30173
rect 4365 30101 4411 30139
rect 4365 30067 4371 30101
rect 4405 30067 4411 30101
rect 4365 30020 4411 30067
rect 4461 30245 4507 30292
rect 4461 30211 4467 30245
rect 4501 30211 4507 30245
rect 4461 30173 4507 30211
rect 4461 30139 4467 30173
rect 4501 30139 4507 30173
rect 4461 30101 4507 30139
rect 4461 30067 4467 30101
rect 4501 30067 4507 30101
rect 4461 30020 4507 30067
rect 4557 30245 4603 30292
rect 4557 30211 4563 30245
rect 4597 30211 4603 30245
rect 4557 30173 4603 30211
rect 4557 30139 4563 30173
rect 4597 30139 4603 30173
rect 4557 30101 4603 30139
rect 4557 30067 4563 30101
rect 4597 30067 4603 30101
rect 4557 30020 4603 30067
rect 4653 30245 4699 30292
rect 4653 30211 4659 30245
rect 4693 30211 4699 30245
rect 4653 30173 4699 30211
rect 4653 30139 4659 30173
rect 4693 30139 4699 30173
rect 4653 30101 4699 30139
rect 4653 30067 4659 30101
rect 4693 30067 4699 30101
rect 4653 30020 4699 30067
rect 4749 30245 4795 30292
rect 4749 30211 4755 30245
rect 4789 30211 4795 30245
rect 4749 30173 4795 30211
rect 4749 30139 4755 30173
rect 4789 30139 4795 30173
rect 4749 30101 4795 30139
rect 4749 30067 4755 30101
rect 4789 30067 4795 30101
rect 4749 30020 4795 30067
rect 4845 30245 4891 30292
rect 4845 30211 4851 30245
rect 4885 30211 4891 30245
rect 4845 30173 4891 30211
rect 4845 30139 4851 30173
rect 4885 30139 4891 30173
rect 4845 30101 4891 30139
rect 4845 30067 4851 30101
rect 4885 30067 4891 30101
rect 4845 30020 4891 30067
rect 4941 30245 4987 30292
rect 4941 30211 4947 30245
rect 4981 30211 4987 30245
rect 4941 30173 4987 30211
rect 4941 30139 4947 30173
rect 4981 30139 4987 30173
rect 4941 30101 4987 30139
rect 4941 30067 4947 30101
rect 4981 30067 4987 30101
rect 4941 30020 4987 30067
rect 5055 30276 5101 30314
rect 5055 30242 5061 30276
rect 5095 30242 5101 30276
rect 5055 30204 5101 30242
rect 5055 30170 5061 30204
rect 5095 30173 5101 30204
rect 5274 30173 5550 30174
rect 5095 30170 5550 30173
rect 5055 30143 5550 30170
rect 5055 30132 5303 30143
rect 5055 30098 5061 30132
rect 5095 30109 5303 30132
rect 5337 30109 5395 30143
rect 5429 30109 5487 30143
rect 5521 30109 5550 30143
rect 5095 30098 5550 30109
rect 5055 30078 5550 30098
rect 5055 30060 5101 30078
rect 5055 30026 5061 30060
rect 5095 30026 5101 30060
rect 2466 29845 3837 29879
rect 2466 29712 2500 29845
rect 2658 29712 2692 29845
rect 2850 29712 2884 29845
rect 3042 29712 3076 29845
rect 3234 29712 3268 29845
rect 3426 29712 3460 29845
rect 3671 29755 3681 29807
rect 3733 29755 3743 29807
rect 3679 29754 3691 29755
rect 3725 29754 3737 29755
rect 3679 29748 3737 29754
rect 3534 29719 3580 29742
rect 2460 29677 2506 29712
rect 2460 29643 2466 29677
rect 2500 29643 2506 29677
rect 2460 29608 2506 29643
rect 2556 29677 2602 29712
rect 2556 29643 2562 29677
rect 2596 29643 2602 29677
rect 2556 29608 2602 29643
rect 2652 29677 2698 29712
rect 2652 29643 2658 29677
rect 2692 29643 2698 29677
rect 2652 29608 2698 29643
rect 2748 29677 2794 29712
rect 2748 29643 2754 29677
rect 2788 29643 2794 29677
rect 2748 29608 2794 29643
rect 2844 29677 2890 29712
rect 2844 29643 2850 29677
rect 2884 29643 2890 29677
rect 2844 29608 2890 29643
rect 2940 29677 2986 29712
rect 2940 29643 2946 29677
rect 2980 29643 2986 29677
rect 2940 29608 2986 29643
rect 3036 29677 3082 29712
rect 3036 29643 3042 29677
rect 3076 29643 3082 29677
rect 3036 29608 3082 29643
rect 3132 29677 3178 29712
rect 3132 29643 3138 29677
rect 3172 29643 3178 29677
rect 3132 29608 3178 29643
rect 3228 29677 3274 29712
rect 3228 29643 3234 29677
rect 3268 29643 3274 29677
rect 3228 29608 3274 29643
rect 3324 29677 3370 29712
rect 3324 29643 3330 29677
rect 3364 29643 3370 29677
rect 3324 29608 3370 29643
rect 3420 29677 3466 29712
rect 3420 29643 3426 29677
rect 3460 29643 3466 29677
rect 3420 29608 3466 29643
rect 3534 29685 3540 29719
rect 3574 29717 3580 29719
rect 3803 29717 3837 29845
rect 3574 29716 3680 29717
rect 3734 29716 3837 29717
rect 3574 29704 3687 29716
rect 3574 29685 3647 29704
rect 3534 29647 3647 29685
rect 3534 29613 3540 29647
rect 3574 29628 3647 29647
rect 3681 29628 3687 29704
rect 3574 29617 3687 29628
rect 3574 29613 3580 29617
rect 3641 29616 3687 29617
rect 3729 29704 3837 29716
rect 3987 29879 4021 30020
rect 4179 29879 4213 30020
rect 4371 29879 4405 30020
rect 4563 29879 4597 30020
rect 4755 29879 4789 30020
rect 4947 29879 4981 30020
rect 5055 29982 5101 30026
rect 5683 29933 5743 31186
rect 5177 29899 5743 29933
rect 5177 29879 5211 29899
rect 3987 29845 5211 29879
rect 3987 29712 4021 29845
rect 4179 29712 4213 29845
rect 4371 29712 4405 29845
rect 4563 29712 4597 29845
rect 4755 29712 4789 29845
rect 4947 29712 4981 29845
rect 5438 29841 5512 29842
rect 5326 29839 5400 29840
rect 5326 29787 5337 29839
rect 5389 29787 5400 29839
rect 5438 29789 5449 29841
rect 5501 29789 5512 29841
rect 5438 29788 5512 29789
rect 5326 29786 5400 29787
rect 5055 29719 5101 29742
rect 3729 29628 3735 29704
rect 3769 29628 3837 29704
rect 3729 29617 3837 29628
rect 3729 29616 3775 29617
rect 2450 29577 2516 29580
rect 2447 29525 2457 29577
rect 2509 29525 2519 29577
rect 2450 29520 2516 29525
rect 2562 29468 2596 29608
rect 2642 29577 2708 29580
rect 2638 29525 2648 29577
rect 2700 29525 2710 29577
rect 2642 29520 2708 29525
rect 2754 29468 2788 29608
rect 2834 29577 2900 29580
rect 2830 29525 2840 29577
rect 2892 29525 2902 29577
rect 2834 29520 2900 29525
rect 2946 29468 2980 29608
rect 3026 29577 3092 29580
rect 3022 29525 3032 29577
rect 3084 29525 3094 29577
rect 3026 29520 3092 29525
rect 3138 29468 3172 29608
rect 3218 29576 3284 29580
rect 3215 29524 3225 29576
rect 3277 29524 3287 29576
rect 3218 29520 3284 29524
rect 3330 29468 3364 29608
rect 3410 29576 3476 29580
rect 3407 29524 3417 29576
rect 3469 29524 3479 29576
rect 3534 29575 3580 29613
rect 3534 29541 3540 29575
rect 3574 29541 3580 29575
rect 3410 29520 3476 29524
rect 2282 29434 3364 29468
rect 3534 29358 3580 29541
rect 3803 29468 3837 29617
rect 3981 29677 4027 29712
rect 3981 29643 3987 29677
rect 4021 29643 4027 29677
rect 3981 29608 4027 29643
rect 4077 29677 4123 29712
rect 4077 29643 4083 29677
rect 4117 29643 4123 29677
rect 4077 29608 4123 29643
rect 4173 29677 4219 29712
rect 4173 29643 4179 29677
rect 4213 29643 4219 29677
rect 4173 29608 4219 29643
rect 4269 29677 4315 29712
rect 4269 29643 4275 29677
rect 4309 29643 4315 29677
rect 4269 29608 4315 29643
rect 4365 29677 4411 29712
rect 4365 29643 4371 29677
rect 4405 29643 4411 29677
rect 4365 29608 4411 29643
rect 4461 29677 4507 29712
rect 4461 29643 4467 29677
rect 4501 29643 4507 29677
rect 4461 29608 4507 29643
rect 4557 29677 4603 29712
rect 4557 29643 4563 29677
rect 4597 29643 4603 29677
rect 4557 29608 4603 29643
rect 4653 29677 4699 29712
rect 4653 29643 4659 29677
rect 4693 29643 4699 29677
rect 4653 29608 4699 29643
rect 4749 29677 4795 29712
rect 4749 29643 4755 29677
rect 4789 29643 4795 29677
rect 4749 29608 4795 29643
rect 4845 29677 4891 29712
rect 4845 29643 4851 29677
rect 4885 29643 4891 29677
rect 4845 29608 4891 29643
rect 4941 29677 4987 29712
rect 4941 29643 4947 29677
rect 4981 29643 4987 29677
rect 4941 29608 4987 29643
rect 5055 29685 5061 29719
rect 5095 29685 5101 29719
rect 5055 29647 5101 29685
rect 5055 29613 5061 29647
rect 5095 29630 5101 29647
rect 5095 29613 5550 29630
rect 3971 29577 4037 29580
rect 3968 29525 3978 29577
rect 4030 29525 4040 29577
rect 3971 29520 4037 29525
rect 4083 29468 4117 29608
rect 4163 29577 4229 29580
rect 4159 29525 4169 29577
rect 4221 29525 4231 29577
rect 4163 29520 4229 29525
rect 4275 29468 4309 29608
rect 4355 29577 4421 29580
rect 4351 29525 4361 29577
rect 4413 29525 4423 29577
rect 4355 29520 4421 29525
rect 4467 29468 4501 29608
rect 4547 29577 4613 29580
rect 4543 29525 4553 29577
rect 4605 29525 4615 29577
rect 4547 29520 4613 29525
rect 4659 29468 4693 29608
rect 4739 29576 4805 29580
rect 4736 29524 4746 29576
rect 4798 29524 4808 29576
rect 4739 29520 4805 29524
rect 4851 29468 4885 29608
rect 5055 29599 5550 29613
rect 4931 29576 4997 29580
rect 4928 29524 4938 29576
rect 4990 29524 5000 29576
rect 5055 29575 5303 29599
rect 5055 29541 5061 29575
rect 5095 29565 5303 29575
rect 5337 29565 5395 29599
rect 5429 29565 5487 29599
rect 5521 29565 5550 29599
rect 5095 29541 5550 29565
rect 5055 29534 5550 29541
rect 4931 29520 4997 29524
rect 3803 29434 4885 29468
rect 5055 29359 5101 29534
rect 129 29151 1211 29185
rect 129 28588 163 29151
rect 294 29041 304 29093
rect 356 29041 366 29093
rect 409 29001 443 29151
rect 487 29041 497 29093
rect 549 29041 559 29093
rect 601 29001 635 29151
rect 678 29041 688 29093
rect 740 29041 750 29093
rect 793 29001 827 29151
rect 870 29041 880 29093
rect 932 29041 942 29093
rect 985 29001 1019 29151
rect 1062 29041 1072 29093
rect 1124 29041 1134 29093
rect 1177 29001 1211 29151
rect 1254 29041 1264 29093
rect 1316 29041 1326 29093
rect 1381 29057 1427 29221
rect 2282 29155 3364 29189
rect 1381 29023 1387 29057
rect 1421 29023 1427 29057
rect 1512 29034 1522 29094
rect 1578 29034 1792 29094
rect 1852 29034 1862 29094
rect 307 28954 353 29001
rect 307 28920 313 28954
rect 347 28920 353 28954
rect 307 28882 353 28920
rect 307 28848 313 28882
rect 347 28848 353 28882
rect 307 28810 353 28848
rect 307 28776 313 28810
rect 347 28776 353 28810
rect 307 28729 353 28776
rect 403 28954 449 29001
rect 403 28920 409 28954
rect 443 28920 449 28954
rect 403 28882 449 28920
rect 403 28848 409 28882
rect 443 28848 449 28882
rect 403 28810 449 28848
rect 403 28776 409 28810
rect 443 28776 449 28810
rect 403 28729 449 28776
rect 499 28954 545 29001
rect 499 28920 505 28954
rect 539 28920 545 28954
rect 499 28882 545 28920
rect 499 28848 505 28882
rect 539 28848 545 28882
rect 499 28810 545 28848
rect 499 28776 505 28810
rect 539 28776 545 28810
rect 499 28729 545 28776
rect 595 28954 641 29001
rect 595 28920 601 28954
rect 635 28920 641 28954
rect 595 28882 641 28920
rect 595 28848 601 28882
rect 635 28848 641 28882
rect 595 28810 641 28848
rect 595 28776 601 28810
rect 635 28776 641 28810
rect 595 28729 641 28776
rect 691 28954 737 29001
rect 691 28920 697 28954
rect 731 28920 737 28954
rect 691 28882 737 28920
rect 691 28848 697 28882
rect 731 28848 737 28882
rect 691 28810 737 28848
rect 691 28776 697 28810
rect 731 28776 737 28810
rect 691 28729 737 28776
rect 787 28954 833 29001
rect 787 28920 793 28954
rect 827 28920 833 28954
rect 787 28882 833 28920
rect 787 28848 793 28882
rect 827 28848 833 28882
rect 787 28810 833 28848
rect 787 28776 793 28810
rect 827 28776 833 28810
rect 787 28729 833 28776
rect 883 28954 929 29001
rect 883 28920 889 28954
rect 923 28920 929 28954
rect 883 28882 929 28920
rect 883 28848 889 28882
rect 923 28848 929 28882
rect 883 28810 929 28848
rect 883 28776 889 28810
rect 923 28776 929 28810
rect 883 28729 929 28776
rect 979 28954 1025 29001
rect 979 28920 985 28954
rect 1019 28920 1025 28954
rect 979 28882 1025 28920
rect 979 28848 985 28882
rect 1019 28848 1025 28882
rect 979 28810 1025 28848
rect 979 28776 985 28810
rect 1019 28776 1025 28810
rect 979 28729 1025 28776
rect 1075 28954 1121 29001
rect 1075 28920 1081 28954
rect 1115 28920 1121 28954
rect 1075 28882 1121 28920
rect 1075 28848 1081 28882
rect 1115 28848 1121 28882
rect 1075 28810 1121 28848
rect 1075 28776 1081 28810
rect 1115 28776 1121 28810
rect 1075 28729 1121 28776
rect 1171 28954 1217 29001
rect 1171 28920 1177 28954
rect 1211 28920 1217 28954
rect 1171 28882 1217 28920
rect 1171 28848 1177 28882
rect 1211 28848 1217 28882
rect 1171 28810 1217 28848
rect 1171 28776 1177 28810
rect 1211 28776 1217 28810
rect 1171 28729 1217 28776
rect 1267 28954 1313 29001
rect 1267 28920 1273 28954
rect 1307 28920 1313 28954
rect 1267 28882 1313 28920
rect 1267 28848 1273 28882
rect 1307 28848 1313 28882
rect 1267 28810 1313 28848
rect 1267 28776 1273 28810
rect 1307 28776 1313 28810
rect 1267 28729 1313 28776
rect 1381 28985 1427 29023
rect 1381 28951 1387 28985
rect 1421 28951 1427 28985
rect 1381 28913 1427 28951
rect 1381 28879 1387 28913
rect 1421 28879 1427 28913
rect 1381 28841 1427 28879
rect 1381 28807 1387 28841
rect 1421 28807 1427 28841
rect 1381 28797 1427 28807
rect 1381 28795 2160 28797
rect 1381 28769 2056 28795
rect 1381 28744 1387 28769
rect 1380 28735 1387 28744
rect 1421 28735 2056 28769
rect 0 28554 163 28588
rect 129 28177 163 28554
rect 313 28588 347 28729
rect 505 28588 539 28729
rect 697 28588 731 28729
rect 889 28588 923 28729
rect 1081 28588 1115 28729
rect 1273 28588 1307 28729
rect 1380 28687 2056 28735
rect 2190 28687 2200 28795
rect 1380 28685 2160 28687
rect 2282 28592 2316 29155
rect 2447 29045 2457 29097
rect 2509 29045 2519 29097
rect 2562 29005 2596 29155
rect 2640 29045 2650 29097
rect 2702 29045 2712 29097
rect 2754 29005 2788 29155
rect 2831 29045 2841 29097
rect 2893 29045 2903 29097
rect 2946 29005 2980 29155
rect 3023 29045 3033 29097
rect 3085 29045 3095 29097
rect 3138 29005 3172 29155
rect 3215 29045 3225 29097
rect 3277 29045 3287 29097
rect 3330 29005 3364 29155
rect 3407 29045 3417 29097
rect 3469 29045 3479 29097
rect 3534 29061 3580 29269
rect 3534 29027 3540 29061
rect 3574 29027 3580 29061
rect 2460 28958 2506 29005
rect 2460 28924 2466 28958
rect 2500 28924 2506 28958
rect 2460 28886 2506 28924
rect 2460 28852 2466 28886
rect 2500 28852 2506 28886
rect 2460 28814 2506 28852
rect 2460 28780 2466 28814
rect 2500 28780 2506 28814
rect 2460 28733 2506 28780
rect 2556 28958 2602 29005
rect 2556 28924 2562 28958
rect 2596 28924 2602 28958
rect 2556 28886 2602 28924
rect 2556 28852 2562 28886
rect 2596 28852 2602 28886
rect 2556 28814 2602 28852
rect 2556 28780 2562 28814
rect 2596 28780 2602 28814
rect 2556 28733 2602 28780
rect 2652 28958 2698 29005
rect 2652 28924 2658 28958
rect 2692 28924 2698 28958
rect 2652 28886 2698 28924
rect 2652 28852 2658 28886
rect 2692 28852 2698 28886
rect 2652 28814 2698 28852
rect 2652 28780 2658 28814
rect 2692 28780 2698 28814
rect 2652 28733 2698 28780
rect 2748 28958 2794 29005
rect 2748 28924 2754 28958
rect 2788 28924 2794 28958
rect 2748 28886 2794 28924
rect 2748 28852 2754 28886
rect 2788 28852 2794 28886
rect 2748 28814 2794 28852
rect 2748 28780 2754 28814
rect 2788 28780 2794 28814
rect 2748 28733 2794 28780
rect 2844 28958 2890 29005
rect 2844 28924 2850 28958
rect 2884 28924 2890 28958
rect 2844 28886 2890 28924
rect 2844 28852 2850 28886
rect 2884 28852 2890 28886
rect 2844 28814 2890 28852
rect 2844 28780 2850 28814
rect 2884 28780 2890 28814
rect 2844 28733 2890 28780
rect 2940 28958 2986 29005
rect 2940 28924 2946 28958
rect 2980 28924 2986 28958
rect 2940 28886 2986 28924
rect 2940 28852 2946 28886
rect 2980 28852 2986 28886
rect 2940 28814 2986 28852
rect 2940 28780 2946 28814
rect 2980 28780 2986 28814
rect 2940 28733 2986 28780
rect 3036 28958 3082 29005
rect 3036 28924 3042 28958
rect 3076 28924 3082 28958
rect 3036 28886 3082 28924
rect 3036 28852 3042 28886
rect 3076 28852 3082 28886
rect 3036 28814 3082 28852
rect 3036 28780 3042 28814
rect 3076 28780 3082 28814
rect 3036 28733 3082 28780
rect 3132 28958 3178 29005
rect 3132 28924 3138 28958
rect 3172 28924 3178 28958
rect 3132 28886 3178 28924
rect 3132 28852 3138 28886
rect 3172 28852 3178 28886
rect 3132 28814 3178 28852
rect 3132 28780 3138 28814
rect 3172 28780 3178 28814
rect 3132 28733 3178 28780
rect 3228 28958 3274 29005
rect 3228 28924 3234 28958
rect 3268 28924 3274 28958
rect 3228 28886 3274 28924
rect 3228 28852 3234 28886
rect 3268 28852 3274 28886
rect 3228 28814 3274 28852
rect 3228 28780 3234 28814
rect 3268 28780 3274 28814
rect 3228 28733 3274 28780
rect 3324 28958 3370 29005
rect 3324 28924 3330 28958
rect 3364 28924 3370 28958
rect 3324 28886 3370 28924
rect 3324 28852 3330 28886
rect 3364 28852 3370 28886
rect 3324 28814 3370 28852
rect 3324 28780 3330 28814
rect 3364 28780 3370 28814
rect 3324 28733 3370 28780
rect 3420 28958 3466 29005
rect 3420 28924 3426 28958
rect 3460 28924 3466 28958
rect 3420 28886 3466 28924
rect 3420 28852 3426 28886
rect 3460 28852 3466 28886
rect 3420 28814 3466 28852
rect 3420 28780 3426 28814
rect 3460 28780 3466 28814
rect 3420 28733 3466 28780
rect 3534 28989 3580 29027
rect 3534 28955 3540 28989
rect 3574 28955 3580 28989
rect 3534 28917 3580 28955
rect 3534 28883 3540 28917
rect 3574 28883 3580 28917
rect 3534 28845 3580 28883
rect 3534 28811 3540 28845
rect 3574 28811 3580 28845
rect 3534 28773 3580 28811
rect 3534 28739 3540 28773
rect 3574 28739 3580 28773
rect 2101 28588 2316 28592
rect 313 28558 2316 28588
rect 313 28554 2141 28558
rect 313 28421 347 28554
rect 505 28421 539 28554
rect 697 28421 731 28554
rect 889 28421 923 28554
rect 1081 28421 1115 28554
rect 1273 28421 1307 28554
rect 1381 28428 1608 28451
rect 307 28386 353 28421
rect 307 28352 313 28386
rect 347 28352 353 28386
rect 307 28317 353 28352
rect 403 28386 449 28421
rect 403 28352 409 28386
rect 443 28352 449 28386
rect 403 28317 449 28352
rect 499 28386 545 28421
rect 499 28352 505 28386
rect 539 28352 545 28386
rect 499 28317 545 28352
rect 595 28386 641 28421
rect 595 28352 601 28386
rect 635 28352 641 28386
rect 595 28317 641 28352
rect 691 28386 737 28421
rect 691 28352 697 28386
rect 731 28352 737 28386
rect 691 28317 737 28352
rect 787 28386 833 28421
rect 787 28352 793 28386
rect 827 28352 833 28386
rect 787 28317 833 28352
rect 883 28386 929 28421
rect 883 28352 889 28386
rect 923 28352 929 28386
rect 883 28317 929 28352
rect 979 28386 1025 28421
rect 979 28352 985 28386
rect 1019 28352 1025 28386
rect 979 28317 1025 28352
rect 1075 28386 1121 28421
rect 1075 28352 1081 28386
rect 1115 28352 1121 28386
rect 1075 28317 1121 28352
rect 1171 28386 1217 28421
rect 1171 28352 1177 28386
rect 1211 28352 1217 28386
rect 1171 28317 1217 28352
rect 1267 28386 1313 28421
rect 1267 28352 1273 28386
rect 1307 28352 1313 28386
rect 1267 28317 1313 28352
rect 1381 28394 1387 28428
rect 1421 28394 1608 28428
rect 1381 28356 1608 28394
rect 1381 28322 1387 28356
rect 1421 28331 1608 28356
rect 1421 28322 1427 28331
rect 1560 28329 1608 28331
rect 1598 28327 1608 28329
rect 1720 28327 1730 28451
rect 297 28286 363 28289
rect 294 28234 304 28286
rect 356 28234 366 28286
rect 297 28229 363 28234
rect 409 28177 443 28317
rect 489 28286 555 28289
rect 485 28234 495 28286
rect 547 28234 557 28286
rect 489 28229 555 28234
rect 601 28177 635 28317
rect 681 28286 747 28289
rect 677 28234 687 28286
rect 739 28234 749 28286
rect 681 28229 747 28234
rect 793 28177 827 28317
rect 873 28286 939 28289
rect 869 28234 879 28286
rect 931 28234 941 28286
rect 873 28229 939 28234
rect 985 28177 1019 28317
rect 1065 28285 1131 28289
rect 1062 28233 1072 28285
rect 1124 28233 1134 28285
rect 1065 28229 1131 28233
rect 1177 28177 1211 28317
rect 1257 28285 1323 28289
rect 1254 28233 1264 28285
rect 1316 28233 1326 28285
rect 1381 28284 1427 28322
rect 1920 28289 1930 28291
rect 1381 28250 1387 28284
rect 1421 28250 1427 28284
rect 1257 28229 1323 28233
rect 129 28143 1211 28177
rect 1381 28107 1427 28250
rect 1458 28233 1468 28289
rect 1524 28235 1930 28289
rect 1986 28235 1996 28291
rect 1524 28233 1986 28235
rect 2282 28181 2316 28558
rect 2466 28592 2500 28733
rect 2658 28592 2692 28733
rect 2850 28592 2884 28733
rect 3042 28592 3076 28733
rect 3234 28592 3268 28733
rect 3426 28592 3460 28733
rect 3534 28695 3580 28739
rect 3803 29155 4885 29189
rect 3803 28592 3837 29155
rect 3968 29045 3978 29097
rect 4030 29045 4040 29097
rect 4083 29005 4117 29155
rect 4161 29045 4171 29097
rect 4223 29045 4233 29097
rect 4275 29005 4309 29155
rect 4352 29045 4362 29097
rect 4414 29045 4424 29097
rect 4467 29005 4501 29155
rect 4544 29045 4554 29097
rect 4606 29045 4616 29097
rect 4659 29005 4693 29155
rect 4736 29045 4746 29097
rect 4798 29045 4808 29097
rect 4851 29005 4885 29155
rect 4928 29045 4938 29097
rect 4990 29045 5000 29097
rect 5055 29061 5101 29266
rect 5055 29027 5061 29061
rect 5095 29027 5101 29061
rect 3981 28958 4027 29005
rect 3981 28924 3987 28958
rect 4021 28924 4027 28958
rect 3981 28886 4027 28924
rect 3981 28852 3987 28886
rect 4021 28852 4027 28886
rect 3981 28814 4027 28852
rect 3981 28780 3987 28814
rect 4021 28780 4027 28814
rect 3981 28733 4027 28780
rect 4077 28958 4123 29005
rect 4077 28924 4083 28958
rect 4117 28924 4123 28958
rect 4077 28886 4123 28924
rect 4077 28852 4083 28886
rect 4117 28852 4123 28886
rect 4077 28814 4123 28852
rect 4077 28780 4083 28814
rect 4117 28780 4123 28814
rect 4077 28733 4123 28780
rect 4173 28958 4219 29005
rect 4173 28924 4179 28958
rect 4213 28924 4219 28958
rect 4173 28886 4219 28924
rect 4173 28852 4179 28886
rect 4213 28852 4219 28886
rect 4173 28814 4219 28852
rect 4173 28780 4179 28814
rect 4213 28780 4219 28814
rect 4173 28733 4219 28780
rect 4269 28958 4315 29005
rect 4269 28924 4275 28958
rect 4309 28924 4315 28958
rect 4269 28886 4315 28924
rect 4269 28852 4275 28886
rect 4309 28852 4315 28886
rect 4269 28814 4315 28852
rect 4269 28780 4275 28814
rect 4309 28780 4315 28814
rect 4269 28733 4315 28780
rect 4365 28958 4411 29005
rect 4365 28924 4371 28958
rect 4405 28924 4411 28958
rect 4365 28886 4411 28924
rect 4365 28852 4371 28886
rect 4405 28852 4411 28886
rect 4365 28814 4411 28852
rect 4365 28780 4371 28814
rect 4405 28780 4411 28814
rect 4365 28733 4411 28780
rect 4461 28958 4507 29005
rect 4461 28924 4467 28958
rect 4501 28924 4507 28958
rect 4461 28886 4507 28924
rect 4461 28852 4467 28886
rect 4501 28852 4507 28886
rect 4461 28814 4507 28852
rect 4461 28780 4467 28814
rect 4501 28780 4507 28814
rect 4461 28733 4507 28780
rect 4557 28958 4603 29005
rect 4557 28924 4563 28958
rect 4597 28924 4603 28958
rect 4557 28886 4603 28924
rect 4557 28852 4563 28886
rect 4597 28852 4603 28886
rect 4557 28814 4603 28852
rect 4557 28780 4563 28814
rect 4597 28780 4603 28814
rect 4557 28733 4603 28780
rect 4653 28958 4699 29005
rect 4653 28924 4659 28958
rect 4693 28924 4699 28958
rect 4653 28886 4699 28924
rect 4653 28852 4659 28886
rect 4693 28852 4699 28886
rect 4653 28814 4699 28852
rect 4653 28780 4659 28814
rect 4693 28780 4699 28814
rect 4653 28733 4699 28780
rect 4749 28958 4795 29005
rect 4749 28924 4755 28958
rect 4789 28924 4795 28958
rect 4749 28886 4795 28924
rect 4749 28852 4755 28886
rect 4789 28852 4795 28886
rect 4749 28814 4795 28852
rect 4749 28780 4755 28814
rect 4789 28780 4795 28814
rect 4749 28733 4795 28780
rect 4845 28958 4891 29005
rect 4845 28924 4851 28958
rect 4885 28924 4891 28958
rect 4845 28886 4891 28924
rect 4845 28852 4851 28886
rect 4885 28852 4891 28886
rect 4845 28814 4891 28852
rect 4845 28780 4851 28814
rect 4885 28780 4891 28814
rect 4845 28733 4891 28780
rect 4941 28958 4987 29005
rect 4941 28924 4947 28958
rect 4981 28924 4987 28958
rect 4941 28886 4987 28924
rect 4941 28852 4947 28886
rect 4981 28852 4987 28886
rect 4941 28814 4987 28852
rect 4941 28780 4947 28814
rect 4981 28780 4987 28814
rect 4941 28733 4987 28780
rect 5055 28989 5101 29027
rect 5055 28955 5061 28989
rect 5095 28955 5101 28989
rect 5055 28917 5101 28955
rect 5055 28883 5061 28917
rect 5095 28886 5101 28917
rect 5274 28886 5550 28887
rect 5095 28883 5550 28886
rect 5055 28856 5550 28883
rect 5055 28845 5303 28856
rect 5055 28811 5061 28845
rect 5095 28822 5303 28845
rect 5337 28822 5395 28856
rect 5429 28822 5487 28856
rect 5521 28822 5550 28856
rect 5095 28811 5550 28822
rect 5055 28791 5550 28811
rect 5055 28773 5101 28791
rect 5055 28739 5061 28773
rect 5095 28739 5101 28773
rect 2466 28558 3837 28592
rect 2466 28425 2500 28558
rect 2658 28425 2692 28558
rect 2850 28425 2884 28558
rect 3042 28425 3076 28558
rect 3234 28425 3268 28558
rect 3426 28425 3460 28558
rect 3671 28468 3681 28520
rect 3733 28468 3743 28520
rect 3679 28467 3691 28468
rect 3725 28467 3737 28468
rect 3679 28461 3737 28467
rect 3534 28432 3580 28455
rect 2460 28390 2506 28425
rect 2460 28356 2466 28390
rect 2500 28356 2506 28390
rect 2460 28321 2506 28356
rect 2556 28390 2602 28425
rect 2556 28356 2562 28390
rect 2596 28356 2602 28390
rect 2556 28321 2602 28356
rect 2652 28390 2698 28425
rect 2652 28356 2658 28390
rect 2692 28356 2698 28390
rect 2652 28321 2698 28356
rect 2748 28390 2794 28425
rect 2748 28356 2754 28390
rect 2788 28356 2794 28390
rect 2748 28321 2794 28356
rect 2844 28390 2890 28425
rect 2844 28356 2850 28390
rect 2884 28356 2890 28390
rect 2844 28321 2890 28356
rect 2940 28390 2986 28425
rect 2940 28356 2946 28390
rect 2980 28356 2986 28390
rect 2940 28321 2986 28356
rect 3036 28390 3082 28425
rect 3036 28356 3042 28390
rect 3076 28356 3082 28390
rect 3036 28321 3082 28356
rect 3132 28390 3178 28425
rect 3132 28356 3138 28390
rect 3172 28356 3178 28390
rect 3132 28321 3178 28356
rect 3228 28390 3274 28425
rect 3228 28356 3234 28390
rect 3268 28356 3274 28390
rect 3228 28321 3274 28356
rect 3324 28390 3370 28425
rect 3324 28356 3330 28390
rect 3364 28356 3370 28390
rect 3324 28321 3370 28356
rect 3420 28390 3466 28425
rect 3420 28356 3426 28390
rect 3460 28356 3466 28390
rect 3420 28321 3466 28356
rect 3534 28398 3540 28432
rect 3574 28430 3580 28432
rect 3803 28430 3837 28558
rect 3574 28429 3680 28430
rect 3734 28429 3837 28430
rect 3574 28417 3687 28429
rect 3574 28398 3647 28417
rect 3534 28360 3647 28398
rect 3534 28326 3540 28360
rect 3574 28341 3647 28360
rect 3681 28341 3687 28417
rect 3574 28330 3687 28341
rect 3574 28326 3580 28330
rect 3641 28329 3687 28330
rect 3729 28417 3837 28429
rect 3987 28592 4021 28733
rect 4179 28592 4213 28733
rect 4371 28592 4405 28733
rect 4563 28592 4597 28733
rect 4755 28592 4789 28733
rect 4947 28592 4981 28733
rect 5055 28695 5101 28739
rect 5683 28646 5743 29899
rect 5177 28612 5743 28646
rect 5177 28592 5211 28612
rect 3987 28558 5211 28592
rect 3987 28425 4021 28558
rect 4179 28425 4213 28558
rect 4371 28425 4405 28558
rect 4563 28425 4597 28558
rect 4755 28425 4789 28558
rect 4947 28425 4981 28558
rect 5438 28554 5512 28555
rect 5326 28552 5400 28553
rect 5326 28500 5337 28552
rect 5389 28500 5400 28552
rect 5438 28502 5449 28554
rect 5501 28502 5512 28554
rect 5438 28501 5512 28502
rect 5326 28499 5400 28500
rect 5055 28432 5101 28455
rect 3729 28341 3735 28417
rect 3769 28341 3837 28417
rect 3729 28330 3837 28341
rect 3729 28329 3775 28330
rect 2450 28290 2516 28293
rect 2447 28238 2457 28290
rect 2509 28238 2519 28290
rect 2450 28233 2516 28238
rect 2562 28181 2596 28321
rect 2642 28290 2708 28293
rect 2638 28238 2648 28290
rect 2700 28238 2710 28290
rect 2642 28233 2708 28238
rect 2754 28181 2788 28321
rect 2834 28290 2900 28293
rect 2830 28238 2840 28290
rect 2892 28238 2902 28290
rect 2834 28233 2900 28238
rect 2946 28181 2980 28321
rect 3026 28290 3092 28293
rect 3022 28238 3032 28290
rect 3084 28238 3094 28290
rect 3026 28233 3092 28238
rect 3138 28181 3172 28321
rect 3218 28289 3284 28293
rect 3215 28237 3225 28289
rect 3277 28237 3287 28289
rect 3218 28233 3284 28237
rect 3330 28181 3364 28321
rect 3410 28289 3476 28293
rect 3407 28237 3417 28289
rect 3469 28237 3479 28289
rect 3534 28288 3580 28326
rect 3534 28254 3540 28288
rect 3574 28254 3580 28288
rect 3410 28233 3476 28237
rect 2282 28147 3364 28181
rect 3534 28071 3580 28254
rect 3803 28181 3837 28330
rect 3981 28390 4027 28425
rect 3981 28356 3987 28390
rect 4021 28356 4027 28390
rect 3981 28321 4027 28356
rect 4077 28390 4123 28425
rect 4077 28356 4083 28390
rect 4117 28356 4123 28390
rect 4077 28321 4123 28356
rect 4173 28390 4219 28425
rect 4173 28356 4179 28390
rect 4213 28356 4219 28390
rect 4173 28321 4219 28356
rect 4269 28390 4315 28425
rect 4269 28356 4275 28390
rect 4309 28356 4315 28390
rect 4269 28321 4315 28356
rect 4365 28390 4411 28425
rect 4365 28356 4371 28390
rect 4405 28356 4411 28390
rect 4365 28321 4411 28356
rect 4461 28390 4507 28425
rect 4461 28356 4467 28390
rect 4501 28356 4507 28390
rect 4461 28321 4507 28356
rect 4557 28390 4603 28425
rect 4557 28356 4563 28390
rect 4597 28356 4603 28390
rect 4557 28321 4603 28356
rect 4653 28390 4699 28425
rect 4653 28356 4659 28390
rect 4693 28356 4699 28390
rect 4653 28321 4699 28356
rect 4749 28390 4795 28425
rect 4749 28356 4755 28390
rect 4789 28356 4795 28390
rect 4749 28321 4795 28356
rect 4845 28390 4891 28425
rect 4845 28356 4851 28390
rect 4885 28356 4891 28390
rect 4845 28321 4891 28356
rect 4941 28390 4987 28425
rect 4941 28356 4947 28390
rect 4981 28356 4987 28390
rect 4941 28321 4987 28356
rect 5055 28398 5061 28432
rect 5095 28398 5101 28432
rect 5055 28360 5101 28398
rect 5055 28326 5061 28360
rect 5095 28343 5101 28360
rect 5095 28326 5550 28343
rect 3971 28290 4037 28293
rect 3968 28238 3978 28290
rect 4030 28238 4040 28290
rect 3971 28233 4037 28238
rect 4083 28181 4117 28321
rect 4163 28290 4229 28293
rect 4159 28238 4169 28290
rect 4221 28238 4231 28290
rect 4163 28233 4229 28238
rect 4275 28181 4309 28321
rect 4355 28290 4421 28293
rect 4351 28238 4361 28290
rect 4413 28238 4423 28290
rect 4355 28233 4421 28238
rect 4467 28181 4501 28321
rect 4547 28290 4613 28293
rect 4543 28238 4553 28290
rect 4605 28238 4615 28290
rect 4547 28233 4613 28238
rect 4659 28181 4693 28321
rect 4739 28289 4805 28293
rect 4736 28237 4746 28289
rect 4798 28237 4808 28289
rect 4739 28233 4805 28237
rect 4851 28181 4885 28321
rect 5055 28312 5550 28326
rect 4931 28289 4997 28293
rect 4928 28237 4938 28289
rect 4990 28237 5000 28289
rect 5055 28288 5303 28312
rect 5055 28254 5061 28288
rect 5095 28278 5303 28288
rect 5337 28278 5395 28312
rect 5429 28278 5487 28312
rect 5521 28278 5550 28312
rect 5095 28254 5550 28278
rect 5055 28247 5550 28254
rect 4931 28233 4997 28237
rect 3803 28147 4885 28181
rect 5055 28072 5101 28247
rect 129 27864 1211 27898
rect 129 27301 163 27864
rect 294 27754 304 27806
rect 356 27754 366 27806
rect 409 27714 443 27864
rect 487 27754 497 27806
rect 549 27754 559 27806
rect 601 27714 635 27864
rect 678 27754 688 27806
rect 740 27754 750 27806
rect 793 27714 827 27864
rect 870 27754 880 27806
rect 932 27754 942 27806
rect 985 27714 1019 27864
rect 1062 27754 1072 27806
rect 1124 27754 1134 27806
rect 1177 27714 1211 27864
rect 1254 27754 1264 27806
rect 1316 27754 1326 27806
rect 1381 27770 1427 27934
rect 2282 27868 3364 27902
rect 1381 27736 1387 27770
rect 1421 27736 1427 27770
rect 1512 27747 1522 27807
rect 1578 27747 1792 27807
rect 1852 27747 1862 27807
rect 307 27667 353 27714
rect 307 27633 313 27667
rect 347 27633 353 27667
rect 307 27595 353 27633
rect 307 27561 313 27595
rect 347 27561 353 27595
rect 307 27523 353 27561
rect 307 27489 313 27523
rect 347 27489 353 27523
rect 307 27442 353 27489
rect 403 27667 449 27714
rect 403 27633 409 27667
rect 443 27633 449 27667
rect 403 27595 449 27633
rect 403 27561 409 27595
rect 443 27561 449 27595
rect 403 27523 449 27561
rect 403 27489 409 27523
rect 443 27489 449 27523
rect 403 27442 449 27489
rect 499 27667 545 27714
rect 499 27633 505 27667
rect 539 27633 545 27667
rect 499 27595 545 27633
rect 499 27561 505 27595
rect 539 27561 545 27595
rect 499 27523 545 27561
rect 499 27489 505 27523
rect 539 27489 545 27523
rect 499 27442 545 27489
rect 595 27667 641 27714
rect 595 27633 601 27667
rect 635 27633 641 27667
rect 595 27595 641 27633
rect 595 27561 601 27595
rect 635 27561 641 27595
rect 595 27523 641 27561
rect 595 27489 601 27523
rect 635 27489 641 27523
rect 595 27442 641 27489
rect 691 27667 737 27714
rect 691 27633 697 27667
rect 731 27633 737 27667
rect 691 27595 737 27633
rect 691 27561 697 27595
rect 731 27561 737 27595
rect 691 27523 737 27561
rect 691 27489 697 27523
rect 731 27489 737 27523
rect 691 27442 737 27489
rect 787 27667 833 27714
rect 787 27633 793 27667
rect 827 27633 833 27667
rect 787 27595 833 27633
rect 787 27561 793 27595
rect 827 27561 833 27595
rect 787 27523 833 27561
rect 787 27489 793 27523
rect 827 27489 833 27523
rect 787 27442 833 27489
rect 883 27667 929 27714
rect 883 27633 889 27667
rect 923 27633 929 27667
rect 883 27595 929 27633
rect 883 27561 889 27595
rect 923 27561 929 27595
rect 883 27523 929 27561
rect 883 27489 889 27523
rect 923 27489 929 27523
rect 883 27442 929 27489
rect 979 27667 1025 27714
rect 979 27633 985 27667
rect 1019 27633 1025 27667
rect 979 27595 1025 27633
rect 979 27561 985 27595
rect 1019 27561 1025 27595
rect 979 27523 1025 27561
rect 979 27489 985 27523
rect 1019 27489 1025 27523
rect 979 27442 1025 27489
rect 1075 27667 1121 27714
rect 1075 27633 1081 27667
rect 1115 27633 1121 27667
rect 1075 27595 1121 27633
rect 1075 27561 1081 27595
rect 1115 27561 1121 27595
rect 1075 27523 1121 27561
rect 1075 27489 1081 27523
rect 1115 27489 1121 27523
rect 1075 27442 1121 27489
rect 1171 27667 1217 27714
rect 1171 27633 1177 27667
rect 1211 27633 1217 27667
rect 1171 27595 1217 27633
rect 1171 27561 1177 27595
rect 1211 27561 1217 27595
rect 1171 27523 1217 27561
rect 1171 27489 1177 27523
rect 1211 27489 1217 27523
rect 1171 27442 1217 27489
rect 1267 27667 1313 27714
rect 1267 27633 1273 27667
rect 1307 27633 1313 27667
rect 1267 27595 1313 27633
rect 1267 27561 1273 27595
rect 1307 27561 1313 27595
rect 1267 27523 1313 27561
rect 1267 27489 1273 27523
rect 1307 27489 1313 27523
rect 1267 27442 1313 27489
rect 1381 27698 1427 27736
rect 1381 27664 1387 27698
rect 1421 27664 1427 27698
rect 1381 27626 1427 27664
rect 1381 27592 1387 27626
rect 1421 27592 1427 27626
rect 1381 27554 1427 27592
rect 1381 27520 1387 27554
rect 1421 27520 1427 27554
rect 1381 27510 1427 27520
rect 1381 27508 2160 27510
rect 1381 27482 2056 27508
rect 1381 27457 1387 27482
rect 1380 27448 1387 27457
rect 1421 27448 2056 27482
rect 0 27267 163 27301
rect 129 26890 163 27267
rect 313 27301 347 27442
rect 505 27301 539 27442
rect 697 27301 731 27442
rect 889 27301 923 27442
rect 1081 27301 1115 27442
rect 1273 27301 1307 27442
rect 1380 27400 2056 27448
rect 2190 27400 2200 27508
rect 1380 27398 2160 27400
rect 2282 27305 2316 27868
rect 2447 27758 2457 27810
rect 2509 27758 2519 27810
rect 2562 27718 2596 27868
rect 2640 27758 2650 27810
rect 2702 27758 2712 27810
rect 2754 27718 2788 27868
rect 2831 27758 2841 27810
rect 2893 27758 2903 27810
rect 2946 27718 2980 27868
rect 3023 27758 3033 27810
rect 3085 27758 3095 27810
rect 3138 27718 3172 27868
rect 3215 27758 3225 27810
rect 3277 27758 3287 27810
rect 3330 27718 3364 27868
rect 3407 27758 3417 27810
rect 3469 27758 3479 27810
rect 3534 27774 3580 27982
rect 3534 27740 3540 27774
rect 3574 27740 3580 27774
rect 2460 27671 2506 27718
rect 2460 27637 2466 27671
rect 2500 27637 2506 27671
rect 2460 27599 2506 27637
rect 2460 27565 2466 27599
rect 2500 27565 2506 27599
rect 2460 27527 2506 27565
rect 2460 27493 2466 27527
rect 2500 27493 2506 27527
rect 2460 27446 2506 27493
rect 2556 27671 2602 27718
rect 2556 27637 2562 27671
rect 2596 27637 2602 27671
rect 2556 27599 2602 27637
rect 2556 27565 2562 27599
rect 2596 27565 2602 27599
rect 2556 27527 2602 27565
rect 2556 27493 2562 27527
rect 2596 27493 2602 27527
rect 2556 27446 2602 27493
rect 2652 27671 2698 27718
rect 2652 27637 2658 27671
rect 2692 27637 2698 27671
rect 2652 27599 2698 27637
rect 2652 27565 2658 27599
rect 2692 27565 2698 27599
rect 2652 27527 2698 27565
rect 2652 27493 2658 27527
rect 2692 27493 2698 27527
rect 2652 27446 2698 27493
rect 2748 27671 2794 27718
rect 2748 27637 2754 27671
rect 2788 27637 2794 27671
rect 2748 27599 2794 27637
rect 2748 27565 2754 27599
rect 2788 27565 2794 27599
rect 2748 27527 2794 27565
rect 2748 27493 2754 27527
rect 2788 27493 2794 27527
rect 2748 27446 2794 27493
rect 2844 27671 2890 27718
rect 2844 27637 2850 27671
rect 2884 27637 2890 27671
rect 2844 27599 2890 27637
rect 2844 27565 2850 27599
rect 2884 27565 2890 27599
rect 2844 27527 2890 27565
rect 2844 27493 2850 27527
rect 2884 27493 2890 27527
rect 2844 27446 2890 27493
rect 2940 27671 2986 27718
rect 2940 27637 2946 27671
rect 2980 27637 2986 27671
rect 2940 27599 2986 27637
rect 2940 27565 2946 27599
rect 2980 27565 2986 27599
rect 2940 27527 2986 27565
rect 2940 27493 2946 27527
rect 2980 27493 2986 27527
rect 2940 27446 2986 27493
rect 3036 27671 3082 27718
rect 3036 27637 3042 27671
rect 3076 27637 3082 27671
rect 3036 27599 3082 27637
rect 3036 27565 3042 27599
rect 3076 27565 3082 27599
rect 3036 27527 3082 27565
rect 3036 27493 3042 27527
rect 3076 27493 3082 27527
rect 3036 27446 3082 27493
rect 3132 27671 3178 27718
rect 3132 27637 3138 27671
rect 3172 27637 3178 27671
rect 3132 27599 3178 27637
rect 3132 27565 3138 27599
rect 3172 27565 3178 27599
rect 3132 27527 3178 27565
rect 3132 27493 3138 27527
rect 3172 27493 3178 27527
rect 3132 27446 3178 27493
rect 3228 27671 3274 27718
rect 3228 27637 3234 27671
rect 3268 27637 3274 27671
rect 3228 27599 3274 27637
rect 3228 27565 3234 27599
rect 3268 27565 3274 27599
rect 3228 27527 3274 27565
rect 3228 27493 3234 27527
rect 3268 27493 3274 27527
rect 3228 27446 3274 27493
rect 3324 27671 3370 27718
rect 3324 27637 3330 27671
rect 3364 27637 3370 27671
rect 3324 27599 3370 27637
rect 3324 27565 3330 27599
rect 3364 27565 3370 27599
rect 3324 27527 3370 27565
rect 3324 27493 3330 27527
rect 3364 27493 3370 27527
rect 3324 27446 3370 27493
rect 3420 27671 3466 27718
rect 3420 27637 3426 27671
rect 3460 27637 3466 27671
rect 3420 27599 3466 27637
rect 3420 27565 3426 27599
rect 3460 27565 3466 27599
rect 3420 27527 3466 27565
rect 3420 27493 3426 27527
rect 3460 27493 3466 27527
rect 3420 27446 3466 27493
rect 3534 27702 3580 27740
rect 3534 27668 3540 27702
rect 3574 27668 3580 27702
rect 3534 27630 3580 27668
rect 3534 27596 3540 27630
rect 3574 27596 3580 27630
rect 3534 27558 3580 27596
rect 3534 27524 3540 27558
rect 3574 27524 3580 27558
rect 3534 27486 3580 27524
rect 3534 27452 3540 27486
rect 3574 27452 3580 27486
rect 2101 27301 2316 27305
rect 313 27271 2316 27301
rect 313 27267 2141 27271
rect 313 27134 347 27267
rect 505 27134 539 27267
rect 697 27134 731 27267
rect 889 27134 923 27267
rect 1081 27134 1115 27267
rect 1273 27134 1307 27267
rect 1381 27141 1608 27164
rect 307 27099 353 27134
rect 307 27065 313 27099
rect 347 27065 353 27099
rect 307 27030 353 27065
rect 403 27099 449 27134
rect 403 27065 409 27099
rect 443 27065 449 27099
rect 403 27030 449 27065
rect 499 27099 545 27134
rect 499 27065 505 27099
rect 539 27065 545 27099
rect 499 27030 545 27065
rect 595 27099 641 27134
rect 595 27065 601 27099
rect 635 27065 641 27099
rect 595 27030 641 27065
rect 691 27099 737 27134
rect 691 27065 697 27099
rect 731 27065 737 27099
rect 691 27030 737 27065
rect 787 27099 833 27134
rect 787 27065 793 27099
rect 827 27065 833 27099
rect 787 27030 833 27065
rect 883 27099 929 27134
rect 883 27065 889 27099
rect 923 27065 929 27099
rect 883 27030 929 27065
rect 979 27099 1025 27134
rect 979 27065 985 27099
rect 1019 27065 1025 27099
rect 979 27030 1025 27065
rect 1075 27099 1121 27134
rect 1075 27065 1081 27099
rect 1115 27065 1121 27099
rect 1075 27030 1121 27065
rect 1171 27099 1217 27134
rect 1171 27065 1177 27099
rect 1211 27065 1217 27099
rect 1171 27030 1217 27065
rect 1267 27099 1313 27134
rect 1267 27065 1273 27099
rect 1307 27065 1313 27099
rect 1267 27030 1313 27065
rect 1381 27107 1387 27141
rect 1421 27107 1608 27141
rect 1381 27069 1608 27107
rect 1381 27035 1387 27069
rect 1421 27044 1608 27069
rect 1421 27035 1427 27044
rect 1560 27042 1608 27044
rect 1598 27040 1608 27042
rect 1720 27040 1730 27164
rect 297 26999 363 27002
rect 294 26947 304 26999
rect 356 26947 366 26999
rect 297 26942 363 26947
rect 409 26890 443 27030
rect 489 26999 555 27002
rect 485 26947 495 26999
rect 547 26947 557 26999
rect 489 26942 555 26947
rect 601 26890 635 27030
rect 681 26999 747 27002
rect 677 26947 687 26999
rect 739 26947 749 26999
rect 681 26942 747 26947
rect 793 26890 827 27030
rect 873 26999 939 27002
rect 869 26947 879 26999
rect 931 26947 941 26999
rect 873 26942 939 26947
rect 985 26890 1019 27030
rect 1065 26998 1131 27002
rect 1062 26946 1072 26998
rect 1124 26946 1134 26998
rect 1065 26942 1131 26946
rect 1177 26890 1211 27030
rect 1257 26998 1323 27002
rect 1254 26946 1264 26998
rect 1316 26946 1326 26998
rect 1381 26997 1427 27035
rect 1920 27002 1930 27004
rect 1381 26963 1387 26997
rect 1421 26963 1427 26997
rect 1257 26942 1323 26946
rect 129 26856 1211 26890
rect 1381 26820 1427 26963
rect 1458 26946 1468 27002
rect 1524 26948 1930 27002
rect 1986 26948 1996 27004
rect 1524 26946 1986 26948
rect 2282 26894 2316 27271
rect 2466 27305 2500 27446
rect 2658 27305 2692 27446
rect 2850 27305 2884 27446
rect 3042 27305 3076 27446
rect 3234 27305 3268 27446
rect 3426 27305 3460 27446
rect 3534 27408 3580 27452
rect 3803 27868 4885 27902
rect 3803 27305 3837 27868
rect 3968 27758 3978 27810
rect 4030 27758 4040 27810
rect 4083 27718 4117 27868
rect 4161 27758 4171 27810
rect 4223 27758 4233 27810
rect 4275 27718 4309 27868
rect 4352 27758 4362 27810
rect 4414 27758 4424 27810
rect 4467 27718 4501 27868
rect 4544 27758 4554 27810
rect 4606 27758 4616 27810
rect 4659 27718 4693 27868
rect 4736 27758 4746 27810
rect 4798 27758 4808 27810
rect 4851 27718 4885 27868
rect 4928 27758 4938 27810
rect 4990 27758 5000 27810
rect 5055 27774 5101 27979
rect 5055 27740 5061 27774
rect 5095 27740 5101 27774
rect 3981 27671 4027 27718
rect 3981 27637 3987 27671
rect 4021 27637 4027 27671
rect 3981 27599 4027 27637
rect 3981 27565 3987 27599
rect 4021 27565 4027 27599
rect 3981 27527 4027 27565
rect 3981 27493 3987 27527
rect 4021 27493 4027 27527
rect 3981 27446 4027 27493
rect 4077 27671 4123 27718
rect 4077 27637 4083 27671
rect 4117 27637 4123 27671
rect 4077 27599 4123 27637
rect 4077 27565 4083 27599
rect 4117 27565 4123 27599
rect 4077 27527 4123 27565
rect 4077 27493 4083 27527
rect 4117 27493 4123 27527
rect 4077 27446 4123 27493
rect 4173 27671 4219 27718
rect 4173 27637 4179 27671
rect 4213 27637 4219 27671
rect 4173 27599 4219 27637
rect 4173 27565 4179 27599
rect 4213 27565 4219 27599
rect 4173 27527 4219 27565
rect 4173 27493 4179 27527
rect 4213 27493 4219 27527
rect 4173 27446 4219 27493
rect 4269 27671 4315 27718
rect 4269 27637 4275 27671
rect 4309 27637 4315 27671
rect 4269 27599 4315 27637
rect 4269 27565 4275 27599
rect 4309 27565 4315 27599
rect 4269 27527 4315 27565
rect 4269 27493 4275 27527
rect 4309 27493 4315 27527
rect 4269 27446 4315 27493
rect 4365 27671 4411 27718
rect 4365 27637 4371 27671
rect 4405 27637 4411 27671
rect 4365 27599 4411 27637
rect 4365 27565 4371 27599
rect 4405 27565 4411 27599
rect 4365 27527 4411 27565
rect 4365 27493 4371 27527
rect 4405 27493 4411 27527
rect 4365 27446 4411 27493
rect 4461 27671 4507 27718
rect 4461 27637 4467 27671
rect 4501 27637 4507 27671
rect 4461 27599 4507 27637
rect 4461 27565 4467 27599
rect 4501 27565 4507 27599
rect 4461 27527 4507 27565
rect 4461 27493 4467 27527
rect 4501 27493 4507 27527
rect 4461 27446 4507 27493
rect 4557 27671 4603 27718
rect 4557 27637 4563 27671
rect 4597 27637 4603 27671
rect 4557 27599 4603 27637
rect 4557 27565 4563 27599
rect 4597 27565 4603 27599
rect 4557 27527 4603 27565
rect 4557 27493 4563 27527
rect 4597 27493 4603 27527
rect 4557 27446 4603 27493
rect 4653 27671 4699 27718
rect 4653 27637 4659 27671
rect 4693 27637 4699 27671
rect 4653 27599 4699 27637
rect 4653 27565 4659 27599
rect 4693 27565 4699 27599
rect 4653 27527 4699 27565
rect 4653 27493 4659 27527
rect 4693 27493 4699 27527
rect 4653 27446 4699 27493
rect 4749 27671 4795 27718
rect 4749 27637 4755 27671
rect 4789 27637 4795 27671
rect 4749 27599 4795 27637
rect 4749 27565 4755 27599
rect 4789 27565 4795 27599
rect 4749 27527 4795 27565
rect 4749 27493 4755 27527
rect 4789 27493 4795 27527
rect 4749 27446 4795 27493
rect 4845 27671 4891 27718
rect 4845 27637 4851 27671
rect 4885 27637 4891 27671
rect 4845 27599 4891 27637
rect 4845 27565 4851 27599
rect 4885 27565 4891 27599
rect 4845 27527 4891 27565
rect 4845 27493 4851 27527
rect 4885 27493 4891 27527
rect 4845 27446 4891 27493
rect 4941 27671 4987 27718
rect 4941 27637 4947 27671
rect 4981 27637 4987 27671
rect 4941 27599 4987 27637
rect 4941 27565 4947 27599
rect 4981 27565 4987 27599
rect 4941 27527 4987 27565
rect 4941 27493 4947 27527
rect 4981 27493 4987 27527
rect 4941 27446 4987 27493
rect 5055 27702 5101 27740
rect 5055 27668 5061 27702
rect 5095 27668 5101 27702
rect 5055 27630 5101 27668
rect 5055 27596 5061 27630
rect 5095 27599 5101 27630
rect 5274 27599 5550 27600
rect 5095 27596 5550 27599
rect 5055 27569 5550 27596
rect 5055 27558 5303 27569
rect 5055 27524 5061 27558
rect 5095 27535 5303 27558
rect 5337 27535 5395 27569
rect 5429 27535 5487 27569
rect 5521 27535 5550 27569
rect 5095 27524 5550 27535
rect 5055 27504 5550 27524
rect 5055 27486 5101 27504
rect 5055 27452 5061 27486
rect 5095 27452 5101 27486
rect 2466 27271 3837 27305
rect 2466 27138 2500 27271
rect 2658 27138 2692 27271
rect 2850 27138 2884 27271
rect 3042 27138 3076 27271
rect 3234 27138 3268 27271
rect 3426 27138 3460 27271
rect 3671 27181 3681 27233
rect 3733 27181 3743 27233
rect 3679 27180 3691 27181
rect 3725 27180 3737 27181
rect 3679 27174 3737 27180
rect 3534 27145 3580 27168
rect 2460 27103 2506 27138
rect 2460 27069 2466 27103
rect 2500 27069 2506 27103
rect 2460 27034 2506 27069
rect 2556 27103 2602 27138
rect 2556 27069 2562 27103
rect 2596 27069 2602 27103
rect 2556 27034 2602 27069
rect 2652 27103 2698 27138
rect 2652 27069 2658 27103
rect 2692 27069 2698 27103
rect 2652 27034 2698 27069
rect 2748 27103 2794 27138
rect 2748 27069 2754 27103
rect 2788 27069 2794 27103
rect 2748 27034 2794 27069
rect 2844 27103 2890 27138
rect 2844 27069 2850 27103
rect 2884 27069 2890 27103
rect 2844 27034 2890 27069
rect 2940 27103 2986 27138
rect 2940 27069 2946 27103
rect 2980 27069 2986 27103
rect 2940 27034 2986 27069
rect 3036 27103 3082 27138
rect 3036 27069 3042 27103
rect 3076 27069 3082 27103
rect 3036 27034 3082 27069
rect 3132 27103 3178 27138
rect 3132 27069 3138 27103
rect 3172 27069 3178 27103
rect 3132 27034 3178 27069
rect 3228 27103 3274 27138
rect 3228 27069 3234 27103
rect 3268 27069 3274 27103
rect 3228 27034 3274 27069
rect 3324 27103 3370 27138
rect 3324 27069 3330 27103
rect 3364 27069 3370 27103
rect 3324 27034 3370 27069
rect 3420 27103 3466 27138
rect 3420 27069 3426 27103
rect 3460 27069 3466 27103
rect 3420 27034 3466 27069
rect 3534 27111 3540 27145
rect 3574 27143 3580 27145
rect 3803 27143 3837 27271
rect 3574 27142 3680 27143
rect 3734 27142 3837 27143
rect 3574 27130 3687 27142
rect 3574 27111 3647 27130
rect 3534 27073 3647 27111
rect 3534 27039 3540 27073
rect 3574 27054 3647 27073
rect 3681 27054 3687 27130
rect 3574 27043 3687 27054
rect 3574 27039 3580 27043
rect 3641 27042 3687 27043
rect 3729 27130 3837 27142
rect 3987 27305 4021 27446
rect 4179 27305 4213 27446
rect 4371 27305 4405 27446
rect 4563 27305 4597 27446
rect 4755 27305 4789 27446
rect 4947 27305 4981 27446
rect 5055 27408 5101 27452
rect 5683 27359 5743 28612
rect 5177 27325 5743 27359
rect 5177 27305 5211 27325
rect 3987 27271 5211 27305
rect 3987 27138 4021 27271
rect 4179 27138 4213 27271
rect 4371 27138 4405 27271
rect 4563 27138 4597 27271
rect 4755 27138 4789 27271
rect 4947 27138 4981 27271
rect 5438 27267 5512 27268
rect 5326 27265 5400 27266
rect 5326 27213 5337 27265
rect 5389 27213 5400 27265
rect 5438 27215 5449 27267
rect 5501 27215 5512 27267
rect 5438 27214 5512 27215
rect 5326 27212 5400 27213
rect 5055 27145 5101 27168
rect 3729 27054 3735 27130
rect 3769 27054 3837 27130
rect 3729 27043 3837 27054
rect 3729 27042 3775 27043
rect 2450 27003 2516 27006
rect 2447 26951 2457 27003
rect 2509 26951 2519 27003
rect 2450 26946 2516 26951
rect 2562 26894 2596 27034
rect 2642 27003 2708 27006
rect 2638 26951 2648 27003
rect 2700 26951 2710 27003
rect 2642 26946 2708 26951
rect 2754 26894 2788 27034
rect 2834 27003 2900 27006
rect 2830 26951 2840 27003
rect 2892 26951 2902 27003
rect 2834 26946 2900 26951
rect 2946 26894 2980 27034
rect 3026 27003 3092 27006
rect 3022 26951 3032 27003
rect 3084 26951 3094 27003
rect 3026 26946 3092 26951
rect 3138 26894 3172 27034
rect 3218 27002 3284 27006
rect 3215 26950 3225 27002
rect 3277 26950 3287 27002
rect 3218 26946 3284 26950
rect 3330 26894 3364 27034
rect 3410 27002 3476 27006
rect 3407 26950 3417 27002
rect 3469 26950 3479 27002
rect 3534 27001 3580 27039
rect 3534 26967 3540 27001
rect 3574 26967 3580 27001
rect 3410 26946 3476 26950
rect 2282 26860 3364 26894
rect 3534 26784 3580 26967
rect 3803 26894 3837 27043
rect 3981 27103 4027 27138
rect 3981 27069 3987 27103
rect 4021 27069 4027 27103
rect 3981 27034 4027 27069
rect 4077 27103 4123 27138
rect 4077 27069 4083 27103
rect 4117 27069 4123 27103
rect 4077 27034 4123 27069
rect 4173 27103 4219 27138
rect 4173 27069 4179 27103
rect 4213 27069 4219 27103
rect 4173 27034 4219 27069
rect 4269 27103 4315 27138
rect 4269 27069 4275 27103
rect 4309 27069 4315 27103
rect 4269 27034 4315 27069
rect 4365 27103 4411 27138
rect 4365 27069 4371 27103
rect 4405 27069 4411 27103
rect 4365 27034 4411 27069
rect 4461 27103 4507 27138
rect 4461 27069 4467 27103
rect 4501 27069 4507 27103
rect 4461 27034 4507 27069
rect 4557 27103 4603 27138
rect 4557 27069 4563 27103
rect 4597 27069 4603 27103
rect 4557 27034 4603 27069
rect 4653 27103 4699 27138
rect 4653 27069 4659 27103
rect 4693 27069 4699 27103
rect 4653 27034 4699 27069
rect 4749 27103 4795 27138
rect 4749 27069 4755 27103
rect 4789 27069 4795 27103
rect 4749 27034 4795 27069
rect 4845 27103 4891 27138
rect 4845 27069 4851 27103
rect 4885 27069 4891 27103
rect 4845 27034 4891 27069
rect 4941 27103 4987 27138
rect 4941 27069 4947 27103
rect 4981 27069 4987 27103
rect 4941 27034 4987 27069
rect 5055 27111 5061 27145
rect 5095 27111 5101 27145
rect 5055 27073 5101 27111
rect 5055 27039 5061 27073
rect 5095 27056 5101 27073
rect 5095 27039 5550 27056
rect 3971 27003 4037 27006
rect 3968 26951 3978 27003
rect 4030 26951 4040 27003
rect 3971 26946 4037 26951
rect 4083 26894 4117 27034
rect 4163 27003 4229 27006
rect 4159 26951 4169 27003
rect 4221 26951 4231 27003
rect 4163 26946 4229 26951
rect 4275 26894 4309 27034
rect 4355 27003 4421 27006
rect 4351 26951 4361 27003
rect 4413 26951 4423 27003
rect 4355 26946 4421 26951
rect 4467 26894 4501 27034
rect 4547 27003 4613 27006
rect 4543 26951 4553 27003
rect 4605 26951 4615 27003
rect 4547 26946 4613 26951
rect 4659 26894 4693 27034
rect 4739 27002 4805 27006
rect 4736 26950 4746 27002
rect 4798 26950 4808 27002
rect 4739 26946 4805 26950
rect 4851 26894 4885 27034
rect 5055 27025 5550 27039
rect 4931 27002 4997 27006
rect 4928 26950 4938 27002
rect 4990 26950 5000 27002
rect 5055 27001 5303 27025
rect 5055 26967 5061 27001
rect 5095 26991 5303 27001
rect 5337 26991 5395 27025
rect 5429 26991 5487 27025
rect 5521 26991 5550 27025
rect 5095 26967 5550 26991
rect 5055 26960 5550 26967
rect 4931 26946 4997 26950
rect 3803 26860 4885 26894
rect 5055 26785 5101 26960
rect 129 26577 1211 26611
rect 129 26014 163 26577
rect 294 26467 304 26519
rect 356 26467 366 26519
rect 409 26427 443 26577
rect 487 26467 497 26519
rect 549 26467 559 26519
rect 601 26427 635 26577
rect 678 26467 688 26519
rect 740 26467 750 26519
rect 793 26427 827 26577
rect 870 26467 880 26519
rect 932 26467 942 26519
rect 985 26427 1019 26577
rect 1062 26467 1072 26519
rect 1124 26467 1134 26519
rect 1177 26427 1211 26577
rect 1254 26467 1264 26519
rect 1316 26467 1326 26519
rect 1381 26483 1427 26647
rect 2282 26581 3364 26615
rect 1381 26449 1387 26483
rect 1421 26449 1427 26483
rect 1512 26460 1522 26520
rect 1578 26460 1792 26520
rect 1852 26460 1862 26520
rect 307 26380 353 26427
rect 307 26346 313 26380
rect 347 26346 353 26380
rect 307 26308 353 26346
rect 307 26274 313 26308
rect 347 26274 353 26308
rect 307 26236 353 26274
rect 307 26202 313 26236
rect 347 26202 353 26236
rect 307 26155 353 26202
rect 403 26380 449 26427
rect 403 26346 409 26380
rect 443 26346 449 26380
rect 403 26308 449 26346
rect 403 26274 409 26308
rect 443 26274 449 26308
rect 403 26236 449 26274
rect 403 26202 409 26236
rect 443 26202 449 26236
rect 403 26155 449 26202
rect 499 26380 545 26427
rect 499 26346 505 26380
rect 539 26346 545 26380
rect 499 26308 545 26346
rect 499 26274 505 26308
rect 539 26274 545 26308
rect 499 26236 545 26274
rect 499 26202 505 26236
rect 539 26202 545 26236
rect 499 26155 545 26202
rect 595 26380 641 26427
rect 595 26346 601 26380
rect 635 26346 641 26380
rect 595 26308 641 26346
rect 595 26274 601 26308
rect 635 26274 641 26308
rect 595 26236 641 26274
rect 595 26202 601 26236
rect 635 26202 641 26236
rect 595 26155 641 26202
rect 691 26380 737 26427
rect 691 26346 697 26380
rect 731 26346 737 26380
rect 691 26308 737 26346
rect 691 26274 697 26308
rect 731 26274 737 26308
rect 691 26236 737 26274
rect 691 26202 697 26236
rect 731 26202 737 26236
rect 691 26155 737 26202
rect 787 26380 833 26427
rect 787 26346 793 26380
rect 827 26346 833 26380
rect 787 26308 833 26346
rect 787 26274 793 26308
rect 827 26274 833 26308
rect 787 26236 833 26274
rect 787 26202 793 26236
rect 827 26202 833 26236
rect 787 26155 833 26202
rect 883 26380 929 26427
rect 883 26346 889 26380
rect 923 26346 929 26380
rect 883 26308 929 26346
rect 883 26274 889 26308
rect 923 26274 929 26308
rect 883 26236 929 26274
rect 883 26202 889 26236
rect 923 26202 929 26236
rect 883 26155 929 26202
rect 979 26380 1025 26427
rect 979 26346 985 26380
rect 1019 26346 1025 26380
rect 979 26308 1025 26346
rect 979 26274 985 26308
rect 1019 26274 1025 26308
rect 979 26236 1025 26274
rect 979 26202 985 26236
rect 1019 26202 1025 26236
rect 979 26155 1025 26202
rect 1075 26380 1121 26427
rect 1075 26346 1081 26380
rect 1115 26346 1121 26380
rect 1075 26308 1121 26346
rect 1075 26274 1081 26308
rect 1115 26274 1121 26308
rect 1075 26236 1121 26274
rect 1075 26202 1081 26236
rect 1115 26202 1121 26236
rect 1075 26155 1121 26202
rect 1171 26380 1217 26427
rect 1171 26346 1177 26380
rect 1211 26346 1217 26380
rect 1171 26308 1217 26346
rect 1171 26274 1177 26308
rect 1211 26274 1217 26308
rect 1171 26236 1217 26274
rect 1171 26202 1177 26236
rect 1211 26202 1217 26236
rect 1171 26155 1217 26202
rect 1267 26380 1313 26427
rect 1267 26346 1273 26380
rect 1307 26346 1313 26380
rect 1267 26308 1313 26346
rect 1267 26274 1273 26308
rect 1307 26274 1313 26308
rect 1267 26236 1313 26274
rect 1267 26202 1273 26236
rect 1307 26202 1313 26236
rect 1267 26155 1313 26202
rect 1381 26411 1427 26449
rect 1381 26377 1387 26411
rect 1421 26377 1427 26411
rect 1381 26339 1427 26377
rect 1381 26305 1387 26339
rect 1421 26305 1427 26339
rect 1381 26267 1427 26305
rect 1381 26233 1387 26267
rect 1421 26233 1427 26267
rect 1381 26223 1427 26233
rect 1381 26221 2160 26223
rect 1381 26195 2056 26221
rect 1381 26170 1387 26195
rect 1380 26161 1387 26170
rect 1421 26161 2056 26195
rect 0 25980 163 26014
rect 129 25603 163 25980
rect 313 26014 347 26155
rect 505 26014 539 26155
rect 697 26014 731 26155
rect 889 26014 923 26155
rect 1081 26014 1115 26155
rect 1273 26014 1307 26155
rect 1380 26113 2056 26161
rect 2190 26113 2200 26221
rect 1380 26111 2160 26113
rect 2282 26018 2316 26581
rect 2447 26471 2457 26523
rect 2509 26471 2519 26523
rect 2562 26431 2596 26581
rect 2640 26471 2650 26523
rect 2702 26471 2712 26523
rect 2754 26431 2788 26581
rect 2831 26471 2841 26523
rect 2893 26471 2903 26523
rect 2946 26431 2980 26581
rect 3023 26471 3033 26523
rect 3085 26471 3095 26523
rect 3138 26431 3172 26581
rect 3215 26471 3225 26523
rect 3277 26471 3287 26523
rect 3330 26431 3364 26581
rect 3407 26471 3417 26523
rect 3469 26471 3479 26523
rect 3534 26487 3580 26695
rect 3534 26453 3540 26487
rect 3574 26453 3580 26487
rect 2460 26384 2506 26431
rect 2460 26350 2466 26384
rect 2500 26350 2506 26384
rect 2460 26312 2506 26350
rect 2460 26278 2466 26312
rect 2500 26278 2506 26312
rect 2460 26240 2506 26278
rect 2460 26206 2466 26240
rect 2500 26206 2506 26240
rect 2460 26159 2506 26206
rect 2556 26384 2602 26431
rect 2556 26350 2562 26384
rect 2596 26350 2602 26384
rect 2556 26312 2602 26350
rect 2556 26278 2562 26312
rect 2596 26278 2602 26312
rect 2556 26240 2602 26278
rect 2556 26206 2562 26240
rect 2596 26206 2602 26240
rect 2556 26159 2602 26206
rect 2652 26384 2698 26431
rect 2652 26350 2658 26384
rect 2692 26350 2698 26384
rect 2652 26312 2698 26350
rect 2652 26278 2658 26312
rect 2692 26278 2698 26312
rect 2652 26240 2698 26278
rect 2652 26206 2658 26240
rect 2692 26206 2698 26240
rect 2652 26159 2698 26206
rect 2748 26384 2794 26431
rect 2748 26350 2754 26384
rect 2788 26350 2794 26384
rect 2748 26312 2794 26350
rect 2748 26278 2754 26312
rect 2788 26278 2794 26312
rect 2748 26240 2794 26278
rect 2748 26206 2754 26240
rect 2788 26206 2794 26240
rect 2748 26159 2794 26206
rect 2844 26384 2890 26431
rect 2844 26350 2850 26384
rect 2884 26350 2890 26384
rect 2844 26312 2890 26350
rect 2844 26278 2850 26312
rect 2884 26278 2890 26312
rect 2844 26240 2890 26278
rect 2844 26206 2850 26240
rect 2884 26206 2890 26240
rect 2844 26159 2890 26206
rect 2940 26384 2986 26431
rect 2940 26350 2946 26384
rect 2980 26350 2986 26384
rect 2940 26312 2986 26350
rect 2940 26278 2946 26312
rect 2980 26278 2986 26312
rect 2940 26240 2986 26278
rect 2940 26206 2946 26240
rect 2980 26206 2986 26240
rect 2940 26159 2986 26206
rect 3036 26384 3082 26431
rect 3036 26350 3042 26384
rect 3076 26350 3082 26384
rect 3036 26312 3082 26350
rect 3036 26278 3042 26312
rect 3076 26278 3082 26312
rect 3036 26240 3082 26278
rect 3036 26206 3042 26240
rect 3076 26206 3082 26240
rect 3036 26159 3082 26206
rect 3132 26384 3178 26431
rect 3132 26350 3138 26384
rect 3172 26350 3178 26384
rect 3132 26312 3178 26350
rect 3132 26278 3138 26312
rect 3172 26278 3178 26312
rect 3132 26240 3178 26278
rect 3132 26206 3138 26240
rect 3172 26206 3178 26240
rect 3132 26159 3178 26206
rect 3228 26384 3274 26431
rect 3228 26350 3234 26384
rect 3268 26350 3274 26384
rect 3228 26312 3274 26350
rect 3228 26278 3234 26312
rect 3268 26278 3274 26312
rect 3228 26240 3274 26278
rect 3228 26206 3234 26240
rect 3268 26206 3274 26240
rect 3228 26159 3274 26206
rect 3324 26384 3370 26431
rect 3324 26350 3330 26384
rect 3364 26350 3370 26384
rect 3324 26312 3370 26350
rect 3324 26278 3330 26312
rect 3364 26278 3370 26312
rect 3324 26240 3370 26278
rect 3324 26206 3330 26240
rect 3364 26206 3370 26240
rect 3324 26159 3370 26206
rect 3420 26384 3466 26431
rect 3420 26350 3426 26384
rect 3460 26350 3466 26384
rect 3420 26312 3466 26350
rect 3420 26278 3426 26312
rect 3460 26278 3466 26312
rect 3420 26240 3466 26278
rect 3420 26206 3426 26240
rect 3460 26206 3466 26240
rect 3420 26159 3466 26206
rect 3534 26415 3580 26453
rect 3534 26381 3540 26415
rect 3574 26381 3580 26415
rect 3534 26343 3580 26381
rect 3534 26309 3540 26343
rect 3574 26309 3580 26343
rect 3534 26271 3580 26309
rect 3534 26237 3540 26271
rect 3574 26237 3580 26271
rect 3534 26199 3580 26237
rect 3534 26165 3540 26199
rect 3574 26165 3580 26199
rect 2101 26014 2316 26018
rect 313 25984 2316 26014
rect 313 25980 2141 25984
rect 313 25847 347 25980
rect 505 25847 539 25980
rect 697 25847 731 25980
rect 889 25847 923 25980
rect 1081 25847 1115 25980
rect 1273 25847 1307 25980
rect 1381 25854 1608 25877
rect 307 25812 353 25847
rect 307 25778 313 25812
rect 347 25778 353 25812
rect 307 25743 353 25778
rect 403 25812 449 25847
rect 403 25778 409 25812
rect 443 25778 449 25812
rect 403 25743 449 25778
rect 499 25812 545 25847
rect 499 25778 505 25812
rect 539 25778 545 25812
rect 499 25743 545 25778
rect 595 25812 641 25847
rect 595 25778 601 25812
rect 635 25778 641 25812
rect 595 25743 641 25778
rect 691 25812 737 25847
rect 691 25778 697 25812
rect 731 25778 737 25812
rect 691 25743 737 25778
rect 787 25812 833 25847
rect 787 25778 793 25812
rect 827 25778 833 25812
rect 787 25743 833 25778
rect 883 25812 929 25847
rect 883 25778 889 25812
rect 923 25778 929 25812
rect 883 25743 929 25778
rect 979 25812 1025 25847
rect 979 25778 985 25812
rect 1019 25778 1025 25812
rect 979 25743 1025 25778
rect 1075 25812 1121 25847
rect 1075 25778 1081 25812
rect 1115 25778 1121 25812
rect 1075 25743 1121 25778
rect 1171 25812 1217 25847
rect 1171 25778 1177 25812
rect 1211 25778 1217 25812
rect 1171 25743 1217 25778
rect 1267 25812 1313 25847
rect 1267 25778 1273 25812
rect 1307 25778 1313 25812
rect 1267 25743 1313 25778
rect 1381 25820 1387 25854
rect 1421 25820 1608 25854
rect 1381 25782 1608 25820
rect 1381 25748 1387 25782
rect 1421 25757 1608 25782
rect 1421 25748 1427 25757
rect 1560 25755 1608 25757
rect 1598 25753 1608 25755
rect 1720 25753 1730 25877
rect 297 25712 363 25715
rect 294 25660 304 25712
rect 356 25660 366 25712
rect 297 25655 363 25660
rect 409 25603 443 25743
rect 489 25712 555 25715
rect 485 25660 495 25712
rect 547 25660 557 25712
rect 489 25655 555 25660
rect 601 25603 635 25743
rect 681 25712 747 25715
rect 677 25660 687 25712
rect 739 25660 749 25712
rect 681 25655 747 25660
rect 793 25603 827 25743
rect 873 25712 939 25715
rect 869 25660 879 25712
rect 931 25660 941 25712
rect 873 25655 939 25660
rect 985 25603 1019 25743
rect 1065 25711 1131 25715
rect 1062 25659 1072 25711
rect 1124 25659 1134 25711
rect 1065 25655 1131 25659
rect 1177 25603 1211 25743
rect 1257 25711 1323 25715
rect 1254 25659 1264 25711
rect 1316 25659 1326 25711
rect 1381 25710 1427 25748
rect 1920 25715 1930 25717
rect 1381 25676 1387 25710
rect 1421 25676 1427 25710
rect 1257 25655 1323 25659
rect 129 25569 1211 25603
rect 1381 25533 1427 25676
rect 1458 25659 1468 25715
rect 1524 25661 1930 25715
rect 1986 25661 1996 25717
rect 1524 25659 1986 25661
rect 2282 25607 2316 25984
rect 2466 26018 2500 26159
rect 2658 26018 2692 26159
rect 2850 26018 2884 26159
rect 3042 26018 3076 26159
rect 3234 26018 3268 26159
rect 3426 26018 3460 26159
rect 3534 26121 3580 26165
rect 3803 26581 4885 26615
rect 3803 26018 3837 26581
rect 3968 26471 3978 26523
rect 4030 26471 4040 26523
rect 4083 26431 4117 26581
rect 4161 26471 4171 26523
rect 4223 26471 4233 26523
rect 4275 26431 4309 26581
rect 4352 26471 4362 26523
rect 4414 26471 4424 26523
rect 4467 26431 4501 26581
rect 4544 26471 4554 26523
rect 4606 26471 4616 26523
rect 4659 26431 4693 26581
rect 4736 26471 4746 26523
rect 4798 26471 4808 26523
rect 4851 26431 4885 26581
rect 4928 26471 4938 26523
rect 4990 26471 5000 26523
rect 5055 26487 5101 26692
rect 5055 26453 5061 26487
rect 5095 26453 5101 26487
rect 3981 26384 4027 26431
rect 3981 26350 3987 26384
rect 4021 26350 4027 26384
rect 3981 26312 4027 26350
rect 3981 26278 3987 26312
rect 4021 26278 4027 26312
rect 3981 26240 4027 26278
rect 3981 26206 3987 26240
rect 4021 26206 4027 26240
rect 3981 26159 4027 26206
rect 4077 26384 4123 26431
rect 4077 26350 4083 26384
rect 4117 26350 4123 26384
rect 4077 26312 4123 26350
rect 4077 26278 4083 26312
rect 4117 26278 4123 26312
rect 4077 26240 4123 26278
rect 4077 26206 4083 26240
rect 4117 26206 4123 26240
rect 4077 26159 4123 26206
rect 4173 26384 4219 26431
rect 4173 26350 4179 26384
rect 4213 26350 4219 26384
rect 4173 26312 4219 26350
rect 4173 26278 4179 26312
rect 4213 26278 4219 26312
rect 4173 26240 4219 26278
rect 4173 26206 4179 26240
rect 4213 26206 4219 26240
rect 4173 26159 4219 26206
rect 4269 26384 4315 26431
rect 4269 26350 4275 26384
rect 4309 26350 4315 26384
rect 4269 26312 4315 26350
rect 4269 26278 4275 26312
rect 4309 26278 4315 26312
rect 4269 26240 4315 26278
rect 4269 26206 4275 26240
rect 4309 26206 4315 26240
rect 4269 26159 4315 26206
rect 4365 26384 4411 26431
rect 4365 26350 4371 26384
rect 4405 26350 4411 26384
rect 4365 26312 4411 26350
rect 4365 26278 4371 26312
rect 4405 26278 4411 26312
rect 4365 26240 4411 26278
rect 4365 26206 4371 26240
rect 4405 26206 4411 26240
rect 4365 26159 4411 26206
rect 4461 26384 4507 26431
rect 4461 26350 4467 26384
rect 4501 26350 4507 26384
rect 4461 26312 4507 26350
rect 4461 26278 4467 26312
rect 4501 26278 4507 26312
rect 4461 26240 4507 26278
rect 4461 26206 4467 26240
rect 4501 26206 4507 26240
rect 4461 26159 4507 26206
rect 4557 26384 4603 26431
rect 4557 26350 4563 26384
rect 4597 26350 4603 26384
rect 4557 26312 4603 26350
rect 4557 26278 4563 26312
rect 4597 26278 4603 26312
rect 4557 26240 4603 26278
rect 4557 26206 4563 26240
rect 4597 26206 4603 26240
rect 4557 26159 4603 26206
rect 4653 26384 4699 26431
rect 4653 26350 4659 26384
rect 4693 26350 4699 26384
rect 4653 26312 4699 26350
rect 4653 26278 4659 26312
rect 4693 26278 4699 26312
rect 4653 26240 4699 26278
rect 4653 26206 4659 26240
rect 4693 26206 4699 26240
rect 4653 26159 4699 26206
rect 4749 26384 4795 26431
rect 4749 26350 4755 26384
rect 4789 26350 4795 26384
rect 4749 26312 4795 26350
rect 4749 26278 4755 26312
rect 4789 26278 4795 26312
rect 4749 26240 4795 26278
rect 4749 26206 4755 26240
rect 4789 26206 4795 26240
rect 4749 26159 4795 26206
rect 4845 26384 4891 26431
rect 4845 26350 4851 26384
rect 4885 26350 4891 26384
rect 4845 26312 4891 26350
rect 4845 26278 4851 26312
rect 4885 26278 4891 26312
rect 4845 26240 4891 26278
rect 4845 26206 4851 26240
rect 4885 26206 4891 26240
rect 4845 26159 4891 26206
rect 4941 26384 4987 26431
rect 4941 26350 4947 26384
rect 4981 26350 4987 26384
rect 4941 26312 4987 26350
rect 4941 26278 4947 26312
rect 4981 26278 4987 26312
rect 4941 26240 4987 26278
rect 4941 26206 4947 26240
rect 4981 26206 4987 26240
rect 4941 26159 4987 26206
rect 5055 26415 5101 26453
rect 5055 26381 5061 26415
rect 5095 26381 5101 26415
rect 5055 26343 5101 26381
rect 5055 26309 5061 26343
rect 5095 26312 5101 26343
rect 5274 26312 5550 26313
rect 5095 26309 5550 26312
rect 5055 26282 5550 26309
rect 5055 26271 5303 26282
rect 5055 26237 5061 26271
rect 5095 26248 5303 26271
rect 5337 26248 5395 26282
rect 5429 26248 5487 26282
rect 5521 26248 5550 26282
rect 5095 26237 5550 26248
rect 5055 26217 5550 26237
rect 5055 26199 5101 26217
rect 5055 26165 5061 26199
rect 5095 26165 5101 26199
rect 2466 25984 3837 26018
rect 2466 25851 2500 25984
rect 2658 25851 2692 25984
rect 2850 25851 2884 25984
rect 3042 25851 3076 25984
rect 3234 25851 3268 25984
rect 3426 25851 3460 25984
rect 3671 25894 3681 25946
rect 3733 25894 3743 25946
rect 3679 25893 3691 25894
rect 3725 25893 3737 25894
rect 3679 25887 3737 25893
rect 3534 25858 3580 25881
rect 2460 25816 2506 25851
rect 2460 25782 2466 25816
rect 2500 25782 2506 25816
rect 2460 25747 2506 25782
rect 2556 25816 2602 25851
rect 2556 25782 2562 25816
rect 2596 25782 2602 25816
rect 2556 25747 2602 25782
rect 2652 25816 2698 25851
rect 2652 25782 2658 25816
rect 2692 25782 2698 25816
rect 2652 25747 2698 25782
rect 2748 25816 2794 25851
rect 2748 25782 2754 25816
rect 2788 25782 2794 25816
rect 2748 25747 2794 25782
rect 2844 25816 2890 25851
rect 2844 25782 2850 25816
rect 2884 25782 2890 25816
rect 2844 25747 2890 25782
rect 2940 25816 2986 25851
rect 2940 25782 2946 25816
rect 2980 25782 2986 25816
rect 2940 25747 2986 25782
rect 3036 25816 3082 25851
rect 3036 25782 3042 25816
rect 3076 25782 3082 25816
rect 3036 25747 3082 25782
rect 3132 25816 3178 25851
rect 3132 25782 3138 25816
rect 3172 25782 3178 25816
rect 3132 25747 3178 25782
rect 3228 25816 3274 25851
rect 3228 25782 3234 25816
rect 3268 25782 3274 25816
rect 3228 25747 3274 25782
rect 3324 25816 3370 25851
rect 3324 25782 3330 25816
rect 3364 25782 3370 25816
rect 3324 25747 3370 25782
rect 3420 25816 3466 25851
rect 3420 25782 3426 25816
rect 3460 25782 3466 25816
rect 3420 25747 3466 25782
rect 3534 25824 3540 25858
rect 3574 25856 3580 25858
rect 3803 25856 3837 25984
rect 3574 25855 3680 25856
rect 3734 25855 3837 25856
rect 3574 25843 3687 25855
rect 3574 25824 3647 25843
rect 3534 25786 3647 25824
rect 3534 25752 3540 25786
rect 3574 25767 3647 25786
rect 3681 25767 3687 25843
rect 3574 25756 3687 25767
rect 3574 25752 3580 25756
rect 3641 25755 3687 25756
rect 3729 25843 3837 25855
rect 3987 26018 4021 26159
rect 4179 26018 4213 26159
rect 4371 26018 4405 26159
rect 4563 26018 4597 26159
rect 4755 26018 4789 26159
rect 4947 26018 4981 26159
rect 5055 26121 5101 26165
rect 5683 26072 5743 27325
rect 5177 26038 5743 26072
rect 5177 26018 5211 26038
rect 3987 25984 5211 26018
rect 3987 25851 4021 25984
rect 4179 25851 4213 25984
rect 4371 25851 4405 25984
rect 4563 25851 4597 25984
rect 4755 25851 4789 25984
rect 4947 25851 4981 25984
rect 5438 25980 5512 25981
rect 5326 25978 5400 25979
rect 5326 25926 5337 25978
rect 5389 25926 5400 25978
rect 5438 25928 5449 25980
rect 5501 25928 5512 25980
rect 5438 25927 5512 25928
rect 5326 25925 5400 25926
rect 5055 25858 5101 25881
rect 3729 25767 3735 25843
rect 3769 25767 3837 25843
rect 3729 25756 3837 25767
rect 3729 25755 3775 25756
rect 2450 25716 2516 25719
rect 2447 25664 2457 25716
rect 2509 25664 2519 25716
rect 2450 25659 2516 25664
rect 2562 25607 2596 25747
rect 2642 25716 2708 25719
rect 2638 25664 2648 25716
rect 2700 25664 2710 25716
rect 2642 25659 2708 25664
rect 2754 25607 2788 25747
rect 2834 25716 2900 25719
rect 2830 25664 2840 25716
rect 2892 25664 2902 25716
rect 2834 25659 2900 25664
rect 2946 25607 2980 25747
rect 3026 25716 3092 25719
rect 3022 25664 3032 25716
rect 3084 25664 3094 25716
rect 3026 25659 3092 25664
rect 3138 25607 3172 25747
rect 3218 25715 3284 25719
rect 3215 25663 3225 25715
rect 3277 25663 3287 25715
rect 3218 25659 3284 25663
rect 3330 25607 3364 25747
rect 3410 25715 3476 25719
rect 3407 25663 3417 25715
rect 3469 25663 3479 25715
rect 3534 25714 3580 25752
rect 3534 25680 3540 25714
rect 3574 25680 3580 25714
rect 3410 25659 3476 25663
rect 2282 25573 3364 25607
rect 3534 25497 3580 25680
rect 3803 25607 3837 25756
rect 3981 25816 4027 25851
rect 3981 25782 3987 25816
rect 4021 25782 4027 25816
rect 3981 25747 4027 25782
rect 4077 25816 4123 25851
rect 4077 25782 4083 25816
rect 4117 25782 4123 25816
rect 4077 25747 4123 25782
rect 4173 25816 4219 25851
rect 4173 25782 4179 25816
rect 4213 25782 4219 25816
rect 4173 25747 4219 25782
rect 4269 25816 4315 25851
rect 4269 25782 4275 25816
rect 4309 25782 4315 25816
rect 4269 25747 4315 25782
rect 4365 25816 4411 25851
rect 4365 25782 4371 25816
rect 4405 25782 4411 25816
rect 4365 25747 4411 25782
rect 4461 25816 4507 25851
rect 4461 25782 4467 25816
rect 4501 25782 4507 25816
rect 4461 25747 4507 25782
rect 4557 25816 4603 25851
rect 4557 25782 4563 25816
rect 4597 25782 4603 25816
rect 4557 25747 4603 25782
rect 4653 25816 4699 25851
rect 4653 25782 4659 25816
rect 4693 25782 4699 25816
rect 4653 25747 4699 25782
rect 4749 25816 4795 25851
rect 4749 25782 4755 25816
rect 4789 25782 4795 25816
rect 4749 25747 4795 25782
rect 4845 25816 4891 25851
rect 4845 25782 4851 25816
rect 4885 25782 4891 25816
rect 4845 25747 4891 25782
rect 4941 25816 4987 25851
rect 4941 25782 4947 25816
rect 4981 25782 4987 25816
rect 4941 25747 4987 25782
rect 5055 25824 5061 25858
rect 5095 25824 5101 25858
rect 5055 25786 5101 25824
rect 5055 25752 5061 25786
rect 5095 25769 5101 25786
rect 5095 25752 5550 25769
rect 3971 25716 4037 25719
rect 3968 25664 3978 25716
rect 4030 25664 4040 25716
rect 3971 25659 4037 25664
rect 4083 25607 4117 25747
rect 4163 25716 4229 25719
rect 4159 25664 4169 25716
rect 4221 25664 4231 25716
rect 4163 25659 4229 25664
rect 4275 25607 4309 25747
rect 4355 25716 4421 25719
rect 4351 25664 4361 25716
rect 4413 25664 4423 25716
rect 4355 25659 4421 25664
rect 4467 25607 4501 25747
rect 4547 25716 4613 25719
rect 4543 25664 4553 25716
rect 4605 25664 4615 25716
rect 4547 25659 4613 25664
rect 4659 25607 4693 25747
rect 4739 25715 4805 25719
rect 4736 25663 4746 25715
rect 4798 25663 4808 25715
rect 4739 25659 4805 25663
rect 4851 25607 4885 25747
rect 5055 25738 5550 25752
rect 4931 25715 4997 25719
rect 4928 25663 4938 25715
rect 4990 25663 5000 25715
rect 5055 25714 5303 25738
rect 5055 25680 5061 25714
rect 5095 25704 5303 25714
rect 5337 25704 5395 25738
rect 5429 25704 5487 25738
rect 5521 25704 5550 25738
rect 5095 25680 5550 25704
rect 5055 25673 5550 25680
rect 4931 25659 4997 25663
rect 3803 25573 4885 25607
rect 5055 25498 5101 25673
rect 129 25290 1211 25324
rect 129 24727 163 25290
rect 294 25180 304 25232
rect 356 25180 366 25232
rect 409 25140 443 25290
rect 487 25180 497 25232
rect 549 25180 559 25232
rect 601 25140 635 25290
rect 678 25180 688 25232
rect 740 25180 750 25232
rect 793 25140 827 25290
rect 870 25180 880 25232
rect 932 25180 942 25232
rect 985 25140 1019 25290
rect 1062 25180 1072 25232
rect 1124 25180 1134 25232
rect 1177 25140 1211 25290
rect 1254 25180 1264 25232
rect 1316 25180 1326 25232
rect 1381 25196 1427 25360
rect 2282 25294 3364 25328
rect 1381 25162 1387 25196
rect 1421 25162 1427 25196
rect 1512 25173 1522 25233
rect 1578 25173 1792 25233
rect 1852 25173 1862 25233
rect 307 25093 353 25140
rect 307 25059 313 25093
rect 347 25059 353 25093
rect 307 25021 353 25059
rect 307 24987 313 25021
rect 347 24987 353 25021
rect 307 24949 353 24987
rect 307 24915 313 24949
rect 347 24915 353 24949
rect 307 24868 353 24915
rect 403 25093 449 25140
rect 403 25059 409 25093
rect 443 25059 449 25093
rect 403 25021 449 25059
rect 403 24987 409 25021
rect 443 24987 449 25021
rect 403 24949 449 24987
rect 403 24915 409 24949
rect 443 24915 449 24949
rect 403 24868 449 24915
rect 499 25093 545 25140
rect 499 25059 505 25093
rect 539 25059 545 25093
rect 499 25021 545 25059
rect 499 24987 505 25021
rect 539 24987 545 25021
rect 499 24949 545 24987
rect 499 24915 505 24949
rect 539 24915 545 24949
rect 499 24868 545 24915
rect 595 25093 641 25140
rect 595 25059 601 25093
rect 635 25059 641 25093
rect 595 25021 641 25059
rect 595 24987 601 25021
rect 635 24987 641 25021
rect 595 24949 641 24987
rect 595 24915 601 24949
rect 635 24915 641 24949
rect 595 24868 641 24915
rect 691 25093 737 25140
rect 691 25059 697 25093
rect 731 25059 737 25093
rect 691 25021 737 25059
rect 691 24987 697 25021
rect 731 24987 737 25021
rect 691 24949 737 24987
rect 691 24915 697 24949
rect 731 24915 737 24949
rect 691 24868 737 24915
rect 787 25093 833 25140
rect 787 25059 793 25093
rect 827 25059 833 25093
rect 787 25021 833 25059
rect 787 24987 793 25021
rect 827 24987 833 25021
rect 787 24949 833 24987
rect 787 24915 793 24949
rect 827 24915 833 24949
rect 787 24868 833 24915
rect 883 25093 929 25140
rect 883 25059 889 25093
rect 923 25059 929 25093
rect 883 25021 929 25059
rect 883 24987 889 25021
rect 923 24987 929 25021
rect 883 24949 929 24987
rect 883 24915 889 24949
rect 923 24915 929 24949
rect 883 24868 929 24915
rect 979 25093 1025 25140
rect 979 25059 985 25093
rect 1019 25059 1025 25093
rect 979 25021 1025 25059
rect 979 24987 985 25021
rect 1019 24987 1025 25021
rect 979 24949 1025 24987
rect 979 24915 985 24949
rect 1019 24915 1025 24949
rect 979 24868 1025 24915
rect 1075 25093 1121 25140
rect 1075 25059 1081 25093
rect 1115 25059 1121 25093
rect 1075 25021 1121 25059
rect 1075 24987 1081 25021
rect 1115 24987 1121 25021
rect 1075 24949 1121 24987
rect 1075 24915 1081 24949
rect 1115 24915 1121 24949
rect 1075 24868 1121 24915
rect 1171 25093 1217 25140
rect 1171 25059 1177 25093
rect 1211 25059 1217 25093
rect 1171 25021 1217 25059
rect 1171 24987 1177 25021
rect 1211 24987 1217 25021
rect 1171 24949 1217 24987
rect 1171 24915 1177 24949
rect 1211 24915 1217 24949
rect 1171 24868 1217 24915
rect 1267 25093 1313 25140
rect 1267 25059 1273 25093
rect 1307 25059 1313 25093
rect 1267 25021 1313 25059
rect 1267 24987 1273 25021
rect 1307 24987 1313 25021
rect 1267 24949 1313 24987
rect 1267 24915 1273 24949
rect 1307 24915 1313 24949
rect 1267 24868 1313 24915
rect 1381 25124 1427 25162
rect 1381 25090 1387 25124
rect 1421 25090 1427 25124
rect 1381 25052 1427 25090
rect 1381 25018 1387 25052
rect 1421 25018 1427 25052
rect 1381 24980 1427 25018
rect 1381 24946 1387 24980
rect 1421 24946 1427 24980
rect 1381 24936 1427 24946
rect 1381 24934 2160 24936
rect 1381 24908 2056 24934
rect 1381 24883 1387 24908
rect 1380 24874 1387 24883
rect 1421 24874 2056 24908
rect 0 24693 163 24727
rect 129 24316 163 24693
rect 313 24727 347 24868
rect 505 24727 539 24868
rect 697 24727 731 24868
rect 889 24727 923 24868
rect 1081 24727 1115 24868
rect 1273 24727 1307 24868
rect 1380 24826 2056 24874
rect 2190 24826 2200 24934
rect 1380 24824 2160 24826
rect 2282 24731 2316 25294
rect 2447 25184 2457 25236
rect 2509 25184 2519 25236
rect 2562 25144 2596 25294
rect 2640 25184 2650 25236
rect 2702 25184 2712 25236
rect 2754 25144 2788 25294
rect 2831 25184 2841 25236
rect 2893 25184 2903 25236
rect 2946 25144 2980 25294
rect 3023 25184 3033 25236
rect 3085 25184 3095 25236
rect 3138 25144 3172 25294
rect 3215 25184 3225 25236
rect 3277 25184 3287 25236
rect 3330 25144 3364 25294
rect 3407 25184 3417 25236
rect 3469 25184 3479 25236
rect 3534 25200 3580 25408
rect 3534 25166 3540 25200
rect 3574 25166 3580 25200
rect 2460 25097 2506 25144
rect 2460 25063 2466 25097
rect 2500 25063 2506 25097
rect 2460 25025 2506 25063
rect 2460 24991 2466 25025
rect 2500 24991 2506 25025
rect 2460 24953 2506 24991
rect 2460 24919 2466 24953
rect 2500 24919 2506 24953
rect 2460 24872 2506 24919
rect 2556 25097 2602 25144
rect 2556 25063 2562 25097
rect 2596 25063 2602 25097
rect 2556 25025 2602 25063
rect 2556 24991 2562 25025
rect 2596 24991 2602 25025
rect 2556 24953 2602 24991
rect 2556 24919 2562 24953
rect 2596 24919 2602 24953
rect 2556 24872 2602 24919
rect 2652 25097 2698 25144
rect 2652 25063 2658 25097
rect 2692 25063 2698 25097
rect 2652 25025 2698 25063
rect 2652 24991 2658 25025
rect 2692 24991 2698 25025
rect 2652 24953 2698 24991
rect 2652 24919 2658 24953
rect 2692 24919 2698 24953
rect 2652 24872 2698 24919
rect 2748 25097 2794 25144
rect 2748 25063 2754 25097
rect 2788 25063 2794 25097
rect 2748 25025 2794 25063
rect 2748 24991 2754 25025
rect 2788 24991 2794 25025
rect 2748 24953 2794 24991
rect 2748 24919 2754 24953
rect 2788 24919 2794 24953
rect 2748 24872 2794 24919
rect 2844 25097 2890 25144
rect 2844 25063 2850 25097
rect 2884 25063 2890 25097
rect 2844 25025 2890 25063
rect 2844 24991 2850 25025
rect 2884 24991 2890 25025
rect 2844 24953 2890 24991
rect 2844 24919 2850 24953
rect 2884 24919 2890 24953
rect 2844 24872 2890 24919
rect 2940 25097 2986 25144
rect 2940 25063 2946 25097
rect 2980 25063 2986 25097
rect 2940 25025 2986 25063
rect 2940 24991 2946 25025
rect 2980 24991 2986 25025
rect 2940 24953 2986 24991
rect 2940 24919 2946 24953
rect 2980 24919 2986 24953
rect 2940 24872 2986 24919
rect 3036 25097 3082 25144
rect 3036 25063 3042 25097
rect 3076 25063 3082 25097
rect 3036 25025 3082 25063
rect 3036 24991 3042 25025
rect 3076 24991 3082 25025
rect 3036 24953 3082 24991
rect 3036 24919 3042 24953
rect 3076 24919 3082 24953
rect 3036 24872 3082 24919
rect 3132 25097 3178 25144
rect 3132 25063 3138 25097
rect 3172 25063 3178 25097
rect 3132 25025 3178 25063
rect 3132 24991 3138 25025
rect 3172 24991 3178 25025
rect 3132 24953 3178 24991
rect 3132 24919 3138 24953
rect 3172 24919 3178 24953
rect 3132 24872 3178 24919
rect 3228 25097 3274 25144
rect 3228 25063 3234 25097
rect 3268 25063 3274 25097
rect 3228 25025 3274 25063
rect 3228 24991 3234 25025
rect 3268 24991 3274 25025
rect 3228 24953 3274 24991
rect 3228 24919 3234 24953
rect 3268 24919 3274 24953
rect 3228 24872 3274 24919
rect 3324 25097 3370 25144
rect 3324 25063 3330 25097
rect 3364 25063 3370 25097
rect 3324 25025 3370 25063
rect 3324 24991 3330 25025
rect 3364 24991 3370 25025
rect 3324 24953 3370 24991
rect 3324 24919 3330 24953
rect 3364 24919 3370 24953
rect 3324 24872 3370 24919
rect 3420 25097 3466 25144
rect 3420 25063 3426 25097
rect 3460 25063 3466 25097
rect 3420 25025 3466 25063
rect 3420 24991 3426 25025
rect 3460 24991 3466 25025
rect 3420 24953 3466 24991
rect 3420 24919 3426 24953
rect 3460 24919 3466 24953
rect 3420 24872 3466 24919
rect 3534 25128 3580 25166
rect 3534 25094 3540 25128
rect 3574 25094 3580 25128
rect 3534 25056 3580 25094
rect 3534 25022 3540 25056
rect 3574 25022 3580 25056
rect 3534 24984 3580 25022
rect 3534 24950 3540 24984
rect 3574 24950 3580 24984
rect 3534 24912 3580 24950
rect 3534 24878 3540 24912
rect 3574 24878 3580 24912
rect 2101 24727 2316 24731
rect 313 24697 2316 24727
rect 313 24693 2141 24697
rect 313 24560 347 24693
rect 505 24560 539 24693
rect 697 24560 731 24693
rect 889 24560 923 24693
rect 1081 24560 1115 24693
rect 1273 24560 1307 24693
rect 1381 24567 1608 24590
rect 307 24525 353 24560
rect 307 24491 313 24525
rect 347 24491 353 24525
rect 307 24456 353 24491
rect 403 24525 449 24560
rect 403 24491 409 24525
rect 443 24491 449 24525
rect 403 24456 449 24491
rect 499 24525 545 24560
rect 499 24491 505 24525
rect 539 24491 545 24525
rect 499 24456 545 24491
rect 595 24525 641 24560
rect 595 24491 601 24525
rect 635 24491 641 24525
rect 595 24456 641 24491
rect 691 24525 737 24560
rect 691 24491 697 24525
rect 731 24491 737 24525
rect 691 24456 737 24491
rect 787 24525 833 24560
rect 787 24491 793 24525
rect 827 24491 833 24525
rect 787 24456 833 24491
rect 883 24525 929 24560
rect 883 24491 889 24525
rect 923 24491 929 24525
rect 883 24456 929 24491
rect 979 24525 1025 24560
rect 979 24491 985 24525
rect 1019 24491 1025 24525
rect 979 24456 1025 24491
rect 1075 24525 1121 24560
rect 1075 24491 1081 24525
rect 1115 24491 1121 24525
rect 1075 24456 1121 24491
rect 1171 24525 1217 24560
rect 1171 24491 1177 24525
rect 1211 24491 1217 24525
rect 1171 24456 1217 24491
rect 1267 24525 1313 24560
rect 1267 24491 1273 24525
rect 1307 24491 1313 24525
rect 1267 24456 1313 24491
rect 1381 24533 1387 24567
rect 1421 24533 1608 24567
rect 1381 24495 1608 24533
rect 1381 24461 1387 24495
rect 1421 24470 1608 24495
rect 1421 24461 1427 24470
rect 1560 24468 1608 24470
rect 1598 24466 1608 24468
rect 1720 24466 1730 24590
rect 297 24425 363 24428
rect 294 24373 304 24425
rect 356 24373 366 24425
rect 297 24368 363 24373
rect 409 24316 443 24456
rect 489 24425 555 24428
rect 485 24373 495 24425
rect 547 24373 557 24425
rect 489 24368 555 24373
rect 601 24316 635 24456
rect 681 24425 747 24428
rect 677 24373 687 24425
rect 739 24373 749 24425
rect 681 24368 747 24373
rect 793 24316 827 24456
rect 873 24425 939 24428
rect 869 24373 879 24425
rect 931 24373 941 24425
rect 873 24368 939 24373
rect 985 24316 1019 24456
rect 1065 24424 1131 24428
rect 1062 24372 1072 24424
rect 1124 24372 1134 24424
rect 1065 24368 1131 24372
rect 1177 24316 1211 24456
rect 1257 24424 1323 24428
rect 1254 24372 1264 24424
rect 1316 24372 1326 24424
rect 1381 24423 1427 24461
rect 1920 24428 1930 24430
rect 1381 24389 1387 24423
rect 1421 24389 1427 24423
rect 1257 24368 1323 24372
rect 129 24282 1211 24316
rect 1381 24246 1427 24389
rect 1458 24372 1468 24428
rect 1524 24374 1930 24428
rect 1986 24374 1996 24430
rect 1524 24372 1986 24374
rect 2282 24320 2316 24697
rect 2466 24731 2500 24872
rect 2658 24731 2692 24872
rect 2850 24731 2884 24872
rect 3042 24731 3076 24872
rect 3234 24731 3268 24872
rect 3426 24731 3460 24872
rect 3534 24834 3580 24878
rect 3803 25294 4885 25328
rect 3803 24731 3837 25294
rect 3968 25184 3978 25236
rect 4030 25184 4040 25236
rect 4083 25144 4117 25294
rect 4161 25184 4171 25236
rect 4223 25184 4233 25236
rect 4275 25144 4309 25294
rect 4352 25184 4362 25236
rect 4414 25184 4424 25236
rect 4467 25144 4501 25294
rect 4544 25184 4554 25236
rect 4606 25184 4616 25236
rect 4659 25144 4693 25294
rect 4736 25184 4746 25236
rect 4798 25184 4808 25236
rect 4851 25144 4885 25294
rect 4928 25184 4938 25236
rect 4990 25184 5000 25236
rect 5055 25200 5101 25405
rect 5055 25166 5061 25200
rect 5095 25166 5101 25200
rect 3981 25097 4027 25144
rect 3981 25063 3987 25097
rect 4021 25063 4027 25097
rect 3981 25025 4027 25063
rect 3981 24991 3987 25025
rect 4021 24991 4027 25025
rect 3981 24953 4027 24991
rect 3981 24919 3987 24953
rect 4021 24919 4027 24953
rect 3981 24872 4027 24919
rect 4077 25097 4123 25144
rect 4077 25063 4083 25097
rect 4117 25063 4123 25097
rect 4077 25025 4123 25063
rect 4077 24991 4083 25025
rect 4117 24991 4123 25025
rect 4077 24953 4123 24991
rect 4077 24919 4083 24953
rect 4117 24919 4123 24953
rect 4077 24872 4123 24919
rect 4173 25097 4219 25144
rect 4173 25063 4179 25097
rect 4213 25063 4219 25097
rect 4173 25025 4219 25063
rect 4173 24991 4179 25025
rect 4213 24991 4219 25025
rect 4173 24953 4219 24991
rect 4173 24919 4179 24953
rect 4213 24919 4219 24953
rect 4173 24872 4219 24919
rect 4269 25097 4315 25144
rect 4269 25063 4275 25097
rect 4309 25063 4315 25097
rect 4269 25025 4315 25063
rect 4269 24991 4275 25025
rect 4309 24991 4315 25025
rect 4269 24953 4315 24991
rect 4269 24919 4275 24953
rect 4309 24919 4315 24953
rect 4269 24872 4315 24919
rect 4365 25097 4411 25144
rect 4365 25063 4371 25097
rect 4405 25063 4411 25097
rect 4365 25025 4411 25063
rect 4365 24991 4371 25025
rect 4405 24991 4411 25025
rect 4365 24953 4411 24991
rect 4365 24919 4371 24953
rect 4405 24919 4411 24953
rect 4365 24872 4411 24919
rect 4461 25097 4507 25144
rect 4461 25063 4467 25097
rect 4501 25063 4507 25097
rect 4461 25025 4507 25063
rect 4461 24991 4467 25025
rect 4501 24991 4507 25025
rect 4461 24953 4507 24991
rect 4461 24919 4467 24953
rect 4501 24919 4507 24953
rect 4461 24872 4507 24919
rect 4557 25097 4603 25144
rect 4557 25063 4563 25097
rect 4597 25063 4603 25097
rect 4557 25025 4603 25063
rect 4557 24991 4563 25025
rect 4597 24991 4603 25025
rect 4557 24953 4603 24991
rect 4557 24919 4563 24953
rect 4597 24919 4603 24953
rect 4557 24872 4603 24919
rect 4653 25097 4699 25144
rect 4653 25063 4659 25097
rect 4693 25063 4699 25097
rect 4653 25025 4699 25063
rect 4653 24991 4659 25025
rect 4693 24991 4699 25025
rect 4653 24953 4699 24991
rect 4653 24919 4659 24953
rect 4693 24919 4699 24953
rect 4653 24872 4699 24919
rect 4749 25097 4795 25144
rect 4749 25063 4755 25097
rect 4789 25063 4795 25097
rect 4749 25025 4795 25063
rect 4749 24991 4755 25025
rect 4789 24991 4795 25025
rect 4749 24953 4795 24991
rect 4749 24919 4755 24953
rect 4789 24919 4795 24953
rect 4749 24872 4795 24919
rect 4845 25097 4891 25144
rect 4845 25063 4851 25097
rect 4885 25063 4891 25097
rect 4845 25025 4891 25063
rect 4845 24991 4851 25025
rect 4885 24991 4891 25025
rect 4845 24953 4891 24991
rect 4845 24919 4851 24953
rect 4885 24919 4891 24953
rect 4845 24872 4891 24919
rect 4941 25097 4987 25144
rect 4941 25063 4947 25097
rect 4981 25063 4987 25097
rect 4941 25025 4987 25063
rect 4941 24991 4947 25025
rect 4981 24991 4987 25025
rect 4941 24953 4987 24991
rect 4941 24919 4947 24953
rect 4981 24919 4987 24953
rect 4941 24872 4987 24919
rect 5055 25128 5101 25166
rect 5055 25094 5061 25128
rect 5095 25094 5101 25128
rect 5055 25056 5101 25094
rect 5055 25022 5061 25056
rect 5095 25025 5101 25056
rect 5274 25025 5550 25026
rect 5095 25022 5550 25025
rect 5055 24995 5550 25022
rect 5055 24984 5303 24995
rect 5055 24950 5061 24984
rect 5095 24961 5303 24984
rect 5337 24961 5395 24995
rect 5429 24961 5487 24995
rect 5521 24961 5550 24995
rect 5095 24950 5550 24961
rect 5055 24930 5550 24950
rect 5055 24912 5101 24930
rect 5055 24878 5061 24912
rect 5095 24878 5101 24912
rect 2466 24697 3837 24731
rect 2466 24564 2500 24697
rect 2658 24564 2692 24697
rect 2850 24564 2884 24697
rect 3042 24564 3076 24697
rect 3234 24564 3268 24697
rect 3426 24564 3460 24697
rect 3671 24607 3681 24659
rect 3733 24607 3743 24659
rect 3679 24606 3691 24607
rect 3725 24606 3737 24607
rect 3679 24600 3737 24606
rect 3534 24571 3580 24594
rect 2460 24529 2506 24564
rect 2460 24495 2466 24529
rect 2500 24495 2506 24529
rect 2460 24460 2506 24495
rect 2556 24529 2602 24564
rect 2556 24495 2562 24529
rect 2596 24495 2602 24529
rect 2556 24460 2602 24495
rect 2652 24529 2698 24564
rect 2652 24495 2658 24529
rect 2692 24495 2698 24529
rect 2652 24460 2698 24495
rect 2748 24529 2794 24564
rect 2748 24495 2754 24529
rect 2788 24495 2794 24529
rect 2748 24460 2794 24495
rect 2844 24529 2890 24564
rect 2844 24495 2850 24529
rect 2884 24495 2890 24529
rect 2844 24460 2890 24495
rect 2940 24529 2986 24564
rect 2940 24495 2946 24529
rect 2980 24495 2986 24529
rect 2940 24460 2986 24495
rect 3036 24529 3082 24564
rect 3036 24495 3042 24529
rect 3076 24495 3082 24529
rect 3036 24460 3082 24495
rect 3132 24529 3178 24564
rect 3132 24495 3138 24529
rect 3172 24495 3178 24529
rect 3132 24460 3178 24495
rect 3228 24529 3274 24564
rect 3228 24495 3234 24529
rect 3268 24495 3274 24529
rect 3228 24460 3274 24495
rect 3324 24529 3370 24564
rect 3324 24495 3330 24529
rect 3364 24495 3370 24529
rect 3324 24460 3370 24495
rect 3420 24529 3466 24564
rect 3420 24495 3426 24529
rect 3460 24495 3466 24529
rect 3420 24460 3466 24495
rect 3534 24537 3540 24571
rect 3574 24569 3580 24571
rect 3803 24569 3837 24697
rect 3574 24568 3680 24569
rect 3734 24568 3837 24569
rect 3574 24556 3687 24568
rect 3574 24537 3647 24556
rect 3534 24499 3647 24537
rect 3534 24465 3540 24499
rect 3574 24480 3647 24499
rect 3681 24480 3687 24556
rect 3574 24469 3687 24480
rect 3574 24465 3580 24469
rect 3641 24468 3687 24469
rect 3729 24556 3837 24568
rect 3987 24731 4021 24872
rect 4179 24731 4213 24872
rect 4371 24731 4405 24872
rect 4563 24731 4597 24872
rect 4755 24731 4789 24872
rect 4947 24731 4981 24872
rect 5055 24834 5101 24878
rect 5683 24785 5743 26038
rect 5177 24751 5743 24785
rect 5177 24731 5211 24751
rect 3987 24697 5211 24731
rect 3987 24564 4021 24697
rect 4179 24564 4213 24697
rect 4371 24564 4405 24697
rect 4563 24564 4597 24697
rect 4755 24564 4789 24697
rect 4947 24564 4981 24697
rect 5438 24693 5512 24694
rect 5326 24691 5400 24692
rect 5326 24639 5337 24691
rect 5389 24639 5400 24691
rect 5438 24641 5449 24693
rect 5501 24641 5512 24693
rect 5438 24640 5512 24641
rect 5326 24638 5400 24639
rect 5055 24571 5101 24594
rect 3729 24480 3735 24556
rect 3769 24480 3837 24556
rect 3729 24469 3837 24480
rect 3729 24468 3775 24469
rect 2450 24429 2516 24432
rect 2447 24377 2457 24429
rect 2509 24377 2519 24429
rect 2450 24372 2516 24377
rect 2562 24320 2596 24460
rect 2642 24429 2708 24432
rect 2638 24377 2648 24429
rect 2700 24377 2710 24429
rect 2642 24372 2708 24377
rect 2754 24320 2788 24460
rect 2834 24429 2900 24432
rect 2830 24377 2840 24429
rect 2892 24377 2902 24429
rect 2834 24372 2900 24377
rect 2946 24320 2980 24460
rect 3026 24429 3092 24432
rect 3022 24377 3032 24429
rect 3084 24377 3094 24429
rect 3026 24372 3092 24377
rect 3138 24320 3172 24460
rect 3218 24428 3284 24432
rect 3215 24376 3225 24428
rect 3277 24376 3287 24428
rect 3218 24372 3284 24376
rect 3330 24320 3364 24460
rect 3410 24428 3476 24432
rect 3407 24376 3417 24428
rect 3469 24376 3479 24428
rect 3534 24427 3580 24465
rect 3534 24393 3540 24427
rect 3574 24393 3580 24427
rect 3410 24372 3476 24376
rect 2282 24286 3364 24320
rect 3534 24210 3580 24393
rect 3803 24320 3837 24469
rect 3981 24529 4027 24564
rect 3981 24495 3987 24529
rect 4021 24495 4027 24529
rect 3981 24460 4027 24495
rect 4077 24529 4123 24564
rect 4077 24495 4083 24529
rect 4117 24495 4123 24529
rect 4077 24460 4123 24495
rect 4173 24529 4219 24564
rect 4173 24495 4179 24529
rect 4213 24495 4219 24529
rect 4173 24460 4219 24495
rect 4269 24529 4315 24564
rect 4269 24495 4275 24529
rect 4309 24495 4315 24529
rect 4269 24460 4315 24495
rect 4365 24529 4411 24564
rect 4365 24495 4371 24529
rect 4405 24495 4411 24529
rect 4365 24460 4411 24495
rect 4461 24529 4507 24564
rect 4461 24495 4467 24529
rect 4501 24495 4507 24529
rect 4461 24460 4507 24495
rect 4557 24529 4603 24564
rect 4557 24495 4563 24529
rect 4597 24495 4603 24529
rect 4557 24460 4603 24495
rect 4653 24529 4699 24564
rect 4653 24495 4659 24529
rect 4693 24495 4699 24529
rect 4653 24460 4699 24495
rect 4749 24529 4795 24564
rect 4749 24495 4755 24529
rect 4789 24495 4795 24529
rect 4749 24460 4795 24495
rect 4845 24529 4891 24564
rect 4845 24495 4851 24529
rect 4885 24495 4891 24529
rect 4845 24460 4891 24495
rect 4941 24529 4987 24564
rect 4941 24495 4947 24529
rect 4981 24495 4987 24529
rect 4941 24460 4987 24495
rect 5055 24537 5061 24571
rect 5095 24537 5101 24571
rect 5055 24499 5101 24537
rect 5055 24465 5061 24499
rect 5095 24482 5101 24499
rect 5095 24465 5550 24482
rect 3971 24429 4037 24432
rect 3968 24377 3978 24429
rect 4030 24377 4040 24429
rect 3971 24372 4037 24377
rect 4083 24320 4117 24460
rect 4163 24429 4229 24432
rect 4159 24377 4169 24429
rect 4221 24377 4231 24429
rect 4163 24372 4229 24377
rect 4275 24320 4309 24460
rect 4355 24429 4421 24432
rect 4351 24377 4361 24429
rect 4413 24377 4423 24429
rect 4355 24372 4421 24377
rect 4467 24320 4501 24460
rect 4547 24429 4613 24432
rect 4543 24377 4553 24429
rect 4605 24377 4615 24429
rect 4547 24372 4613 24377
rect 4659 24320 4693 24460
rect 4739 24428 4805 24432
rect 4736 24376 4746 24428
rect 4798 24376 4808 24428
rect 4739 24372 4805 24376
rect 4851 24320 4885 24460
rect 5055 24451 5550 24465
rect 4931 24428 4997 24432
rect 4928 24376 4938 24428
rect 4990 24376 5000 24428
rect 5055 24427 5303 24451
rect 5055 24393 5061 24427
rect 5095 24417 5303 24427
rect 5337 24417 5395 24451
rect 5429 24417 5487 24451
rect 5521 24417 5550 24451
rect 5095 24393 5550 24417
rect 5055 24386 5550 24393
rect 4931 24372 4997 24376
rect 3803 24286 4885 24320
rect 5055 24211 5101 24386
rect 129 24003 1211 24037
rect 129 23440 163 24003
rect 294 23893 304 23945
rect 356 23893 366 23945
rect 409 23853 443 24003
rect 487 23893 497 23945
rect 549 23893 559 23945
rect 601 23853 635 24003
rect 678 23893 688 23945
rect 740 23893 750 23945
rect 793 23853 827 24003
rect 870 23893 880 23945
rect 932 23893 942 23945
rect 985 23853 1019 24003
rect 1062 23893 1072 23945
rect 1124 23893 1134 23945
rect 1177 23853 1211 24003
rect 1254 23893 1264 23945
rect 1316 23893 1326 23945
rect 1381 23909 1427 24073
rect 2282 24007 3364 24041
rect 1381 23875 1387 23909
rect 1421 23875 1427 23909
rect 1512 23886 1522 23946
rect 1578 23886 1792 23946
rect 1852 23886 1862 23946
rect 307 23806 353 23853
rect 307 23772 313 23806
rect 347 23772 353 23806
rect 307 23734 353 23772
rect 307 23700 313 23734
rect 347 23700 353 23734
rect 307 23662 353 23700
rect 307 23628 313 23662
rect 347 23628 353 23662
rect 307 23581 353 23628
rect 403 23806 449 23853
rect 403 23772 409 23806
rect 443 23772 449 23806
rect 403 23734 449 23772
rect 403 23700 409 23734
rect 443 23700 449 23734
rect 403 23662 449 23700
rect 403 23628 409 23662
rect 443 23628 449 23662
rect 403 23581 449 23628
rect 499 23806 545 23853
rect 499 23772 505 23806
rect 539 23772 545 23806
rect 499 23734 545 23772
rect 499 23700 505 23734
rect 539 23700 545 23734
rect 499 23662 545 23700
rect 499 23628 505 23662
rect 539 23628 545 23662
rect 499 23581 545 23628
rect 595 23806 641 23853
rect 595 23772 601 23806
rect 635 23772 641 23806
rect 595 23734 641 23772
rect 595 23700 601 23734
rect 635 23700 641 23734
rect 595 23662 641 23700
rect 595 23628 601 23662
rect 635 23628 641 23662
rect 595 23581 641 23628
rect 691 23806 737 23853
rect 691 23772 697 23806
rect 731 23772 737 23806
rect 691 23734 737 23772
rect 691 23700 697 23734
rect 731 23700 737 23734
rect 691 23662 737 23700
rect 691 23628 697 23662
rect 731 23628 737 23662
rect 691 23581 737 23628
rect 787 23806 833 23853
rect 787 23772 793 23806
rect 827 23772 833 23806
rect 787 23734 833 23772
rect 787 23700 793 23734
rect 827 23700 833 23734
rect 787 23662 833 23700
rect 787 23628 793 23662
rect 827 23628 833 23662
rect 787 23581 833 23628
rect 883 23806 929 23853
rect 883 23772 889 23806
rect 923 23772 929 23806
rect 883 23734 929 23772
rect 883 23700 889 23734
rect 923 23700 929 23734
rect 883 23662 929 23700
rect 883 23628 889 23662
rect 923 23628 929 23662
rect 883 23581 929 23628
rect 979 23806 1025 23853
rect 979 23772 985 23806
rect 1019 23772 1025 23806
rect 979 23734 1025 23772
rect 979 23700 985 23734
rect 1019 23700 1025 23734
rect 979 23662 1025 23700
rect 979 23628 985 23662
rect 1019 23628 1025 23662
rect 979 23581 1025 23628
rect 1075 23806 1121 23853
rect 1075 23772 1081 23806
rect 1115 23772 1121 23806
rect 1075 23734 1121 23772
rect 1075 23700 1081 23734
rect 1115 23700 1121 23734
rect 1075 23662 1121 23700
rect 1075 23628 1081 23662
rect 1115 23628 1121 23662
rect 1075 23581 1121 23628
rect 1171 23806 1217 23853
rect 1171 23772 1177 23806
rect 1211 23772 1217 23806
rect 1171 23734 1217 23772
rect 1171 23700 1177 23734
rect 1211 23700 1217 23734
rect 1171 23662 1217 23700
rect 1171 23628 1177 23662
rect 1211 23628 1217 23662
rect 1171 23581 1217 23628
rect 1267 23806 1313 23853
rect 1267 23772 1273 23806
rect 1307 23772 1313 23806
rect 1267 23734 1313 23772
rect 1267 23700 1273 23734
rect 1307 23700 1313 23734
rect 1267 23662 1313 23700
rect 1267 23628 1273 23662
rect 1307 23628 1313 23662
rect 1267 23581 1313 23628
rect 1381 23837 1427 23875
rect 1381 23803 1387 23837
rect 1421 23803 1427 23837
rect 1381 23765 1427 23803
rect 1381 23731 1387 23765
rect 1421 23731 1427 23765
rect 1381 23693 1427 23731
rect 1381 23659 1387 23693
rect 1421 23659 1427 23693
rect 1381 23649 1427 23659
rect 1381 23647 2160 23649
rect 1381 23621 2056 23647
rect 1381 23596 1387 23621
rect 1380 23587 1387 23596
rect 1421 23587 2056 23621
rect 0 23406 163 23440
rect 129 23029 163 23406
rect 313 23440 347 23581
rect 505 23440 539 23581
rect 697 23440 731 23581
rect 889 23440 923 23581
rect 1081 23440 1115 23581
rect 1273 23440 1307 23581
rect 1380 23539 2056 23587
rect 2190 23539 2200 23647
rect 1380 23537 2160 23539
rect 2282 23444 2316 24007
rect 2447 23897 2457 23949
rect 2509 23897 2519 23949
rect 2562 23857 2596 24007
rect 2640 23897 2650 23949
rect 2702 23897 2712 23949
rect 2754 23857 2788 24007
rect 2831 23897 2841 23949
rect 2893 23897 2903 23949
rect 2946 23857 2980 24007
rect 3023 23897 3033 23949
rect 3085 23897 3095 23949
rect 3138 23857 3172 24007
rect 3215 23897 3225 23949
rect 3277 23897 3287 23949
rect 3330 23857 3364 24007
rect 3407 23897 3417 23949
rect 3469 23897 3479 23949
rect 3534 23913 3580 24121
rect 3534 23879 3540 23913
rect 3574 23879 3580 23913
rect 2460 23810 2506 23857
rect 2460 23776 2466 23810
rect 2500 23776 2506 23810
rect 2460 23738 2506 23776
rect 2460 23704 2466 23738
rect 2500 23704 2506 23738
rect 2460 23666 2506 23704
rect 2460 23632 2466 23666
rect 2500 23632 2506 23666
rect 2460 23585 2506 23632
rect 2556 23810 2602 23857
rect 2556 23776 2562 23810
rect 2596 23776 2602 23810
rect 2556 23738 2602 23776
rect 2556 23704 2562 23738
rect 2596 23704 2602 23738
rect 2556 23666 2602 23704
rect 2556 23632 2562 23666
rect 2596 23632 2602 23666
rect 2556 23585 2602 23632
rect 2652 23810 2698 23857
rect 2652 23776 2658 23810
rect 2692 23776 2698 23810
rect 2652 23738 2698 23776
rect 2652 23704 2658 23738
rect 2692 23704 2698 23738
rect 2652 23666 2698 23704
rect 2652 23632 2658 23666
rect 2692 23632 2698 23666
rect 2652 23585 2698 23632
rect 2748 23810 2794 23857
rect 2748 23776 2754 23810
rect 2788 23776 2794 23810
rect 2748 23738 2794 23776
rect 2748 23704 2754 23738
rect 2788 23704 2794 23738
rect 2748 23666 2794 23704
rect 2748 23632 2754 23666
rect 2788 23632 2794 23666
rect 2748 23585 2794 23632
rect 2844 23810 2890 23857
rect 2844 23776 2850 23810
rect 2884 23776 2890 23810
rect 2844 23738 2890 23776
rect 2844 23704 2850 23738
rect 2884 23704 2890 23738
rect 2844 23666 2890 23704
rect 2844 23632 2850 23666
rect 2884 23632 2890 23666
rect 2844 23585 2890 23632
rect 2940 23810 2986 23857
rect 2940 23776 2946 23810
rect 2980 23776 2986 23810
rect 2940 23738 2986 23776
rect 2940 23704 2946 23738
rect 2980 23704 2986 23738
rect 2940 23666 2986 23704
rect 2940 23632 2946 23666
rect 2980 23632 2986 23666
rect 2940 23585 2986 23632
rect 3036 23810 3082 23857
rect 3036 23776 3042 23810
rect 3076 23776 3082 23810
rect 3036 23738 3082 23776
rect 3036 23704 3042 23738
rect 3076 23704 3082 23738
rect 3036 23666 3082 23704
rect 3036 23632 3042 23666
rect 3076 23632 3082 23666
rect 3036 23585 3082 23632
rect 3132 23810 3178 23857
rect 3132 23776 3138 23810
rect 3172 23776 3178 23810
rect 3132 23738 3178 23776
rect 3132 23704 3138 23738
rect 3172 23704 3178 23738
rect 3132 23666 3178 23704
rect 3132 23632 3138 23666
rect 3172 23632 3178 23666
rect 3132 23585 3178 23632
rect 3228 23810 3274 23857
rect 3228 23776 3234 23810
rect 3268 23776 3274 23810
rect 3228 23738 3274 23776
rect 3228 23704 3234 23738
rect 3268 23704 3274 23738
rect 3228 23666 3274 23704
rect 3228 23632 3234 23666
rect 3268 23632 3274 23666
rect 3228 23585 3274 23632
rect 3324 23810 3370 23857
rect 3324 23776 3330 23810
rect 3364 23776 3370 23810
rect 3324 23738 3370 23776
rect 3324 23704 3330 23738
rect 3364 23704 3370 23738
rect 3324 23666 3370 23704
rect 3324 23632 3330 23666
rect 3364 23632 3370 23666
rect 3324 23585 3370 23632
rect 3420 23810 3466 23857
rect 3420 23776 3426 23810
rect 3460 23776 3466 23810
rect 3420 23738 3466 23776
rect 3420 23704 3426 23738
rect 3460 23704 3466 23738
rect 3420 23666 3466 23704
rect 3420 23632 3426 23666
rect 3460 23632 3466 23666
rect 3420 23585 3466 23632
rect 3534 23841 3580 23879
rect 3534 23807 3540 23841
rect 3574 23807 3580 23841
rect 3534 23769 3580 23807
rect 3534 23735 3540 23769
rect 3574 23735 3580 23769
rect 3534 23697 3580 23735
rect 3534 23663 3540 23697
rect 3574 23663 3580 23697
rect 3534 23625 3580 23663
rect 3534 23591 3540 23625
rect 3574 23591 3580 23625
rect 2101 23440 2316 23444
rect 313 23410 2316 23440
rect 313 23406 2141 23410
rect 313 23273 347 23406
rect 505 23273 539 23406
rect 697 23273 731 23406
rect 889 23273 923 23406
rect 1081 23273 1115 23406
rect 1273 23273 1307 23406
rect 1381 23280 1608 23303
rect 307 23238 353 23273
rect 307 23204 313 23238
rect 347 23204 353 23238
rect 307 23169 353 23204
rect 403 23238 449 23273
rect 403 23204 409 23238
rect 443 23204 449 23238
rect 403 23169 449 23204
rect 499 23238 545 23273
rect 499 23204 505 23238
rect 539 23204 545 23238
rect 499 23169 545 23204
rect 595 23238 641 23273
rect 595 23204 601 23238
rect 635 23204 641 23238
rect 595 23169 641 23204
rect 691 23238 737 23273
rect 691 23204 697 23238
rect 731 23204 737 23238
rect 691 23169 737 23204
rect 787 23238 833 23273
rect 787 23204 793 23238
rect 827 23204 833 23238
rect 787 23169 833 23204
rect 883 23238 929 23273
rect 883 23204 889 23238
rect 923 23204 929 23238
rect 883 23169 929 23204
rect 979 23238 1025 23273
rect 979 23204 985 23238
rect 1019 23204 1025 23238
rect 979 23169 1025 23204
rect 1075 23238 1121 23273
rect 1075 23204 1081 23238
rect 1115 23204 1121 23238
rect 1075 23169 1121 23204
rect 1171 23238 1217 23273
rect 1171 23204 1177 23238
rect 1211 23204 1217 23238
rect 1171 23169 1217 23204
rect 1267 23238 1313 23273
rect 1267 23204 1273 23238
rect 1307 23204 1313 23238
rect 1267 23169 1313 23204
rect 1381 23246 1387 23280
rect 1421 23246 1608 23280
rect 1381 23208 1608 23246
rect 1381 23174 1387 23208
rect 1421 23183 1608 23208
rect 1421 23174 1427 23183
rect 1560 23181 1608 23183
rect 1598 23179 1608 23181
rect 1720 23179 1730 23303
rect 297 23138 363 23141
rect 294 23086 304 23138
rect 356 23086 366 23138
rect 297 23081 363 23086
rect 409 23029 443 23169
rect 489 23138 555 23141
rect 485 23086 495 23138
rect 547 23086 557 23138
rect 489 23081 555 23086
rect 601 23029 635 23169
rect 681 23138 747 23141
rect 677 23086 687 23138
rect 739 23086 749 23138
rect 681 23081 747 23086
rect 793 23029 827 23169
rect 873 23138 939 23141
rect 869 23086 879 23138
rect 931 23086 941 23138
rect 873 23081 939 23086
rect 985 23029 1019 23169
rect 1065 23137 1131 23141
rect 1062 23085 1072 23137
rect 1124 23085 1134 23137
rect 1065 23081 1131 23085
rect 1177 23029 1211 23169
rect 1257 23137 1323 23141
rect 1254 23085 1264 23137
rect 1316 23085 1326 23137
rect 1381 23136 1427 23174
rect 1920 23141 1930 23143
rect 1381 23102 1387 23136
rect 1421 23102 1427 23136
rect 1257 23081 1323 23085
rect 129 22995 1211 23029
rect 1381 22959 1427 23102
rect 1458 23085 1468 23141
rect 1524 23087 1930 23141
rect 1986 23087 1996 23143
rect 1524 23085 1986 23087
rect 2282 23033 2316 23410
rect 2466 23444 2500 23585
rect 2658 23444 2692 23585
rect 2850 23444 2884 23585
rect 3042 23444 3076 23585
rect 3234 23444 3268 23585
rect 3426 23444 3460 23585
rect 3534 23547 3580 23591
rect 3803 24007 4885 24041
rect 3803 23444 3837 24007
rect 3968 23897 3978 23949
rect 4030 23897 4040 23949
rect 4083 23857 4117 24007
rect 4161 23897 4171 23949
rect 4223 23897 4233 23949
rect 4275 23857 4309 24007
rect 4352 23897 4362 23949
rect 4414 23897 4424 23949
rect 4467 23857 4501 24007
rect 4544 23897 4554 23949
rect 4606 23897 4616 23949
rect 4659 23857 4693 24007
rect 4736 23897 4746 23949
rect 4798 23897 4808 23949
rect 4851 23857 4885 24007
rect 4928 23897 4938 23949
rect 4990 23897 5000 23949
rect 5055 23913 5101 24118
rect 5055 23879 5061 23913
rect 5095 23879 5101 23913
rect 3981 23810 4027 23857
rect 3981 23776 3987 23810
rect 4021 23776 4027 23810
rect 3981 23738 4027 23776
rect 3981 23704 3987 23738
rect 4021 23704 4027 23738
rect 3981 23666 4027 23704
rect 3981 23632 3987 23666
rect 4021 23632 4027 23666
rect 3981 23585 4027 23632
rect 4077 23810 4123 23857
rect 4077 23776 4083 23810
rect 4117 23776 4123 23810
rect 4077 23738 4123 23776
rect 4077 23704 4083 23738
rect 4117 23704 4123 23738
rect 4077 23666 4123 23704
rect 4077 23632 4083 23666
rect 4117 23632 4123 23666
rect 4077 23585 4123 23632
rect 4173 23810 4219 23857
rect 4173 23776 4179 23810
rect 4213 23776 4219 23810
rect 4173 23738 4219 23776
rect 4173 23704 4179 23738
rect 4213 23704 4219 23738
rect 4173 23666 4219 23704
rect 4173 23632 4179 23666
rect 4213 23632 4219 23666
rect 4173 23585 4219 23632
rect 4269 23810 4315 23857
rect 4269 23776 4275 23810
rect 4309 23776 4315 23810
rect 4269 23738 4315 23776
rect 4269 23704 4275 23738
rect 4309 23704 4315 23738
rect 4269 23666 4315 23704
rect 4269 23632 4275 23666
rect 4309 23632 4315 23666
rect 4269 23585 4315 23632
rect 4365 23810 4411 23857
rect 4365 23776 4371 23810
rect 4405 23776 4411 23810
rect 4365 23738 4411 23776
rect 4365 23704 4371 23738
rect 4405 23704 4411 23738
rect 4365 23666 4411 23704
rect 4365 23632 4371 23666
rect 4405 23632 4411 23666
rect 4365 23585 4411 23632
rect 4461 23810 4507 23857
rect 4461 23776 4467 23810
rect 4501 23776 4507 23810
rect 4461 23738 4507 23776
rect 4461 23704 4467 23738
rect 4501 23704 4507 23738
rect 4461 23666 4507 23704
rect 4461 23632 4467 23666
rect 4501 23632 4507 23666
rect 4461 23585 4507 23632
rect 4557 23810 4603 23857
rect 4557 23776 4563 23810
rect 4597 23776 4603 23810
rect 4557 23738 4603 23776
rect 4557 23704 4563 23738
rect 4597 23704 4603 23738
rect 4557 23666 4603 23704
rect 4557 23632 4563 23666
rect 4597 23632 4603 23666
rect 4557 23585 4603 23632
rect 4653 23810 4699 23857
rect 4653 23776 4659 23810
rect 4693 23776 4699 23810
rect 4653 23738 4699 23776
rect 4653 23704 4659 23738
rect 4693 23704 4699 23738
rect 4653 23666 4699 23704
rect 4653 23632 4659 23666
rect 4693 23632 4699 23666
rect 4653 23585 4699 23632
rect 4749 23810 4795 23857
rect 4749 23776 4755 23810
rect 4789 23776 4795 23810
rect 4749 23738 4795 23776
rect 4749 23704 4755 23738
rect 4789 23704 4795 23738
rect 4749 23666 4795 23704
rect 4749 23632 4755 23666
rect 4789 23632 4795 23666
rect 4749 23585 4795 23632
rect 4845 23810 4891 23857
rect 4845 23776 4851 23810
rect 4885 23776 4891 23810
rect 4845 23738 4891 23776
rect 4845 23704 4851 23738
rect 4885 23704 4891 23738
rect 4845 23666 4891 23704
rect 4845 23632 4851 23666
rect 4885 23632 4891 23666
rect 4845 23585 4891 23632
rect 4941 23810 4987 23857
rect 4941 23776 4947 23810
rect 4981 23776 4987 23810
rect 4941 23738 4987 23776
rect 4941 23704 4947 23738
rect 4981 23704 4987 23738
rect 4941 23666 4987 23704
rect 4941 23632 4947 23666
rect 4981 23632 4987 23666
rect 4941 23585 4987 23632
rect 5055 23841 5101 23879
rect 5055 23807 5061 23841
rect 5095 23807 5101 23841
rect 5055 23769 5101 23807
rect 5055 23735 5061 23769
rect 5095 23738 5101 23769
rect 5274 23738 5550 23739
rect 5095 23735 5550 23738
rect 5055 23708 5550 23735
rect 5055 23697 5303 23708
rect 5055 23663 5061 23697
rect 5095 23674 5303 23697
rect 5337 23674 5395 23708
rect 5429 23674 5487 23708
rect 5521 23674 5550 23708
rect 5095 23663 5550 23674
rect 5055 23643 5550 23663
rect 5055 23625 5101 23643
rect 5055 23591 5061 23625
rect 5095 23591 5101 23625
rect 2466 23410 3837 23444
rect 2466 23277 2500 23410
rect 2658 23277 2692 23410
rect 2850 23277 2884 23410
rect 3042 23277 3076 23410
rect 3234 23277 3268 23410
rect 3426 23277 3460 23410
rect 3671 23320 3681 23372
rect 3733 23320 3743 23372
rect 3679 23319 3691 23320
rect 3725 23319 3737 23320
rect 3679 23313 3737 23319
rect 3534 23284 3580 23307
rect 2460 23242 2506 23277
rect 2460 23208 2466 23242
rect 2500 23208 2506 23242
rect 2460 23173 2506 23208
rect 2556 23242 2602 23277
rect 2556 23208 2562 23242
rect 2596 23208 2602 23242
rect 2556 23173 2602 23208
rect 2652 23242 2698 23277
rect 2652 23208 2658 23242
rect 2692 23208 2698 23242
rect 2652 23173 2698 23208
rect 2748 23242 2794 23277
rect 2748 23208 2754 23242
rect 2788 23208 2794 23242
rect 2748 23173 2794 23208
rect 2844 23242 2890 23277
rect 2844 23208 2850 23242
rect 2884 23208 2890 23242
rect 2844 23173 2890 23208
rect 2940 23242 2986 23277
rect 2940 23208 2946 23242
rect 2980 23208 2986 23242
rect 2940 23173 2986 23208
rect 3036 23242 3082 23277
rect 3036 23208 3042 23242
rect 3076 23208 3082 23242
rect 3036 23173 3082 23208
rect 3132 23242 3178 23277
rect 3132 23208 3138 23242
rect 3172 23208 3178 23242
rect 3132 23173 3178 23208
rect 3228 23242 3274 23277
rect 3228 23208 3234 23242
rect 3268 23208 3274 23242
rect 3228 23173 3274 23208
rect 3324 23242 3370 23277
rect 3324 23208 3330 23242
rect 3364 23208 3370 23242
rect 3324 23173 3370 23208
rect 3420 23242 3466 23277
rect 3420 23208 3426 23242
rect 3460 23208 3466 23242
rect 3420 23173 3466 23208
rect 3534 23250 3540 23284
rect 3574 23282 3580 23284
rect 3803 23282 3837 23410
rect 3574 23281 3680 23282
rect 3734 23281 3837 23282
rect 3574 23269 3687 23281
rect 3574 23250 3647 23269
rect 3534 23212 3647 23250
rect 3534 23178 3540 23212
rect 3574 23193 3647 23212
rect 3681 23193 3687 23269
rect 3574 23182 3687 23193
rect 3574 23178 3580 23182
rect 3641 23181 3687 23182
rect 3729 23269 3837 23281
rect 3987 23444 4021 23585
rect 4179 23444 4213 23585
rect 4371 23444 4405 23585
rect 4563 23444 4597 23585
rect 4755 23444 4789 23585
rect 4947 23444 4981 23585
rect 5055 23547 5101 23591
rect 5683 23498 5743 24751
rect 5177 23464 5743 23498
rect 5177 23444 5211 23464
rect 3987 23410 5211 23444
rect 3987 23277 4021 23410
rect 4179 23277 4213 23410
rect 4371 23277 4405 23410
rect 4563 23277 4597 23410
rect 4755 23277 4789 23410
rect 4947 23277 4981 23410
rect 5438 23406 5512 23407
rect 5326 23404 5400 23405
rect 5326 23352 5337 23404
rect 5389 23352 5400 23404
rect 5438 23354 5449 23406
rect 5501 23354 5512 23406
rect 5438 23353 5512 23354
rect 5326 23351 5400 23352
rect 5055 23284 5101 23307
rect 3729 23193 3735 23269
rect 3769 23193 3837 23269
rect 3729 23182 3837 23193
rect 3729 23181 3775 23182
rect 2450 23142 2516 23145
rect 2447 23090 2457 23142
rect 2509 23090 2519 23142
rect 2450 23085 2516 23090
rect 2562 23033 2596 23173
rect 2642 23142 2708 23145
rect 2638 23090 2648 23142
rect 2700 23090 2710 23142
rect 2642 23085 2708 23090
rect 2754 23033 2788 23173
rect 2834 23142 2900 23145
rect 2830 23090 2840 23142
rect 2892 23090 2902 23142
rect 2834 23085 2900 23090
rect 2946 23033 2980 23173
rect 3026 23142 3092 23145
rect 3022 23090 3032 23142
rect 3084 23090 3094 23142
rect 3026 23085 3092 23090
rect 3138 23033 3172 23173
rect 3218 23141 3284 23145
rect 3215 23089 3225 23141
rect 3277 23089 3287 23141
rect 3218 23085 3284 23089
rect 3330 23033 3364 23173
rect 3410 23141 3476 23145
rect 3407 23089 3417 23141
rect 3469 23089 3479 23141
rect 3534 23140 3580 23178
rect 3534 23106 3540 23140
rect 3574 23106 3580 23140
rect 3410 23085 3476 23089
rect 2282 22999 3364 23033
rect 3534 22923 3580 23106
rect 3803 23033 3837 23182
rect 3981 23242 4027 23277
rect 3981 23208 3987 23242
rect 4021 23208 4027 23242
rect 3981 23173 4027 23208
rect 4077 23242 4123 23277
rect 4077 23208 4083 23242
rect 4117 23208 4123 23242
rect 4077 23173 4123 23208
rect 4173 23242 4219 23277
rect 4173 23208 4179 23242
rect 4213 23208 4219 23242
rect 4173 23173 4219 23208
rect 4269 23242 4315 23277
rect 4269 23208 4275 23242
rect 4309 23208 4315 23242
rect 4269 23173 4315 23208
rect 4365 23242 4411 23277
rect 4365 23208 4371 23242
rect 4405 23208 4411 23242
rect 4365 23173 4411 23208
rect 4461 23242 4507 23277
rect 4461 23208 4467 23242
rect 4501 23208 4507 23242
rect 4461 23173 4507 23208
rect 4557 23242 4603 23277
rect 4557 23208 4563 23242
rect 4597 23208 4603 23242
rect 4557 23173 4603 23208
rect 4653 23242 4699 23277
rect 4653 23208 4659 23242
rect 4693 23208 4699 23242
rect 4653 23173 4699 23208
rect 4749 23242 4795 23277
rect 4749 23208 4755 23242
rect 4789 23208 4795 23242
rect 4749 23173 4795 23208
rect 4845 23242 4891 23277
rect 4845 23208 4851 23242
rect 4885 23208 4891 23242
rect 4845 23173 4891 23208
rect 4941 23242 4987 23277
rect 4941 23208 4947 23242
rect 4981 23208 4987 23242
rect 4941 23173 4987 23208
rect 5055 23250 5061 23284
rect 5095 23250 5101 23284
rect 5055 23212 5101 23250
rect 5055 23178 5061 23212
rect 5095 23195 5101 23212
rect 5095 23178 5550 23195
rect 3971 23142 4037 23145
rect 3968 23090 3978 23142
rect 4030 23090 4040 23142
rect 3971 23085 4037 23090
rect 4083 23033 4117 23173
rect 4163 23142 4229 23145
rect 4159 23090 4169 23142
rect 4221 23090 4231 23142
rect 4163 23085 4229 23090
rect 4275 23033 4309 23173
rect 4355 23142 4421 23145
rect 4351 23090 4361 23142
rect 4413 23090 4423 23142
rect 4355 23085 4421 23090
rect 4467 23033 4501 23173
rect 4547 23142 4613 23145
rect 4543 23090 4553 23142
rect 4605 23090 4615 23142
rect 4547 23085 4613 23090
rect 4659 23033 4693 23173
rect 4739 23141 4805 23145
rect 4736 23089 4746 23141
rect 4798 23089 4808 23141
rect 4739 23085 4805 23089
rect 4851 23033 4885 23173
rect 5055 23164 5550 23178
rect 4931 23141 4997 23145
rect 4928 23089 4938 23141
rect 4990 23089 5000 23141
rect 5055 23140 5303 23164
rect 5055 23106 5061 23140
rect 5095 23130 5303 23140
rect 5337 23130 5395 23164
rect 5429 23130 5487 23164
rect 5521 23130 5550 23164
rect 5095 23106 5550 23130
rect 5055 23099 5550 23106
rect 4931 23085 4997 23089
rect 3803 22999 4885 23033
rect 5055 22924 5101 23099
rect 129 22716 1211 22750
rect 129 22153 163 22716
rect 294 22606 304 22658
rect 356 22606 366 22658
rect 409 22566 443 22716
rect 487 22606 497 22658
rect 549 22606 559 22658
rect 601 22566 635 22716
rect 678 22606 688 22658
rect 740 22606 750 22658
rect 793 22566 827 22716
rect 870 22606 880 22658
rect 932 22606 942 22658
rect 985 22566 1019 22716
rect 1062 22606 1072 22658
rect 1124 22606 1134 22658
rect 1177 22566 1211 22716
rect 1254 22606 1264 22658
rect 1316 22606 1326 22658
rect 1381 22622 1427 22786
rect 2282 22720 3364 22754
rect 1381 22588 1387 22622
rect 1421 22588 1427 22622
rect 1512 22599 1522 22659
rect 1578 22599 1792 22659
rect 1852 22599 1862 22659
rect 307 22519 353 22566
rect 307 22485 313 22519
rect 347 22485 353 22519
rect 307 22447 353 22485
rect 307 22413 313 22447
rect 347 22413 353 22447
rect 307 22375 353 22413
rect 307 22341 313 22375
rect 347 22341 353 22375
rect 307 22294 353 22341
rect 403 22519 449 22566
rect 403 22485 409 22519
rect 443 22485 449 22519
rect 403 22447 449 22485
rect 403 22413 409 22447
rect 443 22413 449 22447
rect 403 22375 449 22413
rect 403 22341 409 22375
rect 443 22341 449 22375
rect 403 22294 449 22341
rect 499 22519 545 22566
rect 499 22485 505 22519
rect 539 22485 545 22519
rect 499 22447 545 22485
rect 499 22413 505 22447
rect 539 22413 545 22447
rect 499 22375 545 22413
rect 499 22341 505 22375
rect 539 22341 545 22375
rect 499 22294 545 22341
rect 595 22519 641 22566
rect 595 22485 601 22519
rect 635 22485 641 22519
rect 595 22447 641 22485
rect 595 22413 601 22447
rect 635 22413 641 22447
rect 595 22375 641 22413
rect 595 22341 601 22375
rect 635 22341 641 22375
rect 595 22294 641 22341
rect 691 22519 737 22566
rect 691 22485 697 22519
rect 731 22485 737 22519
rect 691 22447 737 22485
rect 691 22413 697 22447
rect 731 22413 737 22447
rect 691 22375 737 22413
rect 691 22341 697 22375
rect 731 22341 737 22375
rect 691 22294 737 22341
rect 787 22519 833 22566
rect 787 22485 793 22519
rect 827 22485 833 22519
rect 787 22447 833 22485
rect 787 22413 793 22447
rect 827 22413 833 22447
rect 787 22375 833 22413
rect 787 22341 793 22375
rect 827 22341 833 22375
rect 787 22294 833 22341
rect 883 22519 929 22566
rect 883 22485 889 22519
rect 923 22485 929 22519
rect 883 22447 929 22485
rect 883 22413 889 22447
rect 923 22413 929 22447
rect 883 22375 929 22413
rect 883 22341 889 22375
rect 923 22341 929 22375
rect 883 22294 929 22341
rect 979 22519 1025 22566
rect 979 22485 985 22519
rect 1019 22485 1025 22519
rect 979 22447 1025 22485
rect 979 22413 985 22447
rect 1019 22413 1025 22447
rect 979 22375 1025 22413
rect 979 22341 985 22375
rect 1019 22341 1025 22375
rect 979 22294 1025 22341
rect 1075 22519 1121 22566
rect 1075 22485 1081 22519
rect 1115 22485 1121 22519
rect 1075 22447 1121 22485
rect 1075 22413 1081 22447
rect 1115 22413 1121 22447
rect 1075 22375 1121 22413
rect 1075 22341 1081 22375
rect 1115 22341 1121 22375
rect 1075 22294 1121 22341
rect 1171 22519 1217 22566
rect 1171 22485 1177 22519
rect 1211 22485 1217 22519
rect 1171 22447 1217 22485
rect 1171 22413 1177 22447
rect 1211 22413 1217 22447
rect 1171 22375 1217 22413
rect 1171 22341 1177 22375
rect 1211 22341 1217 22375
rect 1171 22294 1217 22341
rect 1267 22519 1313 22566
rect 1267 22485 1273 22519
rect 1307 22485 1313 22519
rect 1267 22447 1313 22485
rect 1267 22413 1273 22447
rect 1307 22413 1313 22447
rect 1267 22375 1313 22413
rect 1267 22341 1273 22375
rect 1307 22341 1313 22375
rect 1267 22294 1313 22341
rect 1381 22550 1427 22588
rect 1381 22516 1387 22550
rect 1421 22516 1427 22550
rect 1381 22478 1427 22516
rect 1381 22444 1387 22478
rect 1421 22444 1427 22478
rect 1381 22406 1427 22444
rect 1381 22372 1387 22406
rect 1421 22372 1427 22406
rect 1381 22362 1427 22372
rect 1381 22360 2160 22362
rect 1381 22334 2056 22360
rect 1381 22309 1387 22334
rect 1380 22300 1387 22309
rect 1421 22300 2056 22334
rect 0 22119 163 22153
rect 129 21742 163 22119
rect 313 22153 347 22294
rect 505 22153 539 22294
rect 697 22153 731 22294
rect 889 22153 923 22294
rect 1081 22153 1115 22294
rect 1273 22153 1307 22294
rect 1380 22252 2056 22300
rect 2190 22252 2200 22360
rect 1380 22250 2160 22252
rect 2282 22157 2316 22720
rect 2447 22610 2457 22662
rect 2509 22610 2519 22662
rect 2562 22570 2596 22720
rect 2640 22610 2650 22662
rect 2702 22610 2712 22662
rect 2754 22570 2788 22720
rect 2831 22610 2841 22662
rect 2893 22610 2903 22662
rect 2946 22570 2980 22720
rect 3023 22610 3033 22662
rect 3085 22610 3095 22662
rect 3138 22570 3172 22720
rect 3215 22610 3225 22662
rect 3277 22610 3287 22662
rect 3330 22570 3364 22720
rect 3407 22610 3417 22662
rect 3469 22610 3479 22662
rect 3534 22626 3580 22834
rect 3534 22592 3540 22626
rect 3574 22592 3580 22626
rect 2460 22523 2506 22570
rect 2460 22489 2466 22523
rect 2500 22489 2506 22523
rect 2460 22451 2506 22489
rect 2460 22417 2466 22451
rect 2500 22417 2506 22451
rect 2460 22379 2506 22417
rect 2460 22345 2466 22379
rect 2500 22345 2506 22379
rect 2460 22298 2506 22345
rect 2556 22523 2602 22570
rect 2556 22489 2562 22523
rect 2596 22489 2602 22523
rect 2556 22451 2602 22489
rect 2556 22417 2562 22451
rect 2596 22417 2602 22451
rect 2556 22379 2602 22417
rect 2556 22345 2562 22379
rect 2596 22345 2602 22379
rect 2556 22298 2602 22345
rect 2652 22523 2698 22570
rect 2652 22489 2658 22523
rect 2692 22489 2698 22523
rect 2652 22451 2698 22489
rect 2652 22417 2658 22451
rect 2692 22417 2698 22451
rect 2652 22379 2698 22417
rect 2652 22345 2658 22379
rect 2692 22345 2698 22379
rect 2652 22298 2698 22345
rect 2748 22523 2794 22570
rect 2748 22489 2754 22523
rect 2788 22489 2794 22523
rect 2748 22451 2794 22489
rect 2748 22417 2754 22451
rect 2788 22417 2794 22451
rect 2748 22379 2794 22417
rect 2748 22345 2754 22379
rect 2788 22345 2794 22379
rect 2748 22298 2794 22345
rect 2844 22523 2890 22570
rect 2844 22489 2850 22523
rect 2884 22489 2890 22523
rect 2844 22451 2890 22489
rect 2844 22417 2850 22451
rect 2884 22417 2890 22451
rect 2844 22379 2890 22417
rect 2844 22345 2850 22379
rect 2884 22345 2890 22379
rect 2844 22298 2890 22345
rect 2940 22523 2986 22570
rect 2940 22489 2946 22523
rect 2980 22489 2986 22523
rect 2940 22451 2986 22489
rect 2940 22417 2946 22451
rect 2980 22417 2986 22451
rect 2940 22379 2986 22417
rect 2940 22345 2946 22379
rect 2980 22345 2986 22379
rect 2940 22298 2986 22345
rect 3036 22523 3082 22570
rect 3036 22489 3042 22523
rect 3076 22489 3082 22523
rect 3036 22451 3082 22489
rect 3036 22417 3042 22451
rect 3076 22417 3082 22451
rect 3036 22379 3082 22417
rect 3036 22345 3042 22379
rect 3076 22345 3082 22379
rect 3036 22298 3082 22345
rect 3132 22523 3178 22570
rect 3132 22489 3138 22523
rect 3172 22489 3178 22523
rect 3132 22451 3178 22489
rect 3132 22417 3138 22451
rect 3172 22417 3178 22451
rect 3132 22379 3178 22417
rect 3132 22345 3138 22379
rect 3172 22345 3178 22379
rect 3132 22298 3178 22345
rect 3228 22523 3274 22570
rect 3228 22489 3234 22523
rect 3268 22489 3274 22523
rect 3228 22451 3274 22489
rect 3228 22417 3234 22451
rect 3268 22417 3274 22451
rect 3228 22379 3274 22417
rect 3228 22345 3234 22379
rect 3268 22345 3274 22379
rect 3228 22298 3274 22345
rect 3324 22523 3370 22570
rect 3324 22489 3330 22523
rect 3364 22489 3370 22523
rect 3324 22451 3370 22489
rect 3324 22417 3330 22451
rect 3364 22417 3370 22451
rect 3324 22379 3370 22417
rect 3324 22345 3330 22379
rect 3364 22345 3370 22379
rect 3324 22298 3370 22345
rect 3420 22523 3466 22570
rect 3420 22489 3426 22523
rect 3460 22489 3466 22523
rect 3420 22451 3466 22489
rect 3420 22417 3426 22451
rect 3460 22417 3466 22451
rect 3420 22379 3466 22417
rect 3420 22345 3426 22379
rect 3460 22345 3466 22379
rect 3420 22298 3466 22345
rect 3534 22554 3580 22592
rect 3534 22520 3540 22554
rect 3574 22520 3580 22554
rect 3534 22482 3580 22520
rect 3534 22448 3540 22482
rect 3574 22448 3580 22482
rect 3534 22410 3580 22448
rect 3534 22376 3540 22410
rect 3574 22376 3580 22410
rect 3534 22338 3580 22376
rect 3534 22304 3540 22338
rect 3574 22304 3580 22338
rect 2101 22153 2316 22157
rect 313 22123 2316 22153
rect 313 22119 2141 22123
rect 313 21986 347 22119
rect 505 21986 539 22119
rect 697 21986 731 22119
rect 889 21986 923 22119
rect 1081 21986 1115 22119
rect 1273 21986 1307 22119
rect 1381 21993 1608 22016
rect 307 21951 353 21986
rect 307 21917 313 21951
rect 347 21917 353 21951
rect 307 21882 353 21917
rect 403 21951 449 21986
rect 403 21917 409 21951
rect 443 21917 449 21951
rect 403 21882 449 21917
rect 499 21951 545 21986
rect 499 21917 505 21951
rect 539 21917 545 21951
rect 499 21882 545 21917
rect 595 21951 641 21986
rect 595 21917 601 21951
rect 635 21917 641 21951
rect 595 21882 641 21917
rect 691 21951 737 21986
rect 691 21917 697 21951
rect 731 21917 737 21951
rect 691 21882 737 21917
rect 787 21951 833 21986
rect 787 21917 793 21951
rect 827 21917 833 21951
rect 787 21882 833 21917
rect 883 21951 929 21986
rect 883 21917 889 21951
rect 923 21917 929 21951
rect 883 21882 929 21917
rect 979 21951 1025 21986
rect 979 21917 985 21951
rect 1019 21917 1025 21951
rect 979 21882 1025 21917
rect 1075 21951 1121 21986
rect 1075 21917 1081 21951
rect 1115 21917 1121 21951
rect 1075 21882 1121 21917
rect 1171 21951 1217 21986
rect 1171 21917 1177 21951
rect 1211 21917 1217 21951
rect 1171 21882 1217 21917
rect 1267 21951 1313 21986
rect 1267 21917 1273 21951
rect 1307 21917 1313 21951
rect 1267 21882 1313 21917
rect 1381 21959 1387 21993
rect 1421 21959 1608 21993
rect 1381 21921 1608 21959
rect 1381 21887 1387 21921
rect 1421 21896 1608 21921
rect 1421 21887 1427 21896
rect 1560 21894 1608 21896
rect 1598 21892 1608 21894
rect 1720 21892 1730 22016
rect 297 21851 363 21854
rect 294 21799 304 21851
rect 356 21799 366 21851
rect 297 21794 363 21799
rect 409 21742 443 21882
rect 489 21851 555 21854
rect 485 21799 495 21851
rect 547 21799 557 21851
rect 489 21794 555 21799
rect 601 21742 635 21882
rect 681 21851 747 21854
rect 677 21799 687 21851
rect 739 21799 749 21851
rect 681 21794 747 21799
rect 793 21742 827 21882
rect 873 21851 939 21854
rect 869 21799 879 21851
rect 931 21799 941 21851
rect 873 21794 939 21799
rect 985 21742 1019 21882
rect 1065 21850 1131 21854
rect 1062 21798 1072 21850
rect 1124 21798 1134 21850
rect 1065 21794 1131 21798
rect 1177 21742 1211 21882
rect 1257 21850 1323 21854
rect 1254 21798 1264 21850
rect 1316 21798 1326 21850
rect 1381 21849 1427 21887
rect 1920 21854 1930 21856
rect 1381 21815 1387 21849
rect 1421 21815 1427 21849
rect 1257 21794 1323 21798
rect 129 21708 1211 21742
rect 1381 21672 1427 21815
rect 1458 21798 1468 21854
rect 1524 21800 1930 21854
rect 1986 21800 1996 21856
rect 1524 21798 1986 21800
rect 2282 21746 2316 22123
rect 2466 22157 2500 22298
rect 2658 22157 2692 22298
rect 2850 22157 2884 22298
rect 3042 22157 3076 22298
rect 3234 22157 3268 22298
rect 3426 22157 3460 22298
rect 3534 22260 3580 22304
rect 3803 22720 4885 22754
rect 3803 22157 3837 22720
rect 3968 22610 3978 22662
rect 4030 22610 4040 22662
rect 4083 22570 4117 22720
rect 4161 22610 4171 22662
rect 4223 22610 4233 22662
rect 4275 22570 4309 22720
rect 4352 22610 4362 22662
rect 4414 22610 4424 22662
rect 4467 22570 4501 22720
rect 4544 22610 4554 22662
rect 4606 22610 4616 22662
rect 4659 22570 4693 22720
rect 4736 22610 4746 22662
rect 4798 22610 4808 22662
rect 4851 22570 4885 22720
rect 4928 22610 4938 22662
rect 4990 22610 5000 22662
rect 5055 22626 5101 22831
rect 5055 22592 5061 22626
rect 5095 22592 5101 22626
rect 3981 22523 4027 22570
rect 3981 22489 3987 22523
rect 4021 22489 4027 22523
rect 3981 22451 4027 22489
rect 3981 22417 3987 22451
rect 4021 22417 4027 22451
rect 3981 22379 4027 22417
rect 3981 22345 3987 22379
rect 4021 22345 4027 22379
rect 3981 22298 4027 22345
rect 4077 22523 4123 22570
rect 4077 22489 4083 22523
rect 4117 22489 4123 22523
rect 4077 22451 4123 22489
rect 4077 22417 4083 22451
rect 4117 22417 4123 22451
rect 4077 22379 4123 22417
rect 4077 22345 4083 22379
rect 4117 22345 4123 22379
rect 4077 22298 4123 22345
rect 4173 22523 4219 22570
rect 4173 22489 4179 22523
rect 4213 22489 4219 22523
rect 4173 22451 4219 22489
rect 4173 22417 4179 22451
rect 4213 22417 4219 22451
rect 4173 22379 4219 22417
rect 4173 22345 4179 22379
rect 4213 22345 4219 22379
rect 4173 22298 4219 22345
rect 4269 22523 4315 22570
rect 4269 22489 4275 22523
rect 4309 22489 4315 22523
rect 4269 22451 4315 22489
rect 4269 22417 4275 22451
rect 4309 22417 4315 22451
rect 4269 22379 4315 22417
rect 4269 22345 4275 22379
rect 4309 22345 4315 22379
rect 4269 22298 4315 22345
rect 4365 22523 4411 22570
rect 4365 22489 4371 22523
rect 4405 22489 4411 22523
rect 4365 22451 4411 22489
rect 4365 22417 4371 22451
rect 4405 22417 4411 22451
rect 4365 22379 4411 22417
rect 4365 22345 4371 22379
rect 4405 22345 4411 22379
rect 4365 22298 4411 22345
rect 4461 22523 4507 22570
rect 4461 22489 4467 22523
rect 4501 22489 4507 22523
rect 4461 22451 4507 22489
rect 4461 22417 4467 22451
rect 4501 22417 4507 22451
rect 4461 22379 4507 22417
rect 4461 22345 4467 22379
rect 4501 22345 4507 22379
rect 4461 22298 4507 22345
rect 4557 22523 4603 22570
rect 4557 22489 4563 22523
rect 4597 22489 4603 22523
rect 4557 22451 4603 22489
rect 4557 22417 4563 22451
rect 4597 22417 4603 22451
rect 4557 22379 4603 22417
rect 4557 22345 4563 22379
rect 4597 22345 4603 22379
rect 4557 22298 4603 22345
rect 4653 22523 4699 22570
rect 4653 22489 4659 22523
rect 4693 22489 4699 22523
rect 4653 22451 4699 22489
rect 4653 22417 4659 22451
rect 4693 22417 4699 22451
rect 4653 22379 4699 22417
rect 4653 22345 4659 22379
rect 4693 22345 4699 22379
rect 4653 22298 4699 22345
rect 4749 22523 4795 22570
rect 4749 22489 4755 22523
rect 4789 22489 4795 22523
rect 4749 22451 4795 22489
rect 4749 22417 4755 22451
rect 4789 22417 4795 22451
rect 4749 22379 4795 22417
rect 4749 22345 4755 22379
rect 4789 22345 4795 22379
rect 4749 22298 4795 22345
rect 4845 22523 4891 22570
rect 4845 22489 4851 22523
rect 4885 22489 4891 22523
rect 4845 22451 4891 22489
rect 4845 22417 4851 22451
rect 4885 22417 4891 22451
rect 4845 22379 4891 22417
rect 4845 22345 4851 22379
rect 4885 22345 4891 22379
rect 4845 22298 4891 22345
rect 4941 22523 4987 22570
rect 4941 22489 4947 22523
rect 4981 22489 4987 22523
rect 4941 22451 4987 22489
rect 4941 22417 4947 22451
rect 4981 22417 4987 22451
rect 4941 22379 4987 22417
rect 4941 22345 4947 22379
rect 4981 22345 4987 22379
rect 4941 22298 4987 22345
rect 5055 22554 5101 22592
rect 5055 22520 5061 22554
rect 5095 22520 5101 22554
rect 5055 22482 5101 22520
rect 5055 22448 5061 22482
rect 5095 22451 5101 22482
rect 5274 22451 5550 22452
rect 5095 22448 5550 22451
rect 5055 22421 5550 22448
rect 5055 22410 5303 22421
rect 5055 22376 5061 22410
rect 5095 22387 5303 22410
rect 5337 22387 5395 22421
rect 5429 22387 5487 22421
rect 5521 22387 5550 22421
rect 5095 22376 5550 22387
rect 5055 22356 5550 22376
rect 5055 22338 5101 22356
rect 5055 22304 5061 22338
rect 5095 22304 5101 22338
rect 2466 22123 3837 22157
rect 2466 21990 2500 22123
rect 2658 21990 2692 22123
rect 2850 21990 2884 22123
rect 3042 21990 3076 22123
rect 3234 21990 3268 22123
rect 3426 21990 3460 22123
rect 3671 22033 3681 22085
rect 3733 22033 3743 22085
rect 3679 22032 3691 22033
rect 3725 22032 3737 22033
rect 3679 22026 3737 22032
rect 3534 21997 3580 22020
rect 2460 21955 2506 21990
rect 2460 21921 2466 21955
rect 2500 21921 2506 21955
rect 2460 21886 2506 21921
rect 2556 21955 2602 21990
rect 2556 21921 2562 21955
rect 2596 21921 2602 21955
rect 2556 21886 2602 21921
rect 2652 21955 2698 21990
rect 2652 21921 2658 21955
rect 2692 21921 2698 21955
rect 2652 21886 2698 21921
rect 2748 21955 2794 21990
rect 2748 21921 2754 21955
rect 2788 21921 2794 21955
rect 2748 21886 2794 21921
rect 2844 21955 2890 21990
rect 2844 21921 2850 21955
rect 2884 21921 2890 21955
rect 2844 21886 2890 21921
rect 2940 21955 2986 21990
rect 2940 21921 2946 21955
rect 2980 21921 2986 21955
rect 2940 21886 2986 21921
rect 3036 21955 3082 21990
rect 3036 21921 3042 21955
rect 3076 21921 3082 21955
rect 3036 21886 3082 21921
rect 3132 21955 3178 21990
rect 3132 21921 3138 21955
rect 3172 21921 3178 21955
rect 3132 21886 3178 21921
rect 3228 21955 3274 21990
rect 3228 21921 3234 21955
rect 3268 21921 3274 21955
rect 3228 21886 3274 21921
rect 3324 21955 3370 21990
rect 3324 21921 3330 21955
rect 3364 21921 3370 21955
rect 3324 21886 3370 21921
rect 3420 21955 3466 21990
rect 3420 21921 3426 21955
rect 3460 21921 3466 21955
rect 3420 21886 3466 21921
rect 3534 21963 3540 21997
rect 3574 21995 3580 21997
rect 3803 21995 3837 22123
rect 3574 21994 3680 21995
rect 3734 21994 3837 21995
rect 3574 21982 3687 21994
rect 3574 21963 3647 21982
rect 3534 21925 3647 21963
rect 3534 21891 3540 21925
rect 3574 21906 3647 21925
rect 3681 21906 3687 21982
rect 3574 21895 3687 21906
rect 3574 21891 3580 21895
rect 3641 21894 3687 21895
rect 3729 21982 3837 21994
rect 3987 22157 4021 22298
rect 4179 22157 4213 22298
rect 4371 22157 4405 22298
rect 4563 22157 4597 22298
rect 4755 22157 4789 22298
rect 4947 22157 4981 22298
rect 5055 22260 5101 22304
rect 5683 22211 5743 23464
rect 5177 22177 5743 22211
rect 5177 22157 5211 22177
rect 3987 22123 5211 22157
rect 3987 21990 4021 22123
rect 4179 21990 4213 22123
rect 4371 21990 4405 22123
rect 4563 21990 4597 22123
rect 4755 21990 4789 22123
rect 4947 21990 4981 22123
rect 5438 22119 5512 22120
rect 5326 22117 5400 22118
rect 5326 22065 5337 22117
rect 5389 22065 5400 22117
rect 5438 22067 5449 22119
rect 5501 22067 5512 22119
rect 5438 22066 5512 22067
rect 5326 22064 5400 22065
rect 5055 21997 5101 22020
rect 3729 21906 3735 21982
rect 3769 21906 3837 21982
rect 3729 21895 3837 21906
rect 3729 21894 3775 21895
rect 2450 21855 2516 21858
rect 2447 21803 2457 21855
rect 2509 21803 2519 21855
rect 2450 21798 2516 21803
rect 2562 21746 2596 21886
rect 2642 21855 2708 21858
rect 2638 21803 2648 21855
rect 2700 21803 2710 21855
rect 2642 21798 2708 21803
rect 2754 21746 2788 21886
rect 2834 21855 2900 21858
rect 2830 21803 2840 21855
rect 2892 21803 2902 21855
rect 2834 21798 2900 21803
rect 2946 21746 2980 21886
rect 3026 21855 3092 21858
rect 3022 21803 3032 21855
rect 3084 21803 3094 21855
rect 3026 21798 3092 21803
rect 3138 21746 3172 21886
rect 3218 21854 3284 21858
rect 3215 21802 3225 21854
rect 3277 21802 3287 21854
rect 3218 21798 3284 21802
rect 3330 21746 3364 21886
rect 3410 21854 3476 21858
rect 3407 21802 3417 21854
rect 3469 21802 3479 21854
rect 3534 21853 3580 21891
rect 3534 21819 3540 21853
rect 3574 21819 3580 21853
rect 3410 21798 3476 21802
rect 2282 21712 3364 21746
rect 3534 21636 3580 21819
rect 3803 21746 3837 21895
rect 3981 21955 4027 21990
rect 3981 21921 3987 21955
rect 4021 21921 4027 21955
rect 3981 21886 4027 21921
rect 4077 21955 4123 21990
rect 4077 21921 4083 21955
rect 4117 21921 4123 21955
rect 4077 21886 4123 21921
rect 4173 21955 4219 21990
rect 4173 21921 4179 21955
rect 4213 21921 4219 21955
rect 4173 21886 4219 21921
rect 4269 21955 4315 21990
rect 4269 21921 4275 21955
rect 4309 21921 4315 21955
rect 4269 21886 4315 21921
rect 4365 21955 4411 21990
rect 4365 21921 4371 21955
rect 4405 21921 4411 21955
rect 4365 21886 4411 21921
rect 4461 21955 4507 21990
rect 4461 21921 4467 21955
rect 4501 21921 4507 21955
rect 4461 21886 4507 21921
rect 4557 21955 4603 21990
rect 4557 21921 4563 21955
rect 4597 21921 4603 21955
rect 4557 21886 4603 21921
rect 4653 21955 4699 21990
rect 4653 21921 4659 21955
rect 4693 21921 4699 21955
rect 4653 21886 4699 21921
rect 4749 21955 4795 21990
rect 4749 21921 4755 21955
rect 4789 21921 4795 21955
rect 4749 21886 4795 21921
rect 4845 21955 4891 21990
rect 4845 21921 4851 21955
rect 4885 21921 4891 21955
rect 4845 21886 4891 21921
rect 4941 21955 4987 21990
rect 4941 21921 4947 21955
rect 4981 21921 4987 21955
rect 4941 21886 4987 21921
rect 5055 21963 5061 21997
rect 5095 21963 5101 21997
rect 5055 21925 5101 21963
rect 5055 21891 5061 21925
rect 5095 21908 5101 21925
rect 5095 21891 5550 21908
rect 3971 21855 4037 21858
rect 3968 21803 3978 21855
rect 4030 21803 4040 21855
rect 3971 21798 4037 21803
rect 4083 21746 4117 21886
rect 4163 21855 4229 21858
rect 4159 21803 4169 21855
rect 4221 21803 4231 21855
rect 4163 21798 4229 21803
rect 4275 21746 4309 21886
rect 4355 21855 4421 21858
rect 4351 21803 4361 21855
rect 4413 21803 4423 21855
rect 4355 21798 4421 21803
rect 4467 21746 4501 21886
rect 4547 21855 4613 21858
rect 4543 21803 4553 21855
rect 4605 21803 4615 21855
rect 4547 21798 4613 21803
rect 4659 21746 4693 21886
rect 4739 21854 4805 21858
rect 4736 21802 4746 21854
rect 4798 21802 4808 21854
rect 4739 21798 4805 21802
rect 4851 21746 4885 21886
rect 5055 21877 5550 21891
rect 4931 21854 4997 21858
rect 4928 21802 4938 21854
rect 4990 21802 5000 21854
rect 5055 21853 5303 21877
rect 5055 21819 5061 21853
rect 5095 21843 5303 21853
rect 5337 21843 5395 21877
rect 5429 21843 5487 21877
rect 5521 21843 5550 21877
rect 5095 21819 5550 21843
rect 5055 21812 5550 21819
rect 4931 21798 4997 21802
rect 3803 21712 4885 21746
rect 5055 21637 5101 21812
rect 129 21429 1211 21463
rect 129 20866 163 21429
rect 294 21319 304 21371
rect 356 21319 366 21371
rect 409 21279 443 21429
rect 487 21319 497 21371
rect 549 21319 559 21371
rect 601 21279 635 21429
rect 678 21319 688 21371
rect 740 21319 750 21371
rect 793 21279 827 21429
rect 870 21319 880 21371
rect 932 21319 942 21371
rect 985 21279 1019 21429
rect 1062 21319 1072 21371
rect 1124 21319 1134 21371
rect 1177 21279 1211 21429
rect 1254 21319 1264 21371
rect 1316 21319 1326 21371
rect 1381 21335 1427 21499
rect 2282 21433 3364 21467
rect 1381 21301 1387 21335
rect 1421 21301 1427 21335
rect 1512 21312 1522 21372
rect 1578 21312 1792 21372
rect 1852 21312 1862 21372
rect 307 21232 353 21279
rect 307 21198 313 21232
rect 347 21198 353 21232
rect 307 21160 353 21198
rect 307 21126 313 21160
rect 347 21126 353 21160
rect 307 21088 353 21126
rect 307 21054 313 21088
rect 347 21054 353 21088
rect 307 21007 353 21054
rect 403 21232 449 21279
rect 403 21198 409 21232
rect 443 21198 449 21232
rect 403 21160 449 21198
rect 403 21126 409 21160
rect 443 21126 449 21160
rect 403 21088 449 21126
rect 403 21054 409 21088
rect 443 21054 449 21088
rect 403 21007 449 21054
rect 499 21232 545 21279
rect 499 21198 505 21232
rect 539 21198 545 21232
rect 499 21160 545 21198
rect 499 21126 505 21160
rect 539 21126 545 21160
rect 499 21088 545 21126
rect 499 21054 505 21088
rect 539 21054 545 21088
rect 499 21007 545 21054
rect 595 21232 641 21279
rect 595 21198 601 21232
rect 635 21198 641 21232
rect 595 21160 641 21198
rect 595 21126 601 21160
rect 635 21126 641 21160
rect 595 21088 641 21126
rect 595 21054 601 21088
rect 635 21054 641 21088
rect 595 21007 641 21054
rect 691 21232 737 21279
rect 691 21198 697 21232
rect 731 21198 737 21232
rect 691 21160 737 21198
rect 691 21126 697 21160
rect 731 21126 737 21160
rect 691 21088 737 21126
rect 691 21054 697 21088
rect 731 21054 737 21088
rect 691 21007 737 21054
rect 787 21232 833 21279
rect 787 21198 793 21232
rect 827 21198 833 21232
rect 787 21160 833 21198
rect 787 21126 793 21160
rect 827 21126 833 21160
rect 787 21088 833 21126
rect 787 21054 793 21088
rect 827 21054 833 21088
rect 787 21007 833 21054
rect 883 21232 929 21279
rect 883 21198 889 21232
rect 923 21198 929 21232
rect 883 21160 929 21198
rect 883 21126 889 21160
rect 923 21126 929 21160
rect 883 21088 929 21126
rect 883 21054 889 21088
rect 923 21054 929 21088
rect 883 21007 929 21054
rect 979 21232 1025 21279
rect 979 21198 985 21232
rect 1019 21198 1025 21232
rect 979 21160 1025 21198
rect 979 21126 985 21160
rect 1019 21126 1025 21160
rect 979 21088 1025 21126
rect 979 21054 985 21088
rect 1019 21054 1025 21088
rect 979 21007 1025 21054
rect 1075 21232 1121 21279
rect 1075 21198 1081 21232
rect 1115 21198 1121 21232
rect 1075 21160 1121 21198
rect 1075 21126 1081 21160
rect 1115 21126 1121 21160
rect 1075 21088 1121 21126
rect 1075 21054 1081 21088
rect 1115 21054 1121 21088
rect 1075 21007 1121 21054
rect 1171 21232 1217 21279
rect 1171 21198 1177 21232
rect 1211 21198 1217 21232
rect 1171 21160 1217 21198
rect 1171 21126 1177 21160
rect 1211 21126 1217 21160
rect 1171 21088 1217 21126
rect 1171 21054 1177 21088
rect 1211 21054 1217 21088
rect 1171 21007 1217 21054
rect 1267 21232 1313 21279
rect 1267 21198 1273 21232
rect 1307 21198 1313 21232
rect 1267 21160 1313 21198
rect 1267 21126 1273 21160
rect 1307 21126 1313 21160
rect 1267 21088 1313 21126
rect 1267 21054 1273 21088
rect 1307 21054 1313 21088
rect 1267 21007 1313 21054
rect 1381 21263 1427 21301
rect 1381 21229 1387 21263
rect 1421 21229 1427 21263
rect 1381 21191 1427 21229
rect 1381 21157 1387 21191
rect 1421 21157 1427 21191
rect 1381 21119 1427 21157
rect 1381 21085 1387 21119
rect 1421 21085 1427 21119
rect 1381 21075 1427 21085
rect 1381 21073 2160 21075
rect 1381 21047 2056 21073
rect 1381 21022 1387 21047
rect 1380 21013 1387 21022
rect 1421 21013 2056 21047
rect 0 20832 163 20866
rect 129 20455 163 20832
rect 313 20866 347 21007
rect 505 20866 539 21007
rect 697 20866 731 21007
rect 889 20866 923 21007
rect 1081 20866 1115 21007
rect 1273 20866 1307 21007
rect 1380 20965 2056 21013
rect 2190 20965 2200 21073
rect 1380 20963 2160 20965
rect 2282 20870 2316 21433
rect 2447 21323 2457 21375
rect 2509 21323 2519 21375
rect 2562 21283 2596 21433
rect 2640 21323 2650 21375
rect 2702 21323 2712 21375
rect 2754 21283 2788 21433
rect 2831 21323 2841 21375
rect 2893 21323 2903 21375
rect 2946 21283 2980 21433
rect 3023 21323 3033 21375
rect 3085 21323 3095 21375
rect 3138 21283 3172 21433
rect 3215 21323 3225 21375
rect 3277 21323 3287 21375
rect 3330 21283 3364 21433
rect 3407 21323 3417 21375
rect 3469 21323 3479 21375
rect 3534 21339 3580 21547
rect 3534 21305 3540 21339
rect 3574 21305 3580 21339
rect 2460 21236 2506 21283
rect 2460 21202 2466 21236
rect 2500 21202 2506 21236
rect 2460 21164 2506 21202
rect 2460 21130 2466 21164
rect 2500 21130 2506 21164
rect 2460 21092 2506 21130
rect 2460 21058 2466 21092
rect 2500 21058 2506 21092
rect 2460 21011 2506 21058
rect 2556 21236 2602 21283
rect 2556 21202 2562 21236
rect 2596 21202 2602 21236
rect 2556 21164 2602 21202
rect 2556 21130 2562 21164
rect 2596 21130 2602 21164
rect 2556 21092 2602 21130
rect 2556 21058 2562 21092
rect 2596 21058 2602 21092
rect 2556 21011 2602 21058
rect 2652 21236 2698 21283
rect 2652 21202 2658 21236
rect 2692 21202 2698 21236
rect 2652 21164 2698 21202
rect 2652 21130 2658 21164
rect 2692 21130 2698 21164
rect 2652 21092 2698 21130
rect 2652 21058 2658 21092
rect 2692 21058 2698 21092
rect 2652 21011 2698 21058
rect 2748 21236 2794 21283
rect 2748 21202 2754 21236
rect 2788 21202 2794 21236
rect 2748 21164 2794 21202
rect 2748 21130 2754 21164
rect 2788 21130 2794 21164
rect 2748 21092 2794 21130
rect 2748 21058 2754 21092
rect 2788 21058 2794 21092
rect 2748 21011 2794 21058
rect 2844 21236 2890 21283
rect 2844 21202 2850 21236
rect 2884 21202 2890 21236
rect 2844 21164 2890 21202
rect 2844 21130 2850 21164
rect 2884 21130 2890 21164
rect 2844 21092 2890 21130
rect 2844 21058 2850 21092
rect 2884 21058 2890 21092
rect 2844 21011 2890 21058
rect 2940 21236 2986 21283
rect 2940 21202 2946 21236
rect 2980 21202 2986 21236
rect 2940 21164 2986 21202
rect 2940 21130 2946 21164
rect 2980 21130 2986 21164
rect 2940 21092 2986 21130
rect 2940 21058 2946 21092
rect 2980 21058 2986 21092
rect 2940 21011 2986 21058
rect 3036 21236 3082 21283
rect 3036 21202 3042 21236
rect 3076 21202 3082 21236
rect 3036 21164 3082 21202
rect 3036 21130 3042 21164
rect 3076 21130 3082 21164
rect 3036 21092 3082 21130
rect 3036 21058 3042 21092
rect 3076 21058 3082 21092
rect 3036 21011 3082 21058
rect 3132 21236 3178 21283
rect 3132 21202 3138 21236
rect 3172 21202 3178 21236
rect 3132 21164 3178 21202
rect 3132 21130 3138 21164
rect 3172 21130 3178 21164
rect 3132 21092 3178 21130
rect 3132 21058 3138 21092
rect 3172 21058 3178 21092
rect 3132 21011 3178 21058
rect 3228 21236 3274 21283
rect 3228 21202 3234 21236
rect 3268 21202 3274 21236
rect 3228 21164 3274 21202
rect 3228 21130 3234 21164
rect 3268 21130 3274 21164
rect 3228 21092 3274 21130
rect 3228 21058 3234 21092
rect 3268 21058 3274 21092
rect 3228 21011 3274 21058
rect 3324 21236 3370 21283
rect 3324 21202 3330 21236
rect 3364 21202 3370 21236
rect 3324 21164 3370 21202
rect 3324 21130 3330 21164
rect 3364 21130 3370 21164
rect 3324 21092 3370 21130
rect 3324 21058 3330 21092
rect 3364 21058 3370 21092
rect 3324 21011 3370 21058
rect 3420 21236 3466 21283
rect 3420 21202 3426 21236
rect 3460 21202 3466 21236
rect 3420 21164 3466 21202
rect 3420 21130 3426 21164
rect 3460 21130 3466 21164
rect 3420 21092 3466 21130
rect 3420 21058 3426 21092
rect 3460 21058 3466 21092
rect 3420 21011 3466 21058
rect 3534 21267 3580 21305
rect 3534 21233 3540 21267
rect 3574 21233 3580 21267
rect 3534 21195 3580 21233
rect 3534 21161 3540 21195
rect 3574 21161 3580 21195
rect 3534 21123 3580 21161
rect 3534 21089 3540 21123
rect 3574 21089 3580 21123
rect 3534 21051 3580 21089
rect 3534 21017 3540 21051
rect 3574 21017 3580 21051
rect 2101 20866 2316 20870
rect 313 20836 2316 20866
rect 313 20832 2141 20836
rect 313 20699 347 20832
rect 505 20699 539 20832
rect 697 20699 731 20832
rect 889 20699 923 20832
rect 1081 20699 1115 20832
rect 1273 20699 1307 20832
rect 1381 20706 1608 20729
rect 307 20664 353 20699
rect 307 20630 313 20664
rect 347 20630 353 20664
rect 307 20595 353 20630
rect 403 20664 449 20699
rect 403 20630 409 20664
rect 443 20630 449 20664
rect 403 20595 449 20630
rect 499 20664 545 20699
rect 499 20630 505 20664
rect 539 20630 545 20664
rect 499 20595 545 20630
rect 595 20664 641 20699
rect 595 20630 601 20664
rect 635 20630 641 20664
rect 595 20595 641 20630
rect 691 20664 737 20699
rect 691 20630 697 20664
rect 731 20630 737 20664
rect 691 20595 737 20630
rect 787 20664 833 20699
rect 787 20630 793 20664
rect 827 20630 833 20664
rect 787 20595 833 20630
rect 883 20664 929 20699
rect 883 20630 889 20664
rect 923 20630 929 20664
rect 883 20595 929 20630
rect 979 20664 1025 20699
rect 979 20630 985 20664
rect 1019 20630 1025 20664
rect 979 20595 1025 20630
rect 1075 20664 1121 20699
rect 1075 20630 1081 20664
rect 1115 20630 1121 20664
rect 1075 20595 1121 20630
rect 1171 20664 1217 20699
rect 1171 20630 1177 20664
rect 1211 20630 1217 20664
rect 1171 20595 1217 20630
rect 1267 20664 1313 20699
rect 1267 20630 1273 20664
rect 1307 20630 1313 20664
rect 1267 20595 1313 20630
rect 1381 20672 1387 20706
rect 1421 20672 1608 20706
rect 1381 20634 1608 20672
rect 1381 20600 1387 20634
rect 1421 20609 1608 20634
rect 1421 20600 1427 20609
rect 1560 20607 1608 20609
rect 1598 20605 1608 20607
rect 1720 20605 1730 20729
rect 297 20564 363 20567
rect 294 20512 304 20564
rect 356 20512 366 20564
rect 297 20507 363 20512
rect 409 20455 443 20595
rect 489 20564 555 20567
rect 485 20512 495 20564
rect 547 20512 557 20564
rect 489 20507 555 20512
rect 601 20455 635 20595
rect 681 20564 747 20567
rect 677 20512 687 20564
rect 739 20512 749 20564
rect 681 20507 747 20512
rect 793 20455 827 20595
rect 873 20564 939 20567
rect 869 20512 879 20564
rect 931 20512 941 20564
rect 873 20507 939 20512
rect 985 20455 1019 20595
rect 1065 20563 1131 20567
rect 1062 20511 1072 20563
rect 1124 20511 1134 20563
rect 1065 20507 1131 20511
rect 1177 20455 1211 20595
rect 1257 20563 1323 20567
rect 1254 20511 1264 20563
rect 1316 20511 1326 20563
rect 1381 20562 1427 20600
rect 1920 20567 1930 20569
rect 1381 20528 1387 20562
rect 1421 20528 1427 20562
rect 1257 20507 1323 20511
rect 129 20421 1211 20455
rect 1381 20385 1427 20528
rect 1458 20511 1468 20567
rect 1524 20513 1930 20567
rect 1986 20513 1996 20569
rect 1524 20511 1986 20513
rect 2282 20459 2316 20836
rect 2466 20870 2500 21011
rect 2658 20870 2692 21011
rect 2850 20870 2884 21011
rect 3042 20870 3076 21011
rect 3234 20870 3268 21011
rect 3426 20870 3460 21011
rect 3534 20973 3580 21017
rect 3803 21433 4885 21467
rect 3803 20870 3837 21433
rect 3968 21323 3978 21375
rect 4030 21323 4040 21375
rect 4083 21283 4117 21433
rect 4161 21323 4171 21375
rect 4223 21323 4233 21375
rect 4275 21283 4309 21433
rect 4352 21323 4362 21375
rect 4414 21323 4424 21375
rect 4467 21283 4501 21433
rect 4544 21323 4554 21375
rect 4606 21323 4616 21375
rect 4659 21283 4693 21433
rect 4736 21323 4746 21375
rect 4798 21323 4808 21375
rect 4851 21283 4885 21433
rect 4928 21323 4938 21375
rect 4990 21323 5000 21375
rect 5055 21339 5101 21544
rect 5055 21305 5061 21339
rect 5095 21305 5101 21339
rect 3981 21236 4027 21283
rect 3981 21202 3987 21236
rect 4021 21202 4027 21236
rect 3981 21164 4027 21202
rect 3981 21130 3987 21164
rect 4021 21130 4027 21164
rect 3981 21092 4027 21130
rect 3981 21058 3987 21092
rect 4021 21058 4027 21092
rect 3981 21011 4027 21058
rect 4077 21236 4123 21283
rect 4077 21202 4083 21236
rect 4117 21202 4123 21236
rect 4077 21164 4123 21202
rect 4077 21130 4083 21164
rect 4117 21130 4123 21164
rect 4077 21092 4123 21130
rect 4077 21058 4083 21092
rect 4117 21058 4123 21092
rect 4077 21011 4123 21058
rect 4173 21236 4219 21283
rect 4173 21202 4179 21236
rect 4213 21202 4219 21236
rect 4173 21164 4219 21202
rect 4173 21130 4179 21164
rect 4213 21130 4219 21164
rect 4173 21092 4219 21130
rect 4173 21058 4179 21092
rect 4213 21058 4219 21092
rect 4173 21011 4219 21058
rect 4269 21236 4315 21283
rect 4269 21202 4275 21236
rect 4309 21202 4315 21236
rect 4269 21164 4315 21202
rect 4269 21130 4275 21164
rect 4309 21130 4315 21164
rect 4269 21092 4315 21130
rect 4269 21058 4275 21092
rect 4309 21058 4315 21092
rect 4269 21011 4315 21058
rect 4365 21236 4411 21283
rect 4365 21202 4371 21236
rect 4405 21202 4411 21236
rect 4365 21164 4411 21202
rect 4365 21130 4371 21164
rect 4405 21130 4411 21164
rect 4365 21092 4411 21130
rect 4365 21058 4371 21092
rect 4405 21058 4411 21092
rect 4365 21011 4411 21058
rect 4461 21236 4507 21283
rect 4461 21202 4467 21236
rect 4501 21202 4507 21236
rect 4461 21164 4507 21202
rect 4461 21130 4467 21164
rect 4501 21130 4507 21164
rect 4461 21092 4507 21130
rect 4461 21058 4467 21092
rect 4501 21058 4507 21092
rect 4461 21011 4507 21058
rect 4557 21236 4603 21283
rect 4557 21202 4563 21236
rect 4597 21202 4603 21236
rect 4557 21164 4603 21202
rect 4557 21130 4563 21164
rect 4597 21130 4603 21164
rect 4557 21092 4603 21130
rect 4557 21058 4563 21092
rect 4597 21058 4603 21092
rect 4557 21011 4603 21058
rect 4653 21236 4699 21283
rect 4653 21202 4659 21236
rect 4693 21202 4699 21236
rect 4653 21164 4699 21202
rect 4653 21130 4659 21164
rect 4693 21130 4699 21164
rect 4653 21092 4699 21130
rect 4653 21058 4659 21092
rect 4693 21058 4699 21092
rect 4653 21011 4699 21058
rect 4749 21236 4795 21283
rect 4749 21202 4755 21236
rect 4789 21202 4795 21236
rect 4749 21164 4795 21202
rect 4749 21130 4755 21164
rect 4789 21130 4795 21164
rect 4749 21092 4795 21130
rect 4749 21058 4755 21092
rect 4789 21058 4795 21092
rect 4749 21011 4795 21058
rect 4845 21236 4891 21283
rect 4845 21202 4851 21236
rect 4885 21202 4891 21236
rect 4845 21164 4891 21202
rect 4845 21130 4851 21164
rect 4885 21130 4891 21164
rect 4845 21092 4891 21130
rect 4845 21058 4851 21092
rect 4885 21058 4891 21092
rect 4845 21011 4891 21058
rect 4941 21236 4987 21283
rect 4941 21202 4947 21236
rect 4981 21202 4987 21236
rect 4941 21164 4987 21202
rect 4941 21130 4947 21164
rect 4981 21130 4987 21164
rect 4941 21092 4987 21130
rect 4941 21058 4947 21092
rect 4981 21058 4987 21092
rect 4941 21011 4987 21058
rect 5055 21267 5101 21305
rect 5055 21233 5061 21267
rect 5095 21233 5101 21267
rect 5055 21195 5101 21233
rect 5055 21161 5061 21195
rect 5095 21164 5101 21195
rect 5274 21164 5550 21165
rect 5095 21161 5550 21164
rect 5055 21134 5550 21161
rect 5055 21123 5303 21134
rect 5055 21089 5061 21123
rect 5095 21100 5303 21123
rect 5337 21100 5395 21134
rect 5429 21100 5487 21134
rect 5521 21100 5550 21134
rect 5095 21089 5550 21100
rect 5055 21069 5550 21089
rect 5055 21051 5101 21069
rect 5055 21017 5061 21051
rect 5095 21017 5101 21051
rect 2466 20836 3837 20870
rect 2466 20703 2500 20836
rect 2658 20703 2692 20836
rect 2850 20703 2884 20836
rect 3042 20703 3076 20836
rect 3234 20703 3268 20836
rect 3426 20703 3460 20836
rect 3671 20746 3681 20798
rect 3733 20746 3743 20798
rect 3679 20745 3691 20746
rect 3725 20745 3737 20746
rect 3679 20739 3737 20745
rect 3534 20710 3580 20733
rect 2460 20668 2506 20703
rect 2460 20634 2466 20668
rect 2500 20634 2506 20668
rect 2460 20599 2506 20634
rect 2556 20668 2602 20703
rect 2556 20634 2562 20668
rect 2596 20634 2602 20668
rect 2556 20599 2602 20634
rect 2652 20668 2698 20703
rect 2652 20634 2658 20668
rect 2692 20634 2698 20668
rect 2652 20599 2698 20634
rect 2748 20668 2794 20703
rect 2748 20634 2754 20668
rect 2788 20634 2794 20668
rect 2748 20599 2794 20634
rect 2844 20668 2890 20703
rect 2844 20634 2850 20668
rect 2884 20634 2890 20668
rect 2844 20599 2890 20634
rect 2940 20668 2986 20703
rect 2940 20634 2946 20668
rect 2980 20634 2986 20668
rect 2940 20599 2986 20634
rect 3036 20668 3082 20703
rect 3036 20634 3042 20668
rect 3076 20634 3082 20668
rect 3036 20599 3082 20634
rect 3132 20668 3178 20703
rect 3132 20634 3138 20668
rect 3172 20634 3178 20668
rect 3132 20599 3178 20634
rect 3228 20668 3274 20703
rect 3228 20634 3234 20668
rect 3268 20634 3274 20668
rect 3228 20599 3274 20634
rect 3324 20668 3370 20703
rect 3324 20634 3330 20668
rect 3364 20634 3370 20668
rect 3324 20599 3370 20634
rect 3420 20668 3466 20703
rect 3420 20634 3426 20668
rect 3460 20634 3466 20668
rect 3420 20599 3466 20634
rect 3534 20676 3540 20710
rect 3574 20708 3580 20710
rect 3803 20708 3837 20836
rect 3574 20707 3680 20708
rect 3734 20707 3837 20708
rect 3574 20695 3687 20707
rect 3574 20676 3647 20695
rect 3534 20638 3647 20676
rect 3534 20604 3540 20638
rect 3574 20619 3647 20638
rect 3681 20619 3687 20695
rect 3574 20608 3687 20619
rect 3574 20604 3580 20608
rect 3641 20607 3687 20608
rect 3729 20695 3837 20707
rect 3987 20870 4021 21011
rect 4179 20870 4213 21011
rect 4371 20870 4405 21011
rect 4563 20870 4597 21011
rect 4755 20870 4789 21011
rect 4947 20870 4981 21011
rect 5055 20973 5101 21017
rect 5683 20924 5743 22177
rect 5177 20890 5743 20924
rect 5177 20870 5211 20890
rect 3987 20836 5211 20870
rect 3987 20703 4021 20836
rect 4179 20703 4213 20836
rect 4371 20703 4405 20836
rect 4563 20703 4597 20836
rect 4755 20703 4789 20836
rect 4947 20703 4981 20836
rect 5438 20832 5512 20833
rect 5326 20830 5400 20831
rect 5326 20778 5337 20830
rect 5389 20778 5400 20830
rect 5438 20780 5449 20832
rect 5501 20780 5512 20832
rect 5438 20779 5512 20780
rect 5326 20777 5400 20778
rect 5055 20710 5101 20733
rect 3729 20619 3735 20695
rect 3769 20619 3837 20695
rect 3729 20608 3837 20619
rect 3729 20607 3775 20608
rect 2450 20568 2516 20571
rect 2447 20516 2457 20568
rect 2509 20516 2519 20568
rect 2450 20511 2516 20516
rect 2562 20459 2596 20599
rect 2642 20568 2708 20571
rect 2638 20516 2648 20568
rect 2700 20516 2710 20568
rect 2642 20511 2708 20516
rect 2754 20459 2788 20599
rect 2834 20568 2900 20571
rect 2830 20516 2840 20568
rect 2892 20516 2902 20568
rect 2834 20511 2900 20516
rect 2946 20459 2980 20599
rect 3026 20568 3092 20571
rect 3022 20516 3032 20568
rect 3084 20516 3094 20568
rect 3026 20511 3092 20516
rect 3138 20459 3172 20599
rect 3218 20567 3284 20571
rect 3215 20515 3225 20567
rect 3277 20515 3287 20567
rect 3218 20511 3284 20515
rect 3330 20459 3364 20599
rect 3410 20567 3476 20571
rect 3407 20515 3417 20567
rect 3469 20515 3479 20567
rect 3534 20566 3580 20604
rect 3534 20532 3540 20566
rect 3574 20532 3580 20566
rect 3410 20511 3476 20515
rect 2282 20425 3364 20459
rect 3534 20349 3580 20532
rect 3803 20459 3837 20608
rect 3981 20668 4027 20703
rect 3981 20634 3987 20668
rect 4021 20634 4027 20668
rect 3981 20599 4027 20634
rect 4077 20668 4123 20703
rect 4077 20634 4083 20668
rect 4117 20634 4123 20668
rect 4077 20599 4123 20634
rect 4173 20668 4219 20703
rect 4173 20634 4179 20668
rect 4213 20634 4219 20668
rect 4173 20599 4219 20634
rect 4269 20668 4315 20703
rect 4269 20634 4275 20668
rect 4309 20634 4315 20668
rect 4269 20599 4315 20634
rect 4365 20668 4411 20703
rect 4365 20634 4371 20668
rect 4405 20634 4411 20668
rect 4365 20599 4411 20634
rect 4461 20668 4507 20703
rect 4461 20634 4467 20668
rect 4501 20634 4507 20668
rect 4461 20599 4507 20634
rect 4557 20668 4603 20703
rect 4557 20634 4563 20668
rect 4597 20634 4603 20668
rect 4557 20599 4603 20634
rect 4653 20668 4699 20703
rect 4653 20634 4659 20668
rect 4693 20634 4699 20668
rect 4653 20599 4699 20634
rect 4749 20668 4795 20703
rect 4749 20634 4755 20668
rect 4789 20634 4795 20668
rect 4749 20599 4795 20634
rect 4845 20668 4891 20703
rect 4845 20634 4851 20668
rect 4885 20634 4891 20668
rect 4845 20599 4891 20634
rect 4941 20668 4987 20703
rect 4941 20634 4947 20668
rect 4981 20634 4987 20668
rect 4941 20599 4987 20634
rect 5055 20676 5061 20710
rect 5095 20676 5101 20710
rect 5055 20638 5101 20676
rect 5055 20604 5061 20638
rect 5095 20621 5101 20638
rect 5095 20604 5550 20621
rect 3971 20568 4037 20571
rect 3968 20516 3978 20568
rect 4030 20516 4040 20568
rect 3971 20511 4037 20516
rect 4083 20459 4117 20599
rect 4163 20568 4229 20571
rect 4159 20516 4169 20568
rect 4221 20516 4231 20568
rect 4163 20511 4229 20516
rect 4275 20459 4309 20599
rect 4355 20568 4421 20571
rect 4351 20516 4361 20568
rect 4413 20516 4423 20568
rect 4355 20511 4421 20516
rect 4467 20459 4501 20599
rect 4547 20568 4613 20571
rect 4543 20516 4553 20568
rect 4605 20516 4615 20568
rect 4547 20511 4613 20516
rect 4659 20459 4693 20599
rect 4739 20567 4805 20571
rect 4736 20515 4746 20567
rect 4798 20515 4808 20567
rect 4739 20511 4805 20515
rect 4851 20459 4885 20599
rect 5055 20590 5550 20604
rect 4931 20567 4997 20571
rect 4928 20515 4938 20567
rect 4990 20515 5000 20567
rect 5055 20566 5303 20590
rect 5055 20532 5061 20566
rect 5095 20556 5303 20566
rect 5337 20556 5395 20590
rect 5429 20556 5487 20590
rect 5521 20556 5550 20590
rect 5095 20532 5550 20556
rect 5055 20525 5550 20532
rect 4931 20511 4997 20515
rect 3803 20425 4885 20459
rect 5055 20350 5101 20525
rect 129 20142 1211 20176
rect 129 19579 163 20142
rect 294 20032 304 20084
rect 356 20032 366 20084
rect 409 19992 443 20142
rect 487 20032 497 20084
rect 549 20032 559 20084
rect 601 19992 635 20142
rect 678 20032 688 20084
rect 740 20032 750 20084
rect 793 19992 827 20142
rect 870 20032 880 20084
rect 932 20032 942 20084
rect 985 19992 1019 20142
rect 1062 20032 1072 20084
rect 1124 20032 1134 20084
rect 1177 19992 1211 20142
rect 1254 20032 1264 20084
rect 1316 20032 1326 20084
rect 1381 20048 1427 20212
rect 2282 20146 3364 20180
rect 1381 20014 1387 20048
rect 1421 20014 1427 20048
rect 1512 20025 1522 20085
rect 1578 20025 1792 20085
rect 1852 20025 1862 20085
rect 307 19945 353 19992
rect 307 19911 313 19945
rect 347 19911 353 19945
rect 307 19873 353 19911
rect 307 19839 313 19873
rect 347 19839 353 19873
rect 307 19801 353 19839
rect 307 19767 313 19801
rect 347 19767 353 19801
rect 307 19720 353 19767
rect 403 19945 449 19992
rect 403 19911 409 19945
rect 443 19911 449 19945
rect 403 19873 449 19911
rect 403 19839 409 19873
rect 443 19839 449 19873
rect 403 19801 449 19839
rect 403 19767 409 19801
rect 443 19767 449 19801
rect 403 19720 449 19767
rect 499 19945 545 19992
rect 499 19911 505 19945
rect 539 19911 545 19945
rect 499 19873 545 19911
rect 499 19839 505 19873
rect 539 19839 545 19873
rect 499 19801 545 19839
rect 499 19767 505 19801
rect 539 19767 545 19801
rect 499 19720 545 19767
rect 595 19945 641 19992
rect 595 19911 601 19945
rect 635 19911 641 19945
rect 595 19873 641 19911
rect 595 19839 601 19873
rect 635 19839 641 19873
rect 595 19801 641 19839
rect 595 19767 601 19801
rect 635 19767 641 19801
rect 595 19720 641 19767
rect 691 19945 737 19992
rect 691 19911 697 19945
rect 731 19911 737 19945
rect 691 19873 737 19911
rect 691 19839 697 19873
rect 731 19839 737 19873
rect 691 19801 737 19839
rect 691 19767 697 19801
rect 731 19767 737 19801
rect 691 19720 737 19767
rect 787 19945 833 19992
rect 787 19911 793 19945
rect 827 19911 833 19945
rect 787 19873 833 19911
rect 787 19839 793 19873
rect 827 19839 833 19873
rect 787 19801 833 19839
rect 787 19767 793 19801
rect 827 19767 833 19801
rect 787 19720 833 19767
rect 883 19945 929 19992
rect 883 19911 889 19945
rect 923 19911 929 19945
rect 883 19873 929 19911
rect 883 19839 889 19873
rect 923 19839 929 19873
rect 883 19801 929 19839
rect 883 19767 889 19801
rect 923 19767 929 19801
rect 883 19720 929 19767
rect 979 19945 1025 19992
rect 979 19911 985 19945
rect 1019 19911 1025 19945
rect 979 19873 1025 19911
rect 979 19839 985 19873
rect 1019 19839 1025 19873
rect 979 19801 1025 19839
rect 979 19767 985 19801
rect 1019 19767 1025 19801
rect 979 19720 1025 19767
rect 1075 19945 1121 19992
rect 1075 19911 1081 19945
rect 1115 19911 1121 19945
rect 1075 19873 1121 19911
rect 1075 19839 1081 19873
rect 1115 19839 1121 19873
rect 1075 19801 1121 19839
rect 1075 19767 1081 19801
rect 1115 19767 1121 19801
rect 1075 19720 1121 19767
rect 1171 19945 1217 19992
rect 1171 19911 1177 19945
rect 1211 19911 1217 19945
rect 1171 19873 1217 19911
rect 1171 19839 1177 19873
rect 1211 19839 1217 19873
rect 1171 19801 1217 19839
rect 1171 19767 1177 19801
rect 1211 19767 1217 19801
rect 1171 19720 1217 19767
rect 1267 19945 1313 19992
rect 1267 19911 1273 19945
rect 1307 19911 1313 19945
rect 1267 19873 1313 19911
rect 1267 19839 1273 19873
rect 1307 19839 1313 19873
rect 1267 19801 1313 19839
rect 1267 19767 1273 19801
rect 1307 19767 1313 19801
rect 1267 19720 1313 19767
rect 1381 19976 1427 20014
rect 1381 19942 1387 19976
rect 1421 19942 1427 19976
rect 1381 19904 1427 19942
rect 1381 19870 1387 19904
rect 1421 19870 1427 19904
rect 1381 19832 1427 19870
rect 1381 19798 1387 19832
rect 1421 19798 1427 19832
rect 1381 19788 1427 19798
rect 1381 19786 2160 19788
rect 1381 19760 2056 19786
rect 1381 19735 1387 19760
rect 1380 19726 1387 19735
rect 1421 19726 2056 19760
rect 0 19545 163 19579
rect 129 19168 163 19545
rect 313 19579 347 19720
rect 505 19579 539 19720
rect 697 19579 731 19720
rect 889 19579 923 19720
rect 1081 19579 1115 19720
rect 1273 19579 1307 19720
rect 1380 19678 2056 19726
rect 2190 19678 2200 19786
rect 1380 19676 2160 19678
rect 2282 19583 2316 20146
rect 2447 20036 2457 20088
rect 2509 20036 2519 20088
rect 2562 19996 2596 20146
rect 2640 20036 2650 20088
rect 2702 20036 2712 20088
rect 2754 19996 2788 20146
rect 2831 20036 2841 20088
rect 2893 20036 2903 20088
rect 2946 19996 2980 20146
rect 3023 20036 3033 20088
rect 3085 20036 3095 20088
rect 3138 19996 3172 20146
rect 3215 20036 3225 20088
rect 3277 20036 3287 20088
rect 3330 19996 3364 20146
rect 3407 20036 3417 20088
rect 3469 20036 3479 20088
rect 3534 20052 3580 20260
rect 3534 20018 3540 20052
rect 3574 20018 3580 20052
rect 2460 19949 2506 19996
rect 2460 19915 2466 19949
rect 2500 19915 2506 19949
rect 2460 19877 2506 19915
rect 2460 19843 2466 19877
rect 2500 19843 2506 19877
rect 2460 19805 2506 19843
rect 2460 19771 2466 19805
rect 2500 19771 2506 19805
rect 2460 19724 2506 19771
rect 2556 19949 2602 19996
rect 2556 19915 2562 19949
rect 2596 19915 2602 19949
rect 2556 19877 2602 19915
rect 2556 19843 2562 19877
rect 2596 19843 2602 19877
rect 2556 19805 2602 19843
rect 2556 19771 2562 19805
rect 2596 19771 2602 19805
rect 2556 19724 2602 19771
rect 2652 19949 2698 19996
rect 2652 19915 2658 19949
rect 2692 19915 2698 19949
rect 2652 19877 2698 19915
rect 2652 19843 2658 19877
rect 2692 19843 2698 19877
rect 2652 19805 2698 19843
rect 2652 19771 2658 19805
rect 2692 19771 2698 19805
rect 2652 19724 2698 19771
rect 2748 19949 2794 19996
rect 2748 19915 2754 19949
rect 2788 19915 2794 19949
rect 2748 19877 2794 19915
rect 2748 19843 2754 19877
rect 2788 19843 2794 19877
rect 2748 19805 2794 19843
rect 2748 19771 2754 19805
rect 2788 19771 2794 19805
rect 2748 19724 2794 19771
rect 2844 19949 2890 19996
rect 2844 19915 2850 19949
rect 2884 19915 2890 19949
rect 2844 19877 2890 19915
rect 2844 19843 2850 19877
rect 2884 19843 2890 19877
rect 2844 19805 2890 19843
rect 2844 19771 2850 19805
rect 2884 19771 2890 19805
rect 2844 19724 2890 19771
rect 2940 19949 2986 19996
rect 2940 19915 2946 19949
rect 2980 19915 2986 19949
rect 2940 19877 2986 19915
rect 2940 19843 2946 19877
rect 2980 19843 2986 19877
rect 2940 19805 2986 19843
rect 2940 19771 2946 19805
rect 2980 19771 2986 19805
rect 2940 19724 2986 19771
rect 3036 19949 3082 19996
rect 3036 19915 3042 19949
rect 3076 19915 3082 19949
rect 3036 19877 3082 19915
rect 3036 19843 3042 19877
rect 3076 19843 3082 19877
rect 3036 19805 3082 19843
rect 3036 19771 3042 19805
rect 3076 19771 3082 19805
rect 3036 19724 3082 19771
rect 3132 19949 3178 19996
rect 3132 19915 3138 19949
rect 3172 19915 3178 19949
rect 3132 19877 3178 19915
rect 3132 19843 3138 19877
rect 3172 19843 3178 19877
rect 3132 19805 3178 19843
rect 3132 19771 3138 19805
rect 3172 19771 3178 19805
rect 3132 19724 3178 19771
rect 3228 19949 3274 19996
rect 3228 19915 3234 19949
rect 3268 19915 3274 19949
rect 3228 19877 3274 19915
rect 3228 19843 3234 19877
rect 3268 19843 3274 19877
rect 3228 19805 3274 19843
rect 3228 19771 3234 19805
rect 3268 19771 3274 19805
rect 3228 19724 3274 19771
rect 3324 19949 3370 19996
rect 3324 19915 3330 19949
rect 3364 19915 3370 19949
rect 3324 19877 3370 19915
rect 3324 19843 3330 19877
rect 3364 19843 3370 19877
rect 3324 19805 3370 19843
rect 3324 19771 3330 19805
rect 3364 19771 3370 19805
rect 3324 19724 3370 19771
rect 3420 19949 3466 19996
rect 3420 19915 3426 19949
rect 3460 19915 3466 19949
rect 3420 19877 3466 19915
rect 3420 19843 3426 19877
rect 3460 19843 3466 19877
rect 3420 19805 3466 19843
rect 3420 19771 3426 19805
rect 3460 19771 3466 19805
rect 3420 19724 3466 19771
rect 3534 19980 3580 20018
rect 3534 19946 3540 19980
rect 3574 19946 3580 19980
rect 3534 19908 3580 19946
rect 3534 19874 3540 19908
rect 3574 19874 3580 19908
rect 3534 19836 3580 19874
rect 3534 19802 3540 19836
rect 3574 19802 3580 19836
rect 3534 19764 3580 19802
rect 3534 19730 3540 19764
rect 3574 19730 3580 19764
rect 2101 19579 2316 19583
rect 313 19549 2316 19579
rect 313 19545 2141 19549
rect 313 19412 347 19545
rect 505 19412 539 19545
rect 697 19412 731 19545
rect 889 19412 923 19545
rect 1081 19412 1115 19545
rect 1273 19412 1307 19545
rect 1381 19419 1608 19442
rect 307 19377 353 19412
rect 307 19343 313 19377
rect 347 19343 353 19377
rect 307 19308 353 19343
rect 403 19377 449 19412
rect 403 19343 409 19377
rect 443 19343 449 19377
rect 403 19308 449 19343
rect 499 19377 545 19412
rect 499 19343 505 19377
rect 539 19343 545 19377
rect 499 19308 545 19343
rect 595 19377 641 19412
rect 595 19343 601 19377
rect 635 19343 641 19377
rect 595 19308 641 19343
rect 691 19377 737 19412
rect 691 19343 697 19377
rect 731 19343 737 19377
rect 691 19308 737 19343
rect 787 19377 833 19412
rect 787 19343 793 19377
rect 827 19343 833 19377
rect 787 19308 833 19343
rect 883 19377 929 19412
rect 883 19343 889 19377
rect 923 19343 929 19377
rect 883 19308 929 19343
rect 979 19377 1025 19412
rect 979 19343 985 19377
rect 1019 19343 1025 19377
rect 979 19308 1025 19343
rect 1075 19377 1121 19412
rect 1075 19343 1081 19377
rect 1115 19343 1121 19377
rect 1075 19308 1121 19343
rect 1171 19377 1217 19412
rect 1171 19343 1177 19377
rect 1211 19343 1217 19377
rect 1171 19308 1217 19343
rect 1267 19377 1313 19412
rect 1267 19343 1273 19377
rect 1307 19343 1313 19377
rect 1267 19308 1313 19343
rect 1381 19385 1387 19419
rect 1421 19385 1608 19419
rect 1381 19347 1608 19385
rect 1381 19313 1387 19347
rect 1421 19322 1608 19347
rect 1421 19313 1427 19322
rect 1560 19320 1608 19322
rect 1598 19318 1608 19320
rect 1720 19318 1730 19442
rect 297 19277 363 19280
rect 294 19225 304 19277
rect 356 19225 366 19277
rect 297 19220 363 19225
rect 409 19168 443 19308
rect 489 19277 555 19280
rect 485 19225 495 19277
rect 547 19225 557 19277
rect 489 19220 555 19225
rect 601 19168 635 19308
rect 681 19277 747 19280
rect 677 19225 687 19277
rect 739 19225 749 19277
rect 681 19220 747 19225
rect 793 19168 827 19308
rect 873 19277 939 19280
rect 869 19225 879 19277
rect 931 19225 941 19277
rect 873 19220 939 19225
rect 985 19168 1019 19308
rect 1065 19276 1131 19280
rect 1062 19224 1072 19276
rect 1124 19224 1134 19276
rect 1065 19220 1131 19224
rect 1177 19168 1211 19308
rect 1257 19276 1323 19280
rect 1254 19224 1264 19276
rect 1316 19224 1326 19276
rect 1381 19275 1427 19313
rect 1920 19280 1930 19282
rect 1381 19241 1387 19275
rect 1421 19241 1427 19275
rect 1257 19220 1323 19224
rect 129 19134 1211 19168
rect 1381 19098 1427 19241
rect 1458 19224 1468 19280
rect 1524 19226 1930 19280
rect 1986 19226 1996 19282
rect 1524 19224 1986 19226
rect 2282 19172 2316 19549
rect 2466 19583 2500 19724
rect 2658 19583 2692 19724
rect 2850 19583 2884 19724
rect 3042 19583 3076 19724
rect 3234 19583 3268 19724
rect 3426 19583 3460 19724
rect 3534 19686 3580 19730
rect 3803 20146 4885 20180
rect 3803 19583 3837 20146
rect 3968 20036 3978 20088
rect 4030 20036 4040 20088
rect 4083 19996 4117 20146
rect 4161 20036 4171 20088
rect 4223 20036 4233 20088
rect 4275 19996 4309 20146
rect 4352 20036 4362 20088
rect 4414 20036 4424 20088
rect 4467 19996 4501 20146
rect 4544 20036 4554 20088
rect 4606 20036 4616 20088
rect 4659 19996 4693 20146
rect 4736 20036 4746 20088
rect 4798 20036 4808 20088
rect 4851 19996 4885 20146
rect 4928 20036 4938 20088
rect 4990 20036 5000 20088
rect 5055 20052 5101 20257
rect 5055 20018 5061 20052
rect 5095 20018 5101 20052
rect 3981 19949 4027 19996
rect 3981 19915 3987 19949
rect 4021 19915 4027 19949
rect 3981 19877 4027 19915
rect 3981 19843 3987 19877
rect 4021 19843 4027 19877
rect 3981 19805 4027 19843
rect 3981 19771 3987 19805
rect 4021 19771 4027 19805
rect 3981 19724 4027 19771
rect 4077 19949 4123 19996
rect 4077 19915 4083 19949
rect 4117 19915 4123 19949
rect 4077 19877 4123 19915
rect 4077 19843 4083 19877
rect 4117 19843 4123 19877
rect 4077 19805 4123 19843
rect 4077 19771 4083 19805
rect 4117 19771 4123 19805
rect 4077 19724 4123 19771
rect 4173 19949 4219 19996
rect 4173 19915 4179 19949
rect 4213 19915 4219 19949
rect 4173 19877 4219 19915
rect 4173 19843 4179 19877
rect 4213 19843 4219 19877
rect 4173 19805 4219 19843
rect 4173 19771 4179 19805
rect 4213 19771 4219 19805
rect 4173 19724 4219 19771
rect 4269 19949 4315 19996
rect 4269 19915 4275 19949
rect 4309 19915 4315 19949
rect 4269 19877 4315 19915
rect 4269 19843 4275 19877
rect 4309 19843 4315 19877
rect 4269 19805 4315 19843
rect 4269 19771 4275 19805
rect 4309 19771 4315 19805
rect 4269 19724 4315 19771
rect 4365 19949 4411 19996
rect 4365 19915 4371 19949
rect 4405 19915 4411 19949
rect 4365 19877 4411 19915
rect 4365 19843 4371 19877
rect 4405 19843 4411 19877
rect 4365 19805 4411 19843
rect 4365 19771 4371 19805
rect 4405 19771 4411 19805
rect 4365 19724 4411 19771
rect 4461 19949 4507 19996
rect 4461 19915 4467 19949
rect 4501 19915 4507 19949
rect 4461 19877 4507 19915
rect 4461 19843 4467 19877
rect 4501 19843 4507 19877
rect 4461 19805 4507 19843
rect 4461 19771 4467 19805
rect 4501 19771 4507 19805
rect 4461 19724 4507 19771
rect 4557 19949 4603 19996
rect 4557 19915 4563 19949
rect 4597 19915 4603 19949
rect 4557 19877 4603 19915
rect 4557 19843 4563 19877
rect 4597 19843 4603 19877
rect 4557 19805 4603 19843
rect 4557 19771 4563 19805
rect 4597 19771 4603 19805
rect 4557 19724 4603 19771
rect 4653 19949 4699 19996
rect 4653 19915 4659 19949
rect 4693 19915 4699 19949
rect 4653 19877 4699 19915
rect 4653 19843 4659 19877
rect 4693 19843 4699 19877
rect 4653 19805 4699 19843
rect 4653 19771 4659 19805
rect 4693 19771 4699 19805
rect 4653 19724 4699 19771
rect 4749 19949 4795 19996
rect 4749 19915 4755 19949
rect 4789 19915 4795 19949
rect 4749 19877 4795 19915
rect 4749 19843 4755 19877
rect 4789 19843 4795 19877
rect 4749 19805 4795 19843
rect 4749 19771 4755 19805
rect 4789 19771 4795 19805
rect 4749 19724 4795 19771
rect 4845 19949 4891 19996
rect 4845 19915 4851 19949
rect 4885 19915 4891 19949
rect 4845 19877 4891 19915
rect 4845 19843 4851 19877
rect 4885 19843 4891 19877
rect 4845 19805 4891 19843
rect 4845 19771 4851 19805
rect 4885 19771 4891 19805
rect 4845 19724 4891 19771
rect 4941 19949 4987 19996
rect 4941 19915 4947 19949
rect 4981 19915 4987 19949
rect 4941 19877 4987 19915
rect 4941 19843 4947 19877
rect 4981 19843 4987 19877
rect 4941 19805 4987 19843
rect 4941 19771 4947 19805
rect 4981 19771 4987 19805
rect 4941 19724 4987 19771
rect 5055 19980 5101 20018
rect 5055 19946 5061 19980
rect 5095 19946 5101 19980
rect 5055 19908 5101 19946
rect 5055 19874 5061 19908
rect 5095 19877 5101 19908
rect 5274 19877 5550 19878
rect 5095 19874 5550 19877
rect 5055 19847 5550 19874
rect 5055 19836 5303 19847
rect 5055 19802 5061 19836
rect 5095 19813 5303 19836
rect 5337 19813 5395 19847
rect 5429 19813 5487 19847
rect 5521 19813 5550 19847
rect 5095 19802 5550 19813
rect 5055 19782 5550 19802
rect 5055 19764 5101 19782
rect 5055 19730 5061 19764
rect 5095 19730 5101 19764
rect 2466 19549 3837 19583
rect 2466 19416 2500 19549
rect 2658 19416 2692 19549
rect 2850 19416 2884 19549
rect 3042 19416 3076 19549
rect 3234 19416 3268 19549
rect 3426 19416 3460 19549
rect 3671 19459 3681 19511
rect 3733 19459 3743 19511
rect 3679 19458 3691 19459
rect 3725 19458 3737 19459
rect 3679 19452 3737 19458
rect 3534 19423 3580 19446
rect 2460 19381 2506 19416
rect 2460 19347 2466 19381
rect 2500 19347 2506 19381
rect 2460 19312 2506 19347
rect 2556 19381 2602 19416
rect 2556 19347 2562 19381
rect 2596 19347 2602 19381
rect 2556 19312 2602 19347
rect 2652 19381 2698 19416
rect 2652 19347 2658 19381
rect 2692 19347 2698 19381
rect 2652 19312 2698 19347
rect 2748 19381 2794 19416
rect 2748 19347 2754 19381
rect 2788 19347 2794 19381
rect 2748 19312 2794 19347
rect 2844 19381 2890 19416
rect 2844 19347 2850 19381
rect 2884 19347 2890 19381
rect 2844 19312 2890 19347
rect 2940 19381 2986 19416
rect 2940 19347 2946 19381
rect 2980 19347 2986 19381
rect 2940 19312 2986 19347
rect 3036 19381 3082 19416
rect 3036 19347 3042 19381
rect 3076 19347 3082 19381
rect 3036 19312 3082 19347
rect 3132 19381 3178 19416
rect 3132 19347 3138 19381
rect 3172 19347 3178 19381
rect 3132 19312 3178 19347
rect 3228 19381 3274 19416
rect 3228 19347 3234 19381
rect 3268 19347 3274 19381
rect 3228 19312 3274 19347
rect 3324 19381 3370 19416
rect 3324 19347 3330 19381
rect 3364 19347 3370 19381
rect 3324 19312 3370 19347
rect 3420 19381 3466 19416
rect 3420 19347 3426 19381
rect 3460 19347 3466 19381
rect 3420 19312 3466 19347
rect 3534 19389 3540 19423
rect 3574 19421 3580 19423
rect 3803 19421 3837 19549
rect 3574 19420 3680 19421
rect 3734 19420 3837 19421
rect 3574 19408 3687 19420
rect 3574 19389 3647 19408
rect 3534 19351 3647 19389
rect 3534 19317 3540 19351
rect 3574 19332 3647 19351
rect 3681 19332 3687 19408
rect 3574 19321 3687 19332
rect 3574 19317 3580 19321
rect 3641 19320 3687 19321
rect 3729 19408 3837 19420
rect 3987 19583 4021 19724
rect 4179 19583 4213 19724
rect 4371 19583 4405 19724
rect 4563 19583 4597 19724
rect 4755 19583 4789 19724
rect 4947 19583 4981 19724
rect 5055 19686 5101 19730
rect 5683 19637 5743 20890
rect 5177 19603 5743 19637
rect 5177 19583 5211 19603
rect 3987 19549 5211 19583
rect 3987 19416 4021 19549
rect 4179 19416 4213 19549
rect 4371 19416 4405 19549
rect 4563 19416 4597 19549
rect 4755 19416 4789 19549
rect 4947 19416 4981 19549
rect 5438 19545 5512 19546
rect 5326 19543 5400 19544
rect 5326 19491 5337 19543
rect 5389 19491 5400 19543
rect 5438 19493 5449 19545
rect 5501 19493 5512 19545
rect 5438 19492 5512 19493
rect 5326 19490 5400 19491
rect 5055 19423 5101 19446
rect 3729 19332 3735 19408
rect 3769 19332 3837 19408
rect 3729 19321 3837 19332
rect 3729 19320 3775 19321
rect 2450 19281 2516 19284
rect 2447 19229 2457 19281
rect 2509 19229 2519 19281
rect 2450 19224 2516 19229
rect 2562 19172 2596 19312
rect 2642 19281 2708 19284
rect 2638 19229 2648 19281
rect 2700 19229 2710 19281
rect 2642 19224 2708 19229
rect 2754 19172 2788 19312
rect 2834 19281 2900 19284
rect 2830 19229 2840 19281
rect 2892 19229 2902 19281
rect 2834 19224 2900 19229
rect 2946 19172 2980 19312
rect 3026 19281 3092 19284
rect 3022 19229 3032 19281
rect 3084 19229 3094 19281
rect 3026 19224 3092 19229
rect 3138 19172 3172 19312
rect 3218 19280 3284 19284
rect 3215 19228 3225 19280
rect 3277 19228 3287 19280
rect 3218 19224 3284 19228
rect 3330 19172 3364 19312
rect 3410 19280 3476 19284
rect 3407 19228 3417 19280
rect 3469 19228 3479 19280
rect 3534 19279 3580 19317
rect 3534 19245 3540 19279
rect 3574 19245 3580 19279
rect 3410 19224 3476 19228
rect 2282 19138 3364 19172
rect 3534 19062 3580 19245
rect 3803 19172 3837 19321
rect 3981 19381 4027 19416
rect 3981 19347 3987 19381
rect 4021 19347 4027 19381
rect 3981 19312 4027 19347
rect 4077 19381 4123 19416
rect 4077 19347 4083 19381
rect 4117 19347 4123 19381
rect 4077 19312 4123 19347
rect 4173 19381 4219 19416
rect 4173 19347 4179 19381
rect 4213 19347 4219 19381
rect 4173 19312 4219 19347
rect 4269 19381 4315 19416
rect 4269 19347 4275 19381
rect 4309 19347 4315 19381
rect 4269 19312 4315 19347
rect 4365 19381 4411 19416
rect 4365 19347 4371 19381
rect 4405 19347 4411 19381
rect 4365 19312 4411 19347
rect 4461 19381 4507 19416
rect 4461 19347 4467 19381
rect 4501 19347 4507 19381
rect 4461 19312 4507 19347
rect 4557 19381 4603 19416
rect 4557 19347 4563 19381
rect 4597 19347 4603 19381
rect 4557 19312 4603 19347
rect 4653 19381 4699 19416
rect 4653 19347 4659 19381
rect 4693 19347 4699 19381
rect 4653 19312 4699 19347
rect 4749 19381 4795 19416
rect 4749 19347 4755 19381
rect 4789 19347 4795 19381
rect 4749 19312 4795 19347
rect 4845 19381 4891 19416
rect 4845 19347 4851 19381
rect 4885 19347 4891 19381
rect 4845 19312 4891 19347
rect 4941 19381 4987 19416
rect 4941 19347 4947 19381
rect 4981 19347 4987 19381
rect 4941 19312 4987 19347
rect 5055 19389 5061 19423
rect 5095 19389 5101 19423
rect 5055 19351 5101 19389
rect 5055 19317 5061 19351
rect 5095 19334 5101 19351
rect 5095 19317 5550 19334
rect 3971 19281 4037 19284
rect 3968 19229 3978 19281
rect 4030 19229 4040 19281
rect 3971 19224 4037 19229
rect 4083 19172 4117 19312
rect 4163 19281 4229 19284
rect 4159 19229 4169 19281
rect 4221 19229 4231 19281
rect 4163 19224 4229 19229
rect 4275 19172 4309 19312
rect 4355 19281 4421 19284
rect 4351 19229 4361 19281
rect 4413 19229 4423 19281
rect 4355 19224 4421 19229
rect 4467 19172 4501 19312
rect 4547 19281 4613 19284
rect 4543 19229 4553 19281
rect 4605 19229 4615 19281
rect 4547 19224 4613 19229
rect 4659 19172 4693 19312
rect 4739 19280 4805 19284
rect 4736 19228 4746 19280
rect 4798 19228 4808 19280
rect 4739 19224 4805 19228
rect 4851 19172 4885 19312
rect 5055 19303 5550 19317
rect 4931 19280 4997 19284
rect 4928 19228 4938 19280
rect 4990 19228 5000 19280
rect 5055 19279 5303 19303
rect 5055 19245 5061 19279
rect 5095 19269 5303 19279
rect 5337 19269 5395 19303
rect 5429 19269 5487 19303
rect 5521 19269 5550 19303
rect 5095 19245 5550 19269
rect 5055 19238 5550 19245
rect 4931 19224 4997 19228
rect 3803 19138 4885 19172
rect 5055 19063 5101 19238
rect 129 18855 1211 18889
rect 129 18292 163 18855
rect 294 18745 304 18797
rect 356 18745 366 18797
rect 409 18705 443 18855
rect 487 18745 497 18797
rect 549 18745 559 18797
rect 601 18705 635 18855
rect 678 18745 688 18797
rect 740 18745 750 18797
rect 793 18705 827 18855
rect 870 18745 880 18797
rect 932 18745 942 18797
rect 985 18705 1019 18855
rect 1062 18745 1072 18797
rect 1124 18745 1134 18797
rect 1177 18705 1211 18855
rect 1254 18745 1264 18797
rect 1316 18745 1326 18797
rect 1381 18761 1427 18925
rect 2282 18859 3364 18893
rect 1381 18727 1387 18761
rect 1421 18727 1427 18761
rect 1512 18738 1522 18798
rect 1578 18738 1792 18798
rect 1852 18738 1862 18798
rect 307 18658 353 18705
rect 307 18624 313 18658
rect 347 18624 353 18658
rect 307 18586 353 18624
rect 307 18552 313 18586
rect 347 18552 353 18586
rect 307 18514 353 18552
rect 307 18480 313 18514
rect 347 18480 353 18514
rect 307 18433 353 18480
rect 403 18658 449 18705
rect 403 18624 409 18658
rect 443 18624 449 18658
rect 403 18586 449 18624
rect 403 18552 409 18586
rect 443 18552 449 18586
rect 403 18514 449 18552
rect 403 18480 409 18514
rect 443 18480 449 18514
rect 403 18433 449 18480
rect 499 18658 545 18705
rect 499 18624 505 18658
rect 539 18624 545 18658
rect 499 18586 545 18624
rect 499 18552 505 18586
rect 539 18552 545 18586
rect 499 18514 545 18552
rect 499 18480 505 18514
rect 539 18480 545 18514
rect 499 18433 545 18480
rect 595 18658 641 18705
rect 595 18624 601 18658
rect 635 18624 641 18658
rect 595 18586 641 18624
rect 595 18552 601 18586
rect 635 18552 641 18586
rect 595 18514 641 18552
rect 595 18480 601 18514
rect 635 18480 641 18514
rect 595 18433 641 18480
rect 691 18658 737 18705
rect 691 18624 697 18658
rect 731 18624 737 18658
rect 691 18586 737 18624
rect 691 18552 697 18586
rect 731 18552 737 18586
rect 691 18514 737 18552
rect 691 18480 697 18514
rect 731 18480 737 18514
rect 691 18433 737 18480
rect 787 18658 833 18705
rect 787 18624 793 18658
rect 827 18624 833 18658
rect 787 18586 833 18624
rect 787 18552 793 18586
rect 827 18552 833 18586
rect 787 18514 833 18552
rect 787 18480 793 18514
rect 827 18480 833 18514
rect 787 18433 833 18480
rect 883 18658 929 18705
rect 883 18624 889 18658
rect 923 18624 929 18658
rect 883 18586 929 18624
rect 883 18552 889 18586
rect 923 18552 929 18586
rect 883 18514 929 18552
rect 883 18480 889 18514
rect 923 18480 929 18514
rect 883 18433 929 18480
rect 979 18658 1025 18705
rect 979 18624 985 18658
rect 1019 18624 1025 18658
rect 979 18586 1025 18624
rect 979 18552 985 18586
rect 1019 18552 1025 18586
rect 979 18514 1025 18552
rect 979 18480 985 18514
rect 1019 18480 1025 18514
rect 979 18433 1025 18480
rect 1075 18658 1121 18705
rect 1075 18624 1081 18658
rect 1115 18624 1121 18658
rect 1075 18586 1121 18624
rect 1075 18552 1081 18586
rect 1115 18552 1121 18586
rect 1075 18514 1121 18552
rect 1075 18480 1081 18514
rect 1115 18480 1121 18514
rect 1075 18433 1121 18480
rect 1171 18658 1217 18705
rect 1171 18624 1177 18658
rect 1211 18624 1217 18658
rect 1171 18586 1217 18624
rect 1171 18552 1177 18586
rect 1211 18552 1217 18586
rect 1171 18514 1217 18552
rect 1171 18480 1177 18514
rect 1211 18480 1217 18514
rect 1171 18433 1217 18480
rect 1267 18658 1313 18705
rect 1267 18624 1273 18658
rect 1307 18624 1313 18658
rect 1267 18586 1313 18624
rect 1267 18552 1273 18586
rect 1307 18552 1313 18586
rect 1267 18514 1313 18552
rect 1267 18480 1273 18514
rect 1307 18480 1313 18514
rect 1267 18433 1313 18480
rect 1381 18689 1427 18727
rect 1381 18655 1387 18689
rect 1421 18655 1427 18689
rect 1381 18617 1427 18655
rect 1381 18583 1387 18617
rect 1421 18583 1427 18617
rect 1381 18545 1427 18583
rect 1381 18511 1387 18545
rect 1421 18511 1427 18545
rect 1381 18501 1427 18511
rect 1381 18499 2160 18501
rect 1381 18473 2056 18499
rect 1381 18448 1387 18473
rect 1380 18439 1387 18448
rect 1421 18439 2056 18473
rect 0 18258 163 18292
rect 129 17881 163 18258
rect 313 18292 347 18433
rect 505 18292 539 18433
rect 697 18292 731 18433
rect 889 18292 923 18433
rect 1081 18292 1115 18433
rect 1273 18292 1307 18433
rect 1380 18391 2056 18439
rect 2190 18391 2200 18499
rect 1380 18389 2160 18391
rect 2282 18296 2316 18859
rect 2447 18749 2457 18801
rect 2509 18749 2519 18801
rect 2562 18709 2596 18859
rect 2640 18749 2650 18801
rect 2702 18749 2712 18801
rect 2754 18709 2788 18859
rect 2831 18749 2841 18801
rect 2893 18749 2903 18801
rect 2946 18709 2980 18859
rect 3023 18749 3033 18801
rect 3085 18749 3095 18801
rect 3138 18709 3172 18859
rect 3215 18749 3225 18801
rect 3277 18749 3287 18801
rect 3330 18709 3364 18859
rect 3407 18749 3417 18801
rect 3469 18749 3479 18801
rect 3534 18765 3580 18973
rect 3534 18731 3540 18765
rect 3574 18731 3580 18765
rect 2460 18662 2506 18709
rect 2460 18628 2466 18662
rect 2500 18628 2506 18662
rect 2460 18590 2506 18628
rect 2460 18556 2466 18590
rect 2500 18556 2506 18590
rect 2460 18518 2506 18556
rect 2460 18484 2466 18518
rect 2500 18484 2506 18518
rect 2460 18437 2506 18484
rect 2556 18662 2602 18709
rect 2556 18628 2562 18662
rect 2596 18628 2602 18662
rect 2556 18590 2602 18628
rect 2556 18556 2562 18590
rect 2596 18556 2602 18590
rect 2556 18518 2602 18556
rect 2556 18484 2562 18518
rect 2596 18484 2602 18518
rect 2556 18437 2602 18484
rect 2652 18662 2698 18709
rect 2652 18628 2658 18662
rect 2692 18628 2698 18662
rect 2652 18590 2698 18628
rect 2652 18556 2658 18590
rect 2692 18556 2698 18590
rect 2652 18518 2698 18556
rect 2652 18484 2658 18518
rect 2692 18484 2698 18518
rect 2652 18437 2698 18484
rect 2748 18662 2794 18709
rect 2748 18628 2754 18662
rect 2788 18628 2794 18662
rect 2748 18590 2794 18628
rect 2748 18556 2754 18590
rect 2788 18556 2794 18590
rect 2748 18518 2794 18556
rect 2748 18484 2754 18518
rect 2788 18484 2794 18518
rect 2748 18437 2794 18484
rect 2844 18662 2890 18709
rect 2844 18628 2850 18662
rect 2884 18628 2890 18662
rect 2844 18590 2890 18628
rect 2844 18556 2850 18590
rect 2884 18556 2890 18590
rect 2844 18518 2890 18556
rect 2844 18484 2850 18518
rect 2884 18484 2890 18518
rect 2844 18437 2890 18484
rect 2940 18662 2986 18709
rect 2940 18628 2946 18662
rect 2980 18628 2986 18662
rect 2940 18590 2986 18628
rect 2940 18556 2946 18590
rect 2980 18556 2986 18590
rect 2940 18518 2986 18556
rect 2940 18484 2946 18518
rect 2980 18484 2986 18518
rect 2940 18437 2986 18484
rect 3036 18662 3082 18709
rect 3036 18628 3042 18662
rect 3076 18628 3082 18662
rect 3036 18590 3082 18628
rect 3036 18556 3042 18590
rect 3076 18556 3082 18590
rect 3036 18518 3082 18556
rect 3036 18484 3042 18518
rect 3076 18484 3082 18518
rect 3036 18437 3082 18484
rect 3132 18662 3178 18709
rect 3132 18628 3138 18662
rect 3172 18628 3178 18662
rect 3132 18590 3178 18628
rect 3132 18556 3138 18590
rect 3172 18556 3178 18590
rect 3132 18518 3178 18556
rect 3132 18484 3138 18518
rect 3172 18484 3178 18518
rect 3132 18437 3178 18484
rect 3228 18662 3274 18709
rect 3228 18628 3234 18662
rect 3268 18628 3274 18662
rect 3228 18590 3274 18628
rect 3228 18556 3234 18590
rect 3268 18556 3274 18590
rect 3228 18518 3274 18556
rect 3228 18484 3234 18518
rect 3268 18484 3274 18518
rect 3228 18437 3274 18484
rect 3324 18662 3370 18709
rect 3324 18628 3330 18662
rect 3364 18628 3370 18662
rect 3324 18590 3370 18628
rect 3324 18556 3330 18590
rect 3364 18556 3370 18590
rect 3324 18518 3370 18556
rect 3324 18484 3330 18518
rect 3364 18484 3370 18518
rect 3324 18437 3370 18484
rect 3420 18662 3466 18709
rect 3420 18628 3426 18662
rect 3460 18628 3466 18662
rect 3420 18590 3466 18628
rect 3420 18556 3426 18590
rect 3460 18556 3466 18590
rect 3420 18518 3466 18556
rect 3420 18484 3426 18518
rect 3460 18484 3466 18518
rect 3420 18437 3466 18484
rect 3534 18693 3580 18731
rect 3534 18659 3540 18693
rect 3574 18659 3580 18693
rect 3534 18621 3580 18659
rect 3534 18587 3540 18621
rect 3574 18587 3580 18621
rect 3534 18549 3580 18587
rect 3534 18515 3540 18549
rect 3574 18515 3580 18549
rect 3534 18477 3580 18515
rect 3534 18443 3540 18477
rect 3574 18443 3580 18477
rect 2101 18292 2316 18296
rect 313 18262 2316 18292
rect 313 18258 2141 18262
rect 313 18125 347 18258
rect 505 18125 539 18258
rect 697 18125 731 18258
rect 889 18125 923 18258
rect 1081 18125 1115 18258
rect 1273 18125 1307 18258
rect 1381 18132 1608 18155
rect 307 18090 353 18125
rect 307 18056 313 18090
rect 347 18056 353 18090
rect 307 18021 353 18056
rect 403 18090 449 18125
rect 403 18056 409 18090
rect 443 18056 449 18090
rect 403 18021 449 18056
rect 499 18090 545 18125
rect 499 18056 505 18090
rect 539 18056 545 18090
rect 499 18021 545 18056
rect 595 18090 641 18125
rect 595 18056 601 18090
rect 635 18056 641 18090
rect 595 18021 641 18056
rect 691 18090 737 18125
rect 691 18056 697 18090
rect 731 18056 737 18090
rect 691 18021 737 18056
rect 787 18090 833 18125
rect 787 18056 793 18090
rect 827 18056 833 18090
rect 787 18021 833 18056
rect 883 18090 929 18125
rect 883 18056 889 18090
rect 923 18056 929 18090
rect 883 18021 929 18056
rect 979 18090 1025 18125
rect 979 18056 985 18090
rect 1019 18056 1025 18090
rect 979 18021 1025 18056
rect 1075 18090 1121 18125
rect 1075 18056 1081 18090
rect 1115 18056 1121 18090
rect 1075 18021 1121 18056
rect 1171 18090 1217 18125
rect 1171 18056 1177 18090
rect 1211 18056 1217 18090
rect 1171 18021 1217 18056
rect 1267 18090 1313 18125
rect 1267 18056 1273 18090
rect 1307 18056 1313 18090
rect 1267 18021 1313 18056
rect 1381 18098 1387 18132
rect 1421 18098 1608 18132
rect 1381 18060 1608 18098
rect 1381 18026 1387 18060
rect 1421 18035 1608 18060
rect 1421 18026 1427 18035
rect 1560 18033 1608 18035
rect 1598 18031 1608 18033
rect 1720 18031 1730 18155
rect 297 17990 363 17993
rect 294 17938 304 17990
rect 356 17938 366 17990
rect 297 17933 363 17938
rect 409 17881 443 18021
rect 489 17990 555 17993
rect 485 17938 495 17990
rect 547 17938 557 17990
rect 489 17933 555 17938
rect 601 17881 635 18021
rect 681 17990 747 17993
rect 677 17938 687 17990
rect 739 17938 749 17990
rect 681 17933 747 17938
rect 793 17881 827 18021
rect 873 17990 939 17993
rect 869 17938 879 17990
rect 931 17938 941 17990
rect 873 17933 939 17938
rect 985 17881 1019 18021
rect 1065 17989 1131 17993
rect 1062 17937 1072 17989
rect 1124 17937 1134 17989
rect 1065 17933 1131 17937
rect 1177 17881 1211 18021
rect 1257 17989 1323 17993
rect 1254 17937 1264 17989
rect 1316 17937 1326 17989
rect 1381 17988 1427 18026
rect 1920 17993 1930 17995
rect 1381 17954 1387 17988
rect 1421 17954 1427 17988
rect 1257 17933 1323 17937
rect 129 17847 1211 17881
rect 1381 17811 1427 17954
rect 1458 17937 1468 17993
rect 1524 17939 1930 17993
rect 1986 17939 1996 17995
rect 1524 17937 1986 17939
rect 2282 17885 2316 18262
rect 2466 18296 2500 18437
rect 2658 18296 2692 18437
rect 2850 18296 2884 18437
rect 3042 18296 3076 18437
rect 3234 18296 3268 18437
rect 3426 18296 3460 18437
rect 3534 18399 3580 18443
rect 3803 18859 4885 18893
rect 3803 18296 3837 18859
rect 3968 18749 3978 18801
rect 4030 18749 4040 18801
rect 4083 18709 4117 18859
rect 4161 18749 4171 18801
rect 4223 18749 4233 18801
rect 4275 18709 4309 18859
rect 4352 18749 4362 18801
rect 4414 18749 4424 18801
rect 4467 18709 4501 18859
rect 4544 18749 4554 18801
rect 4606 18749 4616 18801
rect 4659 18709 4693 18859
rect 4736 18749 4746 18801
rect 4798 18749 4808 18801
rect 4851 18709 4885 18859
rect 4928 18749 4938 18801
rect 4990 18749 5000 18801
rect 5055 18765 5101 18970
rect 5055 18731 5061 18765
rect 5095 18731 5101 18765
rect 3981 18662 4027 18709
rect 3981 18628 3987 18662
rect 4021 18628 4027 18662
rect 3981 18590 4027 18628
rect 3981 18556 3987 18590
rect 4021 18556 4027 18590
rect 3981 18518 4027 18556
rect 3981 18484 3987 18518
rect 4021 18484 4027 18518
rect 3981 18437 4027 18484
rect 4077 18662 4123 18709
rect 4077 18628 4083 18662
rect 4117 18628 4123 18662
rect 4077 18590 4123 18628
rect 4077 18556 4083 18590
rect 4117 18556 4123 18590
rect 4077 18518 4123 18556
rect 4077 18484 4083 18518
rect 4117 18484 4123 18518
rect 4077 18437 4123 18484
rect 4173 18662 4219 18709
rect 4173 18628 4179 18662
rect 4213 18628 4219 18662
rect 4173 18590 4219 18628
rect 4173 18556 4179 18590
rect 4213 18556 4219 18590
rect 4173 18518 4219 18556
rect 4173 18484 4179 18518
rect 4213 18484 4219 18518
rect 4173 18437 4219 18484
rect 4269 18662 4315 18709
rect 4269 18628 4275 18662
rect 4309 18628 4315 18662
rect 4269 18590 4315 18628
rect 4269 18556 4275 18590
rect 4309 18556 4315 18590
rect 4269 18518 4315 18556
rect 4269 18484 4275 18518
rect 4309 18484 4315 18518
rect 4269 18437 4315 18484
rect 4365 18662 4411 18709
rect 4365 18628 4371 18662
rect 4405 18628 4411 18662
rect 4365 18590 4411 18628
rect 4365 18556 4371 18590
rect 4405 18556 4411 18590
rect 4365 18518 4411 18556
rect 4365 18484 4371 18518
rect 4405 18484 4411 18518
rect 4365 18437 4411 18484
rect 4461 18662 4507 18709
rect 4461 18628 4467 18662
rect 4501 18628 4507 18662
rect 4461 18590 4507 18628
rect 4461 18556 4467 18590
rect 4501 18556 4507 18590
rect 4461 18518 4507 18556
rect 4461 18484 4467 18518
rect 4501 18484 4507 18518
rect 4461 18437 4507 18484
rect 4557 18662 4603 18709
rect 4557 18628 4563 18662
rect 4597 18628 4603 18662
rect 4557 18590 4603 18628
rect 4557 18556 4563 18590
rect 4597 18556 4603 18590
rect 4557 18518 4603 18556
rect 4557 18484 4563 18518
rect 4597 18484 4603 18518
rect 4557 18437 4603 18484
rect 4653 18662 4699 18709
rect 4653 18628 4659 18662
rect 4693 18628 4699 18662
rect 4653 18590 4699 18628
rect 4653 18556 4659 18590
rect 4693 18556 4699 18590
rect 4653 18518 4699 18556
rect 4653 18484 4659 18518
rect 4693 18484 4699 18518
rect 4653 18437 4699 18484
rect 4749 18662 4795 18709
rect 4749 18628 4755 18662
rect 4789 18628 4795 18662
rect 4749 18590 4795 18628
rect 4749 18556 4755 18590
rect 4789 18556 4795 18590
rect 4749 18518 4795 18556
rect 4749 18484 4755 18518
rect 4789 18484 4795 18518
rect 4749 18437 4795 18484
rect 4845 18662 4891 18709
rect 4845 18628 4851 18662
rect 4885 18628 4891 18662
rect 4845 18590 4891 18628
rect 4845 18556 4851 18590
rect 4885 18556 4891 18590
rect 4845 18518 4891 18556
rect 4845 18484 4851 18518
rect 4885 18484 4891 18518
rect 4845 18437 4891 18484
rect 4941 18662 4987 18709
rect 4941 18628 4947 18662
rect 4981 18628 4987 18662
rect 4941 18590 4987 18628
rect 4941 18556 4947 18590
rect 4981 18556 4987 18590
rect 4941 18518 4987 18556
rect 4941 18484 4947 18518
rect 4981 18484 4987 18518
rect 4941 18437 4987 18484
rect 5055 18693 5101 18731
rect 5055 18659 5061 18693
rect 5095 18659 5101 18693
rect 5055 18621 5101 18659
rect 5055 18587 5061 18621
rect 5095 18590 5101 18621
rect 5274 18590 5550 18591
rect 5095 18587 5550 18590
rect 5055 18560 5550 18587
rect 5055 18549 5303 18560
rect 5055 18515 5061 18549
rect 5095 18526 5303 18549
rect 5337 18526 5395 18560
rect 5429 18526 5487 18560
rect 5521 18526 5550 18560
rect 5095 18515 5550 18526
rect 5055 18495 5550 18515
rect 5055 18477 5101 18495
rect 5055 18443 5061 18477
rect 5095 18443 5101 18477
rect 2466 18262 3837 18296
rect 2466 18129 2500 18262
rect 2658 18129 2692 18262
rect 2850 18129 2884 18262
rect 3042 18129 3076 18262
rect 3234 18129 3268 18262
rect 3426 18129 3460 18262
rect 3671 18172 3681 18224
rect 3733 18172 3743 18224
rect 3679 18171 3691 18172
rect 3725 18171 3737 18172
rect 3679 18165 3737 18171
rect 3534 18136 3580 18159
rect 2460 18094 2506 18129
rect 2460 18060 2466 18094
rect 2500 18060 2506 18094
rect 2460 18025 2506 18060
rect 2556 18094 2602 18129
rect 2556 18060 2562 18094
rect 2596 18060 2602 18094
rect 2556 18025 2602 18060
rect 2652 18094 2698 18129
rect 2652 18060 2658 18094
rect 2692 18060 2698 18094
rect 2652 18025 2698 18060
rect 2748 18094 2794 18129
rect 2748 18060 2754 18094
rect 2788 18060 2794 18094
rect 2748 18025 2794 18060
rect 2844 18094 2890 18129
rect 2844 18060 2850 18094
rect 2884 18060 2890 18094
rect 2844 18025 2890 18060
rect 2940 18094 2986 18129
rect 2940 18060 2946 18094
rect 2980 18060 2986 18094
rect 2940 18025 2986 18060
rect 3036 18094 3082 18129
rect 3036 18060 3042 18094
rect 3076 18060 3082 18094
rect 3036 18025 3082 18060
rect 3132 18094 3178 18129
rect 3132 18060 3138 18094
rect 3172 18060 3178 18094
rect 3132 18025 3178 18060
rect 3228 18094 3274 18129
rect 3228 18060 3234 18094
rect 3268 18060 3274 18094
rect 3228 18025 3274 18060
rect 3324 18094 3370 18129
rect 3324 18060 3330 18094
rect 3364 18060 3370 18094
rect 3324 18025 3370 18060
rect 3420 18094 3466 18129
rect 3420 18060 3426 18094
rect 3460 18060 3466 18094
rect 3420 18025 3466 18060
rect 3534 18102 3540 18136
rect 3574 18134 3580 18136
rect 3803 18134 3837 18262
rect 3574 18133 3680 18134
rect 3734 18133 3837 18134
rect 3574 18121 3687 18133
rect 3574 18102 3647 18121
rect 3534 18064 3647 18102
rect 3534 18030 3540 18064
rect 3574 18045 3647 18064
rect 3681 18045 3687 18121
rect 3574 18034 3687 18045
rect 3574 18030 3580 18034
rect 3641 18033 3687 18034
rect 3729 18121 3837 18133
rect 3987 18296 4021 18437
rect 4179 18296 4213 18437
rect 4371 18296 4405 18437
rect 4563 18296 4597 18437
rect 4755 18296 4789 18437
rect 4947 18296 4981 18437
rect 5055 18399 5101 18443
rect 5683 18350 5743 19603
rect 5177 18316 5743 18350
rect 5177 18296 5211 18316
rect 3987 18262 5211 18296
rect 3987 18129 4021 18262
rect 4179 18129 4213 18262
rect 4371 18129 4405 18262
rect 4563 18129 4597 18262
rect 4755 18129 4789 18262
rect 4947 18129 4981 18262
rect 5438 18258 5512 18259
rect 5326 18256 5400 18257
rect 5326 18204 5337 18256
rect 5389 18204 5400 18256
rect 5438 18206 5449 18258
rect 5501 18206 5512 18258
rect 5438 18205 5512 18206
rect 5326 18203 5400 18204
rect 5055 18136 5101 18159
rect 3729 18045 3735 18121
rect 3769 18045 3837 18121
rect 3729 18034 3837 18045
rect 3729 18033 3775 18034
rect 2450 17994 2516 17997
rect 2447 17942 2457 17994
rect 2509 17942 2519 17994
rect 2450 17937 2516 17942
rect 2562 17885 2596 18025
rect 2642 17994 2708 17997
rect 2638 17942 2648 17994
rect 2700 17942 2710 17994
rect 2642 17937 2708 17942
rect 2754 17885 2788 18025
rect 2834 17994 2900 17997
rect 2830 17942 2840 17994
rect 2892 17942 2902 17994
rect 2834 17937 2900 17942
rect 2946 17885 2980 18025
rect 3026 17994 3092 17997
rect 3022 17942 3032 17994
rect 3084 17942 3094 17994
rect 3026 17937 3092 17942
rect 3138 17885 3172 18025
rect 3218 17993 3284 17997
rect 3215 17941 3225 17993
rect 3277 17941 3287 17993
rect 3218 17937 3284 17941
rect 3330 17885 3364 18025
rect 3410 17993 3476 17997
rect 3407 17941 3417 17993
rect 3469 17941 3479 17993
rect 3534 17992 3580 18030
rect 3534 17958 3540 17992
rect 3574 17958 3580 17992
rect 3410 17937 3476 17941
rect 2282 17851 3364 17885
rect 3534 17775 3580 17958
rect 3803 17885 3837 18034
rect 3981 18094 4027 18129
rect 3981 18060 3987 18094
rect 4021 18060 4027 18094
rect 3981 18025 4027 18060
rect 4077 18094 4123 18129
rect 4077 18060 4083 18094
rect 4117 18060 4123 18094
rect 4077 18025 4123 18060
rect 4173 18094 4219 18129
rect 4173 18060 4179 18094
rect 4213 18060 4219 18094
rect 4173 18025 4219 18060
rect 4269 18094 4315 18129
rect 4269 18060 4275 18094
rect 4309 18060 4315 18094
rect 4269 18025 4315 18060
rect 4365 18094 4411 18129
rect 4365 18060 4371 18094
rect 4405 18060 4411 18094
rect 4365 18025 4411 18060
rect 4461 18094 4507 18129
rect 4461 18060 4467 18094
rect 4501 18060 4507 18094
rect 4461 18025 4507 18060
rect 4557 18094 4603 18129
rect 4557 18060 4563 18094
rect 4597 18060 4603 18094
rect 4557 18025 4603 18060
rect 4653 18094 4699 18129
rect 4653 18060 4659 18094
rect 4693 18060 4699 18094
rect 4653 18025 4699 18060
rect 4749 18094 4795 18129
rect 4749 18060 4755 18094
rect 4789 18060 4795 18094
rect 4749 18025 4795 18060
rect 4845 18094 4891 18129
rect 4845 18060 4851 18094
rect 4885 18060 4891 18094
rect 4845 18025 4891 18060
rect 4941 18094 4987 18129
rect 4941 18060 4947 18094
rect 4981 18060 4987 18094
rect 4941 18025 4987 18060
rect 5055 18102 5061 18136
rect 5095 18102 5101 18136
rect 5055 18064 5101 18102
rect 5055 18030 5061 18064
rect 5095 18047 5101 18064
rect 5095 18030 5550 18047
rect 3971 17994 4037 17997
rect 3968 17942 3978 17994
rect 4030 17942 4040 17994
rect 3971 17937 4037 17942
rect 4083 17885 4117 18025
rect 4163 17994 4229 17997
rect 4159 17942 4169 17994
rect 4221 17942 4231 17994
rect 4163 17937 4229 17942
rect 4275 17885 4309 18025
rect 4355 17994 4421 17997
rect 4351 17942 4361 17994
rect 4413 17942 4423 17994
rect 4355 17937 4421 17942
rect 4467 17885 4501 18025
rect 4547 17994 4613 17997
rect 4543 17942 4553 17994
rect 4605 17942 4615 17994
rect 4547 17937 4613 17942
rect 4659 17885 4693 18025
rect 4739 17993 4805 17997
rect 4736 17941 4746 17993
rect 4798 17941 4808 17993
rect 4739 17937 4805 17941
rect 4851 17885 4885 18025
rect 5055 18016 5550 18030
rect 4931 17993 4997 17997
rect 4928 17941 4938 17993
rect 4990 17941 5000 17993
rect 5055 17992 5303 18016
rect 5055 17958 5061 17992
rect 5095 17982 5303 17992
rect 5337 17982 5395 18016
rect 5429 17982 5487 18016
rect 5521 17982 5550 18016
rect 5095 17958 5550 17982
rect 5055 17951 5550 17958
rect 4931 17937 4997 17941
rect 3803 17851 4885 17885
rect 5055 17776 5101 17951
rect 129 17568 1211 17602
rect 129 17005 163 17568
rect 294 17458 304 17510
rect 356 17458 366 17510
rect 409 17418 443 17568
rect 487 17458 497 17510
rect 549 17458 559 17510
rect 601 17418 635 17568
rect 678 17458 688 17510
rect 740 17458 750 17510
rect 793 17418 827 17568
rect 870 17458 880 17510
rect 932 17458 942 17510
rect 985 17418 1019 17568
rect 1062 17458 1072 17510
rect 1124 17458 1134 17510
rect 1177 17418 1211 17568
rect 1254 17458 1264 17510
rect 1316 17458 1326 17510
rect 1381 17474 1427 17638
rect 2282 17572 3364 17606
rect 1381 17440 1387 17474
rect 1421 17440 1427 17474
rect 1512 17451 1522 17511
rect 1578 17451 1792 17511
rect 1852 17451 1862 17511
rect 307 17371 353 17418
rect 307 17337 313 17371
rect 347 17337 353 17371
rect 307 17299 353 17337
rect 307 17265 313 17299
rect 347 17265 353 17299
rect 307 17227 353 17265
rect 307 17193 313 17227
rect 347 17193 353 17227
rect 307 17146 353 17193
rect 403 17371 449 17418
rect 403 17337 409 17371
rect 443 17337 449 17371
rect 403 17299 449 17337
rect 403 17265 409 17299
rect 443 17265 449 17299
rect 403 17227 449 17265
rect 403 17193 409 17227
rect 443 17193 449 17227
rect 403 17146 449 17193
rect 499 17371 545 17418
rect 499 17337 505 17371
rect 539 17337 545 17371
rect 499 17299 545 17337
rect 499 17265 505 17299
rect 539 17265 545 17299
rect 499 17227 545 17265
rect 499 17193 505 17227
rect 539 17193 545 17227
rect 499 17146 545 17193
rect 595 17371 641 17418
rect 595 17337 601 17371
rect 635 17337 641 17371
rect 595 17299 641 17337
rect 595 17265 601 17299
rect 635 17265 641 17299
rect 595 17227 641 17265
rect 595 17193 601 17227
rect 635 17193 641 17227
rect 595 17146 641 17193
rect 691 17371 737 17418
rect 691 17337 697 17371
rect 731 17337 737 17371
rect 691 17299 737 17337
rect 691 17265 697 17299
rect 731 17265 737 17299
rect 691 17227 737 17265
rect 691 17193 697 17227
rect 731 17193 737 17227
rect 691 17146 737 17193
rect 787 17371 833 17418
rect 787 17337 793 17371
rect 827 17337 833 17371
rect 787 17299 833 17337
rect 787 17265 793 17299
rect 827 17265 833 17299
rect 787 17227 833 17265
rect 787 17193 793 17227
rect 827 17193 833 17227
rect 787 17146 833 17193
rect 883 17371 929 17418
rect 883 17337 889 17371
rect 923 17337 929 17371
rect 883 17299 929 17337
rect 883 17265 889 17299
rect 923 17265 929 17299
rect 883 17227 929 17265
rect 883 17193 889 17227
rect 923 17193 929 17227
rect 883 17146 929 17193
rect 979 17371 1025 17418
rect 979 17337 985 17371
rect 1019 17337 1025 17371
rect 979 17299 1025 17337
rect 979 17265 985 17299
rect 1019 17265 1025 17299
rect 979 17227 1025 17265
rect 979 17193 985 17227
rect 1019 17193 1025 17227
rect 979 17146 1025 17193
rect 1075 17371 1121 17418
rect 1075 17337 1081 17371
rect 1115 17337 1121 17371
rect 1075 17299 1121 17337
rect 1075 17265 1081 17299
rect 1115 17265 1121 17299
rect 1075 17227 1121 17265
rect 1075 17193 1081 17227
rect 1115 17193 1121 17227
rect 1075 17146 1121 17193
rect 1171 17371 1217 17418
rect 1171 17337 1177 17371
rect 1211 17337 1217 17371
rect 1171 17299 1217 17337
rect 1171 17265 1177 17299
rect 1211 17265 1217 17299
rect 1171 17227 1217 17265
rect 1171 17193 1177 17227
rect 1211 17193 1217 17227
rect 1171 17146 1217 17193
rect 1267 17371 1313 17418
rect 1267 17337 1273 17371
rect 1307 17337 1313 17371
rect 1267 17299 1313 17337
rect 1267 17265 1273 17299
rect 1307 17265 1313 17299
rect 1267 17227 1313 17265
rect 1267 17193 1273 17227
rect 1307 17193 1313 17227
rect 1267 17146 1313 17193
rect 1381 17402 1427 17440
rect 1381 17368 1387 17402
rect 1421 17368 1427 17402
rect 1381 17330 1427 17368
rect 1381 17296 1387 17330
rect 1421 17296 1427 17330
rect 1381 17258 1427 17296
rect 1381 17224 1387 17258
rect 1421 17224 1427 17258
rect 1381 17214 1427 17224
rect 1381 17212 2160 17214
rect 1381 17186 2056 17212
rect 1381 17161 1387 17186
rect 1380 17152 1387 17161
rect 1421 17152 2056 17186
rect 0 16971 163 17005
rect 129 16594 163 16971
rect 313 17005 347 17146
rect 505 17005 539 17146
rect 697 17005 731 17146
rect 889 17005 923 17146
rect 1081 17005 1115 17146
rect 1273 17005 1307 17146
rect 1380 17104 2056 17152
rect 2190 17104 2200 17212
rect 1380 17102 2160 17104
rect 2282 17009 2316 17572
rect 2447 17462 2457 17514
rect 2509 17462 2519 17514
rect 2562 17422 2596 17572
rect 2640 17462 2650 17514
rect 2702 17462 2712 17514
rect 2754 17422 2788 17572
rect 2831 17462 2841 17514
rect 2893 17462 2903 17514
rect 2946 17422 2980 17572
rect 3023 17462 3033 17514
rect 3085 17462 3095 17514
rect 3138 17422 3172 17572
rect 3215 17462 3225 17514
rect 3277 17462 3287 17514
rect 3330 17422 3364 17572
rect 3407 17462 3417 17514
rect 3469 17462 3479 17514
rect 3534 17478 3580 17686
rect 3534 17444 3540 17478
rect 3574 17444 3580 17478
rect 2460 17375 2506 17422
rect 2460 17341 2466 17375
rect 2500 17341 2506 17375
rect 2460 17303 2506 17341
rect 2460 17269 2466 17303
rect 2500 17269 2506 17303
rect 2460 17231 2506 17269
rect 2460 17197 2466 17231
rect 2500 17197 2506 17231
rect 2460 17150 2506 17197
rect 2556 17375 2602 17422
rect 2556 17341 2562 17375
rect 2596 17341 2602 17375
rect 2556 17303 2602 17341
rect 2556 17269 2562 17303
rect 2596 17269 2602 17303
rect 2556 17231 2602 17269
rect 2556 17197 2562 17231
rect 2596 17197 2602 17231
rect 2556 17150 2602 17197
rect 2652 17375 2698 17422
rect 2652 17341 2658 17375
rect 2692 17341 2698 17375
rect 2652 17303 2698 17341
rect 2652 17269 2658 17303
rect 2692 17269 2698 17303
rect 2652 17231 2698 17269
rect 2652 17197 2658 17231
rect 2692 17197 2698 17231
rect 2652 17150 2698 17197
rect 2748 17375 2794 17422
rect 2748 17341 2754 17375
rect 2788 17341 2794 17375
rect 2748 17303 2794 17341
rect 2748 17269 2754 17303
rect 2788 17269 2794 17303
rect 2748 17231 2794 17269
rect 2748 17197 2754 17231
rect 2788 17197 2794 17231
rect 2748 17150 2794 17197
rect 2844 17375 2890 17422
rect 2844 17341 2850 17375
rect 2884 17341 2890 17375
rect 2844 17303 2890 17341
rect 2844 17269 2850 17303
rect 2884 17269 2890 17303
rect 2844 17231 2890 17269
rect 2844 17197 2850 17231
rect 2884 17197 2890 17231
rect 2844 17150 2890 17197
rect 2940 17375 2986 17422
rect 2940 17341 2946 17375
rect 2980 17341 2986 17375
rect 2940 17303 2986 17341
rect 2940 17269 2946 17303
rect 2980 17269 2986 17303
rect 2940 17231 2986 17269
rect 2940 17197 2946 17231
rect 2980 17197 2986 17231
rect 2940 17150 2986 17197
rect 3036 17375 3082 17422
rect 3036 17341 3042 17375
rect 3076 17341 3082 17375
rect 3036 17303 3082 17341
rect 3036 17269 3042 17303
rect 3076 17269 3082 17303
rect 3036 17231 3082 17269
rect 3036 17197 3042 17231
rect 3076 17197 3082 17231
rect 3036 17150 3082 17197
rect 3132 17375 3178 17422
rect 3132 17341 3138 17375
rect 3172 17341 3178 17375
rect 3132 17303 3178 17341
rect 3132 17269 3138 17303
rect 3172 17269 3178 17303
rect 3132 17231 3178 17269
rect 3132 17197 3138 17231
rect 3172 17197 3178 17231
rect 3132 17150 3178 17197
rect 3228 17375 3274 17422
rect 3228 17341 3234 17375
rect 3268 17341 3274 17375
rect 3228 17303 3274 17341
rect 3228 17269 3234 17303
rect 3268 17269 3274 17303
rect 3228 17231 3274 17269
rect 3228 17197 3234 17231
rect 3268 17197 3274 17231
rect 3228 17150 3274 17197
rect 3324 17375 3370 17422
rect 3324 17341 3330 17375
rect 3364 17341 3370 17375
rect 3324 17303 3370 17341
rect 3324 17269 3330 17303
rect 3364 17269 3370 17303
rect 3324 17231 3370 17269
rect 3324 17197 3330 17231
rect 3364 17197 3370 17231
rect 3324 17150 3370 17197
rect 3420 17375 3466 17422
rect 3420 17341 3426 17375
rect 3460 17341 3466 17375
rect 3420 17303 3466 17341
rect 3420 17269 3426 17303
rect 3460 17269 3466 17303
rect 3420 17231 3466 17269
rect 3420 17197 3426 17231
rect 3460 17197 3466 17231
rect 3420 17150 3466 17197
rect 3534 17406 3580 17444
rect 3534 17372 3540 17406
rect 3574 17372 3580 17406
rect 3534 17334 3580 17372
rect 3534 17300 3540 17334
rect 3574 17300 3580 17334
rect 3534 17262 3580 17300
rect 3534 17228 3540 17262
rect 3574 17228 3580 17262
rect 3534 17190 3580 17228
rect 3534 17156 3540 17190
rect 3574 17156 3580 17190
rect 2101 17005 2316 17009
rect 313 16975 2316 17005
rect 313 16971 2141 16975
rect 313 16838 347 16971
rect 505 16838 539 16971
rect 697 16838 731 16971
rect 889 16838 923 16971
rect 1081 16838 1115 16971
rect 1273 16838 1307 16971
rect 1381 16845 1608 16868
rect 307 16803 353 16838
rect 307 16769 313 16803
rect 347 16769 353 16803
rect 307 16734 353 16769
rect 403 16803 449 16838
rect 403 16769 409 16803
rect 443 16769 449 16803
rect 403 16734 449 16769
rect 499 16803 545 16838
rect 499 16769 505 16803
rect 539 16769 545 16803
rect 499 16734 545 16769
rect 595 16803 641 16838
rect 595 16769 601 16803
rect 635 16769 641 16803
rect 595 16734 641 16769
rect 691 16803 737 16838
rect 691 16769 697 16803
rect 731 16769 737 16803
rect 691 16734 737 16769
rect 787 16803 833 16838
rect 787 16769 793 16803
rect 827 16769 833 16803
rect 787 16734 833 16769
rect 883 16803 929 16838
rect 883 16769 889 16803
rect 923 16769 929 16803
rect 883 16734 929 16769
rect 979 16803 1025 16838
rect 979 16769 985 16803
rect 1019 16769 1025 16803
rect 979 16734 1025 16769
rect 1075 16803 1121 16838
rect 1075 16769 1081 16803
rect 1115 16769 1121 16803
rect 1075 16734 1121 16769
rect 1171 16803 1217 16838
rect 1171 16769 1177 16803
rect 1211 16769 1217 16803
rect 1171 16734 1217 16769
rect 1267 16803 1313 16838
rect 1267 16769 1273 16803
rect 1307 16769 1313 16803
rect 1267 16734 1313 16769
rect 1381 16811 1387 16845
rect 1421 16811 1608 16845
rect 1381 16773 1608 16811
rect 1381 16739 1387 16773
rect 1421 16748 1608 16773
rect 1421 16739 1427 16748
rect 1560 16746 1608 16748
rect 1598 16744 1608 16746
rect 1720 16744 1730 16868
rect 297 16703 363 16706
rect 294 16651 304 16703
rect 356 16651 366 16703
rect 297 16646 363 16651
rect 409 16594 443 16734
rect 489 16703 555 16706
rect 485 16651 495 16703
rect 547 16651 557 16703
rect 489 16646 555 16651
rect 601 16594 635 16734
rect 681 16703 747 16706
rect 677 16651 687 16703
rect 739 16651 749 16703
rect 681 16646 747 16651
rect 793 16594 827 16734
rect 873 16703 939 16706
rect 869 16651 879 16703
rect 931 16651 941 16703
rect 873 16646 939 16651
rect 985 16594 1019 16734
rect 1065 16702 1131 16706
rect 1062 16650 1072 16702
rect 1124 16650 1134 16702
rect 1065 16646 1131 16650
rect 1177 16594 1211 16734
rect 1257 16702 1323 16706
rect 1254 16650 1264 16702
rect 1316 16650 1326 16702
rect 1381 16701 1427 16739
rect 1920 16706 1930 16708
rect 1381 16667 1387 16701
rect 1421 16667 1427 16701
rect 1257 16646 1323 16650
rect 129 16560 1211 16594
rect 1381 16524 1427 16667
rect 1458 16650 1468 16706
rect 1524 16652 1930 16706
rect 1986 16652 1996 16708
rect 1524 16650 1986 16652
rect 2282 16598 2316 16975
rect 2466 17009 2500 17150
rect 2658 17009 2692 17150
rect 2850 17009 2884 17150
rect 3042 17009 3076 17150
rect 3234 17009 3268 17150
rect 3426 17009 3460 17150
rect 3534 17112 3580 17156
rect 3803 17572 4885 17606
rect 3803 17009 3837 17572
rect 3968 17462 3978 17514
rect 4030 17462 4040 17514
rect 4083 17422 4117 17572
rect 4161 17462 4171 17514
rect 4223 17462 4233 17514
rect 4275 17422 4309 17572
rect 4352 17462 4362 17514
rect 4414 17462 4424 17514
rect 4467 17422 4501 17572
rect 4544 17462 4554 17514
rect 4606 17462 4616 17514
rect 4659 17422 4693 17572
rect 4736 17462 4746 17514
rect 4798 17462 4808 17514
rect 4851 17422 4885 17572
rect 4928 17462 4938 17514
rect 4990 17462 5000 17514
rect 5055 17478 5101 17683
rect 5055 17444 5061 17478
rect 5095 17444 5101 17478
rect 3981 17375 4027 17422
rect 3981 17341 3987 17375
rect 4021 17341 4027 17375
rect 3981 17303 4027 17341
rect 3981 17269 3987 17303
rect 4021 17269 4027 17303
rect 3981 17231 4027 17269
rect 3981 17197 3987 17231
rect 4021 17197 4027 17231
rect 3981 17150 4027 17197
rect 4077 17375 4123 17422
rect 4077 17341 4083 17375
rect 4117 17341 4123 17375
rect 4077 17303 4123 17341
rect 4077 17269 4083 17303
rect 4117 17269 4123 17303
rect 4077 17231 4123 17269
rect 4077 17197 4083 17231
rect 4117 17197 4123 17231
rect 4077 17150 4123 17197
rect 4173 17375 4219 17422
rect 4173 17341 4179 17375
rect 4213 17341 4219 17375
rect 4173 17303 4219 17341
rect 4173 17269 4179 17303
rect 4213 17269 4219 17303
rect 4173 17231 4219 17269
rect 4173 17197 4179 17231
rect 4213 17197 4219 17231
rect 4173 17150 4219 17197
rect 4269 17375 4315 17422
rect 4269 17341 4275 17375
rect 4309 17341 4315 17375
rect 4269 17303 4315 17341
rect 4269 17269 4275 17303
rect 4309 17269 4315 17303
rect 4269 17231 4315 17269
rect 4269 17197 4275 17231
rect 4309 17197 4315 17231
rect 4269 17150 4315 17197
rect 4365 17375 4411 17422
rect 4365 17341 4371 17375
rect 4405 17341 4411 17375
rect 4365 17303 4411 17341
rect 4365 17269 4371 17303
rect 4405 17269 4411 17303
rect 4365 17231 4411 17269
rect 4365 17197 4371 17231
rect 4405 17197 4411 17231
rect 4365 17150 4411 17197
rect 4461 17375 4507 17422
rect 4461 17341 4467 17375
rect 4501 17341 4507 17375
rect 4461 17303 4507 17341
rect 4461 17269 4467 17303
rect 4501 17269 4507 17303
rect 4461 17231 4507 17269
rect 4461 17197 4467 17231
rect 4501 17197 4507 17231
rect 4461 17150 4507 17197
rect 4557 17375 4603 17422
rect 4557 17341 4563 17375
rect 4597 17341 4603 17375
rect 4557 17303 4603 17341
rect 4557 17269 4563 17303
rect 4597 17269 4603 17303
rect 4557 17231 4603 17269
rect 4557 17197 4563 17231
rect 4597 17197 4603 17231
rect 4557 17150 4603 17197
rect 4653 17375 4699 17422
rect 4653 17341 4659 17375
rect 4693 17341 4699 17375
rect 4653 17303 4699 17341
rect 4653 17269 4659 17303
rect 4693 17269 4699 17303
rect 4653 17231 4699 17269
rect 4653 17197 4659 17231
rect 4693 17197 4699 17231
rect 4653 17150 4699 17197
rect 4749 17375 4795 17422
rect 4749 17341 4755 17375
rect 4789 17341 4795 17375
rect 4749 17303 4795 17341
rect 4749 17269 4755 17303
rect 4789 17269 4795 17303
rect 4749 17231 4795 17269
rect 4749 17197 4755 17231
rect 4789 17197 4795 17231
rect 4749 17150 4795 17197
rect 4845 17375 4891 17422
rect 4845 17341 4851 17375
rect 4885 17341 4891 17375
rect 4845 17303 4891 17341
rect 4845 17269 4851 17303
rect 4885 17269 4891 17303
rect 4845 17231 4891 17269
rect 4845 17197 4851 17231
rect 4885 17197 4891 17231
rect 4845 17150 4891 17197
rect 4941 17375 4987 17422
rect 4941 17341 4947 17375
rect 4981 17341 4987 17375
rect 4941 17303 4987 17341
rect 4941 17269 4947 17303
rect 4981 17269 4987 17303
rect 4941 17231 4987 17269
rect 4941 17197 4947 17231
rect 4981 17197 4987 17231
rect 4941 17150 4987 17197
rect 5055 17406 5101 17444
rect 5055 17372 5061 17406
rect 5095 17372 5101 17406
rect 5055 17334 5101 17372
rect 5055 17300 5061 17334
rect 5095 17303 5101 17334
rect 5274 17303 5550 17304
rect 5095 17300 5550 17303
rect 5055 17273 5550 17300
rect 5055 17262 5303 17273
rect 5055 17228 5061 17262
rect 5095 17239 5303 17262
rect 5337 17239 5395 17273
rect 5429 17239 5487 17273
rect 5521 17239 5550 17273
rect 5095 17228 5550 17239
rect 5055 17208 5550 17228
rect 5055 17190 5101 17208
rect 5055 17156 5061 17190
rect 5095 17156 5101 17190
rect 2466 16975 3837 17009
rect 2466 16842 2500 16975
rect 2658 16842 2692 16975
rect 2850 16842 2884 16975
rect 3042 16842 3076 16975
rect 3234 16842 3268 16975
rect 3426 16842 3460 16975
rect 3671 16885 3681 16937
rect 3733 16885 3743 16937
rect 3679 16884 3691 16885
rect 3725 16884 3737 16885
rect 3679 16878 3737 16884
rect 3534 16849 3580 16872
rect 2460 16807 2506 16842
rect 2460 16773 2466 16807
rect 2500 16773 2506 16807
rect 2460 16738 2506 16773
rect 2556 16807 2602 16842
rect 2556 16773 2562 16807
rect 2596 16773 2602 16807
rect 2556 16738 2602 16773
rect 2652 16807 2698 16842
rect 2652 16773 2658 16807
rect 2692 16773 2698 16807
rect 2652 16738 2698 16773
rect 2748 16807 2794 16842
rect 2748 16773 2754 16807
rect 2788 16773 2794 16807
rect 2748 16738 2794 16773
rect 2844 16807 2890 16842
rect 2844 16773 2850 16807
rect 2884 16773 2890 16807
rect 2844 16738 2890 16773
rect 2940 16807 2986 16842
rect 2940 16773 2946 16807
rect 2980 16773 2986 16807
rect 2940 16738 2986 16773
rect 3036 16807 3082 16842
rect 3036 16773 3042 16807
rect 3076 16773 3082 16807
rect 3036 16738 3082 16773
rect 3132 16807 3178 16842
rect 3132 16773 3138 16807
rect 3172 16773 3178 16807
rect 3132 16738 3178 16773
rect 3228 16807 3274 16842
rect 3228 16773 3234 16807
rect 3268 16773 3274 16807
rect 3228 16738 3274 16773
rect 3324 16807 3370 16842
rect 3324 16773 3330 16807
rect 3364 16773 3370 16807
rect 3324 16738 3370 16773
rect 3420 16807 3466 16842
rect 3420 16773 3426 16807
rect 3460 16773 3466 16807
rect 3420 16738 3466 16773
rect 3534 16815 3540 16849
rect 3574 16847 3580 16849
rect 3803 16847 3837 16975
rect 3574 16846 3680 16847
rect 3734 16846 3837 16847
rect 3574 16834 3687 16846
rect 3574 16815 3647 16834
rect 3534 16777 3647 16815
rect 3534 16743 3540 16777
rect 3574 16758 3647 16777
rect 3681 16758 3687 16834
rect 3574 16747 3687 16758
rect 3574 16743 3580 16747
rect 3641 16746 3687 16747
rect 3729 16834 3837 16846
rect 3987 17009 4021 17150
rect 4179 17009 4213 17150
rect 4371 17009 4405 17150
rect 4563 17009 4597 17150
rect 4755 17009 4789 17150
rect 4947 17009 4981 17150
rect 5055 17112 5101 17156
rect 5683 17063 5743 18316
rect 5177 17029 5743 17063
rect 5177 17009 5211 17029
rect 3987 16975 5211 17009
rect 3987 16842 4021 16975
rect 4179 16842 4213 16975
rect 4371 16842 4405 16975
rect 4563 16842 4597 16975
rect 4755 16842 4789 16975
rect 4947 16842 4981 16975
rect 5438 16971 5512 16972
rect 5326 16969 5400 16970
rect 5326 16917 5337 16969
rect 5389 16917 5400 16969
rect 5438 16919 5449 16971
rect 5501 16919 5512 16971
rect 5438 16918 5512 16919
rect 5326 16916 5400 16917
rect 5055 16849 5101 16872
rect 3729 16758 3735 16834
rect 3769 16758 3837 16834
rect 3729 16747 3837 16758
rect 3729 16746 3775 16747
rect 2450 16707 2516 16710
rect 2447 16655 2457 16707
rect 2509 16655 2519 16707
rect 2450 16650 2516 16655
rect 2562 16598 2596 16738
rect 2642 16707 2708 16710
rect 2638 16655 2648 16707
rect 2700 16655 2710 16707
rect 2642 16650 2708 16655
rect 2754 16598 2788 16738
rect 2834 16707 2900 16710
rect 2830 16655 2840 16707
rect 2892 16655 2902 16707
rect 2834 16650 2900 16655
rect 2946 16598 2980 16738
rect 3026 16707 3092 16710
rect 3022 16655 3032 16707
rect 3084 16655 3094 16707
rect 3026 16650 3092 16655
rect 3138 16598 3172 16738
rect 3218 16706 3284 16710
rect 3215 16654 3225 16706
rect 3277 16654 3287 16706
rect 3218 16650 3284 16654
rect 3330 16598 3364 16738
rect 3410 16706 3476 16710
rect 3407 16654 3417 16706
rect 3469 16654 3479 16706
rect 3534 16705 3580 16743
rect 3534 16671 3540 16705
rect 3574 16671 3580 16705
rect 3410 16650 3476 16654
rect 2282 16564 3364 16598
rect 3534 16488 3580 16671
rect 3803 16598 3837 16747
rect 3981 16807 4027 16842
rect 3981 16773 3987 16807
rect 4021 16773 4027 16807
rect 3981 16738 4027 16773
rect 4077 16807 4123 16842
rect 4077 16773 4083 16807
rect 4117 16773 4123 16807
rect 4077 16738 4123 16773
rect 4173 16807 4219 16842
rect 4173 16773 4179 16807
rect 4213 16773 4219 16807
rect 4173 16738 4219 16773
rect 4269 16807 4315 16842
rect 4269 16773 4275 16807
rect 4309 16773 4315 16807
rect 4269 16738 4315 16773
rect 4365 16807 4411 16842
rect 4365 16773 4371 16807
rect 4405 16773 4411 16807
rect 4365 16738 4411 16773
rect 4461 16807 4507 16842
rect 4461 16773 4467 16807
rect 4501 16773 4507 16807
rect 4461 16738 4507 16773
rect 4557 16807 4603 16842
rect 4557 16773 4563 16807
rect 4597 16773 4603 16807
rect 4557 16738 4603 16773
rect 4653 16807 4699 16842
rect 4653 16773 4659 16807
rect 4693 16773 4699 16807
rect 4653 16738 4699 16773
rect 4749 16807 4795 16842
rect 4749 16773 4755 16807
rect 4789 16773 4795 16807
rect 4749 16738 4795 16773
rect 4845 16807 4891 16842
rect 4845 16773 4851 16807
rect 4885 16773 4891 16807
rect 4845 16738 4891 16773
rect 4941 16807 4987 16842
rect 4941 16773 4947 16807
rect 4981 16773 4987 16807
rect 4941 16738 4987 16773
rect 5055 16815 5061 16849
rect 5095 16815 5101 16849
rect 5055 16777 5101 16815
rect 5055 16743 5061 16777
rect 5095 16760 5101 16777
rect 5095 16743 5550 16760
rect 3971 16707 4037 16710
rect 3968 16655 3978 16707
rect 4030 16655 4040 16707
rect 3971 16650 4037 16655
rect 4083 16598 4117 16738
rect 4163 16707 4229 16710
rect 4159 16655 4169 16707
rect 4221 16655 4231 16707
rect 4163 16650 4229 16655
rect 4275 16598 4309 16738
rect 4355 16707 4421 16710
rect 4351 16655 4361 16707
rect 4413 16655 4423 16707
rect 4355 16650 4421 16655
rect 4467 16598 4501 16738
rect 4547 16707 4613 16710
rect 4543 16655 4553 16707
rect 4605 16655 4615 16707
rect 4547 16650 4613 16655
rect 4659 16598 4693 16738
rect 4739 16706 4805 16710
rect 4736 16654 4746 16706
rect 4798 16654 4808 16706
rect 4739 16650 4805 16654
rect 4851 16598 4885 16738
rect 5055 16729 5550 16743
rect 4931 16706 4997 16710
rect 4928 16654 4938 16706
rect 4990 16654 5000 16706
rect 5055 16705 5303 16729
rect 5055 16671 5061 16705
rect 5095 16695 5303 16705
rect 5337 16695 5395 16729
rect 5429 16695 5487 16729
rect 5521 16695 5550 16729
rect 5095 16671 5550 16695
rect 5055 16664 5550 16671
rect 4931 16650 4997 16654
rect 3803 16564 4885 16598
rect 5055 16489 5101 16664
rect 129 16281 1211 16315
rect 129 15718 163 16281
rect 294 16171 304 16223
rect 356 16171 366 16223
rect 409 16131 443 16281
rect 487 16171 497 16223
rect 549 16171 559 16223
rect 601 16131 635 16281
rect 678 16171 688 16223
rect 740 16171 750 16223
rect 793 16131 827 16281
rect 870 16171 880 16223
rect 932 16171 942 16223
rect 985 16131 1019 16281
rect 1062 16171 1072 16223
rect 1124 16171 1134 16223
rect 1177 16131 1211 16281
rect 1254 16171 1264 16223
rect 1316 16171 1326 16223
rect 1381 16187 1427 16351
rect 2282 16285 3364 16319
rect 1381 16153 1387 16187
rect 1421 16153 1427 16187
rect 1512 16164 1522 16224
rect 1578 16164 1792 16224
rect 1852 16164 1862 16224
rect 307 16084 353 16131
rect 307 16050 313 16084
rect 347 16050 353 16084
rect 307 16012 353 16050
rect 307 15978 313 16012
rect 347 15978 353 16012
rect 307 15940 353 15978
rect 307 15906 313 15940
rect 347 15906 353 15940
rect 307 15859 353 15906
rect 403 16084 449 16131
rect 403 16050 409 16084
rect 443 16050 449 16084
rect 403 16012 449 16050
rect 403 15978 409 16012
rect 443 15978 449 16012
rect 403 15940 449 15978
rect 403 15906 409 15940
rect 443 15906 449 15940
rect 403 15859 449 15906
rect 499 16084 545 16131
rect 499 16050 505 16084
rect 539 16050 545 16084
rect 499 16012 545 16050
rect 499 15978 505 16012
rect 539 15978 545 16012
rect 499 15940 545 15978
rect 499 15906 505 15940
rect 539 15906 545 15940
rect 499 15859 545 15906
rect 595 16084 641 16131
rect 595 16050 601 16084
rect 635 16050 641 16084
rect 595 16012 641 16050
rect 595 15978 601 16012
rect 635 15978 641 16012
rect 595 15940 641 15978
rect 595 15906 601 15940
rect 635 15906 641 15940
rect 595 15859 641 15906
rect 691 16084 737 16131
rect 691 16050 697 16084
rect 731 16050 737 16084
rect 691 16012 737 16050
rect 691 15978 697 16012
rect 731 15978 737 16012
rect 691 15940 737 15978
rect 691 15906 697 15940
rect 731 15906 737 15940
rect 691 15859 737 15906
rect 787 16084 833 16131
rect 787 16050 793 16084
rect 827 16050 833 16084
rect 787 16012 833 16050
rect 787 15978 793 16012
rect 827 15978 833 16012
rect 787 15940 833 15978
rect 787 15906 793 15940
rect 827 15906 833 15940
rect 787 15859 833 15906
rect 883 16084 929 16131
rect 883 16050 889 16084
rect 923 16050 929 16084
rect 883 16012 929 16050
rect 883 15978 889 16012
rect 923 15978 929 16012
rect 883 15940 929 15978
rect 883 15906 889 15940
rect 923 15906 929 15940
rect 883 15859 929 15906
rect 979 16084 1025 16131
rect 979 16050 985 16084
rect 1019 16050 1025 16084
rect 979 16012 1025 16050
rect 979 15978 985 16012
rect 1019 15978 1025 16012
rect 979 15940 1025 15978
rect 979 15906 985 15940
rect 1019 15906 1025 15940
rect 979 15859 1025 15906
rect 1075 16084 1121 16131
rect 1075 16050 1081 16084
rect 1115 16050 1121 16084
rect 1075 16012 1121 16050
rect 1075 15978 1081 16012
rect 1115 15978 1121 16012
rect 1075 15940 1121 15978
rect 1075 15906 1081 15940
rect 1115 15906 1121 15940
rect 1075 15859 1121 15906
rect 1171 16084 1217 16131
rect 1171 16050 1177 16084
rect 1211 16050 1217 16084
rect 1171 16012 1217 16050
rect 1171 15978 1177 16012
rect 1211 15978 1217 16012
rect 1171 15940 1217 15978
rect 1171 15906 1177 15940
rect 1211 15906 1217 15940
rect 1171 15859 1217 15906
rect 1267 16084 1313 16131
rect 1267 16050 1273 16084
rect 1307 16050 1313 16084
rect 1267 16012 1313 16050
rect 1267 15978 1273 16012
rect 1307 15978 1313 16012
rect 1267 15940 1313 15978
rect 1267 15906 1273 15940
rect 1307 15906 1313 15940
rect 1267 15859 1313 15906
rect 1381 16115 1427 16153
rect 1381 16081 1387 16115
rect 1421 16081 1427 16115
rect 1381 16043 1427 16081
rect 1381 16009 1387 16043
rect 1421 16009 1427 16043
rect 1381 15971 1427 16009
rect 1381 15937 1387 15971
rect 1421 15937 1427 15971
rect 1381 15927 1427 15937
rect 1381 15925 2160 15927
rect 1381 15899 2056 15925
rect 1381 15874 1387 15899
rect 1380 15865 1387 15874
rect 1421 15865 2056 15899
rect 0 15684 163 15718
rect 129 15307 163 15684
rect 313 15718 347 15859
rect 505 15718 539 15859
rect 697 15718 731 15859
rect 889 15718 923 15859
rect 1081 15718 1115 15859
rect 1273 15718 1307 15859
rect 1380 15817 2056 15865
rect 2190 15817 2200 15925
rect 1380 15815 2160 15817
rect 2282 15722 2316 16285
rect 2447 16175 2457 16227
rect 2509 16175 2519 16227
rect 2562 16135 2596 16285
rect 2640 16175 2650 16227
rect 2702 16175 2712 16227
rect 2754 16135 2788 16285
rect 2831 16175 2841 16227
rect 2893 16175 2903 16227
rect 2946 16135 2980 16285
rect 3023 16175 3033 16227
rect 3085 16175 3095 16227
rect 3138 16135 3172 16285
rect 3215 16175 3225 16227
rect 3277 16175 3287 16227
rect 3330 16135 3364 16285
rect 3407 16175 3417 16227
rect 3469 16175 3479 16227
rect 3534 16191 3580 16399
rect 3534 16157 3540 16191
rect 3574 16157 3580 16191
rect 2460 16088 2506 16135
rect 2460 16054 2466 16088
rect 2500 16054 2506 16088
rect 2460 16016 2506 16054
rect 2460 15982 2466 16016
rect 2500 15982 2506 16016
rect 2460 15944 2506 15982
rect 2460 15910 2466 15944
rect 2500 15910 2506 15944
rect 2460 15863 2506 15910
rect 2556 16088 2602 16135
rect 2556 16054 2562 16088
rect 2596 16054 2602 16088
rect 2556 16016 2602 16054
rect 2556 15982 2562 16016
rect 2596 15982 2602 16016
rect 2556 15944 2602 15982
rect 2556 15910 2562 15944
rect 2596 15910 2602 15944
rect 2556 15863 2602 15910
rect 2652 16088 2698 16135
rect 2652 16054 2658 16088
rect 2692 16054 2698 16088
rect 2652 16016 2698 16054
rect 2652 15982 2658 16016
rect 2692 15982 2698 16016
rect 2652 15944 2698 15982
rect 2652 15910 2658 15944
rect 2692 15910 2698 15944
rect 2652 15863 2698 15910
rect 2748 16088 2794 16135
rect 2748 16054 2754 16088
rect 2788 16054 2794 16088
rect 2748 16016 2794 16054
rect 2748 15982 2754 16016
rect 2788 15982 2794 16016
rect 2748 15944 2794 15982
rect 2748 15910 2754 15944
rect 2788 15910 2794 15944
rect 2748 15863 2794 15910
rect 2844 16088 2890 16135
rect 2844 16054 2850 16088
rect 2884 16054 2890 16088
rect 2844 16016 2890 16054
rect 2844 15982 2850 16016
rect 2884 15982 2890 16016
rect 2844 15944 2890 15982
rect 2844 15910 2850 15944
rect 2884 15910 2890 15944
rect 2844 15863 2890 15910
rect 2940 16088 2986 16135
rect 2940 16054 2946 16088
rect 2980 16054 2986 16088
rect 2940 16016 2986 16054
rect 2940 15982 2946 16016
rect 2980 15982 2986 16016
rect 2940 15944 2986 15982
rect 2940 15910 2946 15944
rect 2980 15910 2986 15944
rect 2940 15863 2986 15910
rect 3036 16088 3082 16135
rect 3036 16054 3042 16088
rect 3076 16054 3082 16088
rect 3036 16016 3082 16054
rect 3036 15982 3042 16016
rect 3076 15982 3082 16016
rect 3036 15944 3082 15982
rect 3036 15910 3042 15944
rect 3076 15910 3082 15944
rect 3036 15863 3082 15910
rect 3132 16088 3178 16135
rect 3132 16054 3138 16088
rect 3172 16054 3178 16088
rect 3132 16016 3178 16054
rect 3132 15982 3138 16016
rect 3172 15982 3178 16016
rect 3132 15944 3178 15982
rect 3132 15910 3138 15944
rect 3172 15910 3178 15944
rect 3132 15863 3178 15910
rect 3228 16088 3274 16135
rect 3228 16054 3234 16088
rect 3268 16054 3274 16088
rect 3228 16016 3274 16054
rect 3228 15982 3234 16016
rect 3268 15982 3274 16016
rect 3228 15944 3274 15982
rect 3228 15910 3234 15944
rect 3268 15910 3274 15944
rect 3228 15863 3274 15910
rect 3324 16088 3370 16135
rect 3324 16054 3330 16088
rect 3364 16054 3370 16088
rect 3324 16016 3370 16054
rect 3324 15982 3330 16016
rect 3364 15982 3370 16016
rect 3324 15944 3370 15982
rect 3324 15910 3330 15944
rect 3364 15910 3370 15944
rect 3324 15863 3370 15910
rect 3420 16088 3466 16135
rect 3420 16054 3426 16088
rect 3460 16054 3466 16088
rect 3420 16016 3466 16054
rect 3420 15982 3426 16016
rect 3460 15982 3466 16016
rect 3420 15944 3466 15982
rect 3420 15910 3426 15944
rect 3460 15910 3466 15944
rect 3420 15863 3466 15910
rect 3534 16119 3580 16157
rect 3534 16085 3540 16119
rect 3574 16085 3580 16119
rect 3534 16047 3580 16085
rect 3534 16013 3540 16047
rect 3574 16013 3580 16047
rect 3534 15975 3580 16013
rect 3534 15941 3540 15975
rect 3574 15941 3580 15975
rect 3534 15903 3580 15941
rect 3534 15869 3540 15903
rect 3574 15869 3580 15903
rect 2101 15718 2316 15722
rect 313 15688 2316 15718
rect 313 15684 2141 15688
rect 313 15551 347 15684
rect 505 15551 539 15684
rect 697 15551 731 15684
rect 889 15551 923 15684
rect 1081 15551 1115 15684
rect 1273 15551 1307 15684
rect 1381 15558 1608 15581
rect 307 15516 353 15551
rect 307 15482 313 15516
rect 347 15482 353 15516
rect 307 15447 353 15482
rect 403 15516 449 15551
rect 403 15482 409 15516
rect 443 15482 449 15516
rect 403 15447 449 15482
rect 499 15516 545 15551
rect 499 15482 505 15516
rect 539 15482 545 15516
rect 499 15447 545 15482
rect 595 15516 641 15551
rect 595 15482 601 15516
rect 635 15482 641 15516
rect 595 15447 641 15482
rect 691 15516 737 15551
rect 691 15482 697 15516
rect 731 15482 737 15516
rect 691 15447 737 15482
rect 787 15516 833 15551
rect 787 15482 793 15516
rect 827 15482 833 15516
rect 787 15447 833 15482
rect 883 15516 929 15551
rect 883 15482 889 15516
rect 923 15482 929 15516
rect 883 15447 929 15482
rect 979 15516 1025 15551
rect 979 15482 985 15516
rect 1019 15482 1025 15516
rect 979 15447 1025 15482
rect 1075 15516 1121 15551
rect 1075 15482 1081 15516
rect 1115 15482 1121 15516
rect 1075 15447 1121 15482
rect 1171 15516 1217 15551
rect 1171 15482 1177 15516
rect 1211 15482 1217 15516
rect 1171 15447 1217 15482
rect 1267 15516 1313 15551
rect 1267 15482 1273 15516
rect 1307 15482 1313 15516
rect 1267 15447 1313 15482
rect 1381 15524 1387 15558
rect 1421 15524 1608 15558
rect 1381 15486 1608 15524
rect 1381 15452 1387 15486
rect 1421 15461 1608 15486
rect 1421 15452 1427 15461
rect 1560 15459 1608 15461
rect 1598 15457 1608 15459
rect 1720 15457 1730 15581
rect 297 15416 363 15419
rect 294 15364 304 15416
rect 356 15364 366 15416
rect 297 15359 363 15364
rect 409 15307 443 15447
rect 489 15416 555 15419
rect 485 15364 495 15416
rect 547 15364 557 15416
rect 489 15359 555 15364
rect 601 15307 635 15447
rect 681 15416 747 15419
rect 677 15364 687 15416
rect 739 15364 749 15416
rect 681 15359 747 15364
rect 793 15307 827 15447
rect 873 15416 939 15419
rect 869 15364 879 15416
rect 931 15364 941 15416
rect 873 15359 939 15364
rect 985 15307 1019 15447
rect 1065 15415 1131 15419
rect 1062 15363 1072 15415
rect 1124 15363 1134 15415
rect 1065 15359 1131 15363
rect 1177 15307 1211 15447
rect 1257 15415 1323 15419
rect 1254 15363 1264 15415
rect 1316 15363 1326 15415
rect 1381 15414 1427 15452
rect 1920 15419 1930 15421
rect 1381 15380 1387 15414
rect 1421 15380 1427 15414
rect 1257 15359 1323 15363
rect 129 15273 1211 15307
rect 1381 15237 1427 15380
rect 1458 15363 1468 15419
rect 1524 15365 1930 15419
rect 1986 15365 1996 15421
rect 1524 15363 1986 15365
rect 2282 15311 2316 15688
rect 2466 15722 2500 15863
rect 2658 15722 2692 15863
rect 2850 15722 2884 15863
rect 3042 15722 3076 15863
rect 3234 15722 3268 15863
rect 3426 15722 3460 15863
rect 3534 15825 3580 15869
rect 3803 16285 4885 16319
rect 3803 15722 3837 16285
rect 3968 16175 3978 16227
rect 4030 16175 4040 16227
rect 4083 16135 4117 16285
rect 4161 16175 4171 16227
rect 4223 16175 4233 16227
rect 4275 16135 4309 16285
rect 4352 16175 4362 16227
rect 4414 16175 4424 16227
rect 4467 16135 4501 16285
rect 4544 16175 4554 16227
rect 4606 16175 4616 16227
rect 4659 16135 4693 16285
rect 4736 16175 4746 16227
rect 4798 16175 4808 16227
rect 4851 16135 4885 16285
rect 4928 16175 4938 16227
rect 4990 16175 5000 16227
rect 5055 16191 5101 16396
rect 5055 16157 5061 16191
rect 5095 16157 5101 16191
rect 3981 16088 4027 16135
rect 3981 16054 3987 16088
rect 4021 16054 4027 16088
rect 3981 16016 4027 16054
rect 3981 15982 3987 16016
rect 4021 15982 4027 16016
rect 3981 15944 4027 15982
rect 3981 15910 3987 15944
rect 4021 15910 4027 15944
rect 3981 15863 4027 15910
rect 4077 16088 4123 16135
rect 4077 16054 4083 16088
rect 4117 16054 4123 16088
rect 4077 16016 4123 16054
rect 4077 15982 4083 16016
rect 4117 15982 4123 16016
rect 4077 15944 4123 15982
rect 4077 15910 4083 15944
rect 4117 15910 4123 15944
rect 4077 15863 4123 15910
rect 4173 16088 4219 16135
rect 4173 16054 4179 16088
rect 4213 16054 4219 16088
rect 4173 16016 4219 16054
rect 4173 15982 4179 16016
rect 4213 15982 4219 16016
rect 4173 15944 4219 15982
rect 4173 15910 4179 15944
rect 4213 15910 4219 15944
rect 4173 15863 4219 15910
rect 4269 16088 4315 16135
rect 4269 16054 4275 16088
rect 4309 16054 4315 16088
rect 4269 16016 4315 16054
rect 4269 15982 4275 16016
rect 4309 15982 4315 16016
rect 4269 15944 4315 15982
rect 4269 15910 4275 15944
rect 4309 15910 4315 15944
rect 4269 15863 4315 15910
rect 4365 16088 4411 16135
rect 4365 16054 4371 16088
rect 4405 16054 4411 16088
rect 4365 16016 4411 16054
rect 4365 15982 4371 16016
rect 4405 15982 4411 16016
rect 4365 15944 4411 15982
rect 4365 15910 4371 15944
rect 4405 15910 4411 15944
rect 4365 15863 4411 15910
rect 4461 16088 4507 16135
rect 4461 16054 4467 16088
rect 4501 16054 4507 16088
rect 4461 16016 4507 16054
rect 4461 15982 4467 16016
rect 4501 15982 4507 16016
rect 4461 15944 4507 15982
rect 4461 15910 4467 15944
rect 4501 15910 4507 15944
rect 4461 15863 4507 15910
rect 4557 16088 4603 16135
rect 4557 16054 4563 16088
rect 4597 16054 4603 16088
rect 4557 16016 4603 16054
rect 4557 15982 4563 16016
rect 4597 15982 4603 16016
rect 4557 15944 4603 15982
rect 4557 15910 4563 15944
rect 4597 15910 4603 15944
rect 4557 15863 4603 15910
rect 4653 16088 4699 16135
rect 4653 16054 4659 16088
rect 4693 16054 4699 16088
rect 4653 16016 4699 16054
rect 4653 15982 4659 16016
rect 4693 15982 4699 16016
rect 4653 15944 4699 15982
rect 4653 15910 4659 15944
rect 4693 15910 4699 15944
rect 4653 15863 4699 15910
rect 4749 16088 4795 16135
rect 4749 16054 4755 16088
rect 4789 16054 4795 16088
rect 4749 16016 4795 16054
rect 4749 15982 4755 16016
rect 4789 15982 4795 16016
rect 4749 15944 4795 15982
rect 4749 15910 4755 15944
rect 4789 15910 4795 15944
rect 4749 15863 4795 15910
rect 4845 16088 4891 16135
rect 4845 16054 4851 16088
rect 4885 16054 4891 16088
rect 4845 16016 4891 16054
rect 4845 15982 4851 16016
rect 4885 15982 4891 16016
rect 4845 15944 4891 15982
rect 4845 15910 4851 15944
rect 4885 15910 4891 15944
rect 4845 15863 4891 15910
rect 4941 16088 4987 16135
rect 4941 16054 4947 16088
rect 4981 16054 4987 16088
rect 4941 16016 4987 16054
rect 4941 15982 4947 16016
rect 4981 15982 4987 16016
rect 4941 15944 4987 15982
rect 4941 15910 4947 15944
rect 4981 15910 4987 15944
rect 4941 15863 4987 15910
rect 5055 16119 5101 16157
rect 5055 16085 5061 16119
rect 5095 16085 5101 16119
rect 5055 16047 5101 16085
rect 5055 16013 5061 16047
rect 5095 16016 5101 16047
rect 5274 16016 5550 16017
rect 5095 16013 5550 16016
rect 5055 15986 5550 16013
rect 5055 15975 5303 15986
rect 5055 15941 5061 15975
rect 5095 15952 5303 15975
rect 5337 15952 5395 15986
rect 5429 15952 5487 15986
rect 5521 15952 5550 15986
rect 5095 15941 5550 15952
rect 5055 15921 5550 15941
rect 5055 15903 5101 15921
rect 5055 15869 5061 15903
rect 5095 15869 5101 15903
rect 2466 15688 3837 15722
rect 2466 15555 2500 15688
rect 2658 15555 2692 15688
rect 2850 15555 2884 15688
rect 3042 15555 3076 15688
rect 3234 15555 3268 15688
rect 3426 15555 3460 15688
rect 3671 15598 3681 15650
rect 3733 15598 3743 15650
rect 3679 15597 3691 15598
rect 3725 15597 3737 15598
rect 3679 15591 3737 15597
rect 3534 15562 3580 15585
rect 2460 15520 2506 15555
rect 2460 15486 2466 15520
rect 2500 15486 2506 15520
rect 2460 15451 2506 15486
rect 2556 15520 2602 15555
rect 2556 15486 2562 15520
rect 2596 15486 2602 15520
rect 2556 15451 2602 15486
rect 2652 15520 2698 15555
rect 2652 15486 2658 15520
rect 2692 15486 2698 15520
rect 2652 15451 2698 15486
rect 2748 15520 2794 15555
rect 2748 15486 2754 15520
rect 2788 15486 2794 15520
rect 2748 15451 2794 15486
rect 2844 15520 2890 15555
rect 2844 15486 2850 15520
rect 2884 15486 2890 15520
rect 2844 15451 2890 15486
rect 2940 15520 2986 15555
rect 2940 15486 2946 15520
rect 2980 15486 2986 15520
rect 2940 15451 2986 15486
rect 3036 15520 3082 15555
rect 3036 15486 3042 15520
rect 3076 15486 3082 15520
rect 3036 15451 3082 15486
rect 3132 15520 3178 15555
rect 3132 15486 3138 15520
rect 3172 15486 3178 15520
rect 3132 15451 3178 15486
rect 3228 15520 3274 15555
rect 3228 15486 3234 15520
rect 3268 15486 3274 15520
rect 3228 15451 3274 15486
rect 3324 15520 3370 15555
rect 3324 15486 3330 15520
rect 3364 15486 3370 15520
rect 3324 15451 3370 15486
rect 3420 15520 3466 15555
rect 3420 15486 3426 15520
rect 3460 15486 3466 15520
rect 3420 15451 3466 15486
rect 3534 15528 3540 15562
rect 3574 15560 3580 15562
rect 3803 15560 3837 15688
rect 3574 15559 3680 15560
rect 3734 15559 3837 15560
rect 3574 15547 3687 15559
rect 3574 15528 3647 15547
rect 3534 15490 3647 15528
rect 3534 15456 3540 15490
rect 3574 15471 3647 15490
rect 3681 15471 3687 15547
rect 3574 15460 3687 15471
rect 3574 15456 3580 15460
rect 3641 15459 3687 15460
rect 3729 15547 3837 15559
rect 3987 15722 4021 15863
rect 4179 15722 4213 15863
rect 4371 15722 4405 15863
rect 4563 15722 4597 15863
rect 4755 15722 4789 15863
rect 4947 15722 4981 15863
rect 5055 15825 5101 15869
rect 5683 15776 5743 17029
rect 5177 15742 5743 15776
rect 5177 15722 5211 15742
rect 3987 15688 5211 15722
rect 3987 15555 4021 15688
rect 4179 15555 4213 15688
rect 4371 15555 4405 15688
rect 4563 15555 4597 15688
rect 4755 15555 4789 15688
rect 4947 15555 4981 15688
rect 5438 15684 5512 15685
rect 5326 15682 5400 15683
rect 5326 15630 5337 15682
rect 5389 15630 5400 15682
rect 5438 15632 5449 15684
rect 5501 15632 5512 15684
rect 5438 15631 5512 15632
rect 5326 15629 5400 15630
rect 5055 15562 5101 15585
rect 3729 15471 3735 15547
rect 3769 15471 3837 15547
rect 3729 15460 3837 15471
rect 3729 15459 3775 15460
rect 2450 15420 2516 15423
rect 2447 15368 2457 15420
rect 2509 15368 2519 15420
rect 2450 15363 2516 15368
rect 2562 15311 2596 15451
rect 2642 15420 2708 15423
rect 2638 15368 2648 15420
rect 2700 15368 2710 15420
rect 2642 15363 2708 15368
rect 2754 15311 2788 15451
rect 2834 15420 2900 15423
rect 2830 15368 2840 15420
rect 2892 15368 2902 15420
rect 2834 15363 2900 15368
rect 2946 15311 2980 15451
rect 3026 15420 3092 15423
rect 3022 15368 3032 15420
rect 3084 15368 3094 15420
rect 3026 15363 3092 15368
rect 3138 15311 3172 15451
rect 3218 15419 3284 15423
rect 3215 15367 3225 15419
rect 3277 15367 3287 15419
rect 3218 15363 3284 15367
rect 3330 15311 3364 15451
rect 3410 15419 3476 15423
rect 3407 15367 3417 15419
rect 3469 15367 3479 15419
rect 3534 15418 3580 15456
rect 3534 15384 3540 15418
rect 3574 15384 3580 15418
rect 3410 15363 3476 15367
rect 2282 15277 3364 15311
rect 3534 15201 3580 15384
rect 3803 15311 3837 15460
rect 3981 15520 4027 15555
rect 3981 15486 3987 15520
rect 4021 15486 4027 15520
rect 3981 15451 4027 15486
rect 4077 15520 4123 15555
rect 4077 15486 4083 15520
rect 4117 15486 4123 15520
rect 4077 15451 4123 15486
rect 4173 15520 4219 15555
rect 4173 15486 4179 15520
rect 4213 15486 4219 15520
rect 4173 15451 4219 15486
rect 4269 15520 4315 15555
rect 4269 15486 4275 15520
rect 4309 15486 4315 15520
rect 4269 15451 4315 15486
rect 4365 15520 4411 15555
rect 4365 15486 4371 15520
rect 4405 15486 4411 15520
rect 4365 15451 4411 15486
rect 4461 15520 4507 15555
rect 4461 15486 4467 15520
rect 4501 15486 4507 15520
rect 4461 15451 4507 15486
rect 4557 15520 4603 15555
rect 4557 15486 4563 15520
rect 4597 15486 4603 15520
rect 4557 15451 4603 15486
rect 4653 15520 4699 15555
rect 4653 15486 4659 15520
rect 4693 15486 4699 15520
rect 4653 15451 4699 15486
rect 4749 15520 4795 15555
rect 4749 15486 4755 15520
rect 4789 15486 4795 15520
rect 4749 15451 4795 15486
rect 4845 15520 4891 15555
rect 4845 15486 4851 15520
rect 4885 15486 4891 15520
rect 4845 15451 4891 15486
rect 4941 15520 4987 15555
rect 4941 15486 4947 15520
rect 4981 15486 4987 15520
rect 4941 15451 4987 15486
rect 5055 15528 5061 15562
rect 5095 15528 5101 15562
rect 5055 15490 5101 15528
rect 5055 15456 5061 15490
rect 5095 15473 5101 15490
rect 5095 15456 5550 15473
rect 3971 15420 4037 15423
rect 3968 15368 3978 15420
rect 4030 15368 4040 15420
rect 3971 15363 4037 15368
rect 4083 15311 4117 15451
rect 4163 15420 4229 15423
rect 4159 15368 4169 15420
rect 4221 15368 4231 15420
rect 4163 15363 4229 15368
rect 4275 15311 4309 15451
rect 4355 15420 4421 15423
rect 4351 15368 4361 15420
rect 4413 15368 4423 15420
rect 4355 15363 4421 15368
rect 4467 15311 4501 15451
rect 4547 15420 4613 15423
rect 4543 15368 4553 15420
rect 4605 15368 4615 15420
rect 4547 15363 4613 15368
rect 4659 15311 4693 15451
rect 4739 15419 4805 15423
rect 4736 15367 4746 15419
rect 4798 15367 4808 15419
rect 4739 15363 4805 15367
rect 4851 15311 4885 15451
rect 5055 15442 5550 15456
rect 4931 15419 4997 15423
rect 4928 15367 4938 15419
rect 4990 15367 5000 15419
rect 5055 15418 5303 15442
rect 5055 15384 5061 15418
rect 5095 15408 5303 15418
rect 5337 15408 5395 15442
rect 5429 15408 5487 15442
rect 5521 15408 5550 15442
rect 5095 15384 5550 15408
rect 5055 15377 5550 15384
rect 4931 15363 4997 15367
rect 3803 15277 4885 15311
rect 5055 15202 5101 15377
rect 129 14994 1211 15028
rect 129 14431 163 14994
rect 294 14884 304 14936
rect 356 14884 366 14936
rect 409 14844 443 14994
rect 487 14884 497 14936
rect 549 14884 559 14936
rect 601 14844 635 14994
rect 678 14884 688 14936
rect 740 14884 750 14936
rect 793 14844 827 14994
rect 870 14884 880 14936
rect 932 14884 942 14936
rect 985 14844 1019 14994
rect 1062 14884 1072 14936
rect 1124 14884 1134 14936
rect 1177 14844 1211 14994
rect 1254 14884 1264 14936
rect 1316 14884 1326 14936
rect 1381 14900 1427 15064
rect 2282 14998 3364 15032
rect 1381 14866 1387 14900
rect 1421 14866 1427 14900
rect 1512 14877 1522 14937
rect 1578 14877 1792 14937
rect 1852 14877 1862 14937
rect 307 14797 353 14844
rect 307 14763 313 14797
rect 347 14763 353 14797
rect 307 14725 353 14763
rect 307 14691 313 14725
rect 347 14691 353 14725
rect 307 14653 353 14691
rect 307 14619 313 14653
rect 347 14619 353 14653
rect 307 14572 353 14619
rect 403 14797 449 14844
rect 403 14763 409 14797
rect 443 14763 449 14797
rect 403 14725 449 14763
rect 403 14691 409 14725
rect 443 14691 449 14725
rect 403 14653 449 14691
rect 403 14619 409 14653
rect 443 14619 449 14653
rect 403 14572 449 14619
rect 499 14797 545 14844
rect 499 14763 505 14797
rect 539 14763 545 14797
rect 499 14725 545 14763
rect 499 14691 505 14725
rect 539 14691 545 14725
rect 499 14653 545 14691
rect 499 14619 505 14653
rect 539 14619 545 14653
rect 499 14572 545 14619
rect 595 14797 641 14844
rect 595 14763 601 14797
rect 635 14763 641 14797
rect 595 14725 641 14763
rect 595 14691 601 14725
rect 635 14691 641 14725
rect 595 14653 641 14691
rect 595 14619 601 14653
rect 635 14619 641 14653
rect 595 14572 641 14619
rect 691 14797 737 14844
rect 691 14763 697 14797
rect 731 14763 737 14797
rect 691 14725 737 14763
rect 691 14691 697 14725
rect 731 14691 737 14725
rect 691 14653 737 14691
rect 691 14619 697 14653
rect 731 14619 737 14653
rect 691 14572 737 14619
rect 787 14797 833 14844
rect 787 14763 793 14797
rect 827 14763 833 14797
rect 787 14725 833 14763
rect 787 14691 793 14725
rect 827 14691 833 14725
rect 787 14653 833 14691
rect 787 14619 793 14653
rect 827 14619 833 14653
rect 787 14572 833 14619
rect 883 14797 929 14844
rect 883 14763 889 14797
rect 923 14763 929 14797
rect 883 14725 929 14763
rect 883 14691 889 14725
rect 923 14691 929 14725
rect 883 14653 929 14691
rect 883 14619 889 14653
rect 923 14619 929 14653
rect 883 14572 929 14619
rect 979 14797 1025 14844
rect 979 14763 985 14797
rect 1019 14763 1025 14797
rect 979 14725 1025 14763
rect 979 14691 985 14725
rect 1019 14691 1025 14725
rect 979 14653 1025 14691
rect 979 14619 985 14653
rect 1019 14619 1025 14653
rect 979 14572 1025 14619
rect 1075 14797 1121 14844
rect 1075 14763 1081 14797
rect 1115 14763 1121 14797
rect 1075 14725 1121 14763
rect 1075 14691 1081 14725
rect 1115 14691 1121 14725
rect 1075 14653 1121 14691
rect 1075 14619 1081 14653
rect 1115 14619 1121 14653
rect 1075 14572 1121 14619
rect 1171 14797 1217 14844
rect 1171 14763 1177 14797
rect 1211 14763 1217 14797
rect 1171 14725 1217 14763
rect 1171 14691 1177 14725
rect 1211 14691 1217 14725
rect 1171 14653 1217 14691
rect 1171 14619 1177 14653
rect 1211 14619 1217 14653
rect 1171 14572 1217 14619
rect 1267 14797 1313 14844
rect 1267 14763 1273 14797
rect 1307 14763 1313 14797
rect 1267 14725 1313 14763
rect 1267 14691 1273 14725
rect 1307 14691 1313 14725
rect 1267 14653 1313 14691
rect 1267 14619 1273 14653
rect 1307 14619 1313 14653
rect 1267 14572 1313 14619
rect 1381 14828 1427 14866
rect 1381 14794 1387 14828
rect 1421 14794 1427 14828
rect 1381 14756 1427 14794
rect 1381 14722 1387 14756
rect 1421 14722 1427 14756
rect 1381 14684 1427 14722
rect 1381 14650 1387 14684
rect 1421 14650 1427 14684
rect 1381 14640 1427 14650
rect 1381 14638 2160 14640
rect 1381 14612 2056 14638
rect 1381 14587 1387 14612
rect 1380 14578 1387 14587
rect 1421 14578 2056 14612
rect 0 14397 163 14431
rect 129 14020 163 14397
rect 313 14431 347 14572
rect 505 14431 539 14572
rect 697 14431 731 14572
rect 889 14431 923 14572
rect 1081 14431 1115 14572
rect 1273 14431 1307 14572
rect 1380 14530 2056 14578
rect 2190 14530 2200 14638
rect 1380 14528 2160 14530
rect 2282 14435 2316 14998
rect 2447 14888 2457 14940
rect 2509 14888 2519 14940
rect 2562 14848 2596 14998
rect 2640 14888 2650 14940
rect 2702 14888 2712 14940
rect 2754 14848 2788 14998
rect 2831 14888 2841 14940
rect 2893 14888 2903 14940
rect 2946 14848 2980 14998
rect 3023 14888 3033 14940
rect 3085 14888 3095 14940
rect 3138 14848 3172 14998
rect 3215 14888 3225 14940
rect 3277 14888 3287 14940
rect 3330 14848 3364 14998
rect 3407 14888 3417 14940
rect 3469 14888 3479 14940
rect 3534 14904 3580 15112
rect 3534 14870 3540 14904
rect 3574 14870 3580 14904
rect 2460 14801 2506 14848
rect 2460 14767 2466 14801
rect 2500 14767 2506 14801
rect 2460 14729 2506 14767
rect 2460 14695 2466 14729
rect 2500 14695 2506 14729
rect 2460 14657 2506 14695
rect 2460 14623 2466 14657
rect 2500 14623 2506 14657
rect 2460 14576 2506 14623
rect 2556 14801 2602 14848
rect 2556 14767 2562 14801
rect 2596 14767 2602 14801
rect 2556 14729 2602 14767
rect 2556 14695 2562 14729
rect 2596 14695 2602 14729
rect 2556 14657 2602 14695
rect 2556 14623 2562 14657
rect 2596 14623 2602 14657
rect 2556 14576 2602 14623
rect 2652 14801 2698 14848
rect 2652 14767 2658 14801
rect 2692 14767 2698 14801
rect 2652 14729 2698 14767
rect 2652 14695 2658 14729
rect 2692 14695 2698 14729
rect 2652 14657 2698 14695
rect 2652 14623 2658 14657
rect 2692 14623 2698 14657
rect 2652 14576 2698 14623
rect 2748 14801 2794 14848
rect 2748 14767 2754 14801
rect 2788 14767 2794 14801
rect 2748 14729 2794 14767
rect 2748 14695 2754 14729
rect 2788 14695 2794 14729
rect 2748 14657 2794 14695
rect 2748 14623 2754 14657
rect 2788 14623 2794 14657
rect 2748 14576 2794 14623
rect 2844 14801 2890 14848
rect 2844 14767 2850 14801
rect 2884 14767 2890 14801
rect 2844 14729 2890 14767
rect 2844 14695 2850 14729
rect 2884 14695 2890 14729
rect 2844 14657 2890 14695
rect 2844 14623 2850 14657
rect 2884 14623 2890 14657
rect 2844 14576 2890 14623
rect 2940 14801 2986 14848
rect 2940 14767 2946 14801
rect 2980 14767 2986 14801
rect 2940 14729 2986 14767
rect 2940 14695 2946 14729
rect 2980 14695 2986 14729
rect 2940 14657 2986 14695
rect 2940 14623 2946 14657
rect 2980 14623 2986 14657
rect 2940 14576 2986 14623
rect 3036 14801 3082 14848
rect 3036 14767 3042 14801
rect 3076 14767 3082 14801
rect 3036 14729 3082 14767
rect 3036 14695 3042 14729
rect 3076 14695 3082 14729
rect 3036 14657 3082 14695
rect 3036 14623 3042 14657
rect 3076 14623 3082 14657
rect 3036 14576 3082 14623
rect 3132 14801 3178 14848
rect 3132 14767 3138 14801
rect 3172 14767 3178 14801
rect 3132 14729 3178 14767
rect 3132 14695 3138 14729
rect 3172 14695 3178 14729
rect 3132 14657 3178 14695
rect 3132 14623 3138 14657
rect 3172 14623 3178 14657
rect 3132 14576 3178 14623
rect 3228 14801 3274 14848
rect 3228 14767 3234 14801
rect 3268 14767 3274 14801
rect 3228 14729 3274 14767
rect 3228 14695 3234 14729
rect 3268 14695 3274 14729
rect 3228 14657 3274 14695
rect 3228 14623 3234 14657
rect 3268 14623 3274 14657
rect 3228 14576 3274 14623
rect 3324 14801 3370 14848
rect 3324 14767 3330 14801
rect 3364 14767 3370 14801
rect 3324 14729 3370 14767
rect 3324 14695 3330 14729
rect 3364 14695 3370 14729
rect 3324 14657 3370 14695
rect 3324 14623 3330 14657
rect 3364 14623 3370 14657
rect 3324 14576 3370 14623
rect 3420 14801 3466 14848
rect 3420 14767 3426 14801
rect 3460 14767 3466 14801
rect 3420 14729 3466 14767
rect 3420 14695 3426 14729
rect 3460 14695 3466 14729
rect 3420 14657 3466 14695
rect 3420 14623 3426 14657
rect 3460 14623 3466 14657
rect 3420 14576 3466 14623
rect 3534 14832 3580 14870
rect 3534 14798 3540 14832
rect 3574 14798 3580 14832
rect 3534 14760 3580 14798
rect 3534 14726 3540 14760
rect 3574 14726 3580 14760
rect 3534 14688 3580 14726
rect 3534 14654 3540 14688
rect 3574 14654 3580 14688
rect 3534 14616 3580 14654
rect 3534 14582 3540 14616
rect 3574 14582 3580 14616
rect 2101 14431 2316 14435
rect 313 14401 2316 14431
rect 313 14397 2141 14401
rect 313 14264 347 14397
rect 505 14264 539 14397
rect 697 14264 731 14397
rect 889 14264 923 14397
rect 1081 14264 1115 14397
rect 1273 14264 1307 14397
rect 1381 14271 1608 14294
rect 307 14229 353 14264
rect 307 14195 313 14229
rect 347 14195 353 14229
rect 307 14160 353 14195
rect 403 14229 449 14264
rect 403 14195 409 14229
rect 443 14195 449 14229
rect 403 14160 449 14195
rect 499 14229 545 14264
rect 499 14195 505 14229
rect 539 14195 545 14229
rect 499 14160 545 14195
rect 595 14229 641 14264
rect 595 14195 601 14229
rect 635 14195 641 14229
rect 595 14160 641 14195
rect 691 14229 737 14264
rect 691 14195 697 14229
rect 731 14195 737 14229
rect 691 14160 737 14195
rect 787 14229 833 14264
rect 787 14195 793 14229
rect 827 14195 833 14229
rect 787 14160 833 14195
rect 883 14229 929 14264
rect 883 14195 889 14229
rect 923 14195 929 14229
rect 883 14160 929 14195
rect 979 14229 1025 14264
rect 979 14195 985 14229
rect 1019 14195 1025 14229
rect 979 14160 1025 14195
rect 1075 14229 1121 14264
rect 1075 14195 1081 14229
rect 1115 14195 1121 14229
rect 1075 14160 1121 14195
rect 1171 14229 1217 14264
rect 1171 14195 1177 14229
rect 1211 14195 1217 14229
rect 1171 14160 1217 14195
rect 1267 14229 1313 14264
rect 1267 14195 1273 14229
rect 1307 14195 1313 14229
rect 1267 14160 1313 14195
rect 1381 14237 1387 14271
rect 1421 14237 1608 14271
rect 1381 14199 1608 14237
rect 1381 14165 1387 14199
rect 1421 14174 1608 14199
rect 1421 14165 1427 14174
rect 1560 14172 1608 14174
rect 1598 14170 1608 14172
rect 1720 14170 1730 14294
rect 297 14129 363 14132
rect 294 14077 304 14129
rect 356 14077 366 14129
rect 297 14072 363 14077
rect 409 14020 443 14160
rect 489 14129 555 14132
rect 485 14077 495 14129
rect 547 14077 557 14129
rect 489 14072 555 14077
rect 601 14020 635 14160
rect 681 14129 747 14132
rect 677 14077 687 14129
rect 739 14077 749 14129
rect 681 14072 747 14077
rect 793 14020 827 14160
rect 873 14129 939 14132
rect 869 14077 879 14129
rect 931 14077 941 14129
rect 873 14072 939 14077
rect 985 14020 1019 14160
rect 1065 14128 1131 14132
rect 1062 14076 1072 14128
rect 1124 14076 1134 14128
rect 1065 14072 1131 14076
rect 1177 14020 1211 14160
rect 1257 14128 1323 14132
rect 1254 14076 1264 14128
rect 1316 14076 1326 14128
rect 1381 14127 1427 14165
rect 1920 14132 1930 14134
rect 1381 14093 1387 14127
rect 1421 14093 1427 14127
rect 1257 14072 1323 14076
rect 129 13986 1211 14020
rect 1381 13950 1427 14093
rect 1458 14076 1468 14132
rect 1524 14078 1930 14132
rect 1986 14078 1996 14134
rect 1524 14076 1986 14078
rect 2282 14024 2316 14401
rect 2466 14435 2500 14576
rect 2658 14435 2692 14576
rect 2850 14435 2884 14576
rect 3042 14435 3076 14576
rect 3234 14435 3268 14576
rect 3426 14435 3460 14576
rect 3534 14538 3580 14582
rect 3803 14998 4885 15032
rect 3803 14435 3837 14998
rect 3968 14888 3978 14940
rect 4030 14888 4040 14940
rect 4083 14848 4117 14998
rect 4161 14888 4171 14940
rect 4223 14888 4233 14940
rect 4275 14848 4309 14998
rect 4352 14888 4362 14940
rect 4414 14888 4424 14940
rect 4467 14848 4501 14998
rect 4544 14888 4554 14940
rect 4606 14888 4616 14940
rect 4659 14848 4693 14998
rect 4736 14888 4746 14940
rect 4798 14888 4808 14940
rect 4851 14848 4885 14998
rect 4928 14888 4938 14940
rect 4990 14888 5000 14940
rect 5055 14904 5101 15109
rect 5055 14870 5061 14904
rect 5095 14870 5101 14904
rect 3981 14801 4027 14848
rect 3981 14767 3987 14801
rect 4021 14767 4027 14801
rect 3981 14729 4027 14767
rect 3981 14695 3987 14729
rect 4021 14695 4027 14729
rect 3981 14657 4027 14695
rect 3981 14623 3987 14657
rect 4021 14623 4027 14657
rect 3981 14576 4027 14623
rect 4077 14801 4123 14848
rect 4077 14767 4083 14801
rect 4117 14767 4123 14801
rect 4077 14729 4123 14767
rect 4077 14695 4083 14729
rect 4117 14695 4123 14729
rect 4077 14657 4123 14695
rect 4077 14623 4083 14657
rect 4117 14623 4123 14657
rect 4077 14576 4123 14623
rect 4173 14801 4219 14848
rect 4173 14767 4179 14801
rect 4213 14767 4219 14801
rect 4173 14729 4219 14767
rect 4173 14695 4179 14729
rect 4213 14695 4219 14729
rect 4173 14657 4219 14695
rect 4173 14623 4179 14657
rect 4213 14623 4219 14657
rect 4173 14576 4219 14623
rect 4269 14801 4315 14848
rect 4269 14767 4275 14801
rect 4309 14767 4315 14801
rect 4269 14729 4315 14767
rect 4269 14695 4275 14729
rect 4309 14695 4315 14729
rect 4269 14657 4315 14695
rect 4269 14623 4275 14657
rect 4309 14623 4315 14657
rect 4269 14576 4315 14623
rect 4365 14801 4411 14848
rect 4365 14767 4371 14801
rect 4405 14767 4411 14801
rect 4365 14729 4411 14767
rect 4365 14695 4371 14729
rect 4405 14695 4411 14729
rect 4365 14657 4411 14695
rect 4365 14623 4371 14657
rect 4405 14623 4411 14657
rect 4365 14576 4411 14623
rect 4461 14801 4507 14848
rect 4461 14767 4467 14801
rect 4501 14767 4507 14801
rect 4461 14729 4507 14767
rect 4461 14695 4467 14729
rect 4501 14695 4507 14729
rect 4461 14657 4507 14695
rect 4461 14623 4467 14657
rect 4501 14623 4507 14657
rect 4461 14576 4507 14623
rect 4557 14801 4603 14848
rect 4557 14767 4563 14801
rect 4597 14767 4603 14801
rect 4557 14729 4603 14767
rect 4557 14695 4563 14729
rect 4597 14695 4603 14729
rect 4557 14657 4603 14695
rect 4557 14623 4563 14657
rect 4597 14623 4603 14657
rect 4557 14576 4603 14623
rect 4653 14801 4699 14848
rect 4653 14767 4659 14801
rect 4693 14767 4699 14801
rect 4653 14729 4699 14767
rect 4653 14695 4659 14729
rect 4693 14695 4699 14729
rect 4653 14657 4699 14695
rect 4653 14623 4659 14657
rect 4693 14623 4699 14657
rect 4653 14576 4699 14623
rect 4749 14801 4795 14848
rect 4749 14767 4755 14801
rect 4789 14767 4795 14801
rect 4749 14729 4795 14767
rect 4749 14695 4755 14729
rect 4789 14695 4795 14729
rect 4749 14657 4795 14695
rect 4749 14623 4755 14657
rect 4789 14623 4795 14657
rect 4749 14576 4795 14623
rect 4845 14801 4891 14848
rect 4845 14767 4851 14801
rect 4885 14767 4891 14801
rect 4845 14729 4891 14767
rect 4845 14695 4851 14729
rect 4885 14695 4891 14729
rect 4845 14657 4891 14695
rect 4845 14623 4851 14657
rect 4885 14623 4891 14657
rect 4845 14576 4891 14623
rect 4941 14801 4987 14848
rect 4941 14767 4947 14801
rect 4981 14767 4987 14801
rect 4941 14729 4987 14767
rect 4941 14695 4947 14729
rect 4981 14695 4987 14729
rect 4941 14657 4987 14695
rect 4941 14623 4947 14657
rect 4981 14623 4987 14657
rect 4941 14576 4987 14623
rect 5055 14832 5101 14870
rect 5055 14798 5061 14832
rect 5095 14798 5101 14832
rect 5055 14760 5101 14798
rect 5055 14726 5061 14760
rect 5095 14729 5101 14760
rect 5274 14729 5550 14730
rect 5095 14726 5550 14729
rect 5055 14699 5550 14726
rect 5055 14688 5303 14699
rect 5055 14654 5061 14688
rect 5095 14665 5303 14688
rect 5337 14665 5395 14699
rect 5429 14665 5487 14699
rect 5521 14665 5550 14699
rect 5095 14654 5550 14665
rect 5055 14634 5550 14654
rect 5055 14616 5101 14634
rect 5055 14582 5061 14616
rect 5095 14582 5101 14616
rect 2466 14401 3837 14435
rect 2466 14268 2500 14401
rect 2658 14268 2692 14401
rect 2850 14268 2884 14401
rect 3042 14268 3076 14401
rect 3234 14268 3268 14401
rect 3426 14268 3460 14401
rect 3671 14311 3681 14363
rect 3733 14311 3743 14363
rect 3679 14310 3691 14311
rect 3725 14310 3737 14311
rect 3679 14304 3737 14310
rect 3534 14275 3580 14298
rect 2460 14233 2506 14268
rect 2460 14199 2466 14233
rect 2500 14199 2506 14233
rect 2460 14164 2506 14199
rect 2556 14233 2602 14268
rect 2556 14199 2562 14233
rect 2596 14199 2602 14233
rect 2556 14164 2602 14199
rect 2652 14233 2698 14268
rect 2652 14199 2658 14233
rect 2692 14199 2698 14233
rect 2652 14164 2698 14199
rect 2748 14233 2794 14268
rect 2748 14199 2754 14233
rect 2788 14199 2794 14233
rect 2748 14164 2794 14199
rect 2844 14233 2890 14268
rect 2844 14199 2850 14233
rect 2884 14199 2890 14233
rect 2844 14164 2890 14199
rect 2940 14233 2986 14268
rect 2940 14199 2946 14233
rect 2980 14199 2986 14233
rect 2940 14164 2986 14199
rect 3036 14233 3082 14268
rect 3036 14199 3042 14233
rect 3076 14199 3082 14233
rect 3036 14164 3082 14199
rect 3132 14233 3178 14268
rect 3132 14199 3138 14233
rect 3172 14199 3178 14233
rect 3132 14164 3178 14199
rect 3228 14233 3274 14268
rect 3228 14199 3234 14233
rect 3268 14199 3274 14233
rect 3228 14164 3274 14199
rect 3324 14233 3370 14268
rect 3324 14199 3330 14233
rect 3364 14199 3370 14233
rect 3324 14164 3370 14199
rect 3420 14233 3466 14268
rect 3420 14199 3426 14233
rect 3460 14199 3466 14233
rect 3420 14164 3466 14199
rect 3534 14241 3540 14275
rect 3574 14273 3580 14275
rect 3803 14273 3837 14401
rect 3574 14272 3680 14273
rect 3734 14272 3837 14273
rect 3574 14260 3687 14272
rect 3574 14241 3647 14260
rect 3534 14203 3647 14241
rect 3534 14169 3540 14203
rect 3574 14184 3647 14203
rect 3681 14184 3687 14260
rect 3574 14173 3687 14184
rect 3574 14169 3580 14173
rect 3641 14172 3687 14173
rect 3729 14260 3837 14272
rect 3987 14435 4021 14576
rect 4179 14435 4213 14576
rect 4371 14435 4405 14576
rect 4563 14435 4597 14576
rect 4755 14435 4789 14576
rect 4947 14435 4981 14576
rect 5055 14538 5101 14582
rect 5683 14489 5743 15742
rect 5177 14455 5743 14489
rect 5177 14435 5211 14455
rect 3987 14401 5211 14435
rect 3987 14268 4021 14401
rect 4179 14268 4213 14401
rect 4371 14268 4405 14401
rect 4563 14268 4597 14401
rect 4755 14268 4789 14401
rect 4947 14268 4981 14401
rect 5438 14397 5512 14398
rect 5326 14395 5400 14396
rect 5326 14343 5337 14395
rect 5389 14343 5400 14395
rect 5438 14345 5449 14397
rect 5501 14345 5512 14397
rect 5438 14344 5512 14345
rect 5326 14342 5400 14343
rect 5055 14275 5101 14298
rect 3729 14184 3735 14260
rect 3769 14184 3837 14260
rect 3729 14173 3837 14184
rect 3729 14172 3775 14173
rect 2450 14133 2516 14136
rect 2447 14081 2457 14133
rect 2509 14081 2519 14133
rect 2450 14076 2516 14081
rect 2562 14024 2596 14164
rect 2642 14133 2708 14136
rect 2638 14081 2648 14133
rect 2700 14081 2710 14133
rect 2642 14076 2708 14081
rect 2754 14024 2788 14164
rect 2834 14133 2900 14136
rect 2830 14081 2840 14133
rect 2892 14081 2902 14133
rect 2834 14076 2900 14081
rect 2946 14024 2980 14164
rect 3026 14133 3092 14136
rect 3022 14081 3032 14133
rect 3084 14081 3094 14133
rect 3026 14076 3092 14081
rect 3138 14024 3172 14164
rect 3218 14132 3284 14136
rect 3215 14080 3225 14132
rect 3277 14080 3287 14132
rect 3218 14076 3284 14080
rect 3330 14024 3364 14164
rect 3410 14132 3476 14136
rect 3407 14080 3417 14132
rect 3469 14080 3479 14132
rect 3534 14131 3580 14169
rect 3534 14097 3540 14131
rect 3574 14097 3580 14131
rect 3410 14076 3476 14080
rect 2282 13990 3364 14024
rect 3534 13914 3580 14097
rect 3803 14024 3837 14173
rect 3981 14233 4027 14268
rect 3981 14199 3987 14233
rect 4021 14199 4027 14233
rect 3981 14164 4027 14199
rect 4077 14233 4123 14268
rect 4077 14199 4083 14233
rect 4117 14199 4123 14233
rect 4077 14164 4123 14199
rect 4173 14233 4219 14268
rect 4173 14199 4179 14233
rect 4213 14199 4219 14233
rect 4173 14164 4219 14199
rect 4269 14233 4315 14268
rect 4269 14199 4275 14233
rect 4309 14199 4315 14233
rect 4269 14164 4315 14199
rect 4365 14233 4411 14268
rect 4365 14199 4371 14233
rect 4405 14199 4411 14233
rect 4365 14164 4411 14199
rect 4461 14233 4507 14268
rect 4461 14199 4467 14233
rect 4501 14199 4507 14233
rect 4461 14164 4507 14199
rect 4557 14233 4603 14268
rect 4557 14199 4563 14233
rect 4597 14199 4603 14233
rect 4557 14164 4603 14199
rect 4653 14233 4699 14268
rect 4653 14199 4659 14233
rect 4693 14199 4699 14233
rect 4653 14164 4699 14199
rect 4749 14233 4795 14268
rect 4749 14199 4755 14233
rect 4789 14199 4795 14233
rect 4749 14164 4795 14199
rect 4845 14233 4891 14268
rect 4845 14199 4851 14233
rect 4885 14199 4891 14233
rect 4845 14164 4891 14199
rect 4941 14233 4987 14268
rect 4941 14199 4947 14233
rect 4981 14199 4987 14233
rect 4941 14164 4987 14199
rect 5055 14241 5061 14275
rect 5095 14241 5101 14275
rect 5055 14203 5101 14241
rect 5055 14169 5061 14203
rect 5095 14186 5101 14203
rect 5095 14169 5550 14186
rect 3971 14133 4037 14136
rect 3968 14081 3978 14133
rect 4030 14081 4040 14133
rect 3971 14076 4037 14081
rect 4083 14024 4117 14164
rect 4163 14133 4229 14136
rect 4159 14081 4169 14133
rect 4221 14081 4231 14133
rect 4163 14076 4229 14081
rect 4275 14024 4309 14164
rect 4355 14133 4421 14136
rect 4351 14081 4361 14133
rect 4413 14081 4423 14133
rect 4355 14076 4421 14081
rect 4467 14024 4501 14164
rect 4547 14133 4613 14136
rect 4543 14081 4553 14133
rect 4605 14081 4615 14133
rect 4547 14076 4613 14081
rect 4659 14024 4693 14164
rect 4739 14132 4805 14136
rect 4736 14080 4746 14132
rect 4798 14080 4808 14132
rect 4739 14076 4805 14080
rect 4851 14024 4885 14164
rect 5055 14155 5550 14169
rect 4931 14132 4997 14136
rect 4928 14080 4938 14132
rect 4990 14080 5000 14132
rect 5055 14131 5303 14155
rect 5055 14097 5061 14131
rect 5095 14121 5303 14131
rect 5337 14121 5395 14155
rect 5429 14121 5487 14155
rect 5521 14121 5550 14155
rect 5095 14097 5550 14121
rect 5055 14090 5550 14097
rect 4931 14076 4997 14080
rect 3803 13990 4885 14024
rect 5055 13915 5101 14090
rect 129 13707 1211 13741
rect 129 13144 163 13707
rect 294 13597 304 13649
rect 356 13597 366 13649
rect 409 13557 443 13707
rect 487 13597 497 13649
rect 549 13597 559 13649
rect 601 13557 635 13707
rect 678 13597 688 13649
rect 740 13597 750 13649
rect 793 13557 827 13707
rect 870 13597 880 13649
rect 932 13597 942 13649
rect 985 13557 1019 13707
rect 1062 13597 1072 13649
rect 1124 13597 1134 13649
rect 1177 13557 1211 13707
rect 1254 13597 1264 13649
rect 1316 13597 1326 13649
rect 1381 13613 1427 13777
rect 2282 13711 3364 13745
rect 1381 13579 1387 13613
rect 1421 13579 1427 13613
rect 1512 13590 1522 13650
rect 1578 13590 1792 13650
rect 1852 13590 1862 13650
rect 307 13510 353 13557
rect 307 13476 313 13510
rect 347 13476 353 13510
rect 307 13438 353 13476
rect 307 13404 313 13438
rect 347 13404 353 13438
rect 307 13366 353 13404
rect 307 13332 313 13366
rect 347 13332 353 13366
rect 307 13285 353 13332
rect 403 13510 449 13557
rect 403 13476 409 13510
rect 443 13476 449 13510
rect 403 13438 449 13476
rect 403 13404 409 13438
rect 443 13404 449 13438
rect 403 13366 449 13404
rect 403 13332 409 13366
rect 443 13332 449 13366
rect 403 13285 449 13332
rect 499 13510 545 13557
rect 499 13476 505 13510
rect 539 13476 545 13510
rect 499 13438 545 13476
rect 499 13404 505 13438
rect 539 13404 545 13438
rect 499 13366 545 13404
rect 499 13332 505 13366
rect 539 13332 545 13366
rect 499 13285 545 13332
rect 595 13510 641 13557
rect 595 13476 601 13510
rect 635 13476 641 13510
rect 595 13438 641 13476
rect 595 13404 601 13438
rect 635 13404 641 13438
rect 595 13366 641 13404
rect 595 13332 601 13366
rect 635 13332 641 13366
rect 595 13285 641 13332
rect 691 13510 737 13557
rect 691 13476 697 13510
rect 731 13476 737 13510
rect 691 13438 737 13476
rect 691 13404 697 13438
rect 731 13404 737 13438
rect 691 13366 737 13404
rect 691 13332 697 13366
rect 731 13332 737 13366
rect 691 13285 737 13332
rect 787 13510 833 13557
rect 787 13476 793 13510
rect 827 13476 833 13510
rect 787 13438 833 13476
rect 787 13404 793 13438
rect 827 13404 833 13438
rect 787 13366 833 13404
rect 787 13332 793 13366
rect 827 13332 833 13366
rect 787 13285 833 13332
rect 883 13510 929 13557
rect 883 13476 889 13510
rect 923 13476 929 13510
rect 883 13438 929 13476
rect 883 13404 889 13438
rect 923 13404 929 13438
rect 883 13366 929 13404
rect 883 13332 889 13366
rect 923 13332 929 13366
rect 883 13285 929 13332
rect 979 13510 1025 13557
rect 979 13476 985 13510
rect 1019 13476 1025 13510
rect 979 13438 1025 13476
rect 979 13404 985 13438
rect 1019 13404 1025 13438
rect 979 13366 1025 13404
rect 979 13332 985 13366
rect 1019 13332 1025 13366
rect 979 13285 1025 13332
rect 1075 13510 1121 13557
rect 1075 13476 1081 13510
rect 1115 13476 1121 13510
rect 1075 13438 1121 13476
rect 1075 13404 1081 13438
rect 1115 13404 1121 13438
rect 1075 13366 1121 13404
rect 1075 13332 1081 13366
rect 1115 13332 1121 13366
rect 1075 13285 1121 13332
rect 1171 13510 1217 13557
rect 1171 13476 1177 13510
rect 1211 13476 1217 13510
rect 1171 13438 1217 13476
rect 1171 13404 1177 13438
rect 1211 13404 1217 13438
rect 1171 13366 1217 13404
rect 1171 13332 1177 13366
rect 1211 13332 1217 13366
rect 1171 13285 1217 13332
rect 1267 13510 1313 13557
rect 1267 13476 1273 13510
rect 1307 13476 1313 13510
rect 1267 13438 1313 13476
rect 1267 13404 1273 13438
rect 1307 13404 1313 13438
rect 1267 13366 1313 13404
rect 1267 13332 1273 13366
rect 1307 13332 1313 13366
rect 1267 13285 1313 13332
rect 1381 13541 1427 13579
rect 1381 13507 1387 13541
rect 1421 13507 1427 13541
rect 1381 13469 1427 13507
rect 1381 13435 1387 13469
rect 1421 13435 1427 13469
rect 1381 13397 1427 13435
rect 1381 13363 1387 13397
rect 1421 13363 1427 13397
rect 1381 13353 1427 13363
rect 1381 13351 2160 13353
rect 1381 13325 2056 13351
rect 1381 13300 1387 13325
rect 1380 13291 1387 13300
rect 1421 13291 2056 13325
rect 0 13110 163 13144
rect 129 12733 163 13110
rect 313 13144 347 13285
rect 505 13144 539 13285
rect 697 13144 731 13285
rect 889 13144 923 13285
rect 1081 13144 1115 13285
rect 1273 13144 1307 13285
rect 1380 13243 2056 13291
rect 2190 13243 2200 13351
rect 1380 13241 2160 13243
rect 2282 13148 2316 13711
rect 2447 13601 2457 13653
rect 2509 13601 2519 13653
rect 2562 13561 2596 13711
rect 2640 13601 2650 13653
rect 2702 13601 2712 13653
rect 2754 13561 2788 13711
rect 2831 13601 2841 13653
rect 2893 13601 2903 13653
rect 2946 13561 2980 13711
rect 3023 13601 3033 13653
rect 3085 13601 3095 13653
rect 3138 13561 3172 13711
rect 3215 13601 3225 13653
rect 3277 13601 3287 13653
rect 3330 13561 3364 13711
rect 3407 13601 3417 13653
rect 3469 13601 3479 13653
rect 3534 13617 3580 13825
rect 3534 13583 3540 13617
rect 3574 13583 3580 13617
rect 2460 13514 2506 13561
rect 2460 13480 2466 13514
rect 2500 13480 2506 13514
rect 2460 13442 2506 13480
rect 2460 13408 2466 13442
rect 2500 13408 2506 13442
rect 2460 13370 2506 13408
rect 2460 13336 2466 13370
rect 2500 13336 2506 13370
rect 2460 13289 2506 13336
rect 2556 13514 2602 13561
rect 2556 13480 2562 13514
rect 2596 13480 2602 13514
rect 2556 13442 2602 13480
rect 2556 13408 2562 13442
rect 2596 13408 2602 13442
rect 2556 13370 2602 13408
rect 2556 13336 2562 13370
rect 2596 13336 2602 13370
rect 2556 13289 2602 13336
rect 2652 13514 2698 13561
rect 2652 13480 2658 13514
rect 2692 13480 2698 13514
rect 2652 13442 2698 13480
rect 2652 13408 2658 13442
rect 2692 13408 2698 13442
rect 2652 13370 2698 13408
rect 2652 13336 2658 13370
rect 2692 13336 2698 13370
rect 2652 13289 2698 13336
rect 2748 13514 2794 13561
rect 2748 13480 2754 13514
rect 2788 13480 2794 13514
rect 2748 13442 2794 13480
rect 2748 13408 2754 13442
rect 2788 13408 2794 13442
rect 2748 13370 2794 13408
rect 2748 13336 2754 13370
rect 2788 13336 2794 13370
rect 2748 13289 2794 13336
rect 2844 13514 2890 13561
rect 2844 13480 2850 13514
rect 2884 13480 2890 13514
rect 2844 13442 2890 13480
rect 2844 13408 2850 13442
rect 2884 13408 2890 13442
rect 2844 13370 2890 13408
rect 2844 13336 2850 13370
rect 2884 13336 2890 13370
rect 2844 13289 2890 13336
rect 2940 13514 2986 13561
rect 2940 13480 2946 13514
rect 2980 13480 2986 13514
rect 2940 13442 2986 13480
rect 2940 13408 2946 13442
rect 2980 13408 2986 13442
rect 2940 13370 2986 13408
rect 2940 13336 2946 13370
rect 2980 13336 2986 13370
rect 2940 13289 2986 13336
rect 3036 13514 3082 13561
rect 3036 13480 3042 13514
rect 3076 13480 3082 13514
rect 3036 13442 3082 13480
rect 3036 13408 3042 13442
rect 3076 13408 3082 13442
rect 3036 13370 3082 13408
rect 3036 13336 3042 13370
rect 3076 13336 3082 13370
rect 3036 13289 3082 13336
rect 3132 13514 3178 13561
rect 3132 13480 3138 13514
rect 3172 13480 3178 13514
rect 3132 13442 3178 13480
rect 3132 13408 3138 13442
rect 3172 13408 3178 13442
rect 3132 13370 3178 13408
rect 3132 13336 3138 13370
rect 3172 13336 3178 13370
rect 3132 13289 3178 13336
rect 3228 13514 3274 13561
rect 3228 13480 3234 13514
rect 3268 13480 3274 13514
rect 3228 13442 3274 13480
rect 3228 13408 3234 13442
rect 3268 13408 3274 13442
rect 3228 13370 3274 13408
rect 3228 13336 3234 13370
rect 3268 13336 3274 13370
rect 3228 13289 3274 13336
rect 3324 13514 3370 13561
rect 3324 13480 3330 13514
rect 3364 13480 3370 13514
rect 3324 13442 3370 13480
rect 3324 13408 3330 13442
rect 3364 13408 3370 13442
rect 3324 13370 3370 13408
rect 3324 13336 3330 13370
rect 3364 13336 3370 13370
rect 3324 13289 3370 13336
rect 3420 13514 3466 13561
rect 3420 13480 3426 13514
rect 3460 13480 3466 13514
rect 3420 13442 3466 13480
rect 3420 13408 3426 13442
rect 3460 13408 3466 13442
rect 3420 13370 3466 13408
rect 3420 13336 3426 13370
rect 3460 13336 3466 13370
rect 3420 13289 3466 13336
rect 3534 13545 3580 13583
rect 3534 13511 3540 13545
rect 3574 13511 3580 13545
rect 3534 13473 3580 13511
rect 3534 13439 3540 13473
rect 3574 13439 3580 13473
rect 3534 13401 3580 13439
rect 3534 13367 3540 13401
rect 3574 13367 3580 13401
rect 3534 13329 3580 13367
rect 3534 13295 3540 13329
rect 3574 13295 3580 13329
rect 2101 13144 2316 13148
rect 313 13114 2316 13144
rect 313 13110 2141 13114
rect 313 12977 347 13110
rect 505 12977 539 13110
rect 697 12977 731 13110
rect 889 12977 923 13110
rect 1081 12977 1115 13110
rect 1273 12977 1307 13110
rect 1381 12984 1608 13007
rect 307 12942 353 12977
rect 307 12908 313 12942
rect 347 12908 353 12942
rect 307 12873 353 12908
rect 403 12942 449 12977
rect 403 12908 409 12942
rect 443 12908 449 12942
rect 403 12873 449 12908
rect 499 12942 545 12977
rect 499 12908 505 12942
rect 539 12908 545 12942
rect 499 12873 545 12908
rect 595 12942 641 12977
rect 595 12908 601 12942
rect 635 12908 641 12942
rect 595 12873 641 12908
rect 691 12942 737 12977
rect 691 12908 697 12942
rect 731 12908 737 12942
rect 691 12873 737 12908
rect 787 12942 833 12977
rect 787 12908 793 12942
rect 827 12908 833 12942
rect 787 12873 833 12908
rect 883 12942 929 12977
rect 883 12908 889 12942
rect 923 12908 929 12942
rect 883 12873 929 12908
rect 979 12942 1025 12977
rect 979 12908 985 12942
rect 1019 12908 1025 12942
rect 979 12873 1025 12908
rect 1075 12942 1121 12977
rect 1075 12908 1081 12942
rect 1115 12908 1121 12942
rect 1075 12873 1121 12908
rect 1171 12942 1217 12977
rect 1171 12908 1177 12942
rect 1211 12908 1217 12942
rect 1171 12873 1217 12908
rect 1267 12942 1313 12977
rect 1267 12908 1273 12942
rect 1307 12908 1313 12942
rect 1267 12873 1313 12908
rect 1381 12950 1387 12984
rect 1421 12950 1608 12984
rect 1381 12912 1608 12950
rect 1381 12878 1387 12912
rect 1421 12887 1608 12912
rect 1421 12878 1427 12887
rect 1560 12885 1608 12887
rect 1598 12883 1608 12885
rect 1720 12883 1730 13007
rect 297 12842 363 12845
rect 294 12790 304 12842
rect 356 12790 366 12842
rect 297 12785 363 12790
rect 409 12733 443 12873
rect 489 12842 555 12845
rect 485 12790 495 12842
rect 547 12790 557 12842
rect 489 12785 555 12790
rect 601 12733 635 12873
rect 681 12842 747 12845
rect 677 12790 687 12842
rect 739 12790 749 12842
rect 681 12785 747 12790
rect 793 12733 827 12873
rect 873 12842 939 12845
rect 869 12790 879 12842
rect 931 12790 941 12842
rect 873 12785 939 12790
rect 985 12733 1019 12873
rect 1065 12841 1131 12845
rect 1062 12789 1072 12841
rect 1124 12789 1134 12841
rect 1065 12785 1131 12789
rect 1177 12733 1211 12873
rect 1257 12841 1323 12845
rect 1254 12789 1264 12841
rect 1316 12789 1326 12841
rect 1381 12840 1427 12878
rect 1920 12845 1930 12847
rect 1381 12806 1387 12840
rect 1421 12806 1427 12840
rect 1257 12785 1323 12789
rect 129 12699 1211 12733
rect 1381 12663 1427 12806
rect 1458 12789 1468 12845
rect 1524 12791 1930 12845
rect 1986 12791 1996 12847
rect 1524 12789 1986 12791
rect 2282 12737 2316 13114
rect 2466 13148 2500 13289
rect 2658 13148 2692 13289
rect 2850 13148 2884 13289
rect 3042 13148 3076 13289
rect 3234 13148 3268 13289
rect 3426 13148 3460 13289
rect 3534 13251 3580 13295
rect 3803 13711 4885 13745
rect 3803 13148 3837 13711
rect 3968 13601 3978 13653
rect 4030 13601 4040 13653
rect 4083 13561 4117 13711
rect 4161 13601 4171 13653
rect 4223 13601 4233 13653
rect 4275 13561 4309 13711
rect 4352 13601 4362 13653
rect 4414 13601 4424 13653
rect 4467 13561 4501 13711
rect 4544 13601 4554 13653
rect 4606 13601 4616 13653
rect 4659 13561 4693 13711
rect 4736 13601 4746 13653
rect 4798 13601 4808 13653
rect 4851 13561 4885 13711
rect 4928 13601 4938 13653
rect 4990 13601 5000 13653
rect 5055 13617 5101 13822
rect 5055 13583 5061 13617
rect 5095 13583 5101 13617
rect 3981 13514 4027 13561
rect 3981 13480 3987 13514
rect 4021 13480 4027 13514
rect 3981 13442 4027 13480
rect 3981 13408 3987 13442
rect 4021 13408 4027 13442
rect 3981 13370 4027 13408
rect 3981 13336 3987 13370
rect 4021 13336 4027 13370
rect 3981 13289 4027 13336
rect 4077 13514 4123 13561
rect 4077 13480 4083 13514
rect 4117 13480 4123 13514
rect 4077 13442 4123 13480
rect 4077 13408 4083 13442
rect 4117 13408 4123 13442
rect 4077 13370 4123 13408
rect 4077 13336 4083 13370
rect 4117 13336 4123 13370
rect 4077 13289 4123 13336
rect 4173 13514 4219 13561
rect 4173 13480 4179 13514
rect 4213 13480 4219 13514
rect 4173 13442 4219 13480
rect 4173 13408 4179 13442
rect 4213 13408 4219 13442
rect 4173 13370 4219 13408
rect 4173 13336 4179 13370
rect 4213 13336 4219 13370
rect 4173 13289 4219 13336
rect 4269 13514 4315 13561
rect 4269 13480 4275 13514
rect 4309 13480 4315 13514
rect 4269 13442 4315 13480
rect 4269 13408 4275 13442
rect 4309 13408 4315 13442
rect 4269 13370 4315 13408
rect 4269 13336 4275 13370
rect 4309 13336 4315 13370
rect 4269 13289 4315 13336
rect 4365 13514 4411 13561
rect 4365 13480 4371 13514
rect 4405 13480 4411 13514
rect 4365 13442 4411 13480
rect 4365 13408 4371 13442
rect 4405 13408 4411 13442
rect 4365 13370 4411 13408
rect 4365 13336 4371 13370
rect 4405 13336 4411 13370
rect 4365 13289 4411 13336
rect 4461 13514 4507 13561
rect 4461 13480 4467 13514
rect 4501 13480 4507 13514
rect 4461 13442 4507 13480
rect 4461 13408 4467 13442
rect 4501 13408 4507 13442
rect 4461 13370 4507 13408
rect 4461 13336 4467 13370
rect 4501 13336 4507 13370
rect 4461 13289 4507 13336
rect 4557 13514 4603 13561
rect 4557 13480 4563 13514
rect 4597 13480 4603 13514
rect 4557 13442 4603 13480
rect 4557 13408 4563 13442
rect 4597 13408 4603 13442
rect 4557 13370 4603 13408
rect 4557 13336 4563 13370
rect 4597 13336 4603 13370
rect 4557 13289 4603 13336
rect 4653 13514 4699 13561
rect 4653 13480 4659 13514
rect 4693 13480 4699 13514
rect 4653 13442 4699 13480
rect 4653 13408 4659 13442
rect 4693 13408 4699 13442
rect 4653 13370 4699 13408
rect 4653 13336 4659 13370
rect 4693 13336 4699 13370
rect 4653 13289 4699 13336
rect 4749 13514 4795 13561
rect 4749 13480 4755 13514
rect 4789 13480 4795 13514
rect 4749 13442 4795 13480
rect 4749 13408 4755 13442
rect 4789 13408 4795 13442
rect 4749 13370 4795 13408
rect 4749 13336 4755 13370
rect 4789 13336 4795 13370
rect 4749 13289 4795 13336
rect 4845 13514 4891 13561
rect 4845 13480 4851 13514
rect 4885 13480 4891 13514
rect 4845 13442 4891 13480
rect 4845 13408 4851 13442
rect 4885 13408 4891 13442
rect 4845 13370 4891 13408
rect 4845 13336 4851 13370
rect 4885 13336 4891 13370
rect 4845 13289 4891 13336
rect 4941 13514 4987 13561
rect 4941 13480 4947 13514
rect 4981 13480 4987 13514
rect 4941 13442 4987 13480
rect 4941 13408 4947 13442
rect 4981 13408 4987 13442
rect 4941 13370 4987 13408
rect 4941 13336 4947 13370
rect 4981 13336 4987 13370
rect 4941 13289 4987 13336
rect 5055 13545 5101 13583
rect 5055 13511 5061 13545
rect 5095 13511 5101 13545
rect 5055 13473 5101 13511
rect 5055 13439 5061 13473
rect 5095 13442 5101 13473
rect 5274 13442 5550 13443
rect 5095 13439 5550 13442
rect 5055 13412 5550 13439
rect 5055 13401 5303 13412
rect 5055 13367 5061 13401
rect 5095 13378 5303 13401
rect 5337 13378 5395 13412
rect 5429 13378 5487 13412
rect 5521 13378 5550 13412
rect 5095 13367 5550 13378
rect 5055 13347 5550 13367
rect 5055 13329 5101 13347
rect 5055 13295 5061 13329
rect 5095 13295 5101 13329
rect 2466 13114 3837 13148
rect 2466 12981 2500 13114
rect 2658 12981 2692 13114
rect 2850 12981 2884 13114
rect 3042 12981 3076 13114
rect 3234 12981 3268 13114
rect 3426 12981 3460 13114
rect 3671 13024 3681 13076
rect 3733 13024 3743 13076
rect 3679 13023 3691 13024
rect 3725 13023 3737 13024
rect 3679 13017 3737 13023
rect 3534 12988 3580 13011
rect 2460 12946 2506 12981
rect 2460 12912 2466 12946
rect 2500 12912 2506 12946
rect 2460 12877 2506 12912
rect 2556 12946 2602 12981
rect 2556 12912 2562 12946
rect 2596 12912 2602 12946
rect 2556 12877 2602 12912
rect 2652 12946 2698 12981
rect 2652 12912 2658 12946
rect 2692 12912 2698 12946
rect 2652 12877 2698 12912
rect 2748 12946 2794 12981
rect 2748 12912 2754 12946
rect 2788 12912 2794 12946
rect 2748 12877 2794 12912
rect 2844 12946 2890 12981
rect 2844 12912 2850 12946
rect 2884 12912 2890 12946
rect 2844 12877 2890 12912
rect 2940 12946 2986 12981
rect 2940 12912 2946 12946
rect 2980 12912 2986 12946
rect 2940 12877 2986 12912
rect 3036 12946 3082 12981
rect 3036 12912 3042 12946
rect 3076 12912 3082 12946
rect 3036 12877 3082 12912
rect 3132 12946 3178 12981
rect 3132 12912 3138 12946
rect 3172 12912 3178 12946
rect 3132 12877 3178 12912
rect 3228 12946 3274 12981
rect 3228 12912 3234 12946
rect 3268 12912 3274 12946
rect 3228 12877 3274 12912
rect 3324 12946 3370 12981
rect 3324 12912 3330 12946
rect 3364 12912 3370 12946
rect 3324 12877 3370 12912
rect 3420 12946 3466 12981
rect 3420 12912 3426 12946
rect 3460 12912 3466 12946
rect 3420 12877 3466 12912
rect 3534 12954 3540 12988
rect 3574 12986 3580 12988
rect 3803 12986 3837 13114
rect 3574 12985 3680 12986
rect 3734 12985 3837 12986
rect 3574 12973 3687 12985
rect 3574 12954 3647 12973
rect 3534 12916 3647 12954
rect 3534 12882 3540 12916
rect 3574 12897 3647 12916
rect 3681 12897 3687 12973
rect 3574 12886 3687 12897
rect 3574 12882 3580 12886
rect 3641 12885 3687 12886
rect 3729 12973 3837 12985
rect 3987 13148 4021 13289
rect 4179 13148 4213 13289
rect 4371 13148 4405 13289
rect 4563 13148 4597 13289
rect 4755 13148 4789 13289
rect 4947 13148 4981 13289
rect 5055 13251 5101 13295
rect 5683 13202 5743 14455
rect 5177 13168 5743 13202
rect 5177 13148 5211 13168
rect 3987 13114 5211 13148
rect 3987 12981 4021 13114
rect 4179 12981 4213 13114
rect 4371 12981 4405 13114
rect 4563 12981 4597 13114
rect 4755 12981 4789 13114
rect 4947 12981 4981 13114
rect 5438 13110 5512 13111
rect 5326 13108 5400 13109
rect 5326 13056 5337 13108
rect 5389 13056 5400 13108
rect 5438 13058 5449 13110
rect 5501 13058 5512 13110
rect 5438 13057 5512 13058
rect 5326 13055 5400 13056
rect 5055 12988 5101 13011
rect 3729 12897 3735 12973
rect 3769 12897 3837 12973
rect 3729 12886 3837 12897
rect 3729 12885 3775 12886
rect 2450 12846 2516 12849
rect 2447 12794 2457 12846
rect 2509 12794 2519 12846
rect 2450 12789 2516 12794
rect 2562 12737 2596 12877
rect 2642 12846 2708 12849
rect 2638 12794 2648 12846
rect 2700 12794 2710 12846
rect 2642 12789 2708 12794
rect 2754 12737 2788 12877
rect 2834 12846 2900 12849
rect 2830 12794 2840 12846
rect 2892 12794 2902 12846
rect 2834 12789 2900 12794
rect 2946 12737 2980 12877
rect 3026 12846 3092 12849
rect 3022 12794 3032 12846
rect 3084 12794 3094 12846
rect 3026 12789 3092 12794
rect 3138 12737 3172 12877
rect 3218 12845 3284 12849
rect 3215 12793 3225 12845
rect 3277 12793 3287 12845
rect 3218 12789 3284 12793
rect 3330 12737 3364 12877
rect 3410 12845 3476 12849
rect 3407 12793 3417 12845
rect 3469 12793 3479 12845
rect 3534 12844 3580 12882
rect 3534 12810 3540 12844
rect 3574 12810 3580 12844
rect 3410 12789 3476 12793
rect 2282 12703 3364 12737
rect 3534 12627 3580 12810
rect 3803 12737 3837 12886
rect 3981 12946 4027 12981
rect 3981 12912 3987 12946
rect 4021 12912 4027 12946
rect 3981 12877 4027 12912
rect 4077 12946 4123 12981
rect 4077 12912 4083 12946
rect 4117 12912 4123 12946
rect 4077 12877 4123 12912
rect 4173 12946 4219 12981
rect 4173 12912 4179 12946
rect 4213 12912 4219 12946
rect 4173 12877 4219 12912
rect 4269 12946 4315 12981
rect 4269 12912 4275 12946
rect 4309 12912 4315 12946
rect 4269 12877 4315 12912
rect 4365 12946 4411 12981
rect 4365 12912 4371 12946
rect 4405 12912 4411 12946
rect 4365 12877 4411 12912
rect 4461 12946 4507 12981
rect 4461 12912 4467 12946
rect 4501 12912 4507 12946
rect 4461 12877 4507 12912
rect 4557 12946 4603 12981
rect 4557 12912 4563 12946
rect 4597 12912 4603 12946
rect 4557 12877 4603 12912
rect 4653 12946 4699 12981
rect 4653 12912 4659 12946
rect 4693 12912 4699 12946
rect 4653 12877 4699 12912
rect 4749 12946 4795 12981
rect 4749 12912 4755 12946
rect 4789 12912 4795 12946
rect 4749 12877 4795 12912
rect 4845 12946 4891 12981
rect 4845 12912 4851 12946
rect 4885 12912 4891 12946
rect 4845 12877 4891 12912
rect 4941 12946 4987 12981
rect 4941 12912 4947 12946
rect 4981 12912 4987 12946
rect 4941 12877 4987 12912
rect 5055 12954 5061 12988
rect 5095 12954 5101 12988
rect 5055 12916 5101 12954
rect 5055 12882 5061 12916
rect 5095 12899 5101 12916
rect 5095 12882 5550 12899
rect 3971 12846 4037 12849
rect 3968 12794 3978 12846
rect 4030 12794 4040 12846
rect 3971 12789 4037 12794
rect 4083 12737 4117 12877
rect 4163 12846 4229 12849
rect 4159 12794 4169 12846
rect 4221 12794 4231 12846
rect 4163 12789 4229 12794
rect 4275 12737 4309 12877
rect 4355 12846 4421 12849
rect 4351 12794 4361 12846
rect 4413 12794 4423 12846
rect 4355 12789 4421 12794
rect 4467 12737 4501 12877
rect 4547 12846 4613 12849
rect 4543 12794 4553 12846
rect 4605 12794 4615 12846
rect 4547 12789 4613 12794
rect 4659 12737 4693 12877
rect 4739 12845 4805 12849
rect 4736 12793 4746 12845
rect 4798 12793 4808 12845
rect 4739 12789 4805 12793
rect 4851 12737 4885 12877
rect 5055 12868 5550 12882
rect 4931 12845 4997 12849
rect 4928 12793 4938 12845
rect 4990 12793 5000 12845
rect 5055 12844 5303 12868
rect 5055 12810 5061 12844
rect 5095 12834 5303 12844
rect 5337 12834 5395 12868
rect 5429 12834 5487 12868
rect 5521 12834 5550 12868
rect 5095 12810 5550 12834
rect 5055 12803 5550 12810
rect 4931 12789 4997 12793
rect 3803 12703 4885 12737
rect 5055 12628 5101 12803
rect 129 12420 1211 12454
rect 129 11857 163 12420
rect 294 12310 304 12362
rect 356 12310 366 12362
rect 409 12270 443 12420
rect 487 12310 497 12362
rect 549 12310 559 12362
rect 601 12270 635 12420
rect 678 12310 688 12362
rect 740 12310 750 12362
rect 793 12270 827 12420
rect 870 12310 880 12362
rect 932 12310 942 12362
rect 985 12270 1019 12420
rect 1062 12310 1072 12362
rect 1124 12310 1134 12362
rect 1177 12270 1211 12420
rect 1254 12310 1264 12362
rect 1316 12310 1326 12362
rect 1381 12326 1427 12490
rect 2282 12424 3364 12458
rect 1381 12292 1387 12326
rect 1421 12292 1427 12326
rect 1512 12303 1522 12363
rect 1578 12303 1792 12363
rect 1852 12303 1862 12363
rect 307 12223 353 12270
rect 307 12189 313 12223
rect 347 12189 353 12223
rect 307 12151 353 12189
rect 307 12117 313 12151
rect 347 12117 353 12151
rect 307 12079 353 12117
rect 307 12045 313 12079
rect 347 12045 353 12079
rect 307 11998 353 12045
rect 403 12223 449 12270
rect 403 12189 409 12223
rect 443 12189 449 12223
rect 403 12151 449 12189
rect 403 12117 409 12151
rect 443 12117 449 12151
rect 403 12079 449 12117
rect 403 12045 409 12079
rect 443 12045 449 12079
rect 403 11998 449 12045
rect 499 12223 545 12270
rect 499 12189 505 12223
rect 539 12189 545 12223
rect 499 12151 545 12189
rect 499 12117 505 12151
rect 539 12117 545 12151
rect 499 12079 545 12117
rect 499 12045 505 12079
rect 539 12045 545 12079
rect 499 11998 545 12045
rect 595 12223 641 12270
rect 595 12189 601 12223
rect 635 12189 641 12223
rect 595 12151 641 12189
rect 595 12117 601 12151
rect 635 12117 641 12151
rect 595 12079 641 12117
rect 595 12045 601 12079
rect 635 12045 641 12079
rect 595 11998 641 12045
rect 691 12223 737 12270
rect 691 12189 697 12223
rect 731 12189 737 12223
rect 691 12151 737 12189
rect 691 12117 697 12151
rect 731 12117 737 12151
rect 691 12079 737 12117
rect 691 12045 697 12079
rect 731 12045 737 12079
rect 691 11998 737 12045
rect 787 12223 833 12270
rect 787 12189 793 12223
rect 827 12189 833 12223
rect 787 12151 833 12189
rect 787 12117 793 12151
rect 827 12117 833 12151
rect 787 12079 833 12117
rect 787 12045 793 12079
rect 827 12045 833 12079
rect 787 11998 833 12045
rect 883 12223 929 12270
rect 883 12189 889 12223
rect 923 12189 929 12223
rect 883 12151 929 12189
rect 883 12117 889 12151
rect 923 12117 929 12151
rect 883 12079 929 12117
rect 883 12045 889 12079
rect 923 12045 929 12079
rect 883 11998 929 12045
rect 979 12223 1025 12270
rect 979 12189 985 12223
rect 1019 12189 1025 12223
rect 979 12151 1025 12189
rect 979 12117 985 12151
rect 1019 12117 1025 12151
rect 979 12079 1025 12117
rect 979 12045 985 12079
rect 1019 12045 1025 12079
rect 979 11998 1025 12045
rect 1075 12223 1121 12270
rect 1075 12189 1081 12223
rect 1115 12189 1121 12223
rect 1075 12151 1121 12189
rect 1075 12117 1081 12151
rect 1115 12117 1121 12151
rect 1075 12079 1121 12117
rect 1075 12045 1081 12079
rect 1115 12045 1121 12079
rect 1075 11998 1121 12045
rect 1171 12223 1217 12270
rect 1171 12189 1177 12223
rect 1211 12189 1217 12223
rect 1171 12151 1217 12189
rect 1171 12117 1177 12151
rect 1211 12117 1217 12151
rect 1171 12079 1217 12117
rect 1171 12045 1177 12079
rect 1211 12045 1217 12079
rect 1171 11998 1217 12045
rect 1267 12223 1313 12270
rect 1267 12189 1273 12223
rect 1307 12189 1313 12223
rect 1267 12151 1313 12189
rect 1267 12117 1273 12151
rect 1307 12117 1313 12151
rect 1267 12079 1313 12117
rect 1267 12045 1273 12079
rect 1307 12045 1313 12079
rect 1267 11998 1313 12045
rect 1381 12254 1427 12292
rect 1381 12220 1387 12254
rect 1421 12220 1427 12254
rect 1381 12182 1427 12220
rect 1381 12148 1387 12182
rect 1421 12148 1427 12182
rect 1381 12110 1427 12148
rect 1381 12076 1387 12110
rect 1421 12076 1427 12110
rect 1381 12066 1427 12076
rect 1381 12064 2160 12066
rect 1381 12038 2056 12064
rect 1381 12013 1387 12038
rect 1380 12004 1387 12013
rect 1421 12004 2056 12038
rect 0 11823 163 11857
rect 129 11446 163 11823
rect 313 11857 347 11998
rect 505 11857 539 11998
rect 697 11857 731 11998
rect 889 11857 923 11998
rect 1081 11857 1115 11998
rect 1273 11857 1307 11998
rect 1380 11956 2056 12004
rect 2190 11956 2200 12064
rect 1380 11954 2160 11956
rect 2282 11861 2316 12424
rect 2447 12314 2457 12366
rect 2509 12314 2519 12366
rect 2562 12274 2596 12424
rect 2640 12314 2650 12366
rect 2702 12314 2712 12366
rect 2754 12274 2788 12424
rect 2831 12314 2841 12366
rect 2893 12314 2903 12366
rect 2946 12274 2980 12424
rect 3023 12314 3033 12366
rect 3085 12314 3095 12366
rect 3138 12274 3172 12424
rect 3215 12314 3225 12366
rect 3277 12314 3287 12366
rect 3330 12274 3364 12424
rect 3407 12314 3417 12366
rect 3469 12314 3479 12366
rect 3534 12330 3580 12538
rect 3534 12296 3540 12330
rect 3574 12296 3580 12330
rect 2460 12227 2506 12274
rect 2460 12193 2466 12227
rect 2500 12193 2506 12227
rect 2460 12155 2506 12193
rect 2460 12121 2466 12155
rect 2500 12121 2506 12155
rect 2460 12083 2506 12121
rect 2460 12049 2466 12083
rect 2500 12049 2506 12083
rect 2460 12002 2506 12049
rect 2556 12227 2602 12274
rect 2556 12193 2562 12227
rect 2596 12193 2602 12227
rect 2556 12155 2602 12193
rect 2556 12121 2562 12155
rect 2596 12121 2602 12155
rect 2556 12083 2602 12121
rect 2556 12049 2562 12083
rect 2596 12049 2602 12083
rect 2556 12002 2602 12049
rect 2652 12227 2698 12274
rect 2652 12193 2658 12227
rect 2692 12193 2698 12227
rect 2652 12155 2698 12193
rect 2652 12121 2658 12155
rect 2692 12121 2698 12155
rect 2652 12083 2698 12121
rect 2652 12049 2658 12083
rect 2692 12049 2698 12083
rect 2652 12002 2698 12049
rect 2748 12227 2794 12274
rect 2748 12193 2754 12227
rect 2788 12193 2794 12227
rect 2748 12155 2794 12193
rect 2748 12121 2754 12155
rect 2788 12121 2794 12155
rect 2748 12083 2794 12121
rect 2748 12049 2754 12083
rect 2788 12049 2794 12083
rect 2748 12002 2794 12049
rect 2844 12227 2890 12274
rect 2844 12193 2850 12227
rect 2884 12193 2890 12227
rect 2844 12155 2890 12193
rect 2844 12121 2850 12155
rect 2884 12121 2890 12155
rect 2844 12083 2890 12121
rect 2844 12049 2850 12083
rect 2884 12049 2890 12083
rect 2844 12002 2890 12049
rect 2940 12227 2986 12274
rect 2940 12193 2946 12227
rect 2980 12193 2986 12227
rect 2940 12155 2986 12193
rect 2940 12121 2946 12155
rect 2980 12121 2986 12155
rect 2940 12083 2986 12121
rect 2940 12049 2946 12083
rect 2980 12049 2986 12083
rect 2940 12002 2986 12049
rect 3036 12227 3082 12274
rect 3036 12193 3042 12227
rect 3076 12193 3082 12227
rect 3036 12155 3082 12193
rect 3036 12121 3042 12155
rect 3076 12121 3082 12155
rect 3036 12083 3082 12121
rect 3036 12049 3042 12083
rect 3076 12049 3082 12083
rect 3036 12002 3082 12049
rect 3132 12227 3178 12274
rect 3132 12193 3138 12227
rect 3172 12193 3178 12227
rect 3132 12155 3178 12193
rect 3132 12121 3138 12155
rect 3172 12121 3178 12155
rect 3132 12083 3178 12121
rect 3132 12049 3138 12083
rect 3172 12049 3178 12083
rect 3132 12002 3178 12049
rect 3228 12227 3274 12274
rect 3228 12193 3234 12227
rect 3268 12193 3274 12227
rect 3228 12155 3274 12193
rect 3228 12121 3234 12155
rect 3268 12121 3274 12155
rect 3228 12083 3274 12121
rect 3228 12049 3234 12083
rect 3268 12049 3274 12083
rect 3228 12002 3274 12049
rect 3324 12227 3370 12274
rect 3324 12193 3330 12227
rect 3364 12193 3370 12227
rect 3324 12155 3370 12193
rect 3324 12121 3330 12155
rect 3364 12121 3370 12155
rect 3324 12083 3370 12121
rect 3324 12049 3330 12083
rect 3364 12049 3370 12083
rect 3324 12002 3370 12049
rect 3420 12227 3466 12274
rect 3420 12193 3426 12227
rect 3460 12193 3466 12227
rect 3420 12155 3466 12193
rect 3420 12121 3426 12155
rect 3460 12121 3466 12155
rect 3420 12083 3466 12121
rect 3420 12049 3426 12083
rect 3460 12049 3466 12083
rect 3420 12002 3466 12049
rect 3534 12258 3580 12296
rect 3534 12224 3540 12258
rect 3574 12224 3580 12258
rect 3534 12186 3580 12224
rect 3534 12152 3540 12186
rect 3574 12152 3580 12186
rect 3534 12114 3580 12152
rect 3534 12080 3540 12114
rect 3574 12080 3580 12114
rect 3534 12042 3580 12080
rect 3534 12008 3540 12042
rect 3574 12008 3580 12042
rect 2101 11857 2316 11861
rect 313 11827 2316 11857
rect 313 11823 2141 11827
rect 313 11690 347 11823
rect 505 11690 539 11823
rect 697 11690 731 11823
rect 889 11690 923 11823
rect 1081 11690 1115 11823
rect 1273 11690 1307 11823
rect 1381 11697 1608 11720
rect 307 11655 353 11690
rect 307 11621 313 11655
rect 347 11621 353 11655
rect 307 11586 353 11621
rect 403 11655 449 11690
rect 403 11621 409 11655
rect 443 11621 449 11655
rect 403 11586 449 11621
rect 499 11655 545 11690
rect 499 11621 505 11655
rect 539 11621 545 11655
rect 499 11586 545 11621
rect 595 11655 641 11690
rect 595 11621 601 11655
rect 635 11621 641 11655
rect 595 11586 641 11621
rect 691 11655 737 11690
rect 691 11621 697 11655
rect 731 11621 737 11655
rect 691 11586 737 11621
rect 787 11655 833 11690
rect 787 11621 793 11655
rect 827 11621 833 11655
rect 787 11586 833 11621
rect 883 11655 929 11690
rect 883 11621 889 11655
rect 923 11621 929 11655
rect 883 11586 929 11621
rect 979 11655 1025 11690
rect 979 11621 985 11655
rect 1019 11621 1025 11655
rect 979 11586 1025 11621
rect 1075 11655 1121 11690
rect 1075 11621 1081 11655
rect 1115 11621 1121 11655
rect 1075 11586 1121 11621
rect 1171 11655 1217 11690
rect 1171 11621 1177 11655
rect 1211 11621 1217 11655
rect 1171 11586 1217 11621
rect 1267 11655 1313 11690
rect 1267 11621 1273 11655
rect 1307 11621 1313 11655
rect 1267 11586 1313 11621
rect 1381 11663 1387 11697
rect 1421 11663 1608 11697
rect 1381 11625 1608 11663
rect 1381 11591 1387 11625
rect 1421 11600 1608 11625
rect 1421 11591 1427 11600
rect 1560 11598 1608 11600
rect 1598 11596 1608 11598
rect 1720 11596 1730 11720
rect 297 11555 363 11558
rect 294 11503 304 11555
rect 356 11503 366 11555
rect 297 11498 363 11503
rect 409 11446 443 11586
rect 489 11555 555 11558
rect 485 11503 495 11555
rect 547 11503 557 11555
rect 489 11498 555 11503
rect 601 11446 635 11586
rect 681 11555 747 11558
rect 677 11503 687 11555
rect 739 11503 749 11555
rect 681 11498 747 11503
rect 793 11446 827 11586
rect 873 11555 939 11558
rect 869 11503 879 11555
rect 931 11503 941 11555
rect 873 11498 939 11503
rect 985 11446 1019 11586
rect 1065 11554 1131 11558
rect 1062 11502 1072 11554
rect 1124 11502 1134 11554
rect 1065 11498 1131 11502
rect 1177 11446 1211 11586
rect 1257 11554 1323 11558
rect 1254 11502 1264 11554
rect 1316 11502 1326 11554
rect 1381 11553 1427 11591
rect 1920 11558 1930 11560
rect 1381 11519 1387 11553
rect 1421 11519 1427 11553
rect 1257 11498 1323 11502
rect 129 11412 1211 11446
rect 1381 11376 1427 11519
rect 1458 11502 1468 11558
rect 1524 11504 1930 11558
rect 1986 11504 1996 11560
rect 1524 11502 1986 11504
rect 2282 11450 2316 11827
rect 2466 11861 2500 12002
rect 2658 11861 2692 12002
rect 2850 11861 2884 12002
rect 3042 11861 3076 12002
rect 3234 11861 3268 12002
rect 3426 11861 3460 12002
rect 3534 11964 3580 12008
rect 3803 12424 4885 12458
rect 3803 11861 3837 12424
rect 3968 12314 3978 12366
rect 4030 12314 4040 12366
rect 4083 12274 4117 12424
rect 4161 12314 4171 12366
rect 4223 12314 4233 12366
rect 4275 12274 4309 12424
rect 4352 12314 4362 12366
rect 4414 12314 4424 12366
rect 4467 12274 4501 12424
rect 4544 12314 4554 12366
rect 4606 12314 4616 12366
rect 4659 12274 4693 12424
rect 4736 12314 4746 12366
rect 4798 12314 4808 12366
rect 4851 12274 4885 12424
rect 4928 12314 4938 12366
rect 4990 12314 5000 12366
rect 5055 12330 5101 12535
rect 5055 12296 5061 12330
rect 5095 12296 5101 12330
rect 3981 12227 4027 12274
rect 3981 12193 3987 12227
rect 4021 12193 4027 12227
rect 3981 12155 4027 12193
rect 3981 12121 3987 12155
rect 4021 12121 4027 12155
rect 3981 12083 4027 12121
rect 3981 12049 3987 12083
rect 4021 12049 4027 12083
rect 3981 12002 4027 12049
rect 4077 12227 4123 12274
rect 4077 12193 4083 12227
rect 4117 12193 4123 12227
rect 4077 12155 4123 12193
rect 4077 12121 4083 12155
rect 4117 12121 4123 12155
rect 4077 12083 4123 12121
rect 4077 12049 4083 12083
rect 4117 12049 4123 12083
rect 4077 12002 4123 12049
rect 4173 12227 4219 12274
rect 4173 12193 4179 12227
rect 4213 12193 4219 12227
rect 4173 12155 4219 12193
rect 4173 12121 4179 12155
rect 4213 12121 4219 12155
rect 4173 12083 4219 12121
rect 4173 12049 4179 12083
rect 4213 12049 4219 12083
rect 4173 12002 4219 12049
rect 4269 12227 4315 12274
rect 4269 12193 4275 12227
rect 4309 12193 4315 12227
rect 4269 12155 4315 12193
rect 4269 12121 4275 12155
rect 4309 12121 4315 12155
rect 4269 12083 4315 12121
rect 4269 12049 4275 12083
rect 4309 12049 4315 12083
rect 4269 12002 4315 12049
rect 4365 12227 4411 12274
rect 4365 12193 4371 12227
rect 4405 12193 4411 12227
rect 4365 12155 4411 12193
rect 4365 12121 4371 12155
rect 4405 12121 4411 12155
rect 4365 12083 4411 12121
rect 4365 12049 4371 12083
rect 4405 12049 4411 12083
rect 4365 12002 4411 12049
rect 4461 12227 4507 12274
rect 4461 12193 4467 12227
rect 4501 12193 4507 12227
rect 4461 12155 4507 12193
rect 4461 12121 4467 12155
rect 4501 12121 4507 12155
rect 4461 12083 4507 12121
rect 4461 12049 4467 12083
rect 4501 12049 4507 12083
rect 4461 12002 4507 12049
rect 4557 12227 4603 12274
rect 4557 12193 4563 12227
rect 4597 12193 4603 12227
rect 4557 12155 4603 12193
rect 4557 12121 4563 12155
rect 4597 12121 4603 12155
rect 4557 12083 4603 12121
rect 4557 12049 4563 12083
rect 4597 12049 4603 12083
rect 4557 12002 4603 12049
rect 4653 12227 4699 12274
rect 4653 12193 4659 12227
rect 4693 12193 4699 12227
rect 4653 12155 4699 12193
rect 4653 12121 4659 12155
rect 4693 12121 4699 12155
rect 4653 12083 4699 12121
rect 4653 12049 4659 12083
rect 4693 12049 4699 12083
rect 4653 12002 4699 12049
rect 4749 12227 4795 12274
rect 4749 12193 4755 12227
rect 4789 12193 4795 12227
rect 4749 12155 4795 12193
rect 4749 12121 4755 12155
rect 4789 12121 4795 12155
rect 4749 12083 4795 12121
rect 4749 12049 4755 12083
rect 4789 12049 4795 12083
rect 4749 12002 4795 12049
rect 4845 12227 4891 12274
rect 4845 12193 4851 12227
rect 4885 12193 4891 12227
rect 4845 12155 4891 12193
rect 4845 12121 4851 12155
rect 4885 12121 4891 12155
rect 4845 12083 4891 12121
rect 4845 12049 4851 12083
rect 4885 12049 4891 12083
rect 4845 12002 4891 12049
rect 4941 12227 4987 12274
rect 4941 12193 4947 12227
rect 4981 12193 4987 12227
rect 4941 12155 4987 12193
rect 4941 12121 4947 12155
rect 4981 12121 4987 12155
rect 4941 12083 4987 12121
rect 4941 12049 4947 12083
rect 4981 12049 4987 12083
rect 4941 12002 4987 12049
rect 5055 12258 5101 12296
rect 5055 12224 5061 12258
rect 5095 12224 5101 12258
rect 5055 12186 5101 12224
rect 5055 12152 5061 12186
rect 5095 12155 5101 12186
rect 5274 12155 5550 12156
rect 5095 12152 5550 12155
rect 5055 12125 5550 12152
rect 5055 12114 5303 12125
rect 5055 12080 5061 12114
rect 5095 12091 5303 12114
rect 5337 12091 5395 12125
rect 5429 12091 5487 12125
rect 5521 12091 5550 12125
rect 5095 12080 5550 12091
rect 5055 12060 5550 12080
rect 5055 12042 5101 12060
rect 5055 12008 5061 12042
rect 5095 12008 5101 12042
rect 2466 11827 3837 11861
rect 2466 11694 2500 11827
rect 2658 11694 2692 11827
rect 2850 11694 2884 11827
rect 3042 11694 3076 11827
rect 3234 11694 3268 11827
rect 3426 11694 3460 11827
rect 3671 11737 3681 11789
rect 3733 11737 3743 11789
rect 3679 11736 3691 11737
rect 3725 11736 3737 11737
rect 3679 11730 3737 11736
rect 3534 11701 3580 11724
rect 2460 11659 2506 11694
rect 2460 11625 2466 11659
rect 2500 11625 2506 11659
rect 2460 11590 2506 11625
rect 2556 11659 2602 11694
rect 2556 11625 2562 11659
rect 2596 11625 2602 11659
rect 2556 11590 2602 11625
rect 2652 11659 2698 11694
rect 2652 11625 2658 11659
rect 2692 11625 2698 11659
rect 2652 11590 2698 11625
rect 2748 11659 2794 11694
rect 2748 11625 2754 11659
rect 2788 11625 2794 11659
rect 2748 11590 2794 11625
rect 2844 11659 2890 11694
rect 2844 11625 2850 11659
rect 2884 11625 2890 11659
rect 2844 11590 2890 11625
rect 2940 11659 2986 11694
rect 2940 11625 2946 11659
rect 2980 11625 2986 11659
rect 2940 11590 2986 11625
rect 3036 11659 3082 11694
rect 3036 11625 3042 11659
rect 3076 11625 3082 11659
rect 3036 11590 3082 11625
rect 3132 11659 3178 11694
rect 3132 11625 3138 11659
rect 3172 11625 3178 11659
rect 3132 11590 3178 11625
rect 3228 11659 3274 11694
rect 3228 11625 3234 11659
rect 3268 11625 3274 11659
rect 3228 11590 3274 11625
rect 3324 11659 3370 11694
rect 3324 11625 3330 11659
rect 3364 11625 3370 11659
rect 3324 11590 3370 11625
rect 3420 11659 3466 11694
rect 3420 11625 3426 11659
rect 3460 11625 3466 11659
rect 3420 11590 3466 11625
rect 3534 11667 3540 11701
rect 3574 11699 3580 11701
rect 3803 11699 3837 11827
rect 3574 11698 3680 11699
rect 3734 11698 3837 11699
rect 3574 11686 3687 11698
rect 3574 11667 3647 11686
rect 3534 11629 3647 11667
rect 3534 11595 3540 11629
rect 3574 11610 3647 11629
rect 3681 11610 3687 11686
rect 3574 11599 3687 11610
rect 3574 11595 3580 11599
rect 3641 11598 3687 11599
rect 3729 11686 3837 11698
rect 3987 11861 4021 12002
rect 4179 11861 4213 12002
rect 4371 11861 4405 12002
rect 4563 11861 4597 12002
rect 4755 11861 4789 12002
rect 4947 11861 4981 12002
rect 5055 11964 5101 12008
rect 5683 11915 5743 13168
rect 5177 11881 5743 11915
rect 5177 11861 5211 11881
rect 3987 11827 5211 11861
rect 3987 11694 4021 11827
rect 4179 11694 4213 11827
rect 4371 11694 4405 11827
rect 4563 11694 4597 11827
rect 4755 11694 4789 11827
rect 4947 11694 4981 11827
rect 5438 11823 5512 11824
rect 5326 11821 5400 11822
rect 5326 11769 5337 11821
rect 5389 11769 5400 11821
rect 5438 11771 5449 11823
rect 5501 11771 5512 11823
rect 5438 11770 5512 11771
rect 5326 11768 5400 11769
rect 5055 11701 5101 11724
rect 3729 11610 3735 11686
rect 3769 11610 3837 11686
rect 3729 11599 3837 11610
rect 3729 11598 3775 11599
rect 2450 11559 2516 11562
rect 2447 11507 2457 11559
rect 2509 11507 2519 11559
rect 2450 11502 2516 11507
rect 2562 11450 2596 11590
rect 2642 11559 2708 11562
rect 2638 11507 2648 11559
rect 2700 11507 2710 11559
rect 2642 11502 2708 11507
rect 2754 11450 2788 11590
rect 2834 11559 2900 11562
rect 2830 11507 2840 11559
rect 2892 11507 2902 11559
rect 2834 11502 2900 11507
rect 2946 11450 2980 11590
rect 3026 11559 3092 11562
rect 3022 11507 3032 11559
rect 3084 11507 3094 11559
rect 3026 11502 3092 11507
rect 3138 11450 3172 11590
rect 3218 11558 3284 11562
rect 3215 11506 3225 11558
rect 3277 11506 3287 11558
rect 3218 11502 3284 11506
rect 3330 11450 3364 11590
rect 3410 11558 3476 11562
rect 3407 11506 3417 11558
rect 3469 11506 3479 11558
rect 3534 11557 3580 11595
rect 3534 11523 3540 11557
rect 3574 11523 3580 11557
rect 3410 11502 3476 11506
rect 2282 11416 3364 11450
rect 3534 11340 3580 11523
rect 3803 11450 3837 11599
rect 3981 11659 4027 11694
rect 3981 11625 3987 11659
rect 4021 11625 4027 11659
rect 3981 11590 4027 11625
rect 4077 11659 4123 11694
rect 4077 11625 4083 11659
rect 4117 11625 4123 11659
rect 4077 11590 4123 11625
rect 4173 11659 4219 11694
rect 4173 11625 4179 11659
rect 4213 11625 4219 11659
rect 4173 11590 4219 11625
rect 4269 11659 4315 11694
rect 4269 11625 4275 11659
rect 4309 11625 4315 11659
rect 4269 11590 4315 11625
rect 4365 11659 4411 11694
rect 4365 11625 4371 11659
rect 4405 11625 4411 11659
rect 4365 11590 4411 11625
rect 4461 11659 4507 11694
rect 4461 11625 4467 11659
rect 4501 11625 4507 11659
rect 4461 11590 4507 11625
rect 4557 11659 4603 11694
rect 4557 11625 4563 11659
rect 4597 11625 4603 11659
rect 4557 11590 4603 11625
rect 4653 11659 4699 11694
rect 4653 11625 4659 11659
rect 4693 11625 4699 11659
rect 4653 11590 4699 11625
rect 4749 11659 4795 11694
rect 4749 11625 4755 11659
rect 4789 11625 4795 11659
rect 4749 11590 4795 11625
rect 4845 11659 4891 11694
rect 4845 11625 4851 11659
rect 4885 11625 4891 11659
rect 4845 11590 4891 11625
rect 4941 11659 4987 11694
rect 4941 11625 4947 11659
rect 4981 11625 4987 11659
rect 4941 11590 4987 11625
rect 5055 11667 5061 11701
rect 5095 11667 5101 11701
rect 5055 11629 5101 11667
rect 5055 11595 5061 11629
rect 5095 11612 5101 11629
rect 5095 11595 5550 11612
rect 3971 11559 4037 11562
rect 3968 11507 3978 11559
rect 4030 11507 4040 11559
rect 3971 11502 4037 11507
rect 4083 11450 4117 11590
rect 4163 11559 4229 11562
rect 4159 11507 4169 11559
rect 4221 11507 4231 11559
rect 4163 11502 4229 11507
rect 4275 11450 4309 11590
rect 4355 11559 4421 11562
rect 4351 11507 4361 11559
rect 4413 11507 4423 11559
rect 4355 11502 4421 11507
rect 4467 11450 4501 11590
rect 4547 11559 4613 11562
rect 4543 11507 4553 11559
rect 4605 11507 4615 11559
rect 4547 11502 4613 11507
rect 4659 11450 4693 11590
rect 4739 11558 4805 11562
rect 4736 11506 4746 11558
rect 4798 11506 4808 11558
rect 4739 11502 4805 11506
rect 4851 11450 4885 11590
rect 5055 11581 5550 11595
rect 4931 11558 4997 11562
rect 4928 11506 4938 11558
rect 4990 11506 5000 11558
rect 5055 11557 5303 11581
rect 5055 11523 5061 11557
rect 5095 11547 5303 11557
rect 5337 11547 5395 11581
rect 5429 11547 5487 11581
rect 5521 11547 5550 11581
rect 5095 11523 5550 11547
rect 5055 11516 5550 11523
rect 4931 11502 4997 11506
rect 3803 11416 4885 11450
rect 5055 11341 5101 11516
rect 129 11133 1211 11167
rect 129 10570 163 11133
rect 294 11023 304 11075
rect 356 11023 366 11075
rect 409 10983 443 11133
rect 487 11023 497 11075
rect 549 11023 559 11075
rect 601 10983 635 11133
rect 678 11023 688 11075
rect 740 11023 750 11075
rect 793 10983 827 11133
rect 870 11023 880 11075
rect 932 11023 942 11075
rect 985 10983 1019 11133
rect 1062 11023 1072 11075
rect 1124 11023 1134 11075
rect 1177 10983 1211 11133
rect 1254 11023 1264 11075
rect 1316 11023 1326 11075
rect 1381 11039 1427 11203
rect 2282 11137 3364 11171
rect 1381 11005 1387 11039
rect 1421 11005 1427 11039
rect 1512 11016 1522 11076
rect 1578 11016 1792 11076
rect 1852 11016 1862 11076
rect 307 10936 353 10983
rect 307 10902 313 10936
rect 347 10902 353 10936
rect 307 10864 353 10902
rect 307 10830 313 10864
rect 347 10830 353 10864
rect 307 10792 353 10830
rect 307 10758 313 10792
rect 347 10758 353 10792
rect 307 10711 353 10758
rect 403 10936 449 10983
rect 403 10902 409 10936
rect 443 10902 449 10936
rect 403 10864 449 10902
rect 403 10830 409 10864
rect 443 10830 449 10864
rect 403 10792 449 10830
rect 403 10758 409 10792
rect 443 10758 449 10792
rect 403 10711 449 10758
rect 499 10936 545 10983
rect 499 10902 505 10936
rect 539 10902 545 10936
rect 499 10864 545 10902
rect 499 10830 505 10864
rect 539 10830 545 10864
rect 499 10792 545 10830
rect 499 10758 505 10792
rect 539 10758 545 10792
rect 499 10711 545 10758
rect 595 10936 641 10983
rect 595 10902 601 10936
rect 635 10902 641 10936
rect 595 10864 641 10902
rect 595 10830 601 10864
rect 635 10830 641 10864
rect 595 10792 641 10830
rect 595 10758 601 10792
rect 635 10758 641 10792
rect 595 10711 641 10758
rect 691 10936 737 10983
rect 691 10902 697 10936
rect 731 10902 737 10936
rect 691 10864 737 10902
rect 691 10830 697 10864
rect 731 10830 737 10864
rect 691 10792 737 10830
rect 691 10758 697 10792
rect 731 10758 737 10792
rect 691 10711 737 10758
rect 787 10936 833 10983
rect 787 10902 793 10936
rect 827 10902 833 10936
rect 787 10864 833 10902
rect 787 10830 793 10864
rect 827 10830 833 10864
rect 787 10792 833 10830
rect 787 10758 793 10792
rect 827 10758 833 10792
rect 787 10711 833 10758
rect 883 10936 929 10983
rect 883 10902 889 10936
rect 923 10902 929 10936
rect 883 10864 929 10902
rect 883 10830 889 10864
rect 923 10830 929 10864
rect 883 10792 929 10830
rect 883 10758 889 10792
rect 923 10758 929 10792
rect 883 10711 929 10758
rect 979 10936 1025 10983
rect 979 10902 985 10936
rect 1019 10902 1025 10936
rect 979 10864 1025 10902
rect 979 10830 985 10864
rect 1019 10830 1025 10864
rect 979 10792 1025 10830
rect 979 10758 985 10792
rect 1019 10758 1025 10792
rect 979 10711 1025 10758
rect 1075 10936 1121 10983
rect 1075 10902 1081 10936
rect 1115 10902 1121 10936
rect 1075 10864 1121 10902
rect 1075 10830 1081 10864
rect 1115 10830 1121 10864
rect 1075 10792 1121 10830
rect 1075 10758 1081 10792
rect 1115 10758 1121 10792
rect 1075 10711 1121 10758
rect 1171 10936 1217 10983
rect 1171 10902 1177 10936
rect 1211 10902 1217 10936
rect 1171 10864 1217 10902
rect 1171 10830 1177 10864
rect 1211 10830 1217 10864
rect 1171 10792 1217 10830
rect 1171 10758 1177 10792
rect 1211 10758 1217 10792
rect 1171 10711 1217 10758
rect 1267 10936 1313 10983
rect 1267 10902 1273 10936
rect 1307 10902 1313 10936
rect 1267 10864 1313 10902
rect 1267 10830 1273 10864
rect 1307 10830 1313 10864
rect 1267 10792 1313 10830
rect 1267 10758 1273 10792
rect 1307 10758 1313 10792
rect 1267 10711 1313 10758
rect 1381 10967 1427 11005
rect 1381 10933 1387 10967
rect 1421 10933 1427 10967
rect 1381 10895 1427 10933
rect 1381 10861 1387 10895
rect 1421 10861 1427 10895
rect 1381 10823 1427 10861
rect 1381 10789 1387 10823
rect 1421 10789 1427 10823
rect 1381 10779 1427 10789
rect 1381 10777 2160 10779
rect 1381 10751 2056 10777
rect 1381 10726 1387 10751
rect 1380 10717 1387 10726
rect 1421 10717 2056 10751
rect 0 10536 163 10570
rect 129 10159 163 10536
rect 313 10570 347 10711
rect 505 10570 539 10711
rect 697 10570 731 10711
rect 889 10570 923 10711
rect 1081 10570 1115 10711
rect 1273 10570 1307 10711
rect 1380 10669 2056 10717
rect 2190 10669 2200 10777
rect 1380 10667 2160 10669
rect 2282 10574 2316 11137
rect 2447 11027 2457 11079
rect 2509 11027 2519 11079
rect 2562 10987 2596 11137
rect 2640 11027 2650 11079
rect 2702 11027 2712 11079
rect 2754 10987 2788 11137
rect 2831 11027 2841 11079
rect 2893 11027 2903 11079
rect 2946 10987 2980 11137
rect 3023 11027 3033 11079
rect 3085 11027 3095 11079
rect 3138 10987 3172 11137
rect 3215 11027 3225 11079
rect 3277 11027 3287 11079
rect 3330 10987 3364 11137
rect 3407 11027 3417 11079
rect 3469 11027 3479 11079
rect 3534 11043 3580 11251
rect 3534 11009 3540 11043
rect 3574 11009 3580 11043
rect 2460 10940 2506 10987
rect 2460 10906 2466 10940
rect 2500 10906 2506 10940
rect 2460 10868 2506 10906
rect 2460 10834 2466 10868
rect 2500 10834 2506 10868
rect 2460 10796 2506 10834
rect 2460 10762 2466 10796
rect 2500 10762 2506 10796
rect 2460 10715 2506 10762
rect 2556 10940 2602 10987
rect 2556 10906 2562 10940
rect 2596 10906 2602 10940
rect 2556 10868 2602 10906
rect 2556 10834 2562 10868
rect 2596 10834 2602 10868
rect 2556 10796 2602 10834
rect 2556 10762 2562 10796
rect 2596 10762 2602 10796
rect 2556 10715 2602 10762
rect 2652 10940 2698 10987
rect 2652 10906 2658 10940
rect 2692 10906 2698 10940
rect 2652 10868 2698 10906
rect 2652 10834 2658 10868
rect 2692 10834 2698 10868
rect 2652 10796 2698 10834
rect 2652 10762 2658 10796
rect 2692 10762 2698 10796
rect 2652 10715 2698 10762
rect 2748 10940 2794 10987
rect 2748 10906 2754 10940
rect 2788 10906 2794 10940
rect 2748 10868 2794 10906
rect 2748 10834 2754 10868
rect 2788 10834 2794 10868
rect 2748 10796 2794 10834
rect 2748 10762 2754 10796
rect 2788 10762 2794 10796
rect 2748 10715 2794 10762
rect 2844 10940 2890 10987
rect 2844 10906 2850 10940
rect 2884 10906 2890 10940
rect 2844 10868 2890 10906
rect 2844 10834 2850 10868
rect 2884 10834 2890 10868
rect 2844 10796 2890 10834
rect 2844 10762 2850 10796
rect 2884 10762 2890 10796
rect 2844 10715 2890 10762
rect 2940 10940 2986 10987
rect 2940 10906 2946 10940
rect 2980 10906 2986 10940
rect 2940 10868 2986 10906
rect 2940 10834 2946 10868
rect 2980 10834 2986 10868
rect 2940 10796 2986 10834
rect 2940 10762 2946 10796
rect 2980 10762 2986 10796
rect 2940 10715 2986 10762
rect 3036 10940 3082 10987
rect 3036 10906 3042 10940
rect 3076 10906 3082 10940
rect 3036 10868 3082 10906
rect 3036 10834 3042 10868
rect 3076 10834 3082 10868
rect 3036 10796 3082 10834
rect 3036 10762 3042 10796
rect 3076 10762 3082 10796
rect 3036 10715 3082 10762
rect 3132 10940 3178 10987
rect 3132 10906 3138 10940
rect 3172 10906 3178 10940
rect 3132 10868 3178 10906
rect 3132 10834 3138 10868
rect 3172 10834 3178 10868
rect 3132 10796 3178 10834
rect 3132 10762 3138 10796
rect 3172 10762 3178 10796
rect 3132 10715 3178 10762
rect 3228 10940 3274 10987
rect 3228 10906 3234 10940
rect 3268 10906 3274 10940
rect 3228 10868 3274 10906
rect 3228 10834 3234 10868
rect 3268 10834 3274 10868
rect 3228 10796 3274 10834
rect 3228 10762 3234 10796
rect 3268 10762 3274 10796
rect 3228 10715 3274 10762
rect 3324 10940 3370 10987
rect 3324 10906 3330 10940
rect 3364 10906 3370 10940
rect 3324 10868 3370 10906
rect 3324 10834 3330 10868
rect 3364 10834 3370 10868
rect 3324 10796 3370 10834
rect 3324 10762 3330 10796
rect 3364 10762 3370 10796
rect 3324 10715 3370 10762
rect 3420 10940 3466 10987
rect 3420 10906 3426 10940
rect 3460 10906 3466 10940
rect 3420 10868 3466 10906
rect 3420 10834 3426 10868
rect 3460 10834 3466 10868
rect 3420 10796 3466 10834
rect 3420 10762 3426 10796
rect 3460 10762 3466 10796
rect 3420 10715 3466 10762
rect 3534 10971 3580 11009
rect 3534 10937 3540 10971
rect 3574 10937 3580 10971
rect 3534 10899 3580 10937
rect 3534 10865 3540 10899
rect 3574 10865 3580 10899
rect 3534 10827 3580 10865
rect 3534 10793 3540 10827
rect 3574 10793 3580 10827
rect 3534 10755 3580 10793
rect 3534 10721 3540 10755
rect 3574 10721 3580 10755
rect 2101 10570 2316 10574
rect 313 10540 2316 10570
rect 313 10536 2141 10540
rect 313 10403 347 10536
rect 505 10403 539 10536
rect 697 10403 731 10536
rect 889 10403 923 10536
rect 1081 10403 1115 10536
rect 1273 10403 1307 10536
rect 1381 10410 1608 10433
rect 307 10368 353 10403
rect 307 10334 313 10368
rect 347 10334 353 10368
rect 307 10299 353 10334
rect 403 10368 449 10403
rect 403 10334 409 10368
rect 443 10334 449 10368
rect 403 10299 449 10334
rect 499 10368 545 10403
rect 499 10334 505 10368
rect 539 10334 545 10368
rect 499 10299 545 10334
rect 595 10368 641 10403
rect 595 10334 601 10368
rect 635 10334 641 10368
rect 595 10299 641 10334
rect 691 10368 737 10403
rect 691 10334 697 10368
rect 731 10334 737 10368
rect 691 10299 737 10334
rect 787 10368 833 10403
rect 787 10334 793 10368
rect 827 10334 833 10368
rect 787 10299 833 10334
rect 883 10368 929 10403
rect 883 10334 889 10368
rect 923 10334 929 10368
rect 883 10299 929 10334
rect 979 10368 1025 10403
rect 979 10334 985 10368
rect 1019 10334 1025 10368
rect 979 10299 1025 10334
rect 1075 10368 1121 10403
rect 1075 10334 1081 10368
rect 1115 10334 1121 10368
rect 1075 10299 1121 10334
rect 1171 10368 1217 10403
rect 1171 10334 1177 10368
rect 1211 10334 1217 10368
rect 1171 10299 1217 10334
rect 1267 10368 1313 10403
rect 1267 10334 1273 10368
rect 1307 10334 1313 10368
rect 1267 10299 1313 10334
rect 1381 10376 1387 10410
rect 1421 10376 1608 10410
rect 1381 10338 1608 10376
rect 1381 10304 1387 10338
rect 1421 10313 1608 10338
rect 1421 10304 1427 10313
rect 1560 10311 1608 10313
rect 1598 10309 1608 10311
rect 1720 10309 1730 10433
rect 297 10268 363 10271
rect 294 10216 304 10268
rect 356 10216 366 10268
rect 297 10211 363 10216
rect 409 10159 443 10299
rect 489 10268 555 10271
rect 485 10216 495 10268
rect 547 10216 557 10268
rect 489 10211 555 10216
rect 601 10159 635 10299
rect 681 10268 747 10271
rect 677 10216 687 10268
rect 739 10216 749 10268
rect 681 10211 747 10216
rect 793 10159 827 10299
rect 873 10268 939 10271
rect 869 10216 879 10268
rect 931 10216 941 10268
rect 873 10211 939 10216
rect 985 10159 1019 10299
rect 1065 10267 1131 10271
rect 1062 10215 1072 10267
rect 1124 10215 1134 10267
rect 1065 10211 1131 10215
rect 1177 10159 1211 10299
rect 1257 10267 1323 10271
rect 1254 10215 1264 10267
rect 1316 10215 1326 10267
rect 1381 10266 1427 10304
rect 1920 10271 1930 10273
rect 1381 10232 1387 10266
rect 1421 10232 1427 10266
rect 1257 10211 1323 10215
rect 129 10125 1211 10159
rect 1381 10089 1427 10232
rect 1458 10215 1468 10271
rect 1524 10217 1930 10271
rect 1986 10217 1996 10273
rect 1524 10215 1986 10217
rect 2282 10163 2316 10540
rect 2466 10574 2500 10715
rect 2658 10574 2692 10715
rect 2850 10574 2884 10715
rect 3042 10574 3076 10715
rect 3234 10574 3268 10715
rect 3426 10574 3460 10715
rect 3534 10677 3580 10721
rect 3803 11137 4885 11171
rect 3803 10574 3837 11137
rect 3968 11027 3978 11079
rect 4030 11027 4040 11079
rect 4083 10987 4117 11137
rect 4161 11027 4171 11079
rect 4223 11027 4233 11079
rect 4275 10987 4309 11137
rect 4352 11027 4362 11079
rect 4414 11027 4424 11079
rect 4467 10987 4501 11137
rect 4544 11027 4554 11079
rect 4606 11027 4616 11079
rect 4659 10987 4693 11137
rect 4736 11027 4746 11079
rect 4798 11027 4808 11079
rect 4851 10987 4885 11137
rect 4928 11027 4938 11079
rect 4990 11027 5000 11079
rect 5055 11043 5101 11248
rect 5055 11009 5061 11043
rect 5095 11009 5101 11043
rect 3981 10940 4027 10987
rect 3981 10906 3987 10940
rect 4021 10906 4027 10940
rect 3981 10868 4027 10906
rect 3981 10834 3987 10868
rect 4021 10834 4027 10868
rect 3981 10796 4027 10834
rect 3981 10762 3987 10796
rect 4021 10762 4027 10796
rect 3981 10715 4027 10762
rect 4077 10940 4123 10987
rect 4077 10906 4083 10940
rect 4117 10906 4123 10940
rect 4077 10868 4123 10906
rect 4077 10834 4083 10868
rect 4117 10834 4123 10868
rect 4077 10796 4123 10834
rect 4077 10762 4083 10796
rect 4117 10762 4123 10796
rect 4077 10715 4123 10762
rect 4173 10940 4219 10987
rect 4173 10906 4179 10940
rect 4213 10906 4219 10940
rect 4173 10868 4219 10906
rect 4173 10834 4179 10868
rect 4213 10834 4219 10868
rect 4173 10796 4219 10834
rect 4173 10762 4179 10796
rect 4213 10762 4219 10796
rect 4173 10715 4219 10762
rect 4269 10940 4315 10987
rect 4269 10906 4275 10940
rect 4309 10906 4315 10940
rect 4269 10868 4315 10906
rect 4269 10834 4275 10868
rect 4309 10834 4315 10868
rect 4269 10796 4315 10834
rect 4269 10762 4275 10796
rect 4309 10762 4315 10796
rect 4269 10715 4315 10762
rect 4365 10940 4411 10987
rect 4365 10906 4371 10940
rect 4405 10906 4411 10940
rect 4365 10868 4411 10906
rect 4365 10834 4371 10868
rect 4405 10834 4411 10868
rect 4365 10796 4411 10834
rect 4365 10762 4371 10796
rect 4405 10762 4411 10796
rect 4365 10715 4411 10762
rect 4461 10940 4507 10987
rect 4461 10906 4467 10940
rect 4501 10906 4507 10940
rect 4461 10868 4507 10906
rect 4461 10834 4467 10868
rect 4501 10834 4507 10868
rect 4461 10796 4507 10834
rect 4461 10762 4467 10796
rect 4501 10762 4507 10796
rect 4461 10715 4507 10762
rect 4557 10940 4603 10987
rect 4557 10906 4563 10940
rect 4597 10906 4603 10940
rect 4557 10868 4603 10906
rect 4557 10834 4563 10868
rect 4597 10834 4603 10868
rect 4557 10796 4603 10834
rect 4557 10762 4563 10796
rect 4597 10762 4603 10796
rect 4557 10715 4603 10762
rect 4653 10940 4699 10987
rect 4653 10906 4659 10940
rect 4693 10906 4699 10940
rect 4653 10868 4699 10906
rect 4653 10834 4659 10868
rect 4693 10834 4699 10868
rect 4653 10796 4699 10834
rect 4653 10762 4659 10796
rect 4693 10762 4699 10796
rect 4653 10715 4699 10762
rect 4749 10940 4795 10987
rect 4749 10906 4755 10940
rect 4789 10906 4795 10940
rect 4749 10868 4795 10906
rect 4749 10834 4755 10868
rect 4789 10834 4795 10868
rect 4749 10796 4795 10834
rect 4749 10762 4755 10796
rect 4789 10762 4795 10796
rect 4749 10715 4795 10762
rect 4845 10940 4891 10987
rect 4845 10906 4851 10940
rect 4885 10906 4891 10940
rect 4845 10868 4891 10906
rect 4845 10834 4851 10868
rect 4885 10834 4891 10868
rect 4845 10796 4891 10834
rect 4845 10762 4851 10796
rect 4885 10762 4891 10796
rect 4845 10715 4891 10762
rect 4941 10940 4987 10987
rect 4941 10906 4947 10940
rect 4981 10906 4987 10940
rect 4941 10868 4987 10906
rect 4941 10834 4947 10868
rect 4981 10834 4987 10868
rect 4941 10796 4987 10834
rect 4941 10762 4947 10796
rect 4981 10762 4987 10796
rect 4941 10715 4987 10762
rect 5055 10971 5101 11009
rect 5055 10937 5061 10971
rect 5095 10937 5101 10971
rect 5055 10899 5101 10937
rect 5055 10865 5061 10899
rect 5095 10868 5101 10899
rect 5274 10868 5550 10869
rect 5095 10865 5550 10868
rect 5055 10838 5550 10865
rect 5055 10827 5303 10838
rect 5055 10793 5061 10827
rect 5095 10804 5303 10827
rect 5337 10804 5395 10838
rect 5429 10804 5487 10838
rect 5521 10804 5550 10838
rect 5095 10793 5550 10804
rect 5055 10773 5550 10793
rect 5055 10755 5101 10773
rect 5055 10721 5061 10755
rect 5095 10721 5101 10755
rect 2466 10540 3837 10574
rect 2466 10407 2500 10540
rect 2658 10407 2692 10540
rect 2850 10407 2884 10540
rect 3042 10407 3076 10540
rect 3234 10407 3268 10540
rect 3426 10407 3460 10540
rect 3671 10450 3681 10502
rect 3733 10450 3743 10502
rect 3679 10449 3691 10450
rect 3725 10449 3737 10450
rect 3679 10443 3737 10449
rect 3534 10414 3580 10437
rect 2460 10372 2506 10407
rect 2460 10338 2466 10372
rect 2500 10338 2506 10372
rect 2460 10303 2506 10338
rect 2556 10372 2602 10407
rect 2556 10338 2562 10372
rect 2596 10338 2602 10372
rect 2556 10303 2602 10338
rect 2652 10372 2698 10407
rect 2652 10338 2658 10372
rect 2692 10338 2698 10372
rect 2652 10303 2698 10338
rect 2748 10372 2794 10407
rect 2748 10338 2754 10372
rect 2788 10338 2794 10372
rect 2748 10303 2794 10338
rect 2844 10372 2890 10407
rect 2844 10338 2850 10372
rect 2884 10338 2890 10372
rect 2844 10303 2890 10338
rect 2940 10372 2986 10407
rect 2940 10338 2946 10372
rect 2980 10338 2986 10372
rect 2940 10303 2986 10338
rect 3036 10372 3082 10407
rect 3036 10338 3042 10372
rect 3076 10338 3082 10372
rect 3036 10303 3082 10338
rect 3132 10372 3178 10407
rect 3132 10338 3138 10372
rect 3172 10338 3178 10372
rect 3132 10303 3178 10338
rect 3228 10372 3274 10407
rect 3228 10338 3234 10372
rect 3268 10338 3274 10372
rect 3228 10303 3274 10338
rect 3324 10372 3370 10407
rect 3324 10338 3330 10372
rect 3364 10338 3370 10372
rect 3324 10303 3370 10338
rect 3420 10372 3466 10407
rect 3420 10338 3426 10372
rect 3460 10338 3466 10372
rect 3420 10303 3466 10338
rect 3534 10380 3540 10414
rect 3574 10412 3580 10414
rect 3803 10412 3837 10540
rect 3574 10411 3680 10412
rect 3734 10411 3837 10412
rect 3574 10399 3687 10411
rect 3574 10380 3647 10399
rect 3534 10342 3647 10380
rect 3534 10308 3540 10342
rect 3574 10323 3647 10342
rect 3681 10323 3687 10399
rect 3574 10312 3687 10323
rect 3574 10308 3580 10312
rect 3641 10311 3687 10312
rect 3729 10399 3837 10411
rect 3987 10574 4021 10715
rect 4179 10574 4213 10715
rect 4371 10574 4405 10715
rect 4563 10574 4597 10715
rect 4755 10574 4789 10715
rect 4947 10574 4981 10715
rect 5055 10677 5101 10721
rect 5683 10628 5743 11881
rect 5177 10594 5743 10628
rect 5177 10574 5211 10594
rect 3987 10540 5211 10574
rect 3987 10407 4021 10540
rect 4179 10407 4213 10540
rect 4371 10407 4405 10540
rect 4563 10407 4597 10540
rect 4755 10407 4789 10540
rect 4947 10407 4981 10540
rect 5438 10536 5512 10537
rect 5326 10534 5400 10535
rect 5326 10482 5337 10534
rect 5389 10482 5400 10534
rect 5438 10484 5449 10536
rect 5501 10484 5512 10536
rect 5438 10483 5512 10484
rect 5326 10481 5400 10482
rect 5055 10414 5101 10437
rect 3729 10323 3735 10399
rect 3769 10323 3837 10399
rect 3729 10312 3837 10323
rect 3729 10311 3775 10312
rect 2450 10272 2516 10275
rect 2447 10220 2457 10272
rect 2509 10220 2519 10272
rect 2450 10215 2516 10220
rect 2562 10163 2596 10303
rect 2642 10272 2708 10275
rect 2638 10220 2648 10272
rect 2700 10220 2710 10272
rect 2642 10215 2708 10220
rect 2754 10163 2788 10303
rect 2834 10272 2900 10275
rect 2830 10220 2840 10272
rect 2892 10220 2902 10272
rect 2834 10215 2900 10220
rect 2946 10163 2980 10303
rect 3026 10272 3092 10275
rect 3022 10220 3032 10272
rect 3084 10220 3094 10272
rect 3026 10215 3092 10220
rect 3138 10163 3172 10303
rect 3218 10271 3284 10275
rect 3215 10219 3225 10271
rect 3277 10219 3287 10271
rect 3218 10215 3284 10219
rect 3330 10163 3364 10303
rect 3410 10271 3476 10275
rect 3407 10219 3417 10271
rect 3469 10219 3479 10271
rect 3534 10270 3580 10308
rect 3534 10236 3540 10270
rect 3574 10236 3580 10270
rect 3410 10215 3476 10219
rect 2282 10129 3364 10163
rect 3534 10053 3580 10236
rect 3803 10163 3837 10312
rect 3981 10372 4027 10407
rect 3981 10338 3987 10372
rect 4021 10338 4027 10372
rect 3981 10303 4027 10338
rect 4077 10372 4123 10407
rect 4077 10338 4083 10372
rect 4117 10338 4123 10372
rect 4077 10303 4123 10338
rect 4173 10372 4219 10407
rect 4173 10338 4179 10372
rect 4213 10338 4219 10372
rect 4173 10303 4219 10338
rect 4269 10372 4315 10407
rect 4269 10338 4275 10372
rect 4309 10338 4315 10372
rect 4269 10303 4315 10338
rect 4365 10372 4411 10407
rect 4365 10338 4371 10372
rect 4405 10338 4411 10372
rect 4365 10303 4411 10338
rect 4461 10372 4507 10407
rect 4461 10338 4467 10372
rect 4501 10338 4507 10372
rect 4461 10303 4507 10338
rect 4557 10372 4603 10407
rect 4557 10338 4563 10372
rect 4597 10338 4603 10372
rect 4557 10303 4603 10338
rect 4653 10372 4699 10407
rect 4653 10338 4659 10372
rect 4693 10338 4699 10372
rect 4653 10303 4699 10338
rect 4749 10372 4795 10407
rect 4749 10338 4755 10372
rect 4789 10338 4795 10372
rect 4749 10303 4795 10338
rect 4845 10372 4891 10407
rect 4845 10338 4851 10372
rect 4885 10338 4891 10372
rect 4845 10303 4891 10338
rect 4941 10372 4987 10407
rect 4941 10338 4947 10372
rect 4981 10338 4987 10372
rect 4941 10303 4987 10338
rect 5055 10380 5061 10414
rect 5095 10380 5101 10414
rect 5055 10342 5101 10380
rect 5055 10308 5061 10342
rect 5095 10325 5101 10342
rect 5095 10308 5550 10325
rect 3971 10272 4037 10275
rect 3968 10220 3978 10272
rect 4030 10220 4040 10272
rect 3971 10215 4037 10220
rect 4083 10163 4117 10303
rect 4163 10272 4229 10275
rect 4159 10220 4169 10272
rect 4221 10220 4231 10272
rect 4163 10215 4229 10220
rect 4275 10163 4309 10303
rect 4355 10272 4421 10275
rect 4351 10220 4361 10272
rect 4413 10220 4423 10272
rect 4355 10215 4421 10220
rect 4467 10163 4501 10303
rect 4547 10272 4613 10275
rect 4543 10220 4553 10272
rect 4605 10220 4615 10272
rect 4547 10215 4613 10220
rect 4659 10163 4693 10303
rect 4739 10271 4805 10275
rect 4736 10219 4746 10271
rect 4798 10219 4808 10271
rect 4739 10215 4805 10219
rect 4851 10163 4885 10303
rect 5055 10294 5550 10308
rect 4931 10271 4997 10275
rect 4928 10219 4938 10271
rect 4990 10219 5000 10271
rect 5055 10270 5303 10294
rect 5055 10236 5061 10270
rect 5095 10260 5303 10270
rect 5337 10260 5395 10294
rect 5429 10260 5487 10294
rect 5521 10260 5550 10294
rect 5095 10236 5550 10260
rect 5055 10229 5550 10236
rect 4931 10215 4997 10219
rect 3803 10129 4885 10163
rect 5055 10054 5101 10229
rect 129 9846 1211 9880
rect 129 9283 163 9846
rect 294 9736 304 9788
rect 356 9736 366 9788
rect 409 9696 443 9846
rect 487 9736 497 9788
rect 549 9736 559 9788
rect 601 9696 635 9846
rect 678 9736 688 9788
rect 740 9736 750 9788
rect 793 9696 827 9846
rect 870 9736 880 9788
rect 932 9736 942 9788
rect 985 9696 1019 9846
rect 1062 9736 1072 9788
rect 1124 9736 1134 9788
rect 1177 9696 1211 9846
rect 1254 9736 1264 9788
rect 1316 9736 1326 9788
rect 1381 9752 1427 9916
rect 2282 9850 3364 9884
rect 1381 9718 1387 9752
rect 1421 9718 1427 9752
rect 1512 9729 1522 9789
rect 1578 9729 1792 9789
rect 1852 9729 1862 9789
rect 307 9649 353 9696
rect 307 9615 313 9649
rect 347 9615 353 9649
rect 307 9577 353 9615
rect 307 9543 313 9577
rect 347 9543 353 9577
rect 307 9505 353 9543
rect 307 9471 313 9505
rect 347 9471 353 9505
rect 307 9424 353 9471
rect 403 9649 449 9696
rect 403 9615 409 9649
rect 443 9615 449 9649
rect 403 9577 449 9615
rect 403 9543 409 9577
rect 443 9543 449 9577
rect 403 9505 449 9543
rect 403 9471 409 9505
rect 443 9471 449 9505
rect 403 9424 449 9471
rect 499 9649 545 9696
rect 499 9615 505 9649
rect 539 9615 545 9649
rect 499 9577 545 9615
rect 499 9543 505 9577
rect 539 9543 545 9577
rect 499 9505 545 9543
rect 499 9471 505 9505
rect 539 9471 545 9505
rect 499 9424 545 9471
rect 595 9649 641 9696
rect 595 9615 601 9649
rect 635 9615 641 9649
rect 595 9577 641 9615
rect 595 9543 601 9577
rect 635 9543 641 9577
rect 595 9505 641 9543
rect 595 9471 601 9505
rect 635 9471 641 9505
rect 595 9424 641 9471
rect 691 9649 737 9696
rect 691 9615 697 9649
rect 731 9615 737 9649
rect 691 9577 737 9615
rect 691 9543 697 9577
rect 731 9543 737 9577
rect 691 9505 737 9543
rect 691 9471 697 9505
rect 731 9471 737 9505
rect 691 9424 737 9471
rect 787 9649 833 9696
rect 787 9615 793 9649
rect 827 9615 833 9649
rect 787 9577 833 9615
rect 787 9543 793 9577
rect 827 9543 833 9577
rect 787 9505 833 9543
rect 787 9471 793 9505
rect 827 9471 833 9505
rect 787 9424 833 9471
rect 883 9649 929 9696
rect 883 9615 889 9649
rect 923 9615 929 9649
rect 883 9577 929 9615
rect 883 9543 889 9577
rect 923 9543 929 9577
rect 883 9505 929 9543
rect 883 9471 889 9505
rect 923 9471 929 9505
rect 883 9424 929 9471
rect 979 9649 1025 9696
rect 979 9615 985 9649
rect 1019 9615 1025 9649
rect 979 9577 1025 9615
rect 979 9543 985 9577
rect 1019 9543 1025 9577
rect 979 9505 1025 9543
rect 979 9471 985 9505
rect 1019 9471 1025 9505
rect 979 9424 1025 9471
rect 1075 9649 1121 9696
rect 1075 9615 1081 9649
rect 1115 9615 1121 9649
rect 1075 9577 1121 9615
rect 1075 9543 1081 9577
rect 1115 9543 1121 9577
rect 1075 9505 1121 9543
rect 1075 9471 1081 9505
rect 1115 9471 1121 9505
rect 1075 9424 1121 9471
rect 1171 9649 1217 9696
rect 1171 9615 1177 9649
rect 1211 9615 1217 9649
rect 1171 9577 1217 9615
rect 1171 9543 1177 9577
rect 1211 9543 1217 9577
rect 1171 9505 1217 9543
rect 1171 9471 1177 9505
rect 1211 9471 1217 9505
rect 1171 9424 1217 9471
rect 1267 9649 1313 9696
rect 1267 9615 1273 9649
rect 1307 9615 1313 9649
rect 1267 9577 1313 9615
rect 1267 9543 1273 9577
rect 1307 9543 1313 9577
rect 1267 9505 1313 9543
rect 1267 9471 1273 9505
rect 1307 9471 1313 9505
rect 1267 9424 1313 9471
rect 1381 9680 1427 9718
rect 1381 9646 1387 9680
rect 1421 9646 1427 9680
rect 1381 9608 1427 9646
rect 1381 9574 1387 9608
rect 1421 9574 1427 9608
rect 1381 9536 1427 9574
rect 1381 9502 1387 9536
rect 1421 9502 1427 9536
rect 1381 9492 1427 9502
rect 1381 9490 2160 9492
rect 1381 9464 2056 9490
rect 1381 9439 1387 9464
rect 1380 9430 1387 9439
rect 1421 9430 2056 9464
rect 0 9249 163 9283
rect 129 8872 163 9249
rect 313 9283 347 9424
rect 505 9283 539 9424
rect 697 9283 731 9424
rect 889 9283 923 9424
rect 1081 9283 1115 9424
rect 1273 9283 1307 9424
rect 1380 9382 2056 9430
rect 2190 9382 2200 9490
rect 1380 9380 2160 9382
rect 2282 9287 2316 9850
rect 2447 9740 2457 9792
rect 2509 9740 2519 9792
rect 2562 9700 2596 9850
rect 2640 9740 2650 9792
rect 2702 9740 2712 9792
rect 2754 9700 2788 9850
rect 2831 9740 2841 9792
rect 2893 9740 2903 9792
rect 2946 9700 2980 9850
rect 3023 9740 3033 9792
rect 3085 9740 3095 9792
rect 3138 9700 3172 9850
rect 3215 9740 3225 9792
rect 3277 9740 3287 9792
rect 3330 9700 3364 9850
rect 3407 9740 3417 9792
rect 3469 9740 3479 9792
rect 3534 9756 3580 9964
rect 3534 9722 3540 9756
rect 3574 9722 3580 9756
rect 2460 9653 2506 9700
rect 2460 9619 2466 9653
rect 2500 9619 2506 9653
rect 2460 9581 2506 9619
rect 2460 9547 2466 9581
rect 2500 9547 2506 9581
rect 2460 9509 2506 9547
rect 2460 9475 2466 9509
rect 2500 9475 2506 9509
rect 2460 9428 2506 9475
rect 2556 9653 2602 9700
rect 2556 9619 2562 9653
rect 2596 9619 2602 9653
rect 2556 9581 2602 9619
rect 2556 9547 2562 9581
rect 2596 9547 2602 9581
rect 2556 9509 2602 9547
rect 2556 9475 2562 9509
rect 2596 9475 2602 9509
rect 2556 9428 2602 9475
rect 2652 9653 2698 9700
rect 2652 9619 2658 9653
rect 2692 9619 2698 9653
rect 2652 9581 2698 9619
rect 2652 9547 2658 9581
rect 2692 9547 2698 9581
rect 2652 9509 2698 9547
rect 2652 9475 2658 9509
rect 2692 9475 2698 9509
rect 2652 9428 2698 9475
rect 2748 9653 2794 9700
rect 2748 9619 2754 9653
rect 2788 9619 2794 9653
rect 2748 9581 2794 9619
rect 2748 9547 2754 9581
rect 2788 9547 2794 9581
rect 2748 9509 2794 9547
rect 2748 9475 2754 9509
rect 2788 9475 2794 9509
rect 2748 9428 2794 9475
rect 2844 9653 2890 9700
rect 2844 9619 2850 9653
rect 2884 9619 2890 9653
rect 2844 9581 2890 9619
rect 2844 9547 2850 9581
rect 2884 9547 2890 9581
rect 2844 9509 2890 9547
rect 2844 9475 2850 9509
rect 2884 9475 2890 9509
rect 2844 9428 2890 9475
rect 2940 9653 2986 9700
rect 2940 9619 2946 9653
rect 2980 9619 2986 9653
rect 2940 9581 2986 9619
rect 2940 9547 2946 9581
rect 2980 9547 2986 9581
rect 2940 9509 2986 9547
rect 2940 9475 2946 9509
rect 2980 9475 2986 9509
rect 2940 9428 2986 9475
rect 3036 9653 3082 9700
rect 3036 9619 3042 9653
rect 3076 9619 3082 9653
rect 3036 9581 3082 9619
rect 3036 9547 3042 9581
rect 3076 9547 3082 9581
rect 3036 9509 3082 9547
rect 3036 9475 3042 9509
rect 3076 9475 3082 9509
rect 3036 9428 3082 9475
rect 3132 9653 3178 9700
rect 3132 9619 3138 9653
rect 3172 9619 3178 9653
rect 3132 9581 3178 9619
rect 3132 9547 3138 9581
rect 3172 9547 3178 9581
rect 3132 9509 3178 9547
rect 3132 9475 3138 9509
rect 3172 9475 3178 9509
rect 3132 9428 3178 9475
rect 3228 9653 3274 9700
rect 3228 9619 3234 9653
rect 3268 9619 3274 9653
rect 3228 9581 3274 9619
rect 3228 9547 3234 9581
rect 3268 9547 3274 9581
rect 3228 9509 3274 9547
rect 3228 9475 3234 9509
rect 3268 9475 3274 9509
rect 3228 9428 3274 9475
rect 3324 9653 3370 9700
rect 3324 9619 3330 9653
rect 3364 9619 3370 9653
rect 3324 9581 3370 9619
rect 3324 9547 3330 9581
rect 3364 9547 3370 9581
rect 3324 9509 3370 9547
rect 3324 9475 3330 9509
rect 3364 9475 3370 9509
rect 3324 9428 3370 9475
rect 3420 9653 3466 9700
rect 3420 9619 3426 9653
rect 3460 9619 3466 9653
rect 3420 9581 3466 9619
rect 3420 9547 3426 9581
rect 3460 9547 3466 9581
rect 3420 9509 3466 9547
rect 3420 9475 3426 9509
rect 3460 9475 3466 9509
rect 3420 9428 3466 9475
rect 3534 9684 3580 9722
rect 3534 9650 3540 9684
rect 3574 9650 3580 9684
rect 3534 9612 3580 9650
rect 3534 9578 3540 9612
rect 3574 9578 3580 9612
rect 3534 9540 3580 9578
rect 3534 9506 3540 9540
rect 3574 9506 3580 9540
rect 3534 9468 3580 9506
rect 3534 9434 3540 9468
rect 3574 9434 3580 9468
rect 2101 9283 2316 9287
rect 313 9253 2316 9283
rect 313 9249 2141 9253
rect 313 9116 347 9249
rect 505 9116 539 9249
rect 697 9116 731 9249
rect 889 9116 923 9249
rect 1081 9116 1115 9249
rect 1273 9116 1307 9249
rect 1381 9123 1608 9146
rect 307 9081 353 9116
rect 307 9047 313 9081
rect 347 9047 353 9081
rect 307 9012 353 9047
rect 403 9081 449 9116
rect 403 9047 409 9081
rect 443 9047 449 9081
rect 403 9012 449 9047
rect 499 9081 545 9116
rect 499 9047 505 9081
rect 539 9047 545 9081
rect 499 9012 545 9047
rect 595 9081 641 9116
rect 595 9047 601 9081
rect 635 9047 641 9081
rect 595 9012 641 9047
rect 691 9081 737 9116
rect 691 9047 697 9081
rect 731 9047 737 9081
rect 691 9012 737 9047
rect 787 9081 833 9116
rect 787 9047 793 9081
rect 827 9047 833 9081
rect 787 9012 833 9047
rect 883 9081 929 9116
rect 883 9047 889 9081
rect 923 9047 929 9081
rect 883 9012 929 9047
rect 979 9081 1025 9116
rect 979 9047 985 9081
rect 1019 9047 1025 9081
rect 979 9012 1025 9047
rect 1075 9081 1121 9116
rect 1075 9047 1081 9081
rect 1115 9047 1121 9081
rect 1075 9012 1121 9047
rect 1171 9081 1217 9116
rect 1171 9047 1177 9081
rect 1211 9047 1217 9081
rect 1171 9012 1217 9047
rect 1267 9081 1313 9116
rect 1267 9047 1273 9081
rect 1307 9047 1313 9081
rect 1267 9012 1313 9047
rect 1381 9089 1387 9123
rect 1421 9089 1608 9123
rect 1381 9051 1608 9089
rect 1381 9017 1387 9051
rect 1421 9026 1608 9051
rect 1421 9017 1427 9026
rect 1560 9024 1608 9026
rect 1598 9022 1608 9024
rect 1720 9022 1730 9146
rect 297 8981 363 8984
rect 294 8929 304 8981
rect 356 8929 366 8981
rect 297 8924 363 8929
rect 409 8872 443 9012
rect 489 8981 555 8984
rect 485 8929 495 8981
rect 547 8929 557 8981
rect 489 8924 555 8929
rect 601 8872 635 9012
rect 681 8981 747 8984
rect 677 8929 687 8981
rect 739 8929 749 8981
rect 681 8924 747 8929
rect 793 8872 827 9012
rect 873 8981 939 8984
rect 869 8929 879 8981
rect 931 8929 941 8981
rect 873 8924 939 8929
rect 985 8872 1019 9012
rect 1065 8980 1131 8984
rect 1062 8928 1072 8980
rect 1124 8928 1134 8980
rect 1065 8924 1131 8928
rect 1177 8872 1211 9012
rect 1257 8980 1323 8984
rect 1254 8928 1264 8980
rect 1316 8928 1326 8980
rect 1381 8979 1427 9017
rect 1920 8984 1930 8986
rect 1381 8945 1387 8979
rect 1421 8945 1427 8979
rect 1257 8924 1323 8928
rect 129 8838 1211 8872
rect 1381 8802 1427 8945
rect 1458 8928 1468 8984
rect 1524 8930 1930 8984
rect 1986 8930 1996 8986
rect 1524 8928 1986 8930
rect 2282 8876 2316 9253
rect 2466 9287 2500 9428
rect 2658 9287 2692 9428
rect 2850 9287 2884 9428
rect 3042 9287 3076 9428
rect 3234 9287 3268 9428
rect 3426 9287 3460 9428
rect 3534 9390 3580 9434
rect 3803 9850 4885 9884
rect 3803 9287 3837 9850
rect 3968 9740 3978 9792
rect 4030 9740 4040 9792
rect 4083 9700 4117 9850
rect 4161 9740 4171 9792
rect 4223 9740 4233 9792
rect 4275 9700 4309 9850
rect 4352 9740 4362 9792
rect 4414 9740 4424 9792
rect 4467 9700 4501 9850
rect 4544 9740 4554 9792
rect 4606 9740 4616 9792
rect 4659 9700 4693 9850
rect 4736 9740 4746 9792
rect 4798 9740 4808 9792
rect 4851 9700 4885 9850
rect 4928 9740 4938 9792
rect 4990 9740 5000 9792
rect 5055 9756 5101 9961
rect 5055 9722 5061 9756
rect 5095 9722 5101 9756
rect 3981 9653 4027 9700
rect 3981 9619 3987 9653
rect 4021 9619 4027 9653
rect 3981 9581 4027 9619
rect 3981 9547 3987 9581
rect 4021 9547 4027 9581
rect 3981 9509 4027 9547
rect 3981 9475 3987 9509
rect 4021 9475 4027 9509
rect 3981 9428 4027 9475
rect 4077 9653 4123 9700
rect 4077 9619 4083 9653
rect 4117 9619 4123 9653
rect 4077 9581 4123 9619
rect 4077 9547 4083 9581
rect 4117 9547 4123 9581
rect 4077 9509 4123 9547
rect 4077 9475 4083 9509
rect 4117 9475 4123 9509
rect 4077 9428 4123 9475
rect 4173 9653 4219 9700
rect 4173 9619 4179 9653
rect 4213 9619 4219 9653
rect 4173 9581 4219 9619
rect 4173 9547 4179 9581
rect 4213 9547 4219 9581
rect 4173 9509 4219 9547
rect 4173 9475 4179 9509
rect 4213 9475 4219 9509
rect 4173 9428 4219 9475
rect 4269 9653 4315 9700
rect 4269 9619 4275 9653
rect 4309 9619 4315 9653
rect 4269 9581 4315 9619
rect 4269 9547 4275 9581
rect 4309 9547 4315 9581
rect 4269 9509 4315 9547
rect 4269 9475 4275 9509
rect 4309 9475 4315 9509
rect 4269 9428 4315 9475
rect 4365 9653 4411 9700
rect 4365 9619 4371 9653
rect 4405 9619 4411 9653
rect 4365 9581 4411 9619
rect 4365 9547 4371 9581
rect 4405 9547 4411 9581
rect 4365 9509 4411 9547
rect 4365 9475 4371 9509
rect 4405 9475 4411 9509
rect 4365 9428 4411 9475
rect 4461 9653 4507 9700
rect 4461 9619 4467 9653
rect 4501 9619 4507 9653
rect 4461 9581 4507 9619
rect 4461 9547 4467 9581
rect 4501 9547 4507 9581
rect 4461 9509 4507 9547
rect 4461 9475 4467 9509
rect 4501 9475 4507 9509
rect 4461 9428 4507 9475
rect 4557 9653 4603 9700
rect 4557 9619 4563 9653
rect 4597 9619 4603 9653
rect 4557 9581 4603 9619
rect 4557 9547 4563 9581
rect 4597 9547 4603 9581
rect 4557 9509 4603 9547
rect 4557 9475 4563 9509
rect 4597 9475 4603 9509
rect 4557 9428 4603 9475
rect 4653 9653 4699 9700
rect 4653 9619 4659 9653
rect 4693 9619 4699 9653
rect 4653 9581 4699 9619
rect 4653 9547 4659 9581
rect 4693 9547 4699 9581
rect 4653 9509 4699 9547
rect 4653 9475 4659 9509
rect 4693 9475 4699 9509
rect 4653 9428 4699 9475
rect 4749 9653 4795 9700
rect 4749 9619 4755 9653
rect 4789 9619 4795 9653
rect 4749 9581 4795 9619
rect 4749 9547 4755 9581
rect 4789 9547 4795 9581
rect 4749 9509 4795 9547
rect 4749 9475 4755 9509
rect 4789 9475 4795 9509
rect 4749 9428 4795 9475
rect 4845 9653 4891 9700
rect 4845 9619 4851 9653
rect 4885 9619 4891 9653
rect 4845 9581 4891 9619
rect 4845 9547 4851 9581
rect 4885 9547 4891 9581
rect 4845 9509 4891 9547
rect 4845 9475 4851 9509
rect 4885 9475 4891 9509
rect 4845 9428 4891 9475
rect 4941 9653 4987 9700
rect 4941 9619 4947 9653
rect 4981 9619 4987 9653
rect 4941 9581 4987 9619
rect 4941 9547 4947 9581
rect 4981 9547 4987 9581
rect 4941 9509 4987 9547
rect 4941 9475 4947 9509
rect 4981 9475 4987 9509
rect 4941 9428 4987 9475
rect 5055 9684 5101 9722
rect 5055 9650 5061 9684
rect 5095 9650 5101 9684
rect 5055 9612 5101 9650
rect 5055 9578 5061 9612
rect 5095 9581 5101 9612
rect 5274 9581 5550 9582
rect 5095 9578 5550 9581
rect 5055 9551 5550 9578
rect 5055 9540 5303 9551
rect 5055 9506 5061 9540
rect 5095 9517 5303 9540
rect 5337 9517 5395 9551
rect 5429 9517 5487 9551
rect 5521 9517 5550 9551
rect 5095 9506 5550 9517
rect 5055 9486 5550 9506
rect 5055 9468 5101 9486
rect 5055 9434 5061 9468
rect 5095 9434 5101 9468
rect 2466 9253 3837 9287
rect 2466 9120 2500 9253
rect 2658 9120 2692 9253
rect 2850 9120 2884 9253
rect 3042 9120 3076 9253
rect 3234 9120 3268 9253
rect 3426 9120 3460 9253
rect 3671 9163 3681 9215
rect 3733 9163 3743 9215
rect 3679 9162 3691 9163
rect 3725 9162 3737 9163
rect 3679 9156 3737 9162
rect 3534 9127 3580 9150
rect 2460 9085 2506 9120
rect 2460 9051 2466 9085
rect 2500 9051 2506 9085
rect 2460 9016 2506 9051
rect 2556 9085 2602 9120
rect 2556 9051 2562 9085
rect 2596 9051 2602 9085
rect 2556 9016 2602 9051
rect 2652 9085 2698 9120
rect 2652 9051 2658 9085
rect 2692 9051 2698 9085
rect 2652 9016 2698 9051
rect 2748 9085 2794 9120
rect 2748 9051 2754 9085
rect 2788 9051 2794 9085
rect 2748 9016 2794 9051
rect 2844 9085 2890 9120
rect 2844 9051 2850 9085
rect 2884 9051 2890 9085
rect 2844 9016 2890 9051
rect 2940 9085 2986 9120
rect 2940 9051 2946 9085
rect 2980 9051 2986 9085
rect 2940 9016 2986 9051
rect 3036 9085 3082 9120
rect 3036 9051 3042 9085
rect 3076 9051 3082 9085
rect 3036 9016 3082 9051
rect 3132 9085 3178 9120
rect 3132 9051 3138 9085
rect 3172 9051 3178 9085
rect 3132 9016 3178 9051
rect 3228 9085 3274 9120
rect 3228 9051 3234 9085
rect 3268 9051 3274 9085
rect 3228 9016 3274 9051
rect 3324 9085 3370 9120
rect 3324 9051 3330 9085
rect 3364 9051 3370 9085
rect 3324 9016 3370 9051
rect 3420 9085 3466 9120
rect 3420 9051 3426 9085
rect 3460 9051 3466 9085
rect 3420 9016 3466 9051
rect 3534 9093 3540 9127
rect 3574 9125 3580 9127
rect 3803 9125 3837 9253
rect 3574 9124 3680 9125
rect 3734 9124 3837 9125
rect 3574 9112 3687 9124
rect 3574 9093 3647 9112
rect 3534 9055 3647 9093
rect 3534 9021 3540 9055
rect 3574 9036 3647 9055
rect 3681 9036 3687 9112
rect 3574 9025 3687 9036
rect 3574 9021 3580 9025
rect 3641 9024 3687 9025
rect 3729 9112 3837 9124
rect 3987 9287 4021 9428
rect 4179 9287 4213 9428
rect 4371 9287 4405 9428
rect 4563 9287 4597 9428
rect 4755 9287 4789 9428
rect 4947 9287 4981 9428
rect 5055 9390 5101 9434
rect 5683 9341 5743 10594
rect 5177 9307 5743 9341
rect 5177 9287 5211 9307
rect 3987 9253 5211 9287
rect 3987 9120 4021 9253
rect 4179 9120 4213 9253
rect 4371 9120 4405 9253
rect 4563 9120 4597 9253
rect 4755 9120 4789 9253
rect 4947 9120 4981 9253
rect 5438 9249 5512 9250
rect 5326 9247 5400 9248
rect 5326 9195 5337 9247
rect 5389 9195 5400 9247
rect 5438 9197 5449 9249
rect 5501 9197 5512 9249
rect 5438 9196 5512 9197
rect 5326 9194 5400 9195
rect 5055 9127 5101 9150
rect 3729 9036 3735 9112
rect 3769 9036 3837 9112
rect 3729 9025 3837 9036
rect 3729 9024 3775 9025
rect 2450 8985 2516 8988
rect 2447 8933 2457 8985
rect 2509 8933 2519 8985
rect 2450 8928 2516 8933
rect 2562 8876 2596 9016
rect 2642 8985 2708 8988
rect 2638 8933 2648 8985
rect 2700 8933 2710 8985
rect 2642 8928 2708 8933
rect 2754 8876 2788 9016
rect 2834 8985 2900 8988
rect 2830 8933 2840 8985
rect 2892 8933 2902 8985
rect 2834 8928 2900 8933
rect 2946 8876 2980 9016
rect 3026 8985 3092 8988
rect 3022 8933 3032 8985
rect 3084 8933 3094 8985
rect 3026 8928 3092 8933
rect 3138 8876 3172 9016
rect 3218 8984 3284 8988
rect 3215 8932 3225 8984
rect 3277 8932 3287 8984
rect 3218 8928 3284 8932
rect 3330 8876 3364 9016
rect 3410 8984 3476 8988
rect 3407 8932 3417 8984
rect 3469 8932 3479 8984
rect 3534 8983 3580 9021
rect 3534 8949 3540 8983
rect 3574 8949 3580 8983
rect 3410 8928 3476 8932
rect 2282 8842 3364 8876
rect 3534 8766 3580 8949
rect 3803 8876 3837 9025
rect 3981 9085 4027 9120
rect 3981 9051 3987 9085
rect 4021 9051 4027 9085
rect 3981 9016 4027 9051
rect 4077 9085 4123 9120
rect 4077 9051 4083 9085
rect 4117 9051 4123 9085
rect 4077 9016 4123 9051
rect 4173 9085 4219 9120
rect 4173 9051 4179 9085
rect 4213 9051 4219 9085
rect 4173 9016 4219 9051
rect 4269 9085 4315 9120
rect 4269 9051 4275 9085
rect 4309 9051 4315 9085
rect 4269 9016 4315 9051
rect 4365 9085 4411 9120
rect 4365 9051 4371 9085
rect 4405 9051 4411 9085
rect 4365 9016 4411 9051
rect 4461 9085 4507 9120
rect 4461 9051 4467 9085
rect 4501 9051 4507 9085
rect 4461 9016 4507 9051
rect 4557 9085 4603 9120
rect 4557 9051 4563 9085
rect 4597 9051 4603 9085
rect 4557 9016 4603 9051
rect 4653 9085 4699 9120
rect 4653 9051 4659 9085
rect 4693 9051 4699 9085
rect 4653 9016 4699 9051
rect 4749 9085 4795 9120
rect 4749 9051 4755 9085
rect 4789 9051 4795 9085
rect 4749 9016 4795 9051
rect 4845 9085 4891 9120
rect 4845 9051 4851 9085
rect 4885 9051 4891 9085
rect 4845 9016 4891 9051
rect 4941 9085 4987 9120
rect 4941 9051 4947 9085
rect 4981 9051 4987 9085
rect 4941 9016 4987 9051
rect 5055 9093 5061 9127
rect 5095 9093 5101 9127
rect 5055 9055 5101 9093
rect 5055 9021 5061 9055
rect 5095 9038 5101 9055
rect 5095 9021 5550 9038
rect 3971 8985 4037 8988
rect 3968 8933 3978 8985
rect 4030 8933 4040 8985
rect 3971 8928 4037 8933
rect 4083 8876 4117 9016
rect 4163 8985 4229 8988
rect 4159 8933 4169 8985
rect 4221 8933 4231 8985
rect 4163 8928 4229 8933
rect 4275 8876 4309 9016
rect 4355 8985 4421 8988
rect 4351 8933 4361 8985
rect 4413 8933 4423 8985
rect 4355 8928 4421 8933
rect 4467 8876 4501 9016
rect 4547 8985 4613 8988
rect 4543 8933 4553 8985
rect 4605 8933 4615 8985
rect 4547 8928 4613 8933
rect 4659 8876 4693 9016
rect 4739 8984 4805 8988
rect 4736 8932 4746 8984
rect 4798 8932 4808 8984
rect 4739 8928 4805 8932
rect 4851 8876 4885 9016
rect 5055 9007 5550 9021
rect 4931 8984 4997 8988
rect 4928 8932 4938 8984
rect 4990 8932 5000 8984
rect 5055 8983 5303 9007
rect 5055 8949 5061 8983
rect 5095 8973 5303 8983
rect 5337 8973 5395 9007
rect 5429 8973 5487 9007
rect 5521 8973 5550 9007
rect 5095 8949 5550 8973
rect 5055 8942 5550 8949
rect 4931 8928 4997 8932
rect 3803 8842 4885 8876
rect 5055 8767 5101 8942
rect 129 8559 1211 8593
rect 129 7996 163 8559
rect 294 8449 304 8501
rect 356 8449 366 8501
rect 409 8409 443 8559
rect 487 8449 497 8501
rect 549 8449 559 8501
rect 601 8409 635 8559
rect 678 8449 688 8501
rect 740 8449 750 8501
rect 793 8409 827 8559
rect 870 8449 880 8501
rect 932 8449 942 8501
rect 985 8409 1019 8559
rect 1062 8449 1072 8501
rect 1124 8449 1134 8501
rect 1177 8409 1211 8559
rect 1254 8449 1264 8501
rect 1316 8449 1326 8501
rect 1381 8465 1427 8629
rect 2282 8563 3364 8597
rect 1381 8431 1387 8465
rect 1421 8431 1427 8465
rect 1512 8442 1522 8502
rect 1578 8442 1792 8502
rect 1852 8442 1862 8502
rect 307 8362 353 8409
rect 307 8328 313 8362
rect 347 8328 353 8362
rect 307 8290 353 8328
rect 307 8256 313 8290
rect 347 8256 353 8290
rect 307 8218 353 8256
rect 307 8184 313 8218
rect 347 8184 353 8218
rect 307 8137 353 8184
rect 403 8362 449 8409
rect 403 8328 409 8362
rect 443 8328 449 8362
rect 403 8290 449 8328
rect 403 8256 409 8290
rect 443 8256 449 8290
rect 403 8218 449 8256
rect 403 8184 409 8218
rect 443 8184 449 8218
rect 403 8137 449 8184
rect 499 8362 545 8409
rect 499 8328 505 8362
rect 539 8328 545 8362
rect 499 8290 545 8328
rect 499 8256 505 8290
rect 539 8256 545 8290
rect 499 8218 545 8256
rect 499 8184 505 8218
rect 539 8184 545 8218
rect 499 8137 545 8184
rect 595 8362 641 8409
rect 595 8328 601 8362
rect 635 8328 641 8362
rect 595 8290 641 8328
rect 595 8256 601 8290
rect 635 8256 641 8290
rect 595 8218 641 8256
rect 595 8184 601 8218
rect 635 8184 641 8218
rect 595 8137 641 8184
rect 691 8362 737 8409
rect 691 8328 697 8362
rect 731 8328 737 8362
rect 691 8290 737 8328
rect 691 8256 697 8290
rect 731 8256 737 8290
rect 691 8218 737 8256
rect 691 8184 697 8218
rect 731 8184 737 8218
rect 691 8137 737 8184
rect 787 8362 833 8409
rect 787 8328 793 8362
rect 827 8328 833 8362
rect 787 8290 833 8328
rect 787 8256 793 8290
rect 827 8256 833 8290
rect 787 8218 833 8256
rect 787 8184 793 8218
rect 827 8184 833 8218
rect 787 8137 833 8184
rect 883 8362 929 8409
rect 883 8328 889 8362
rect 923 8328 929 8362
rect 883 8290 929 8328
rect 883 8256 889 8290
rect 923 8256 929 8290
rect 883 8218 929 8256
rect 883 8184 889 8218
rect 923 8184 929 8218
rect 883 8137 929 8184
rect 979 8362 1025 8409
rect 979 8328 985 8362
rect 1019 8328 1025 8362
rect 979 8290 1025 8328
rect 979 8256 985 8290
rect 1019 8256 1025 8290
rect 979 8218 1025 8256
rect 979 8184 985 8218
rect 1019 8184 1025 8218
rect 979 8137 1025 8184
rect 1075 8362 1121 8409
rect 1075 8328 1081 8362
rect 1115 8328 1121 8362
rect 1075 8290 1121 8328
rect 1075 8256 1081 8290
rect 1115 8256 1121 8290
rect 1075 8218 1121 8256
rect 1075 8184 1081 8218
rect 1115 8184 1121 8218
rect 1075 8137 1121 8184
rect 1171 8362 1217 8409
rect 1171 8328 1177 8362
rect 1211 8328 1217 8362
rect 1171 8290 1217 8328
rect 1171 8256 1177 8290
rect 1211 8256 1217 8290
rect 1171 8218 1217 8256
rect 1171 8184 1177 8218
rect 1211 8184 1217 8218
rect 1171 8137 1217 8184
rect 1267 8362 1313 8409
rect 1267 8328 1273 8362
rect 1307 8328 1313 8362
rect 1267 8290 1313 8328
rect 1267 8256 1273 8290
rect 1307 8256 1313 8290
rect 1267 8218 1313 8256
rect 1267 8184 1273 8218
rect 1307 8184 1313 8218
rect 1267 8137 1313 8184
rect 1381 8393 1427 8431
rect 1381 8359 1387 8393
rect 1421 8359 1427 8393
rect 1381 8321 1427 8359
rect 1381 8287 1387 8321
rect 1421 8287 1427 8321
rect 1381 8249 1427 8287
rect 1381 8215 1387 8249
rect 1421 8215 1427 8249
rect 1381 8205 1427 8215
rect 1381 8203 2160 8205
rect 1381 8177 2056 8203
rect 1381 8152 1387 8177
rect 1380 8143 1387 8152
rect 1421 8143 2056 8177
rect 0 7962 163 7996
rect 129 7585 163 7962
rect 313 7996 347 8137
rect 505 7996 539 8137
rect 697 7996 731 8137
rect 889 7996 923 8137
rect 1081 7996 1115 8137
rect 1273 7996 1307 8137
rect 1380 8095 2056 8143
rect 2190 8095 2200 8203
rect 1380 8093 2160 8095
rect 2282 8000 2316 8563
rect 2447 8453 2457 8505
rect 2509 8453 2519 8505
rect 2562 8413 2596 8563
rect 2640 8453 2650 8505
rect 2702 8453 2712 8505
rect 2754 8413 2788 8563
rect 2831 8453 2841 8505
rect 2893 8453 2903 8505
rect 2946 8413 2980 8563
rect 3023 8453 3033 8505
rect 3085 8453 3095 8505
rect 3138 8413 3172 8563
rect 3215 8453 3225 8505
rect 3277 8453 3287 8505
rect 3330 8413 3364 8563
rect 3407 8453 3417 8505
rect 3469 8453 3479 8505
rect 3534 8469 3580 8677
rect 3534 8435 3540 8469
rect 3574 8435 3580 8469
rect 2460 8366 2506 8413
rect 2460 8332 2466 8366
rect 2500 8332 2506 8366
rect 2460 8294 2506 8332
rect 2460 8260 2466 8294
rect 2500 8260 2506 8294
rect 2460 8222 2506 8260
rect 2460 8188 2466 8222
rect 2500 8188 2506 8222
rect 2460 8141 2506 8188
rect 2556 8366 2602 8413
rect 2556 8332 2562 8366
rect 2596 8332 2602 8366
rect 2556 8294 2602 8332
rect 2556 8260 2562 8294
rect 2596 8260 2602 8294
rect 2556 8222 2602 8260
rect 2556 8188 2562 8222
rect 2596 8188 2602 8222
rect 2556 8141 2602 8188
rect 2652 8366 2698 8413
rect 2652 8332 2658 8366
rect 2692 8332 2698 8366
rect 2652 8294 2698 8332
rect 2652 8260 2658 8294
rect 2692 8260 2698 8294
rect 2652 8222 2698 8260
rect 2652 8188 2658 8222
rect 2692 8188 2698 8222
rect 2652 8141 2698 8188
rect 2748 8366 2794 8413
rect 2748 8332 2754 8366
rect 2788 8332 2794 8366
rect 2748 8294 2794 8332
rect 2748 8260 2754 8294
rect 2788 8260 2794 8294
rect 2748 8222 2794 8260
rect 2748 8188 2754 8222
rect 2788 8188 2794 8222
rect 2748 8141 2794 8188
rect 2844 8366 2890 8413
rect 2844 8332 2850 8366
rect 2884 8332 2890 8366
rect 2844 8294 2890 8332
rect 2844 8260 2850 8294
rect 2884 8260 2890 8294
rect 2844 8222 2890 8260
rect 2844 8188 2850 8222
rect 2884 8188 2890 8222
rect 2844 8141 2890 8188
rect 2940 8366 2986 8413
rect 2940 8332 2946 8366
rect 2980 8332 2986 8366
rect 2940 8294 2986 8332
rect 2940 8260 2946 8294
rect 2980 8260 2986 8294
rect 2940 8222 2986 8260
rect 2940 8188 2946 8222
rect 2980 8188 2986 8222
rect 2940 8141 2986 8188
rect 3036 8366 3082 8413
rect 3036 8332 3042 8366
rect 3076 8332 3082 8366
rect 3036 8294 3082 8332
rect 3036 8260 3042 8294
rect 3076 8260 3082 8294
rect 3036 8222 3082 8260
rect 3036 8188 3042 8222
rect 3076 8188 3082 8222
rect 3036 8141 3082 8188
rect 3132 8366 3178 8413
rect 3132 8332 3138 8366
rect 3172 8332 3178 8366
rect 3132 8294 3178 8332
rect 3132 8260 3138 8294
rect 3172 8260 3178 8294
rect 3132 8222 3178 8260
rect 3132 8188 3138 8222
rect 3172 8188 3178 8222
rect 3132 8141 3178 8188
rect 3228 8366 3274 8413
rect 3228 8332 3234 8366
rect 3268 8332 3274 8366
rect 3228 8294 3274 8332
rect 3228 8260 3234 8294
rect 3268 8260 3274 8294
rect 3228 8222 3274 8260
rect 3228 8188 3234 8222
rect 3268 8188 3274 8222
rect 3228 8141 3274 8188
rect 3324 8366 3370 8413
rect 3324 8332 3330 8366
rect 3364 8332 3370 8366
rect 3324 8294 3370 8332
rect 3324 8260 3330 8294
rect 3364 8260 3370 8294
rect 3324 8222 3370 8260
rect 3324 8188 3330 8222
rect 3364 8188 3370 8222
rect 3324 8141 3370 8188
rect 3420 8366 3466 8413
rect 3420 8332 3426 8366
rect 3460 8332 3466 8366
rect 3420 8294 3466 8332
rect 3420 8260 3426 8294
rect 3460 8260 3466 8294
rect 3420 8222 3466 8260
rect 3420 8188 3426 8222
rect 3460 8188 3466 8222
rect 3420 8141 3466 8188
rect 3534 8397 3580 8435
rect 3534 8363 3540 8397
rect 3574 8363 3580 8397
rect 3534 8325 3580 8363
rect 3534 8291 3540 8325
rect 3574 8291 3580 8325
rect 3534 8253 3580 8291
rect 3534 8219 3540 8253
rect 3574 8219 3580 8253
rect 3534 8181 3580 8219
rect 3534 8147 3540 8181
rect 3574 8147 3580 8181
rect 2101 7996 2316 8000
rect 313 7966 2316 7996
rect 313 7962 2141 7966
rect 313 7829 347 7962
rect 505 7829 539 7962
rect 697 7829 731 7962
rect 889 7829 923 7962
rect 1081 7829 1115 7962
rect 1273 7829 1307 7962
rect 1381 7836 1608 7859
rect 307 7794 353 7829
rect 307 7760 313 7794
rect 347 7760 353 7794
rect 307 7725 353 7760
rect 403 7794 449 7829
rect 403 7760 409 7794
rect 443 7760 449 7794
rect 403 7725 449 7760
rect 499 7794 545 7829
rect 499 7760 505 7794
rect 539 7760 545 7794
rect 499 7725 545 7760
rect 595 7794 641 7829
rect 595 7760 601 7794
rect 635 7760 641 7794
rect 595 7725 641 7760
rect 691 7794 737 7829
rect 691 7760 697 7794
rect 731 7760 737 7794
rect 691 7725 737 7760
rect 787 7794 833 7829
rect 787 7760 793 7794
rect 827 7760 833 7794
rect 787 7725 833 7760
rect 883 7794 929 7829
rect 883 7760 889 7794
rect 923 7760 929 7794
rect 883 7725 929 7760
rect 979 7794 1025 7829
rect 979 7760 985 7794
rect 1019 7760 1025 7794
rect 979 7725 1025 7760
rect 1075 7794 1121 7829
rect 1075 7760 1081 7794
rect 1115 7760 1121 7794
rect 1075 7725 1121 7760
rect 1171 7794 1217 7829
rect 1171 7760 1177 7794
rect 1211 7760 1217 7794
rect 1171 7725 1217 7760
rect 1267 7794 1313 7829
rect 1267 7760 1273 7794
rect 1307 7760 1313 7794
rect 1267 7725 1313 7760
rect 1381 7802 1387 7836
rect 1421 7802 1608 7836
rect 1381 7764 1608 7802
rect 1381 7730 1387 7764
rect 1421 7739 1608 7764
rect 1421 7730 1427 7739
rect 1560 7737 1608 7739
rect 1598 7735 1608 7737
rect 1720 7735 1730 7859
rect 297 7694 363 7697
rect 294 7642 304 7694
rect 356 7642 366 7694
rect 297 7637 363 7642
rect 409 7585 443 7725
rect 489 7694 555 7697
rect 485 7642 495 7694
rect 547 7642 557 7694
rect 489 7637 555 7642
rect 601 7585 635 7725
rect 681 7694 747 7697
rect 677 7642 687 7694
rect 739 7642 749 7694
rect 681 7637 747 7642
rect 793 7585 827 7725
rect 873 7694 939 7697
rect 869 7642 879 7694
rect 931 7642 941 7694
rect 873 7637 939 7642
rect 985 7585 1019 7725
rect 1065 7693 1131 7697
rect 1062 7641 1072 7693
rect 1124 7641 1134 7693
rect 1065 7637 1131 7641
rect 1177 7585 1211 7725
rect 1257 7693 1323 7697
rect 1254 7641 1264 7693
rect 1316 7641 1326 7693
rect 1381 7692 1427 7730
rect 1920 7697 1930 7699
rect 1381 7658 1387 7692
rect 1421 7658 1427 7692
rect 1257 7637 1323 7641
rect 129 7551 1211 7585
rect 1381 7515 1427 7658
rect 1458 7641 1468 7697
rect 1524 7643 1930 7697
rect 1986 7643 1996 7699
rect 1524 7641 1986 7643
rect 2282 7589 2316 7966
rect 2466 8000 2500 8141
rect 2658 8000 2692 8141
rect 2850 8000 2884 8141
rect 3042 8000 3076 8141
rect 3234 8000 3268 8141
rect 3426 8000 3460 8141
rect 3534 8103 3580 8147
rect 3803 8563 4885 8597
rect 3803 8000 3837 8563
rect 3968 8453 3978 8505
rect 4030 8453 4040 8505
rect 4083 8413 4117 8563
rect 4161 8453 4171 8505
rect 4223 8453 4233 8505
rect 4275 8413 4309 8563
rect 4352 8453 4362 8505
rect 4414 8453 4424 8505
rect 4467 8413 4501 8563
rect 4544 8453 4554 8505
rect 4606 8453 4616 8505
rect 4659 8413 4693 8563
rect 4736 8453 4746 8505
rect 4798 8453 4808 8505
rect 4851 8413 4885 8563
rect 4928 8453 4938 8505
rect 4990 8453 5000 8505
rect 5055 8469 5101 8674
rect 5055 8435 5061 8469
rect 5095 8435 5101 8469
rect 3981 8366 4027 8413
rect 3981 8332 3987 8366
rect 4021 8332 4027 8366
rect 3981 8294 4027 8332
rect 3981 8260 3987 8294
rect 4021 8260 4027 8294
rect 3981 8222 4027 8260
rect 3981 8188 3987 8222
rect 4021 8188 4027 8222
rect 3981 8141 4027 8188
rect 4077 8366 4123 8413
rect 4077 8332 4083 8366
rect 4117 8332 4123 8366
rect 4077 8294 4123 8332
rect 4077 8260 4083 8294
rect 4117 8260 4123 8294
rect 4077 8222 4123 8260
rect 4077 8188 4083 8222
rect 4117 8188 4123 8222
rect 4077 8141 4123 8188
rect 4173 8366 4219 8413
rect 4173 8332 4179 8366
rect 4213 8332 4219 8366
rect 4173 8294 4219 8332
rect 4173 8260 4179 8294
rect 4213 8260 4219 8294
rect 4173 8222 4219 8260
rect 4173 8188 4179 8222
rect 4213 8188 4219 8222
rect 4173 8141 4219 8188
rect 4269 8366 4315 8413
rect 4269 8332 4275 8366
rect 4309 8332 4315 8366
rect 4269 8294 4315 8332
rect 4269 8260 4275 8294
rect 4309 8260 4315 8294
rect 4269 8222 4315 8260
rect 4269 8188 4275 8222
rect 4309 8188 4315 8222
rect 4269 8141 4315 8188
rect 4365 8366 4411 8413
rect 4365 8332 4371 8366
rect 4405 8332 4411 8366
rect 4365 8294 4411 8332
rect 4365 8260 4371 8294
rect 4405 8260 4411 8294
rect 4365 8222 4411 8260
rect 4365 8188 4371 8222
rect 4405 8188 4411 8222
rect 4365 8141 4411 8188
rect 4461 8366 4507 8413
rect 4461 8332 4467 8366
rect 4501 8332 4507 8366
rect 4461 8294 4507 8332
rect 4461 8260 4467 8294
rect 4501 8260 4507 8294
rect 4461 8222 4507 8260
rect 4461 8188 4467 8222
rect 4501 8188 4507 8222
rect 4461 8141 4507 8188
rect 4557 8366 4603 8413
rect 4557 8332 4563 8366
rect 4597 8332 4603 8366
rect 4557 8294 4603 8332
rect 4557 8260 4563 8294
rect 4597 8260 4603 8294
rect 4557 8222 4603 8260
rect 4557 8188 4563 8222
rect 4597 8188 4603 8222
rect 4557 8141 4603 8188
rect 4653 8366 4699 8413
rect 4653 8332 4659 8366
rect 4693 8332 4699 8366
rect 4653 8294 4699 8332
rect 4653 8260 4659 8294
rect 4693 8260 4699 8294
rect 4653 8222 4699 8260
rect 4653 8188 4659 8222
rect 4693 8188 4699 8222
rect 4653 8141 4699 8188
rect 4749 8366 4795 8413
rect 4749 8332 4755 8366
rect 4789 8332 4795 8366
rect 4749 8294 4795 8332
rect 4749 8260 4755 8294
rect 4789 8260 4795 8294
rect 4749 8222 4795 8260
rect 4749 8188 4755 8222
rect 4789 8188 4795 8222
rect 4749 8141 4795 8188
rect 4845 8366 4891 8413
rect 4845 8332 4851 8366
rect 4885 8332 4891 8366
rect 4845 8294 4891 8332
rect 4845 8260 4851 8294
rect 4885 8260 4891 8294
rect 4845 8222 4891 8260
rect 4845 8188 4851 8222
rect 4885 8188 4891 8222
rect 4845 8141 4891 8188
rect 4941 8366 4987 8413
rect 4941 8332 4947 8366
rect 4981 8332 4987 8366
rect 4941 8294 4987 8332
rect 4941 8260 4947 8294
rect 4981 8260 4987 8294
rect 4941 8222 4987 8260
rect 4941 8188 4947 8222
rect 4981 8188 4987 8222
rect 4941 8141 4987 8188
rect 5055 8397 5101 8435
rect 5055 8363 5061 8397
rect 5095 8363 5101 8397
rect 5055 8325 5101 8363
rect 5055 8291 5061 8325
rect 5095 8294 5101 8325
rect 5274 8294 5550 8295
rect 5095 8291 5550 8294
rect 5055 8264 5550 8291
rect 5055 8253 5303 8264
rect 5055 8219 5061 8253
rect 5095 8230 5303 8253
rect 5337 8230 5395 8264
rect 5429 8230 5487 8264
rect 5521 8230 5550 8264
rect 5095 8219 5550 8230
rect 5055 8199 5550 8219
rect 5055 8181 5101 8199
rect 5055 8147 5061 8181
rect 5095 8147 5101 8181
rect 2466 7966 3837 8000
rect 2466 7833 2500 7966
rect 2658 7833 2692 7966
rect 2850 7833 2884 7966
rect 3042 7833 3076 7966
rect 3234 7833 3268 7966
rect 3426 7833 3460 7966
rect 3671 7876 3681 7928
rect 3733 7876 3743 7928
rect 3679 7875 3691 7876
rect 3725 7875 3737 7876
rect 3679 7869 3737 7875
rect 3534 7840 3580 7863
rect 2460 7798 2506 7833
rect 2460 7764 2466 7798
rect 2500 7764 2506 7798
rect 2460 7729 2506 7764
rect 2556 7798 2602 7833
rect 2556 7764 2562 7798
rect 2596 7764 2602 7798
rect 2556 7729 2602 7764
rect 2652 7798 2698 7833
rect 2652 7764 2658 7798
rect 2692 7764 2698 7798
rect 2652 7729 2698 7764
rect 2748 7798 2794 7833
rect 2748 7764 2754 7798
rect 2788 7764 2794 7798
rect 2748 7729 2794 7764
rect 2844 7798 2890 7833
rect 2844 7764 2850 7798
rect 2884 7764 2890 7798
rect 2844 7729 2890 7764
rect 2940 7798 2986 7833
rect 2940 7764 2946 7798
rect 2980 7764 2986 7798
rect 2940 7729 2986 7764
rect 3036 7798 3082 7833
rect 3036 7764 3042 7798
rect 3076 7764 3082 7798
rect 3036 7729 3082 7764
rect 3132 7798 3178 7833
rect 3132 7764 3138 7798
rect 3172 7764 3178 7798
rect 3132 7729 3178 7764
rect 3228 7798 3274 7833
rect 3228 7764 3234 7798
rect 3268 7764 3274 7798
rect 3228 7729 3274 7764
rect 3324 7798 3370 7833
rect 3324 7764 3330 7798
rect 3364 7764 3370 7798
rect 3324 7729 3370 7764
rect 3420 7798 3466 7833
rect 3420 7764 3426 7798
rect 3460 7764 3466 7798
rect 3420 7729 3466 7764
rect 3534 7806 3540 7840
rect 3574 7838 3580 7840
rect 3803 7838 3837 7966
rect 3574 7837 3680 7838
rect 3734 7837 3837 7838
rect 3574 7825 3687 7837
rect 3574 7806 3647 7825
rect 3534 7768 3647 7806
rect 3534 7734 3540 7768
rect 3574 7749 3647 7768
rect 3681 7749 3687 7825
rect 3574 7738 3687 7749
rect 3574 7734 3580 7738
rect 3641 7737 3687 7738
rect 3729 7825 3837 7837
rect 3987 8000 4021 8141
rect 4179 8000 4213 8141
rect 4371 8000 4405 8141
rect 4563 8000 4597 8141
rect 4755 8000 4789 8141
rect 4947 8000 4981 8141
rect 5055 8103 5101 8147
rect 5683 8054 5743 9307
rect 5177 8020 5743 8054
rect 5177 8000 5211 8020
rect 3987 7966 5211 8000
rect 3987 7833 4021 7966
rect 4179 7833 4213 7966
rect 4371 7833 4405 7966
rect 4563 7833 4597 7966
rect 4755 7833 4789 7966
rect 4947 7833 4981 7966
rect 5438 7962 5512 7963
rect 5326 7960 5400 7961
rect 5326 7908 5337 7960
rect 5389 7908 5400 7960
rect 5438 7910 5449 7962
rect 5501 7910 5512 7962
rect 5438 7909 5512 7910
rect 5326 7907 5400 7908
rect 5055 7840 5101 7863
rect 3729 7749 3735 7825
rect 3769 7749 3837 7825
rect 3729 7738 3837 7749
rect 3729 7737 3775 7738
rect 2450 7698 2516 7701
rect 2447 7646 2457 7698
rect 2509 7646 2519 7698
rect 2450 7641 2516 7646
rect 2562 7589 2596 7729
rect 2642 7698 2708 7701
rect 2638 7646 2648 7698
rect 2700 7646 2710 7698
rect 2642 7641 2708 7646
rect 2754 7589 2788 7729
rect 2834 7698 2900 7701
rect 2830 7646 2840 7698
rect 2892 7646 2902 7698
rect 2834 7641 2900 7646
rect 2946 7589 2980 7729
rect 3026 7698 3092 7701
rect 3022 7646 3032 7698
rect 3084 7646 3094 7698
rect 3026 7641 3092 7646
rect 3138 7589 3172 7729
rect 3218 7697 3284 7701
rect 3215 7645 3225 7697
rect 3277 7645 3287 7697
rect 3218 7641 3284 7645
rect 3330 7589 3364 7729
rect 3410 7697 3476 7701
rect 3407 7645 3417 7697
rect 3469 7645 3479 7697
rect 3534 7696 3580 7734
rect 3534 7662 3540 7696
rect 3574 7662 3580 7696
rect 3410 7641 3476 7645
rect 2282 7555 3364 7589
rect 3534 7479 3580 7662
rect 3803 7589 3837 7738
rect 3981 7798 4027 7833
rect 3981 7764 3987 7798
rect 4021 7764 4027 7798
rect 3981 7729 4027 7764
rect 4077 7798 4123 7833
rect 4077 7764 4083 7798
rect 4117 7764 4123 7798
rect 4077 7729 4123 7764
rect 4173 7798 4219 7833
rect 4173 7764 4179 7798
rect 4213 7764 4219 7798
rect 4173 7729 4219 7764
rect 4269 7798 4315 7833
rect 4269 7764 4275 7798
rect 4309 7764 4315 7798
rect 4269 7729 4315 7764
rect 4365 7798 4411 7833
rect 4365 7764 4371 7798
rect 4405 7764 4411 7798
rect 4365 7729 4411 7764
rect 4461 7798 4507 7833
rect 4461 7764 4467 7798
rect 4501 7764 4507 7798
rect 4461 7729 4507 7764
rect 4557 7798 4603 7833
rect 4557 7764 4563 7798
rect 4597 7764 4603 7798
rect 4557 7729 4603 7764
rect 4653 7798 4699 7833
rect 4653 7764 4659 7798
rect 4693 7764 4699 7798
rect 4653 7729 4699 7764
rect 4749 7798 4795 7833
rect 4749 7764 4755 7798
rect 4789 7764 4795 7798
rect 4749 7729 4795 7764
rect 4845 7798 4891 7833
rect 4845 7764 4851 7798
rect 4885 7764 4891 7798
rect 4845 7729 4891 7764
rect 4941 7798 4987 7833
rect 4941 7764 4947 7798
rect 4981 7764 4987 7798
rect 4941 7729 4987 7764
rect 5055 7806 5061 7840
rect 5095 7806 5101 7840
rect 5055 7768 5101 7806
rect 5055 7734 5061 7768
rect 5095 7751 5101 7768
rect 5095 7734 5550 7751
rect 3971 7698 4037 7701
rect 3968 7646 3978 7698
rect 4030 7646 4040 7698
rect 3971 7641 4037 7646
rect 4083 7589 4117 7729
rect 4163 7698 4229 7701
rect 4159 7646 4169 7698
rect 4221 7646 4231 7698
rect 4163 7641 4229 7646
rect 4275 7589 4309 7729
rect 4355 7698 4421 7701
rect 4351 7646 4361 7698
rect 4413 7646 4423 7698
rect 4355 7641 4421 7646
rect 4467 7589 4501 7729
rect 4547 7698 4613 7701
rect 4543 7646 4553 7698
rect 4605 7646 4615 7698
rect 4547 7641 4613 7646
rect 4659 7589 4693 7729
rect 4739 7697 4805 7701
rect 4736 7645 4746 7697
rect 4798 7645 4808 7697
rect 4739 7641 4805 7645
rect 4851 7589 4885 7729
rect 5055 7720 5550 7734
rect 4931 7697 4997 7701
rect 4928 7645 4938 7697
rect 4990 7645 5000 7697
rect 5055 7696 5303 7720
rect 5055 7662 5061 7696
rect 5095 7686 5303 7696
rect 5337 7686 5395 7720
rect 5429 7686 5487 7720
rect 5521 7686 5550 7720
rect 5095 7662 5550 7686
rect 5055 7655 5550 7662
rect 4931 7641 4997 7645
rect 3803 7555 4885 7589
rect 5055 7480 5101 7655
rect 129 7272 1211 7306
rect 129 6709 163 7272
rect 294 7162 304 7214
rect 356 7162 366 7214
rect 409 7122 443 7272
rect 487 7162 497 7214
rect 549 7162 559 7214
rect 601 7122 635 7272
rect 678 7162 688 7214
rect 740 7162 750 7214
rect 793 7122 827 7272
rect 870 7162 880 7214
rect 932 7162 942 7214
rect 985 7122 1019 7272
rect 1062 7162 1072 7214
rect 1124 7162 1134 7214
rect 1177 7122 1211 7272
rect 1254 7162 1264 7214
rect 1316 7162 1326 7214
rect 1381 7178 1427 7342
rect 2282 7276 3364 7310
rect 1381 7144 1387 7178
rect 1421 7144 1427 7178
rect 1512 7155 1522 7215
rect 1578 7155 1792 7215
rect 1852 7155 1862 7215
rect 307 7075 353 7122
rect 307 7041 313 7075
rect 347 7041 353 7075
rect 307 7003 353 7041
rect 307 6969 313 7003
rect 347 6969 353 7003
rect 307 6931 353 6969
rect 307 6897 313 6931
rect 347 6897 353 6931
rect 307 6850 353 6897
rect 403 7075 449 7122
rect 403 7041 409 7075
rect 443 7041 449 7075
rect 403 7003 449 7041
rect 403 6969 409 7003
rect 443 6969 449 7003
rect 403 6931 449 6969
rect 403 6897 409 6931
rect 443 6897 449 6931
rect 403 6850 449 6897
rect 499 7075 545 7122
rect 499 7041 505 7075
rect 539 7041 545 7075
rect 499 7003 545 7041
rect 499 6969 505 7003
rect 539 6969 545 7003
rect 499 6931 545 6969
rect 499 6897 505 6931
rect 539 6897 545 6931
rect 499 6850 545 6897
rect 595 7075 641 7122
rect 595 7041 601 7075
rect 635 7041 641 7075
rect 595 7003 641 7041
rect 595 6969 601 7003
rect 635 6969 641 7003
rect 595 6931 641 6969
rect 595 6897 601 6931
rect 635 6897 641 6931
rect 595 6850 641 6897
rect 691 7075 737 7122
rect 691 7041 697 7075
rect 731 7041 737 7075
rect 691 7003 737 7041
rect 691 6969 697 7003
rect 731 6969 737 7003
rect 691 6931 737 6969
rect 691 6897 697 6931
rect 731 6897 737 6931
rect 691 6850 737 6897
rect 787 7075 833 7122
rect 787 7041 793 7075
rect 827 7041 833 7075
rect 787 7003 833 7041
rect 787 6969 793 7003
rect 827 6969 833 7003
rect 787 6931 833 6969
rect 787 6897 793 6931
rect 827 6897 833 6931
rect 787 6850 833 6897
rect 883 7075 929 7122
rect 883 7041 889 7075
rect 923 7041 929 7075
rect 883 7003 929 7041
rect 883 6969 889 7003
rect 923 6969 929 7003
rect 883 6931 929 6969
rect 883 6897 889 6931
rect 923 6897 929 6931
rect 883 6850 929 6897
rect 979 7075 1025 7122
rect 979 7041 985 7075
rect 1019 7041 1025 7075
rect 979 7003 1025 7041
rect 979 6969 985 7003
rect 1019 6969 1025 7003
rect 979 6931 1025 6969
rect 979 6897 985 6931
rect 1019 6897 1025 6931
rect 979 6850 1025 6897
rect 1075 7075 1121 7122
rect 1075 7041 1081 7075
rect 1115 7041 1121 7075
rect 1075 7003 1121 7041
rect 1075 6969 1081 7003
rect 1115 6969 1121 7003
rect 1075 6931 1121 6969
rect 1075 6897 1081 6931
rect 1115 6897 1121 6931
rect 1075 6850 1121 6897
rect 1171 7075 1217 7122
rect 1171 7041 1177 7075
rect 1211 7041 1217 7075
rect 1171 7003 1217 7041
rect 1171 6969 1177 7003
rect 1211 6969 1217 7003
rect 1171 6931 1217 6969
rect 1171 6897 1177 6931
rect 1211 6897 1217 6931
rect 1171 6850 1217 6897
rect 1267 7075 1313 7122
rect 1267 7041 1273 7075
rect 1307 7041 1313 7075
rect 1267 7003 1313 7041
rect 1267 6969 1273 7003
rect 1307 6969 1313 7003
rect 1267 6931 1313 6969
rect 1267 6897 1273 6931
rect 1307 6897 1313 6931
rect 1267 6850 1313 6897
rect 1381 7106 1427 7144
rect 1381 7072 1387 7106
rect 1421 7072 1427 7106
rect 1381 7034 1427 7072
rect 1381 7000 1387 7034
rect 1421 7000 1427 7034
rect 1381 6962 1427 7000
rect 1381 6928 1387 6962
rect 1421 6928 1427 6962
rect 1381 6918 1427 6928
rect 1381 6916 2160 6918
rect 1381 6890 2056 6916
rect 1381 6865 1387 6890
rect 1380 6856 1387 6865
rect 1421 6856 2056 6890
rect 0 6675 163 6709
rect 129 6298 163 6675
rect 313 6709 347 6850
rect 505 6709 539 6850
rect 697 6709 731 6850
rect 889 6709 923 6850
rect 1081 6709 1115 6850
rect 1273 6709 1307 6850
rect 1380 6808 2056 6856
rect 2190 6808 2200 6916
rect 1380 6806 2160 6808
rect 2282 6713 2316 7276
rect 2447 7166 2457 7218
rect 2509 7166 2519 7218
rect 2562 7126 2596 7276
rect 2640 7166 2650 7218
rect 2702 7166 2712 7218
rect 2754 7126 2788 7276
rect 2831 7166 2841 7218
rect 2893 7166 2903 7218
rect 2946 7126 2980 7276
rect 3023 7166 3033 7218
rect 3085 7166 3095 7218
rect 3138 7126 3172 7276
rect 3215 7166 3225 7218
rect 3277 7166 3287 7218
rect 3330 7126 3364 7276
rect 3407 7166 3417 7218
rect 3469 7166 3479 7218
rect 3534 7182 3580 7390
rect 3534 7148 3540 7182
rect 3574 7148 3580 7182
rect 2460 7079 2506 7126
rect 2460 7045 2466 7079
rect 2500 7045 2506 7079
rect 2460 7007 2506 7045
rect 2460 6973 2466 7007
rect 2500 6973 2506 7007
rect 2460 6935 2506 6973
rect 2460 6901 2466 6935
rect 2500 6901 2506 6935
rect 2460 6854 2506 6901
rect 2556 7079 2602 7126
rect 2556 7045 2562 7079
rect 2596 7045 2602 7079
rect 2556 7007 2602 7045
rect 2556 6973 2562 7007
rect 2596 6973 2602 7007
rect 2556 6935 2602 6973
rect 2556 6901 2562 6935
rect 2596 6901 2602 6935
rect 2556 6854 2602 6901
rect 2652 7079 2698 7126
rect 2652 7045 2658 7079
rect 2692 7045 2698 7079
rect 2652 7007 2698 7045
rect 2652 6973 2658 7007
rect 2692 6973 2698 7007
rect 2652 6935 2698 6973
rect 2652 6901 2658 6935
rect 2692 6901 2698 6935
rect 2652 6854 2698 6901
rect 2748 7079 2794 7126
rect 2748 7045 2754 7079
rect 2788 7045 2794 7079
rect 2748 7007 2794 7045
rect 2748 6973 2754 7007
rect 2788 6973 2794 7007
rect 2748 6935 2794 6973
rect 2748 6901 2754 6935
rect 2788 6901 2794 6935
rect 2748 6854 2794 6901
rect 2844 7079 2890 7126
rect 2844 7045 2850 7079
rect 2884 7045 2890 7079
rect 2844 7007 2890 7045
rect 2844 6973 2850 7007
rect 2884 6973 2890 7007
rect 2844 6935 2890 6973
rect 2844 6901 2850 6935
rect 2884 6901 2890 6935
rect 2844 6854 2890 6901
rect 2940 7079 2986 7126
rect 2940 7045 2946 7079
rect 2980 7045 2986 7079
rect 2940 7007 2986 7045
rect 2940 6973 2946 7007
rect 2980 6973 2986 7007
rect 2940 6935 2986 6973
rect 2940 6901 2946 6935
rect 2980 6901 2986 6935
rect 2940 6854 2986 6901
rect 3036 7079 3082 7126
rect 3036 7045 3042 7079
rect 3076 7045 3082 7079
rect 3036 7007 3082 7045
rect 3036 6973 3042 7007
rect 3076 6973 3082 7007
rect 3036 6935 3082 6973
rect 3036 6901 3042 6935
rect 3076 6901 3082 6935
rect 3036 6854 3082 6901
rect 3132 7079 3178 7126
rect 3132 7045 3138 7079
rect 3172 7045 3178 7079
rect 3132 7007 3178 7045
rect 3132 6973 3138 7007
rect 3172 6973 3178 7007
rect 3132 6935 3178 6973
rect 3132 6901 3138 6935
rect 3172 6901 3178 6935
rect 3132 6854 3178 6901
rect 3228 7079 3274 7126
rect 3228 7045 3234 7079
rect 3268 7045 3274 7079
rect 3228 7007 3274 7045
rect 3228 6973 3234 7007
rect 3268 6973 3274 7007
rect 3228 6935 3274 6973
rect 3228 6901 3234 6935
rect 3268 6901 3274 6935
rect 3228 6854 3274 6901
rect 3324 7079 3370 7126
rect 3324 7045 3330 7079
rect 3364 7045 3370 7079
rect 3324 7007 3370 7045
rect 3324 6973 3330 7007
rect 3364 6973 3370 7007
rect 3324 6935 3370 6973
rect 3324 6901 3330 6935
rect 3364 6901 3370 6935
rect 3324 6854 3370 6901
rect 3420 7079 3466 7126
rect 3420 7045 3426 7079
rect 3460 7045 3466 7079
rect 3420 7007 3466 7045
rect 3420 6973 3426 7007
rect 3460 6973 3466 7007
rect 3420 6935 3466 6973
rect 3420 6901 3426 6935
rect 3460 6901 3466 6935
rect 3420 6854 3466 6901
rect 3534 7110 3580 7148
rect 3534 7076 3540 7110
rect 3574 7076 3580 7110
rect 3534 7038 3580 7076
rect 3534 7004 3540 7038
rect 3574 7004 3580 7038
rect 3534 6966 3580 7004
rect 3534 6932 3540 6966
rect 3574 6932 3580 6966
rect 3534 6894 3580 6932
rect 3534 6860 3540 6894
rect 3574 6860 3580 6894
rect 2101 6709 2316 6713
rect 313 6679 2316 6709
rect 313 6675 2141 6679
rect 313 6542 347 6675
rect 505 6542 539 6675
rect 697 6542 731 6675
rect 889 6542 923 6675
rect 1081 6542 1115 6675
rect 1273 6542 1307 6675
rect 1381 6549 1608 6572
rect 307 6507 353 6542
rect 307 6473 313 6507
rect 347 6473 353 6507
rect 307 6438 353 6473
rect 403 6507 449 6542
rect 403 6473 409 6507
rect 443 6473 449 6507
rect 403 6438 449 6473
rect 499 6507 545 6542
rect 499 6473 505 6507
rect 539 6473 545 6507
rect 499 6438 545 6473
rect 595 6507 641 6542
rect 595 6473 601 6507
rect 635 6473 641 6507
rect 595 6438 641 6473
rect 691 6507 737 6542
rect 691 6473 697 6507
rect 731 6473 737 6507
rect 691 6438 737 6473
rect 787 6507 833 6542
rect 787 6473 793 6507
rect 827 6473 833 6507
rect 787 6438 833 6473
rect 883 6507 929 6542
rect 883 6473 889 6507
rect 923 6473 929 6507
rect 883 6438 929 6473
rect 979 6507 1025 6542
rect 979 6473 985 6507
rect 1019 6473 1025 6507
rect 979 6438 1025 6473
rect 1075 6507 1121 6542
rect 1075 6473 1081 6507
rect 1115 6473 1121 6507
rect 1075 6438 1121 6473
rect 1171 6507 1217 6542
rect 1171 6473 1177 6507
rect 1211 6473 1217 6507
rect 1171 6438 1217 6473
rect 1267 6507 1313 6542
rect 1267 6473 1273 6507
rect 1307 6473 1313 6507
rect 1267 6438 1313 6473
rect 1381 6515 1387 6549
rect 1421 6515 1608 6549
rect 1381 6477 1608 6515
rect 1381 6443 1387 6477
rect 1421 6452 1608 6477
rect 1421 6443 1427 6452
rect 1560 6450 1608 6452
rect 1598 6448 1608 6450
rect 1720 6448 1730 6572
rect 297 6407 363 6410
rect 294 6355 304 6407
rect 356 6355 366 6407
rect 297 6350 363 6355
rect 409 6298 443 6438
rect 489 6407 555 6410
rect 485 6355 495 6407
rect 547 6355 557 6407
rect 489 6350 555 6355
rect 601 6298 635 6438
rect 681 6407 747 6410
rect 677 6355 687 6407
rect 739 6355 749 6407
rect 681 6350 747 6355
rect 793 6298 827 6438
rect 873 6407 939 6410
rect 869 6355 879 6407
rect 931 6355 941 6407
rect 873 6350 939 6355
rect 985 6298 1019 6438
rect 1065 6406 1131 6410
rect 1062 6354 1072 6406
rect 1124 6354 1134 6406
rect 1065 6350 1131 6354
rect 1177 6298 1211 6438
rect 1257 6406 1323 6410
rect 1254 6354 1264 6406
rect 1316 6354 1326 6406
rect 1381 6405 1427 6443
rect 1920 6410 1930 6412
rect 1381 6371 1387 6405
rect 1421 6371 1427 6405
rect 1257 6350 1323 6354
rect 129 6264 1211 6298
rect 1381 6228 1427 6371
rect 1458 6354 1468 6410
rect 1524 6356 1930 6410
rect 1986 6356 1996 6412
rect 1524 6354 1986 6356
rect 2282 6302 2316 6679
rect 2466 6713 2500 6854
rect 2658 6713 2692 6854
rect 2850 6713 2884 6854
rect 3042 6713 3076 6854
rect 3234 6713 3268 6854
rect 3426 6713 3460 6854
rect 3534 6816 3580 6860
rect 3803 7276 4885 7310
rect 3803 6713 3837 7276
rect 3968 7166 3978 7218
rect 4030 7166 4040 7218
rect 4083 7126 4117 7276
rect 4161 7166 4171 7218
rect 4223 7166 4233 7218
rect 4275 7126 4309 7276
rect 4352 7166 4362 7218
rect 4414 7166 4424 7218
rect 4467 7126 4501 7276
rect 4544 7166 4554 7218
rect 4606 7166 4616 7218
rect 4659 7126 4693 7276
rect 4736 7166 4746 7218
rect 4798 7166 4808 7218
rect 4851 7126 4885 7276
rect 4928 7166 4938 7218
rect 4990 7166 5000 7218
rect 5055 7182 5101 7387
rect 5055 7148 5061 7182
rect 5095 7148 5101 7182
rect 3981 7079 4027 7126
rect 3981 7045 3987 7079
rect 4021 7045 4027 7079
rect 3981 7007 4027 7045
rect 3981 6973 3987 7007
rect 4021 6973 4027 7007
rect 3981 6935 4027 6973
rect 3981 6901 3987 6935
rect 4021 6901 4027 6935
rect 3981 6854 4027 6901
rect 4077 7079 4123 7126
rect 4077 7045 4083 7079
rect 4117 7045 4123 7079
rect 4077 7007 4123 7045
rect 4077 6973 4083 7007
rect 4117 6973 4123 7007
rect 4077 6935 4123 6973
rect 4077 6901 4083 6935
rect 4117 6901 4123 6935
rect 4077 6854 4123 6901
rect 4173 7079 4219 7126
rect 4173 7045 4179 7079
rect 4213 7045 4219 7079
rect 4173 7007 4219 7045
rect 4173 6973 4179 7007
rect 4213 6973 4219 7007
rect 4173 6935 4219 6973
rect 4173 6901 4179 6935
rect 4213 6901 4219 6935
rect 4173 6854 4219 6901
rect 4269 7079 4315 7126
rect 4269 7045 4275 7079
rect 4309 7045 4315 7079
rect 4269 7007 4315 7045
rect 4269 6973 4275 7007
rect 4309 6973 4315 7007
rect 4269 6935 4315 6973
rect 4269 6901 4275 6935
rect 4309 6901 4315 6935
rect 4269 6854 4315 6901
rect 4365 7079 4411 7126
rect 4365 7045 4371 7079
rect 4405 7045 4411 7079
rect 4365 7007 4411 7045
rect 4365 6973 4371 7007
rect 4405 6973 4411 7007
rect 4365 6935 4411 6973
rect 4365 6901 4371 6935
rect 4405 6901 4411 6935
rect 4365 6854 4411 6901
rect 4461 7079 4507 7126
rect 4461 7045 4467 7079
rect 4501 7045 4507 7079
rect 4461 7007 4507 7045
rect 4461 6973 4467 7007
rect 4501 6973 4507 7007
rect 4461 6935 4507 6973
rect 4461 6901 4467 6935
rect 4501 6901 4507 6935
rect 4461 6854 4507 6901
rect 4557 7079 4603 7126
rect 4557 7045 4563 7079
rect 4597 7045 4603 7079
rect 4557 7007 4603 7045
rect 4557 6973 4563 7007
rect 4597 6973 4603 7007
rect 4557 6935 4603 6973
rect 4557 6901 4563 6935
rect 4597 6901 4603 6935
rect 4557 6854 4603 6901
rect 4653 7079 4699 7126
rect 4653 7045 4659 7079
rect 4693 7045 4699 7079
rect 4653 7007 4699 7045
rect 4653 6973 4659 7007
rect 4693 6973 4699 7007
rect 4653 6935 4699 6973
rect 4653 6901 4659 6935
rect 4693 6901 4699 6935
rect 4653 6854 4699 6901
rect 4749 7079 4795 7126
rect 4749 7045 4755 7079
rect 4789 7045 4795 7079
rect 4749 7007 4795 7045
rect 4749 6973 4755 7007
rect 4789 6973 4795 7007
rect 4749 6935 4795 6973
rect 4749 6901 4755 6935
rect 4789 6901 4795 6935
rect 4749 6854 4795 6901
rect 4845 7079 4891 7126
rect 4845 7045 4851 7079
rect 4885 7045 4891 7079
rect 4845 7007 4891 7045
rect 4845 6973 4851 7007
rect 4885 6973 4891 7007
rect 4845 6935 4891 6973
rect 4845 6901 4851 6935
rect 4885 6901 4891 6935
rect 4845 6854 4891 6901
rect 4941 7079 4987 7126
rect 4941 7045 4947 7079
rect 4981 7045 4987 7079
rect 4941 7007 4987 7045
rect 4941 6973 4947 7007
rect 4981 6973 4987 7007
rect 4941 6935 4987 6973
rect 4941 6901 4947 6935
rect 4981 6901 4987 6935
rect 4941 6854 4987 6901
rect 5055 7110 5101 7148
rect 5055 7076 5061 7110
rect 5095 7076 5101 7110
rect 5055 7038 5101 7076
rect 5055 7004 5061 7038
rect 5095 7007 5101 7038
rect 5274 7007 5550 7008
rect 5095 7004 5550 7007
rect 5055 6977 5550 7004
rect 5055 6966 5303 6977
rect 5055 6932 5061 6966
rect 5095 6943 5303 6966
rect 5337 6943 5395 6977
rect 5429 6943 5487 6977
rect 5521 6943 5550 6977
rect 5095 6932 5550 6943
rect 5055 6912 5550 6932
rect 5055 6894 5101 6912
rect 5055 6860 5061 6894
rect 5095 6860 5101 6894
rect 2466 6679 3837 6713
rect 2466 6546 2500 6679
rect 2658 6546 2692 6679
rect 2850 6546 2884 6679
rect 3042 6546 3076 6679
rect 3234 6546 3268 6679
rect 3426 6546 3460 6679
rect 3671 6589 3681 6641
rect 3733 6589 3743 6641
rect 3679 6588 3691 6589
rect 3725 6588 3737 6589
rect 3679 6582 3737 6588
rect 3534 6553 3580 6576
rect 2460 6511 2506 6546
rect 2460 6477 2466 6511
rect 2500 6477 2506 6511
rect 2460 6442 2506 6477
rect 2556 6511 2602 6546
rect 2556 6477 2562 6511
rect 2596 6477 2602 6511
rect 2556 6442 2602 6477
rect 2652 6511 2698 6546
rect 2652 6477 2658 6511
rect 2692 6477 2698 6511
rect 2652 6442 2698 6477
rect 2748 6511 2794 6546
rect 2748 6477 2754 6511
rect 2788 6477 2794 6511
rect 2748 6442 2794 6477
rect 2844 6511 2890 6546
rect 2844 6477 2850 6511
rect 2884 6477 2890 6511
rect 2844 6442 2890 6477
rect 2940 6511 2986 6546
rect 2940 6477 2946 6511
rect 2980 6477 2986 6511
rect 2940 6442 2986 6477
rect 3036 6511 3082 6546
rect 3036 6477 3042 6511
rect 3076 6477 3082 6511
rect 3036 6442 3082 6477
rect 3132 6511 3178 6546
rect 3132 6477 3138 6511
rect 3172 6477 3178 6511
rect 3132 6442 3178 6477
rect 3228 6511 3274 6546
rect 3228 6477 3234 6511
rect 3268 6477 3274 6511
rect 3228 6442 3274 6477
rect 3324 6511 3370 6546
rect 3324 6477 3330 6511
rect 3364 6477 3370 6511
rect 3324 6442 3370 6477
rect 3420 6511 3466 6546
rect 3420 6477 3426 6511
rect 3460 6477 3466 6511
rect 3420 6442 3466 6477
rect 3534 6519 3540 6553
rect 3574 6551 3580 6553
rect 3803 6551 3837 6679
rect 3574 6550 3680 6551
rect 3734 6550 3837 6551
rect 3574 6538 3687 6550
rect 3574 6519 3647 6538
rect 3534 6481 3647 6519
rect 3534 6447 3540 6481
rect 3574 6462 3647 6481
rect 3681 6462 3687 6538
rect 3574 6451 3687 6462
rect 3574 6447 3580 6451
rect 3641 6450 3687 6451
rect 3729 6538 3837 6550
rect 3987 6713 4021 6854
rect 4179 6713 4213 6854
rect 4371 6713 4405 6854
rect 4563 6713 4597 6854
rect 4755 6713 4789 6854
rect 4947 6713 4981 6854
rect 5055 6816 5101 6860
rect 5683 6767 5743 8020
rect 5177 6733 5743 6767
rect 5177 6713 5211 6733
rect 3987 6679 5211 6713
rect 3987 6546 4021 6679
rect 4179 6546 4213 6679
rect 4371 6546 4405 6679
rect 4563 6546 4597 6679
rect 4755 6546 4789 6679
rect 4947 6546 4981 6679
rect 5438 6675 5512 6676
rect 5326 6673 5400 6674
rect 5326 6621 5337 6673
rect 5389 6621 5400 6673
rect 5438 6623 5449 6675
rect 5501 6623 5512 6675
rect 5438 6622 5512 6623
rect 5326 6620 5400 6621
rect 5055 6553 5101 6576
rect 3729 6462 3735 6538
rect 3769 6462 3837 6538
rect 3729 6451 3837 6462
rect 3729 6450 3775 6451
rect 2450 6411 2516 6414
rect 2447 6359 2457 6411
rect 2509 6359 2519 6411
rect 2450 6354 2516 6359
rect 2562 6302 2596 6442
rect 2642 6411 2708 6414
rect 2638 6359 2648 6411
rect 2700 6359 2710 6411
rect 2642 6354 2708 6359
rect 2754 6302 2788 6442
rect 2834 6411 2900 6414
rect 2830 6359 2840 6411
rect 2892 6359 2902 6411
rect 2834 6354 2900 6359
rect 2946 6302 2980 6442
rect 3026 6411 3092 6414
rect 3022 6359 3032 6411
rect 3084 6359 3094 6411
rect 3026 6354 3092 6359
rect 3138 6302 3172 6442
rect 3218 6410 3284 6414
rect 3215 6358 3225 6410
rect 3277 6358 3287 6410
rect 3218 6354 3284 6358
rect 3330 6302 3364 6442
rect 3410 6410 3476 6414
rect 3407 6358 3417 6410
rect 3469 6358 3479 6410
rect 3534 6409 3580 6447
rect 3534 6375 3540 6409
rect 3574 6375 3580 6409
rect 3410 6354 3476 6358
rect 2282 6268 3364 6302
rect 3534 6192 3580 6375
rect 3803 6302 3837 6451
rect 3981 6511 4027 6546
rect 3981 6477 3987 6511
rect 4021 6477 4027 6511
rect 3981 6442 4027 6477
rect 4077 6511 4123 6546
rect 4077 6477 4083 6511
rect 4117 6477 4123 6511
rect 4077 6442 4123 6477
rect 4173 6511 4219 6546
rect 4173 6477 4179 6511
rect 4213 6477 4219 6511
rect 4173 6442 4219 6477
rect 4269 6511 4315 6546
rect 4269 6477 4275 6511
rect 4309 6477 4315 6511
rect 4269 6442 4315 6477
rect 4365 6511 4411 6546
rect 4365 6477 4371 6511
rect 4405 6477 4411 6511
rect 4365 6442 4411 6477
rect 4461 6511 4507 6546
rect 4461 6477 4467 6511
rect 4501 6477 4507 6511
rect 4461 6442 4507 6477
rect 4557 6511 4603 6546
rect 4557 6477 4563 6511
rect 4597 6477 4603 6511
rect 4557 6442 4603 6477
rect 4653 6511 4699 6546
rect 4653 6477 4659 6511
rect 4693 6477 4699 6511
rect 4653 6442 4699 6477
rect 4749 6511 4795 6546
rect 4749 6477 4755 6511
rect 4789 6477 4795 6511
rect 4749 6442 4795 6477
rect 4845 6511 4891 6546
rect 4845 6477 4851 6511
rect 4885 6477 4891 6511
rect 4845 6442 4891 6477
rect 4941 6511 4987 6546
rect 4941 6477 4947 6511
rect 4981 6477 4987 6511
rect 4941 6442 4987 6477
rect 5055 6519 5061 6553
rect 5095 6519 5101 6553
rect 5055 6481 5101 6519
rect 5055 6447 5061 6481
rect 5095 6464 5101 6481
rect 5095 6447 5550 6464
rect 3971 6411 4037 6414
rect 3968 6359 3978 6411
rect 4030 6359 4040 6411
rect 3971 6354 4037 6359
rect 4083 6302 4117 6442
rect 4163 6411 4229 6414
rect 4159 6359 4169 6411
rect 4221 6359 4231 6411
rect 4163 6354 4229 6359
rect 4275 6302 4309 6442
rect 4355 6411 4421 6414
rect 4351 6359 4361 6411
rect 4413 6359 4423 6411
rect 4355 6354 4421 6359
rect 4467 6302 4501 6442
rect 4547 6411 4613 6414
rect 4543 6359 4553 6411
rect 4605 6359 4615 6411
rect 4547 6354 4613 6359
rect 4659 6302 4693 6442
rect 4739 6410 4805 6414
rect 4736 6358 4746 6410
rect 4798 6358 4808 6410
rect 4739 6354 4805 6358
rect 4851 6302 4885 6442
rect 5055 6433 5550 6447
rect 4931 6410 4997 6414
rect 4928 6358 4938 6410
rect 4990 6358 5000 6410
rect 5055 6409 5303 6433
rect 5055 6375 5061 6409
rect 5095 6399 5303 6409
rect 5337 6399 5395 6433
rect 5429 6399 5487 6433
rect 5521 6399 5550 6433
rect 5095 6375 5550 6399
rect 5055 6368 5550 6375
rect 4931 6354 4997 6358
rect 3803 6268 4885 6302
rect 5055 6193 5101 6368
rect 129 5985 1211 6019
rect 129 5422 163 5985
rect 294 5875 304 5927
rect 356 5875 366 5927
rect 409 5835 443 5985
rect 487 5875 497 5927
rect 549 5875 559 5927
rect 601 5835 635 5985
rect 678 5875 688 5927
rect 740 5875 750 5927
rect 793 5835 827 5985
rect 870 5875 880 5927
rect 932 5875 942 5927
rect 985 5835 1019 5985
rect 1062 5875 1072 5927
rect 1124 5875 1134 5927
rect 1177 5835 1211 5985
rect 1254 5875 1264 5927
rect 1316 5875 1326 5927
rect 1381 5891 1427 6055
rect 2282 5989 3364 6023
rect 1381 5857 1387 5891
rect 1421 5857 1427 5891
rect 1512 5868 1522 5928
rect 1578 5868 1792 5928
rect 1852 5868 1862 5928
rect 307 5788 353 5835
rect 307 5754 313 5788
rect 347 5754 353 5788
rect 307 5716 353 5754
rect 307 5682 313 5716
rect 347 5682 353 5716
rect 307 5644 353 5682
rect 307 5610 313 5644
rect 347 5610 353 5644
rect 307 5563 353 5610
rect 403 5788 449 5835
rect 403 5754 409 5788
rect 443 5754 449 5788
rect 403 5716 449 5754
rect 403 5682 409 5716
rect 443 5682 449 5716
rect 403 5644 449 5682
rect 403 5610 409 5644
rect 443 5610 449 5644
rect 403 5563 449 5610
rect 499 5788 545 5835
rect 499 5754 505 5788
rect 539 5754 545 5788
rect 499 5716 545 5754
rect 499 5682 505 5716
rect 539 5682 545 5716
rect 499 5644 545 5682
rect 499 5610 505 5644
rect 539 5610 545 5644
rect 499 5563 545 5610
rect 595 5788 641 5835
rect 595 5754 601 5788
rect 635 5754 641 5788
rect 595 5716 641 5754
rect 595 5682 601 5716
rect 635 5682 641 5716
rect 595 5644 641 5682
rect 595 5610 601 5644
rect 635 5610 641 5644
rect 595 5563 641 5610
rect 691 5788 737 5835
rect 691 5754 697 5788
rect 731 5754 737 5788
rect 691 5716 737 5754
rect 691 5682 697 5716
rect 731 5682 737 5716
rect 691 5644 737 5682
rect 691 5610 697 5644
rect 731 5610 737 5644
rect 691 5563 737 5610
rect 787 5788 833 5835
rect 787 5754 793 5788
rect 827 5754 833 5788
rect 787 5716 833 5754
rect 787 5682 793 5716
rect 827 5682 833 5716
rect 787 5644 833 5682
rect 787 5610 793 5644
rect 827 5610 833 5644
rect 787 5563 833 5610
rect 883 5788 929 5835
rect 883 5754 889 5788
rect 923 5754 929 5788
rect 883 5716 929 5754
rect 883 5682 889 5716
rect 923 5682 929 5716
rect 883 5644 929 5682
rect 883 5610 889 5644
rect 923 5610 929 5644
rect 883 5563 929 5610
rect 979 5788 1025 5835
rect 979 5754 985 5788
rect 1019 5754 1025 5788
rect 979 5716 1025 5754
rect 979 5682 985 5716
rect 1019 5682 1025 5716
rect 979 5644 1025 5682
rect 979 5610 985 5644
rect 1019 5610 1025 5644
rect 979 5563 1025 5610
rect 1075 5788 1121 5835
rect 1075 5754 1081 5788
rect 1115 5754 1121 5788
rect 1075 5716 1121 5754
rect 1075 5682 1081 5716
rect 1115 5682 1121 5716
rect 1075 5644 1121 5682
rect 1075 5610 1081 5644
rect 1115 5610 1121 5644
rect 1075 5563 1121 5610
rect 1171 5788 1217 5835
rect 1171 5754 1177 5788
rect 1211 5754 1217 5788
rect 1171 5716 1217 5754
rect 1171 5682 1177 5716
rect 1211 5682 1217 5716
rect 1171 5644 1217 5682
rect 1171 5610 1177 5644
rect 1211 5610 1217 5644
rect 1171 5563 1217 5610
rect 1267 5788 1313 5835
rect 1267 5754 1273 5788
rect 1307 5754 1313 5788
rect 1267 5716 1313 5754
rect 1267 5682 1273 5716
rect 1307 5682 1313 5716
rect 1267 5644 1313 5682
rect 1267 5610 1273 5644
rect 1307 5610 1313 5644
rect 1267 5563 1313 5610
rect 1381 5819 1427 5857
rect 1381 5785 1387 5819
rect 1421 5785 1427 5819
rect 1381 5747 1427 5785
rect 1381 5713 1387 5747
rect 1421 5713 1427 5747
rect 1381 5675 1427 5713
rect 1381 5641 1387 5675
rect 1421 5641 1427 5675
rect 1381 5631 1427 5641
rect 1381 5629 2160 5631
rect 1381 5603 2056 5629
rect 1381 5578 1387 5603
rect 1380 5569 1387 5578
rect 1421 5569 2056 5603
rect 0 5388 163 5422
rect 129 5011 163 5388
rect 313 5422 347 5563
rect 505 5422 539 5563
rect 697 5422 731 5563
rect 889 5422 923 5563
rect 1081 5422 1115 5563
rect 1273 5422 1307 5563
rect 1380 5521 2056 5569
rect 2190 5521 2200 5629
rect 1380 5519 2160 5521
rect 2282 5426 2316 5989
rect 2447 5879 2457 5931
rect 2509 5879 2519 5931
rect 2562 5839 2596 5989
rect 2640 5879 2650 5931
rect 2702 5879 2712 5931
rect 2754 5839 2788 5989
rect 2831 5879 2841 5931
rect 2893 5879 2903 5931
rect 2946 5839 2980 5989
rect 3023 5879 3033 5931
rect 3085 5879 3095 5931
rect 3138 5839 3172 5989
rect 3215 5879 3225 5931
rect 3277 5879 3287 5931
rect 3330 5839 3364 5989
rect 3407 5879 3417 5931
rect 3469 5879 3479 5931
rect 3534 5895 3580 6103
rect 3534 5861 3540 5895
rect 3574 5861 3580 5895
rect 2460 5792 2506 5839
rect 2460 5758 2466 5792
rect 2500 5758 2506 5792
rect 2460 5720 2506 5758
rect 2460 5686 2466 5720
rect 2500 5686 2506 5720
rect 2460 5648 2506 5686
rect 2460 5614 2466 5648
rect 2500 5614 2506 5648
rect 2460 5567 2506 5614
rect 2556 5792 2602 5839
rect 2556 5758 2562 5792
rect 2596 5758 2602 5792
rect 2556 5720 2602 5758
rect 2556 5686 2562 5720
rect 2596 5686 2602 5720
rect 2556 5648 2602 5686
rect 2556 5614 2562 5648
rect 2596 5614 2602 5648
rect 2556 5567 2602 5614
rect 2652 5792 2698 5839
rect 2652 5758 2658 5792
rect 2692 5758 2698 5792
rect 2652 5720 2698 5758
rect 2652 5686 2658 5720
rect 2692 5686 2698 5720
rect 2652 5648 2698 5686
rect 2652 5614 2658 5648
rect 2692 5614 2698 5648
rect 2652 5567 2698 5614
rect 2748 5792 2794 5839
rect 2748 5758 2754 5792
rect 2788 5758 2794 5792
rect 2748 5720 2794 5758
rect 2748 5686 2754 5720
rect 2788 5686 2794 5720
rect 2748 5648 2794 5686
rect 2748 5614 2754 5648
rect 2788 5614 2794 5648
rect 2748 5567 2794 5614
rect 2844 5792 2890 5839
rect 2844 5758 2850 5792
rect 2884 5758 2890 5792
rect 2844 5720 2890 5758
rect 2844 5686 2850 5720
rect 2884 5686 2890 5720
rect 2844 5648 2890 5686
rect 2844 5614 2850 5648
rect 2884 5614 2890 5648
rect 2844 5567 2890 5614
rect 2940 5792 2986 5839
rect 2940 5758 2946 5792
rect 2980 5758 2986 5792
rect 2940 5720 2986 5758
rect 2940 5686 2946 5720
rect 2980 5686 2986 5720
rect 2940 5648 2986 5686
rect 2940 5614 2946 5648
rect 2980 5614 2986 5648
rect 2940 5567 2986 5614
rect 3036 5792 3082 5839
rect 3036 5758 3042 5792
rect 3076 5758 3082 5792
rect 3036 5720 3082 5758
rect 3036 5686 3042 5720
rect 3076 5686 3082 5720
rect 3036 5648 3082 5686
rect 3036 5614 3042 5648
rect 3076 5614 3082 5648
rect 3036 5567 3082 5614
rect 3132 5792 3178 5839
rect 3132 5758 3138 5792
rect 3172 5758 3178 5792
rect 3132 5720 3178 5758
rect 3132 5686 3138 5720
rect 3172 5686 3178 5720
rect 3132 5648 3178 5686
rect 3132 5614 3138 5648
rect 3172 5614 3178 5648
rect 3132 5567 3178 5614
rect 3228 5792 3274 5839
rect 3228 5758 3234 5792
rect 3268 5758 3274 5792
rect 3228 5720 3274 5758
rect 3228 5686 3234 5720
rect 3268 5686 3274 5720
rect 3228 5648 3274 5686
rect 3228 5614 3234 5648
rect 3268 5614 3274 5648
rect 3228 5567 3274 5614
rect 3324 5792 3370 5839
rect 3324 5758 3330 5792
rect 3364 5758 3370 5792
rect 3324 5720 3370 5758
rect 3324 5686 3330 5720
rect 3364 5686 3370 5720
rect 3324 5648 3370 5686
rect 3324 5614 3330 5648
rect 3364 5614 3370 5648
rect 3324 5567 3370 5614
rect 3420 5792 3466 5839
rect 3420 5758 3426 5792
rect 3460 5758 3466 5792
rect 3420 5720 3466 5758
rect 3420 5686 3426 5720
rect 3460 5686 3466 5720
rect 3420 5648 3466 5686
rect 3420 5614 3426 5648
rect 3460 5614 3466 5648
rect 3420 5567 3466 5614
rect 3534 5823 3580 5861
rect 3534 5789 3540 5823
rect 3574 5789 3580 5823
rect 3534 5751 3580 5789
rect 3534 5717 3540 5751
rect 3574 5717 3580 5751
rect 3534 5679 3580 5717
rect 3534 5645 3540 5679
rect 3574 5645 3580 5679
rect 3534 5607 3580 5645
rect 3534 5573 3540 5607
rect 3574 5573 3580 5607
rect 2101 5422 2316 5426
rect 313 5392 2316 5422
rect 313 5388 2141 5392
rect 313 5255 347 5388
rect 505 5255 539 5388
rect 697 5255 731 5388
rect 889 5255 923 5388
rect 1081 5255 1115 5388
rect 1273 5255 1307 5388
rect 1381 5262 1608 5285
rect 307 5220 353 5255
rect 307 5186 313 5220
rect 347 5186 353 5220
rect 307 5151 353 5186
rect 403 5220 449 5255
rect 403 5186 409 5220
rect 443 5186 449 5220
rect 403 5151 449 5186
rect 499 5220 545 5255
rect 499 5186 505 5220
rect 539 5186 545 5220
rect 499 5151 545 5186
rect 595 5220 641 5255
rect 595 5186 601 5220
rect 635 5186 641 5220
rect 595 5151 641 5186
rect 691 5220 737 5255
rect 691 5186 697 5220
rect 731 5186 737 5220
rect 691 5151 737 5186
rect 787 5220 833 5255
rect 787 5186 793 5220
rect 827 5186 833 5220
rect 787 5151 833 5186
rect 883 5220 929 5255
rect 883 5186 889 5220
rect 923 5186 929 5220
rect 883 5151 929 5186
rect 979 5220 1025 5255
rect 979 5186 985 5220
rect 1019 5186 1025 5220
rect 979 5151 1025 5186
rect 1075 5220 1121 5255
rect 1075 5186 1081 5220
rect 1115 5186 1121 5220
rect 1075 5151 1121 5186
rect 1171 5220 1217 5255
rect 1171 5186 1177 5220
rect 1211 5186 1217 5220
rect 1171 5151 1217 5186
rect 1267 5220 1313 5255
rect 1267 5186 1273 5220
rect 1307 5186 1313 5220
rect 1267 5151 1313 5186
rect 1381 5228 1387 5262
rect 1421 5228 1608 5262
rect 1381 5190 1608 5228
rect 1381 5156 1387 5190
rect 1421 5165 1608 5190
rect 1421 5156 1427 5165
rect 1560 5163 1608 5165
rect 1598 5161 1608 5163
rect 1720 5161 1730 5285
rect 297 5120 363 5123
rect 294 5068 304 5120
rect 356 5068 366 5120
rect 297 5063 363 5068
rect 409 5011 443 5151
rect 489 5120 555 5123
rect 485 5068 495 5120
rect 547 5068 557 5120
rect 489 5063 555 5068
rect 601 5011 635 5151
rect 681 5120 747 5123
rect 677 5068 687 5120
rect 739 5068 749 5120
rect 681 5063 747 5068
rect 793 5011 827 5151
rect 873 5120 939 5123
rect 869 5068 879 5120
rect 931 5068 941 5120
rect 873 5063 939 5068
rect 985 5011 1019 5151
rect 1065 5119 1131 5123
rect 1062 5067 1072 5119
rect 1124 5067 1134 5119
rect 1065 5063 1131 5067
rect 1177 5011 1211 5151
rect 1257 5119 1323 5123
rect 1254 5067 1264 5119
rect 1316 5067 1326 5119
rect 1381 5118 1427 5156
rect 1920 5123 1930 5125
rect 1381 5084 1387 5118
rect 1421 5084 1427 5118
rect 1257 5063 1323 5067
rect 129 4977 1211 5011
rect 1381 4941 1427 5084
rect 1458 5067 1468 5123
rect 1524 5069 1930 5123
rect 1986 5069 1996 5125
rect 1524 5067 1986 5069
rect 2282 5015 2316 5392
rect 2466 5426 2500 5567
rect 2658 5426 2692 5567
rect 2850 5426 2884 5567
rect 3042 5426 3076 5567
rect 3234 5426 3268 5567
rect 3426 5426 3460 5567
rect 3534 5529 3580 5573
rect 3803 5989 4885 6023
rect 3803 5426 3837 5989
rect 3968 5879 3978 5931
rect 4030 5879 4040 5931
rect 4083 5839 4117 5989
rect 4161 5879 4171 5931
rect 4223 5879 4233 5931
rect 4275 5839 4309 5989
rect 4352 5879 4362 5931
rect 4414 5879 4424 5931
rect 4467 5839 4501 5989
rect 4544 5879 4554 5931
rect 4606 5879 4616 5931
rect 4659 5839 4693 5989
rect 4736 5879 4746 5931
rect 4798 5879 4808 5931
rect 4851 5839 4885 5989
rect 4928 5879 4938 5931
rect 4990 5879 5000 5931
rect 5055 5895 5101 6100
rect 5055 5861 5061 5895
rect 5095 5861 5101 5895
rect 3981 5792 4027 5839
rect 3981 5758 3987 5792
rect 4021 5758 4027 5792
rect 3981 5720 4027 5758
rect 3981 5686 3987 5720
rect 4021 5686 4027 5720
rect 3981 5648 4027 5686
rect 3981 5614 3987 5648
rect 4021 5614 4027 5648
rect 3981 5567 4027 5614
rect 4077 5792 4123 5839
rect 4077 5758 4083 5792
rect 4117 5758 4123 5792
rect 4077 5720 4123 5758
rect 4077 5686 4083 5720
rect 4117 5686 4123 5720
rect 4077 5648 4123 5686
rect 4077 5614 4083 5648
rect 4117 5614 4123 5648
rect 4077 5567 4123 5614
rect 4173 5792 4219 5839
rect 4173 5758 4179 5792
rect 4213 5758 4219 5792
rect 4173 5720 4219 5758
rect 4173 5686 4179 5720
rect 4213 5686 4219 5720
rect 4173 5648 4219 5686
rect 4173 5614 4179 5648
rect 4213 5614 4219 5648
rect 4173 5567 4219 5614
rect 4269 5792 4315 5839
rect 4269 5758 4275 5792
rect 4309 5758 4315 5792
rect 4269 5720 4315 5758
rect 4269 5686 4275 5720
rect 4309 5686 4315 5720
rect 4269 5648 4315 5686
rect 4269 5614 4275 5648
rect 4309 5614 4315 5648
rect 4269 5567 4315 5614
rect 4365 5792 4411 5839
rect 4365 5758 4371 5792
rect 4405 5758 4411 5792
rect 4365 5720 4411 5758
rect 4365 5686 4371 5720
rect 4405 5686 4411 5720
rect 4365 5648 4411 5686
rect 4365 5614 4371 5648
rect 4405 5614 4411 5648
rect 4365 5567 4411 5614
rect 4461 5792 4507 5839
rect 4461 5758 4467 5792
rect 4501 5758 4507 5792
rect 4461 5720 4507 5758
rect 4461 5686 4467 5720
rect 4501 5686 4507 5720
rect 4461 5648 4507 5686
rect 4461 5614 4467 5648
rect 4501 5614 4507 5648
rect 4461 5567 4507 5614
rect 4557 5792 4603 5839
rect 4557 5758 4563 5792
rect 4597 5758 4603 5792
rect 4557 5720 4603 5758
rect 4557 5686 4563 5720
rect 4597 5686 4603 5720
rect 4557 5648 4603 5686
rect 4557 5614 4563 5648
rect 4597 5614 4603 5648
rect 4557 5567 4603 5614
rect 4653 5792 4699 5839
rect 4653 5758 4659 5792
rect 4693 5758 4699 5792
rect 4653 5720 4699 5758
rect 4653 5686 4659 5720
rect 4693 5686 4699 5720
rect 4653 5648 4699 5686
rect 4653 5614 4659 5648
rect 4693 5614 4699 5648
rect 4653 5567 4699 5614
rect 4749 5792 4795 5839
rect 4749 5758 4755 5792
rect 4789 5758 4795 5792
rect 4749 5720 4795 5758
rect 4749 5686 4755 5720
rect 4789 5686 4795 5720
rect 4749 5648 4795 5686
rect 4749 5614 4755 5648
rect 4789 5614 4795 5648
rect 4749 5567 4795 5614
rect 4845 5792 4891 5839
rect 4845 5758 4851 5792
rect 4885 5758 4891 5792
rect 4845 5720 4891 5758
rect 4845 5686 4851 5720
rect 4885 5686 4891 5720
rect 4845 5648 4891 5686
rect 4845 5614 4851 5648
rect 4885 5614 4891 5648
rect 4845 5567 4891 5614
rect 4941 5792 4987 5839
rect 4941 5758 4947 5792
rect 4981 5758 4987 5792
rect 4941 5720 4987 5758
rect 4941 5686 4947 5720
rect 4981 5686 4987 5720
rect 4941 5648 4987 5686
rect 4941 5614 4947 5648
rect 4981 5614 4987 5648
rect 4941 5567 4987 5614
rect 5055 5823 5101 5861
rect 5055 5789 5061 5823
rect 5095 5789 5101 5823
rect 5055 5751 5101 5789
rect 5055 5717 5061 5751
rect 5095 5720 5101 5751
rect 5274 5720 5550 5721
rect 5095 5717 5550 5720
rect 5055 5690 5550 5717
rect 5055 5679 5303 5690
rect 5055 5645 5061 5679
rect 5095 5656 5303 5679
rect 5337 5656 5395 5690
rect 5429 5656 5487 5690
rect 5521 5656 5550 5690
rect 5095 5645 5550 5656
rect 5055 5625 5550 5645
rect 5055 5607 5101 5625
rect 5055 5573 5061 5607
rect 5095 5573 5101 5607
rect 2466 5392 3837 5426
rect 2466 5259 2500 5392
rect 2658 5259 2692 5392
rect 2850 5259 2884 5392
rect 3042 5259 3076 5392
rect 3234 5259 3268 5392
rect 3426 5259 3460 5392
rect 3671 5302 3681 5354
rect 3733 5302 3743 5354
rect 3679 5301 3691 5302
rect 3725 5301 3737 5302
rect 3679 5295 3737 5301
rect 3534 5266 3580 5289
rect 2460 5224 2506 5259
rect 2460 5190 2466 5224
rect 2500 5190 2506 5224
rect 2460 5155 2506 5190
rect 2556 5224 2602 5259
rect 2556 5190 2562 5224
rect 2596 5190 2602 5224
rect 2556 5155 2602 5190
rect 2652 5224 2698 5259
rect 2652 5190 2658 5224
rect 2692 5190 2698 5224
rect 2652 5155 2698 5190
rect 2748 5224 2794 5259
rect 2748 5190 2754 5224
rect 2788 5190 2794 5224
rect 2748 5155 2794 5190
rect 2844 5224 2890 5259
rect 2844 5190 2850 5224
rect 2884 5190 2890 5224
rect 2844 5155 2890 5190
rect 2940 5224 2986 5259
rect 2940 5190 2946 5224
rect 2980 5190 2986 5224
rect 2940 5155 2986 5190
rect 3036 5224 3082 5259
rect 3036 5190 3042 5224
rect 3076 5190 3082 5224
rect 3036 5155 3082 5190
rect 3132 5224 3178 5259
rect 3132 5190 3138 5224
rect 3172 5190 3178 5224
rect 3132 5155 3178 5190
rect 3228 5224 3274 5259
rect 3228 5190 3234 5224
rect 3268 5190 3274 5224
rect 3228 5155 3274 5190
rect 3324 5224 3370 5259
rect 3324 5190 3330 5224
rect 3364 5190 3370 5224
rect 3324 5155 3370 5190
rect 3420 5224 3466 5259
rect 3420 5190 3426 5224
rect 3460 5190 3466 5224
rect 3420 5155 3466 5190
rect 3534 5232 3540 5266
rect 3574 5264 3580 5266
rect 3803 5264 3837 5392
rect 3574 5263 3680 5264
rect 3734 5263 3837 5264
rect 3574 5251 3687 5263
rect 3574 5232 3647 5251
rect 3534 5194 3647 5232
rect 3534 5160 3540 5194
rect 3574 5175 3647 5194
rect 3681 5175 3687 5251
rect 3574 5164 3687 5175
rect 3574 5160 3580 5164
rect 3641 5163 3687 5164
rect 3729 5251 3837 5263
rect 3987 5426 4021 5567
rect 4179 5426 4213 5567
rect 4371 5426 4405 5567
rect 4563 5426 4597 5567
rect 4755 5426 4789 5567
rect 4947 5426 4981 5567
rect 5055 5529 5101 5573
rect 5683 5480 5743 6733
rect 5177 5446 5743 5480
rect 5177 5426 5211 5446
rect 3987 5392 5211 5426
rect 3987 5259 4021 5392
rect 4179 5259 4213 5392
rect 4371 5259 4405 5392
rect 4563 5259 4597 5392
rect 4755 5259 4789 5392
rect 4947 5259 4981 5392
rect 5438 5388 5512 5389
rect 5326 5386 5400 5387
rect 5326 5334 5337 5386
rect 5389 5334 5400 5386
rect 5438 5336 5449 5388
rect 5501 5336 5512 5388
rect 5438 5335 5512 5336
rect 5326 5333 5400 5334
rect 5055 5266 5101 5289
rect 3729 5175 3735 5251
rect 3769 5175 3837 5251
rect 3729 5164 3837 5175
rect 3729 5163 3775 5164
rect 2450 5124 2516 5127
rect 2447 5072 2457 5124
rect 2509 5072 2519 5124
rect 2450 5067 2516 5072
rect 2562 5015 2596 5155
rect 2642 5124 2708 5127
rect 2638 5072 2648 5124
rect 2700 5072 2710 5124
rect 2642 5067 2708 5072
rect 2754 5015 2788 5155
rect 2834 5124 2900 5127
rect 2830 5072 2840 5124
rect 2892 5072 2902 5124
rect 2834 5067 2900 5072
rect 2946 5015 2980 5155
rect 3026 5124 3092 5127
rect 3022 5072 3032 5124
rect 3084 5072 3094 5124
rect 3026 5067 3092 5072
rect 3138 5015 3172 5155
rect 3218 5123 3284 5127
rect 3215 5071 3225 5123
rect 3277 5071 3287 5123
rect 3218 5067 3284 5071
rect 3330 5015 3364 5155
rect 3410 5123 3476 5127
rect 3407 5071 3417 5123
rect 3469 5071 3479 5123
rect 3534 5122 3580 5160
rect 3534 5088 3540 5122
rect 3574 5088 3580 5122
rect 3410 5067 3476 5071
rect 2282 4981 3364 5015
rect 3534 4905 3580 5088
rect 3803 5015 3837 5164
rect 3981 5224 4027 5259
rect 3981 5190 3987 5224
rect 4021 5190 4027 5224
rect 3981 5155 4027 5190
rect 4077 5224 4123 5259
rect 4077 5190 4083 5224
rect 4117 5190 4123 5224
rect 4077 5155 4123 5190
rect 4173 5224 4219 5259
rect 4173 5190 4179 5224
rect 4213 5190 4219 5224
rect 4173 5155 4219 5190
rect 4269 5224 4315 5259
rect 4269 5190 4275 5224
rect 4309 5190 4315 5224
rect 4269 5155 4315 5190
rect 4365 5224 4411 5259
rect 4365 5190 4371 5224
rect 4405 5190 4411 5224
rect 4365 5155 4411 5190
rect 4461 5224 4507 5259
rect 4461 5190 4467 5224
rect 4501 5190 4507 5224
rect 4461 5155 4507 5190
rect 4557 5224 4603 5259
rect 4557 5190 4563 5224
rect 4597 5190 4603 5224
rect 4557 5155 4603 5190
rect 4653 5224 4699 5259
rect 4653 5190 4659 5224
rect 4693 5190 4699 5224
rect 4653 5155 4699 5190
rect 4749 5224 4795 5259
rect 4749 5190 4755 5224
rect 4789 5190 4795 5224
rect 4749 5155 4795 5190
rect 4845 5224 4891 5259
rect 4845 5190 4851 5224
rect 4885 5190 4891 5224
rect 4845 5155 4891 5190
rect 4941 5224 4987 5259
rect 4941 5190 4947 5224
rect 4981 5190 4987 5224
rect 4941 5155 4987 5190
rect 5055 5232 5061 5266
rect 5095 5232 5101 5266
rect 5055 5194 5101 5232
rect 5055 5160 5061 5194
rect 5095 5177 5101 5194
rect 5095 5160 5550 5177
rect 3971 5124 4037 5127
rect 3968 5072 3978 5124
rect 4030 5072 4040 5124
rect 3971 5067 4037 5072
rect 4083 5015 4117 5155
rect 4163 5124 4229 5127
rect 4159 5072 4169 5124
rect 4221 5072 4231 5124
rect 4163 5067 4229 5072
rect 4275 5015 4309 5155
rect 4355 5124 4421 5127
rect 4351 5072 4361 5124
rect 4413 5072 4423 5124
rect 4355 5067 4421 5072
rect 4467 5015 4501 5155
rect 4547 5124 4613 5127
rect 4543 5072 4553 5124
rect 4605 5072 4615 5124
rect 4547 5067 4613 5072
rect 4659 5015 4693 5155
rect 4739 5123 4805 5127
rect 4736 5071 4746 5123
rect 4798 5071 4808 5123
rect 4739 5067 4805 5071
rect 4851 5015 4885 5155
rect 5055 5146 5550 5160
rect 4931 5123 4997 5127
rect 4928 5071 4938 5123
rect 4990 5071 5000 5123
rect 5055 5122 5303 5146
rect 5055 5088 5061 5122
rect 5095 5112 5303 5122
rect 5337 5112 5395 5146
rect 5429 5112 5487 5146
rect 5521 5112 5550 5146
rect 5095 5088 5550 5112
rect 5055 5081 5550 5088
rect 4931 5067 4997 5071
rect 3803 4981 4885 5015
rect 5055 4906 5101 5081
rect 129 4698 1211 4732
rect 129 4135 163 4698
rect 294 4588 304 4640
rect 356 4588 366 4640
rect 409 4548 443 4698
rect 487 4588 497 4640
rect 549 4588 559 4640
rect 601 4548 635 4698
rect 678 4588 688 4640
rect 740 4588 750 4640
rect 793 4548 827 4698
rect 870 4588 880 4640
rect 932 4588 942 4640
rect 985 4548 1019 4698
rect 1062 4588 1072 4640
rect 1124 4588 1134 4640
rect 1177 4548 1211 4698
rect 1254 4588 1264 4640
rect 1316 4588 1326 4640
rect 1381 4604 1427 4768
rect 2282 4702 3364 4736
rect 1381 4570 1387 4604
rect 1421 4570 1427 4604
rect 1512 4581 1522 4641
rect 1578 4581 1792 4641
rect 1852 4581 1862 4641
rect 307 4501 353 4548
rect 307 4467 313 4501
rect 347 4467 353 4501
rect 307 4429 353 4467
rect 307 4395 313 4429
rect 347 4395 353 4429
rect 307 4357 353 4395
rect 307 4323 313 4357
rect 347 4323 353 4357
rect 307 4276 353 4323
rect 403 4501 449 4548
rect 403 4467 409 4501
rect 443 4467 449 4501
rect 403 4429 449 4467
rect 403 4395 409 4429
rect 443 4395 449 4429
rect 403 4357 449 4395
rect 403 4323 409 4357
rect 443 4323 449 4357
rect 403 4276 449 4323
rect 499 4501 545 4548
rect 499 4467 505 4501
rect 539 4467 545 4501
rect 499 4429 545 4467
rect 499 4395 505 4429
rect 539 4395 545 4429
rect 499 4357 545 4395
rect 499 4323 505 4357
rect 539 4323 545 4357
rect 499 4276 545 4323
rect 595 4501 641 4548
rect 595 4467 601 4501
rect 635 4467 641 4501
rect 595 4429 641 4467
rect 595 4395 601 4429
rect 635 4395 641 4429
rect 595 4357 641 4395
rect 595 4323 601 4357
rect 635 4323 641 4357
rect 595 4276 641 4323
rect 691 4501 737 4548
rect 691 4467 697 4501
rect 731 4467 737 4501
rect 691 4429 737 4467
rect 691 4395 697 4429
rect 731 4395 737 4429
rect 691 4357 737 4395
rect 691 4323 697 4357
rect 731 4323 737 4357
rect 691 4276 737 4323
rect 787 4501 833 4548
rect 787 4467 793 4501
rect 827 4467 833 4501
rect 787 4429 833 4467
rect 787 4395 793 4429
rect 827 4395 833 4429
rect 787 4357 833 4395
rect 787 4323 793 4357
rect 827 4323 833 4357
rect 787 4276 833 4323
rect 883 4501 929 4548
rect 883 4467 889 4501
rect 923 4467 929 4501
rect 883 4429 929 4467
rect 883 4395 889 4429
rect 923 4395 929 4429
rect 883 4357 929 4395
rect 883 4323 889 4357
rect 923 4323 929 4357
rect 883 4276 929 4323
rect 979 4501 1025 4548
rect 979 4467 985 4501
rect 1019 4467 1025 4501
rect 979 4429 1025 4467
rect 979 4395 985 4429
rect 1019 4395 1025 4429
rect 979 4357 1025 4395
rect 979 4323 985 4357
rect 1019 4323 1025 4357
rect 979 4276 1025 4323
rect 1075 4501 1121 4548
rect 1075 4467 1081 4501
rect 1115 4467 1121 4501
rect 1075 4429 1121 4467
rect 1075 4395 1081 4429
rect 1115 4395 1121 4429
rect 1075 4357 1121 4395
rect 1075 4323 1081 4357
rect 1115 4323 1121 4357
rect 1075 4276 1121 4323
rect 1171 4501 1217 4548
rect 1171 4467 1177 4501
rect 1211 4467 1217 4501
rect 1171 4429 1217 4467
rect 1171 4395 1177 4429
rect 1211 4395 1217 4429
rect 1171 4357 1217 4395
rect 1171 4323 1177 4357
rect 1211 4323 1217 4357
rect 1171 4276 1217 4323
rect 1267 4501 1313 4548
rect 1267 4467 1273 4501
rect 1307 4467 1313 4501
rect 1267 4429 1313 4467
rect 1267 4395 1273 4429
rect 1307 4395 1313 4429
rect 1267 4357 1313 4395
rect 1267 4323 1273 4357
rect 1307 4323 1313 4357
rect 1267 4276 1313 4323
rect 1381 4532 1427 4570
rect 1381 4498 1387 4532
rect 1421 4498 1427 4532
rect 1381 4460 1427 4498
rect 1381 4426 1387 4460
rect 1421 4426 1427 4460
rect 1381 4388 1427 4426
rect 1381 4354 1387 4388
rect 1421 4354 1427 4388
rect 1381 4344 1427 4354
rect 1381 4342 2160 4344
rect 1381 4316 2056 4342
rect 1381 4291 1387 4316
rect 1380 4282 1387 4291
rect 1421 4282 2056 4316
rect 0 4101 163 4135
rect 129 3724 163 4101
rect 313 4135 347 4276
rect 505 4135 539 4276
rect 697 4135 731 4276
rect 889 4135 923 4276
rect 1081 4135 1115 4276
rect 1273 4135 1307 4276
rect 1380 4234 2056 4282
rect 2190 4234 2200 4342
rect 1380 4232 2160 4234
rect 2282 4139 2316 4702
rect 2447 4592 2457 4644
rect 2509 4592 2519 4644
rect 2562 4552 2596 4702
rect 2640 4592 2650 4644
rect 2702 4592 2712 4644
rect 2754 4552 2788 4702
rect 2831 4592 2841 4644
rect 2893 4592 2903 4644
rect 2946 4552 2980 4702
rect 3023 4592 3033 4644
rect 3085 4592 3095 4644
rect 3138 4552 3172 4702
rect 3215 4592 3225 4644
rect 3277 4592 3287 4644
rect 3330 4552 3364 4702
rect 3407 4592 3417 4644
rect 3469 4592 3479 4644
rect 3534 4608 3580 4816
rect 3534 4574 3540 4608
rect 3574 4574 3580 4608
rect 2460 4505 2506 4552
rect 2460 4471 2466 4505
rect 2500 4471 2506 4505
rect 2460 4433 2506 4471
rect 2460 4399 2466 4433
rect 2500 4399 2506 4433
rect 2460 4361 2506 4399
rect 2460 4327 2466 4361
rect 2500 4327 2506 4361
rect 2460 4280 2506 4327
rect 2556 4505 2602 4552
rect 2556 4471 2562 4505
rect 2596 4471 2602 4505
rect 2556 4433 2602 4471
rect 2556 4399 2562 4433
rect 2596 4399 2602 4433
rect 2556 4361 2602 4399
rect 2556 4327 2562 4361
rect 2596 4327 2602 4361
rect 2556 4280 2602 4327
rect 2652 4505 2698 4552
rect 2652 4471 2658 4505
rect 2692 4471 2698 4505
rect 2652 4433 2698 4471
rect 2652 4399 2658 4433
rect 2692 4399 2698 4433
rect 2652 4361 2698 4399
rect 2652 4327 2658 4361
rect 2692 4327 2698 4361
rect 2652 4280 2698 4327
rect 2748 4505 2794 4552
rect 2748 4471 2754 4505
rect 2788 4471 2794 4505
rect 2748 4433 2794 4471
rect 2748 4399 2754 4433
rect 2788 4399 2794 4433
rect 2748 4361 2794 4399
rect 2748 4327 2754 4361
rect 2788 4327 2794 4361
rect 2748 4280 2794 4327
rect 2844 4505 2890 4552
rect 2844 4471 2850 4505
rect 2884 4471 2890 4505
rect 2844 4433 2890 4471
rect 2844 4399 2850 4433
rect 2884 4399 2890 4433
rect 2844 4361 2890 4399
rect 2844 4327 2850 4361
rect 2884 4327 2890 4361
rect 2844 4280 2890 4327
rect 2940 4505 2986 4552
rect 2940 4471 2946 4505
rect 2980 4471 2986 4505
rect 2940 4433 2986 4471
rect 2940 4399 2946 4433
rect 2980 4399 2986 4433
rect 2940 4361 2986 4399
rect 2940 4327 2946 4361
rect 2980 4327 2986 4361
rect 2940 4280 2986 4327
rect 3036 4505 3082 4552
rect 3036 4471 3042 4505
rect 3076 4471 3082 4505
rect 3036 4433 3082 4471
rect 3036 4399 3042 4433
rect 3076 4399 3082 4433
rect 3036 4361 3082 4399
rect 3036 4327 3042 4361
rect 3076 4327 3082 4361
rect 3036 4280 3082 4327
rect 3132 4505 3178 4552
rect 3132 4471 3138 4505
rect 3172 4471 3178 4505
rect 3132 4433 3178 4471
rect 3132 4399 3138 4433
rect 3172 4399 3178 4433
rect 3132 4361 3178 4399
rect 3132 4327 3138 4361
rect 3172 4327 3178 4361
rect 3132 4280 3178 4327
rect 3228 4505 3274 4552
rect 3228 4471 3234 4505
rect 3268 4471 3274 4505
rect 3228 4433 3274 4471
rect 3228 4399 3234 4433
rect 3268 4399 3274 4433
rect 3228 4361 3274 4399
rect 3228 4327 3234 4361
rect 3268 4327 3274 4361
rect 3228 4280 3274 4327
rect 3324 4505 3370 4552
rect 3324 4471 3330 4505
rect 3364 4471 3370 4505
rect 3324 4433 3370 4471
rect 3324 4399 3330 4433
rect 3364 4399 3370 4433
rect 3324 4361 3370 4399
rect 3324 4327 3330 4361
rect 3364 4327 3370 4361
rect 3324 4280 3370 4327
rect 3420 4505 3466 4552
rect 3420 4471 3426 4505
rect 3460 4471 3466 4505
rect 3420 4433 3466 4471
rect 3420 4399 3426 4433
rect 3460 4399 3466 4433
rect 3420 4361 3466 4399
rect 3420 4327 3426 4361
rect 3460 4327 3466 4361
rect 3420 4280 3466 4327
rect 3534 4536 3580 4574
rect 3534 4502 3540 4536
rect 3574 4502 3580 4536
rect 3534 4464 3580 4502
rect 3534 4430 3540 4464
rect 3574 4430 3580 4464
rect 3534 4392 3580 4430
rect 3534 4358 3540 4392
rect 3574 4358 3580 4392
rect 3534 4320 3580 4358
rect 3534 4286 3540 4320
rect 3574 4286 3580 4320
rect 2101 4135 2316 4139
rect 313 4105 2316 4135
rect 313 4101 2141 4105
rect 313 3968 347 4101
rect 505 3968 539 4101
rect 697 3968 731 4101
rect 889 3968 923 4101
rect 1081 3968 1115 4101
rect 1273 3968 1307 4101
rect 1381 3975 1608 3998
rect 307 3933 353 3968
rect 307 3899 313 3933
rect 347 3899 353 3933
rect 307 3864 353 3899
rect 403 3933 449 3968
rect 403 3899 409 3933
rect 443 3899 449 3933
rect 403 3864 449 3899
rect 499 3933 545 3968
rect 499 3899 505 3933
rect 539 3899 545 3933
rect 499 3864 545 3899
rect 595 3933 641 3968
rect 595 3899 601 3933
rect 635 3899 641 3933
rect 595 3864 641 3899
rect 691 3933 737 3968
rect 691 3899 697 3933
rect 731 3899 737 3933
rect 691 3864 737 3899
rect 787 3933 833 3968
rect 787 3899 793 3933
rect 827 3899 833 3933
rect 787 3864 833 3899
rect 883 3933 929 3968
rect 883 3899 889 3933
rect 923 3899 929 3933
rect 883 3864 929 3899
rect 979 3933 1025 3968
rect 979 3899 985 3933
rect 1019 3899 1025 3933
rect 979 3864 1025 3899
rect 1075 3933 1121 3968
rect 1075 3899 1081 3933
rect 1115 3899 1121 3933
rect 1075 3864 1121 3899
rect 1171 3933 1217 3968
rect 1171 3899 1177 3933
rect 1211 3899 1217 3933
rect 1171 3864 1217 3899
rect 1267 3933 1313 3968
rect 1267 3899 1273 3933
rect 1307 3899 1313 3933
rect 1267 3864 1313 3899
rect 1381 3941 1387 3975
rect 1421 3941 1608 3975
rect 1381 3903 1608 3941
rect 1381 3869 1387 3903
rect 1421 3878 1608 3903
rect 1421 3869 1427 3878
rect 1560 3876 1608 3878
rect 1598 3874 1608 3876
rect 1720 3874 1730 3998
rect 297 3833 363 3836
rect 294 3781 304 3833
rect 356 3781 366 3833
rect 297 3776 363 3781
rect 409 3724 443 3864
rect 489 3833 555 3836
rect 485 3781 495 3833
rect 547 3781 557 3833
rect 489 3776 555 3781
rect 601 3724 635 3864
rect 681 3833 747 3836
rect 677 3781 687 3833
rect 739 3781 749 3833
rect 681 3776 747 3781
rect 793 3724 827 3864
rect 873 3833 939 3836
rect 869 3781 879 3833
rect 931 3781 941 3833
rect 873 3776 939 3781
rect 985 3724 1019 3864
rect 1065 3832 1131 3836
rect 1062 3780 1072 3832
rect 1124 3780 1134 3832
rect 1065 3776 1131 3780
rect 1177 3724 1211 3864
rect 1257 3832 1323 3836
rect 1254 3780 1264 3832
rect 1316 3780 1326 3832
rect 1381 3831 1427 3869
rect 1920 3836 1930 3838
rect 1381 3797 1387 3831
rect 1421 3797 1427 3831
rect 1257 3776 1323 3780
rect 129 3690 1211 3724
rect 1381 3654 1427 3797
rect 1458 3780 1468 3836
rect 1524 3782 1930 3836
rect 1986 3782 1996 3838
rect 1524 3780 1986 3782
rect 2282 3728 2316 4105
rect 2466 4139 2500 4280
rect 2658 4139 2692 4280
rect 2850 4139 2884 4280
rect 3042 4139 3076 4280
rect 3234 4139 3268 4280
rect 3426 4139 3460 4280
rect 3534 4242 3580 4286
rect 3803 4702 4885 4736
rect 3803 4139 3837 4702
rect 3968 4592 3978 4644
rect 4030 4592 4040 4644
rect 4083 4552 4117 4702
rect 4161 4592 4171 4644
rect 4223 4592 4233 4644
rect 4275 4552 4309 4702
rect 4352 4592 4362 4644
rect 4414 4592 4424 4644
rect 4467 4552 4501 4702
rect 4544 4592 4554 4644
rect 4606 4592 4616 4644
rect 4659 4552 4693 4702
rect 4736 4592 4746 4644
rect 4798 4592 4808 4644
rect 4851 4552 4885 4702
rect 4928 4592 4938 4644
rect 4990 4592 5000 4644
rect 5055 4608 5101 4813
rect 5055 4574 5061 4608
rect 5095 4574 5101 4608
rect 3981 4505 4027 4552
rect 3981 4471 3987 4505
rect 4021 4471 4027 4505
rect 3981 4433 4027 4471
rect 3981 4399 3987 4433
rect 4021 4399 4027 4433
rect 3981 4361 4027 4399
rect 3981 4327 3987 4361
rect 4021 4327 4027 4361
rect 3981 4280 4027 4327
rect 4077 4505 4123 4552
rect 4077 4471 4083 4505
rect 4117 4471 4123 4505
rect 4077 4433 4123 4471
rect 4077 4399 4083 4433
rect 4117 4399 4123 4433
rect 4077 4361 4123 4399
rect 4077 4327 4083 4361
rect 4117 4327 4123 4361
rect 4077 4280 4123 4327
rect 4173 4505 4219 4552
rect 4173 4471 4179 4505
rect 4213 4471 4219 4505
rect 4173 4433 4219 4471
rect 4173 4399 4179 4433
rect 4213 4399 4219 4433
rect 4173 4361 4219 4399
rect 4173 4327 4179 4361
rect 4213 4327 4219 4361
rect 4173 4280 4219 4327
rect 4269 4505 4315 4552
rect 4269 4471 4275 4505
rect 4309 4471 4315 4505
rect 4269 4433 4315 4471
rect 4269 4399 4275 4433
rect 4309 4399 4315 4433
rect 4269 4361 4315 4399
rect 4269 4327 4275 4361
rect 4309 4327 4315 4361
rect 4269 4280 4315 4327
rect 4365 4505 4411 4552
rect 4365 4471 4371 4505
rect 4405 4471 4411 4505
rect 4365 4433 4411 4471
rect 4365 4399 4371 4433
rect 4405 4399 4411 4433
rect 4365 4361 4411 4399
rect 4365 4327 4371 4361
rect 4405 4327 4411 4361
rect 4365 4280 4411 4327
rect 4461 4505 4507 4552
rect 4461 4471 4467 4505
rect 4501 4471 4507 4505
rect 4461 4433 4507 4471
rect 4461 4399 4467 4433
rect 4501 4399 4507 4433
rect 4461 4361 4507 4399
rect 4461 4327 4467 4361
rect 4501 4327 4507 4361
rect 4461 4280 4507 4327
rect 4557 4505 4603 4552
rect 4557 4471 4563 4505
rect 4597 4471 4603 4505
rect 4557 4433 4603 4471
rect 4557 4399 4563 4433
rect 4597 4399 4603 4433
rect 4557 4361 4603 4399
rect 4557 4327 4563 4361
rect 4597 4327 4603 4361
rect 4557 4280 4603 4327
rect 4653 4505 4699 4552
rect 4653 4471 4659 4505
rect 4693 4471 4699 4505
rect 4653 4433 4699 4471
rect 4653 4399 4659 4433
rect 4693 4399 4699 4433
rect 4653 4361 4699 4399
rect 4653 4327 4659 4361
rect 4693 4327 4699 4361
rect 4653 4280 4699 4327
rect 4749 4505 4795 4552
rect 4749 4471 4755 4505
rect 4789 4471 4795 4505
rect 4749 4433 4795 4471
rect 4749 4399 4755 4433
rect 4789 4399 4795 4433
rect 4749 4361 4795 4399
rect 4749 4327 4755 4361
rect 4789 4327 4795 4361
rect 4749 4280 4795 4327
rect 4845 4505 4891 4552
rect 4845 4471 4851 4505
rect 4885 4471 4891 4505
rect 4845 4433 4891 4471
rect 4845 4399 4851 4433
rect 4885 4399 4891 4433
rect 4845 4361 4891 4399
rect 4845 4327 4851 4361
rect 4885 4327 4891 4361
rect 4845 4280 4891 4327
rect 4941 4505 4987 4552
rect 4941 4471 4947 4505
rect 4981 4471 4987 4505
rect 4941 4433 4987 4471
rect 4941 4399 4947 4433
rect 4981 4399 4987 4433
rect 4941 4361 4987 4399
rect 4941 4327 4947 4361
rect 4981 4327 4987 4361
rect 4941 4280 4987 4327
rect 5055 4536 5101 4574
rect 5055 4502 5061 4536
rect 5095 4502 5101 4536
rect 5055 4464 5101 4502
rect 5055 4430 5061 4464
rect 5095 4433 5101 4464
rect 5274 4433 5550 4434
rect 5095 4430 5550 4433
rect 5055 4403 5550 4430
rect 5055 4392 5303 4403
rect 5055 4358 5061 4392
rect 5095 4369 5303 4392
rect 5337 4369 5395 4403
rect 5429 4369 5487 4403
rect 5521 4369 5550 4403
rect 5095 4358 5550 4369
rect 5055 4338 5550 4358
rect 5055 4320 5101 4338
rect 5055 4286 5061 4320
rect 5095 4286 5101 4320
rect 2466 4105 3837 4139
rect 2466 3972 2500 4105
rect 2658 3972 2692 4105
rect 2850 3972 2884 4105
rect 3042 3972 3076 4105
rect 3234 3972 3268 4105
rect 3426 3972 3460 4105
rect 3671 4015 3681 4067
rect 3733 4015 3743 4067
rect 3679 4014 3691 4015
rect 3725 4014 3737 4015
rect 3679 4008 3737 4014
rect 3534 3979 3580 4002
rect 2460 3937 2506 3972
rect 2460 3903 2466 3937
rect 2500 3903 2506 3937
rect 2460 3868 2506 3903
rect 2556 3937 2602 3972
rect 2556 3903 2562 3937
rect 2596 3903 2602 3937
rect 2556 3868 2602 3903
rect 2652 3937 2698 3972
rect 2652 3903 2658 3937
rect 2692 3903 2698 3937
rect 2652 3868 2698 3903
rect 2748 3937 2794 3972
rect 2748 3903 2754 3937
rect 2788 3903 2794 3937
rect 2748 3868 2794 3903
rect 2844 3937 2890 3972
rect 2844 3903 2850 3937
rect 2884 3903 2890 3937
rect 2844 3868 2890 3903
rect 2940 3937 2986 3972
rect 2940 3903 2946 3937
rect 2980 3903 2986 3937
rect 2940 3868 2986 3903
rect 3036 3937 3082 3972
rect 3036 3903 3042 3937
rect 3076 3903 3082 3937
rect 3036 3868 3082 3903
rect 3132 3937 3178 3972
rect 3132 3903 3138 3937
rect 3172 3903 3178 3937
rect 3132 3868 3178 3903
rect 3228 3937 3274 3972
rect 3228 3903 3234 3937
rect 3268 3903 3274 3937
rect 3228 3868 3274 3903
rect 3324 3937 3370 3972
rect 3324 3903 3330 3937
rect 3364 3903 3370 3937
rect 3324 3868 3370 3903
rect 3420 3937 3466 3972
rect 3420 3903 3426 3937
rect 3460 3903 3466 3937
rect 3420 3868 3466 3903
rect 3534 3945 3540 3979
rect 3574 3977 3580 3979
rect 3803 3977 3837 4105
rect 3574 3976 3680 3977
rect 3734 3976 3837 3977
rect 3574 3964 3687 3976
rect 3574 3945 3647 3964
rect 3534 3907 3647 3945
rect 3534 3873 3540 3907
rect 3574 3888 3647 3907
rect 3681 3888 3687 3964
rect 3574 3877 3687 3888
rect 3574 3873 3580 3877
rect 3641 3876 3687 3877
rect 3729 3964 3837 3976
rect 3987 4139 4021 4280
rect 4179 4139 4213 4280
rect 4371 4139 4405 4280
rect 4563 4139 4597 4280
rect 4755 4139 4789 4280
rect 4947 4139 4981 4280
rect 5055 4242 5101 4286
rect 5683 4193 5743 5446
rect 5177 4159 5743 4193
rect 5177 4139 5211 4159
rect 3987 4105 5211 4139
rect 3987 3972 4021 4105
rect 4179 3972 4213 4105
rect 4371 3972 4405 4105
rect 4563 3972 4597 4105
rect 4755 3972 4789 4105
rect 4947 3972 4981 4105
rect 5438 4101 5512 4102
rect 5326 4099 5400 4100
rect 5326 4047 5337 4099
rect 5389 4047 5400 4099
rect 5438 4049 5449 4101
rect 5501 4049 5512 4101
rect 5438 4048 5512 4049
rect 5326 4046 5400 4047
rect 5055 3979 5101 4002
rect 3729 3888 3735 3964
rect 3769 3888 3837 3964
rect 3729 3877 3837 3888
rect 3729 3876 3775 3877
rect 2450 3837 2516 3840
rect 2447 3785 2457 3837
rect 2509 3785 2519 3837
rect 2450 3780 2516 3785
rect 2562 3728 2596 3868
rect 2642 3837 2708 3840
rect 2638 3785 2648 3837
rect 2700 3785 2710 3837
rect 2642 3780 2708 3785
rect 2754 3728 2788 3868
rect 2834 3837 2900 3840
rect 2830 3785 2840 3837
rect 2892 3785 2902 3837
rect 2834 3780 2900 3785
rect 2946 3728 2980 3868
rect 3026 3837 3092 3840
rect 3022 3785 3032 3837
rect 3084 3785 3094 3837
rect 3026 3780 3092 3785
rect 3138 3728 3172 3868
rect 3218 3836 3284 3840
rect 3215 3784 3225 3836
rect 3277 3784 3287 3836
rect 3218 3780 3284 3784
rect 3330 3728 3364 3868
rect 3410 3836 3476 3840
rect 3407 3784 3417 3836
rect 3469 3784 3479 3836
rect 3534 3835 3580 3873
rect 3534 3801 3540 3835
rect 3574 3801 3580 3835
rect 3410 3780 3476 3784
rect 2282 3694 3364 3728
rect 3534 3618 3580 3801
rect 3803 3728 3837 3877
rect 3981 3937 4027 3972
rect 3981 3903 3987 3937
rect 4021 3903 4027 3937
rect 3981 3868 4027 3903
rect 4077 3937 4123 3972
rect 4077 3903 4083 3937
rect 4117 3903 4123 3937
rect 4077 3868 4123 3903
rect 4173 3937 4219 3972
rect 4173 3903 4179 3937
rect 4213 3903 4219 3937
rect 4173 3868 4219 3903
rect 4269 3937 4315 3972
rect 4269 3903 4275 3937
rect 4309 3903 4315 3937
rect 4269 3868 4315 3903
rect 4365 3937 4411 3972
rect 4365 3903 4371 3937
rect 4405 3903 4411 3937
rect 4365 3868 4411 3903
rect 4461 3937 4507 3972
rect 4461 3903 4467 3937
rect 4501 3903 4507 3937
rect 4461 3868 4507 3903
rect 4557 3937 4603 3972
rect 4557 3903 4563 3937
rect 4597 3903 4603 3937
rect 4557 3868 4603 3903
rect 4653 3937 4699 3972
rect 4653 3903 4659 3937
rect 4693 3903 4699 3937
rect 4653 3868 4699 3903
rect 4749 3937 4795 3972
rect 4749 3903 4755 3937
rect 4789 3903 4795 3937
rect 4749 3868 4795 3903
rect 4845 3937 4891 3972
rect 4845 3903 4851 3937
rect 4885 3903 4891 3937
rect 4845 3868 4891 3903
rect 4941 3937 4987 3972
rect 4941 3903 4947 3937
rect 4981 3903 4987 3937
rect 4941 3868 4987 3903
rect 5055 3945 5061 3979
rect 5095 3945 5101 3979
rect 5055 3907 5101 3945
rect 5055 3873 5061 3907
rect 5095 3890 5101 3907
rect 5095 3873 5550 3890
rect 3971 3837 4037 3840
rect 3968 3785 3978 3837
rect 4030 3785 4040 3837
rect 3971 3780 4037 3785
rect 4083 3728 4117 3868
rect 4163 3837 4229 3840
rect 4159 3785 4169 3837
rect 4221 3785 4231 3837
rect 4163 3780 4229 3785
rect 4275 3728 4309 3868
rect 4355 3837 4421 3840
rect 4351 3785 4361 3837
rect 4413 3785 4423 3837
rect 4355 3780 4421 3785
rect 4467 3728 4501 3868
rect 4547 3837 4613 3840
rect 4543 3785 4553 3837
rect 4605 3785 4615 3837
rect 4547 3780 4613 3785
rect 4659 3728 4693 3868
rect 4739 3836 4805 3840
rect 4736 3784 4746 3836
rect 4798 3784 4808 3836
rect 4739 3780 4805 3784
rect 4851 3728 4885 3868
rect 5055 3859 5550 3873
rect 4931 3836 4997 3840
rect 4928 3784 4938 3836
rect 4990 3784 5000 3836
rect 5055 3835 5303 3859
rect 5055 3801 5061 3835
rect 5095 3825 5303 3835
rect 5337 3825 5395 3859
rect 5429 3825 5487 3859
rect 5521 3825 5550 3859
rect 5095 3801 5550 3825
rect 5055 3794 5550 3801
rect 4931 3780 4997 3784
rect 3803 3694 4885 3728
rect 5055 3619 5101 3794
rect 129 3411 1211 3445
rect 129 2848 163 3411
rect 294 3301 304 3353
rect 356 3301 366 3353
rect 409 3261 443 3411
rect 487 3301 497 3353
rect 549 3301 559 3353
rect 601 3261 635 3411
rect 678 3301 688 3353
rect 740 3301 750 3353
rect 793 3261 827 3411
rect 870 3301 880 3353
rect 932 3301 942 3353
rect 985 3261 1019 3411
rect 1062 3301 1072 3353
rect 1124 3301 1134 3353
rect 1177 3261 1211 3411
rect 1254 3301 1264 3353
rect 1316 3301 1326 3353
rect 1381 3317 1427 3481
rect 2282 3415 3364 3449
rect 1381 3283 1387 3317
rect 1421 3283 1427 3317
rect 1512 3294 1522 3354
rect 1578 3294 1792 3354
rect 1852 3294 1862 3354
rect 307 3214 353 3261
rect 307 3180 313 3214
rect 347 3180 353 3214
rect 307 3142 353 3180
rect 307 3108 313 3142
rect 347 3108 353 3142
rect 307 3070 353 3108
rect 307 3036 313 3070
rect 347 3036 353 3070
rect 307 2989 353 3036
rect 403 3214 449 3261
rect 403 3180 409 3214
rect 443 3180 449 3214
rect 403 3142 449 3180
rect 403 3108 409 3142
rect 443 3108 449 3142
rect 403 3070 449 3108
rect 403 3036 409 3070
rect 443 3036 449 3070
rect 403 2989 449 3036
rect 499 3214 545 3261
rect 499 3180 505 3214
rect 539 3180 545 3214
rect 499 3142 545 3180
rect 499 3108 505 3142
rect 539 3108 545 3142
rect 499 3070 545 3108
rect 499 3036 505 3070
rect 539 3036 545 3070
rect 499 2989 545 3036
rect 595 3214 641 3261
rect 595 3180 601 3214
rect 635 3180 641 3214
rect 595 3142 641 3180
rect 595 3108 601 3142
rect 635 3108 641 3142
rect 595 3070 641 3108
rect 595 3036 601 3070
rect 635 3036 641 3070
rect 595 2989 641 3036
rect 691 3214 737 3261
rect 691 3180 697 3214
rect 731 3180 737 3214
rect 691 3142 737 3180
rect 691 3108 697 3142
rect 731 3108 737 3142
rect 691 3070 737 3108
rect 691 3036 697 3070
rect 731 3036 737 3070
rect 691 2989 737 3036
rect 787 3214 833 3261
rect 787 3180 793 3214
rect 827 3180 833 3214
rect 787 3142 833 3180
rect 787 3108 793 3142
rect 827 3108 833 3142
rect 787 3070 833 3108
rect 787 3036 793 3070
rect 827 3036 833 3070
rect 787 2989 833 3036
rect 883 3214 929 3261
rect 883 3180 889 3214
rect 923 3180 929 3214
rect 883 3142 929 3180
rect 883 3108 889 3142
rect 923 3108 929 3142
rect 883 3070 929 3108
rect 883 3036 889 3070
rect 923 3036 929 3070
rect 883 2989 929 3036
rect 979 3214 1025 3261
rect 979 3180 985 3214
rect 1019 3180 1025 3214
rect 979 3142 1025 3180
rect 979 3108 985 3142
rect 1019 3108 1025 3142
rect 979 3070 1025 3108
rect 979 3036 985 3070
rect 1019 3036 1025 3070
rect 979 2989 1025 3036
rect 1075 3214 1121 3261
rect 1075 3180 1081 3214
rect 1115 3180 1121 3214
rect 1075 3142 1121 3180
rect 1075 3108 1081 3142
rect 1115 3108 1121 3142
rect 1075 3070 1121 3108
rect 1075 3036 1081 3070
rect 1115 3036 1121 3070
rect 1075 2989 1121 3036
rect 1171 3214 1217 3261
rect 1171 3180 1177 3214
rect 1211 3180 1217 3214
rect 1171 3142 1217 3180
rect 1171 3108 1177 3142
rect 1211 3108 1217 3142
rect 1171 3070 1217 3108
rect 1171 3036 1177 3070
rect 1211 3036 1217 3070
rect 1171 2989 1217 3036
rect 1267 3214 1313 3261
rect 1267 3180 1273 3214
rect 1307 3180 1313 3214
rect 1267 3142 1313 3180
rect 1267 3108 1273 3142
rect 1307 3108 1313 3142
rect 1267 3070 1313 3108
rect 1267 3036 1273 3070
rect 1307 3036 1313 3070
rect 1267 2989 1313 3036
rect 1381 3245 1427 3283
rect 1381 3211 1387 3245
rect 1421 3211 1427 3245
rect 1381 3173 1427 3211
rect 1381 3139 1387 3173
rect 1421 3139 1427 3173
rect 1381 3101 1427 3139
rect 1381 3067 1387 3101
rect 1421 3067 1427 3101
rect 1381 3057 1427 3067
rect 1381 3055 2160 3057
rect 1381 3029 2056 3055
rect 1381 3004 1387 3029
rect 1380 2995 1387 3004
rect 1421 2995 2056 3029
rect 0 2814 163 2848
rect 129 2437 163 2814
rect 313 2848 347 2989
rect 505 2848 539 2989
rect 697 2848 731 2989
rect 889 2848 923 2989
rect 1081 2848 1115 2989
rect 1273 2848 1307 2989
rect 1380 2947 2056 2995
rect 2190 2947 2200 3055
rect 1380 2945 2160 2947
rect 2282 2852 2316 3415
rect 2447 3305 2457 3357
rect 2509 3305 2519 3357
rect 2562 3265 2596 3415
rect 2640 3305 2650 3357
rect 2702 3305 2712 3357
rect 2754 3265 2788 3415
rect 2831 3305 2841 3357
rect 2893 3305 2903 3357
rect 2946 3265 2980 3415
rect 3023 3305 3033 3357
rect 3085 3305 3095 3357
rect 3138 3265 3172 3415
rect 3215 3305 3225 3357
rect 3277 3305 3287 3357
rect 3330 3265 3364 3415
rect 3407 3305 3417 3357
rect 3469 3305 3479 3357
rect 3534 3321 3580 3529
rect 3534 3287 3540 3321
rect 3574 3287 3580 3321
rect 2460 3218 2506 3265
rect 2460 3184 2466 3218
rect 2500 3184 2506 3218
rect 2460 3146 2506 3184
rect 2460 3112 2466 3146
rect 2500 3112 2506 3146
rect 2460 3074 2506 3112
rect 2460 3040 2466 3074
rect 2500 3040 2506 3074
rect 2460 2993 2506 3040
rect 2556 3218 2602 3265
rect 2556 3184 2562 3218
rect 2596 3184 2602 3218
rect 2556 3146 2602 3184
rect 2556 3112 2562 3146
rect 2596 3112 2602 3146
rect 2556 3074 2602 3112
rect 2556 3040 2562 3074
rect 2596 3040 2602 3074
rect 2556 2993 2602 3040
rect 2652 3218 2698 3265
rect 2652 3184 2658 3218
rect 2692 3184 2698 3218
rect 2652 3146 2698 3184
rect 2652 3112 2658 3146
rect 2692 3112 2698 3146
rect 2652 3074 2698 3112
rect 2652 3040 2658 3074
rect 2692 3040 2698 3074
rect 2652 2993 2698 3040
rect 2748 3218 2794 3265
rect 2748 3184 2754 3218
rect 2788 3184 2794 3218
rect 2748 3146 2794 3184
rect 2748 3112 2754 3146
rect 2788 3112 2794 3146
rect 2748 3074 2794 3112
rect 2748 3040 2754 3074
rect 2788 3040 2794 3074
rect 2748 2993 2794 3040
rect 2844 3218 2890 3265
rect 2844 3184 2850 3218
rect 2884 3184 2890 3218
rect 2844 3146 2890 3184
rect 2844 3112 2850 3146
rect 2884 3112 2890 3146
rect 2844 3074 2890 3112
rect 2844 3040 2850 3074
rect 2884 3040 2890 3074
rect 2844 2993 2890 3040
rect 2940 3218 2986 3265
rect 2940 3184 2946 3218
rect 2980 3184 2986 3218
rect 2940 3146 2986 3184
rect 2940 3112 2946 3146
rect 2980 3112 2986 3146
rect 2940 3074 2986 3112
rect 2940 3040 2946 3074
rect 2980 3040 2986 3074
rect 2940 2993 2986 3040
rect 3036 3218 3082 3265
rect 3036 3184 3042 3218
rect 3076 3184 3082 3218
rect 3036 3146 3082 3184
rect 3036 3112 3042 3146
rect 3076 3112 3082 3146
rect 3036 3074 3082 3112
rect 3036 3040 3042 3074
rect 3076 3040 3082 3074
rect 3036 2993 3082 3040
rect 3132 3218 3178 3265
rect 3132 3184 3138 3218
rect 3172 3184 3178 3218
rect 3132 3146 3178 3184
rect 3132 3112 3138 3146
rect 3172 3112 3178 3146
rect 3132 3074 3178 3112
rect 3132 3040 3138 3074
rect 3172 3040 3178 3074
rect 3132 2993 3178 3040
rect 3228 3218 3274 3265
rect 3228 3184 3234 3218
rect 3268 3184 3274 3218
rect 3228 3146 3274 3184
rect 3228 3112 3234 3146
rect 3268 3112 3274 3146
rect 3228 3074 3274 3112
rect 3228 3040 3234 3074
rect 3268 3040 3274 3074
rect 3228 2993 3274 3040
rect 3324 3218 3370 3265
rect 3324 3184 3330 3218
rect 3364 3184 3370 3218
rect 3324 3146 3370 3184
rect 3324 3112 3330 3146
rect 3364 3112 3370 3146
rect 3324 3074 3370 3112
rect 3324 3040 3330 3074
rect 3364 3040 3370 3074
rect 3324 2993 3370 3040
rect 3420 3218 3466 3265
rect 3420 3184 3426 3218
rect 3460 3184 3466 3218
rect 3420 3146 3466 3184
rect 3420 3112 3426 3146
rect 3460 3112 3466 3146
rect 3420 3074 3466 3112
rect 3420 3040 3426 3074
rect 3460 3040 3466 3074
rect 3420 2993 3466 3040
rect 3534 3249 3580 3287
rect 3534 3215 3540 3249
rect 3574 3215 3580 3249
rect 3534 3177 3580 3215
rect 3534 3143 3540 3177
rect 3574 3143 3580 3177
rect 3534 3105 3580 3143
rect 3534 3071 3540 3105
rect 3574 3071 3580 3105
rect 3534 3033 3580 3071
rect 3534 2999 3540 3033
rect 3574 2999 3580 3033
rect 2101 2848 2316 2852
rect 313 2818 2316 2848
rect 313 2814 2141 2818
rect 313 2681 347 2814
rect 505 2681 539 2814
rect 697 2681 731 2814
rect 889 2681 923 2814
rect 1081 2681 1115 2814
rect 1273 2681 1307 2814
rect 1381 2688 1608 2711
rect 307 2646 353 2681
rect 307 2612 313 2646
rect 347 2612 353 2646
rect 307 2577 353 2612
rect 403 2646 449 2681
rect 403 2612 409 2646
rect 443 2612 449 2646
rect 403 2577 449 2612
rect 499 2646 545 2681
rect 499 2612 505 2646
rect 539 2612 545 2646
rect 499 2577 545 2612
rect 595 2646 641 2681
rect 595 2612 601 2646
rect 635 2612 641 2646
rect 595 2577 641 2612
rect 691 2646 737 2681
rect 691 2612 697 2646
rect 731 2612 737 2646
rect 691 2577 737 2612
rect 787 2646 833 2681
rect 787 2612 793 2646
rect 827 2612 833 2646
rect 787 2577 833 2612
rect 883 2646 929 2681
rect 883 2612 889 2646
rect 923 2612 929 2646
rect 883 2577 929 2612
rect 979 2646 1025 2681
rect 979 2612 985 2646
rect 1019 2612 1025 2646
rect 979 2577 1025 2612
rect 1075 2646 1121 2681
rect 1075 2612 1081 2646
rect 1115 2612 1121 2646
rect 1075 2577 1121 2612
rect 1171 2646 1217 2681
rect 1171 2612 1177 2646
rect 1211 2612 1217 2646
rect 1171 2577 1217 2612
rect 1267 2646 1313 2681
rect 1267 2612 1273 2646
rect 1307 2612 1313 2646
rect 1267 2577 1313 2612
rect 1381 2654 1387 2688
rect 1421 2654 1608 2688
rect 1381 2616 1608 2654
rect 1381 2582 1387 2616
rect 1421 2591 1608 2616
rect 1421 2582 1427 2591
rect 1560 2589 1608 2591
rect 1598 2587 1608 2589
rect 1720 2587 1730 2711
rect 297 2546 363 2549
rect 294 2494 304 2546
rect 356 2494 366 2546
rect 297 2489 363 2494
rect 409 2437 443 2577
rect 489 2546 555 2549
rect 485 2494 495 2546
rect 547 2494 557 2546
rect 489 2489 555 2494
rect 601 2437 635 2577
rect 681 2546 747 2549
rect 677 2494 687 2546
rect 739 2494 749 2546
rect 681 2489 747 2494
rect 793 2437 827 2577
rect 873 2546 939 2549
rect 869 2494 879 2546
rect 931 2494 941 2546
rect 873 2489 939 2494
rect 985 2437 1019 2577
rect 1065 2545 1131 2549
rect 1062 2493 1072 2545
rect 1124 2493 1134 2545
rect 1065 2489 1131 2493
rect 1177 2437 1211 2577
rect 1257 2545 1323 2549
rect 1254 2493 1264 2545
rect 1316 2493 1326 2545
rect 1381 2544 1427 2582
rect 1920 2549 1930 2551
rect 1381 2510 1387 2544
rect 1421 2510 1427 2544
rect 1257 2489 1323 2493
rect 129 2403 1211 2437
rect 1381 2367 1427 2510
rect 1458 2493 1468 2549
rect 1524 2495 1930 2549
rect 1986 2495 1996 2551
rect 1524 2493 1986 2495
rect 2282 2441 2316 2818
rect 2466 2852 2500 2993
rect 2658 2852 2692 2993
rect 2850 2852 2884 2993
rect 3042 2852 3076 2993
rect 3234 2852 3268 2993
rect 3426 2852 3460 2993
rect 3534 2955 3580 2999
rect 3803 3415 4885 3449
rect 3803 2852 3837 3415
rect 3968 3305 3978 3357
rect 4030 3305 4040 3357
rect 4083 3265 4117 3415
rect 4161 3305 4171 3357
rect 4223 3305 4233 3357
rect 4275 3265 4309 3415
rect 4352 3305 4362 3357
rect 4414 3305 4424 3357
rect 4467 3265 4501 3415
rect 4544 3305 4554 3357
rect 4606 3305 4616 3357
rect 4659 3265 4693 3415
rect 4736 3305 4746 3357
rect 4798 3305 4808 3357
rect 4851 3265 4885 3415
rect 4928 3305 4938 3357
rect 4990 3305 5000 3357
rect 5055 3321 5101 3526
rect 5055 3287 5061 3321
rect 5095 3287 5101 3321
rect 3981 3218 4027 3265
rect 3981 3184 3987 3218
rect 4021 3184 4027 3218
rect 3981 3146 4027 3184
rect 3981 3112 3987 3146
rect 4021 3112 4027 3146
rect 3981 3074 4027 3112
rect 3981 3040 3987 3074
rect 4021 3040 4027 3074
rect 3981 2993 4027 3040
rect 4077 3218 4123 3265
rect 4077 3184 4083 3218
rect 4117 3184 4123 3218
rect 4077 3146 4123 3184
rect 4077 3112 4083 3146
rect 4117 3112 4123 3146
rect 4077 3074 4123 3112
rect 4077 3040 4083 3074
rect 4117 3040 4123 3074
rect 4077 2993 4123 3040
rect 4173 3218 4219 3265
rect 4173 3184 4179 3218
rect 4213 3184 4219 3218
rect 4173 3146 4219 3184
rect 4173 3112 4179 3146
rect 4213 3112 4219 3146
rect 4173 3074 4219 3112
rect 4173 3040 4179 3074
rect 4213 3040 4219 3074
rect 4173 2993 4219 3040
rect 4269 3218 4315 3265
rect 4269 3184 4275 3218
rect 4309 3184 4315 3218
rect 4269 3146 4315 3184
rect 4269 3112 4275 3146
rect 4309 3112 4315 3146
rect 4269 3074 4315 3112
rect 4269 3040 4275 3074
rect 4309 3040 4315 3074
rect 4269 2993 4315 3040
rect 4365 3218 4411 3265
rect 4365 3184 4371 3218
rect 4405 3184 4411 3218
rect 4365 3146 4411 3184
rect 4365 3112 4371 3146
rect 4405 3112 4411 3146
rect 4365 3074 4411 3112
rect 4365 3040 4371 3074
rect 4405 3040 4411 3074
rect 4365 2993 4411 3040
rect 4461 3218 4507 3265
rect 4461 3184 4467 3218
rect 4501 3184 4507 3218
rect 4461 3146 4507 3184
rect 4461 3112 4467 3146
rect 4501 3112 4507 3146
rect 4461 3074 4507 3112
rect 4461 3040 4467 3074
rect 4501 3040 4507 3074
rect 4461 2993 4507 3040
rect 4557 3218 4603 3265
rect 4557 3184 4563 3218
rect 4597 3184 4603 3218
rect 4557 3146 4603 3184
rect 4557 3112 4563 3146
rect 4597 3112 4603 3146
rect 4557 3074 4603 3112
rect 4557 3040 4563 3074
rect 4597 3040 4603 3074
rect 4557 2993 4603 3040
rect 4653 3218 4699 3265
rect 4653 3184 4659 3218
rect 4693 3184 4699 3218
rect 4653 3146 4699 3184
rect 4653 3112 4659 3146
rect 4693 3112 4699 3146
rect 4653 3074 4699 3112
rect 4653 3040 4659 3074
rect 4693 3040 4699 3074
rect 4653 2993 4699 3040
rect 4749 3218 4795 3265
rect 4749 3184 4755 3218
rect 4789 3184 4795 3218
rect 4749 3146 4795 3184
rect 4749 3112 4755 3146
rect 4789 3112 4795 3146
rect 4749 3074 4795 3112
rect 4749 3040 4755 3074
rect 4789 3040 4795 3074
rect 4749 2993 4795 3040
rect 4845 3218 4891 3265
rect 4845 3184 4851 3218
rect 4885 3184 4891 3218
rect 4845 3146 4891 3184
rect 4845 3112 4851 3146
rect 4885 3112 4891 3146
rect 4845 3074 4891 3112
rect 4845 3040 4851 3074
rect 4885 3040 4891 3074
rect 4845 2993 4891 3040
rect 4941 3218 4987 3265
rect 4941 3184 4947 3218
rect 4981 3184 4987 3218
rect 4941 3146 4987 3184
rect 4941 3112 4947 3146
rect 4981 3112 4987 3146
rect 4941 3074 4987 3112
rect 4941 3040 4947 3074
rect 4981 3040 4987 3074
rect 4941 2993 4987 3040
rect 5055 3249 5101 3287
rect 5055 3215 5061 3249
rect 5095 3215 5101 3249
rect 5055 3177 5101 3215
rect 5055 3143 5061 3177
rect 5095 3146 5101 3177
rect 5274 3146 5550 3147
rect 5095 3143 5550 3146
rect 5055 3116 5550 3143
rect 5055 3105 5303 3116
rect 5055 3071 5061 3105
rect 5095 3082 5303 3105
rect 5337 3082 5395 3116
rect 5429 3082 5487 3116
rect 5521 3082 5550 3116
rect 5095 3071 5550 3082
rect 5055 3051 5550 3071
rect 5055 3033 5101 3051
rect 5055 2999 5061 3033
rect 5095 2999 5101 3033
rect 2466 2818 3837 2852
rect 2466 2685 2500 2818
rect 2658 2685 2692 2818
rect 2850 2685 2884 2818
rect 3042 2685 3076 2818
rect 3234 2685 3268 2818
rect 3426 2685 3460 2818
rect 3671 2728 3681 2780
rect 3733 2728 3743 2780
rect 3679 2727 3691 2728
rect 3725 2727 3737 2728
rect 3679 2721 3737 2727
rect 3534 2692 3580 2715
rect 2460 2650 2506 2685
rect 2460 2616 2466 2650
rect 2500 2616 2506 2650
rect 2460 2581 2506 2616
rect 2556 2650 2602 2685
rect 2556 2616 2562 2650
rect 2596 2616 2602 2650
rect 2556 2581 2602 2616
rect 2652 2650 2698 2685
rect 2652 2616 2658 2650
rect 2692 2616 2698 2650
rect 2652 2581 2698 2616
rect 2748 2650 2794 2685
rect 2748 2616 2754 2650
rect 2788 2616 2794 2650
rect 2748 2581 2794 2616
rect 2844 2650 2890 2685
rect 2844 2616 2850 2650
rect 2884 2616 2890 2650
rect 2844 2581 2890 2616
rect 2940 2650 2986 2685
rect 2940 2616 2946 2650
rect 2980 2616 2986 2650
rect 2940 2581 2986 2616
rect 3036 2650 3082 2685
rect 3036 2616 3042 2650
rect 3076 2616 3082 2650
rect 3036 2581 3082 2616
rect 3132 2650 3178 2685
rect 3132 2616 3138 2650
rect 3172 2616 3178 2650
rect 3132 2581 3178 2616
rect 3228 2650 3274 2685
rect 3228 2616 3234 2650
rect 3268 2616 3274 2650
rect 3228 2581 3274 2616
rect 3324 2650 3370 2685
rect 3324 2616 3330 2650
rect 3364 2616 3370 2650
rect 3324 2581 3370 2616
rect 3420 2650 3466 2685
rect 3420 2616 3426 2650
rect 3460 2616 3466 2650
rect 3420 2581 3466 2616
rect 3534 2658 3540 2692
rect 3574 2690 3580 2692
rect 3803 2690 3837 2818
rect 3574 2689 3680 2690
rect 3734 2689 3837 2690
rect 3574 2677 3687 2689
rect 3574 2658 3647 2677
rect 3534 2620 3647 2658
rect 3534 2586 3540 2620
rect 3574 2601 3647 2620
rect 3681 2601 3687 2677
rect 3574 2590 3687 2601
rect 3574 2586 3580 2590
rect 3641 2589 3687 2590
rect 3729 2677 3837 2689
rect 3987 2852 4021 2993
rect 4179 2852 4213 2993
rect 4371 2852 4405 2993
rect 4563 2852 4597 2993
rect 4755 2852 4789 2993
rect 4947 2852 4981 2993
rect 5055 2955 5101 2999
rect 5683 2906 5743 4159
rect 5177 2872 5743 2906
rect 5177 2852 5211 2872
rect 3987 2818 5211 2852
rect 3987 2685 4021 2818
rect 4179 2685 4213 2818
rect 4371 2685 4405 2818
rect 4563 2685 4597 2818
rect 4755 2685 4789 2818
rect 4947 2685 4981 2818
rect 5438 2814 5512 2815
rect 5326 2812 5400 2813
rect 5326 2760 5337 2812
rect 5389 2760 5400 2812
rect 5438 2762 5449 2814
rect 5501 2762 5512 2814
rect 5438 2761 5512 2762
rect 5326 2759 5400 2760
rect 5055 2692 5101 2715
rect 3729 2601 3735 2677
rect 3769 2601 3837 2677
rect 3729 2590 3837 2601
rect 3729 2589 3775 2590
rect 2450 2550 2516 2553
rect 2447 2498 2457 2550
rect 2509 2498 2519 2550
rect 2450 2493 2516 2498
rect 2562 2441 2596 2581
rect 2642 2550 2708 2553
rect 2638 2498 2648 2550
rect 2700 2498 2710 2550
rect 2642 2493 2708 2498
rect 2754 2441 2788 2581
rect 2834 2550 2900 2553
rect 2830 2498 2840 2550
rect 2892 2498 2902 2550
rect 2834 2493 2900 2498
rect 2946 2441 2980 2581
rect 3026 2550 3092 2553
rect 3022 2498 3032 2550
rect 3084 2498 3094 2550
rect 3026 2493 3092 2498
rect 3138 2441 3172 2581
rect 3218 2549 3284 2553
rect 3215 2497 3225 2549
rect 3277 2497 3287 2549
rect 3218 2493 3284 2497
rect 3330 2441 3364 2581
rect 3410 2549 3476 2553
rect 3407 2497 3417 2549
rect 3469 2497 3479 2549
rect 3534 2548 3580 2586
rect 3534 2514 3540 2548
rect 3574 2514 3580 2548
rect 3410 2493 3476 2497
rect 2282 2407 3364 2441
rect 3534 2331 3580 2514
rect 3803 2441 3837 2590
rect 3981 2650 4027 2685
rect 3981 2616 3987 2650
rect 4021 2616 4027 2650
rect 3981 2581 4027 2616
rect 4077 2650 4123 2685
rect 4077 2616 4083 2650
rect 4117 2616 4123 2650
rect 4077 2581 4123 2616
rect 4173 2650 4219 2685
rect 4173 2616 4179 2650
rect 4213 2616 4219 2650
rect 4173 2581 4219 2616
rect 4269 2650 4315 2685
rect 4269 2616 4275 2650
rect 4309 2616 4315 2650
rect 4269 2581 4315 2616
rect 4365 2650 4411 2685
rect 4365 2616 4371 2650
rect 4405 2616 4411 2650
rect 4365 2581 4411 2616
rect 4461 2650 4507 2685
rect 4461 2616 4467 2650
rect 4501 2616 4507 2650
rect 4461 2581 4507 2616
rect 4557 2650 4603 2685
rect 4557 2616 4563 2650
rect 4597 2616 4603 2650
rect 4557 2581 4603 2616
rect 4653 2650 4699 2685
rect 4653 2616 4659 2650
rect 4693 2616 4699 2650
rect 4653 2581 4699 2616
rect 4749 2650 4795 2685
rect 4749 2616 4755 2650
rect 4789 2616 4795 2650
rect 4749 2581 4795 2616
rect 4845 2650 4891 2685
rect 4845 2616 4851 2650
rect 4885 2616 4891 2650
rect 4845 2581 4891 2616
rect 4941 2650 4987 2685
rect 4941 2616 4947 2650
rect 4981 2616 4987 2650
rect 4941 2581 4987 2616
rect 5055 2658 5061 2692
rect 5095 2658 5101 2692
rect 5055 2620 5101 2658
rect 5055 2586 5061 2620
rect 5095 2603 5101 2620
rect 5095 2586 5550 2603
rect 3971 2550 4037 2553
rect 3968 2498 3978 2550
rect 4030 2498 4040 2550
rect 3971 2493 4037 2498
rect 4083 2441 4117 2581
rect 4163 2550 4229 2553
rect 4159 2498 4169 2550
rect 4221 2498 4231 2550
rect 4163 2493 4229 2498
rect 4275 2441 4309 2581
rect 4355 2550 4421 2553
rect 4351 2498 4361 2550
rect 4413 2498 4423 2550
rect 4355 2493 4421 2498
rect 4467 2441 4501 2581
rect 4547 2550 4613 2553
rect 4543 2498 4553 2550
rect 4605 2498 4615 2550
rect 4547 2493 4613 2498
rect 4659 2441 4693 2581
rect 4739 2549 4805 2553
rect 4736 2497 4746 2549
rect 4798 2497 4808 2549
rect 4739 2493 4805 2497
rect 4851 2441 4885 2581
rect 5055 2572 5550 2586
rect 4931 2549 4997 2553
rect 4928 2497 4938 2549
rect 4990 2497 5000 2549
rect 5055 2548 5303 2572
rect 5055 2514 5061 2548
rect 5095 2538 5303 2548
rect 5337 2538 5395 2572
rect 5429 2538 5487 2572
rect 5521 2538 5550 2572
rect 5095 2514 5550 2538
rect 5055 2507 5550 2514
rect 4931 2493 4997 2497
rect 3803 2407 4885 2441
rect 5055 2332 5101 2507
rect 129 2124 1211 2158
rect 129 1561 163 2124
rect 294 2014 304 2066
rect 356 2014 366 2066
rect 409 1974 443 2124
rect 487 2014 497 2066
rect 549 2014 559 2066
rect 601 1974 635 2124
rect 678 2014 688 2066
rect 740 2014 750 2066
rect 793 1974 827 2124
rect 870 2014 880 2066
rect 932 2014 942 2066
rect 985 1974 1019 2124
rect 1062 2014 1072 2066
rect 1124 2014 1134 2066
rect 1177 1974 1211 2124
rect 1254 2014 1264 2066
rect 1316 2014 1326 2066
rect 1381 2030 1427 2194
rect 2282 2128 3364 2162
rect 1381 1996 1387 2030
rect 1421 1996 1427 2030
rect 1512 2007 1522 2067
rect 1578 2007 1792 2067
rect 1852 2007 1862 2067
rect 307 1927 353 1974
rect 307 1893 313 1927
rect 347 1893 353 1927
rect 307 1855 353 1893
rect 307 1821 313 1855
rect 347 1821 353 1855
rect 307 1783 353 1821
rect 307 1749 313 1783
rect 347 1749 353 1783
rect 307 1702 353 1749
rect 403 1927 449 1974
rect 403 1893 409 1927
rect 443 1893 449 1927
rect 403 1855 449 1893
rect 403 1821 409 1855
rect 443 1821 449 1855
rect 403 1783 449 1821
rect 403 1749 409 1783
rect 443 1749 449 1783
rect 403 1702 449 1749
rect 499 1927 545 1974
rect 499 1893 505 1927
rect 539 1893 545 1927
rect 499 1855 545 1893
rect 499 1821 505 1855
rect 539 1821 545 1855
rect 499 1783 545 1821
rect 499 1749 505 1783
rect 539 1749 545 1783
rect 499 1702 545 1749
rect 595 1927 641 1974
rect 595 1893 601 1927
rect 635 1893 641 1927
rect 595 1855 641 1893
rect 595 1821 601 1855
rect 635 1821 641 1855
rect 595 1783 641 1821
rect 595 1749 601 1783
rect 635 1749 641 1783
rect 595 1702 641 1749
rect 691 1927 737 1974
rect 691 1893 697 1927
rect 731 1893 737 1927
rect 691 1855 737 1893
rect 691 1821 697 1855
rect 731 1821 737 1855
rect 691 1783 737 1821
rect 691 1749 697 1783
rect 731 1749 737 1783
rect 691 1702 737 1749
rect 787 1927 833 1974
rect 787 1893 793 1927
rect 827 1893 833 1927
rect 787 1855 833 1893
rect 787 1821 793 1855
rect 827 1821 833 1855
rect 787 1783 833 1821
rect 787 1749 793 1783
rect 827 1749 833 1783
rect 787 1702 833 1749
rect 883 1927 929 1974
rect 883 1893 889 1927
rect 923 1893 929 1927
rect 883 1855 929 1893
rect 883 1821 889 1855
rect 923 1821 929 1855
rect 883 1783 929 1821
rect 883 1749 889 1783
rect 923 1749 929 1783
rect 883 1702 929 1749
rect 979 1927 1025 1974
rect 979 1893 985 1927
rect 1019 1893 1025 1927
rect 979 1855 1025 1893
rect 979 1821 985 1855
rect 1019 1821 1025 1855
rect 979 1783 1025 1821
rect 979 1749 985 1783
rect 1019 1749 1025 1783
rect 979 1702 1025 1749
rect 1075 1927 1121 1974
rect 1075 1893 1081 1927
rect 1115 1893 1121 1927
rect 1075 1855 1121 1893
rect 1075 1821 1081 1855
rect 1115 1821 1121 1855
rect 1075 1783 1121 1821
rect 1075 1749 1081 1783
rect 1115 1749 1121 1783
rect 1075 1702 1121 1749
rect 1171 1927 1217 1974
rect 1171 1893 1177 1927
rect 1211 1893 1217 1927
rect 1171 1855 1217 1893
rect 1171 1821 1177 1855
rect 1211 1821 1217 1855
rect 1171 1783 1217 1821
rect 1171 1749 1177 1783
rect 1211 1749 1217 1783
rect 1171 1702 1217 1749
rect 1267 1927 1313 1974
rect 1267 1893 1273 1927
rect 1307 1893 1313 1927
rect 1267 1855 1313 1893
rect 1267 1821 1273 1855
rect 1307 1821 1313 1855
rect 1267 1783 1313 1821
rect 1267 1749 1273 1783
rect 1307 1749 1313 1783
rect 1267 1702 1313 1749
rect 1381 1958 1427 1996
rect 1381 1924 1387 1958
rect 1421 1924 1427 1958
rect 1381 1886 1427 1924
rect 1381 1852 1387 1886
rect 1421 1852 1427 1886
rect 1381 1814 1427 1852
rect 1381 1780 1387 1814
rect 1421 1780 1427 1814
rect 1381 1770 1427 1780
rect 1381 1768 2160 1770
rect 1381 1742 2056 1768
rect 1381 1717 1387 1742
rect 1380 1708 1387 1717
rect 1421 1708 2056 1742
rect 0 1527 163 1561
rect 129 1150 163 1527
rect 313 1561 347 1702
rect 505 1561 539 1702
rect 697 1561 731 1702
rect 889 1561 923 1702
rect 1081 1561 1115 1702
rect 1273 1561 1307 1702
rect 1380 1660 2056 1708
rect 2190 1660 2200 1768
rect 1380 1658 2160 1660
rect 2282 1565 2316 2128
rect 2447 2018 2457 2070
rect 2509 2018 2519 2070
rect 2562 1978 2596 2128
rect 2640 2018 2650 2070
rect 2702 2018 2712 2070
rect 2754 1978 2788 2128
rect 2831 2018 2841 2070
rect 2893 2018 2903 2070
rect 2946 1978 2980 2128
rect 3023 2018 3033 2070
rect 3085 2018 3095 2070
rect 3138 1978 3172 2128
rect 3215 2018 3225 2070
rect 3277 2018 3287 2070
rect 3330 1978 3364 2128
rect 3407 2018 3417 2070
rect 3469 2018 3479 2070
rect 3534 2034 3580 2242
rect 3534 2000 3540 2034
rect 3574 2000 3580 2034
rect 2460 1931 2506 1978
rect 2460 1897 2466 1931
rect 2500 1897 2506 1931
rect 2460 1859 2506 1897
rect 2460 1825 2466 1859
rect 2500 1825 2506 1859
rect 2460 1787 2506 1825
rect 2460 1753 2466 1787
rect 2500 1753 2506 1787
rect 2460 1706 2506 1753
rect 2556 1931 2602 1978
rect 2556 1897 2562 1931
rect 2596 1897 2602 1931
rect 2556 1859 2602 1897
rect 2556 1825 2562 1859
rect 2596 1825 2602 1859
rect 2556 1787 2602 1825
rect 2556 1753 2562 1787
rect 2596 1753 2602 1787
rect 2556 1706 2602 1753
rect 2652 1931 2698 1978
rect 2652 1897 2658 1931
rect 2692 1897 2698 1931
rect 2652 1859 2698 1897
rect 2652 1825 2658 1859
rect 2692 1825 2698 1859
rect 2652 1787 2698 1825
rect 2652 1753 2658 1787
rect 2692 1753 2698 1787
rect 2652 1706 2698 1753
rect 2748 1931 2794 1978
rect 2748 1897 2754 1931
rect 2788 1897 2794 1931
rect 2748 1859 2794 1897
rect 2748 1825 2754 1859
rect 2788 1825 2794 1859
rect 2748 1787 2794 1825
rect 2748 1753 2754 1787
rect 2788 1753 2794 1787
rect 2748 1706 2794 1753
rect 2844 1931 2890 1978
rect 2844 1897 2850 1931
rect 2884 1897 2890 1931
rect 2844 1859 2890 1897
rect 2844 1825 2850 1859
rect 2884 1825 2890 1859
rect 2844 1787 2890 1825
rect 2844 1753 2850 1787
rect 2884 1753 2890 1787
rect 2844 1706 2890 1753
rect 2940 1931 2986 1978
rect 2940 1897 2946 1931
rect 2980 1897 2986 1931
rect 2940 1859 2986 1897
rect 2940 1825 2946 1859
rect 2980 1825 2986 1859
rect 2940 1787 2986 1825
rect 2940 1753 2946 1787
rect 2980 1753 2986 1787
rect 2940 1706 2986 1753
rect 3036 1931 3082 1978
rect 3036 1897 3042 1931
rect 3076 1897 3082 1931
rect 3036 1859 3082 1897
rect 3036 1825 3042 1859
rect 3076 1825 3082 1859
rect 3036 1787 3082 1825
rect 3036 1753 3042 1787
rect 3076 1753 3082 1787
rect 3036 1706 3082 1753
rect 3132 1931 3178 1978
rect 3132 1897 3138 1931
rect 3172 1897 3178 1931
rect 3132 1859 3178 1897
rect 3132 1825 3138 1859
rect 3172 1825 3178 1859
rect 3132 1787 3178 1825
rect 3132 1753 3138 1787
rect 3172 1753 3178 1787
rect 3132 1706 3178 1753
rect 3228 1931 3274 1978
rect 3228 1897 3234 1931
rect 3268 1897 3274 1931
rect 3228 1859 3274 1897
rect 3228 1825 3234 1859
rect 3268 1825 3274 1859
rect 3228 1787 3274 1825
rect 3228 1753 3234 1787
rect 3268 1753 3274 1787
rect 3228 1706 3274 1753
rect 3324 1931 3370 1978
rect 3324 1897 3330 1931
rect 3364 1897 3370 1931
rect 3324 1859 3370 1897
rect 3324 1825 3330 1859
rect 3364 1825 3370 1859
rect 3324 1787 3370 1825
rect 3324 1753 3330 1787
rect 3364 1753 3370 1787
rect 3324 1706 3370 1753
rect 3420 1931 3466 1978
rect 3420 1897 3426 1931
rect 3460 1897 3466 1931
rect 3420 1859 3466 1897
rect 3420 1825 3426 1859
rect 3460 1825 3466 1859
rect 3420 1787 3466 1825
rect 3420 1753 3426 1787
rect 3460 1753 3466 1787
rect 3420 1706 3466 1753
rect 3534 1962 3580 2000
rect 3534 1928 3540 1962
rect 3574 1928 3580 1962
rect 3534 1890 3580 1928
rect 3534 1856 3540 1890
rect 3574 1856 3580 1890
rect 3534 1818 3580 1856
rect 3534 1784 3540 1818
rect 3574 1784 3580 1818
rect 3534 1746 3580 1784
rect 3534 1712 3540 1746
rect 3574 1712 3580 1746
rect 2101 1561 2316 1565
rect 313 1531 2316 1561
rect 313 1527 2141 1531
rect 313 1394 347 1527
rect 505 1394 539 1527
rect 697 1394 731 1527
rect 889 1394 923 1527
rect 1081 1394 1115 1527
rect 1273 1394 1307 1527
rect 1381 1401 1608 1424
rect 307 1359 353 1394
rect 307 1325 313 1359
rect 347 1325 353 1359
rect 307 1290 353 1325
rect 403 1359 449 1394
rect 403 1325 409 1359
rect 443 1325 449 1359
rect 403 1290 449 1325
rect 499 1359 545 1394
rect 499 1325 505 1359
rect 539 1325 545 1359
rect 499 1290 545 1325
rect 595 1359 641 1394
rect 595 1325 601 1359
rect 635 1325 641 1359
rect 595 1290 641 1325
rect 691 1359 737 1394
rect 691 1325 697 1359
rect 731 1325 737 1359
rect 691 1290 737 1325
rect 787 1359 833 1394
rect 787 1325 793 1359
rect 827 1325 833 1359
rect 787 1290 833 1325
rect 883 1359 929 1394
rect 883 1325 889 1359
rect 923 1325 929 1359
rect 883 1290 929 1325
rect 979 1359 1025 1394
rect 979 1325 985 1359
rect 1019 1325 1025 1359
rect 979 1290 1025 1325
rect 1075 1359 1121 1394
rect 1075 1325 1081 1359
rect 1115 1325 1121 1359
rect 1075 1290 1121 1325
rect 1171 1359 1217 1394
rect 1171 1325 1177 1359
rect 1211 1325 1217 1359
rect 1171 1290 1217 1325
rect 1267 1359 1313 1394
rect 1267 1325 1273 1359
rect 1307 1325 1313 1359
rect 1267 1290 1313 1325
rect 1381 1367 1387 1401
rect 1421 1367 1608 1401
rect 1381 1329 1608 1367
rect 1381 1295 1387 1329
rect 1421 1304 1608 1329
rect 1421 1295 1427 1304
rect 1560 1302 1608 1304
rect 1598 1300 1608 1302
rect 1720 1300 1730 1424
rect 297 1259 363 1262
rect 294 1207 304 1259
rect 356 1207 366 1259
rect 297 1202 363 1207
rect 409 1150 443 1290
rect 489 1259 555 1262
rect 485 1207 495 1259
rect 547 1207 557 1259
rect 489 1202 555 1207
rect 601 1150 635 1290
rect 681 1259 747 1262
rect 677 1207 687 1259
rect 739 1207 749 1259
rect 681 1202 747 1207
rect 793 1150 827 1290
rect 873 1259 939 1262
rect 869 1207 879 1259
rect 931 1207 941 1259
rect 873 1202 939 1207
rect 985 1150 1019 1290
rect 1065 1258 1131 1262
rect 1062 1206 1072 1258
rect 1124 1206 1134 1258
rect 1065 1202 1131 1206
rect 1177 1150 1211 1290
rect 1257 1258 1323 1262
rect 1254 1206 1264 1258
rect 1316 1206 1326 1258
rect 1381 1257 1427 1295
rect 1920 1262 1930 1264
rect 1381 1223 1387 1257
rect 1421 1223 1427 1257
rect 1257 1202 1323 1206
rect 129 1116 1211 1150
rect 1381 1080 1427 1223
rect 1458 1206 1468 1262
rect 1524 1208 1930 1262
rect 1986 1208 1996 1264
rect 1524 1206 1986 1208
rect 2282 1154 2316 1531
rect 2466 1565 2500 1706
rect 2658 1565 2692 1706
rect 2850 1565 2884 1706
rect 3042 1565 3076 1706
rect 3234 1565 3268 1706
rect 3426 1565 3460 1706
rect 3534 1668 3580 1712
rect 3803 2128 4885 2162
rect 3803 1565 3837 2128
rect 3968 2018 3978 2070
rect 4030 2018 4040 2070
rect 4083 1978 4117 2128
rect 4161 2018 4171 2070
rect 4223 2018 4233 2070
rect 4275 1978 4309 2128
rect 4352 2018 4362 2070
rect 4414 2018 4424 2070
rect 4467 1978 4501 2128
rect 4544 2018 4554 2070
rect 4606 2018 4616 2070
rect 4659 1978 4693 2128
rect 4736 2018 4746 2070
rect 4798 2018 4808 2070
rect 4851 1978 4885 2128
rect 4928 2018 4938 2070
rect 4990 2018 5000 2070
rect 5055 2034 5101 2239
rect 5055 2000 5061 2034
rect 5095 2000 5101 2034
rect 3981 1931 4027 1978
rect 3981 1897 3987 1931
rect 4021 1897 4027 1931
rect 3981 1859 4027 1897
rect 3981 1825 3987 1859
rect 4021 1825 4027 1859
rect 3981 1787 4027 1825
rect 3981 1753 3987 1787
rect 4021 1753 4027 1787
rect 3981 1706 4027 1753
rect 4077 1931 4123 1978
rect 4077 1897 4083 1931
rect 4117 1897 4123 1931
rect 4077 1859 4123 1897
rect 4077 1825 4083 1859
rect 4117 1825 4123 1859
rect 4077 1787 4123 1825
rect 4077 1753 4083 1787
rect 4117 1753 4123 1787
rect 4077 1706 4123 1753
rect 4173 1931 4219 1978
rect 4173 1897 4179 1931
rect 4213 1897 4219 1931
rect 4173 1859 4219 1897
rect 4173 1825 4179 1859
rect 4213 1825 4219 1859
rect 4173 1787 4219 1825
rect 4173 1753 4179 1787
rect 4213 1753 4219 1787
rect 4173 1706 4219 1753
rect 4269 1931 4315 1978
rect 4269 1897 4275 1931
rect 4309 1897 4315 1931
rect 4269 1859 4315 1897
rect 4269 1825 4275 1859
rect 4309 1825 4315 1859
rect 4269 1787 4315 1825
rect 4269 1753 4275 1787
rect 4309 1753 4315 1787
rect 4269 1706 4315 1753
rect 4365 1931 4411 1978
rect 4365 1897 4371 1931
rect 4405 1897 4411 1931
rect 4365 1859 4411 1897
rect 4365 1825 4371 1859
rect 4405 1825 4411 1859
rect 4365 1787 4411 1825
rect 4365 1753 4371 1787
rect 4405 1753 4411 1787
rect 4365 1706 4411 1753
rect 4461 1931 4507 1978
rect 4461 1897 4467 1931
rect 4501 1897 4507 1931
rect 4461 1859 4507 1897
rect 4461 1825 4467 1859
rect 4501 1825 4507 1859
rect 4461 1787 4507 1825
rect 4461 1753 4467 1787
rect 4501 1753 4507 1787
rect 4461 1706 4507 1753
rect 4557 1931 4603 1978
rect 4557 1897 4563 1931
rect 4597 1897 4603 1931
rect 4557 1859 4603 1897
rect 4557 1825 4563 1859
rect 4597 1825 4603 1859
rect 4557 1787 4603 1825
rect 4557 1753 4563 1787
rect 4597 1753 4603 1787
rect 4557 1706 4603 1753
rect 4653 1931 4699 1978
rect 4653 1897 4659 1931
rect 4693 1897 4699 1931
rect 4653 1859 4699 1897
rect 4653 1825 4659 1859
rect 4693 1825 4699 1859
rect 4653 1787 4699 1825
rect 4653 1753 4659 1787
rect 4693 1753 4699 1787
rect 4653 1706 4699 1753
rect 4749 1931 4795 1978
rect 4749 1897 4755 1931
rect 4789 1897 4795 1931
rect 4749 1859 4795 1897
rect 4749 1825 4755 1859
rect 4789 1825 4795 1859
rect 4749 1787 4795 1825
rect 4749 1753 4755 1787
rect 4789 1753 4795 1787
rect 4749 1706 4795 1753
rect 4845 1931 4891 1978
rect 4845 1897 4851 1931
rect 4885 1897 4891 1931
rect 4845 1859 4891 1897
rect 4845 1825 4851 1859
rect 4885 1825 4891 1859
rect 4845 1787 4891 1825
rect 4845 1753 4851 1787
rect 4885 1753 4891 1787
rect 4845 1706 4891 1753
rect 4941 1931 4987 1978
rect 4941 1897 4947 1931
rect 4981 1897 4987 1931
rect 4941 1859 4987 1897
rect 4941 1825 4947 1859
rect 4981 1825 4987 1859
rect 4941 1787 4987 1825
rect 4941 1753 4947 1787
rect 4981 1753 4987 1787
rect 4941 1706 4987 1753
rect 5055 1962 5101 2000
rect 5055 1928 5061 1962
rect 5095 1928 5101 1962
rect 5055 1890 5101 1928
rect 5055 1856 5061 1890
rect 5095 1859 5101 1890
rect 5274 1859 5550 1860
rect 5095 1856 5550 1859
rect 5055 1829 5550 1856
rect 5055 1818 5303 1829
rect 5055 1784 5061 1818
rect 5095 1795 5303 1818
rect 5337 1795 5395 1829
rect 5429 1795 5487 1829
rect 5521 1795 5550 1829
rect 5095 1784 5550 1795
rect 5055 1764 5550 1784
rect 5055 1746 5101 1764
rect 5055 1712 5061 1746
rect 5095 1712 5101 1746
rect 2466 1531 3837 1565
rect 2466 1398 2500 1531
rect 2658 1398 2692 1531
rect 2850 1398 2884 1531
rect 3042 1398 3076 1531
rect 3234 1398 3268 1531
rect 3426 1398 3460 1531
rect 3671 1441 3681 1493
rect 3733 1441 3743 1493
rect 3679 1440 3691 1441
rect 3725 1440 3737 1441
rect 3679 1434 3737 1440
rect 3534 1405 3580 1428
rect 2460 1363 2506 1398
rect 2460 1329 2466 1363
rect 2500 1329 2506 1363
rect 2460 1294 2506 1329
rect 2556 1363 2602 1398
rect 2556 1329 2562 1363
rect 2596 1329 2602 1363
rect 2556 1294 2602 1329
rect 2652 1363 2698 1398
rect 2652 1329 2658 1363
rect 2692 1329 2698 1363
rect 2652 1294 2698 1329
rect 2748 1363 2794 1398
rect 2748 1329 2754 1363
rect 2788 1329 2794 1363
rect 2748 1294 2794 1329
rect 2844 1363 2890 1398
rect 2844 1329 2850 1363
rect 2884 1329 2890 1363
rect 2844 1294 2890 1329
rect 2940 1363 2986 1398
rect 2940 1329 2946 1363
rect 2980 1329 2986 1363
rect 2940 1294 2986 1329
rect 3036 1363 3082 1398
rect 3036 1329 3042 1363
rect 3076 1329 3082 1363
rect 3036 1294 3082 1329
rect 3132 1363 3178 1398
rect 3132 1329 3138 1363
rect 3172 1329 3178 1363
rect 3132 1294 3178 1329
rect 3228 1363 3274 1398
rect 3228 1329 3234 1363
rect 3268 1329 3274 1363
rect 3228 1294 3274 1329
rect 3324 1363 3370 1398
rect 3324 1329 3330 1363
rect 3364 1329 3370 1363
rect 3324 1294 3370 1329
rect 3420 1363 3466 1398
rect 3420 1329 3426 1363
rect 3460 1329 3466 1363
rect 3420 1294 3466 1329
rect 3534 1371 3540 1405
rect 3574 1403 3580 1405
rect 3803 1403 3837 1531
rect 3574 1402 3680 1403
rect 3734 1402 3837 1403
rect 3574 1390 3687 1402
rect 3574 1371 3647 1390
rect 3534 1333 3647 1371
rect 3534 1299 3540 1333
rect 3574 1314 3647 1333
rect 3681 1314 3687 1390
rect 3574 1303 3687 1314
rect 3574 1299 3580 1303
rect 3641 1302 3687 1303
rect 3729 1390 3837 1402
rect 3987 1565 4021 1706
rect 4179 1565 4213 1706
rect 4371 1565 4405 1706
rect 4563 1565 4597 1706
rect 4755 1565 4789 1706
rect 4947 1565 4981 1706
rect 5055 1668 5101 1712
rect 5683 1619 5743 2872
rect 5177 1585 5743 1619
rect 5177 1565 5211 1585
rect 5683 1584 5743 1585
rect 3987 1531 5211 1565
rect 3987 1398 4021 1531
rect 4179 1398 4213 1531
rect 4371 1398 4405 1531
rect 4563 1398 4597 1531
rect 4755 1398 4789 1531
rect 4947 1398 4981 1531
rect 5438 1527 5512 1528
rect 5326 1525 5400 1526
rect 5326 1473 5337 1525
rect 5389 1473 5400 1525
rect 5438 1475 5449 1527
rect 5501 1475 5512 1527
rect 5438 1474 5512 1475
rect 5326 1472 5400 1473
rect 5055 1405 5101 1428
rect 3729 1314 3735 1390
rect 3769 1314 3837 1390
rect 3729 1303 3837 1314
rect 3729 1302 3775 1303
rect 2450 1263 2516 1266
rect 2447 1211 2457 1263
rect 2509 1211 2519 1263
rect 2450 1206 2516 1211
rect 2562 1154 2596 1294
rect 2642 1263 2708 1266
rect 2638 1211 2648 1263
rect 2700 1211 2710 1263
rect 2642 1206 2708 1211
rect 2754 1154 2788 1294
rect 2834 1263 2900 1266
rect 2830 1211 2840 1263
rect 2892 1211 2902 1263
rect 2834 1206 2900 1211
rect 2946 1154 2980 1294
rect 3026 1263 3092 1266
rect 3022 1211 3032 1263
rect 3084 1211 3094 1263
rect 3026 1206 3092 1211
rect 3138 1154 3172 1294
rect 3218 1262 3284 1266
rect 3215 1210 3225 1262
rect 3277 1210 3287 1262
rect 3218 1206 3284 1210
rect 3330 1154 3364 1294
rect 3410 1262 3476 1266
rect 3407 1210 3417 1262
rect 3469 1210 3479 1262
rect 3534 1261 3580 1299
rect 3534 1227 3540 1261
rect 3574 1227 3580 1261
rect 3410 1206 3476 1210
rect 2282 1120 3364 1154
rect 3534 1044 3580 1227
rect 3803 1154 3837 1303
rect 3981 1363 4027 1398
rect 3981 1329 3987 1363
rect 4021 1329 4027 1363
rect 3981 1294 4027 1329
rect 4077 1363 4123 1398
rect 4077 1329 4083 1363
rect 4117 1329 4123 1363
rect 4077 1294 4123 1329
rect 4173 1363 4219 1398
rect 4173 1329 4179 1363
rect 4213 1329 4219 1363
rect 4173 1294 4219 1329
rect 4269 1363 4315 1398
rect 4269 1329 4275 1363
rect 4309 1329 4315 1363
rect 4269 1294 4315 1329
rect 4365 1363 4411 1398
rect 4365 1329 4371 1363
rect 4405 1329 4411 1363
rect 4365 1294 4411 1329
rect 4461 1363 4507 1398
rect 4461 1329 4467 1363
rect 4501 1329 4507 1363
rect 4461 1294 4507 1329
rect 4557 1363 4603 1398
rect 4557 1329 4563 1363
rect 4597 1329 4603 1363
rect 4557 1294 4603 1329
rect 4653 1363 4699 1398
rect 4653 1329 4659 1363
rect 4693 1329 4699 1363
rect 4653 1294 4699 1329
rect 4749 1363 4795 1398
rect 4749 1329 4755 1363
rect 4789 1329 4795 1363
rect 4749 1294 4795 1329
rect 4845 1363 4891 1398
rect 4845 1329 4851 1363
rect 4885 1329 4891 1363
rect 4845 1294 4891 1329
rect 4941 1363 4987 1398
rect 4941 1329 4947 1363
rect 4981 1329 4987 1363
rect 4941 1294 4987 1329
rect 5055 1371 5061 1405
rect 5095 1371 5101 1405
rect 5055 1333 5101 1371
rect 5055 1299 5061 1333
rect 5095 1316 5101 1333
rect 5095 1299 5550 1316
rect 3971 1263 4037 1266
rect 3968 1211 3978 1263
rect 4030 1211 4040 1263
rect 3971 1206 4037 1211
rect 4083 1154 4117 1294
rect 4163 1263 4229 1266
rect 4159 1211 4169 1263
rect 4221 1211 4231 1263
rect 4163 1206 4229 1211
rect 4275 1154 4309 1294
rect 4355 1263 4421 1266
rect 4351 1211 4361 1263
rect 4413 1211 4423 1263
rect 4355 1206 4421 1211
rect 4467 1154 4501 1294
rect 4547 1263 4613 1266
rect 4543 1211 4553 1263
rect 4605 1211 4615 1263
rect 4547 1206 4613 1211
rect 4659 1154 4693 1294
rect 4739 1262 4805 1266
rect 4736 1210 4746 1262
rect 4798 1210 4808 1262
rect 4739 1206 4805 1210
rect 4851 1154 4885 1294
rect 5055 1285 5550 1299
rect 4931 1262 4997 1266
rect 4928 1210 4938 1262
rect 4990 1210 5000 1262
rect 5055 1261 5303 1285
rect 5055 1227 5061 1261
rect 5095 1251 5303 1261
rect 5337 1251 5395 1285
rect 5429 1251 5487 1285
rect 5521 1251 5550 1285
rect 5095 1227 5550 1251
rect 5055 1220 5550 1227
rect 4931 1206 4997 1210
rect 3803 1120 4885 1154
rect 5055 1045 5101 1220
<< via1 >>
rect 304 41953 356 41963
rect 304 41919 313 41953
rect 313 41919 347 41953
rect 347 41919 356 41953
rect 304 41911 356 41919
rect 497 41953 549 41963
rect 497 41919 505 41953
rect 505 41919 539 41953
rect 539 41919 549 41953
rect 497 41911 549 41919
rect 688 41953 740 41963
rect 688 41919 697 41953
rect 697 41919 731 41953
rect 731 41919 740 41953
rect 688 41911 740 41919
rect 880 41953 932 41963
rect 880 41919 889 41953
rect 889 41919 923 41953
rect 923 41919 932 41953
rect 880 41911 932 41919
rect 1072 41953 1124 41963
rect 1072 41919 1081 41953
rect 1081 41919 1115 41953
rect 1115 41919 1124 41953
rect 1072 41911 1124 41919
rect 1264 41953 1316 41963
rect 1264 41919 1273 41953
rect 1273 41919 1307 41953
rect 1307 41919 1316 41953
rect 1264 41911 1316 41919
rect 1522 41904 1578 41964
rect 1792 41904 1852 41964
rect 2056 41557 2190 41665
rect 2457 41957 2509 41967
rect 2457 41923 2466 41957
rect 2466 41923 2500 41957
rect 2500 41923 2509 41957
rect 2457 41915 2509 41923
rect 2650 41957 2702 41967
rect 2650 41923 2658 41957
rect 2658 41923 2692 41957
rect 2692 41923 2702 41957
rect 2650 41915 2702 41923
rect 2841 41957 2893 41967
rect 2841 41923 2850 41957
rect 2850 41923 2884 41957
rect 2884 41923 2893 41957
rect 2841 41915 2893 41923
rect 3033 41957 3085 41967
rect 3033 41923 3042 41957
rect 3042 41923 3076 41957
rect 3076 41923 3085 41957
rect 3033 41915 3085 41923
rect 3225 41957 3277 41967
rect 3225 41923 3234 41957
rect 3234 41923 3268 41957
rect 3268 41923 3277 41957
rect 3225 41915 3277 41923
rect 3417 41957 3469 41967
rect 3417 41923 3426 41957
rect 3426 41923 3460 41957
rect 3460 41923 3469 41957
rect 3417 41915 3469 41923
rect 1608 41197 1720 41321
rect 304 41145 356 41156
rect 304 41111 313 41145
rect 313 41111 347 41145
rect 347 41111 356 41145
rect 304 41104 356 41111
rect 495 41145 547 41156
rect 495 41111 505 41145
rect 505 41111 539 41145
rect 539 41111 547 41145
rect 495 41104 547 41111
rect 687 41145 739 41156
rect 687 41111 697 41145
rect 697 41111 731 41145
rect 731 41111 739 41145
rect 687 41104 739 41111
rect 879 41145 931 41156
rect 879 41111 889 41145
rect 889 41111 923 41145
rect 923 41111 931 41145
rect 879 41104 931 41111
rect 1072 41145 1124 41155
rect 1072 41111 1081 41145
rect 1081 41111 1115 41145
rect 1115 41111 1124 41145
rect 1072 41103 1124 41111
rect 1264 41145 1316 41155
rect 1264 41111 1273 41145
rect 1273 41111 1307 41145
rect 1307 41111 1316 41145
rect 1264 41103 1316 41111
rect 1468 41103 1524 41159
rect 1930 41105 1986 41161
rect 3978 41957 4030 41967
rect 3978 41923 3987 41957
rect 3987 41923 4021 41957
rect 4021 41923 4030 41957
rect 3978 41915 4030 41923
rect 4171 41957 4223 41967
rect 4171 41923 4179 41957
rect 4179 41923 4213 41957
rect 4213 41923 4223 41957
rect 4171 41915 4223 41923
rect 4362 41957 4414 41967
rect 4362 41923 4371 41957
rect 4371 41923 4405 41957
rect 4405 41923 4414 41957
rect 4362 41915 4414 41923
rect 4554 41957 4606 41967
rect 4554 41923 4563 41957
rect 4563 41923 4597 41957
rect 4597 41923 4606 41957
rect 4554 41915 4606 41923
rect 4746 41957 4798 41967
rect 4746 41923 4755 41957
rect 4755 41923 4789 41957
rect 4789 41923 4798 41957
rect 4746 41915 4798 41923
rect 4938 41957 4990 41967
rect 4938 41923 4947 41957
rect 4947 41923 4981 41957
rect 4981 41923 4990 41957
rect 4938 41915 4990 41923
rect 3681 41371 3733 41390
rect 3681 41338 3691 41371
rect 3691 41338 3725 41371
rect 3725 41338 3733 41371
rect 5337 41412 5389 41422
rect 5337 41378 5348 41412
rect 5348 41378 5382 41412
rect 5382 41378 5389 41412
rect 5337 41370 5389 41378
rect 5449 41417 5501 41424
rect 5449 41383 5450 41417
rect 5450 41383 5484 41417
rect 5484 41383 5501 41417
rect 5449 41372 5501 41383
rect 2457 41149 2509 41160
rect 2457 41115 2466 41149
rect 2466 41115 2500 41149
rect 2500 41115 2509 41149
rect 2457 41108 2509 41115
rect 2648 41149 2700 41160
rect 2648 41115 2658 41149
rect 2658 41115 2692 41149
rect 2692 41115 2700 41149
rect 2648 41108 2700 41115
rect 2840 41149 2892 41160
rect 2840 41115 2850 41149
rect 2850 41115 2884 41149
rect 2884 41115 2892 41149
rect 2840 41108 2892 41115
rect 3032 41149 3084 41160
rect 3032 41115 3042 41149
rect 3042 41115 3076 41149
rect 3076 41115 3084 41149
rect 3032 41108 3084 41115
rect 3225 41149 3277 41159
rect 3225 41115 3234 41149
rect 3234 41115 3268 41149
rect 3268 41115 3277 41149
rect 3225 41107 3277 41115
rect 3417 41149 3469 41159
rect 3417 41115 3426 41149
rect 3426 41115 3460 41149
rect 3460 41115 3469 41149
rect 3417 41107 3469 41115
rect 3978 41149 4030 41160
rect 3978 41115 3987 41149
rect 3987 41115 4021 41149
rect 4021 41115 4030 41149
rect 3978 41108 4030 41115
rect 4169 41149 4221 41160
rect 4169 41115 4179 41149
rect 4179 41115 4213 41149
rect 4213 41115 4221 41149
rect 4169 41108 4221 41115
rect 4361 41149 4413 41160
rect 4361 41115 4371 41149
rect 4371 41115 4405 41149
rect 4405 41115 4413 41149
rect 4361 41108 4413 41115
rect 4553 41149 4605 41160
rect 4553 41115 4563 41149
rect 4563 41115 4597 41149
rect 4597 41115 4605 41149
rect 4553 41108 4605 41115
rect 4746 41149 4798 41159
rect 4746 41115 4755 41149
rect 4755 41115 4789 41149
rect 4789 41115 4798 41149
rect 4746 41107 4798 41115
rect 4938 41149 4990 41159
rect 4938 41115 4947 41149
rect 4947 41115 4981 41149
rect 4981 41115 4990 41149
rect 4938 41107 4990 41115
rect 304 40666 356 40676
rect 304 40632 313 40666
rect 313 40632 347 40666
rect 347 40632 356 40666
rect 304 40624 356 40632
rect 497 40666 549 40676
rect 497 40632 505 40666
rect 505 40632 539 40666
rect 539 40632 549 40666
rect 497 40624 549 40632
rect 688 40666 740 40676
rect 688 40632 697 40666
rect 697 40632 731 40666
rect 731 40632 740 40666
rect 688 40624 740 40632
rect 880 40666 932 40676
rect 880 40632 889 40666
rect 889 40632 923 40666
rect 923 40632 932 40666
rect 880 40624 932 40632
rect 1072 40666 1124 40676
rect 1072 40632 1081 40666
rect 1081 40632 1115 40666
rect 1115 40632 1124 40666
rect 1072 40624 1124 40632
rect 1264 40666 1316 40676
rect 1264 40632 1273 40666
rect 1273 40632 1307 40666
rect 1307 40632 1316 40666
rect 1264 40624 1316 40632
rect 1522 40617 1578 40677
rect 1792 40617 1852 40677
rect 2056 40270 2190 40378
rect 2457 40670 2509 40680
rect 2457 40636 2466 40670
rect 2466 40636 2500 40670
rect 2500 40636 2509 40670
rect 2457 40628 2509 40636
rect 2650 40670 2702 40680
rect 2650 40636 2658 40670
rect 2658 40636 2692 40670
rect 2692 40636 2702 40670
rect 2650 40628 2702 40636
rect 2841 40670 2893 40680
rect 2841 40636 2850 40670
rect 2850 40636 2884 40670
rect 2884 40636 2893 40670
rect 2841 40628 2893 40636
rect 3033 40670 3085 40680
rect 3033 40636 3042 40670
rect 3042 40636 3076 40670
rect 3076 40636 3085 40670
rect 3033 40628 3085 40636
rect 3225 40670 3277 40680
rect 3225 40636 3234 40670
rect 3234 40636 3268 40670
rect 3268 40636 3277 40670
rect 3225 40628 3277 40636
rect 3417 40670 3469 40680
rect 3417 40636 3426 40670
rect 3426 40636 3460 40670
rect 3460 40636 3469 40670
rect 3417 40628 3469 40636
rect 1608 39910 1720 40034
rect 304 39858 356 39869
rect 304 39824 313 39858
rect 313 39824 347 39858
rect 347 39824 356 39858
rect 304 39817 356 39824
rect 495 39858 547 39869
rect 495 39824 505 39858
rect 505 39824 539 39858
rect 539 39824 547 39858
rect 495 39817 547 39824
rect 687 39858 739 39869
rect 687 39824 697 39858
rect 697 39824 731 39858
rect 731 39824 739 39858
rect 687 39817 739 39824
rect 879 39858 931 39869
rect 879 39824 889 39858
rect 889 39824 923 39858
rect 923 39824 931 39858
rect 879 39817 931 39824
rect 1072 39858 1124 39868
rect 1072 39824 1081 39858
rect 1081 39824 1115 39858
rect 1115 39824 1124 39858
rect 1072 39816 1124 39824
rect 1264 39858 1316 39868
rect 1264 39824 1273 39858
rect 1273 39824 1307 39858
rect 1307 39824 1316 39858
rect 1264 39816 1316 39824
rect 1468 39816 1524 39872
rect 1930 39818 1986 39874
rect 3978 40670 4030 40680
rect 3978 40636 3987 40670
rect 3987 40636 4021 40670
rect 4021 40636 4030 40670
rect 3978 40628 4030 40636
rect 4171 40670 4223 40680
rect 4171 40636 4179 40670
rect 4179 40636 4213 40670
rect 4213 40636 4223 40670
rect 4171 40628 4223 40636
rect 4362 40670 4414 40680
rect 4362 40636 4371 40670
rect 4371 40636 4405 40670
rect 4405 40636 4414 40670
rect 4362 40628 4414 40636
rect 4554 40670 4606 40680
rect 4554 40636 4563 40670
rect 4563 40636 4597 40670
rect 4597 40636 4606 40670
rect 4554 40628 4606 40636
rect 4746 40670 4798 40680
rect 4746 40636 4755 40670
rect 4755 40636 4789 40670
rect 4789 40636 4798 40670
rect 4746 40628 4798 40636
rect 4938 40670 4990 40680
rect 4938 40636 4947 40670
rect 4947 40636 4981 40670
rect 4981 40636 4990 40670
rect 4938 40628 4990 40636
rect 3681 40084 3733 40103
rect 3681 40051 3691 40084
rect 3691 40051 3725 40084
rect 3725 40051 3733 40084
rect 5337 40125 5389 40135
rect 5337 40091 5348 40125
rect 5348 40091 5382 40125
rect 5382 40091 5389 40125
rect 5337 40083 5389 40091
rect 5449 40130 5501 40137
rect 5449 40096 5450 40130
rect 5450 40096 5484 40130
rect 5484 40096 5501 40130
rect 5449 40085 5501 40096
rect 2457 39862 2509 39873
rect 2457 39828 2466 39862
rect 2466 39828 2500 39862
rect 2500 39828 2509 39862
rect 2457 39821 2509 39828
rect 2648 39862 2700 39873
rect 2648 39828 2658 39862
rect 2658 39828 2692 39862
rect 2692 39828 2700 39862
rect 2648 39821 2700 39828
rect 2840 39862 2892 39873
rect 2840 39828 2850 39862
rect 2850 39828 2884 39862
rect 2884 39828 2892 39862
rect 2840 39821 2892 39828
rect 3032 39862 3084 39873
rect 3032 39828 3042 39862
rect 3042 39828 3076 39862
rect 3076 39828 3084 39862
rect 3032 39821 3084 39828
rect 3225 39862 3277 39872
rect 3225 39828 3234 39862
rect 3234 39828 3268 39862
rect 3268 39828 3277 39862
rect 3225 39820 3277 39828
rect 3417 39862 3469 39872
rect 3417 39828 3426 39862
rect 3426 39828 3460 39862
rect 3460 39828 3469 39862
rect 3417 39820 3469 39828
rect 3978 39862 4030 39873
rect 3978 39828 3987 39862
rect 3987 39828 4021 39862
rect 4021 39828 4030 39862
rect 3978 39821 4030 39828
rect 4169 39862 4221 39873
rect 4169 39828 4179 39862
rect 4179 39828 4213 39862
rect 4213 39828 4221 39862
rect 4169 39821 4221 39828
rect 4361 39862 4413 39873
rect 4361 39828 4371 39862
rect 4371 39828 4405 39862
rect 4405 39828 4413 39862
rect 4361 39821 4413 39828
rect 4553 39862 4605 39873
rect 4553 39828 4563 39862
rect 4563 39828 4597 39862
rect 4597 39828 4605 39862
rect 4553 39821 4605 39828
rect 4746 39862 4798 39872
rect 4746 39828 4755 39862
rect 4755 39828 4789 39862
rect 4789 39828 4798 39862
rect 4746 39820 4798 39828
rect 4938 39862 4990 39872
rect 4938 39828 4947 39862
rect 4947 39828 4981 39862
rect 4981 39828 4990 39862
rect 4938 39820 4990 39828
rect 304 39379 356 39389
rect 304 39345 313 39379
rect 313 39345 347 39379
rect 347 39345 356 39379
rect 304 39337 356 39345
rect 497 39379 549 39389
rect 497 39345 505 39379
rect 505 39345 539 39379
rect 539 39345 549 39379
rect 497 39337 549 39345
rect 688 39379 740 39389
rect 688 39345 697 39379
rect 697 39345 731 39379
rect 731 39345 740 39379
rect 688 39337 740 39345
rect 880 39379 932 39389
rect 880 39345 889 39379
rect 889 39345 923 39379
rect 923 39345 932 39379
rect 880 39337 932 39345
rect 1072 39379 1124 39389
rect 1072 39345 1081 39379
rect 1081 39345 1115 39379
rect 1115 39345 1124 39379
rect 1072 39337 1124 39345
rect 1264 39379 1316 39389
rect 1264 39345 1273 39379
rect 1273 39345 1307 39379
rect 1307 39345 1316 39379
rect 1264 39337 1316 39345
rect 1522 39330 1578 39390
rect 1792 39330 1852 39390
rect 2056 38983 2190 39091
rect 2457 39383 2509 39393
rect 2457 39349 2466 39383
rect 2466 39349 2500 39383
rect 2500 39349 2509 39383
rect 2457 39341 2509 39349
rect 2650 39383 2702 39393
rect 2650 39349 2658 39383
rect 2658 39349 2692 39383
rect 2692 39349 2702 39383
rect 2650 39341 2702 39349
rect 2841 39383 2893 39393
rect 2841 39349 2850 39383
rect 2850 39349 2884 39383
rect 2884 39349 2893 39383
rect 2841 39341 2893 39349
rect 3033 39383 3085 39393
rect 3033 39349 3042 39383
rect 3042 39349 3076 39383
rect 3076 39349 3085 39383
rect 3033 39341 3085 39349
rect 3225 39383 3277 39393
rect 3225 39349 3234 39383
rect 3234 39349 3268 39383
rect 3268 39349 3277 39383
rect 3225 39341 3277 39349
rect 3417 39383 3469 39393
rect 3417 39349 3426 39383
rect 3426 39349 3460 39383
rect 3460 39349 3469 39383
rect 3417 39341 3469 39349
rect 1608 38623 1720 38747
rect 304 38571 356 38582
rect 304 38537 313 38571
rect 313 38537 347 38571
rect 347 38537 356 38571
rect 304 38530 356 38537
rect 495 38571 547 38582
rect 495 38537 505 38571
rect 505 38537 539 38571
rect 539 38537 547 38571
rect 495 38530 547 38537
rect 687 38571 739 38582
rect 687 38537 697 38571
rect 697 38537 731 38571
rect 731 38537 739 38571
rect 687 38530 739 38537
rect 879 38571 931 38582
rect 879 38537 889 38571
rect 889 38537 923 38571
rect 923 38537 931 38571
rect 879 38530 931 38537
rect 1072 38571 1124 38581
rect 1072 38537 1081 38571
rect 1081 38537 1115 38571
rect 1115 38537 1124 38571
rect 1072 38529 1124 38537
rect 1264 38571 1316 38581
rect 1264 38537 1273 38571
rect 1273 38537 1307 38571
rect 1307 38537 1316 38571
rect 1264 38529 1316 38537
rect 1468 38529 1524 38585
rect 1930 38531 1986 38587
rect 3978 39383 4030 39393
rect 3978 39349 3987 39383
rect 3987 39349 4021 39383
rect 4021 39349 4030 39383
rect 3978 39341 4030 39349
rect 4171 39383 4223 39393
rect 4171 39349 4179 39383
rect 4179 39349 4213 39383
rect 4213 39349 4223 39383
rect 4171 39341 4223 39349
rect 4362 39383 4414 39393
rect 4362 39349 4371 39383
rect 4371 39349 4405 39383
rect 4405 39349 4414 39383
rect 4362 39341 4414 39349
rect 4554 39383 4606 39393
rect 4554 39349 4563 39383
rect 4563 39349 4597 39383
rect 4597 39349 4606 39383
rect 4554 39341 4606 39349
rect 4746 39383 4798 39393
rect 4746 39349 4755 39383
rect 4755 39349 4789 39383
rect 4789 39349 4798 39383
rect 4746 39341 4798 39349
rect 4938 39383 4990 39393
rect 4938 39349 4947 39383
rect 4947 39349 4981 39383
rect 4981 39349 4990 39383
rect 4938 39341 4990 39349
rect 3681 38797 3733 38816
rect 3681 38764 3691 38797
rect 3691 38764 3725 38797
rect 3725 38764 3733 38797
rect 5337 38838 5389 38848
rect 5337 38804 5348 38838
rect 5348 38804 5382 38838
rect 5382 38804 5389 38838
rect 5337 38796 5389 38804
rect 5449 38843 5501 38850
rect 5449 38809 5450 38843
rect 5450 38809 5484 38843
rect 5484 38809 5501 38843
rect 5449 38798 5501 38809
rect 2457 38575 2509 38586
rect 2457 38541 2466 38575
rect 2466 38541 2500 38575
rect 2500 38541 2509 38575
rect 2457 38534 2509 38541
rect 2648 38575 2700 38586
rect 2648 38541 2658 38575
rect 2658 38541 2692 38575
rect 2692 38541 2700 38575
rect 2648 38534 2700 38541
rect 2840 38575 2892 38586
rect 2840 38541 2850 38575
rect 2850 38541 2884 38575
rect 2884 38541 2892 38575
rect 2840 38534 2892 38541
rect 3032 38575 3084 38586
rect 3032 38541 3042 38575
rect 3042 38541 3076 38575
rect 3076 38541 3084 38575
rect 3032 38534 3084 38541
rect 3225 38575 3277 38585
rect 3225 38541 3234 38575
rect 3234 38541 3268 38575
rect 3268 38541 3277 38575
rect 3225 38533 3277 38541
rect 3417 38575 3469 38585
rect 3417 38541 3426 38575
rect 3426 38541 3460 38575
rect 3460 38541 3469 38575
rect 3417 38533 3469 38541
rect 3978 38575 4030 38586
rect 3978 38541 3987 38575
rect 3987 38541 4021 38575
rect 4021 38541 4030 38575
rect 3978 38534 4030 38541
rect 4169 38575 4221 38586
rect 4169 38541 4179 38575
rect 4179 38541 4213 38575
rect 4213 38541 4221 38575
rect 4169 38534 4221 38541
rect 4361 38575 4413 38586
rect 4361 38541 4371 38575
rect 4371 38541 4405 38575
rect 4405 38541 4413 38575
rect 4361 38534 4413 38541
rect 4553 38575 4605 38586
rect 4553 38541 4563 38575
rect 4563 38541 4597 38575
rect 4597 38541 4605 38575
rect 4553 38534 4605 38541
rect 4746 38575 4798 38585
rect 4746 38541 4755 38575
rect 4755 38541 4789 38575
rect 4789 38541 4798 38575
rect 4746 38533 4798 38541
rect 4938 38575 4990 38585
rect 4938 38541 4947 38575
rect 4947 38541 4981 38575
rect 4981 38541 4990 38575
rect 4938 38533 4990 38541
rect 304 38092 356 38102
rect 304 38058 313 38092
rect 313 38058 347 38092
rect 347 38058 356 38092
rect 304 38050 356 38058
rect 497 38092 549 38102
rect 497 38058 505 38092
rect 505 38058 539 38092
rect 539 38058 549 38092
rect 497 38050 549 38058
rect 688 38092 740 38102
rect 688 38058 697 38092
rect 697 38058 731 38092
rect 731 38058 740 38092
rect 688 38050 740 38058
rect 880 38092 932 38102
rect 880 38058 889 38092
rect 889 38058 923 38092
rect 923 38058 932 38092
rect 880 38050 932 38058
rect 1072 38092 1124 38102
rect 1072 38058 1081 38092
rect 1081 38058 1115 38092
rect 1115 38058 1124 38092
rect 1072 38050 1124 38058
rect 1264 38092 1316 38102
rect 1264 38058 1273 38092
rect 1273 38058 1307 38092
rect 1307 38058 1316 38092
rect 1264 38050 1316 38058
rect 1522 38043 1578 38103
rect 1792 38043 1852 38103
rect 2056 37696 2190 37804
rect 2457 38096 2509 38106
rect 2457 38062 2466 38096
rect 2466 38062 2500 38096
rect 2500 38062 2509 38096
rect 2457 38054 2509 38062
rect 2650 38096 2702 38106
rect 2650 38062 2658 38096
rect 2658 38062 2692 38096
rect 2692 38062 2702 38096
rect 2650 38054 2702 38062
rect 2841 38096 2893 38106
rect 2841 38062 2850 38096
rect 2850 38062 2884 38096
rect 2884 38062 2893 38096
rect 2841 38054 2893 38062
rect 3033 38096 3085 38106
rect 3033 38062 3042 38096
rect 3042 38062 3076 38096
rect 3076 38062 3085 38096
rect 3033 38054 3085 38062
rect 3225 38096 3277 38106
rect 3225 38062 3234 38096
rect 3234 38062 3268 38096
rect 3268 38062 3277 38096
rect 3225 38054 3277 38062
rect 3417 38096 3469 38106
rect 3417 38062 3426 38096
rect 3426 38062 3460 38096
rect 3460 38062 3469 38096
rect 3417 38054 3469 38062
rect 1608 37336 1720 37460
rect 304 37284 356 37295
rect 304 37250 313 37284
rect 313 37250 347 37284
rect 347 37250 356 37284
rect 304 37243 356 37250
rect 495 37284 547 37295
rect 495 37250 505 37284
rect 505 37250 539 37284
rect 539 37250 547 37284
rect 495 37243 547 37250
rect 687 37284 739 37295
rect 687 37250 697 37284
rect 697 37250 731 37284
rect 731 37250 739 37284
rect 687 37243 739 37250
rect 879 37284 931 37295
rect 879 37250 889 37284
rect 889 37250 923 37284
rect 923 37250 931 37284
rect 879 37243 931 37250
rect 1072 37284 1124 37294
rect 1072 37250 1081 37284
rect 1081 37250 1115 37284
rect 1115 37250 1124 37284
rect 1072 37242 1124 37250
rect 1264 37284 1316 37294
rect 1264 37250 1273 37284
rect 1273 37250 1307 37284
rect 1307 37250 1316 37284
rect 1264 37242 1316 37250
rect 1468 37242 1524 37298
rect 1930 37244 1986 37300
rect 3978 38096 4030 38106
rect 3978 38062 3987 38096
rect 3987 38062 4021 38096
rect 4021 38062 4030 38096
rect 3978 38054 4030 38062
rect 4171 38096 4223 38106
rect 4171 38062 4179 38096
rect 4179 38062 4213 38096
rect 4213 38062 4223 38096
rect 4171 38054 4223 38062
rect 4362 38096 4414 38106
rect 4362 38062 4371 38096
rect 4371 38062 4405 38096
rect 4405 38062 4414 38096
rect 4362 38054 4414 38062
rect 4554 38096 4606 38106
rect 4554 38062 4563 38096
rect 4563 38062 4597 38096
rect 4597 38062 4606 38096
rect 4554 38054 4606 38062
rect 4746 38096 4798 38106
rect 4746 38062 4755 38096
rect 4755 38062 4789 38096
rect 4789 38062 4798 38096
rect 4746 38054 4798 38062
rect 4938 38096 4990 38106
rect 4938 38062 4947 38096
rect 4947 38062 4981 38096
rect 4981 38062 4990 38096
rect 4938 38054 4990 38062
rect 3681 37510 3733 37529
rect 3681 37477 3691 37510
rect 3691 37477 3725 37510
rect 3725 37477 3733 37510
rect 5337 37551 5389 37561
rect 5337 37517 5348 37551
rect 5348 37517 5382 37551
rect 5382 37517 5389 37551
rect 5337 37509 5389 37517
rect 5449 37556 5501 37563
rect 5449 37522 5450 37556
rect 5450 37522 5484 37556
rect 5484 37522 5501 37556
rect 5449 37511 5501 37522
rect 2457 37288 2509 37299
rect 2457 37254 2466 37288
rect 2466 37254 2500 37288
rect 2500 37254 2509 37288
rect 2457 37247 2509 37254
rect 2648 37288 2700 37299
rect 2648 37254 2658 37288
rect 2658 37254 2692 37288
rect 2692 37254 2700 37288
rect 2648 37247 2700 37254
rect 2840 37288 2892 37299
rect 2840 37254 2850 37288
rect 2850 37254 2884 37288
rect 2884 37254 2892 37288
rect 2840 37247 2892 37254
rect 3032 37288 3084 37299
rect 3032 37254 3042 37288
rect 3042 37254 3076 37288
rect 3076 37254 3084 37288
rect 3032 37247 3084 37254
rect 3225 37288 3277 37298
rect 3225 37254 3234 37288
rect 3234 37254 3268 37288
rect 3268 37254 3277 37288
rect 3225 37246 3277 37254
rect 3417 37288 3469 37298
rect 3417 37254 3426 37288
rect 3426 37254 3460 37288
rect 3460 37254 3469 37288
rect 3417 37246 3469 37254
rect 3978 37288 4030 37299
rect 3978 37254 3987 37288
rect 3987 37254 4021 37288
rect 4021 37254 4030 37288
rect 3978 37247 4030 37254
rect 4169 37288 4221 37299
rect 4169 37254 4179 37288
rect 4179 37254 4213 37288
rect 4213 37254 4221 37288
rect 4169 37247 4221 37254
rect 4361 37288 4413 37299
rect 4361 37254 4371 37288
rect 4371 37254 4405 37288
rect 4405 37254 4413 37288
rect 4361 37247 4413 37254
rect 4553 37288 4605 37299
rect 4553 37254 4563 37288
rect 4563 37254 4597 37288
rect 4597 37254 4605 37288
rect 4553 37247 4605 37254
rect 4746 37288 4798 37298
rect 4746 37254 4755 37288
rect 4755 37254 4789 37288
rect 4789 37254 4798 37288
rect 4746 37246 4798 37254
rect 4938 37288 4990 37298
rect 4938 37254 4947 37288
rect 4947 37254 4981 37288
rect 4981 37254 4990 37288
rect 4938 37246 4990 37254
rect 304 36805 356 36815
rect 304 36771 313 36805
rect 313 36771 347 36805
rect 347 36771 356 36805
rect 304 36763 356 36771
rect 497 36805 549 36815
rect 497 36771 505 36805
rect 505 36771 539 36805
rect 539 36771 549 36805
rect 497 36763 549 36771
rect 688 36805 740 36815
rect 688 36771 697 36805
rect 697 36771 731 36805
rect 731 36771 740 36805
rect 688 36763 740 36771
rect 880 36805 932 36815
rect 880 36771 889 36805
rect 889 36771 923 36805
rect 923 36771 932 36805
rect 880 36763 932 36771
rect 1072 36805 1124 36815
rect 1072 36771 1081 36805
rect 1081 36771 1115 36805
rect 1115 36771 1124 36805
rect 1072 36763 1124 36771
rect 1264 36805 1316 36815
rect 1264 36771 1273 36805
rect 1273 36771 1307 36805
rect 1307 36771 1316 36805
rect 1264 36763 1316 36771
rect 1522 36756 1578 36816
rect 1792 36756 1852 36816
rect 2056 36409 2190 36517
rect 2457 36809 2509 36819
rect 2457 36775 2466 36809
rect 2466 36775 2500 36809
rect 2500 36775 2509 36809
rect 2457 36767 2509 36775
rect 2650 36809 2702 36819
rect 2650 36775 2658 36809
rect 2658 36775 2692 36809
rect 2692 36775 2702 36809
rect 2650 36767 2702 36775
rect 2841 36809 2893 36819
rect 2841 36775 2850 36809
rect 2850 36775 2884 36809
rect 2884 36775 2893 36809
rect 2841 36767 2893 36775
rect 3033 36809 3085 36819
rect 3033 36775 3042 36809
rect 3042 36775 3076 36809
rect 3076 36775 3085 36809
rect 3033 36767 3085 36775
rect 3225 36809 3277 36819
rect 3225 36775 3234 36809
rect 3234 36775 3268 36809
rect 3268 36775 3277 36809
rect 3225 36767 3277 36775
rect 3417 36809 3469 36819
rect 3417 36775 3426 36809
rect 3426 36775 3460 36809
rect 3460 36775 3469 36809
rect 3417 36767 3469 36775
rect 1608 36049 1720 36173
rect 304 35997 356 36008
rect 304 35963 313 35997
rect 313 35963 347 35997
rect 347 35963 356 35997
rect 304 35956 356 35963
rect 495 35997 547 36008
rect 495 35963 505 35997
rect 505 35963 539 35997
rect 539 35963 547 35997
rect 495 35956 547 35963
rect 687 35997 739 36008
rect 687 35963 697 35997
rect 697 35963 731 35997
rect 731 35963 739 35997
rect 687 35956 739 35963
rect 879 35997 931 36008
rect 879 35963 889 35997
rect 889 35963 923 35997
rect 923 35963 931 35997
rect 879 35956 931 35963
rect 1072 35997 1124 36007
rect 1072 35963 1081 35997
rect 1081 35963 1115 35997
rect 1115 35963 1124 35997
rect 1072 35955 1124 35963
rect 1264 35997 1316 36007
rect 1264 35963 1273 35997
rect 1273 35963 1307 35997
rect 1307 35963 1316 35997
rect 1264 35955 1316 35963
rect 1468 35955 1524 36011
rect 1930 35957 1986 36013
rect 3978 36809 4030 36819
rect 3978 36775 3987 36809
rect 3987 36775 4021 36809
rect 4021 36775 4030 36809
rect 3978 36767 4030 36775
rect 4171 36809 4223 36819
rect 4171 36775 4179 36809
rect 4179 36775 4213 36809
rect 4213 36775 4223 36809
rect 4171 36767 4223 36775
rect 4362 36809 4414 36819
rect 4362 36775 4371 36809
rect 4371 36775 4405 36809
rect 4405 36775 4414 36809
rect 4362 36767 4414 36775
rect 4554 36809 4606 36819
rect 4554 36775 4563 36809
rect 4563 36775 4597 36809
rect 4597 36775 4606 36809
rect 4554 36767 4606 36775
rect 4746 36809 4798 36819
rect 4746 36775 4755 36809
rect 4755 36775 4789 36809
rect 4789 36775 4798 36809
rect 4746 36767 4798 36775
rect 4938 36809 4990 36819
rect 4938 36775 4947 36809
rect 4947 36775 4981 36809
rect 4981 36775 4990 36809
rect 4938 36767 4990 36775
rect 3681 36223 3733 36242
rect 3681 36190 3691 36223
rect 3691 36190 3725 36223
rect 3725 36190 3733 36223
rect 5337 36264 5389 36274
rect 5337 36230 5348 36264
rect 5348 36230 5382 36264
rect 5382 36230 5389 36264
rect 5337 36222 5389 36230
rect 5449 36269 5501 36276
rect 5449 36235 5450 36269
rect 5450 36235 5484 36269
rect 5484 36235 5501 36269
rect 5449 36224 5501 36235
rect 2457 36001 2509 36012
rect 2457 35967 2466 36001
rect 2466 35967 2500 36001
rect 2500 35967 2509 36001
rect 2457 35960 2509 35967
rect 2648 36001 2700 36012
rect 2648 35967 2658 36001
rect 2658 35967 2692 36001
rect 2692 35967 2700 36001
rect 2648 35960 2700 35967
rect 2840 36001 2892 36012
rect 2840 35967 2850 36001
rect 2850 35967 2884 36001
rect 2884 35967 2892 36001
rect 2840 35960 2892 35967
rect 3032 36001 3084 36012
rect 3032 35967 3042 36001
rect 3042 35967 3076 36001
rect 3076 35967 3084 36001
rect 3032 35960 3084 35967
rect 3225 36001 3277 36011
rect 3225 35967 3234 36001
rect 3234 35967 3268 36001
rect 3268 35967 3277 36001
rect 3225 35959 3277 35967
rect 3417 36001 3469 36011
rect 3417 35967 3426 36001
rect 3426 35967 3460 36001
rect 3460 35967 3469 36001
rect 3417 35959 3469 35967
rect 3978 36001 4030 36012
rect 3978 35967 3987 36001
rect 3987 35967 4021 36001
rect 4021 35967 4030 36001
rect 3978 35960 4030 35967
rect 4169 36001 4221 36012
rect 4169 35967 4179 36001
rect 4179 35967 4213 36001
rect 4213 35967 4221 36001
rect 4169 35960 4221 35967
rect 4361 36001 4413 36012
rect 4361 35967 4371 36001
rect 4371 35967 4405 36001
rect 4405 35967 4413 36001
rect 4361 35960 4413 35967
rect 4553 36001 4605 36012
rect 4553 35967 4563 36001
rect 4563 35967 4597 36001
rect 4597 35967 4605 36001
rect 4553 35960 4605 35967
rect 4746 36001 4798 36011
rect 4746 35967 4755 36001
rect 4755 35967 4789 36001
rect 4789 35967 4798 36001
rect 4746 35959 4798 35967
rect 4938 36001 4990 36011
rect 4938 35967 4947 36001
rect 4947 35967 4981 36001
rect 4981 35967 4990 36001
rect 4938 35959 4990 35967
rect 304 35518 356 35528
rect 304 35484 313 35518
rect 313 35484 347 35518
rect 347 35484 356 35518
rect 304 35476 356 35484
rect 497 35518 549 35528
rect 497 35484 505 35518
rect 505 35484 539 35518
rect 539 35484 549 35518
rect 497 35476 549 35484
rect 688 35518 740 35528
rect 688 35484 697 35518
rect 697 35484 731 35518
rect 731 35484 740 35518
rect 688 35476 740 35484
rect 880 35518 932 35528
rect 880 35484 889 35518
rect 889 35484 923 35518
rect 923 35484 932 35518
rect 880 35476 932 35484
rect 1072 35518 1124 35528
rect 1072 35484 1081 35518
rect 1081 35484 1115 35518
rect 1115 35484 1124 35518
rect 1072 35476 1124 35484
rect 1264 35518 1316 35528
rect 1264 35484 1273 35518
rect 1273 35484 1307 35518
rect 1307 35484 1316 35518
rect 1264 35476 1316 35484
rect 1522 35469 1578 35529
rect 1792 35469 1852 35529
rect 2056 35122 2190 35230
rect 2457 35522 2509 35532
rect 2457 35488 2466 35522
rect 2466 35488 2500 35522
rect 2500 35488 2509 35522
rect 2457 35480 2509 35488
rect 2650 35522 2702 35532
rect 2650 35488 2658 35522
rect 2658 35488 2692 35522
rect 2692 35488 2702 35522
rect 2650 35480 2702 35488
rect 2841 35522 2893 35532
rect 2841 35488 2850 35522
rect 2850 35488 2884 35522
rect 2884 35488 2893 35522
rect 2841 35480 2893 35488
rect 3033 35522 3085 35532
rect 3033 35488 3042 35522
rect 3042 35488 3076 35522
rect 3076 35488 3085 35522
rect 3033 35480 3085 35488
rect 3225 35522 3277 35532
rect 3225 35488 3234 35522
rect 3234 35488 3268 35522
rect 3268 35488 3277 35522
rect 3225 35480 3277 35488
rect 3417 35522 3469 35532
rect 3417 35488 3426 35522
rect 3426 35488 3460 35522
rect 3460 35488 3469 35522
rect 3417 35480 3469 35488
rect 1608 34762 1720 34886
rect 304 34710 356 34721
rect 304 34676 313 34710
rect 313 34676 347 34710
rect 347 34676 356 34710
rect 304 34669 356 34676
rect 495 34710 547 34721
rect 495 34676 505 34710
rect 505 34676 539 34710
rect 539 34676 547 34710
rect 495 34669 547 34676
rect 687 34710 739 34721
rect 687 34676 697 34710
rect 697 34676 731 34710
rect 731 34676 739 34710
rect 687 34669 739 34676
rect 879 34710 931 34721
rect 879 34676 889 34710
rect 889 34676 923 34710
rect 923 34676 931 34710
rect 879 34669 931 34676
rect 1072 34710 1124 34720
rect 1072 34676 1081 34710
rect 1081 34676 1115 34710
rect 1115 34676 1124 34710
rect 1072 34668 1124 34676
rect 1264 34710 1316 34720
rect 1264 34676 1273 34710
rect 1273 34676 1307 34710
rect 1307 34676 1316 34710
rect 1264 34668 1316 34676
rect 1468 34668 1524 34724
rect 1930 34670 1986 34726
rect 3978 35522 4030 35532
rect 3978 35488 3987 35522
rect 3987 35488 4021 35522
rect 4021 35488 4030 35522
rect 3978 35480 4030 35488
rect 4171 35522 4223 35532
rect 4171 35488 4179 35522
rect 4179 35488 4213 35522
rect 4213 35488 4223 35522
rect 4171 35480 4223 35488
rect 4362 35522 4414 35532
rect 4362 35488 4371 35522
rect 4371 35488 4405 35522
rect 4405 35488 4414 35522
rect 4362 35480 4414 35488
rect 4554 35522 4606 35532
rect 4554 35488 4563 35522
rect 4563 35488 4597 35522
rect 4597 35488 4606 35522
rect 4554 35480 4606 35488
rect 4746 35522 4798 35532
rect 4746 35488 4755 35522
rect 4755 35488 4789 35522
rect 4789 35488 4798 35522
rect 4746 35480 4798 35488
rect 4938 35522 4990 35532
rect 4938 35488 4947 35522
rect 4947 35488 4981 35522
rect 4981 35488 4990 35522
rect 4938 35480 4990 35488
rect 3681 34936 3733 34955
rect 3681 34903 3691 34936
rect 3691 34903 3725 34936
rect 3725 34903 3733 34936
rect 5337 34977 5389 34987
rect 5337 34943 5348 34977
rect 5348 34943 5382 34977
rect 5382 34943 5389 34977
rect 5337 34935 5389 34943
rect 5449 34982 5501 34989
rect 5449 34948 5450 34982
rect 5450 34948 5484 34982
rect 5484 34948 5501 34982
rect 5449 34937 5501 34948
rect 2457 34714 2509 34725
rect 2457 34680 2466 34714
rect 2466 34680 2500 34714
rect 2500 34680 2509 34714
rect 2457 34673 2509 34680
rect 2648 34714 2700 34725
rect 2648 34680 2658 34714
rect 2658 34680 2692 34714
rect 2692 34680 2700 34714
rect 2648 34673 2700 34680
rect 2840 34714 2892 34725
rect 2840 34680 2850 34714
rect 2850 34680 2884 34714
rect 2884 34680 2892 34714
rect 2840 34673 2892 34680
rect 3032 34714 3084 34725
rect 3032 34680 3042 34714
rect 3042 34680 3076 34714
rect 3076 34680 3084 34714
rect 3032 34673 3084 34680
rect 3225 34714 3277 34724
rect 3225 34680 3234 34714
rect 3234 34680 3268 34714
rect 3268 34680 3277 34714
rect 3225 34672 3277 34680
rect 3417 34714 3469 34724
rect 3417 34680 3426 34714
rect 3426 34680 3460 34714
rect 3460 34680 3469 34714
rect 3417 34672 3469 34680
rect 3978 34714 4030 34725
rect 3978 34680 3987 34714
rect 3987 34680 4021 34714
rect 4021 34680 4030 34714
rect 3978 34673 4030 34680
rect 4169 34714 4221 34725
rect 4169 34680 4179 34714
rect 4179 34680 4213 34714
rect 4213 34680 4221 34714
rect 4169 34673 4221 34680
rect 4361 34714 4413 34725
rect 4361 34680 4371 34714
rect 4371 34680 4405 34714
rect 4405 34680 4413 34714
rect 4361 34673 4413 34680
rect 4553 34714 4605 34725
rect 4553 34680 4563 34714
rect 4563 34680 4597 34714
rect 4597 34680 4605 34714
rect 4553 34673 4605 34680
rect 4746 34714 4798 34724
rect 4746 34680 4755 34714
rect 4755 34680 4789 34714
rect 4789 34680 4798 34714
rect 4746 34672 4798 34680
rect 4938 34714 4990 34724
rect 4938 34680 4947 34714
rect 4947 34680 4981 34714
rect 4981 34680 4990 34714
rect 4938 34672 4990 34680
rect 304 34231 356 34241
rect 304 34197 313 34231
rect 313 34197 347 34231
rect 347 34197 356 34231
rect 304 34189 356 34197
rect 497 34231 549 34241
rect 497 34197 505 34231
rect 505 34197 539 34231
rect 539 34197 549 34231
rect 497 34189 549 34197
rect 688 34231 740 34241
rect 688 34197 697 34231
rect 697 34197 731 34231
rect 731 34197 740 34231
rect 688 34189 740 34197
rect 880 34231 932 34241
rect 880 34197 889 34231
rect 889 34197 923 34231
rect 923 34197 932 34231
rect 880 34189 932 34197
rect 1072 34231 1124 34241
rect 1072 34197 1081 34231
rect 1081 34197 1115 34231
rect 1115 34197 1124 34231
rect 1072 34189 1124 34197
rect 1264 34231 1316 34241
rect 1264 34197 1273 34231
rect 1273 34197 1307 34231
rect 1307 34197 1316 34231
rect 1264 34189 1316 34197
rect 1522 34182 1578 34242
rect 1792 34182 1852 34242
rect 2056 33835 2190 33943
rect 2457 34235 2509 34245
rect 2457 34201 2466 34235
rect 2466 34201 2500 34235
rect 2500 34201 2509 34235
rect 2457 34193 2509 34201
rect 2650 34235 2702 34245
rect 2650 34201 2658 34235
rect 2658 34201 2692 34235
rect 2692 34201 2702 34235
rect 2650 34193 2702 34201
rect 2841 34235 2893 34245
rect 2841 34201 2850 34235
rect 2850 34201 2884 34235
rect 2884 34201 2893 34235
rect 2841 34193 2893 34201
rect 3033 34235 3085 34245
rect 3033 34201 3042 34235
rect 3042 34201 3076 34235
rect 3076 34201 3085 34235
rect 3033 34193 3085 34201
rect 3225 34235 3277 34245
rect 3225 34201 3234 34235
rect 3234 34201 3268 34235
rect 3268 34201 3277 34235
rect 3225 34193 3277 34201
rect 3417 34235 3469 34245
rect 3417 34201 3426 34235
rect 3426 34201 3460 34235
rect 3460 34201 3469 34235
rect 3417 34193 3469 34201
rect 1608 33475 1720 33599
rect 304 33423 356 33434
rect 304 33389 313 33423
rect 313 33389 347 33423
rect 347 33389 356 33423
rect 304 33382 356 33389
rect 495 33423 547 33434
rect 495 33389 505 33423
rect 505 33389 539 33423
rect 539 33389 547 33423
rect 495 33382 547 33389
rect 687 33423 739 33434
rect 687 33389 697 33423
rect 697 33389 731 33423
rect 731 33389 739 33423
rect 687 33382 739 33389
rect 879 33423 931 33434
rect 879 33389 889 33423
rect 889 33389 923 33423
rect 923 33389 931 33423
rect 879 33382 931 33389
rect 1072 33423 1124 33433
rect 1072 33389 1081 33423
rect 1081 33389 1115 33423
rect 1115 33389 1124 33423
rect 1072 33381 1124 33389
rect 1264 33423 1316 33433
rect 1264 33389 1273 33423
rect 1273 33389 1307 33423
rect 1307 33389 1316 33423
rect 1264 33381 1316 33389
rect 1468 33381 1524 33437
rect 1930 33383 1986 33439
rect 3978 34235 4030 34245
rect 3978 34201 3987 34235
rect 3987 34201 4021 34235
rect 4021 34201 4030 34235
rect 3978 34193 4030 34201
rect 4171 34235 4223 34245
rect 4171 34201 4179 34235
rect 4179 34201 4213 34235
rect 4213 34201 4223 34235
rect 4171 34193 4223 34201
rect 4362 34235 4414 34245
rect 4362 34201 4371 34235
rect 4371 34201 4405 34235
rect 4405 34201 4414 34235
rect 4362 34193 4414 34201
rect 4554 34235 4606 34245
rect 4554 34201 4563 34235
rect 4563 34201 4597 34235
rect 4597 34201 4606 34235
rect 4554 34193 4606 34201
rect 4746 34235 4798 34245
rect 4746 34201 4755 34235
rect 4755 34201 4789 34235
rect 4789 34201 4798 34235
rect 4746 34193 4798 34201
rect 4938 34235 4990 34245
rect 4938 34201 4947 34235
rect 4947 34201 4981 34235
rect 4981 34201 4990 34235
rect 4938 34193 4990 34201
rect 3681 33649 3733 33668
rect 3681 33616 3691 33649
rect 3691 33616 3725 33649
rect 3725 33616 3733 33649
rect 5337 33690 5389 33700
rect 5337 33656 5348 33690
rect 5348 33656 5382 33690
rect 5382 33656 5389 33690
rect 5337 33648 5389 33656
rect 5449 33695 5501 33702
rect 5449 33661 5450 33695
rect 5450 33661 5484 33695
rect 5484 33661 5501 33695
rect 5449 33650 5501 33661
rect 2457 33427 2509 33438
rect 2457 33393 2466 33427
rect 2466 33393 2500 33427
rect 2500 33393 2509 33427
rect 2457 33386 2509 33393
rect 2648 33427 2700 33438
rect 2648 33393 2658 33427
rect 2658 33393 2692 33427
rect 2692 33393 2700 33427
rect 2648 33386 2700 33393
rect 2840 33427 2892 33438
rect 2840 33393 2850 33427
rect 2850 33393 2884 33427
rect 2884 33393 2892 33427
rect 2840 33386 2892 33393
rect 3032 33427 3084 33438
rect 3032 33393 3042 33427
rect 3042 33393 3076 33427
rect 3076 33393 3084 33427
rect 3032 33386 3084 33393
rect 3225 33427 3277 33437
rect 3225 33393 3234 33427
rect 3234 33393 3268 33427
rect 3268 33393 3277 33427
rect 3225 33385 3277 33393
rect 3417 33427 3469 33437
rect 3417 33393 3426 33427
rect 3426 33393 3460 33427
rect 3460 33393 3469 33427
rect 3417 33385 3469 33393
rect 3978 33427 4030 33438
rect 3978 33393 3987 33427
rect 3987 33393 4021 33427
rect 4021 33393 4030 33427
rect 3978 33386 4030 33393
rect 4169 33427 4221 33438
rect 4169 33393 4179 33427
rect 4179 33393 4213 33427
rect 4213 33393 4221 33427
rect 4169 33386 4221 33393
rect 4361 33427 4413 33438
rect 4361 33393 4371 33427
rect 4371 33393 4405 33427
rect 4405 33393 4413 33427
rect 4361 33386 4413 33393
rect 4553 33427 4605 33438
rect 4553 33393 4563 33427
rect 4563 33393 4597 33427
rect 4597 33393 4605 33427
rect 4553 33386 4605 33393
rect 4746 33427 4798 33437
rect 4746 33393 4755 33427
rect 4755 33393 4789 33427
rect 4789 33393 4798 33427
rect 4746 33385 4798 33393
rect 4938 33427 4990 33437
rect 4938 33393 4947 33427
rect 4947 33393 4981 33427
rect 4981 33393 4990 33427
rect 4938 33385 4990 33393
rect 304 32944 356 32954
rect 304 32910 313 32944
rect 313 32910 347 32944
rect 347 32910 356 32944
rect 304 32902 356 32910
rect 497 32944 549 32954
rect 497 32910 505 32944
rect 505 32910 539 32944
rect 539 32910 549 32944
rect 497 32902 549 32910
rect 688 32944 740 32954
rect 688 32910 697 32944
rect 697 32910 731 32944
rect 731 32910 740 32944
rect 688 32902 740 32910
rect 880 32944 932 32954
rect 880 32910 889 32944
rect 889 32910 923 32944
rect 923 32910 932 32944
rect 880 32902 932 32910
rect 1072 32944 1124 32954
rect 1072 32910 1081 32944
rect 1081 32910 1115 32944
rect 1115 32910 1124 32944
rect 1072 32902 1124 32910
rect 1264 32944 1316 32954
rect 1264 32910 1273 32944
rect 1273 32910 1307 32944
rect 1307 32910 1316 32944
rect 1264 32902 1316 32910
rect 1522 32895 1578 32955
rect 1792 32895 1852 32955
rect 2056 32548 2190 32656
rect 2457 32948 2509 32958
rect 2457 32914 2466 32948
rect 2466 32914 2500 32948
rect 2500 32914 2509 32948
rect 2457 32906 2509 32914
rect 2650 32948 2702 32958
rect 2650 32914 2658 32948
rect 2658 32914 2692 32948
rect 2692 32914 2702 32948
rect 2650 32906 2702 32914
rect 2841 32948 2893 32958
rect 2841 32914 2850 32948
rect 2850 32914 2884 32948
rect 2884 32914 2893 32948
rect 2841 32906 2893 32914
rect 3033 32948 3085 32958
rect 3033 32914 3042 32948
rect 3042 32914 3076 32948
rect 3076 32914 3085 32948
rect 3033 32906 3085 32914
rect 3225 32948 3277 32958
rect 3225 32914 3234 32948
rect 3234 32914 3268 32948
rect 3268 32914 3277 32948
rect 3225 32906 3277 32914
rect 3417 32948 3469 32958
rect 3417 32914 3426 32948
rect 3426 32914 3460 32948
rect 3460 32914 3469 32948
rect 3417 32906 3469 32914
rect 1608 32188 1720 32312
rect 304 32136 356 32147
rect 304 32102 313 32136
rect 313 32102 347 32136
rect 347 32102 356 32136
rect 304 32095 356 32102
rect 495 32136 547 32147
rect 495 32102 505 32136
rect 505 32102 539 32136
rect 539 32102 547 32136
rect 495 32095 547 32102
rect 687 32136 739 32147
rect 687 32102 697 32136
rect 697 32102 731 32136
rect 731 32102 739 32136
rect 687 32095 739 32102
rect 879 32136 931 32147
rect 879 32102 889 32136
rect 889 32102 923 32136
rect 923 32102 931 32136
rect 879 32095 931 32102
rect 1072 32136 1124 32146
rect 1072 32102 1081 32136
rect 1081 32102 1115 32136
rect 1115 32102 1124 32136
rect 1072 32094 1124 32102
rect 1264 32136 1316 32146
rect 1264 32102 1273 32136
rect 1273 32102 1307 32136
rect 1307 32102 1316 32136
rect 1264 32094 1316 32102
rect 1468 32094 1524 32150
rect 1930 32096 1986 32152
rect 3978 32948 4030 32958
rect 3978 32914 3987 32948
rect 3987 32914 4021 32948
rect 4021 32914 4030 32948
rect 3978 32906 4030 32914
rect 4171 32948 4223 32958
rect 4171 32914 4179 32948
rect 4179 32914 4213 32948
rect 4213 32914 4223 32948
rect 4171 32906 4223 32914
rect 4362 32948 4414 32958
rect 4362 32914 4371 32948
rect 4371 32914 4405 32948
rect 4405 32914 4414 32948
rect 4362 32906 4414 32914
rect 4554 32948 4606 32958
rect 4554 32914 4563 32948
rect 4563 32914 4597 32948
rect 4597 32914 4606 32948
rect 4554 32906 4606 32914
rect 4746 32948 4798 32958
rect 4746 32914 4755 32948
rect 4755 32914 4789 32948
rect 4789 32914 4798 32948
rect 4746 32906 4798 32914
rect 4938 32948 4990 32958
rect 4938 32914 4947 32948
rect 4947 32914 4981 32948
rect 4981 32914 4990 32948
rect 4938 32906 4990 32914
rect 3681 32362 3733 32381
rect 3681 32329 3691 32362
rect 3691 32329 3725 32362
rect 3725 32329 3733 32362
rect 5337 32403 5389 32413
rect 5337 32369 5348 32403
rect 5348 32369 5382 32403
rect 5382 32369 5389 32403
rect 5337 32361 5389 32369
rect 5449 32408 5501 32415
rect 5449 32374 5450 32408
rect 5450 32374 5484 32408
rect 5484 32374 5501 32408
rect 5449 32363 5501 32374
rect 2457 32140 2509 32151
rect 2457 32106 2466 32140
rect 2466 32106 2500 32140
rect 2500 32106 2509 32140
rect 2457 32099 2509 32106
rect 2648 32140 2700 32151
rect 2648 32106 2658 32140
rect 2658 32106 2692 32140
rect 2692 32106 2700 32140
rect 2648 32099 2700 32106
rect 2840 32140 2892 32151
rect 2840 32106 2850 32140
rect 2850 32106 2884 32140
rect 2884 32106 2892 32140
rect 2840 32099 2892 32106
rect 3032 32140 3084 32151
rect 3032 32106 3042 32140
rect 3042 32106 3076 32140
rect 3076 32106 3084 32140
rect 3032 32099 3084 32106
rect 3225 32140 3277 32150
rect 3225 32106 3234 32140
rect 3234 32106 3268 32140
rect 3268 32106 3277 32140
rect 3225 32098 3277 32106
rect 3417 32140 3469 32150
rect 3417 32106 3426 32140
rect 3426 32106 3460 32140
rect 3460 32106 3469 32140
rect 3417 32098 3469 32106
rect 3978 32140 4030 32151
rect 3978 32106 3987 32140
rect 3987 32106 4021 32140
rect 4021 32106 4030 32140
rect 3978 32099 4030 32106
rect 4169 32140 4221 32151
rect 4169 32106 4179 32140
rect 4179 32106 4213 32140
rect 4213 32106 4221 32140
rect 4169 32099 4221 32106
rect 4361 32140 4413 32151
rect 4361 32106 4371 32140
rect 4371 32106 4405 32140
rect 4405 32106 4413 32140
rect 4361 32099 4413 32106
rect 4553 32140 4605 32151
rect 4553 32106 4563 32140
rect 4563 32106 4597 32140
rect 4597 32106 4605 32140
rect 4553 32099 4605 32106
rect 4746 32140 4798 32150
rect 4746 32106 4755 32140
rect 4755 32106 4789 32140
rect 4789 32106 4798 32140
rect 4746 32098 4798 32106
rect 4938 32140 4990 32150
rect 4938 32106 4947 32140
rect 4947 32106 4981 32140
rect 4981 32106 4990 32140
rect 4938 32098 4990 32106
rect 304 31657 356 31667
rect 304 31623 313 31657
rect 313 31623 347 31657
rect 347 31623 356 31657
rect 304 31615 356 31623
rect 497 31657 549 31667
rect 497 31623 505 31657
rect 505 31623 539 31657
rect 539 31623 549 31657
rect 497 31615 549 31623
rect 688 31657 740 31667
rect 688 31623 697 31657
rect 697 31623 731 31657
rect 731 31623 740 31657
rect 688 31615 740 31623
rect 880 31657 932 31667
rect 880 31623 889 31657
rect 889 31623 923 31657
rect 923 31623 932 31657
rect 880 31615 932 31623
rect 1072 31657 1124 31667
rect 1072 31623 1081 31657
rect 1081 31623 1115 31657
rect 1115 31623 1124 31657
rect 1072 31615 1124 31623
rect 1264 31657 1316 31667
rect 1264 31623 1273 31657
rect 1273 31623 1307 31657
rect 1307 31623 1316 31657
rect 1264 31615 1316 31623
rect 1522 31608 1578 31668
rect 1792 31608 1852 31668
rect 2056 31261 2190 31369
rect 2457 31661 2509 31671
rect 2457 31627 2466 31661
rect 2466 31627 2500 31661
rect 2500 31627 2509 31661
rect 2457 31619 2509 31627
rect 2650 31661 2702 31671
rect 2650 31627 2658 31661
rect 2658 31627 2692 31661
rect 2692 31627 2702 31661
rect 2650 31619 2702 31627
rect 2841 31661 2893 31671
rect 2841 31627 2850 31661
rect 2850 31627 2884 31661
rect 2884 31627 2893 31661
rect 2841 31619 2893 31627
rect 3033 31661 3085 31671
rect 3033 31627 3042 31661
rect 3042 31627 3076 31661
rect 3076 31627 3085 31661
rect 3033 31619 3085 31627
rect 3225 31661 3277 31671
rect 3225 31627 3234 31661
rect 3234 31627 3268 31661
rect 3268 31627 3277 31661
rect 3225 31619 3277 31627
rect 3417 31661 3469 31671
rect 3417 31627 3426 31661
rect 3426 31627 3460 31661
rect 3460 31627 3469 31661
rect 3417 31619 3469 31627
rect 1608 30901 1720 31025
rect 304 30849 356 30860
rect 304 30815 313 30849
rect 313 30815 347 30849
rect 347 30815 356 30849
rect 304 30808 356 30815
rect 495 30849 547 30860
rect 495 30815 505 30849
rect 505 30815 539 30849
rect 539 30815 547 30849
rect 495 30808 547 30815
rect 687 30849 739 30860
rect 687 30815 697 30849
rect 697 30815 731 30849
rect 731 30815 739 30849
rect 687 30808 739 30815
rect 879 30849 931 30860
rect 879 30815 889 30849
rect 889 30815 923 30849
rect 923 30815 931 30849
rect 879 30808 931 30815
rect 1072 30849 1124 30859
rect 1072 30815 1081 30849
rect 1081 30815 1115 30849
rect 1115 30815 1124 30849
rect 1072 30807 1124 30815
rect 1264 30849 1316 30859
rect 1264 30815 1273 30849
rect 1273 30815 1307 30849
rect 1307 30815 1316 30849
rect 1264 30807 1316 30815
rect 1468 30807 1524 30863
rect 1930 30809 1986 30865
rect 3978 31661 4030 31671
rect 3978 31627 3987 31661
rect 3987 31627 4021 31661
rect 4021 31627 4030 31661
rect 3978 31619 4030 31627
rect 4171 31661 4223 31671
rect 4171 31627 4179 31661
rect 4179 31627 4213 31661
rect 4213 31627 4223 31661
rect 4171 31619 4223 31627
rect 4362 31661 4414 31671
rect 4362 31627 4371 31661
rect 4371 31627 4405 31661
rect 4405 31627 4414 31661
rect 4362 31619 4414 31627
rect 4554 31661 4606 31671
rect 4554 31627 4563 31661
rect 4563 31627 4597 31661
rect 4597 31627 4606 31661
rect 4554 31619 4606 31627
rect 4746 31661 4798 31671
rect 4746 31627 4755 31661
rect 4755 31627 4789 31661
rect 4789 31627 4798 31661
rect 4746 31619 4798 31627
rect 4938 31661 4990 31671
rect 4938 31627 4947 31661
rect 4947 31627 4981 31661
rect 4981 31627 4990 31661
rect 4938 31619 4990 31627
rect 3681 31075 3733 31094
rect 3681 31042 3691 31075
rect 3691 31042 3725 31075
rect 3725 31042 3733 31075
rect 5337 31116 5389 31126
rect 5337 31082 5348 31116
rect 5348 31082 5382 31116
rect 5382 31082 5389 31116
rect 5337 31074 5389 31082
rect 5449 31121 5501 31128
rect 5449 31087 5450 31121
rect 5450 31087 5484 31121
rect 5484 31087 5501 31121
rect 5449 31076 5501 31087
rect 2457 30853 2509 30864
rect 2457 30819 2466 30853
rect 2466 30819 2500 30853
rect 2500 30819 2509 30853
rect 2457 30812 2509 30819
rect 2648 30853 2700 30864
rect 2648 30819 2658 30853
rect 2658 30819 2692 30853
rect 2692 30819 2700 30853
rect 2648 30812 2700 30819
rect 2840 30853 2892 30864
rect 2840 30819 2850 30853
rect 2850 30819 2884 30853
rect 2884 30819 2892 30853
rect 2840 30812 2892 30819
rect 3032 30853 3084 30864
rect 3032 30819 3042 30853
rect 3042 30819 3076 30853
rect 3076 30819 3084 30853
rect 3032 30812 3084 30819
rect 3225 30853 3277 30863
rect 3225 30819 3234 30853
rect 3234 30819 3268 30853
rect 3268 30819 3277 30853
rect 3225 30811 3277 30819
rect 3417 30853 3469 30863
rect 3417 30819 3426 30853
rect 3426 30819 3460 30853
rect 3460 30819 3469 30853
rect 3417 30811 3469 30819
rect 3978 30853 4030 30864
rect 3978 30819 3987 30853
rect 3987 30819 4021 30853
rect 4021 30819 4030 30853
rect 3978 30812 4030 30819
rect 4169 30853 4221 30864
rect 4169 30819 4179 30853
rect 4179 30819 4213 30853
rect 4213 30819 4221 30853
rect 4169 30812 4221 30819
rect 4361 30853 4413 30864
rect 4361 30819 4371 30853
rect 4371 30819 4405 30853
rect 4405 30819 4413 30853
rect 4361 30812 4413 30819
rect 4553 30853 4605 30864
rect 4553 30819 4563 30853
rect 4563 30819 4597 30853
rect 4597 30819 4605 30853
rect 4553 30812 4605 30819
rect 4746 30853 4798 30863
rect 4746 30819 4755 30853
rect 4755 30819 4789 30853
rect 4789 30819 4798 30853
rect 4746 30811 4798 30819
rect 4938 30853 4990 30863
rect 4938 30819 4947 30853
rect 4947 30819 4981 30853
rect 4981 30819 4990 30853
rect 4938 30811 4990 30819
rect 304 30370 356 30380
rect 304 30336 313 30370
rect 313 30336 347 30370
rect 347 30336 356 30370
rect 304 30328 356 30336
rect 497 30370 549 30380
rect 497 30336 505 30370
rect 505 30336 539 30370
rect 539 30336 549 30370
rect 497 30328 549 30336
rect 688 30370 740 30380
rect 688 30336 697 30370
rect 697 30336 731 30370
rect 731 30336 740 30370
rect 688 30328 740 30336
rect 880 30370 932 30380
rect 880 30336 889 30370
rect 889 30336 923 30370
rect 923 30336 932 30370
rect 880 30328 932 30336
rect 1072 30370 1124 30380
rect 1072 30336 1081 30370
rect 1081 30336 1115 30370
rect 1115 30336 1124 30370
rect 1072 30328 1124 30336
rect 1264 30370 1316 30380
rect 1264 30336 1273 30370
rect 1273 30336 1307 30370
rect 1307 30336 1316 30370
rect 1264 30328 1316 30336
rect 1522 30321 1578 30381
rect 1792 30321 1852 30381
rect 2056 29974 2190 30082
rect 2457 30374 2509 30384
rect 2457 30340 2466 30374
rect 2466 30340 2500 30374
rect 2500 30340 2509 30374
rect 2457 30332 2509 30340
rect 2650 30374 2702 30384
rect 2650 30340 2658 30374
rect 2658 30340 2692 30374
rect 2692 30340 2702 30374
rect 2650 30332 2702 30340
rect 2841 30374 2893 30384
rect 2841 30340 2850 30374
rect 2850 30340 2884 30374
rect 2884 30340 2893 30374
rect 2841 30332 2893 30340
rect 3033 30374 3085 30384
rect 3033 30340 3042 30374
rect 3042 30340 3076 30374
rect 3076 30340 3085 30374
rect 3033 30332 3085 30340
rect 3225 30374 3277 30384
rect 3225 30340 3234 30374
rect 3234 30340 3268 30374
rect 3268 30340 3277 30374
rect 3225 30332 3277 30340
rect 3417 30374 3469 30384
rect 3417 30340 3426 30374
rect 3426 30340 3460 30374
rect 3460 30340 3469 30374
rect 3417 30332 3469 30340
rect 1608 29614 1720 29738
rect 304 29562 356 29573
rect 304 29528 313 29562
rect 313 29528 347 29562
rect 347 29528 356 29562
rect 304 29521 356 29528
rect 495 29562 547 29573
rect 495 29528 505 29562
rect 505 29528 539 29562
rect 539 29528 547 29562
rect 495 29521 547 29528
rect 687 29562 739 29573
rect 687 29528 697 29562
rect 697 29528 731 29562
rect 731 29528 739 29562
rect 687 29521 739 29528
rect 879 29562 931 29573
rect 879 29528 889 29562
rect 889 29528 923 29562
rect 923 29528 931 29562
rect 879 29521 931 29528
rect 1072 29562 1124 29572
rect 1072 29528 1081 29562
rect 1081 29528 1115 29562
rect 1115 29528 1124 29562
rect 1072 29520 1124 29528
rect 1264 29562 1316 29572
rect 1264 29528 1273 29562
rect 1273 29528 1307 29562
rect 1307 29528 1316 29562
rect 1264 29520 1316 29528
rect 1468 29520 1524 29576
rect 1930 29522 1986 29578
rect 3978 30374 4030 30384
rect 3978 30340 3987 30374
rect 3987 30340 4021 30374
rect 4021 30340 4030 30374
rect 3978 30332 4030 30340
rect 4171 30374 4223 30384
rect 4171 30340 4179 30374
rect 4179 30340 4213 30374
rect 4213 30340 4223 30374
rect 4171 30332 4223 30340
rect 4362 30374 4414 30384
rect 4362 30340 4371 30374
rect 4371 30340 4405 30374
rect 4405 30340 4414 30374
rect 4362 30332 4414 30340
rect 4554 30374 4606 30384
rect 4554 30340 4563 30374
rect 4563 30340 4597 30374
rect 4597 30340 4606 30374
rect 4554 30332 4606 30340
rect 4746 30374 4798 30384
rect 4746 30340 4755 30374
rect 4755 30340 4789 30374
rect 4789 30340 4798 30374
rect 4746 30332 4798 30340
rect 4938 30374 4990 30384
rect 4938 30340 4947 30374
rect 4947 30340 4981 30374
rect 4981 30340 4990 30374
rect 4938 30332 4990 30340
rect 3681 29788 3733 29807
rect 3681 29755 3691 29788
rect 3691 29755 3725 29788
rect 3725 29755 3733 29788
rect 5337 29829 5389 29839
rect 5337 29795 5348 29829
rect 5348 29795 5382 29829
rect 5382 29795 5389 29829
rect 5337 29787 5389 29795
rect 5449 29834 5501 29841
rect 5449 29800 5450 29834
rect 5450 29800 5484 29834
rect 5484 29800 5501 29834
rect 5449 29789 5501 29800
rect 2457 29566 2509 29577
rect 2457 29532 2466 29566
rect 2466 29532 2500 29566
rect 2500 29532 2509 29566
rect 2457 29525 2509 29532
rect 2648 29566 2700 29577
rect 2648 29532 2658 29566
rect 2658 29532 2692 29566
rect 2692 29532 2700 29566
rect 2648 29525 2700 29532
rect 2840 29566 2892 29577
rect 2840 29532 2850 29566
rect 2850 29532 2884 29566
rect 2884 29532 2892 29566
rect 2840 29525 2892 29532
rect 3032 29566 3084 29577
rect 3032 29532 3042 29566
rect 3042 29532 3076 29566
rect 3076 29532 3084 29566
rect 3032 29525 3084 29532
rect 3225 29566 3277 29576
rect 3225 29532 3234 29566
rect 3234 29532 3268 29566
rect 3268 29532 3277 29566
rect 3225 29524 3277 29532
rect 3417 29566 3469 29576
rect 3417 29532 3426 29566
rect 3426 29532 3460 29566
rect 3460 29532 3469 29566
rect 3417 29524 3469 29532
rect 3978 29566 4030 29577
rect 3978 29532 3987 29566
rect 3987 29532 4021 29566
rect 4021 29532 4030 29566
rect 3978 29525 4030 29532
rect 4169 29566 4221 29577
rect 4169 29532 4179 29566
rect 4179 29532 4213 29566
rect 4213 29532 4221 29566
rect 4169 29525 4221 29532
rect 4361 29566 4413 29577
rect 4361 29532 4371 29566
rect 4371 29532 4405 29566
rect 4405 29532 4413 29566
rect 4361 29525 4413 29532
rect 4553 29566 4605 29577
rect 4553 29532 4563 29566
rect 4563 29532 4597 29566
rect 4597 29532 4605 29566
rect 4553 29525 4605 29532
rect 4746 29566 4798 29576
rect 4746 29532 4755 29566
rect 4755 29532 4789 29566
rect 4789 29532 4798 29566
rect 4746 29524 4798 29532
rect 4938 29566 4990 29576
rect 4938 29532 4947 29566
rect 4947 29532 4981 29566
rect 4981 29532 4990 29566
rect 4938 29524 4990 29532
rect 304 29083 356 29093
rect 304 29049 313 29083
rect 313 29049 347 29083
rect 347 29049 356 29083
rect 304 29041 356 29049
rect 497 29083 549 29093
rect 497 29049 505 29083
rect 505 29049 539 29083
rect 539 29049 549 29083
rect 497 29041 549 29049
rect 688 29083 740 29093
rect 688 29049 697 29083
rect 697 29049 731 29083
rect 731 29049 740 29083
rect 688 29041 740 29049
rect 880 29083 932 29093
rect 880 29049 889 29083
rect 889 29049 923 29083
rect 923 29049 932 29083
rect 880 29041 932 29049
rect 1072 29083 1124 29093
rect 1072 29049 1081 29083
rect 1081 29049 1115 29083
rect 1115 29049 1124 29083
rect 1072 29041 1124 29049
rect 1264 29083 1316 29093
rect 1264 29049 1273 29083
rect 1273 29049 1307 29083
rect 1307 29049 1316 29083
rect 1264 29041 1316 29049
rect 1522 29034 1578 29094
rect 1792 29034 1852 29094
rect 2056 28687 2190 28795
rect 2457 29087 2509 29097
rect 2457 29053 2466 29087
rect 2466 29053 2500 29087
rect 2500 29053 2509 29087
rect 2457 29045 2509 29053
rect 2650 29087 2702 29097
rect 2650 29053 2658 29087
rect 2658 29053 2692 29087
rect 2692 29053 2702 29087
rect 2650 29045 2702 29053
rect 2841 29087 2893 29097
rect 2841 29053 2850 29087
rect 2850 29053 2884 29087
rect 2884 29053 2893 29087
rect 2841 29045 2893 29053
rect 3033 29087 3085 29097
rect 3033 29053 3042 29087
rect 3042 29053 3076 29087
rect 3076 29053 3085 29087
rect 3033 29045 3085 29053
rect 3225 29087 3277 29097
rect 3225 29053 3234 29087
rect 3234 29053 3268 29087
rect 3268 29053 3277 29087
rect 3225 29045 3277 29053
rect 3417 29087 3469 29097
rect 3417 29053 3426 29087
rect 3426 29053 3460 29087
rect 3460 29053 3469 29087
rect 3417 29045 3469 29053
rect 1608 28327 1720 28451
rect 304 28275 356 28286
rect 304 28241 313 28275
rect 313 28241 347 28275
rect 347 28241 356 28275
rect 304 28234 356 28241
rect 495 28275 547 28286
rect 495 28241 505 28275
rect 505 28241 539 28275
rect 539 28241 547 28275
rect 495 28234 547 28241
rect 687 28275 739 28286
rect 687 28241 697 28275
rect 697 28241 731 28275
rect 731 28241 739 28275
rect 687 28234 739 28241
rect 879 28275 931 28286
rect 879 28241 889 28275
rect 889 28241 923 28275
rect 923 28241 931 28275
rect 879 28234 931 28241
rect 1072 28275 1124 28285
rect 1072 28241 1081 28275
rect 1081 28241 1115 28275
rect 1115 28241 1124 28275
rect 1072 28233 1124 28241
rect 1264 28275 1316 28285
rect 1264 28241 1273 28275
rect 1273 28241 1307 28275
rect 1307 28241 1316 28275
rect 1264 28233 1316 28241
rect 1468 28233 1524 28289
rect 1930 28235 1986 28291
rect 3978 29087 4030 29097
rect 3978 29053 3987 29087
rect 3987 29053 4021 29087
rect 4021 29053 4030 29087
rect 3978 29045 4030 29053
rect 4171 29087 4223 29097
rect 4171 29053 4179 29087
rect 4179 29053 4213 29087
rect 4213 29053 4223 29087
rect 4171 29045 4223 29053
rect 4362 29087 4414 29097
rect 4362 29053 4371 29087
rect 4371 29053 4405 29087
rect 4405 29053 4414 29087
rect 4362 29045 4414 29053
rect 4554 29087 4606 29097
rect 4554 29053 4563 29087
rect 4563 29053 4597 29087
rect 4597 29053 4606 29087
rect 4554 29045 4606 29053
rect 4746 29087 4798 29097
rect 4746 29053 4755 29087
rect 4755 29053 4789 29087
rect 4789 29053 4798 29087
rect 4746 29045 4798 29053
rect 4938 29087 4990 29097
rect 4938 29053 4947 29087
rect 4947 29053 4981 29087
rect 4981 29053 4990 29087
rect 4938 29045 4990 29053
rect 3681 28501 3733 28520
rect 3681 28468 3691 28501
rect 3691 28468 3725 28501
rect 3725 28468 3733 28501
rect 5337 28542 5389 28552
rect 5337 28508 5348 28542
rect 5348 28508 5382 28542
rect 5382 28508 5389 28542
rect 5337 28500 5389 28508
rect 5449 28547 5501 28554
rect 5449 28513 5450 28547
rect 5450 28513 5484 28547
rect 5484 28513 5501 28547
rect 5449 28502 5501 28513
rect 2457 28279 2509 28290
rect 2457 28245 2466 28279
rect 2466 28245 2500 28279
rect 2500 28245 2509 28279
rect 2457 28238 2509 28245
rect 2648 28279 2700 28290
rect 2648 28245 2658 28279
rect 2658 28245 2692 28279
rect 2692 28245 2700 28279
rect 2648 28238 2700 28245
rect 2840 28279 2892 28290
rect 2840 28245 2850 28279
rect 2850 28245 2884 28279
rect 2884 28245 2892 28279
rect 2840 28238 2892 28245
rect 3032 28279 3084 28290
rect 3032 28245 3042 28279
rect 3042 28245 3076 28279
rect 3076 28245 3084 28279
rect 3032 28238 3084 28245
rect 3225 28279 3277 28289
rect 3225 28245 3234 28279
rect 3234 28245 3268 28279
rect 3268 28245 3277 28279
rect 3225 28237 3277 28245
rect 3417 28279 3469 28289
rect 3417 28245 3426 28279
rect 3426 28245 3460 28279
rect 3460 28245 3469 28279
rect 3417 28237 3469 28245
rect 3978 28279 4030 28290
rect 3978 28245 3987 28279
rect 3987 28245 4021 28279
rect 4021 28245 4030 28279
rect 3978 28238 4030 28245
rect 4169 28279 4221 28290
rect 4169 28245 4179 28279
rect 4179 28245 4213 28279
rect 4213 28245 4221 28279
rect 4169 28238 4221 28245
rect 4361 28279 4413 28290
rect 4361 28245 4371 28279
rect 4371 28245 4405 28279
rect 4405 28245 4413 28279
rect 4361 28238 4413 28245
rect 4553 28279 4605 28290
rect 4553 28245 4563 28279
rect 4563 28245 4597 28279
rect 4597 28245 4605 28279
rect 4553 28238 4605 28245
rect 4746 28279 4798 28289
rect 4746 28245 4755 28279
rect 4755 28245 4789 28279
rect 4789 28245 4798 28279
rect 4746 28237 4798 28245
rect 4938 28279 4990 28289
rect 4938 28245 4947 28279
rect 4947 28245 4981 28279
rect 4981 28245 4990 28279
rect 4938 28237 4990 28245
rect 304 27796 356 27806
rect 304 27762 313 27796
rect 313 27762 347 27796
rect 347 27762 356 27796
rect 304 27754 356 27762
rect 497 27796 549 27806
rect 497 27762 505 27796
rect 505 27762 539 27796
rect 539 27762 549 27796
rect 497 27754 549 27762
rect 688 27796 740 27806
rect 688 27762 697 27796
rect 697 27762 731 27796
rect 731 27762 740 27796
rect 688 27754 740 27762
rect 880 27796 932 27806
rect 880 27762 889 27796
rect 889 27762 923 27796
rect 923 27762 932 27796
rect 880 27754 932 27762
rect 1072 27796 1124 27806
rect 1072 27762 1081 27796
rect 1081 27762 1115 27796
rect 1115 27762 1124 27796
rect 1072 27754 1124 27762
rect 1264 27796 1316 27806
rect 1264 27762 1273 27796
rect 1273 27762 1307 27796
rect 1307 27762 1316 27796
rect 1264 27754 1316 27762
rect 1522 27747 1578 27807
rect 1792 27747 1852 27807
rect 2056 27400 2190 27508
rect 2457 27800 2509 27810
rect 2457 27766 2466 27800
rect 2466 27766 2500 27800
rect 2500 27766 2509 27800
rect 2457 27758 2509 27766
rect 2650 27800 2702 27810
rect 2650 27766 2658 27800
rect 2658 27766 2692 27800
rect 2692 27766 2702 27800
rect 2650 27758 2702 27766
rect 2841 27800 2893 27810
rect 2841 27766 2850 27800
rect 2850 27766 2884 27800
rect 2884 27766 2893 27800
rect 2841 27758 2893 27766
rect 3033 27800 3085 27810
rect 3033 27766 3042 27800
rect 3042 27766 3076 27800
rect 3076 27766 3085 27800
rect 3033 27758 3085 27766
rect 3225 27800 3277 27810
rect 3225 27766 3234 27800
rect 3234 27766 3268 27800
rect 3268 27766 3277 27800
rect 3225 27758 3277 27766
rect 3417 27800 3469 27810
rect 3417 27766 3426 27800
rect 3426 27766 3460 27800
rect 3460 27766 3469 27800
rect 3417 27758 3469 27766
rect 1608 27040 1720 27164
rect 304 26988 356 26999
rect 304 26954 313 26988
rect 313 26954 347 26988
rect 347 26954 356 26988
rect 304 26947 356 26954
rect 495 26988 547 26999
rect 495 26954 505 26988
rect 505 26954 539 26988
rect 539 26954 547 26988
rect 495 26947 547 26954
rect 687 26988 739 26999
rect 687 26954 697 26988
rect 697 26954 731 26988
rect 731 26954 739 26988
rect 687 26947 739 26954
rect 879 26988 931 26999
rect 879 26954 889 26988
rect 889 26954 923 26988
rect 923 26954 931 26988
rect 879 26947 931 26954
rect 1072 26988 1124 26998
rect 1072 26954 1081 26988
rect 1081 26954 1115 26988
rect 1115 26954 1124 26988
rect 1072 26946 1124 26954
rect 1264 26988 1316 26998
rect 1264 26954 1273 26988
rect 1273 26954 1307 26988
rect 1307 26954 1316 26988
rect 1264 26946 1316 26954
rect 1468 26946 1524 27002
rect 1930 26948 1986 27004
rect 3978 27800 4030 27810
rect 3978 27766 3987 27800
rect 3987 27766 4021 27800
rect 4021 27766 4030 27800
rect 3978 27758 4030 27766
rect 4171 27800 4223 27810
rect 4171 27766 4179 27800
rect 4179 27766 4213 27800
rect 4213 27766 4223 27800
rect 4171 27758 4223 27766
rect 4362 27800 4414 27810
rect 4362 27766 4371 27800
rect 4371 27766 4405 27800
rect 4405 27766 4414 27800
rect 4362 27758 4414 27766
rect 4554 27800 4606 27810
rect 4554 27766 4563 27800
rect 4563 27766 4597 27800
rect 4597 27766 4606 27800
rect 4554 27758 4606 27766
rect 4746 27800 4798 27810
rect 4746 27766 4755 27800
rect 4755 27766 4789 27800
rect 4789 27766 4798 27800
rect 4746 27758 4798 27766
rect 4938 27800 4990 27810
rect 4938 27766 4947 27800
rect 4947 27766 4981 27800
rect 4981 27766 4990 27800
rect 4938 27758 4990 27766
rect 3681 27214 3733 27233
rect 3681 27181 3691 27214
rect 3691 27181 3725 27214
rect 3725 27181 3733 27214
rect 5337 27255 5389 27265
rect 5337 27221 5348 27255
rect 5348 27221 5382 27255
rect 5382 27221 5389 27255
rect 5337 27213 5389 27221
rect 5449 27260 5501 27267
rect 5449 27226 5450 27260
rect 5450 27226 5484 27260
rect 5484 27226 5501 27260
rect 5449 27215 5501 27226
rect 2457 26992 2509 27003
rect 2457 26958 2466 26992
rect 2466 26958 2500 26992
rect 2500 26958 2509 26992
rect 2457 26951 2509 26958
rect 2648 26992 2700 27003
rect 2648 26958 2658 26992
rect 2658 26958 2692 26992
rect 2692 26958 2700 26992
rect 2648 26951 2700 26958
rect 2840 26992 2892 27003
rect 2840 26958 2850 26992
rect 2850 26958 2884 26992
rect 2884 26958 2892 26992
rect 2840 26951 2892 26958
rect 3032 26992 3084 27003
rect 3032 26958 3042 26992
rect 3042 26958 3076 26992
rect 3076 26958 3084 26992
rect 3032 26951 3084 26958
rect 3225 26992 3277 27002
rect 3225 26958 3234 26992
rect 3234 26958 3268 26992
rect 3268 26958 3277 26992
rect 3225 26950 3277 26958
rect 3417 26992 3469 27002
rect 3417 26958 3426 26992
rect 3426 26958 3460 26992
rect 3460 26958 3469 26992
rect 3417 26950 3469 26958
rect 3978 26992 4030 27003
rect 3978 26958 3987 26992
rect 3987 26958 4021 26992
rect 4021 26958 4030 26992
rect 3978 26951 4030 26958
rect 4169 26992 4221 27003
rect 4169 26958 4179 26992
rect 4179 26958 4213 26992
rect 4213 26958 4221 26992
rect 4169 26951 4221 26958
rect 4361 26992 4413 27003
rect 4361 26958 4371 26992
rect 4371 26958 4405 26992
rect 4405 26958 4413 26992
rect 4361 26951 4413 26958
rect 4553 26992 4605 27003
rect 4553 26958 4563 26992
rect 4563 26958 4597 26992
rect 4597 26958 4605 26992
rect 4553 26951 4605 26958
rect 4746 26992 4798 27002
rect 4746 26958 4755 26992
rect 4755 26958 4789 26992
rect 4789 26958 4798 26992
rect 4746 26950 4798 26958
rect 4938 26992 4990 27002
rect 4938 26958 4947 26992
rect 4947 26958 4981 26992
rect 4981 26958 4990 26992
rect 4938 26950 4990 26958
rect 304 26509 356 26519
rect 304 26475 313 26509
rect 313 26475 347 26509
rect 347 26475 356 26509
rect 304 26467 356 26475
rect 497 26509 549 26519
rect 497 26475 505 26509
rect 505 26475 539 26509
rect 539 26475 549 26509
rect 497 26467 549 26475
rect 688 26509 740 26519
rect 688 26475 697 26509
rect 697 26475 731 26509
rect 731 26475 740 26509
rect 688 26467 740 26475
rect 880 26509 932 26519
rect 880 26475 889 26509
rect 889 26475 923 26509
rect 923 26475 932 26509
rect 880 26467 932 26475
rect 1072 26509 1124 26519
rect 1072 26475 1081 26509
rect 1081 26475 1115 26509
rect 1115 26475 1124 26509
rect 1072 26467 1124 26475
rect 1264 26509 1316 26519
rect 1264 26475 1273 26509
rect 1273 26475 1307 26509
rect 1307 26475 1316 26509
rect 1264 26467 1316 26475
rect 1522 26460 1578 26520
rect 1792 26460 1852 26520
rect 2056 26113 2190 26221
rect 2457 26513 2509 26523
rect 2457 26479 2466 26513
rect 2466 26479 2500 26513
rect 2500 26479 2509 26513
rect 2457 26471 2509 26479
rect 2650 26513 2702 26523
rect 2650 26479 2658 26513
rect 2658 26479 2692 26513
rect 2692 26479 2702 26513
rect 2650 26471 2702 26479
rect 2841 26513 2893 26523
rect 2841 26479 2850 26513
rect 2850 26479 2884 26513
rect 2884 26479 2893 26513
rect 2841 26471 2893 26479
rect 3033 26513 3085 26523
rect 3033 26479 3042 26513
rect 3042 26479 3076 26513
rect 3076 26479 3085 26513
rect 3033 26471 3085 26479
rect 3225 26513 3277 26523
rect 3225 26479 3234 26513
rect 3234 26479 3268 26513
rect 3268 26479 3277 26513
rect 3225 26471 3277 26479
rect 3417 26513 3469 26523
rect 3417 26479 3426 26513
rect 3426 26479 3460 26513
rect 3460 26479 3469 26513
rect 3417 26471 3469 26479
rect 1608 25753 1720 25877
rect 304 25701 356 25712
rect 304 25667 313 25701
rect 313 25667 347 25701
rect 347 25667 356 25701
rect 304 25660 356 25667
rect 495 25701 547 25712
rect 495 25667 505 25701
rect 505 25667 539 25701
rect 539 25667 547 25701
rect 495 25660 547 25667
rect 687 25701 739 25712
rect 687 25667 697 25701
rect 697 25667 731 25701
rect 731 25667 739 25701
rect 687 25660 739 25667
rect 879 25701 931 25712
rect 879 25667 889 25701
rect 889 25667 923 25701
rect 923 25667 931 25701
rect 879 25660 931 25667
rect 1072 25701 1124 25711
rect 1072 25667 1081 25701
rect 1081 25667 1115 25701
rect 1115 25667 1124 25701
rect 1072 25659 1124 25667
rect 1264 25701 1316 25711
rect 1264 25667 1273 25701
rect 1273 25667 1307 25701
rect 1307 25667 1316 25701
rect 1264 25659 1316 25667
rect 1468 25659 1524 25715
rect 1930 25661 1986 25717
rect 3978 26513 4030 26523
rect 3978 26479 3987 26513
rect 3987 26479 4021 26513
rect 4021 26479 4030 26513
rect 3978 26471 4030 26479
rect 4171 26513 4223 26523
rect 4171 26479 4179 26513
rect 4179 26479 4213 26513
rect 4213 26479 4223 26513
rect 4171 26471 4223 26479
rect 4362 26513 4414 26523
rect 4362 26479 4371 26513
rect 4371 26479 4405 26513
rect 4405 26479 4414 26513
rect 4362 26471 4414 26479
rect 4554 26513 4606 26523
rect 4554 26479 4563 26513
rect 4563 26479 4597 26513
rect 4597 26479 4606 26513
rect 4554 26471 4606 26479
rect 4746 26513 4798 26523
rect 4746 26479 4755 26513
rect 4755 26479 4789 26513
rect 4789 26479 4798 26513
rect 4746 26471 4798 26479
rect 4938 26513 4990 26523
rect 4938 26479 4947 26513
rect 4947 26479 4981 26513
rect 4981 26479 4990 26513
rect 4938 26471 4990 26479
rect 3681 25927 3733 25946
rect 3681 25894 3691 25927
rect 3691 25894 3725 25927
rect 3725 25894 3733 25927
rect 5337 25968 5389 25978
rect 5337 25934 5348 25968
rect 5348 25934 5382 25968
rect 5382 25934 5389 25968
rect 5337 25926 5389 25934
rect 5449 25973 5501 25980
rect 5449 25939 5450 25973
rect 5450 25939 5484 25973
rect 5484 25939 5501 25973
rect 5449 25928 5501 25939
rect 2457 25705 2509 25716
rect 2457 25671 2466 25705
rect 2466 25671 2500 25705
rect 2500 25671 2509 25705
rect 2457 25664 2509 25671
rect 2648 25705 2700 25716
rect 2648 25671 2658 25705
rect 2658 25671 2692 25705
rect 2692 25671 2700 25705
rect 2648 25664 2700 25671
rect 2840 25705 2892 25716
rect 2840 25671 2850 25705
rect 2850 25671 2884 25705
rect 2884 25671 2892 25705
rect 2840 25664 2892 25671
rect 3032 25705 3084 25716
rect 3032 25671 3042 25705
rect 3042 25671 3076 25705
rect 3076 25671 3084 25705
rect 3032 25664 3084 25671
rect 3225 25705 3277 25715
rect 3225 25671 3234 25705
rect 3234 25671 3268 25705
rect 3268 25671 3277 25705
rect 3225 25663 3277 25671
rect 3417 25705 3469 25715
rect 3417 25671 3426 25705
rect 3426 25671 3460 25705
rect 3460 25671 3469 25705
rect 3417 25663 3469 25671
rect 3978 25705 4030 25716
rect 3978 25671 3987 25705
rect 3987 25671 4021 25705
rect 4021 25671 4030 25705
rect 3978 25664 4030 25671
rect 4169 25705 4221 25716
rect 4169 25671 4179 25705
rect 4179 25671 4213 25705
rect 4213 25671 4221 25705
rect 4169 25664 4221 25671
rect 4361 25705 4413 25716
rect 4361 25671 4371 25705
rect 4371 25671 4405 25705
rect 4405 25671 4413 25705
rect 4361 25664 4413 25671
rect 4553 25705 4605 25716
rect 4553 25671 4563 25705
rect 4563 25671 4597 25705
rect 4597 25671 4605 25705
rect 4553 25664 4605 25671
rect 4746 25705 4798 25715
rect 4746 25671 4755 25705
rect 4755 25671 4789 25705
rect 4789 25671 4798 25705
rect 4746 25663 4798 25671
rect 4938 25705 4990 25715
rect 4938 25671 4947 25705
rect 4947 25671 4981 25705
rect 4981 25671 4990 25705
rect 4938 25663 4990 25671
rect 304 25222 356 25232
rect 304 25188 313 25222
rect 313 25188 347 25222
rect 347 25188 356 25222
rect 304 25180 356 25188
rect 497 25222 549 25232
rect 497 25188 505 25222
rect 505 25188 539 25222
rect 539 25188 549 25222
rect 497 25180 549 25188
rect 688 25222 740 25232
rect 688 25188 697 25222
rect 697 25188 731 25222
rect 731 25188 740 25222
rect 688 25180 740 25188
rect 880 25222 932 25232
rect 880 25188 889 25222
rect 889 25188 923 25222
rect 923 25188 932 25222
rect 880 25180 932 25188
rect 1072 25222 1124 25232
rect 1072 25188 1081 25222
rect 1081 25188 1115 25222
rect 1115 25188 1124 25222
rect 1072 25180 1124 25188
rect 1264 25222 1316 25232
rect 1264 25188 1273 25222
rect 1273 25188 1307 25222
rect 1307 25188 1316 25222
rect 1264 25180 1316 25188
rect 1522 25173 1578 25233
rect 1792 25173 1852 25233
rect 2056 24826 2190 24934
rect 2457 25226 2509 25236
rect 2457 25192 2466 25226
rect 2466 25192 2500 25226
rect 2500 25192 2509 25226
rect 2457 25184 2509 25192
rect 2650 25226 2702 25236
rect 2650 25192 2658 25226
rect 2658 25192 2692 25226
rect 2692 25192 2702 25226
rect 2650 25184 2702 25192
rect 2841 25226 2893 25236
rect 2841 25192 2850 25226
rect 2850 25192 2884 25226
rect 2884 25192 2893 25226
rect 2841 25184 2893 25192
rect 3033 25226 3085 25236
rect 3033 25192 3042 25226
rect 3042 25192 3076 25226
rect 3076 25192 3085 25226
rect 3033 25184 3085 25192
rect 3225 25226 3277 25236
rect 3225 25192 3234 25226
rect 3234 25192 3268 25226
rect 3268 25192 3277 25226
rect 3225 25184 3277 25192
rect 3417 25226 3469 25236
rect 3417 25192 3426 25226
rect 3426 25192 3460 25226
rect 3460 25192 3469 25226
rect 3417 25184 3469 25192
rect 1608 24466 1720 24590
rect 304 24414 356 24425
rect 304 24380 313 24414
rect 313 24380 347 24414
rect 347 24380 356 24414
rect 304 24373 356 24380
rect 495 24414 547 24425
rect 495 24380 505 24414
rect 505 24380 539 24414
rect 539 24380 547 24414
rect 495 24373 547 24380
rect 687 24414 739 24425
rect 687 24380 697 24414
rect 697 24380 731 24414
rect 731 24380 739 24414
rect 687 24373 739 24380
rect 879 24414 931 24425
rect 879 24380 889 24414
rect 889 24380 923 24414
rect 923 24380 931 24414
rect 879 24373 931 24380
rect 1072 24414 1124 24424
rect 1072 24380 1081 24414
rect 1081 24380 1115 24414
rect 1115 24380 1124 24414
rect 1072 24372 1124 24380
rect 1264 24414 1316 24424
rect 1264 24380 1273 24414
rect 1273 24380 1307 24414
rect 1307 24380 1316 24414
rect 1264 24372 1316 24380
rect 1468 24372 1524 24428
rect 1930 24374 1986 24430
rect 3978 25226 4030 25236
rect 3978 25192 3987 25226
rect 3987 25192 4021 25226
rect 4021 25192 4030 25226
rect 3978 25184 4030 25192
rect 4171 25226 4223 25236
rect 4171 25192 4179 25226
rect 4179 25192 4213 25226
rect 4213 25192 4223 25226
rect 4171 25184 4223 25192
rect 4362 25226 4414 25236
rect 4362 25192 4371 25226
rect 4371 25192 4405 25226
rect 4405 25192 4414 25226
rect 4362 25184 4414 25192
rect 4554 25226 4606 25236
rect 4554 25192 4563 25226
rect 4563 25192 4597 25226
rect 4597 25192 4606 25226
rect 4554 25184 4606 25192
rect 4746 25226 4798 25236
rect 4746 25192 4755 25226
rect 4755 25192 4789 25226
rect 4789 25192 4798 25226
rect 4746 25184 4798 25192
rect 4938 25226 4990 25236
rect 4938 25192 4947 25226
rect 4947 25192 4981 25226
rect 4981 25192 4990 25226
rect 4938 25184 4990 25192
rect 3681 24640 3733 24659
rect 3681 24607 3691 24640
rect 3691 24607 3725 24640
rect 3725 24607 3733 24640
rect 5337 24681 5389 24691
rect 5337 24647 5348 24681
rect 5348 24647 5382 24681
rect 5382 24647 5389 24681
rect 5337 24639 5389 24647
rect 5449 24686 5501 24693
rect 5449 24652 5450 24686
rect 5450 24652 5484 24686
rect 5484 24652 5501 24686
rect 5449 24641 5501 24652
rect 2457 24418 2509 24429
rect 2457 24384 2466 24418
rect 2466 24384 2500 24418
rect 2500 24384 2509 24418
rect 2457 24377 2509 24384
rect 2648 24418 2700 24429
rect 2648 24384 2658 24418
rect 2658 24384 2692 24418
rect 2692 24384 2700 24418
rect 2648 24377 2700 24384
rect 2840 24418 2892 24429
rect 2840 24384 2850 24418
rect 2850 24384 2884 24418
rect 2884 24384 2892 24418
rect 2840 24377 2892 24384
rect 3032 24418 3084 24429
rect 3032 24384 3042 24418
rect 3042 24384 3076 24418
rect 3076 24384 3084 24418
rect 3032 24377 3084 24384
rect 3225 24418 3277 24428
rect 3225 24384 3234 24418
rect 3234 24384 3268 24418
rect 3268 24384 3277 24418
rect 3225 24376 3277 24384
rect 3417 24418 3469 24428
rect 3417 24384 3426 24418
rect 3426 24384 3460 24418
rect 3460 24384 3469 24418
rect 3417 24376 3469 24384
rect 3978 24418 4030 24429
rect 3978 24384 3987 24418
rect 3987 24384 4021 24418
rect 4021 24384 4030 24418
rect 3978 24377 4030 24384
rect 4169 24418 4221 24429
rect 4169 24384 4179 24418
rect 4179 24384 4213 24418
rect 4213 24384 4221 24418
rect 4169 24377 4221 24384
rect 4361 24418 4413 24429
rect 4361 24384 4371 24418
rect 4371 24384 4405 24418
rect 4405 24384 4413 24418
rect 4361 24377 4413 24384
rect 4553 24418 4605 24429
rect 4553 24384 4563 24418
rect 4563 24384 4597 24418
rect 4597 24384 4605 24418
rect 4553 24377 4605 24384
rect 4746 24418 4798 24428
rect 4746 24384 4755 24418
rect 4755 24384 4789 24418
rect 4789 24384 4798 24418
rect 4746 24376 4798 24384
rect 4938 24418 4990 24428
rect 4938 24384 4947 24418
rect 4947 24384 4981 24418
rect 4981 24384 4990 24418
rect 4938 24376 4990 24384
rect 304 23935 356 23945
rect 304 23901 313 23935
rect 313 23901 347 23935
rect 347 23901 356 23935
rect 304 23893 356 23901
rect 497 23935 549 23945
rect 497 23901 505 23935
rect 505 23901 539 23935
rect 539 23901 549 23935
rect 497 23893 549 23901
rect 688 23935 740 23945
rect 688 23901 697 23935
rect 697 23901 731 23935
rect 731 23901 740 23935
rect 688 23893 740 23901
rect 880 23935 932 23945
rect 880 23901 889 23935
rect 889 23901 923 23935
rect 923 23901 932 23935
rect 880 23893 932 23901
rect 1072 23935 1124 23945
rect 1072 23901 1081 23935
rect 1081 23901 1115 23935
rect 1115 23901 1124 23935
rect 1072 23893 1124 23901
rect 1264 23935 1316 23945
rect 1264 23901 1273 23935
rect 1273 23901 1307 23935
rect 1307 23901 1316 23935
rect 1264 23893 1316 23901
rect 1522 23886 1578 23946
rect 1792 23886 1852 23946
rect 2056 23539 2190 23647
rect 2457 23939 2509 23949
rect 2457 23905 2466 23939
rect 2466 23905 2500 23939
rect 2500 23905 2509 23939
rect 2457 23897 2509 23905
rect 2650 23939 2702 23949
rect 2650 23905 2658 23939
rect 2658 23905 2692 23939
rect 2692 23905 2702 23939
rect 2650 23897 2702 23905
rect 2841 23939 2893 23949
rect 2841 23905 2850 23939
rect 2850 23905 2884 23939
rect 2884 23905 2893 23939
rect 2841 23897 2893 23905
rect 3033 23939 3085 23949
rect 3033 23905 3042 23939
rect 3042 23905 3076 23939
rect 3076 23905 3085 23939
rect 3033 23897 3085 23905
rect 3225 23939 3277 23949
rect 3225 23905 3234 23939
rect 3234 23905 3268 23939
rect 3268 23905 3277 23939
rect 3225 23897 3277 23905
rect 3417 23939 3469 23949
rect 3417 23905 3426 23939
rect 3426 23905 3460 23939
rect 3460 23905 3469 23939
rect 3417 23897 3469 23905
rect 1608 23179 1720 23303
rect 304 23127 356 23138
rect 304 23093 313 23127
rect 313 23093 347 23127
rect 347 23093 356 23127
rect 304 23086 356 23093
rect 495 23127 547 23138
rect 495 23093 505 23127
rect 505 23093 539 23127
rect 539 23093 547 23127
rect 495 23086 547 23093
rect 687 23127 739 23138
rect 687 23093 697 23127
rect 697 23093 731 23127
rect 731 23093 739 23127
rect 687 23086 739 23093
rect 879 23127 931 23138
rect 879 23093 889 23127
rect 889 23093 923 23127
rect 923 23093 931 23127
rect 879 23086 931 23093
rect 1072 23127 1124 23137
rect 1072 23093 1081 23127
rect 1081 23093 1115 23127
rect 1115 23093 1124 23127
rect 1072 23085 1124 23093
rect 1264 23127 1316 23137
rect 1264 23093 1273 23127
rect 1273 23093 1307 23127
rect 1307 23093 1316 23127
rect 1264 23085 1316 23093
rect 1468 23085 1524 23141
rect 1930 23087 1986 23143
rect 3978 23939 4030 23949
rect 3978 23905 3987 23939
rect 3987 23905 4021 23939
rect 4021 23905 4030 23939
rect 3978 23897 4030 23905
rect 4171 23939 4223 23949
rect 4171 23905 4179 23939
rect 4179 23905 4213 23939
rect 4213 23905 4223 23939
rect 4171 23897 4223 23905
rect 4362 23939 4414 23949
rect 4362 23905 4371 23939
rect 4371 23905 4405 23939
rect 4405 23905 4414 23939
rect 4362 23897 4414 23905
rect 4554 23939 4606 23949
rect 4554 23905 4563 23939
rect 4563 23905 4597 23939
rect 4597 23905 4606 23939
rect 4554 23897 4606 23905
rect 4746 23939 4798 23949
rect 4746 23905 4755 23939
rect 4755 23905 4789 23939
rect 4789 23905 4798 23939
rect 4746 23897 4798 23905
rect 4938 23939 4990 23949
rect 4938 23905 4947 23939
rect 4947 23905 4981 23939
rect 4981 23905 4990 23939
rect 4938 23897 4990 23905
rect 3681 23353 3733 23372
rect 3681 23320 3691 23353
rect 3691 23320 3725 23353
rect 3725 23320 3733 23353
rect 5337 23394 5389 23404
rect 5337 23360 5348 23394
rect 5348 23360 5382 23394
rect 5382 23360 5389 23394
rect 5337 23352 5389 23360
rect 5449 23399 5501 23406
rect 5449 23365 5450 23399
rect 5450 23365 5484 23399
rect 5484 23365 5501 23399
rect 5449 23354 5501 23365
rect 2457 23131 2509 23142
rect 2457 23097 2466 23131
rect 2466 23097 2500 23131
rect 2500 23097 2509 23131
rect 2457 23090 2509 23097
rect 2648 23131 2700 23142
rect 2648 23097 2658 23131
rect 2658 23097 2692 23131
rect 2692 23097 2700 23131
rect 2648 23090 2700 23097
rect 2840 23131 2892 23142
rect 2840 23097 2850 23131
rect 2850 23097 2884 23131
rect 2884 23097 2892 23131
rect 2840 23090 2892 23097
rect 3032 23131 3084 23142
rect 3032 23097 3042 23131
rect 3042 23097 3076 23131
rect 3076 23097 3084 23131
rect 3032 23090 3084 23097
rect 3225 23131 3277 23141
rect 3225 23097 3234 23131
rect 3234 23097 3268 23131
rect 3268 23097 3277 23131
rect 3225 23089 3277 23097
rect 3417 23131 3469 23141
rect 3417 23097 3426 23131
rect 3426 23097 3460 23131
rect 3460 23097 3469 23131
rect 3417 23089 3469 23097
rect 3978 23131 4030 23142
rect 3978 23097 3987 23131
rect 3987 23097 4021 23131
rect 4021 23097 4030 23131
rect 3978 23090 4030 23097
rect 4169 23131 4221 23142
rect 4169 23097 4179 23131
rect 4179 23097 4213 23131
rect 4213 23097 4221 23131
rect 4169 23090 4221 23097
rect 4361 23131 4413 23142
rect 4361 23097 4371 23131
rect 4371 23097 4405 23131
rect 4405 23097 4413 23131
rect 4361 23090 4413 23097
rect 4553 23131 4605 23142
rect 4553 23097 4563 23131
rect 4563 23097 4597 23131
rect 4597 23097 4605 23131
rect 4553 23090 4605 23097
rect 4746 23131 4798 23141
rect 4746 23097 4755 23131
rect 4755 23097 4789 23131
rect 4789 23097 4798 23131
rect 4746 23089 4798 23097
rect 4938 23131 4990 23141
rect 4938 23097 4947 23131
rect 4947 23097 4981 23131
rect 4981 23097 4990 23131
rect 4938 23089 4990 23097
rect 304 22648 356 22658
rect 304 22614 313 22648
rect 313 22614 347 22648
rect 347 22614 356 22648
rect 304 22606 356 22614
rect 497 22648 549 22658
rect 497 22614 505 22648
rect 505 22614 539 22648
rect 539 22614 549 22648
rect 497 22606 549 22614
rect 688 22648 740 22658
rect 688 22614 697 22648
rect 697 22614 731 22648
rect 731 22614 740 22648
rect 688 22606 740 22614
rect 880 22648 932 22658
rect 880 22614 889 22648
rect 889 22614 923 22648
rect 923 22614 932 22648
rect 880 22606 932 22614
rect 1072 22648 1124 22658
rect 1072 22614 1081 22648
rect 1081 22614 1115 22648
rect 1115 22614 1124 22648
rect 1072 22606 1124 22614
rect 1264 22648 1316 22658
rect 1264 22614 1273 22648
rect 1273 22614 1307 22648
rect 1307 22614 1316 22648
rect 1264 22606 1316 22614
rect 1522 22599 1578 22659
rect 1792 22599 1852 22659
rect 2056 22252 2190 22360
rect 2457 22652 2509 22662
rect 2457 22618 2466 22652
rect 2466 22618 2500 22652
rect 2500 22618 2509 22652
rect 2457 22610 2509 22618
rect 2650 22652 2702 22662
rect 2650 22618 2658 22652
rect 2658 22618 2692 22652
rect 2692 22618 2702 22652
rect 2650 22610 2702 22618
rect 2841 22652 2893 22662
rect 2841 22618 2850 22652
rect 2850 22618 2884 22652
rect 2884 22618 2893 22652
rect 2841 22610 2893 22618
rect 3033 22652 3085 22662
rect 3033 22618 3042 22652
rect 3042 22618 3076 22652
rect 3076 22618 3085 22652
rect 3033 22610 3085 22618
rect 3225 22652 3277 22662
rect 3225 22618 3234 22652
rect 3234 22618 3268 22652
rect 3268 22618 3277 22652
rect 3225 22610 3277 22618
rect 3417 22652 3469 22662
rect 3417 22618 3426 22652
rect 3426 22618 3460 22652
rect 3460 22618 3469 22652
rect 3417 22610 3469 22618
rect 1608 21892 1720 22016
rect 304 21840 356 21851
rect 304 21806 313 21840
rect 313 21806 347 21840
rect 347 21806 356 21840
rect 304 21799 356 21806
rect 495 21840 547 21851
rect 495 21806 505 21840
rect 505 21806 539 21840
rect 539 21806 547 21840
rect 495 21799 547 21806
rect 687 21840 739 21851
rect 687 21806 697 21840
rect 697 21806 731 21840
rect 731 21806 739 21840
rect 687 21799 739 21806
rect 879 21840 931 21851
rect 879 21806 889 21840
rect 889 21806 923 21840
rect 923 21806 931 21840
rect 879 21799 931 21806
rect 1072 21840 1124 21850
rect 1072 21806 1081 21840
rect 1081 21806 1115 21840
rect 1115 21806 1124 21840
rect 1072 21798 1124 21806
rect 1264 21840 1316 21850
rect 1264 21806 1273 21840
rect 1273 21806 1307 21840
rect 1307 21806 1316 21840
rect 1264 21798 1316 21806
rect 1468 21798 1524 21854
rect 1930 21800 1986 21856
rect 3978 22652 4030 22662
rect 3978 22618 3987 22652
rect 3987 22618 4021 22652
rect 4021 22618 4030 22652
rect 3978 22610 4030 22618
rect 4171 22652 4223 22662
rect 4171 22618 4179 22652
rect 4179 22618 4213 22652
rect 4213 22618 4223 22652
rect 4171 22610 4223 22618
rect 4362 22652 4414 22662
rect 4362 22618 4371 22652
rect 4371 22618 4405 22652
rect 4405 22618 4414 22652
rect 4362 22610 4414 22618
rect 4554 22652 4606 22662
rect 4554 22618 4563 22652
rect 4563 22618 4597 22652
rect 4597 22618 4606 22652
rect 4554 22610 4606 22618
rect 4746 22652 4798 22662
rect 4746 22618 4755 22652
rect 4755 22618 4789 22652
rect 4789 22618 4798 22652
rect 4746 22610 4798 22618
rect 4938 22652 4990 22662
rect 4938 22618 4947 22652
rect 4947 22618 4981 22652
rect 4981 22618 4990 22652
rect 4938 22610 4990 22618
rect 3681 22066 3733 22085
rect 3681 22033 3691 22066
rect 3691 22033 3725 22066
rect 3725 22033 3733 22066
rect 5337 22107 5389 22117
rect 5337 22073 5348 22107
rect 5348 22073 5382 22107
rect 5382 22073 5389 22107
rect 5337 22065 5389 22073
rect 5449 22112 5501 22119
rect 5449 22078 5450 22112
rect 5450 22078 5484 22112
rect 5484 22078 5501 22112
rect 5449 22067 5501 22078
rect 2457 21844 2509 21855
rect 2457 21810 2466 21844
rect 2466 21810 2500 21844
rect 2500 21810 2509 21844
rect 2457 21803 2509 21810
rect 2648 21844 2700 21855
rect 2648 21810 2658 21844
rect 2658 21810 2692 21844
rect 2692 21810 2700 21844
rect 2648 21803 2700 21810
rect 2840 21844 2892 21855
rect 2840 21810 2850 21844
rect 2850 21810 2884 21844
rect 2884 21810 2892 21844
rect 2840 21803 2892 21810
rect 3032 21844 3084 21855
rect 3032 21810 3042 21844
rect 3042 21810 3076 21844
rect 3076 21810 3084 21844
rect 3032 21803 3084 21810
rect 3225 21844 3277 21854
rect 3225 21810 3234 21844
rect 3234 21810 3268 21844
rect 3268 21810 3277 21844
rect 3225 21802 3277 21810
rect 3417 21844 3469 21854
rect 3417 21810 3426 21844
rect 3426 21810 3460 21844
rect 3460 21810 3469 21844
rect 3417 21802 3469 21810
rect 3978 21844 4030 21855
rect 3978 21810 3987 21844
rect 3987 21810 4021 21844
rect 4021 21810 4030 21844
rect 3978 21803 4030 21810
rect 4169 21844 4221 21855
rect 4169 21810 4179 21844
rect 4179 21810 4213 21844
rect 4213 21810 4221 21844
rect 4169 21803 4221 21810
rect 4361 21844 4413 21855
rect 4361 21810 4371 21844
rect 4371 21810 4405 21844
rect 4405 21810 4413 21844
rect 4361 21803 4413 21810
rect 4553 21844 4605 21855
rect 4553 21810 4563 21844
rect 4563 21810 4597 21844
rect 4597 21810 4605 21844
rect 4553 21803 4605 21810
rect 4746 21844 4798 21854
rect 4746 21810 4755 21844
rect 4755 21810 4789 21844
rect 4789 21810 4798 21844
rect 4746 21802 4798 21810
rect 4938 21844 4990 21854
rect 4938 21810 4947 21844
rect 4947 21810 4981 21844
rect 4981 21810 4990 21844
rect 4938 21802 4990 21810
rect 304 21361 356 21371
rect 304 21327 313 21361
rect 313 21327 347 21361
rect 347 21327 356 21361
rect 304 21319 356 21327
rect 497 21361 549 21371
rect 497 21327 505 21361
rect 505 21327 539 21361
rect 539 21327 549 21361
rect 497 21319 549 21327
rect 688 21361 740 21371
rect 688 21327 697 21361
rect 697 21327 731 21361
rect 731 21327 740 21361
rect 688 21319 740 21327
rect 880 21361 932 21371
rect 880 21327 889 21361
rect 889 21327 923 21361
rect 923 21327 932 21361
rect 880 21319 932 21327
rect 1072 21361 1124 21371
rect 1072 21327 1081 21361
rect 1081 21327 1115 21361
rect 1115 21327 1124 21361
rect 1072 21319 1124 21327
rect 1264 21361 1316 21371
rect 1264 21327 1273 21361
rect 1273 21327 1307 21361
rect 1307 21327 1316 21361
rect 1264 21319 1316 21327
rect 1522 21312 1578 21372
rect 1792 21312 1852 21372
rect 2056 20965 2190 21073
rect 2457 21365 2509 21375
rect 2457 21331 2466 21365
rect 2466 21331 2500 21365
rect 2500 21331 2509 21365
rect 2457 21323 2509 21331
rect 2650 21365 2702 21375
rect 2650 21331 2658 21365
rect 2658 21331 2692 21365
rect 2692 21331 2702 21365
rect 2650 21323 2702 21331
rect 2841 21365 2893 21375
rect 2841 21331 2850 21365
rect 2850 21331 2884 21365
rect 2884 21331 2893 21365
rect 2841 21323 2893 21331
rect 3033 21365 3085 21375
rect 3033 21331 3042 21365
rect 3042 21331 3076 21365
rect 3076 21331 3085 21365
rect 3033 21323 3085 21331
rect 3225 21365 3277 21375
rect 3225 21331 3234 21365
rect 3234 21331 3268 21365
rect 3268 21331 3277 21365
rect 3225 21323 3277 21331
rect 3417 21365 3469 21375
rect 3417 21331 3426 21365
rect 3426 21331 3460 21365
rect 3460 21331 3469 21365
rect 3417 21323 3469 21331
rect 1608 20605 1720 20729
rect 304 20553 356 20564
rect 304 20519 313 20553
rect 313 20519 347 20553
rect 347 20519 356 20553
rect 304 20512 356 20519
rect 495 20553 547 20564
rect 495 20519 505 20553
rect 505 20519 539 20553
rect 539 20519 547 20553
rect 495 20512 547 20519
rect 687 20553 739 20564
rect 687 20519 697 20553
rect 697 20519 731 20553
rect 731 20519 739 20553
rect 687 20512 739 20519
rect 879 20553 931 20564
rect 879 20519 889 20553
rect 889 20519 923 20553
rect 923 20519 931 20553
rect 879 20512 931 20519
rect 1072 20553 1124 20563
rect 1072 20519 1081 20553
rect 1081 20519 1115 20553
rect 1115 20519 1124 20553
rect 1072 20511 1124 20519
rect 1264 20553 1316 20563
rect 1264 20519 1273 20553
rect 1273 20519 1307 20553
rect 1307 20519 1316 20553
rect 1264 20511 1316 20519
rect 1468 20511 1524 20567
rect 1930 20513 1986 20569
rect 3978 21365 4030 21375
rect 3978 21331 3987 21365
rect 3987 21331 4021 21365
rect 4021 21331 4030 21365
rect 3978 21323 4030 21331
rect 4171 21365 4223 21375
rect 4171 21331 4179 21365
rect 4179 21331 4213 21365
rect 4213 21331 4223 21365
rect 4171 21323 4223 21331
rect 4362 21365 4414 21375
rect 4362 21331 4371 21365
rect 4371 21331 4405 21365
rect 4405 21331 4414 21365
rect 4362 21323 4414 21331
rect 4554 21365 4606 21375
rect 4554 21331 4563 21365
rect 4563 21331 4597 21365
rect 4597 21331 4606 21365
rect 4554 21323 4606 21331
rect 4746 21365 4798 21375
rect 4746 21331 4755 21365
rect 4755 21331 4789 21365
rect 4789 21331 4798 21365
rect 4746 21323 4798 21331
rect 4938 21365 4990 21375
rect 4938 21331 4947 21365
rect 4947 21331 4981 21365
rect 4981 21331 4990 21365
rect 4938 21323 4990 21331
rect 3681 20779 3733 20798
rect 3681 20746 3691 20779
rect 3691 20746 3725 20779
rect 3725 20746 3733 20779
rect 5337 20820 5389 20830
rect 5337 20786 5348 20820
rect 5348 20786 5382 20820
rect 5382 20786 5389 20820
rect 5337 20778 5389 20786
rect 5449 20825 5501 20832
rect 5449 20791 5450 20825
rect 5450 20791 5484 20825
rect 5484 20791 5501 20825
rect 5449 20780 5501 20791
rect 2457 20557 2509 20568
rect 2457 20523 2466 20557
rect 2466 20523 2500 20557
rect 2500 20523 2509 20557
rect 2457 20516 2509 20523
rect 2648 20557 2700 20568
rect 2648 20523 2658 20557
rect 2658 20523 2692 20557
rect 2692 20523 2700 20557
rect 2648 20516 2700 20523
rect 2840 20557 2892 20568
rect 2840 20523 2850 20557
rect 2850 20523 2884 20557
rect 2884 20523 2892 20557
rect 2840 20516 2892 20523
rect 3032 20557 3084 20568
rect 3032 20523 3042 20557
rect 3042 20523 3076 20557
rect 3076 20523 3084 20557
rect 3032 20516 3084 20523
rect 3225 20557 3277 20567
rect 3225 20523 3234 20557
rect 3234 20523 3268 20557
rect 3268 20523 3277 20557
rect 3225 20515 3277 20523
rect 3417 20557 3469 20567
rect 3417 20523 3426 20557
rect 3426 20523 3460 20557
rect 3460 20523 3469 20557
rect 3417 20515 3469 20523
rect 3978 20557 4030 20568
rect 3978 20523 3987 20557
rect 3987 20523 4021 20557
rect 4021 20523 4030 20557
rect 3978 20516 4030 20523
rect 4169 20557 4221 20568
rect 4169 20523 4179 20557
rect 4179 20523 4213 20557
rect 4213 20523 4221 20557
rect 4169 20516 4221 20523
rect 4361 20557 4413 20568
rect 4361 20523 4371 20557
rect 4371 20523 4405 20557
rect 4405 20523 4413 20557
rect 4361 20516 4413 20523
rect 4553 20557 4605 20568
rect 4553 20523 4563 20557
rect 4563 20523 4597 20557
rect 4597 20523 4605 20557
rect 4553 20516 4605 20523
rect 4746 20557 4798 20567
rect 4746 20523 4755 20557
rect 4755 20523 4789 20557
rect 4789 20523 4798 20557
rect 4746 20515 4798 20523
rect 4938 20557 4990 20567
rect 4938 20523 4947 20557
rect 4947 20523 4981 20557
rect 4981 20523 4990 20557
rect 4938 20515 4990 20523
rect 304 20074 356 20084
rect 304 20040 313 20074
rect 313 20040 347 20074
rect 347 20040 356 20074
rect 304 20032 356 20040
rect 497 20074 549 20084
rect 497 20040 505 20074
rect 505 20040 539 20074
rect 539 20040 549 20074
rect 497 20032 549 20040
rect 688 20074 740 20084
rect 688 20040 697 20074
rect 697 20040 731 20074
rect 731 20040 740 20074
rect 688 20032 740 20040
rect 880 20074 932 20084
rect 880 20040 889 20074
rect 889 20040 923 20074
rect 923 20040 932 20074
rect 880 20032 932 20040
rect 1072 20074 1124 20084
rect 1072 20040 1081 20074
rect 1081 20040 1115 20074
rect 1115 20040 1124 20074
rect 1072 20032 1124 20040
rect 1264 20074 1316 20084
rect 1264 20040 1273 20074
rect 1273 20040 1307 20074
rect 1307 20040 1316 20074
rect 1264 20032 1316 20040
rect 1522 20025 1578 20085
rect 1792 20025 1852 20085
rect 2056 19678 2190 19786
rect 2457 20078 2509 20088
rect 2457 20044 2466 20078
rect 2466 20044 2500 20078
rect 2500 20044 2509 20078
rect 2457 20036 2509 20044
rect 2650 20078 2702 20088
rect 2650 20044 2658 20078
rect 2658 20044 2692 20078
rect 2692 20044 2702 20078
rect 2650 20036 2702 20044
rect 2841 20078 2893 20088
rect 2841 20044 2850 20078
rect 2850 20044 2884 20078
rect 2884 20044 2893 20078
rect 2841 20036 2893 20044
rect 3033 20078 3085 20088
rect 3033 20044 3042 20078
rect 3042 20044 3076 20078
rect 3076 20044 3085 20078
rect 3033 20036 3085 20044
rect 3225 20078 3277 20088
rect 3225 20044 3234 20078
rect 3234 20044 3268 20078
rect 3268 20044 3277 20078
rect 3225 20036 3277 20044
rect 3417 20078 3469 20088
rect 3417 20044 3426 20078
rect 3426 20044 3460 20078
rect 3460 20044 3469 20078
rect 3417 20036 3469 20044
rect 1608 19318 1720 19442
rect 304 19266 356 19277
rect 304 19232 313 19266
rect 313 19232 347 19266
rect 347 19232 356 19266
rect 304 19225 356 19232
rect 495 19266 547 19277
rect 495 19232 505 19266
rect 505 19232 539 19266
rect 539 19232 547 19266
rect 495 19225 547 19232
rect 687 19266 739 19277
rect 687 19232 697 19266
rect 697 19232 731 19266
rect 731 19232 739 19266
rect 687 19225 739 19232
rect 879 19266 931 19277
rect 879 19232 889 19266
rect 889 19232 923 19266
rect 923 19232 931 19266
rect 879 19225 931 19232
rect 1072 19266 1124 19276
rect 1072 19232 1081 19266
rect 1081 19232 1115 19266
rect 1115 19232 1124 19266
rect 1072 19224 1124 19232
rect 1264 19266 1316 19276
rect 1264 19232 1273 19266
rect 1273 19232 1307 19266
rect 1307 19232 1316 19266
rect 1264 19224 1316 19232
rect 1468 19224 1524 19280
rect 1930 19226 1986 19282
rect 3978 20078 4030 20088
rect 3978 20044 3987 20078
rect 3987 20044 4021 20078
rect 4021 20044 4030 20078
rect 3978 20036 4030 20044
rect 4171 20078 4223 20088
rect 4171 20044 4179 20078
rect 4179 20044 4213 20078
rect 4213 20044 4223 20078
rect 4171 20036 4223 20044
rect 4362 20078 4414 20088
rect 4362 20044 4371 20078
rect 4371 20044 4405 20078
rect 4405 20044 4414 20078
rect 4362 20036 4414 20044
rect 4554 20078 4606 20088
rect 4554 20044 4563 20078
rect 4563 20044 4597 20078
rect 4597 20044 4606 20078
rect 4554 20036 4606 20044
rect 4746 20078 4798 20088
rect 4746 20044 4755 20078
rect 4755 20044 4789 20078
rect 4789 20044 4798 20078
rect 4746 20036 4798 20044
rect 4938 20078 4990 20088
rect 4938 20044 4947 20078
rect 4947 20044 4981 20078
rect 4981 20044 4990 20078
rect 4938 20036 4990 20044
rect 3681 19492 3733 19511
rect 3681 19459 3691 19492
rect 3691 19459 3725 19492
rect 3725 19459 3733 19492
rect 5337 19533 5389 19543
rect 5337 19499 5348 19533
rect 5348 19499 5382 19533
rect 5382 19499 5389 19533
rect 5337 19491 5389 19499
rect 5449 19538 5501 19545
rect 5449 19504 5450 19538
rect 5450 19504 5484 19538
rect 5484 19504 5501 19538
rect 5449 19493 5501 19504
rect 2457 19270 2509 19281
rect 2457 19236 2466 19270
rect 2466 19236 2500 19270
rect 2500 19236 2509 19270
rect 2457 19229 2509 19236
rect 2648 19270 2700 19281
rect 2648 19236 2658 19270
rect 2658 19236 2692 19270
rect 2692 19236 2700 19270
rect 2648 19229 2700 19236
rect 2840 19270 2892 19281
rect 2840 19236 2850 19270
rect 2850 19236 2884 19270
rect 2884 19236 2892 19270
rect 2840 19229 2892 19236
rect 3032 19270 3084 19281
rect 3032 19236 3042 19270
rect 3042 19236 3076 19270
rect 3076 19236 3084 19270
rect 3032 19229 3084 19236
rect 3225 19270 3277 19280
rect 3225 19236 3234 19270
rect 3234 19236 3268 19270
rect 3268 19236 3277 19270
rect 3225 19228 3277 19236
rect 3417 19270 3469 19280
rect 3417 19236 3426 19270
rect 3426 19236 3460 19270
rect 3460 19236 3469 19270
rect 3417 19228 3469 19236
rect 3978 19270 4030 19281
rect 3978 19236 3987 19270
rect 3987 19236 4021 19270
rect 4021 19236 4030 19270
rect 3978 19229 4030 19236
rect 4169 19270 4221 19281
rect 4169 19236 4179 19270
rect 4179 19236 4213 19270
rect 4213 19236 4221 19270
rect 4169 19229 4221 19236
rect 4361 19270 4413 19281
rect 4361 19236 4371 19270
rect 4371 19236 4405 19270
rect 4405 19236 4413 19270
rect 4361 19229 4413 19236
rect 4553 19270 4605 19281
rect 4553 19236 4563 19270
rect 4563 19236 4597 19270
rect 4597 19236 4605 19270
rect 4553 19229 4605 19236
rect 4746 19270 4798 19280
rect 4746 19236 4755 19270
rect 4755 19236 4789 19270
rect 4789 19236 4798 19270
rect 4746 19228 4798 19236
rect 4938 19270 4990 19280
rect 4938 19236 4947 19270
rect 4947 19236 4981 19270
rect 4981 19236 4990 19270
rect 4938 19228 4990 19236
rect 304 18787 356 18797
rect 304 18753 313 18787
rect 313 18753 347 18787
rect 347 18753 356 18787
rect 304 18745 356 18753
rect 497 18787 549 18797
rect 497 18753 505 18787
rect 505 18753 539 18787
rect 539 18753 549 18787
rect 497 18745 549 18753
rect 688 18787 740 18797
rect 688 18753 697 18787
rect 697 18753 731 18787
rect 731 18753 740 18787
rect 688 18745 740 18753
rect 880 18787 932 18797
rect 880 18753 889 18787
rect 889 18753 923 18787
rect 923 18753 932 18787
rect 880 18745 932 18753
rect 1072 18787 1124 18797
rect 1072 18753 1081 18787
rect 1081 18753 1115 18787
rect 1115 18753 1124 18787
rect 1072 18745 1124 18753
rect 1264 18787 1316 18797
rect 1264 18753 1273 18787
rect 1273 18753 1307 18787
rect 1307 18753 1316 18787
rect 1264 18745 1316 18753
rect 1522 18738 1578 18798
rect 1792 18738 1852 18798
rect 2056 18391 2190 18499
rect 2457 18791 2509 18801
rect 2457 18757 2466 18791
rect 2466 18757 2500 18791
rect 2500 18757 2509 18791
rect 2457 18749 2509 18757
rect 2650 18791 2702 18801
rect 2650 18757 2658 18791
rect 2658 18757 2692 18791
rect 2692 18757 2702 18791
rect 2650 18749 2702 18757
rect 2841 18791 2893 18801
rect 2841 18757 2850 18791
rect 2850 18757 2884 18791
rect 2884 18757 2893 18791
rect 2841 18749 2893 18757
rect 3033 18791 3085 18801
rect 3033 18757 3042 18791
rect 3042 18757 3076 18791
rect 3076 18757 3085 18791
rect 3033 18749 3085 18757
rect 3225 18791 3277 18801
rect 3225 18757 3234 18791
rect 3234 18757 3268 18791
rect 3268 18757 3277 18791
rect 3225 18749 3277 18757
rect 3417 18791 3469 18801
rect 3417 18757 3426 18791
rect 3426 18757 3460 18791
rect 3460 18757 3469 18791
rect 3417 18749 3469 18757
rect 1608 18031 1720 18155
rect 304 17979 356 17990
rect 304 17945 313 17979
rect 313 17945 347 17979
rect 347 17945 356 17979
rect 304 17938 356 17945
rect 495 17979 547 17990
rect 495 17945 505 17979
rect 505 17945 539 17979
rect 539 17945 547 17979
rect 495 17938 547 17945
rect 687 17979 739 17990
rect 687 17945 697 17979
rect 697 17945 731 17979
rect 731 17945 739 17979
rect 687 17938 739 17945
rect 879 17979 931 17990
rect 879 17945 889 17979
rect 889 17945 923 17979
rect 923 17945 931 17979
rect 879 17938 931 17945
rect 1072 17979 1124 17989
rect 1072 17945 1081 17979
rect 1081 17945 1115 17979
rect 1115 17945 1124 17979
rect 1072 17937 1124 17945
rect 1264 17979 1316 17989
rect 1264 17945 1273 17979
rect 1273 17945 1307 17979
rect 1307 17945 1316 17979
rect 1264 17937 1316 17945
rect 1468 17937 1524 17993
rect 1930 17939 1986 17995
rect 3978 18791 4030 18801
rect 3978 18757 3987 18791
rect 3987 18757 4021 18791
rect 4021 18757 4030 18791
rect 3978 18749 4030 18757
rect 4171 18791 4223 18801
rect 4171 18757 4179 18791
rect 4179 18757 4213 18791
rect 4213 18757 4223 18791
rect 4171 18749 4223 18757
rect 4362 18791 4414 18801
rect 4362 18757 4371 18791
rect 4371 18757 4405 18791
rect 4405 18757 4414 18791
rect 4362 18749 4414 18757
rect 4554 18791 4606 18801
rect 4554 18757 4563 18791
rect 4563 18757 4597 18791
rect 4597 18757 4606 18791
rect 4554 18749 4606 18757
rect 4746 18791 4798 18801
rect 4746 18757 4755 18791
rect 4755 18757 4789 18791
rect 4789 18757 4798 18791
rect 4746 18749 4798 18757
rect 4938 18791 4990 18801
rect 4938 18757 4947 18791
rect 4947 18757 4981 18791
rect 4981 18757 4990 18791
rect 4938 18749 4990 18757
rect 3681 18205 3733 18224
rect 3681 18172 3691 18205
rect 3691 18172 3725 18205
rect 3725 18172 3733 18205
rect 5337 18246 5389 18256
rect 5337 18212 5348 18246
rect 5348 18212 5382 18246
rect 5382 18212 5389 18246
rect 5337 18204 5389 18212
rect 5449 18251 5501 18258
rect 5449 18217 5450 18251
rect 5450 18217 5484 18251
rect 5484 18217 5501 18251
rect 5449 18206 5501 18217
rect 2457 17983 2509 17994
rect 2457 17949 2466 17983
rect 2466 17949 2500 17983
rect 2500 17949 2509 17983
rect 2457 17942 2509 17949
rect 2648 17983 2700 17994
rect 2648 17949 2658 17983
rect 2658 17949 2692 17983
rect 2692 17949 2700 17983
rect 2648 17942 2700 17949
rect 2840 17983 2892 17994
rect 2840 17949 2850 17983
rect 2850 17949 2884 17983
rect 2884 17949 2892 17983
rect 2840 17942 2892 17949
rect 3032 17983 3084 17994
rect 3032 17949 3042 17983
rect 3042 17949 3076 17983
rect 3076 17949 3084 17983
rect 3032 17942 3084 17949
rect 3225 17983 3277 17993
rect 3225 17949 3234 17983
rect 3234 17949 3268 17983
rect 3268 17949 3277 17983
rect 3225 17941 3277 17949
rect 3417 17983 3469 17993
rect 3417 17949 3426 17983
rect 3426 17949 3460 17983
rect 3460 17949 3469 17983
rect 3417 17941 3469 17949
rect 3978 17983 4030 17994
rect 3978 17949 3987 17983
rect 3987 17949 4021 17983
rect 4021 17949 4030 17983
rect 3978 17942 4030 17949
rect 4169 17983 4221 17994
rect 4169 17949 4179 17983
rect 4179 17949 4213 17983
rect 4213 17949 4221 17983
rect 4169 17942 4221 17949
rect 4361 17983 4413 17994
rect 4361 17949 4371 17983
rect 4371 17949 4405 17983
rect 4405 17949 4413 17983
rect 4361 17942 4413 17949
rect 4553 17983 4605 17994
rect 4553 17949 4563 17983
rect 4563 17949 4597 17983
rect 4597 17949 4605 17983
rect 4553 17942 4605 17949
rect 4746 17983 4798 17993
rect 4746 17949 4755 17983
rect 4755 17949 4789 17983
rect 4789 17949 4798 17983
rect 4746 17941 4798 17949
rect 4938 17983 4990 17993
rect 4938 17949 4947 17983
rect 4947 17949 4981 17983
rect 4981 17949 4990 17983
rect 4938 17941 4990 17949
rect 304 17500 356 17510
rect 304 17466 313 17500
rect 313 17466 347 17500
rect 347 17466 356 17500
rect 304 17458 356 17466
rect 497 17500 549 17510
rect 497 17466 505 17500
rect 505 17466 539 17500
rect 539 17466 549 17500
rect 497 17458 549 17466
rect 688 17500 740 17510
rect 688 17466 697 17500
rect 697 17466 731 17500
rect 731 17466 740 17500
rect 688 17458 740 17466
rect 880 17500 932 17510
rect 880 17466 889 17500
rect 889 17466 923 17500
rect 923 17466 932 17500
rect 880 17458 932 17466
rect 1072 17500 1124 17510
rect 1072 17466 1081 17500
rect 1081 17466 1115 17500
rect 1115 17466 1124 17500
rect 1072 17458 1124 17466
rect 1264 17500 1316 17510
rect 1264 17466 1273 17500
rect 1273 17466 1307 17500
rect 1307 17466 1316 17500
rect 1264 17458 1316 17466
rect 1522 17451 1578 17511
rect 1792 17451 1852 17511
rect 2056 17104 2190 17212
rect 2457 17504 2509 17514
rect 2457 17470 2466 17504
rect 2466 17470 2500 17504
rect 2500 17470 2509 17504
rect 2457 17462 2509 17470
rect 2650 17504 2702 17514
rect 2650 17470 2658 17504
rect 2658 17470 2692 17504
rect 2692 17470 2702 17504
rect 2650 17462 2702 17470
rect 2841 17504 2893 17514
rect 2841 17470 2850 17504
rect 2850 17470 2884 17504
rect 2884 17470 2893 17504
rect 2841 17462 2893 17470
rect 3033 17504 3085 17514
rect 3033 17470 3042 17504
rect 3042 17470 3076 17504
rect 3076 17470 3085 17504
rect 3033 17462 3085 17470
rect 3225 17504 3277 17514
rect 3225 17470 3234 17504
rect 3234 17470 3268 17504
rect 3268 17470 3277 17504
rect 3225 17462 3277 17470
rect 3417 17504 3469 17514
rect 3417 17470 3426 17504
rect 3426 17470 3460 17504
rect 3460 17470 3469 17504
rect 3417 17462 3469 17470
rect 1608 16744 1720 16868
rect 304 16692 356 16703
rect 304 16658 313 16692
rect 313 16658 347 16692
rect 347 16658 356 16692
rect 304 16651 356 16658
rect 495 16692 547 16703
rect 495 16658 505 16692
rect 505 16658 539 16692
rect 539 16658 547 16692
rect 495 16651 547 16658
rect 687 16692 739 16703
rect 687 16658 697 16692
rect 697 16658 731 16692
rect 731 16658 739 16692
rect 687 16651 739 16658
rect 879 16692 931 16703
rect 879 16658 889 16692
rect 889 16658 923 16692
rect 923 16658 931 16692
rect 879 16651 931 16658
rect 1072 16692 1124 16702
rect 1072 16658 1081 16692
rect 1081 16658 1115 16692
rect 1115 16658 1124 16692
rect 1072 16650 1124 16658
rect 1264 16692 1316 16702
rect 1264 16658 1273 16692
rect 1273 16658 1307 16692
rect 1307 16658 1316 16692
rect 1264 16650 1316 16658
rect 1468 16650 1524 16706
rect 1930 16652 1986 16708
rect 3978 17504 4030 17514
rect 3978 17470 3987 17504
rect 3987 17470 4021 17504
rect 4021 17470 4030 17504
rect 3978 17462 4030 17470
rect 4171 17504 4223 17514
rect 4171 17470 4179 17504
rect 4179 17470 4213 17504
rect 4213 17470 4223 17504
rect 4171 17462 4223 17470
rect 4362 17504 4414 17514
rect 4362 17470 4371 17504
rect 4371 17470 4405 17504
rect 4405 17470 4414 17504
rect 4362 17462 4414 17470
rect 4554 17504 4606 17514
rect 4554 17470 4563 17504
rect 4563 17470 4597 17504
rect 4597 17470 4606 17504
rect 4554 17462 4606 17470
rect 4746 17504 4798 17514
rect 4746 17470 4755 17504
rect 4755 17470 4789 17504
rect 4789 17470 4798 17504
rect 4746 17462 4798 17470
rect 4938 17504 4990 17514
rect 4938 17470 4947 17504
rect 4947 17470 4981 17504
rect 4981 17470 4990 17504
rect 4938 17462 4990 17470
rect 3681 16918 3733 16937
rect 3681 16885 3691 16918
rect 3691 16885 3725 16918
rect 3725 16885 3733 16918
rect 5337 16959 5389 16969
rect 5337 16925 5348 16959
rect 5348 16925 5382 16959
rect 5382 16925 5389 16959
rect 5337 16917 5389 16925
rect 5449 16964 5501 16971
rect 5449 16930 5450 16964
rect 5450 16930 5484 16964
rect 5484 16930 5501 16964
rect 5449 16919 5501 16930
rect 2457 16696 2509 16707
rect 2457 16662 2466 16696
rect 2466 16662 2500 16696
rect 2500 16662 2509 16696
rect 2457 16655 2509 16662
rect 2648 16696 2700 16707
rect 2648 16662 2658 16696
rect 2658 16662 2692 16696
rect 2692 16662 2700 16696
rect 2648 16655 2700 16662
rect 2840 16696 2892 16707
rect 2840 16662 2850 16696
rect 2850 16662 2884 16696
rect 2884 16662 2892 16696
rect 2840 16655 2892 16662
rect 3032 16696 3084 16707
rect 3032 16662 3042 16696
rect 3042 16662 3076 16696
rect 3076 16662 3084 16696
rect 3032 16655 3084 16662
rect 3225 16696 3277 16706
rect 3225 16662 3234 16696
rect 3234 16662 3268 16696
rect 3268 16662 3277 16696
rect 3225 16654 3277 16662
rect 3417 16696 3469 16706
rect 3417 16662 3426 16696
rect 3426 16662 3460 16696
rect 3460 16662 3469 16696
rect 3417 16654 3469 16662
rect 3978 16696 4030 16707
rect 3978 16662 3987 16696
rect 3987 16662 4021 16696
rect 4021 16662 4030 16696
rect 3978 16655 4030 16662
rect 4169 16696 4221 16707
rect 4169 16662 4179 16696
rect 4179 16662 4213 16696
rect 4213 16662 4221 16696
rect 4169 16655 4221 16662
rect 4361 16696 4413 16707
rect 4361 16662 4371 16696
rect 4371 16662 4405 16696
rect 4405 16662 4413 16696
rect 4361 16655 4413 16662
rect 4553 16696 4605 16707
rect 4553 16662 4563 16696
rect 4563 16662 4597 16696
rect 4597 16662 4605 16696
rect 4553 16655 4605 16662
rect 4746 16696 4798 16706
rect 4746 16662 4755 16696
rect 4755 16662 4789 16696
rect 4789 16662 4798 16696
rect 4746 16654 4798 16662
rect 4938 16696 4990 16706
rect 4938 16662 4947 16696
rect 4947 16662 4981 16696
rect 4981 16662 4990 16696
rect 4938 16654 4990 16662
rect 304 16213 356 16223
rect 304 16179 313 16213
rect 313 16179 347 16213
rect 347 16179 356 16213
rect 304 16171 356 16179
rect 497 16213 549 16223
rect 497 16179 505 16213
rect 505 16179 539 16213
rect 539 16179 549 16213
rect 497 16171 549 16179
rect 688 16213 740 16223
rect 688 16179 697 16213
rect 697 16179 731 16213
rect 731 16179 740 16213
rect 688 16171 740 16179
rect 880 16213 932 16223
rect 880 16179 889 16213
rect 889 16179 923 16213
rect 923 16179 932 16213
rect 880 16171 932 16179
rect 1072 16213 1124 16223
rect 1072 16179 1081 16213
rect 1081 16179 1115 16213
rect 1115 16179 1124 16213
rect 1072 16171 1124 16179
rect 1264 16213 1316 16223
rect 1264 16179 1273 16213
rect 1273 16179 1307 16213
rect 1307 16179 1316 16213
rect 1264 16171 1316 16179
rect 1522 16164 1578 16224
rect 1792 16164 1852 16224
rect 2056 15817 2190 15925
rect 2457 16217 2509 16227
rect 2457 16183 2466 16217
rect 2466 16183 2500 16217
rect 2500 16183 2509 16217
rect 2457 16175 2509 16183
rect 2650 16217 2702 16227
rect 2650 16183 2658 16217
rect 2658 16183 2692 16217
rect 2692 16183 2702 16217
rect 2650 16175 2702 16183
rect 2841 16217 2893 16227
rect 2841 16183 2850 16217
rect 2850 16183 2884 16217
rect 2884 16183 2893 16217
rect 2841 16175 2893 16183
rect 3033 16217 3085 16227
rect 3033 16183 3042 16217
rect 3042 16183 3076 16217
rect 3076 16183 3085 16217
rect 3033 16175 3085 16183
rect 3225 16217 3277 16227
rect 3225 16183 3234 16217
rect 3234 16183 3268 16217
rect 3268 16183 3277 16217
rect 3225 16175 3277 16183
rect 3417 16217 3469 16227
rect 3417 16183 3426 16217
rect 3426 16183 3460 16217
rect 3460 16183 3469 16217
rect 3417 16175 3469 16183
rect 1608 15457 1720 15581
rect 304 15405 356 15416
rect 304 15371 313 15405
rect 313 15371 347 15405
rect 347 15371 356 15405
rect 304 15364 356 15371
rect 495 15405 547 15416
rect 495 15371 505 15405
rect 505 15371 539 15405
rect 539 15371 547 15405
rect 495 15364 547 15371
rect 687 15405 739 15416
rect 687 15371 697 15405
rect 697 15371 731 15405
rect 731 15371 739 15405
rect 687 15364 739 15371
rect 879 15405 931 15416
rect 879 15371 889 15405
rect 889 15371 923 15405
rect 923 15371 931 15405
rect 879 15364 931 15371
rect 1072 15405 1124 15415
rect 1072 15371 1081 15405
rect 1081 15371 1115 15405
rect 1115 15371 1124 15405
rect 1072 15363 1124 15371
rect 1264 15405 1316 15415
rect 1264 15371 1273 15405
rect 1273 15371 1307 15405
rect 1307 15371 1316 15405
rect 1264 15363 1316 15371
rect 1468 15363 1524 15419
rect 1930 15365 1986 15421
rect 3978 16217 4030 16227
rect 3978 16183 3987 16217
rect 3987 16183 4021 16217
rect 4021 16183 4030 16217
rect 3978 16175 4030 16183
rect 4171 16217 4223 16227
rect 4171 16183 4179 16217
rect 4179 16183 4213 16217
rect 4213 16183 4223 16217
rect 4171 16175 4223 16183
rect 4362 16217 4414 16227
rect 4362 16183 4371 16217
rect 4371 16183 4405 16217
rect 4405 16183 4414 16217
rect 4362 16175 4414 16183
rect 4554 16217 4606 16227
rect 4554 16183 4563 16217
rect 4563 16183 4597 16217
rect 4597 16183 4606 16217
rect 4554 16175 4606 16183
rect 4746 16217 4798 16227
rect 4746 16183 4755 16217
rect 4755 16183 4789 16217
rect 4789 16183 4798 16217
rect 4746 16175 4798 16183
rect 4938 16217 4990 16227
rect 4938 16183 4947 16217
rect 4947 16183 4981 16217
rect 4981 16183 4990 16217
rect 4938 16175 4990 16183
rect 3681 15631 3733 15650
rect 3681 15598 3691 15631
rect 3691 15598 3725 15631
rect 3725 15598 3733 15631
rect 5337 15672 5389 15682
rect 5337 15638 5348 15672
rect 5348 15638 5382 15672
rect 5382 15638 5389 15672
rect 5337 15630 5389 15638
rect 5449 15677 5501 15684
rect 5449 15643 5450 15677
rect 5450 15643 5484 15677
rect 5484 15643 5501 15677
rect 5449 15632 5501 15643
rect 2457 15409 2509 15420
rect 2457 15375 2466 15409
rect 2466 15375 2500 15409
rect 2500 15375 2509 15409
rect 2457 15368 2509 15375
rect 2648 15409 2700 15420
rect 2648 15375 2658 15409
rect 2658 15375 2692 15409
rect 2692 15375 2700 15409
rect 2648 15368 2700 15375
rect 2840 15409 2892 15420
rect 2840 15375 2850 15409
rect 2850 15375 2884 15409
rect 2884 15375 2892 15409
rect 2840 15368 2892 15375
rect 3032 15409 3084 15420
rect 3032 15375 3042 15409
rect 3042 15375 3076 15409
rect 3076 15375 3084 15409
rect 3032 15368 3084 15375
rect 3225 15409 3277 15419
rect 3225 15375 3234 15409
rect 3234 15375 3268 15409
rect 3268 15375 3277 15409
rect 3225 15367 3277 15375
rect 3417 15409 3469 15419
rect 3417 15375 3426 15409
rect 3426 15375 3460 15409
rect 3460 15375 3469 15409
rect 3417 15367 3469 15375
rect 3978 15409 4030 15420
rect 3978 15375 3987 15409
rect 3987 15375 4021 15409
rect 4021 15375 4030 15409
rect 3978 15368 4030 15375
rect 4169 15409 4221 15420
rect 4169 15375 4179 15409
rect 4179 15375 4213 15409
rect 4213 15375 4221 15409
rect 4169 15368 4221 15375
rect 4361 15409 4413 15420
rect 4361 15375 4371 15409
rect 4371 15375 4405 15409
rect 4405 15375 4413 15409
rect 4361 15368 4413 15375
rect 4553 15409 4605 15420
rect 4553 15375 4563 15409
rect 4563 15375 4597 15409
rect 4597 15375 4605 15409
rect 4553 15368 4605 15375
rect 4746 15409 4798 15419
rect 4746 15375 4755 15409
rect 4755 15375 4789 15409
rect 4789 15375 4798 15409
rect 4746 15367 4798 15375
rect 4938 15409 4990 15419
rect 4938 15375 4947 15409
rect 4947 15375 4981 15409
rect 4981 15375 4990 15409
rect 4938 15367 4990 15375
rect 304 14926 356 14936
rect 304 14892 313 14926
rect 313 14892 347 14926
rect 347 14892 356 14926
rect 304 14884 356 14892
rect 497 14926 549 14936
rect 497 14892 505 14926
rect 505 14892 539 14926
rect 539 14892 549 14926
rect 497 14884 549 14892
rect 688 14926 740 14936
rect 688 14892 697 14926
rect 697 14892 731 14926
rect 731 14892 740 14926
rect 688 14884 740 14892
rect 880 14926 932 14936
rect 880 14892 889 14926
rect 889 14892 923 14926
rect 923 14892 932 14926
rect 880 14884 932 14892
rect 1072 14926 1124 14936
rect 1072 14892 1081 14926
rect 1081 14892 1115 14926
rect 1115 14892 1124 14926
rect 1072 14884 1124 14892
rect 1264 14926 1316 14936
rect 1264 14892 1273 14926
rect 1273 14892 1307 14926
rect 1307 14892 1316 14926
rect 1264 14884 1316 14892
rect 1522 14877 1578 14937
rect 1792 14877 1852 14937
rect 2056 14530 2190 14638
rect 2457 14930 2509 14940
rect 2457 14896 2466 14930
rect 2466 14896 2500 14930
rect 2500 14896 2509 14930
rect 2457 14888 2509 14896
rect 2650 14930 2702 14940
rect 2650 14896 2658 14930
rect 2658 14896 2692 14930
rect 2692 14896 2702 14930
rect 2650 14888 2702 14896
rect 2841 14930 2893 14940
rect 2841 14896 2850 14930
rect 2850 14896 2884 14930
rect 2884 14896 2893 14930
rect 2841 14888 2893 14896
rect 3033 14930 3085 14940
rect 3033 14896 3042 14930
rect 3042 14896 3076 14930
rect 3076 14896 3085 14930
rect 3033 14888 3085 14896
rect 3225 14930 3277 14940
rect 3225 14896 3234 14930
rect 3234 14896 3268 14930
rect 3268 14896 3277 14930
rect 3225 14888 3277 14896
rect 3417 14930 3469 14940
rect 3417 14896 3426 14930
rect 3426 14896 3460 14930
rect 3460 14896 3469 14930
rect 3417 14888 3469 14896
rect 1608 14170 1720 14294
rect 304 14118 356 14129
rect 304 14084 313 14118
rect 313 14084 347 14118
rect 347 14084 356 14118
rect 304 14077 356 14084
rect 495 14118 547 14129
rect 495 14084 505 14118
rect 505 14084 539 14118
rect 539 14084 547 14118
rect 495 14077 547 14084
rect 687 14118 739 14129
rect 687 14084 697 14118
rect 697 14084 731 14118
rect 731 14084 739 14118
rect 687 14077 739 14084
rect 879 14118 931 14129
rect 879 14084 889 14118
rect 889 14084 923 14118
rect 923 14084 931 14118
rect 879 14077 931 14084
rect 1072 14118 1124 14128
rect 1072 14084 1081 14118
rect 1081 14084 1115 14118
rect 1115 14084 1124 14118
rect 1072 14076 1124 14084
rect 1264 14118 1316 14128
rect 1264 14084 1273 14118
rect 1273 14084 1307 14118
rect 1307 14084 1316 14118
rect 1264 14076 1316 14084
rect 1468 14076 1524 14132
rect 1930 14078 1986 14134
rect 3978 14930 4030 14940
rect 3978 14896 3987 14930
rect 3987 14896 4021 14930
rect 4021 14896 4030 14930
rect 3978 14888 4030 14896
rect 4171 14930 4223 14940
rect 4171 14896 4179 14930
rect 4179 14896 4213 14930
rect 4213 14896 4223 14930
rect 4171 14888 4223 14896
rect 4362 14930 4414 14940
rect 4362 14896 4371 14930
rect 4371 14896 4405 14930
rect 4405 14896 4414 14930
rect 4362 14888 4414 14896
rect 4554 14930 4606 14940
rect 4554 14896 4563 14930
rect 4563 14896 4597 14930
rect 4597 14896 4606 14930
rect 4554 14888 4606 14896
rect 4746 14930 4798 14940
rect 4746 14896 4755 14930
rect 4755 14896 4789 14930
rect 4789 14896 4798 14930
rect 4746 14888 4798 14896
rect 4938 14930 4990 14940
rect 4938 14896 4947 14930
rect 4947 14896 4981 14930
rect 4981 14896 4990 14930
rect 4938 14888 4990 14896
rect 3681 14344 3733 14363
rect 3681 14311 3691 14344
rect 3691 14311 3725 14344
rect 3725 14311 3733 14344
rect 5337 14385 5389 14395
rect 5337 14351 5348 14385
rect 5348 14351 5382 14385
rect 5382 14351 5389 14385
rect 5337 14343 5389 14351
rect 5449 14390 5501 14397
rect 5449 14356 5450 14390
rect 5450 14356 5484 14390
rect 5484 14356 5501 14390
rect 5449 14345 5501 14356
rect 2457 14122 2509 14133
rect 2457 14088 2466 14122
rect 2466 14088 2500 14122
rect 2500 14088 2509 14122
rect 2457 14081 2509 14088
rect 2648 14122 2700 14133
rect 2648 14088 2658 14122
rect 2658 14088 2692 14122
rect 2692 14088 2700 14122
rect 2648 14081 2700 14088
rect 2840 14122 2892 14133
rect 2840 14088 2850 14122
rect 2850 14088 2884 14122
rect 2884 14088 2892 14122
rect 2840 14081 2892 14088
rect 3032 14122 3084 14133
rect 3032 14088 3042 14122
rect 3042 14088 3076 14122
rect 3076 14088 3084 14122
rect 3032 14081 3084 14088
rect 3225 14122 3277 14132
rect 3225 14088 3234 14122
rect 3234 14088 3268 14122
rect 3268 14088 3277 14122
rect 3225 14080 3277 14088
rect 3417 14122 3469 14132
rect 3417 14088 3426 14122
rect 3426 14088 3460 14122
rect 3460 14088 3469 14122
rect 3417 14080 3469 14088
rect 3978 14122 4030 14133
rect 3978 14088 3987 14122
rect 3987 14088 4021 14122
rect 4021 14088 4030 14122
rect 3978 14081 4030 14088
rect 4169 14122 4221 14133
rect 4169 14088 4179 14122
rect 4179 14088 4213 14122
rect 4213 14088 4221 14122
rect 4169 14081 4221 14088
rect 4361 14122 4413 14133
rect 4361 14088 4371 14122
rect 4371 14088 4405 14122
rect 4405 14088 4413 14122
rect 4361 14081 4413 14088
rect 4553 14122 4605 14133
rect 4553 14088 4563 14122
rect 4563 14088 4597 14122
rect 4597 14088 4605 14122
rect 4553 14081 4605 14088
rect 4746 14122 4798 14132
rect 4746 14088 4755 14122
rect 4755 14088 4789 14122
rect 4789 14088 4798 14122
rect 4746 14080 4798 14088
rect 4938 14122 4990 14132
rect 4938 14088 4947 14122
rect 4947 14088 4981 14122
rect 4981 14088 4990 14122
rect 4938 14080 4990 14088
rect 304 13639 356 13649
rect 304 13605 313 13639
rect 313 13605 347 13639
rect 347 13605 356 13639
rect 304 13597 356 13605
rect 497 13639 549 13649
rect 497 13605 505 13639
rect 505 13605 539 13639
rect 539 13605 549 13639
rect 497 13597 549 13605
rect 688 13639 740 13649
rect 688 13605 697 13639
rect 697 13605 731 13639
rect 731 13605 740 13639
rect 688 13597 740 13605
rect 880 13639 932 13649
rect 880 13605 889 13639
rect 889 13605 923 13639
rect 923 13605 932 13639
rect 880 13597 932 13605
rect 1072 13639 1124 13649
rect 1072 13605 1081 13639
rect 1081 13605 1115 13639
rect 1115 13605 1124 13639
rect 1072 13597 1124 13605
rect 1264 13639 1316 13649
rect 1264 13605 1273 13639
rect 1273 13605 1307 13639
rect 1307 13605 1316 13639
rect 1264 13597 1316 13605
rect 1522 13590 1578 13650
rect 1792 13590 1852 13650
rect 2056 13243 2190 13351
rect 2457 13643 2509 13653
rect 2457 13609 2466 13643
rect 2466 13609 2500 13643
rect 2500 13609 2509 13643
rect 2457 13601 2509 13609
rect 2650 13643 2702 13653
rect 2650 13609 2658 13643
rect 2658 13609 2692 13643
rect 2692 13609 2702 13643
rect 2650 13601 2702 13609
rect 2841 13643 2893 13653
rect 2841 13609 2850 13643
rect 2850 13609 2884 13643
rect 2884 13609 2893 13643
rect 2841 13601 2893 13609
rect 3033 13643 3085 13653
rect 3033 13609 3042 13643
rect 3042 13609 3076 13643
rect 3076 13609 3085 13643
rect 3033 13601 3085 13609
rect 3225 13643 3277 13653
rect 3225 13609 3234 13643
rect 3234 13609 3268 13643
rect 3268 13609 3277 13643
rect 3225 13601 3277 13609
rect 3417 13643 3469 13653
rect 3417 13609 3426 13643
rect 3426 13609 3460 13643
rect 3460 13609 3469 13643
rect 3417 13601 3469 13609
rect 1608 12883 1720 13007
rect 304 12831 356 12842
rect 304 12797 313 12831
rect 313 12797 347 12831
rect 347 12797 356 12831
rect 304 12790 356 12797
rect 495 12831 547 12842
rect 495 12797 505 12831
rect 505 12797 539 12831
rect 539 12797 547 12831
rect 495 12790 547 12797
rect 687 12831 739 12842
rect 687 12797 697 12831
rect 697 12797 731 12831
rect 731 12797 739 12831
rect 687 12790 739 12797
rect 879 12831 931 12842
rect 879 12797 889 12831
rect 889 12797 923 12831
rect 923 12797 931 12831
rect 879 12790 931 12797
rect 1072 12831 1124 12841
rect 1072 12797 1081 12831
rect 1081 12797 1115 12831
rect 1115 12797 1124 12831
rect 1072 12789 1124 12797
rect 1264 12831 1316 12841
rect 1264 12797 1273 12831
rect 1273 12797 1307 12831
rect 1307 12797 1316 12831
rect 1264 12789 1316 12797
rect 1468 12789 1524 12845
rect 1930 12791 1986 12847
rect 3978 13643 4030 13653
rect 3978 13609 3987 13643
rect 3987 13609 4021 13643
rect 4021 13609 4030 13643
rect 3978 13601 4030 13609
rect 4171 13643 4223 13653
rect 4171 13609 4179 13643
rect 4179 13609 4213 13643
rect 4213 13609 4223 13643
rect 4171 13601 4223 13609
rect 4362 13643 4414 13653
rect 4362 13609 4371 13643
rect 4371 13609 4405 13643
rect 4405 13609 4414 13643
rect 4362 13601 4414 13609
rect 4554 13643 4606 13653
rect 4554 13609 4563 13643
rect 4563 13609 4597 13643
rect 4597 13609 4606 13643
rect 4554 13601 4606 13609
rect 4746 13643 4798 13653
rect 4746 13609 4755 13643
rect 4755 13609 4789 13643
rect 4789 13609 4798 13643
rect 4746 13601 4798 13609
rect 4938 13643 4990 13653
rect 4938 13609 4947 13643
rect 4947 13609 4981 13643
rect 4981 13609 4990 13643
rect 4938 13601 4990 13609
rect 3681 13057 3733 13076
rect 3681 13024 3691 13057
rect 3691 13024 3725 13057
rect 3725 13024 3733 13057
rect 5337 13098 5389 13108
rect 5337 13064 5348 13098
rect 5348 13064 5382 13098
rect 5382 13064 5389 13098
rect 5337 13056 5389 13064
rect 5449 13103 5501 13110
rect 5449 13069 5450 13103
rect 5450 13069 5484 13103
rect 5484 13069 5501 13103
rect 5449 13058 5501 13069
rect 2457 12835 2509 12846
rect 2457 12801 2466 12835
rect 2466 12801 2500 12835
rect 2500 12801 2509 12835
rect 2457 12794 2509 12801
rect 2648 12835 2700 12846
rect 2648 12801 2658 12835
rect 2658 12801 2692 12835
rect 2692 12801 2700 12835
rect 2648 12794 2700 12801
rect 2840 12835 2892 12846
rect 2840 12801 2850 12835
rect 2850 12801 2884 12835
rect 2884 12801 2892 12835
rect 2840 12794 2892 12801
rect 3032 12835 3084 12846
rect 3032 12801 3042 12835
rect 3042 12801 3076 12835
rect 3076 12801 3084 12835
rect 3032 12794 3084 12801
rect 3225 12835 3277 12845
rect 3225 12801 3234 12835
rect 3234 12801 3268 12835
rect 3268 12801 3277 12835
rect 3225 12793 3277 12801
rect 3417 12835 3469 12845
rect 3417 12801 3426 12835
rect 3426 12801 3460 12835
rect 3460 12801 3469 12835
rect 3417 12793 3469 12801
rect 3978 12835 4030 12846
rect 3978 12801 3987 12835
rect 3987 12801 4021 12835
rect 4021 12801 4030 12835
rect 3978 12794 4030 12801
rect 4169 12835 4221 12846
rect 4169 12801 4179 12835
rect 4179 12801 4213 12835
rect 4213 12801 4221 12835
rect 4169 12794 4221 12801
rect 4361 12835 4413 12846
rect 4361 12801 4371 12835
rect 4371 12801 4405 12835
rect 4405 12801 4413 12835
rect 4361 12794 4413 12801
rect 4553 12835 4605 12846
rect 4553 12801 4563 12835
rect 4563 12801 4597 12835
rect 4597 12801 4605 12835
rect 4553 12794 4605 12801
rect 4746 12835 4798 12845
rect 4746 12801 4755 12835
rect 4755 12801 4789 12835
rect 4789 12801 4798 12835
rect 4746 12793 4798 12801
rect 4938 12835 4990 12845
rect 4938 12801 4947 12835
rect 4947 12801 4981 12835
rect 4981 12801 4990 12835
rect 4938 12793 4990 12801
rect 304 12352 356 12362
rect 304 12318 313 12352
rect 313 12318 347 12352
rect 347 12318 356 12352
rect 304 12310 356 12318
rect 497 12352 549 12362
rect 497 12318 505 12352
rect 505 12318 539 12352
rect 539 12318 549 12352
rect 497 12310 549 12318
rect 688 12352 740 12362
rect 688 12318 697 12352
rect 697 12318 731 12352
rect 731 12318 740 12352
rect 688 12310 740 12318
rect 880 12352 932 12362
rect 880 12318 889 12352
rect 889 12318 923 12352
rect 923 12318 932 12352
rect 880 12310 932 12318
rect 1072 12352 1124 12362
rect 1072 12318 1081 12352
rect 1081 12318 1115 12352
rect 1115 12318 1124 12352
rect 1072 12310 1124 12318
rect 1264 12352 1316 12362
rect 1264 12318 1273 12352
rect 1273 12318 1307 12352
rect 1307 12318 1316 12352
rect 1264 12310 1316 12318
rect 1522 12303 1578 12363
rect 1792 12303 1852 12363
rect 2056 11956 2190 12064
rect 2457 12356 2509 12366
rect 2457 12322 2466 12356
rect 2466 12322 2500 12356
rect 2500 12322 2509 12356
rect 2457 12314 2509 12322
rect 2650 12356 2702 12366
rect 2650 12322 2658 12356
rect 2658 12322 2692 12356
rect 2692 12322 2702 12356
rect 2650 12314 2702 12322
rect 2841 12356 2893 12366
rect 2841 12322 2850 12356
rect 2850 12322 2884 12356
rect 2884 12322 2893 12356
rect 2841 12314 2893 12322
rect 3033 12356 3085 12366
rect 3033 12322 3042 12356
rect 3042 12322 3076 12356
rect 3076 12322 3085 12356
rect 3033 12314 3085 12322
rect 3225 12356 3277 12366
rect 3225 12322 3234 12356
rect 3234 12322 3268 12356
rect 3268 12322 3277 12356
rect 3225 12314 3277 12322
rect 3417 12356 3469 12366
rect 3417 12322 3426 12356
rect 3426 12322 3460 12356
rect 3460 12322 3469 12356
rect 3417 12314 3469 12322
rect 1608 11596 1720 11720
rect 304 11544 356 11555
rect 304 11510 313 11544
rect 313 11510 347 11544
rect 347 11510 356 11544
rect 304 11503 356 11510
rect 495 11544 547 11555
rect 495 11510 505 11544
rect 505 11510 539 11544
rect 539 11510 547 11544
rect 495 11503 547 11510
rect 687 11544 739 11555
rect 687 11510 697 11544
rect 697 11510 731 11544
rect 731 11510 739 11544
rect 687 11503 739 11510
rect 879 11544 931 11555
rect 879 11510 889 11544
rect 889 11510 923 11544
rect 923 11510 931 11544
rect 879 11503 931 11510
rect 1072 11544 1124 11554
rect 1072 11510 1081 11544
rect 1081 11510 1115 11544
rect 1115 11510 1124 11544
rect 1072 11502 1124 11510
rect 1264 11544 1316 11554
rect 1264 11510 1273 11544
rect 1273 11510 1307 11544
rect 1307 11510 1316 11544
rect 1264 11502 1316 11510
rect 1468 11502 1524 11558
rect 1930 11504 1986 11560
rect 3978 12356 4030 12366
rect 3978 12322 3987 12356
rect 3987 12322 4021 12356
rect 4021 12322 4030 12356
rect 3978 12314 4030 12322
rect 4171 12356 4223 12366
rect 4171 12322 4179 12356
rect 4179 12322 4213 12356
rect 4213 12322 4223 12356
rect 4171 12314 4223 12322
rect 4362 12356 4414 12366
rect 4362 12322 4371 12356
rect 4371 12322 4405 12356
rect 4405 12322 4414 12356
rect 4362 12314 4414 12322
rect 4554 12356 4606 12366
rect 4554 12322 4563 12356
rect 4563 12322 4597 12356
rect 4597 12322 4606 12356
rect 4554 12314 4606 12322
rect 4746 12356 4798 12366
rect 4746 12322 4755 12356
rect 4755 12322 4789 12356
rect 4789 12322 4798 12356
rect 4746 12314 4798 12322
rect 4938 12356 4990 12366
rect 4938 12322 4947 12356
rect 4947 12322 4981 12356
rect 4981 12322 4990 12356
rect 4938 12314 4990 12322
rect 3681 11770 3733 11789
rect 3681 11737 3691 11770
rect 3691 11737 3725 11770
rect 3725 11737 3733 11770
rect 5337 11811 5389 11821
rect 5337 11777 5348 11811
rect 5348 11777 5382 11811
rect 5382 11777 5389 11811
rect 5337 11769 5389 11777
rect 5449 11816 5501 11823
rect 5449 11782 5450 11816
rect 5450 11782 5484 11816
rect 5484 11782 5501 11816
rect 5449 11771 5501 11782
rect 2457 11548 2509 11559
rect 2457 11514 2466 11548
rect 2466 11514 2500 11548
rect 2500 11514 2509 11548
rect 2457 11507 2509 11514
rect 2648 11548 2700 11559
rect 2648 11514 2658 11548
rect 2658 11514 2692 11548
rect 2692 11514 2700 11548
rect 2648 11507 2700 11514
rect 2840 11548 2892 11559
rect 2840 11514 2850 11548
rect 2850 11514 2884 11548
rect 2884 11514 2892 11548
rect 2840 11507 2892 11514
rect 3032 11548 3084 11559
rect 3032 11514 3042 11548
rect 3042 11514 3076 11548
rect 3076 11514 3084 11548
rect 3032 11507 3084 11514
rect 3225 11548 3277 11558
rect 3225 11514 3234 11548
rect 3234 11514 3268 11548
rect 3268 11514 3277 11548
rect 3225 11506 3277 11514
rect 3417 11548 3469 11558
rect 3417 11514 3426 11548
rect 3426 11514 3460 11548
rect 3460 11514 3469 11548
rect 3417 11506 3469 11514
rect 3978 11548 4030 11559
rect 3978 11514 3987 11548
rect 3987 11514 4021 11548
rect 4021 11514 4030 11548
rect 3978 11507 4030 11514
rect 4169 11548 4221 11559
rect 4169 11514 4179 11548
rect 4179 11514 4213 11548
rect 4213 11514 4221 11548
rect 4169 11507 4221 11514
rect 4361 11548 4413 11559
rect 4361 11514 4371 11548
rect 4371 11514 4405 11548
rect 4405 11514 4413 11548
rect 4361 11507 4413 11514
rect 4553 11548 4605 11559
rect 4553 11514 4563 11548
rect 4563 11514 4597 11548
rect 4597 11514 4605 11548
rect 4553 11507 4605 11514
rect 4746 11548 4798 11558
rect 4746 11514 4755 11548
rect 4755 11514 4789 11548
rect 4789 11514 4798 11548
rect 4746 11506 4798 11514
rect 4938 11548 4990 11558
rect 4938 11514 4947 11548
rect 4947 11514 4981 11548
rect 4981 11514 4990 11548
rect 4938 11506 4990 11514
rect 304 11065 356 11075
rect 304 11031 313 11065
rect 313 11031 347 11065
rect 347 11031 356 11065
rect 304 11023 356 11031
rect 497 11065 549 11075
rect 497 11031 505 11065
rect 505 11031 539 11065
rect 539 11031 549 11065
rect 497 11023 549 11031
rect 688 11065 740 11075
rect 688 11031 697 11065
rect 697 11031 731 11065
rect 731 11031 740 11065
rect 688 11023 740 11031
rect 880 11065 932 11075
rect 880 11031 889 11065
rect 889 11031 923 11065
rect 923 11031 932 11065
rect 880 11023 932 11031
rect 1072 11065 1124 11075
rect 1072 11031 1081 11065
rect 1081 11031 1115 11065
rect 1115 11031 1124 11065
rect 1072 11023 1124 11031
rect 1264 11065 1316 11075
rect 1264 11031 1273 11065
rect 1273 11031 1307 11065
rect 1307 11031 1316 11065
rect 1264 11023 1316 11031
rect 1522 11016 1578 11076
rect 1792 11016 1852 11076
rect 2056 10669 2190 10777
rect 2457 11069 2509 11079
rect 2457 11035 2466 11069
rect 2466 11035 2500 11069
rect 2500 11035 2509 11069
rect 2457 11027 2509 11035
rect 2650 11069 2702 11079
rect 2650 11035 2658 11069
rect 2658 11035 2692 11069
rect 2692 11035 2702 11069
rect 2650 11027 2702 11035
rect 2841 11069 2893 11079
rect 2841 11035 2850 11069
rect 2850 11035 2884 11069
rect 2884 11035 2893 11069
rect 2841 11027 2893 11035
rect 3033 11069 3085 11079
rect 3033 11035 3042 11069
rect 3042 11035 3076 11069
rect 3076 11035 3085 11069
rect 3033 11027 3085 11035
rect 3225 11069 3277 11079
rect 3225 11035 3234 11069
rect 3234 11035 3268 11069
rect 3268 11035 3277 11069
rect 3225 11027 3277 11035
rect 3417 11069 3469 11079
rect 3417 11035 3426 11069
rect 3426 11035 3460 11069
rect 3460 11035 3469 11069
rect 3417 11027 3469 11035
rect 1608 10309 1720 10433
rect 304 10257 356 10268
rect 304 10223 313 10257
rect 313 10223 347 10257
rect 347 10223 356 10257
rect 304 10216 356 10223
rect 495 10257 547 10268
rect 495 10223 505 10257
rect 505 10223 539 10257
rect 539 10223 547 10257
rect 495 10216 547 10223
rect 687 10257 739 10268
rect 687 10223 697 10257
rect 697 10223 731 10257
rect 731 10223 739 10257
rect 687 10216 739 10223
rect 879 10257 931 10268
rect 879 10223 889 10257
rect 889 10223 923 10257
rect 923 10223 931 10257
rect 879 10216 931 10223
rect 1072 10257 1124 10267
rect 1072 10223 1081 10257
rect 1081 10223 1115 10257
rect 1115 10223 1124 10257
rect 1072 10215 1124 10223
rect 1264 10257 1316 10267
rect 1264 10223 1273 10257
rect 1273 10223 1307 10257
rect 1307 10223 1316 10257
rect 1264 10215 1316 10223
rect 1468 10215 1524 10271
rect 1930 10217 1986 10273
rect 3978 11069 4030 11079
rect 3978 11035 3987 11069
rect 3987 11035 4021 11069
rect 4021 11035 4030 11069
rect 3978 11027 4030 11035
rect 4171 11069 4223 11079
rect 4171 11035 4179 11069
rect 4179 11035 4213 11069
rect 4213 11035 4223 11069
rect 4171 11027 4223 11035
rect 4362 11069 4414 11079
rect 4362 11035 4371 11069
rect 4371 11035 4405 11069
rect 4405 11035 4414 11069
rect 4362 11027 4414 11035
rect 4554 11069 4606 11079
rect 4554 11035 4563 11069
rect 4563 11035 4597 11069
rect 4597 11035 4606 11069
rect 4554 11027 4606 11035
rect 4746 11069 4798 11079
rect 4746 11035 4755 11069
rect 4755 11035 4789 11069
rect 4789 11035 4798 11069
rect 4746 11027 4798 11035
rect 4938 11069 4990 11079
rect 4938 11035 4947 11069
rect 4947 11035 4981 11069
rect 4981 11035 4990 11069
rect 4938 11027 4990 11035
rect 3681 10483 3733 10502
rect 3681 10450 3691 10483
rect 3691 10450 3725 10483
rect 3725 10450 3733 10483
rect 5337 10524 5389 10534
rect 5337 10490 5348 10524
rect 5348 10490 5382 10524
rect 5382 10490 5389 10524
rect 5337 10482 5389 10490
rect 5449 10529 5501 10536
rect 5449 10495 5450 10529
rect 5450 10495 5484 10529
rect 5484 10495 5501 10529
rect 5449 10484 5501 10495
rect 2457 10261 2509 10272
rect 2457 10227 2466 10261
rect 2466 10227 2500 10261
rect 2500 10227 2509 10261
rect 2457 10220 2509 10227
rect 2648 10261 2700 10272
rect 2648 10227 2658 10261
rect 2658 10227 2692 10261
rect 2692 10227 2700 10261
rect 2648 10220 2700 10227
rect 2840 10261 2892 10272
rect 2840 10227 2850 10261
rect 2850 10227 2884 10261
rect 2884 10227 2892 10261
rect 2840 10220 2892 10227
rect 3032 10261 3084 10272
rect 3032 10227 3042 10261
rect 3042 10227 3076 10261
rect 3076 10227 3084 10261
rect 3032 10220 3084 10227
rect 3225 10261 3277 10271
rect 3225 10227 3234 10261
rect 3234 10227 3268 10261
rect 3268 10227 3277 10261
rect 3225 10219 3277 10227
rect 3417 10261 3469 10271
rect 3417 10227 3426 10261
rect 3426 10227 3460 10261
rect 3460 10227 3469 10261
rect 3417 10219 3469 10227
rect 3978 10261 4030 10272
rect 3978 10227 3987 10261
rect 3987 10227 4021 10261
rect 4021 10227 4030 10261
rect 3978 10220 4030 10227
rect 4169 10261 4221 10272
rect 4169 10227 4179 10261
rect 4179 10227 4213 10261
rect 4213 10227 4221 10261
rect 4169 10220 4221 10227
rect 4361 10261 4413 10272
rect 4361 10227 4371 10261
rect 4371 10227 4405 10261
rect 4405 10227 4413 10261
rect 4361 10220 4413 10227
rect 4553 10261 4605 10272
rect 4553 10227 4563 10261
rect 4563 10227 4597 10261
rect 4597 10227 4605 10261
rect 4553 10220 4605 10227
rect 4746 10261 4798 10271
rect 4746 10227 4755 10261
rect 4755 10227 4789 10261
rect 4789 10227 4798 10261
rect 4746 10219 4798 10227
rect 4938 10261 4990 10271
rect 4938 10227 4947 10261
rect 4947 10227 4981 10261
rect 4981 10227 4990 10261
rect 4938 10219 4990 10227
rect 304 9778 356 9788
rect 304 9744 313 9778
rect 313 9744 347 9778
rect 347 9744 356 9778
rect 304 9736 356 9744
rect 497 9778 549 9788
rect 497 9744 505 9778
rect 505 9744 539 9778
rect 539 9744 549 9778
rect 497 9736 549 9744
rect 688 9778 740 9788
rect 688 9744 697 9778
rect 697 9744 731 9778
rect 731 9744 740 9778
rect 688 9736 740 9744
rect 880 9778 932 9788
rect 880 9744 889 9778
rect 889 9744 923 9778
rect 923 9744 932 9778
rect 880 9736 932 9744
rect 1072 9778 1124 9788
rect 1072 9744 1081 9778
rect 1081 9744 1115 9778
rect 1115 9744 1124 9778
rect 1072 9736 1124 9744
rect 1264 9778 1316 9788
rect 1264 9744 1273 9778
rect 1273 9744 1307 9778
rect 1307 9744 1316 9778
rect 1264 9736 1316 9744
rect 1522 9729 1578 9789
rect 1792 9729 1852 9789
rect 2056 9382 2190 9490
rect 2457 9782 2509 9792
rect 2457 9748 2466 9782
rect 2466 9748 2500 9782
rect 2500 9748 2509 9782
rect 2457 9740 2509 9748
rect 2650 9782 2702 9792
rect 2650 9748 2658 9782
rect 2658 9748 2692 9782
rect 2692 9748 2702 9782
rect 2650 9740 2702 9748
rect 2841 9782 2893 9792
rect 2841 9748 2850 9782
rect 2850 9748 2884 9782
rect 2884 9748 2893 9782
rect 2841 9740 2893 9748
rect 3033 9782 3085 9792
rect 3033 9748 3042 9782
rect 3042 9748 3076 9782
rect 3076 9748 3085 9782
rect 3033 9740 3085 9748
rect 3225 9782 3277 9792
rect 3225 9748 3234 9782
rect 3234 9748 3268 9782
rect 3268 9748 3277 9782
rect 3225 9740 3277 9748
rect 3417 9782 3469 9792
rect 3417 9748 3426 9782
rect 3426 9748 3460 9782
rect 3460 9748 3469 9782
rect 3417 9740 3469 9748
rect 1608 9022 1720 9146
rect 304 8970 356 8981
rect 304 8936 313 8970
rect 313 8936 347 8970
rect 347 8936 356 8970
rect 304 8929 356 8936
rect 495 8970 547 8981
rect 495 8936 505 8970
rect 505 8936 539 8970
rect 539 8936 547 8970
rect 495 8929 547 8936
rect 687 8970 739 8981
rect 687 8936 697 8970
rect 697 8936 731 8970
rect 731 8936 739 8970
rect 687 8929 739 8936
rect 879 8970 931 8981
rect 879 8936 889 8970
rect 889 8936 923 8970
rect 923 8936 931 8970
rect 879 8929 931 8936
rect 1072 8970 1124 8980
rect 1072 8936 1081 8970
rect 1081 8936 1115 8970
rect 1115 8936 1124 8970
rect 1072 8928 1124 8936
rect 1264 8970 1316 8980
rect 1264 8936 1273 8970
rect 1273 8936 1307 8970
rect 1307 8936 1316 8970
rect 1264 8928 1316 8936
rect 1468 8928 1524 8984
rect 1930 8930 1986 8986
rect 3978 9782 4030 9792
rect 3978 9748 3987 9782
rect 3987 9748 4021 9782
rect 4021 9748 4030 9782
rect 3978 9740 4030 9748
rect 4171 9782 4223 9792
rect 4171 9748 4179 9782
rect 4179 9748 4213 9782
rect 4213 9748 4223 9782
rect 4171 9740 4223 9748
rect 4362 9782 4414 9792
rect 4362 9748 4371 9782
rect 4371 9748 4405 9782
rect 4405 9748 4414 9782
rect 4362 9740 4414 9748
rect 4554 9782 4606 9792
rect 4554 9748 4563 9782
rect 4563 9748 4597 9782
rect 4597 9748 4606 9782
rect 4554 9740 4606 9748
rect 4746 9782 4798 9792
rect 4746 9748 4755 9782
rect 4755 9748 4789 9782
rect 4789 9748 4798 9782
rect 4746 9740 4798 9748
rect 4938 9782 4990 9792
rect 4938 9748 4947 9782
rect 4947 9748 4981 9782
rect 4981 9748 4990 9782
rect 4938 9740 4990 9748
rect 3681 9196 3733 9215
rect 3681 9163 3691 9196
rect 3691 9163 3725 9196
rect 3725 9163 3733 9196
rect 5337 9237 5389 9247
rect 5337 9203 5348 9237
rect 5348 9203 5382 9237
rect 5382 9203 5389 9237
rect 5337 9195 5389 9203
rect 5449 9242 5501 9249
rect 5449 9208 5450 9242
rect 5450 9208 5484 9242
rect 5484 9208 5501 9242
rect 5449 9197 5501 9208
rect 2457 8974 2509 8985
rect 2457 8940 2466 8974
rect 2466 8940 2500 8974
rect 2500 8940 2509 8974
rect 2457 8933 2509 8940
rect 2648 8974 2700 8985
rect 2648 8940 2658 8974
rect 2658 8940 2692 8974
rect 2692 8940 2700 8974
rect 2648 8933 2700 8940
rect 2840 8974 2892 8985
rect 2840 8940 2850 8974
rect 2850 8940 2884 8974
rect 2884 8940 2892 8974
rect 2840 8933 2892 8940
rect 3032 8974 3084 8985
rect 3032 8940 3042 8974
rect 3042 8940 3076 8974
rect 3076 8940 3084 8974
rect 3032 8933 3084 8940
rect 3225 8974 3277 8984
rect 3225 8940 3234 8974
rect 3234 8940 3268 8974
rect 3268 8940 3277 8974
rect 3225 8932 3277 8940
rect 3417 8974 3469 8984
rect 3417 8940 3426 8974
rect 3426 8940 3460 8974
rect 3460 8940 3469 8974
rect 3417 8932 3469 8940
rect 3978 8974 4030 8985
rect 3978 8940 3987 8974
rect 3987 8940 4021 8974
rect 4021 8940 4030 8974
rect 3978 8933 4030 8940
rect 4169 8974 4221 8985
rect 4169 8940 4179 8974
rect 4179 8940 4213 8974
rect 4213 8940 4221 8974
rect 4169 8933 4221 8940
rect 4361 8974 4413 8985
rect 4361 8940 4371 8974
rect 4371 8940 4405 8974
rect 4405 8940 4413 8974
rect 4361 8933 4413 8940
rect 4553 8974 4605 8985
rect 4553 8940 4563 8974
rect 4563 8940 4597 8974
rect 4597 8940 4605 8974
rect 4553 8933 4605 8940
rect 4746 8974 4798 8984
rect 4746 8940 4755 8974
rect 4755 8940 4789 8974
rect 4789 8940 4798 8974
rect 4746 8932 4798 8940
rect 4938 8974 4990 8984
rect 4938 8940 4947 8974
rect 4947 8940 4981 8974
rect 4981 8940 4990 8974
rect 4938 8932 4990 8940
rect 304 8491 356 8501
rect 304 8457 313 8491
rect 313 8457 347 8491
rect 347 8457 356 8491
rect 304 8449 356 8457
rect 497 8491 549 8501
rect 497 8457 505 8491
rect 505 8457 539 8491
rect 539 8457 549 8491
rect 497 8449 549 8457
rect 688 8491 740 8501
rect 688 8457 697 8491
rect 697 8457 731 8491
rect 731 8457 740 8491
rect 688 8449 740 8457
rect 880 8491 932 8501
rect 880 8457 889 8491
rect 889 8457 923 8491
rect 923 8457 932 8491
rect 880 8449 932 8457
rect 1072 8491 1124 8501
rect 1072 8457 1081 8491
rect 1081 8457 1115 8491
rect 1115 8457 1124 8491
rect 1072 8449 1124 8457
rect 1264 8491 1316 8501
rect 1264 8457 1273 8491
rect 1273 8457 1307 8491
rect 1307 8457 1316 8491
rect 1264 8449 1316 8457
rect 1522 8442 1578 8502
rect 1792 8442 1852 8502
rect 2056 8095 2190 8203
rect 2457 8495 2509 8505
rect 2457 8461 2466 8495
rect 2466 8461 2500 8495
rect 2500 8461 2509 8495
rect 2457 8453 2509 8461
rect 2650 8495 2702 8505
rect 2650 8461 2658 8495
rect 2658 8461 2692 8495
rect 2692 8461 2702 8495
rect 2650 8453 2702 8461
rect 2841 8495 2893 8505
rect 2841 8461 2850 8495
rect 2850 8461 2884 8495
rect 2884 8461 2893 8495
rect 2841 8453 2893 8461
rect 3033 8495 3085 8505
rect 3033 8461 3042 8495
rect 3042 8461 3076 8495
rect 3076 8461 3085 8495
rect 3033 8453 3085 8461
rect 3225 8495 3277 8505
rect 3225 8461 3234 8495
rect 3234 8461 3268 8495
rect 3268 8461 3277 8495
rect 3225 8453 3277 8461
rect 3417 8495 3469 8505
rect 3417 8461 3426 8495
rect 3426 8461 3460 8495
rect 3460 8461 3469 8495
rect 3417 8453 3469 8461
rect 1608 7735 1720 7859
rect 304 7683 356 7694
rect 304 7649 313 7683
rect 313 7649 347 7683
rect 347 7649 356 7683
rect 304 7642 356 7649
rect 495 7683 547 7694
rect 495 7649 505 7683
rect 505 7649 539 7683
rect 539 7649 547 7683
rect 495 7642 547 7649
rect 687 7683 739 7694
rect 687 7649 697 7683
rect 697 7649 731 7683
rect 731 7649 739 7683
rect 687 7642 739 7649
rect 879 7683 931 7694
rect 879 7649 889 7683
rect 889 7649 923 7683
rect 923 7649 931 7683
rect 879 7642 931 7649
rect 1072 7683 1124 7693
rect 1072 7649 1081 7683
rect 1081 7649 1115 7683
rect 1115 7649 1124 7683
rect 1072 7641 1124 7649
rect 1264 7683 1316 7693
rect 1264 7649 1273 7683
rect 1273 7649 1307 7683
rect 1307 7649 1316 7683
rect 1264 7641 1316 7649
rect 1468 7641 1524 7697
rect 1930 7643 1986 7699
rect 3978 8495 4030 8505
rect 3978 8461 3987 8495
rect 3987 8461 4021 8495
rect 4021 8461 4030 8495
rect 3978 8453 4030 8461
rect 4171 8495 4223 8505
rect 4171 8461 4179 8495
rect 4179 8461 4213 8495
rect 4213 8461 4223 8495
rect 4171 8453 4223 8461
rect 4362 8495 4414 8505
rect 4362 8461 4371 8495
rect 4371 8461 4405 8495
rect 4405 8461 4414 8495
rect 4362 8453 4414 8461
rect 4554 8495 4606 8505
rect 4554 8461 4563 8495
rect 4563 8461 4597 8495
rect 4597 8461 4606 8495
rect 4554 8453 4606 8461
rect 4746 8495 4798 8505
rect 4746 8461 4755 8495
rect 4755 8461 4789 8495
rect 4789 8461 4798 8495
rect 4746 8453 4798 8461
rect 4938 8495 4990 8505
rect 4938 8461 4947 8495
rect 4947 8461 4981 8495
rect 4981 8461 4990 8495
rect 4938 8453 4990 8461
rect 3681 7909 3733 7928
rect 3681 7876 3691 7909
rect 3691 7876 3725 7909
rect 3725 7876 3733 7909
rect 5337 7950 5389 7960
rect 5337 7916 5348 7950
rect 5348 7916 5382 7950
rect 5382 7916 5389 7950
rect 5337 7908 5389 7916
rect 5449 7955 5501 7962
rect 5449 7921 5450 7955
rect 5450 7921 5484 7955
rect 5484 7921 5501 7955
rect 5449 7910 5501 7921
rect 2457 7687 2509 7698
rect 2457 7653 2466 7687
rect 2466 7653 2500 7687
rect 2500 7653 2509 7687
rect 2457 7646 2509 7653
rect 2648 7687 2700 7698
rect 2648 7653 2658 7687
rect 2658 7653 2692 7687
rect 2692 7653 2700 7687
rect 2648 7646 2700 7653
rect 2840 7687 2892 7698
rect 2840 7653 2850 7687
rect 2850 7653 2884 7687
rect 2884 7653 2892 7687
rect 2840 7646 2892 7653
rect 3032 7687 3084 7698
rect 3032 7653 3042 7687
rect 3042 7653 3076 7687
rect 3076 7653 3084 7687
rect 3032 7646 3084 7653
rect 3225 7687 3277 7697
rect 3225 7653 3234 7687
rect 3234 7653 3268 7687
rect 3268 7653 3277 7687
rect 3225 7645 3277 7653
rect 3417 7687 3469 7697
rect 3417 7653 3426 7687
rect 3426 7653 3460 7687
rect 3460 7653 3469 7687
rect 3417 7645 3469 7653
rect 3978 7687 4030 7698
rect 3978 7653 3987 7687
rect 3987 7653 4021 7687
rect 4021 7653 4030 7687
rect 3978 7646 4030 7653
rect 4169 7687 4221 7698
rect 4169 7653 4179 7687
rect 4179 7653 4213 7687
rect 4213 7653 4221 7687
rect 4169 7646 4221 7653
rect 4361 7687 4413 7698
rect 4361 7653 4371 7687
rect 4371 7653 4405 7687
rect 4405 7653 4413 7687
rect 4361 7646 4413 7653
rect 4553 7687 4605 7698
rect 4553 7653 4563 7687
rect 4563 7653 4597 7687
rect 4597 7653 4605 7687
rect 4553 7646 4605 7653
rect 4746 7687 4798 7697
rect 4746 7653 4755 7687
rect 4755 7653 4789 7687
rect 4789 7653 4798 7687
rect 4746 7645 4798 7653
rect 4938 7687 4990 7697
rect 4938 7653 4947 7687
rect 4947 7653 4981 7687
rect 4981 7653 4990 7687
rect 4938 7645 4990 7653
rect 304 7204 356 7214
rect 304 7170 313 7204
rect 313 7170 347 7204
rect 347 7170 356 7204
rect 304 7162 356 7170
rect 497 7204 549 7214
rect 497 7170 505 7204
rect 505 7170 539 7204
rect 539 7170 549 7204
rect 497 7162 549 7170
rect 688 7204 740 7214
rect 688 7170 697 7204
rect 697 7170 731 7204
rect 731 7170 740 7204
rect 688 7162 740 7170
rect 880 7204 932 7214
rect 880 7170 889 7204
rect 889 7170 923 7204
rect 923 7170 932 7204
rect 880 7162 932 7170
rect 1072 7204 1124 7214
rect 1072 7170 1081 7204
rect 1081 7170 1115 7204
rect 1115 7170 1124 7204
rect 1072 7162 1124 7170
rect 1264 7204 1316 7214
rect 1264 7170 1273 7204
rect 1273 7170 1307 7204
rect 1307 7170 1316 7204
rect 1264 7162 1316 7170
rect 1522 7155 1578 7215
rect 1792 7155 1852 7215
rect 2056 6808 2190 6916
rect 2457 7208 2509 7218
rect 2457 7174 2466 7208
rect 2466 7174 2500 7208
rect 2500 7174 2509 7208
rect 2457 7166 2509 7174
rect 2650 7208 2702 7218
rect 2650 7174 2658 7208
rect 2658 7174 2692 7208
rect 2692 7174 2702 7208
rect 2650 7166 2702 7174
rect 2841 7208 2893 7218
rect 2841 7174 2850 7208
rect 2850 7174 2884 7208
rect 2884 7174 2893 7208
rect 2841 7166 2893 7174
rect 3033 7208 3085 7218
rect 3033 7174 3042 7208
rect 3042 7174 3076 7208
rect 3076 7174 3085 7208
rect 3033 7166 3085 7174
rect 3225 7208 3277 7218
rect 3225 7174 3234 7208
rect 3234 7174 3268 7208
rect 3268 7174 3277 7208
rect 3225 7166 3277 7174
rect 3417 7208 3469 7218
rect 3417 7174 3426 7208
rect 3426 7174 3460 7208
rect 3460 7174 3469 7208
rect 3417 7166 3469 7174
rect 1608 6448 1720 6572
rect 304 6396 356 6407
rect 304 6362 313 6396
rect 313 6362 347 6396
rect 347 6362 356 6396
rect 304 6355 356 6362
rect 495 6396 547 6407
rect 495 6362 505 6396
rect 505 6362 539 6396
rect 539 6362 547 6396
rect 495 6355 547 6362
rect 687 6396 739 6407
rect 687 6362 697 6396
rect 697 6362 731 6396
rect 731 6362 739 6396
rect 687 6355 739 6362
rect 879 6396 931 6407
rect 879 6362 889 6396
rect 889 6362 923 6396
rect 923 6362 931 6396
rect 879 6355 931 6362
rect 1072 6396 1124 6406
rect 1072 6362 1081 6396
rect 1081 6362 1115 6396
rect 1115 6362 1124 6396
rect 1072 6354 1124 6362
rect 1264 6396 1316 6406
rect 1264 6362 1273 6396
rect 1273 6362 1307 6396
rect 1307 6362 1316 6396
rect 1264 6354 1316 6362
rect 1468 6354 1524 6410
rect 1930 6356 1986 6412
rect 3978 7208 4030 7218
rect 3978 7174 3987 7208
rect 3987 7174 4021 7208
rect 4021 7174 4030 7208
rect 3978 7166 4030 7174
rect 4171 7208 4223 7218
rect 4171 7174 4179 7208
rect 4179 7174 4213 7208
rect 4213 7174 4223 7208
rect 4171 7166 4223 7174
rect 4362 7208 4414 7218
rect 4362 7174 4371 7208
rect 4371 7174 4405 7208
rect 4405 7174 4414 7208
rect 4362 7166 4414 7174
rect 4554 7208 4606 7218
rect 4554 7174 4563 7208
rect 4563 7174 4597 7208
rect 4597 7174 4606 7208
rect 4554 7166 4606 7174
rect 4746 7208 4798 7218
rect 4746 7174 4755 7208
rect 4755 7174 4789 7208
rect 4789 7174 4798 7208
rect 4746 7166 4798 7174
rect 4938 7208 4990 7218
rect 4938 7174 4947 7208
rect 4947 7174 4981 7208
rect 4981 7174 4990 7208
rect 4938 7166 4990 7174
rect 3681 6622 3733 6641
rect 3681 6589 3691 6622
rect 3691 6589 3725 6622
rect 3725 6589 3733 6622
rect 5337 6663 5389 6673
rect 5337 6629 5348 6663
rect 5348 6629 5382 6663
rect 5382 6629 5389 6663
rect 5337 6621 5389 6629
rect 5449 6668 5501 6675
rect 5449 6634 5450 6668
rect 5450 6634 5484 6668
rect 5484 6634 5501 6668
rect 5449 6623 5501 6634
rect 2457 6400 2509 6411
rect 2457 6366 2466 6400
rect 2466 6366 2500 6400
rect 2500 6366 2509 6400
rect 2457 6359 2509 6366
rect 2648 6400 2700 6411
rect 2648 6366 2658 6400
rect 2658 6366 2692 6400
rect 2692 6366 2700 6400
rect 2648 6359 2700 6366
rect 2840 6400 2892 6411
rect 2840 6366 2850 6400
rect 2850 6366 2884 6400
rect 2884 6366 2892 6400
rect 2840 6359 2892 6366
rect 3032 6400 3084 6411
rect 3032 6366 3042 6400
rect 3042 6366 3076 6400
rect 3076 6366 3084 6400
rect 3032 6359 3084 6366
rect 3225 6400 3277 6410
rect 3225 6366 3234 6400
rect 3234 6366 3268 6400
rect 3268 6366 3277 6400
rect 3225 6358 3277 6366
rect 3417 6400 3469 6410
rect 3417 6366 3426 6400
rect 3426 6366 3460 6400
rect 3460 6366 3469 6400
rect 3417 6358 3469 6366
rect 3978 6400 4030 6411
rect 3978 6366 3987 6400
rect 3987 6366 4021 6400
rect 4021 6366 4030 6400
rect 3978 6359 4030 6366
rect 4169 6400 4221 6411
rect 4169 6366 4179 6400
rect 4179 6366 4213 6400
rect 4213 6366 4221 6400
rect 4169 6359 4221 6366
rect 4361 6400 4413 6411
rect 4361 6366 4371 6400
rect 4371 6366 4405 6400
rect 4405 6366 4413 6400
rect 4361 6359 4413 6366
rect 4553 6400 4605 6411
rect 4553 6366 4563 6400
rect 4563 6366 4597 6400
rect 4597 6366 4605 6400
rect 4553 6359 4605 6366
rect 4746 6400 4798 6410
rect 4746 6366 4755 6400
rect 4755 6366 4789 6400
rect 4789 6366 4798 6400
rect 4746 6358 4798 6366
rect 4938 6400 4990 6410
rect 4938 6366 4947 6400
rect 4947 6366 4981 6400
rect 4981 6366 4990 6400
rect 4938 6358 4990 6366
rect 304 5917 356 5927
rect 304 5883 313 5917
rect 313 5883 347 5917
rect 347 5883 356 5917
rect 304 5875 356 5883
rect 497 5917 549 5927
rect 497 5883 505 5917
rect 505 5883 539 5917
rect 539 5883 549 5917
rect 497 5875 549 5883
rect 688 5917 740 5927
rect 688 5883 697 5917
rect 697 5883 731 5917
rect 731 5883 740 5917
rect 688 5875 740 5883
rect 880 5917 932 5927
rect 880 5883 889 5917
rect 889 5883 923 5917
rect 923 5883 932 5917
rect 880 5875 932 5883
rect 1072 5917 1124 5927
rect 1072 5883 1081 5917
rect 1081 5883 1115 5917
rect 1115 5883 1124 5917
rect 1072 5875 1124 5883
rect 1264 5917 1316 5927
rect 1264 5883 1273 5917
rect 1273 5883 1307 5917
rect 1307 5883 1316 5917
rect 1264 5875 1316 5883
rect 1522 5868 1578 5928
rect 1792 5868 1852 5928
rect 2056 5521 2190 5629
rect 2457 5921 2509 5931
rect 2457 5887 2466 5921
rect 2466 5887 2500 5921
rect 2500 5887 2509 5921
rect 2457 5879 2509 5887
rect 2650 5921 2702 5931
rect 2650 5887 2658 5921
rect 2658 5887 2692 5921
rect 2692 5887 2702 5921
rect 2650 5879 2702 5887
rect 2841 5921 2893 5931
rect 2841 5887 2850 5921
rect 2850 5887 2884 5921
rect 2884 5887 2893 5921
rect 2841 5879 2893 5887
rect 3033 5921 3085 5931
rect 3033 5887 3042 5921
rect 3042 5887 3076 5921
rect 3076 5887 3085 5921
rect 3033 5879 3085 5887
rect 3225 5921 3277 5931
rect 3225 5887 3234 5921
rect 3234 5887 3268 5921
rect 3268 5887 3277 5921
rect 3225 5879 3277 5887
rect 3417 5921 3469 5931
rect 3417 5887 3426 5921
rect 3426 5887 3460 5921
rect 3460 5887 3469 5921
rect 3417 5879 3469 5887
rect 1608 5161 1720 5285
rect 304 5109 356 5120
rect 304 5075 313 5109
rect 313 5075 347 5109
rect 347 5075 356 5109
rect 304 5068 356 5075
rect 495 5109 547 5120
rect 495 5075 505 5109
rect 505 5075 539 5109
rect 539 5075 547 5109
rect 495 5068 547 5075
rect 687 5109 739 5120
rect 687 5075 697 5109
rect 697 5075 731 5109
rect 731 5075 739 5109
rect 687 5068 739 5075
rect 879 5109 931 5120
rect 879 5075 889 5109
rect 889 5075 923 5109
rect 923 5075 931 5109
rect 879 5068 931 5075
rect 1072 5109 1124 5119
rect 1072 5075 1081 5109
rect 1081 5075 1115 5109
rect 1115 5075 1124 5109
rect 1072 5067 1124 5075
rect 1264 5109 1316 5119
rect 1264 5075 1273 5109
rect 1273 5075 1307 5109
rect 1307 5075 1316 5109
rect 1264 5067 1316 5075
rect 1468 5067 1524 5123
rect 1930 5069 1986 5125
rect 3978 5921 4030 5931
rect 3978 5887 3987 5921
rect 3987 5887 4021 5921
rect 4021 5887 4030 5921
rect 3978 5879 4030 5887
rect 4171 5921 4223 5931
rect 4171 5887 4179 5921
rect 4179 5887 4213 5921
rect 4213 5887 4223 5921
rect 4171 5879 4223 5887
rect 4362 5921 4414 5931
rect 4362 5887 4371 5921
rect 4371 5887 4405 5921
rect 4405 5887 4414 5921
rect 4362 5879 4414 5887
rect 4554 5921 4606 5931
rect 4554 5887 4563 5921
rect 4563 5887 4597 5921
rect 4597 5887 4606 5921
rect 4554 5879 4606 5887
rect 4746 5921 4798 5931
rect 4746 5887 4755 5921
rect 4755 5887 4789 5921
rect 4789 5887 4798 5921
rect 4746 5879 4798 5887
rect 4938 5921 4990 5931
rect 4938 5887 4947 5921
rect 4947 5887 4981 5921
rect 4981 5887 4990 5921
rect 4938 5879 4990 5887
rect 3681 5335 3733 5354
rect 3681 5302 3691 5335
rect 3691 5302 3725 5335
rect 3725 5302 3733 5335
rect 5337 5376 5389 5386
rect 5337 5342 5348 5376
rect 5348 5342 5382 5376
rect 5382 5342 5389 5376
rect 5337 5334 5389 5342
rect 5449 5381 5501 5388
rect 5449 5347 5450 5381
rect 5450 5347 5484 5381
rect 5484 5347 5501 5381
rect 5449 5336 5501 5347
rect 2457 5113 2509 5124
rect 2457 5079 2466 5113
rect 2466 5079 2500 5113
rect 2500 5079 2509 5113
rect 2457 5072 2509 5079
rect 2648 5113 2700 5124
rect 2648 5079 2658 5113
rect 2658 5079 2692 5113
rect 2692 5079 2700 5113
rect 2648 5072 2700 5079
rect 2840 5113 2892 5124
rect 2840 5079 2850 5113
rect 2850 5079 2884 5113
rect 2884 5079 2892 5113
rect 2840 5072 2892 5079
rect 3032 5113 3084 5124
rect 3032 5079 3042 5113
rect 3042 5079 3076 5113
rect 3076 5079 3084 5113
rect 3032 5072 3084 5079
rect 3225 5113 3277 5123
rect 3225 5079 3234 5113
rect 3234 5079 3268 5113
rect 3268 5079 3277 5113
rect 3225 5071 3277 5079
rect 3417 5113 3469 5123
rect 3417 5079 3426 5113
rect 3426 5079 3460 5113
rect 3460 5079 3469 5113
rect 3417 5071 3469 5079
rect 3978 5113 4030 5124
rect 3978 5079 3987 5113
rect 3987 5079 4021 5113
rect 4021 5079 4030 5113
rect 3978 5072 4030 5079
rect 4169 5113 4221 5124
rect 4169 5079 4179 5113
rect 4179 5079 4213 5113
rect 4213 5079 4221 5113
rect 4169 5072 4221 5079
rect 4361 5113 4413 5124
rect 4361 5079 4371 5113
rect 4371 5079 4405 5113
rect 4405 5079 4413 5113
rect 4361 5072 4413 5079
rect 4553 5113 4605 5124
rect 4553 5079 4563 5113
rect 4563 5079 4597 5113
rect 4597 5079 4605 5113
rect 4553 5072 4605 5079
rect 4746 5113 4798 5123
rect 4746 5079 4755 5113
rect 4755 5079 4789 5113
rect 4789 5079 4798 5113
rect 4746 5071 4798 5079
rect 4938 5113 4990 5123
rect 4938 5079 4947 5113
rect 4947 5079 4981 5113
rect 4981 5079 4990 5113
rect 4938 5071 4990 5079
rect 304 4630 356 4640
rect 304 4596 313 4630
rect 313 4596 347 4630
rect 347 4596 356 4630
rect 304 4588 356 4596
rect 497 4630 549 4640
rect 497 4596 505 4630
rect 505 4596 539 4630
rect 539 4596 549 4630
rect 497 4588 549 4596
rect 688 4630 740 4640
rect 688 4596 697 4630
rect 697 4596 731 4630
rect 731 4596 740 4630
rect 688 4588 740 4596
rect 880 4630 932 4640
rect 880 4596 889 4630
rect 889 4596 923 4630
rect 923 4596 932 4630
rect 880 4588 932 4596
rect 1072 4630 1124 4640
rect 1072 4596 1081 4630
rect 1081 4596 1115 4630
rect 1115 4596 1124 4630
rect 1072 4588 1124 4596
rect 1264 4630 1316 4640
rect 1264 4596 1273 4630
rect 1273 4596 1307 4630
rect 1307 4596 1316 4630
rect 1264 4588 1316 4596
rect 1522 4581 1578 4641
rect 1792 4581 1852 4641
rect 2056 4234 2190 4342
rect 2457 4634 2509 4644
rect 2457 4600 2466 4634
rect 2466 4600 2500 4634
rect 2500 4600 2509 4634
rect 2457 4592 2509 4600
rect 2650 4634 2702 4644
rect 2650 4600 2658 4634
rect 2658 4600 2692 4634
rect 2692 4600 2702 4634
rect 2650 4592 2702 4600
rect 2841 4634 2893 4644
rect 2841 4600 2850 4634
rect 2850 4600 2884 4634
rect 2884 4600 2893 4634
rect 2841 4592 2893 4600
rect 3033 4634 3085 4644
rect 3033 4600 3042 4634
rect 3042 4600 3076 4634
rect 3076 4600 3085 4634
rect 3033 4592 3085 4600
rect 3225 4634 3277 4644
rect 3225 4600 3234 4634
rect 3234 4600 3268 4634
rect 3268 4600 3277 4634
rect 3225 4592 3277 4600
rect 3417 4634 3469 4644
rect 3417 4600 3426 4634
rect 3426 4600 3460 4634
rect 3460 4600 3469 4634
rect 3417 4592 3469 4600
rect 1608 3874 1720 3998
rect 304 3822 356 3833
rect 304 3788 313 3822
rect 313 3788 347 3822
rect 347 3788 356 3822
rect 304 3781 356 3788
rect 495 3822 547 3833
rect 495 3788 505 3822
rect 505 3788 539 3822
rect 539 3788 547 3822
rect 495 3781 547 3788
rect 687 3822 739 3833
rect 687 3788 697 3822
rect 697 3788 731 3822
rect 731 3788 739 3822
rect 687 3781 739 3788
rect 879 3822 931 3833
rect 879 3788 889 3822
rect 889 3788 923 3822
rect 923 3788 931 3822
rect 879 3781 931 3788
rect 1072 3822 1124 3832
rect 1072 3788 1081 3822
rect 1081 3788 1115 3822
rect 1115 3788 1124 3822
rect 1072 3780 1124 3788
rect 1264 3822 1316 3832
rect 1264 3788 1273 3822
rect 1273 3788 1307 3822
rect 1307 3788 1316 3822
rect 1264 3780 1316 3788
rect 1468 3780 1524 3836
rect 1930 3782 1986 3838
rect 3978 4634 4030 4644
rect 3978 4600 3987 4634
rect 3987 4600 4021 4634
rect 4021 4600 4030 4634
rect 3978 4592 4030 4600
rect 4171 4634 4223 4644
rect 4171 4600 4179 4634
rect 4179 4600 4213 4634
rect 4213 4600 4223 4634
rect 4171 4592 4223 4600
rect 4362 4634 4414 4644
rect 4362 4600 4371 4634
rect 4371 4600 4405 4634
rect 4405 4600 4414 4634
rect 4362 4592 4414 4600
rect 4554 4634 4606 4644
rect 4554 4600 4563 4634
rect 4563 4600 4597 4634
rect 4597 4600 4606 4634
rect 4554 4592 4606 4600
rect 4746 4634 4798 4644
rect 4746 4600 4755 4634
rect 4755 4600 4789 4634
rect 4789 4600 4798 4634
rect 4746 4592 4798 4600
rect 4938 4634 4990 4644
rect 4938 4600 4947 4634
rect 4947 4600 4981 4634
rect 4981 4600 4990 4634
rect 4938 4592 4990 4600
rect 3681 4048 3733 4067
rect 3681 4015 3691 4048
rect 3691 4015 3725 4048
rect 3725 4015 3733 4048
rect 5337 4089 5389 4099
rect 5337 4055 5348 4089
rect 5348 4055 5382 4089
rect 5382 4055 5389 4089
rect 5337 4047 5389 4055
rect 5449 4094 5501 4101
rect 5449 4060 5450 4094
rect 5450 4060 5484 4094
rect 5484 4060 5501 4094
rect 5449 4049 5501 4060
rect 2457 3826 2509 3837
rect 2457 3792 2466 3826
rect 2466 3792 2500 3826
rect 2500 3792 2509 3826
rect 2457 3785 2509 3792
rect 2648 3826 2700 3837
rect 2648 3792 2658 3826
rect 2658 3792 2692 3826
rect 2692 3792 2700 3826
rect 2648 3785 2700 3792
rect 2840 3826 2892 3837
rect 2840 3792 2850 3826
rect 2850 3792 2884 3826
rect 2884 3792 2892 3826
rect 2840 3785 2892 3792
rect 3032 3826 3084 3837
rect 3032 3792 3042 3826
rect 3042 3792 3076 3826
rect 3076 3792 3084 3826
rect 3032 3785 3084 3792
rect 3225 3826 3277 3836
rect 3225 3792 3234 3826
rect 3234 3792 3268 3826
rect 3268 3792 3277 3826
rect 3225 3784 3277 3792
rect 3417 3826 3469 3836
rect 3417 3792 3426 3826
rect 3426 3792 3460 3826
rect 3460 3792 3469 3826
rect 3417 3784 3469 3792
rect 3978 3826 4030 3837
rect 3978 3792 3987 3826
rect 3987 3792 4021 3826
rect 4021 3792 4030 3826
rect 3978 3785 4030 3792
rect 4169 3826 4221 3837
rect 4169 3792 4179 3826
rect 4179 3792 4213 3826
rect 4213 3792 4221 3826
rect 4169 3785 4221 3792
rect 4361 3826 4413 3837
rect 4361 3792 4371 3826
rect 4371 3792 4405 3826
rect 4405 3792 4413 3826
rect 4361 3785 4413 3792
rect 4553 3826 4605 3837
rect 4553 3792 4563 3826
rect 4563 3792 4597 3826
rect 4597 3792 4605 3826
rect 4553 3785 4605 3792
rect 4746 3826 4798 3836
rect 4746 3792 4755 3826
rect 4755 3792 4789 3826
rect 4789 3792 4798 3826
rect 4746 3784 4798 3792
rect 4938 3826 4990 3836
rect 4938 3792 4947 3826
rect 4947 3792 4981 3826
rect 4981 3792 4990 3826
rect 4938 3784 4990 3792
rect 304 3343 356 3353
rect 304 3309 313 3343
rect 313 3309 347 3343
rect 347 3309 356 3343
rect 304 3301 356 3309
rect 497 3343 549 3353
rect 497 3309 505 3343
rect 505 3309 539 3343
rect 539 3309 549 3343
rect 497 3301 549 3309
rect 688 3343 740 3353
rect 688 3309 697 3343
rect 697 3309 731 3343
rect 731 3309 740 3343
rect 688 3301 740 3309
rect 880 3343 932 3353
rect 880 3309 889 3343
rect 889 3309 923 3343
rect 923 3309 932 3343
rect 880 3301 932 3309
rect 1072 3343 1124 3353
rect 1072 3309 1081 3343
rect 1081 3309 1115 3343
rect 1115 3309 1124 3343
rect 1072 3301 1124 3309
rect 1264 3343 1316 3353
rect 1264 3309 1273 3343
rect 1273 3309 1307 3343
rect 1307 3309 1316 3343
rect 1264 3301 1316 3309
rect 1522 3294 1578 3354
rect 1792 3294 1852 3354
rect 2056 2947 2190 3055
rect 2457 3347 2509 3357
rect 2457 3313 2466 3347
rect 2466 3313 2500 3347
rect 2500 3313 2509 3347
rect 2457 3305 2509 3313
rect 2650 3347 2702 3357
rect 2650 3313 2658 3347
rect 2658 3313 2692 3347
rect 2692 3313 2702 3347
rect 2650 3305 2702 3313
rect 2841 3347 2893 3357
rect 2841 3313 2850 3347
rect 2850 3313 2884 3347
rect 2884 3313 2893 3347
rect 2841 3305 2893 3313
rect 3033 3347 3085 3357
rect 3033 3313 3042 3347
rect 3042 3313 3076 3347
rect 3076 3313 3085 3347
rect 3033 3305 3085 3313
rect 3225 3347 3277 3357
rect 3225 3313 3234 3347
rect 3234 3313 3268 3347
rect 3268 3313 3277 3347
rect 3225 3305 3277 3313
rect 3417 3347 3469 3357
rect 3417 3313 3426 3347
rect 3426 3313 3460 3347
rect 3460 3313 3469 3347
rect 3417 3305 3469 3313
rect 1608 2587 1720 2711
rect 304 2535 356 2546
rect 304 2501 313 2535
rect 313 2501 347 2535
rect 347 2501 356 2535
rect 304 2494 356 2501
rect 495 2535 547 2546
rect 495 2501 505 2535
rect 505 2501 539 2535
rect 539 2501 547 2535
rect 495 2494 547 2501
rect 687 2535 739 2546
rect 687 2501 697 2535
rect 697 2501 731 2535
rect 731 2501 739 2535
rect 687 2494 739 2501
rect 879 2535 931 2546
rect 879 2501 889 2535
rect 889 2501 923 2535
rect 923 2501 931 2535
rect 879 2494 931 2501
rect 1072 2535 1124 2545
rect 1072 2501 1081 2535
rect 1081 2501 1115 2535
rect 1115 2501 1124 2535
rect 1072 2493 1124 2501
rect 1264 2535 1316 2545
rect 1264 2501 1273 2535
rect 1273 2501 1307 2535
rect 1307 2501 1316 2535
rect 1264 2493 1316 2501
rect 1468 2493 1524 2549
rect 1930 2495 1986 2551
rect 3978 3347 4030 3357
rect 3978 3313 3987 3347
rect 3987 3313 4021 3347
rect 4021 3313 4030 3347
rect 3978 3305 4030 3313
rect 4171 3347 4223 3357
rect 4171 3313 4179 3347
rect 4179 3313 4213 3347
rect 4213 3313 4223 3347
rect 4171 3305 4223 3313
rect 4362 3347 4414 3357
rect 4362 3313 4371 3347
rect 4371 3313 4405 3347
rect 4405 3313 4414 3347
rect 4362 3305 4414 3313
rect 4554 3347 4606 3357
rect 4554 3313 4563 3347
rect 4563 3313 4597 3347
rect 4597 3313 4606 3347
rect 4554 3305 4606 3313
rect 4746 3347 4798 3357
rect 4746 3313 4755 3347
rect 4755 3313 4789 3347
rect 4789 3313 4798 3347
rect 4746 3305 4798 3313
rect 4938 3347 4990 3357
rect 4938 3313 4947 3347
rect 4947 3313 4981 3347
rect 4981 3313 4990 3347
rect 4938 3305 4990 3313
rect 3681 2761 3733 2780
rect 3681 2728 3691 2761
rect 3691 2728 3725 2761
rect 3725 2728 3733 2761
rect 5337 2802 5389 2812
rect 5337 2768 5348 2802
rect 5348 2768 5382 2802
rect 5382 2768 5389 2802
rect 5337 2760 5389 2768
rect 5449 2807 5501 2814
rect 5449 2773 5450 2807
rect 5450 2773 5484 2807
rect 5484 2773 5501 2807
rect 5449 2762 5501 2773
rect 2457 2539 2509 2550
rect 2457 2505 2466 2539
rect 2466 2505 2500 2539
rect 2500 2505 2509 2539
rect 2457 2498 2509 2505
rect 2648 2539 2700 2550
rect 2648 2505 2658 2539
rect 2658 2505 2692 2539
rect 2692 2505 2700 2539
rect 2648 2498 2700 2505
rect 2840 2539 2892 2550
rect 2840 2505 2850 2539
rect 2850 2505 2884 2539
rect 2884 2505 2892 2539
rect 2840 2498 2892 2505
rect 3032 2539 3084 2550
rect 3032 2505 3042 2539
rect 3042 2505 3076 2539
rect 3076 2505 3084 2539
rect 3032 2498 3084 2505
rect 3225 2539 3277 2549
rect 3225 2505 3234 2539
rect 3234 2505 3268 2539
rect 3268 2505 3277 2539
rect 3225 2497 3277 2505
rect 3417 2539 3469 2549
rect 3417 2505 3426 2539
rect 3426 2505 3460 2539
rect 3460 2505 3469 2539
rect 3417 2497 3469 2505
rect 3978 2539 4030 2550
rect 3978 2505 3987 2539
rect 3987 2505 4021 2539
rect 4021 2505 4030 2539
rect 3978 2498 4030 2505
rect 4169 2539 4221 2550
rect 4169 2505 4179 2539
rect 4179 2505 4213 2539
rect 4213 2505 4221 2539
rect 4169 2498 4221 2505
rect 4361 2539 4413 2550
rect 4361 2505 4371 2539
rect 4371 2505 4405 2539
rect 4405 2505 4413 2539
rect 4361 2498 4413 2505
rect 4553 2539 4605 2550
rect 4553 2505 4563 2539
rect 4563 2505 4597 2539
rect 4597 2505 4605 2539
rect 4553 2498 4605 2505
rect 4746 2539 4798 2549
rect 4746 2505 4755 2539
rect 4755 2505 4789 2539
rect 4789 2505 4798 2539
rect 4746 2497 4798 2505
rect 4938 2539 4990 2549
rect 4938 2505 4947 2539
rect 4947 2505 4981 2539
rect 4981 2505 4990 2539
rect 4938 2497 4990 2505
rect 304 2056 356 2066
rect 304 2022 313 2056
rect 313 2022 347 2056
rect 347 2022 356 2056
rect 304 2014 356 2022
rect 497 2056 549 2066
rect 497 2022 505 2056
rect 505 2022 539 2056
rect 539 2022 549 2056
rect 497 2014 549 2022
rect 688 2056 740 2066
rect 688 2022 697 2056
rect 697 2022 731 2056
rect 731 2022 740 2056
rect 688 2014 740 2022
rect 880 2056 932 2066
rect 880 2022 889 2056
rect 889 2022 923 2056
rect 923 2022 932 2056
rect 880 2014 932 2022
rect 1072 2056 1124 2066
rect 1072 2022 1081 2056
rect 1081 2022 1115 2056
rect 1115 2022 1124 2056
rect 1072 2014 1124 2022
rect 1264 2056 1316 2066
rect 1264 2022 1273 2056
rect 1273 2022 1307 2056
rect 1307 2022 1316 2056
rect 1264 2014 1316 2022
rect 1522 2007 1578 2067
rect 1792 2007 1852 2067
rect 2056 1660 2190 1768
rect 2457 2060 2509 2070
rect 2457 2026 2466 2060
rect 2466 2026 2500 2060
rect 2500 2026 2509 2060
rect 2457 2018 2509 2026
rect 2650 2060 2702 2070
rect 2650 2026 2658 2060
rect 2658 2026 2692 2060
rect 2692 2026 2702 2060
rect 2650 2018 2702 2026
rect 2841 2060 2893 2070
rect 2841 2026 2850 2060
rect 2850 2026 2884 2060
rect 2884 2026 2893 2060
rect 2841 2018 2893 2026
rect 3033 2060 3085 2070
rect 3033 2026 3042 2060
rect 3042 2026 3076 2060
rect 3076 2026 3085 2060
rect 3033 2018 3085 2026
rect 3225 2060 3277 2070
rect 3225 2026 3234 2060
rect 3234 2026 3268 2060
rect 3268 2026 3277 2060
rect 3225 2018 3277 2026
rect 3417 2060 3469 2070
rect 3417 2026 3426 2060
rect 3426 2026 3460 2060
rect 3460 2026 3469 2060
rect 3417 2018 3469 2026
rect 1608 1300 1720 1424
rect 304 1248 356 1259
rect 304 1214 313 1248
rect 313 1214 347 1248
rect 347 1214 356 1248
rect 304 1207 356 1214
rect 495 1248 547 1259
rect 495 1214 505 1248
rect 505 1214 539 1248
rect 539 1214 547 1248
rect 495 1207 547 1214
rect 687 1248 739 1259
rect 687 1214 697 1248
rect 697 1214 731 1248
rect 731 1214 739 1248
rect 687 1207 739 1214
rect 879 1248 931 1259
rect 879 1214 889 1248
rect 889 1214 923 1248
rect 923 1214 931 1248
rect 879 1207 931 1214
rect 1072 1248 1124 1258
rect 1072 1214 1081 1248
rect 1081 1214 1115 1248
rect 1115 1214 1124 1248
rect 1072 1206 1124 1214
rect 1264 1248 1316 1258
rect 1264 1214 1273 1248
rect 1273 1214 1307 1248
rect 1307 1214 1316 1248
rect 1264 1206 1316 1214
rect 1468 1206 1524 1262
rect 1930 1208 1986 1264
rect 3978 2060 4030 2070
rect 3978 2026 3987 2060
rect 3987 2026 4021 2060
rect 4021 2026 4030 2060
rect 3978 2018 4030 2026
rect 4171 2060 4223 2070
rect 4171 2026 4179 2060
rect 4179 2026 4213 2060
rect 4213 2026 4223 2060
rect 4171 2018 4223 2026
rect 4362 2060 4414 2070
rect 4362 2026 4371 2060
rect 4371 2026 4405 2060
rect 4405 2026 4414 2060
rect 4362 2018 4414 2026
rect 4554 2060 4606 2070
rect 4554 2026 4563 2060
rect 4563 2026 4597 2060
rect 4597 2026 4606 2060
rect 4554 2018 4606 2026
rect 4746 2060 4798 2070
rect 4746 2026 4755 2060
rect 4755 2026 4789 2060
rect 4789 2026 4798 2060
rect 4746 2018 4798 2026
rect 4938 2060 4990 2070
rect 4938 2026 4947 2060
rect 4947 2026 4981 2060
rect 4981 2026 4990 2060
rect 4938 2018 4990 2026
rect 3681 1474 3733 1493
rect 3681 1441 3691 1474
rect 3691 1441 3725 1474
rect 3725 1441 3733 1474
rect 5337 1515 5389 1525
rect 5337 1481 5348 1515
rect 5348 1481 5382 1515
rect 5382 1481 5389 1515
rect 5337 1473 5389 1481
rect 5449 1520 5501 1527
rect 5449 1486 5450 1520
rect 5450 1486 5484 1520
rect 5484 1486 5501 1520
rect 5449 1475 5501 1486
rect 2457 1252 2509 1263
rect 2457 1218 2466 1252
rect 2466 1218 2500 1252
rect 2500 1218 2509 1252
rect 2457 1211 2509 1218
rect 2648 1252 2700 1263
rect 2648 1218 2658 1252
rect 2658 1218 2692 1252
rect 2692 1218 2700 1252
rect 2648 1211 2700 1218
rect 2840 1252 2892 1263
rect 2840 1218 2850 1252
rect 2850 1218 2884 1252
rect 2884 1218 2892 1252
rect 2840 1211 2892 1218
rect 3032 1252 3084 1263
rect 3032 1218 3042 1252
rect 3042 1218 3076 1252
rect 3076 1218 3084 1252
rect 3032 1211 3084 1218
rect 3225 1252 3277 1262
rect 3225 1218 3234 1252
rect 3234 1218 3268 1252
rect 3268 1218 3277 1252
rect 3225 1210 3277 1218
rect 3417 1252 3469 1262
rect 3417 1218 3426 1252
rect 3426 1218 3460 1252
rect 3460 1218 3469 1252
rect 3417 1210 3469 1218
rect 3978 1252 4030 1263
rect 3978 1218 3987 1252
rect 3987 1218 4021 1252
rect 4021 1218 4030 1252
rect 3978 1211 4030 1218
rect 4169 1252 4221 1263
rect 4169 1218 4179 1252
rect 4179 1218 4213 1252
rect 4213 1218 4221 1252
rect 4169 1211 4221 1218
rect 4361 1252 4413 1263
rect 4361 1218 4371 1252
rect 4371 1218 4405 1252
rect 4405 1218 4413 1252
rect 4361 1211 4413 1218
rect 4553 1252 4605 1263
rect 4553 1218 4563 1252
rect 4563 1218 4597 1252
rect 4597 1218 4605 1252
rect 4553 1211 4605 1218
rect 4746 1252 4798 1262
rect 4746 1218 4755 1252
rect 4755 1218 4789 1252
rect 4789 1218 4798 1252
rect 4746 1210 4798 1218
rect 4938 1252 4990 1262
rect 4938 1218 4947 1252
rect 4947 1218 4981 1252
rect 4981 1218 4990 1252
rect 4938 1210 4990 1218
<< metal2 >>
rect 304 41963 356 41973
rect 497 41963 549 41973
rect 688 41963 740 41973
rect 880 41963 932 41973
rect 1072 41963 1124 41973
rect 1264 41963 1316 41973
rect 1522 41964 1578 41974
rect 96 41911 304 41963
rect 356 41911 497 41963
rect 549 41911 688 41963
rect 740 41911 880 41963
rect 932 41911 1072 41963
rect 1124 41911 1264 41963
rect 1316 41911 1522 41963
rect 304 41901 356 41911
rect 497 41901 549 41911
rect 688 41901 740 41911
rect 880 41901 932 41911
rect 1072 41901 1124 41911
rect 1264 41901 1316 41911
rect 1522 41894 1578 41904
rect 1610 41331 1722 42210
rect 1608 41321 1722 41331
rect 1720 41197 1722 41321
rect 1608 41187 1722 41197
rect 304 41156 356 41166
rect 495 41156 547 41166
rect 687 41156 739 41166
rect 879 41156 931 41166
rect 1072 41156 1124 41165
rect 1264 41156 1316 41165
rect 1468 41159 1524 41169
rect 96 41104 304 41156
rect 356 41104 495 41156
rect 547 41104 687 41156
rect 739 41104 879 41156
rect 931 41155 1468 41156
rect 931 41104 1072 41155
rect 304 41094 356 41104
rect 495 41094 547 41104
rect 687 41094 739 41104
rect 879 41094 931 41104
rect 1124 41104 1264 41155
rect 1072 41093 1124 41103
rect 1316 41104 1468 41155
rect 1264 41093 1316 41103
rect 1524 41104 1526 41156
rect 1468 41093 1524 41103
rect 304 40676 356 40686
rect 497 40676 549 40686
rect 688 40676 740 40686
rect 880 40676 932 40686
rect 1072 40676 1124 40686
rect 1264 40676 1316 40686
rect 1522 40677 1578 40687
rect 96 40624 304 40676
rect 356 40624 497 40676
rect 549 40624 688 40676
rect 740 40624 880 40676
rect 932 40624 1072 40676
rect 1124 40624 1264 40676
rect 1316 40624 1522 40676
rect 304 40614 356 40624
rect 497 40614 549 40624
rect 688 40614 740 40624
rect 880 40614 932 40624
rect 1072 40614 1124 40624
rect 1264 40614 1316 40624
rect 1522 40607 1578 40617
rect 1610 40044 1722 41187
rect 1608 40034 1722 40044
rect 1720 39910 1722 40034
rect 1608 39900 1722 39910
rect 304 39869 356 39879
rect 495 39869 547 39879
rect 687 39869 739 39879
rect 879 39869 931 39879
rect 1072 39869 1124 39878
rect 1264 39869 1316 39878
rect 1468 39872 1524 39882
rect 96 39817 304 39869
rect 356 39817 495 39869
rect 547 39817 687 39869
rect 739 39817 879 39869
rect 931 39868 1468 39869
rect 931 39817 1072 39868
rect 304 39807 356 39817
rect 495 39807 547 39817
rect 687 39807 739 39817
rect 879 39807 931 39817
rect 1124 39817 1264 39868
rect 1072 39806 1124 39816
rect 1316 39817 1468 39868
rect 1264 39806 1316 39816
rect 1524 39817 1526 39869
rect 1468 39806 1524 39816
rect 304 39389 356 39399
rect 497 39389 549 39399
rect 688 39389 740 39399
rect 880 39389 932 39399
rect 1072 39389 1124 39399
rect 1264 39389 1316 39399
rect 1522 39390 1578 39400
rect 96 39337 304 39389
rect 356 39337 497 39389
rect 549 39337 688 39389
rect 740 39337 880 39389
rect 932 39337 1072 39389
rect 1124 39337 1264 39389
rect 1316 39337 1522 39389
rect 304 39327 356 39337
rect 497 39327 549 39337
rect 688 39327 740 39337
rect 880 39327 932 39337
rect 1072 39327 1124 39337
rect 1264 39327 1316 39337
rect 1522 39320 1578 39330
rect 1610 38757 1722 39900
rect 1608 38747 1722 38757
rect 1720 38623 1722 38747
rect 1608 38613 1722 38623
rect 304 38582 356 38592
rect 495 38582 547 38592
rect 687 38582 739 38592
rect 879 38582 931 38592
rect 1072 38582 1124 38591
rect 1264 38582 1316 38591
rect 1468 38585 1524 38595
rect 96 38530 304 38582
rect 356 38530 495 38582
rect 547 38530 687 38582
rect 739 38530 879 38582
rect 931 38581 1468 38582
rect 931 38530 1072 38581
rect 304 38520 356 38530
rect 495 38520 547 38530
rect 687 38520 739 38530
rect 879 38520 931 38530
rect 1124 38530 1264 38581
rect 1072 38519 1124 38529
rect 1316 38530 1468 38581
rect 1264 38519 1316 38529
rect 1524 38530 1526 38582
rect 1468 38519 1524 38529
rect 304 38102 356 38112
rect 497 38102 549 38112
rect 688 38102 740 38112
rect 880 38102 932 38112
rect 1072 38102 1124 38112
rect 1264 38102 1316 38112
rect 1522 38103 1578 38113
rect 96 38050 304 38102
rect 356 38050 497 38102
rect 549 38050 688 38102
rect 740 38050 880 38102
rect 932 38050 1072 38102
rect 1124 38050 1264 38102
rect 1316 38050 1522 38102
rect 304 38040 356 38050
rect 497 38040 549 38050
rect 688 38040 740 38050
rect 880 38040 932 38050
rect 1072 38040 1124 38050
rect 1264 38040 1316 38050
rect 1522 38033 1578 38043
rect 1610 37470 1722 38613
rect 1608 37460 1722 37470
rect 1720 37336 1722 37460
rect 1608 37326 1722 37336
rect 304 37295 356 37305
rect 495 37295 547 37305
rect 687 37295 739 37305
rect 879 37295 931 37305
rect 1072 37295 1124 37304
rect 1264 37295 1316 37304
rect 1468 37298 1524 37308
rect 96 37243 304 37295
rect 356 37243 495 37295
rect 547 37243 687 37295
rect 739 37243 879 37295
rect 931 37294 1468 37295
rect 931 37243 1072 37294
rect 304 37233 356 37243
rect 495 37233 547 37243
rect 687 37233 739 37243
rect 879 37233 931 37243
rect 1124 37243 1264 37294
rect 1072 37232 1124 37242
rect 1316 37243 1468 37294
rect 1264 37232 1316 37242
rect 1524 37243 1526 37295
rect 1468 37232 1524 37242
rect 304 36815 356 36825
rect 497 36815 549 36825
rect 688 36815 740 36825
rect 880 36815 932 36825
rect 1072 36815 1124 36825
rect 1264 36815 1316 36825
rect 1522 36816 1578 36826
rect 96 36763 304 36815
rect 356 36763 497 36815
rect 549 36763 688 36815
rect 740 36763 880 36815
rect 932 36763 1072 36815
rect 1124 36763 1264 36815
rect 1316 36763 1522 36815
rect 304 36753 356 36763
rect 497 36753 549 36763
rect 688 36753 740 36763
rect 880 36753 932 36763
rect 1072 36753 1124 36763
rect 1264 36753 1316 36763
rect 1522 36746 1578 36756
rect 1610 36183 1722 37326
rect 1608 36173 1722 36183
rect 1720 36049 1722 36173
rect 1608 36039 1722 36049
rect 304 36008 356 36018
rect 495 36008 547 36018
rect 687 36008 739 36018
rect 879 36008 931 36018
rect 1072 36008 1124 36017
rect 1264 36008 1316 36017
rect 1468 36011 1524 36021
rect 96 35956 304 36008
rect 356 35956 495 36008
rect 547 35956 687 36008
rect 739 35956 879 36008
rect 931 36007 1468 36008
rect 931 35956 1072 36007
rect 304 35946 356 35956
rect 495 35946 547 35956
rect 687 35946 739 35956
rect 879 35946 931 35956
rect 1124 35956 1264 36007
rect 1072 35945 1124 35955
rect 1316 35956 1468 36007
rect 1264 35945 1316 35955
rect 1524 35956 1526 36008
rect 1468 35945 1524 35955
rect 304 35528 356 35538
rect 497 35528 549 35538
rect 688 35528 740 35538
rect 880 35528 932 35538
rect 1072 35528 1124 35538
rect 1264 35528 1316 35538
rect 1522 35529 1578 35539
rect 96 35476 304 35528
rect 356 35476 497 35528
rect 549 35476 688 35528
rect 740 35476 880 35528
rect 932 35476 1072 35528
rect 1124 35476 1264 35528
rect 1316 35476 1522 35528
rect 304 35466 356 35476
rect 497 35466 549 35476
rect 688 35466 740 35476
rect 880 35466 932 35476
rect 1072 35466 1124 35476
rect 1264 35466 1316 35476
rect 1522 35459 1578 35469
rect 1610 34896 1722 36039
rect 1608 34886 1722 34896
rect 1720 34762 1722 34886
rect 1608 34752 1722 34762
rect 304 34721 356 34731
rect 495 34721 547 34731
rect 687 34721 739 34731
rect 879 34721 931 34731
rect 1072 34721 1124 34730
rect 1264 34721 1316 34730
rect 1468 34724 1524 34734
rect 96 34669 304 34721
rect 356 34669 495 34721
rect 547 34669 687 34721
rect 739 34669 879 34721
rect 931 34720 1468 34721
rect 931 34669 1072 34720
rect 304 34659 356 34669
rect 495 34659 547 34669
rect 687 34659 739 34669
rect 879 34659 931 34669
rect 1124 34669 1264 34720
rect 1072 34658 1124 34668
rect 1316 34669 1468 34720
rect 1264 34658 1316 34668
rect 1524 34669 1526 34721
rect 1468 34658 1524 34668
rect 304 34241 356 34251
rect 497 34241 549 34251
rect 688 34241 740 34251
rect 880 34241 932 34251
rect 1072 34241 1124 34251
rect 1264 34241 1316 34251
rect 1522 34242 1578 34252
rect 96 34189 304 34241
rect 356 34189 497 34241
rect 549 34189 688 34241
rect 740 34189 880 34241
rect 932 34189 1072 34241
rect 1124 34189 1264 34241
rect 1316 34189 1522 34241
rect 304 34179 356 34189
rect 497 34179 549 34189
rect 688 34179 740 34189
rect 880 34179 932 34189
rect 1072 34179 1124 34189
rect 1264 34179 1316 34189
rect 1522 34172 1578 34182
rect 1610 33609 1722 34752
rect 1608 33599 1722 33609
rect 1720 33475 1722 33599
rect 1608 33465 1722 33475
rect 304 33434 356 33444
rect 495 33434 547 33444
rect 687 33434 739 33444
rect 879 33434 931 33444
rect 1072 33434 1124 33443
rect 1264 33434 1316 33443
rect 1468 33437 1524 33447
rect 96 33382 304 33434
rect 356 33382 495 33434
rect 547 33382 687 33434
rect 739 33382 879 33434
rect 931 33433 1468 33434
rect 931 33382 1072 33433
rect 304 33372 356 33382
rect 495 33372 547 33382
rect 687 33372 739 33382
rect 879 33372 931 33382
rect 1124 33382 1264 33433
rect 1072 33371 1124 33381
rect 1316 33382 1468 33433
rect 1264 33371 1316 33381
rect 1524 33382 1526 33434
rect 1468 33371 1524 33381
rect 304 32954 356 32964
rect 497 32954 549 32964
rect 688 32954 740 32964
rect 880 32954 932 32964
rect 1072 32954 1124 32964
rect 1264 32954 1316 32964
rect 1522 32955 1578 32965
rect 96 32902 304 32954
rect 356 32902 497 32954
rect 549 32902 688 32954
rect 740 32902 880 32954
rect 932 32902 1072 32954
rect 1124 32902 1264 32954
rect 1316 32902 1522 32954
rect 304 32892 356 32902
rect 497 32892 549 32902
rect 688 32892 740 32902
rect 880 32892 932 32902
rect 1072 32892 1124 32902
rect 1264 32892 1316 32902
rect 1522 32885 1578 32895
rect 1610 32322 1722 33465
rect 1608 32312 1722 32322
rect 1720 32188 1722 32312
rect 1608 32178 1722 32188
rect 304 32147 356 32157
rect 495 32147 547 32157
rect 687 32147 739 32157
rect 879 32147 931 32157
rect 1072 32147 1124 32156
rect 1264 32147 1316 32156
rect 1468 32150 1524 32160
rect 96 32095 304 32147
rect 356 32095 495 32147
rect 547 32095 687 32147
rect 739 32095 879 32147
rect 931 32146 1468 32147
rect 931 32095 1072 32146
rect 304 32085 356 32095
rect 495 32085 547 32095
rect 687 32085 739 32095
rect 879 32085 931 32095
rect 1124 32095 1264 32146
rect 1072 32084 1124 32094
rect 1316 32095 1468 32146
rect 1264 32084 1316 32094
rect 1524 32095 1526 32147
rect 1468 32084 1524 32094
rect 304 31667 356 31677
rect 497 31667 549 31677
rect 688 31667 740 31677
rect 880 31667 932 31677
rect 1072 31667 1124 31677
rect 1264 31667 1316 31677
rect 1522 31668 1578 31678
rect 96 31615 304 31667
rect 356 31615 497 31667
rect 549 31615 688 31667
rect 740 31615 880 31667
rect 932 31615 1072 31667
rect 1124 31615 1264 31667
rect 1316 31615 1522 31667
rect 304 31605 356 31615
rect 497 31605 549 31615
rect 688 31605 740 31615
rect 880 31605 932 31615
rect 1072 31605 1124 31615
rect 1264 31605 1316 31615
rect 1522 31598 1578 31608
rect 1610 31035 1722 32178
rect 1608 31025 1722 31035
rect 1720 30901 1722 31025
rect 1608 30891 1722 30901
rect 304 30860 356 30870
rect 495 30860 547 30870
rect 687 30860 739 30870
rect 879 30860 931 30870
rect 1072 30860 1124 30869
rect 1264 30860 1316 30869
rect 1468 30863 1524 30873
rect 96 30808 304 30860
rect 356 30808 495 30860
rect 547 30808 687 30860
rect 739 30808 879 30860
rect 931 30859 1468 30860
rect 931 30808 1072 30859
rect 304 30798 356 30808
rect 495 30798 547 30808
rect 687 30798 739 30808
rect 879 30798 931 30808
rect 1124 30808 1264 30859
rect 1072 30797 1124 30807
rect 1316 30808 1468 30859
rect 1264 30797 1316 30807
rect 1524 30808 1526 30860
rect 1468 30797 1524 30807
rect 304 30380 356 30390
rect 497 30380 549 30390
rect 688 30380 740 30390
rect 880 30380 932 30390
rect 1072 30380 1124 30390
rect 1264 30380 1316 30390
rect 1522 30381 1578 30391
rect 96 30328 304 30380
rect 356 30328 497 30380
rect 549 30328 688 30380
rect 740 30328 880 30380
rect 932 30328 1072 30380
rect 1124 30328 1264 30380
rect 1316 30328 1522 30380
rect 304 30318 356 30328
rect 497 30318 549 30328
rect 688 30318 740 30328
rect 880 30318 932 30328
rect 1072 30318 1124 30328
rect 1264 30318 1316 30328
rect 1522 30311 1578 30321
rect 1610 29748 1722 30891
rect 1608 29738 1722 29748
rect 1720 29614 1722 29738
rect 1608 29604 1722 29614
rect 304 29573 356 29583
rect 495 29573 547 29583
rect 687 29573 739 29583
rect 879 29573 931 29583
rect 1072 29573 1124 29582
rect 1264 29573 1316 29582
rect 1468 29576 1524 29586
rect 96 29521 304 29573
rect 356 29521 495 29573
rect 547 29521 687 29573
rect 739 29521 879 29573
rect 931 29572 1468 29573
rect 931 29521 1072 29572
rect 304 29511 356 29521
rect 495 29511 547 29521
rect 687 29511 739 29521
rect 879 29511 931 29521
rect 1124 29521 1264 29572
rect 1072 29510 1124 29520
rect 1316 29521 1468 29572
rect 1264 29510 1316 29520
rect 1524 29521 1526 29573
rect 1468 29510 1524 29520
rect 304 29093 356 29103
rect 497 29093 549 29103
rect 688 29093 740 29103
rect 880 29093 932 29103
rect 1072 29093 1124 29103
rect 1264 29093 1316 29103
rect 1522 29094 1578 29104
rect 96 29041 304 29093
rect 356 29041 497 29093
rect 549 29041 688 29093
rect 740 29041 880 29093
rect 932 29041 1072 29093
rect 1124 29041 1264 29093
rect 1316 29041 1522 29093
rect 304 29031 356 29041
rect 497 29031 549 29041
rect 688 29031 740 29041
rect 880 29031 932 29041
rect 1072 29031 1124 29041
rect 1264 29031 1316 29041
rect 1522 29024 1578 29034
rect 1610 28461 1722 29604
rect 1608 28451 1722 28461
rect 1720 28327 1722 28451
rect 1608 28317 1722 28327
rect 304 28286 356 28296
rect 495 28286 547 28296
rect 687 28286 739 28296
rect 879 28286 931 28296
rect 1072 28286 1124 28295
rect 1264 28286 1316 28295
rect 1468 28289 1524 28299
rect 96 28234 304 28286
rect 356 28234 495 28286
rect 547 28234 687 28286
rect 739 28234 879 28286
rect 931 28285 1468 28286
rect 931 28234 1072 28285
rect 304 28224 356 28234
rect 495 28224 547 28234
rect 687 28224 739 28234
rect 879 28224 931 28234
rect 1124 28234 1264 28285
rect 1072 28223 1124 28233
rect 1316 28234 1468 28285
rect 1264 28223 1316 28233
rect 1524 28234 1526 28286
rect 1468 28223 1524 28233
rect 304 27806 356 27816
rect 497 27806 549 27816
rect 688 27806 740 27816
rect 880 27806 932 27816
rect 1072 27806 1124 27816
rect 1264 27806 1316 27816
rect 1522 27807 1578 27817
rect 96 27754 304 27806
rect 356 27754 497 27806
rect 549 27754 688 27806
rect 740 27754 880 27806
rect 932 27754 1072 27806
rect 1124 27754 1264 27806
rect 1316 27754 1522 27806
rect 304 27744 356 27754
rect 497 27744 549 27754
rect 688 27744 740 27754
rect 880 27744 932 27754
rect 1072 27744 1124 27754
rect 1264 27744 1316 27754
rect 1522 27737 1578 27747
rect 1610 27174 1722 28317
rect 1608 27164 1722 27174
rect 1720 27040 1722 27164
rect 1608 27030 1722 27040
rect 304 26999 356 27009
rect 495 26999 547 27009
rect 687 26999 739 27009
rect 879 26999 931 27009
rect 1072 26999 1124 27008
rect 1264 26999 1316 27008
rect 1468 27002 1524 27012
rect 96 26947 304 26999
rect 356 26947 495 26999
rect 547 26947 687 26999
rect 739 26947 879 26999
rect 931 26998 1468 26999
rect 931 26947 1072 26998
rect 304 26937 356 26947
rect 495 26937 547 26947
rect 687 26937 739 26947
rect 879 26937 931 26947
rect 1124 26947 1264 26998
rect 1072 26936 1124 26946
rect 1316 26947 1468 26998
rect 1264 26936 1316 26946
rect 1524 26947 1526 26999
rect 1468 26936 1524 26946
rect 304 26519 356 26529
rect 497 26519 549 26529
rect 688 26519 740 26529
rect 880 26519 932 26529
rect 1072 26519 1124 26529
rect 1264 26519 1316 26529
rect 1522 26520 1578 26530
rect 96 26467 304 26519
rect 356 26467 497 26519
rect 549 26467 688 26519
rect 740 26467 880 26519
rect 932 26467 1072 26519
rect 1124 26467 1264 26519
rect 1316 26467 1522 26519
rect 304 26457 356 26467
rect 497 26457 549 26467
rect 688 26457 740 26467
rect 880 26457 932 26467
rect 1072 26457 1124 26467
rect 1264 26457 1316 26467
rect 1522 26450 1578 26460
rect 1610 25887 1722 27030
rect 1608 25877 1722 25887
rect 1720 25753 1722 25877
rect 1608 25743 1722 25753
rect 304 25712 356 25722
rect 495 25712 547 25722
rect 687 25712 739 25722
rect 879 25712 931 25722
rect 1072 25712 1124 25721
rect 1264 25712 1316 25721
rect 1468 25715 1524 25725
rect 96 25660 304 25712
rect 356 25660 495 25712
rect 547 25660 687 25712
rect 739 25660 879 25712
rect 931 25711 1468 25712
rect 931 25660 1072 25711
rect 304 25650 356 25660
rect 495 25650 547 25660
rect 687 25650 739 25660
rect 879 25650 931 25660
rect 1124 25660 1264 25711
rect 1072 25649 1124 25659
rect 1316 25660 1468 25711
rect 1264 25649 1316 25659
rect 1524 25660 1526 25712
rect 1468 25649 1524 25659
rect 304 25232 356 25242
rect 497 25232 549 25242
rect 688 25232 740 25242
rect 880 25232 932 25242
rect 1072 25232 1124 25242
rect 1264 25232 1316 25242
rect 1522 25233 1578 25243
rect 96 25180 304 25232
rect 356 25180 497 25232
rect 549 25180 688 25232
rect 740 25180 880 25232
rect 932 25180 1072 25232
rect 1124 25180 1264 25232
rect 1316 25180 1522 25232
rect 304 25170 356 25180
rect 497 25170 549 25180
rect 688 25170 740 25180
rect 880 25170 932 25180
rect 1072 25170 1124 25180
rect 1264 25170 1316 25180
rect 1522 25163 1578 25173
rect 1610 24600 1722 25743
rect 1608 24590 1722 24600
rect 1720 24466 1722 24590
rect 1608 24456 1722 24466
rect 304 24425 356 24435
rect 495 24425 547 24435
rect 687 24425 739 24435
rect 879 24425 931 24435
rect 1072 24425 1124 24434
rect 1264 24425 1316 24434
rect 1468 24428 1524 24438
rect 96 24373 304 24425
rect 356 24373 495 24425
rect 547 24373 687 24425
rect 739 24373 879 24425
rect 931 24424 1468 24425
rect 931 24373 1072 24424
rect 304 24363 356 24373
rect 495 24363 547 24373
rect 687 24363 739 24373
rect 879 24363 931 24373
rect 1124 24373 1264 24424
rect 1072 24362 1124 24372
rect 1316 24373 1468 24424
rect 1264 24362 1316 24372
rect 1524 24373 1526 24425
rect 1468 24362 1524 24372
rect 304 23945 356 23955
rect 497 23945 549 23955
rect 688 23945 740 23955
rect 880 23945 932 23955
rect 1072 23945 1124 23955
rect 1264 23945 1316 23955
rect 1522 23946 1578 23956
rect 96 23893 304 23945
rect 356 23893 497 23945
rect 549 23893 688 23945
rect 740 23893 880 23945
rect 932 23893 1072 23945
rect 1124 23893 1264 23945
rect 1316 23893 1522 23945
rect 304 23883 356 23893
rect 497 23883 549 23893
rect 688 23883 740 23893
rect 880 23883 932 23893
rect 1072 23883 1124 23893
rect 1264 23883 1316 23893
rect 1522 23876 1578 23886
rect 1610 23313 1722 24456
rect 1608 23303 1722 23313
rect 1720 23179 1722 23303
rect 1608 23169 1722 23179
rect 304 23138 356 23148
rect 495 23138 547 23148
rect 687 23138 739 23148
rect 879 23138 931 23148
rect 1072 23138 1124 23147
rect 1264 23138 1316 23147
rect 1468 23141 1524 23151
rect 96 23086 304 23138
rect 356 23086 495 23138
rect 547 23086 687 23138
rect 739 23086 879 23138
rect 931 23137 1468 23138
rect 931 23086 1072 23137
rect 304 23076 356 23086
rect 495 23076 547 23086
rect 687 23076 739 23086
rect 879 23076 931 23086
rect 1124 23086 1264 23137
rect 1072 23075 1124 23085
rect 1316 23086 1468 23137
rect 1264 23075 1316 23085
rect 1524 23086 1526 23138
rect 1468 23075 1524 23085
rect 304 22658 356 22668
rect 497 22658 549 22668
rect 688 22658 740 22668
rect 880 22658 932 22668
rect 1072 22658 1124 22668
rect 1264 22658 1316 22668
rect 1522 22659 1578 22669
rect 96 22606 304 22658
rect 356 22606 497 22658
rect 549 22606 688 22658
rect 740 22606 880 22658
rect 932 22606 1072 22658
rect 1124 22606 1264 22658
rect 1316 22606 1522 22658
rect 304 22596 356 22606
rect 497 22596 549 22606
rect 688 22596 740 22606
rect 880 22596 932 22606
rect 1072 22596 1124 22606
rect 1264 22596 1316 22606
rect 1522 22589 1578 22599
rect 1610 22026 1722 23169
rect 1608 22016 1722 22026
rect 1720 21892 1722 22016
rect 1608 21882 1722 21892
rect 304 21851 356 21861
rect 495 21851 547 21861
rect 687 21851 739 21861
rect 879 21851 931 21861
rect 1072 21851 1124 21860
rect 1264 21851 1316 21860
rect 1468 21854 1524 21864
rect 96 21799 304 21851
rect 356 21799 495 21851
rect 547 21799 687 21851
rect 739 21799 879 21851
rect 931 21850 1468 21851
rect 931 21799 1072 21850
rect 304 21789 356 21799
rect 495 21789 547 21799
rect 687 21789 739 21799
rect 879 21789 931 21799
rect 1124 21799 1264 21850
rect 1072 21788 1124 21798
rect 1316 21799 1468 21850
rect 1264 21788 1316 21798
rect 1524 21799 1526 21851
rect 1468 21788 1524 21798
rect 304 21371 356 21381
rect 497 21371 549 21381
rect 688 21371 740 21381
rect 880 21371 932 21381
rect 1072 21371 1124 21381
rect 1264 21371 1316 21381
rect 1522 21372 1578 21382
rect 96 21319 304 21371
rect 356 21319 497 21371
rect 549 21319 688 21371
rect 740 21319 880 21371
rect 932 21319 1072 21371
rect 1124 21319 1264 21371
rect 1316 21319 1522 21371
rect 304 21309 356 21319
rect 497 21309 549 21319
rect 688 21309 740 21319
rect 880 21309 932 21319
rect 1072 21309 1124 21319
rect 1264 21309 1316 21319
rect 1522 21302 1578 21312
rect 1610 20739 1722 21882
rect 1608 20729 1722 20739
rect 1720 20605 1722 20729
rect 1608 20595 1722 20605
rect 304 20564 356 20574
rect 495 20564 547 20574
rect 687 20564 739 20574
rect 879 20564 931 20574
rect 1072 20564 1124 20573
rect 1264 20564 1316 20573
rect 1468 20567 1524 20577
rect 96 20512 304 20564
rect 356 20512 495 20564
rect 547 20512 687 20564
rect 739 20512 879 20564
rect 931 20563 1468 20564
rect 931 20512 1072 20563
rect 304 20502 356 20512
rect 495 20502 547 20512
rect 687 20502 739 20512
rect 879 20502 931 20512
rect 1124 20512 1264 20563
rect 1072 20501 1124 20511
rect 1316 20512 1468 20563
rect 1264 20501 1316 20511
rect 1524 20512 1526 20564
rect 1468 20501 1524 20511
rect 304 20084 356 20094
rect 497 20084 549 20094
rect 688 20084 740 20094
rect 880 20084 932 20094
rect 1072 20084 1124 20094
rect 1264 20084 1316 20094
rect 1522 20085 1578 20095
rect 96 20032 304 20084
rect 356 20032 497 20084
rect 549 20032 688 20084
rect 740 20032 880 20084
rect 932 20032 1072 20084
rect 1124 20032 1264 20084
rect 1316 20032 1522 20084
rect 304 20022 356 20032
rect 497 20022 549 20032
rect 688 20022 740 20032
rect 880 20022 932 20032
rect 1072 20022 1124 20032
rect 1264 20022 1316 20032
rect 1522 20015 1578 20025
rect 1610 19452 1722 20595
rect 1608 19442 1722 19452
rect 1720 19318 1722 19442
rect 1608 19308 1722 19318
rect 304 19277 356 19287
rect 495 19277 547 19287
rect 687 19277 739 19287
rect 879 19277 931 19287
rect 1072 19277 1124 19286
rect 1264 19277 1316 19286
rect 1468 19280 1524 19290
rect 96 19225 304 19277
rect 356 19225 495 19277
rect 547 19225 687 19277
rect 739 19225 879 19277
rect 931 19276 1468 19277
rect 931 19225 1072 19276
rect 304 19215 356 19225
rect 495 19215 547 19225
rect 687 19215 739 19225
rect 879 19215 931 19225
rect 1124 19225 1264 19276
rect 1072 19214 1124 19224
rect 1316 19225 1468 19276
rect 1264 19214 1316 19224
rect 1524 19225 1526 19277
rect 1468 19214 1524 19224
rect 304 18797 356 18807
rect 497 18797 549 18807
rect 688 18797 740 18807
rect 880 18797 932 18807
rect 1072 18797 1124 18807
rect 1264 18797 1316 18807
rect 1522 18798 1578 18808
rect 96 18745 304 18797
rect 356 18745 497 18797
rect 549 18745 688 18797
rect 740 18745 880 18797
rect 932 18745 1072 18797
rect 1124 18745 1264 18797
rect 1316 18745 1522 18797
rect 304 18735 356 18745
rect 497 18735 549 18745
rect 688 18735 740 18745
rect 880 18735 932 18745
rect 1072 18735 1124 18745
rect 1264 18735 1316 18745
rect 1522 18728 1578 18738
rect 1610 18165 1722 19308
rect 1608 18155 1722 18165
rect 1720 18031 1722 18155
rect 1608 18021 1722 18031
rect 304 17990 356 18000
rect 495 17990 547 18000
rect 687 17990 739 18000
rect 879 17990 931 18000
rect 1072 17990 1124 17999
rect 1264 17990 1316 17999
rect 1468 17993 1524 18003
rect 96 17938 304 17990
rect 356 17938 495 17990
rect 547 17938 687 17990
rect 739 17938 879 17990
rect 931 17989 1468 17990
rect 931 17938 1072 17989
rect 304 17928 356 17938
rect 495 17928 547 17938
rect 687 17928 739 17938
rect 879 17928 931 17938
rect 1124 17938 1264 17989
rect 1072 17927 1124 17937
rect 1316 17938 1468 17989
rect 1264 17927 1316 17937
rect 1524 17938 1526 17990
rect 1468 17927 1524 17937
rect 304 17510 356 17520
rect 497 17510 549 17520
rect 688 17510 740 17520
rect 880 17510 932 17520
rect 1072 17510 1124 17520
rect 1264 17510 1316 17520
rect 1522 17511 1578 17521
rect 96 17458 304 17510
rect 356 17458 497 17510
rect 549 17458 688 17510
rect 740 17458 880 17510
rect 932 17458 1072 17510
rect 1124 17458 1264 17510
rect 1316 17458 1522 17510
rect 304 17448 356 17458
rect 497 17448 549 17458
rect 688 17448 740 17458
rect 880 17448 932 17458
rect 1072 17448 1124 17458
rect 1264 17448 1316 17458
rect 1522 17441 1578 17451
rect 1610 16878 1722 18021
rect 1608 16868 1722 16878
rect 1720 16744 1722 16868
rect 1608 16734 1722 16744
rect 304 16703 356 16713
rect 495 16703 547 16713
rect 687 16703 739 16713
rect 879 16703 931 16713
rect 1072 16703 1124 16712
rect 1264 16703 1316 16712
rect 1468 16706 1524 16716
rect 96 16651 304 16703
rect 356 16651 495 16703
rect 547 16651 687 16703
rect 739 16651 879 16703
rect 931 16702 1468 16703
rect 931 16651 1072 16702
rect 304 16641 356 16651
rect 495 16641 547 16651
rect 687 16641 739 16651
rect 879 16641 931 16651
rect 1124 16651 1264 16702
rect 1072 16640 1124 16650
rect 1316 16651 1468 16702
rect 1264 16640 1316 16650
rect 1524 16651 1526 16703
rect 1468 16640 1524 16650
rect 304 16223 356 16233
rect 497 16223 549 16233
rect 688 16223 740 16233
rect 880 16223 932 16233
rect 1072 16223 1124 16233
rect 1264 16223 1316 16233
rect 1522 16224 1578 16234
rect 96 16171 304 16223
rect 356 16171 497 16223
rect 549 16171 688 16223
rect 740 16171 880 16223
rect 932 16171 1072 16223
rect 1124 16171 1264 16223
rect 1316 16171 1522 16223
rect 304 16161 356 16171
rect 497 16161 549 16171
rect 688 16161 740 16171
rect 880 16161 932 16171
rect 1072 16161 1124 16171
rect 1264 16161 1316 16171
rect 1522 16154 1578 16164
rect 1610 15591 1722 16734
rect 1608 15581 1722 15591
rect 1720 15457 1722 15581
rect 1608 15447 1722 15457
rect 304 15416 356 15426
rect 495 15416 547 15426
rect 687 15416 739 15426
rect 879 15416 931 15426
rect 1072 15416 1124 15425
rect 1264 15416 1316 15425
rect 1468 15419 1524 15429
rect 96 15364 304 15416
rect 356 15364 495 15416
rect 547 15364 687 15416
rect 739 15364 879 15416
rect 931 15415 1468 15416
rect 931 15364 1072 15415
rect 304 15354 356 15364
rect 495 15354 547 15364
rect 687 15354 739 15364
rect 879 15354 931 15364
rect 1124 15364 1264 15415
rect 1072 15353 1124 15363
rect 1316 15364 1468 15415
rect 1264 15353 1316 15363
rect 1524 15364 1526 15416
rect 1468 15353 1524 15363
rect 304 14936 356 14946
rect 497 14936 549 14946
rect 688 14936 740 14946
rect 880 14936 932 14946
rect 1072 14936 1124 14946
rect 1264 14936 1316 14946
rect 1522 14937 1578 14947
rect 96 14884 304 14936
rect 356 14884 497 14936
rect 549 14884 688 14936
rect 740 14884 880 14936
rect 932 14884 1072 14936
rect 1124 14884 1264 14936
rect 1316 14884 1522 14936
rect 304 14874 356 14884
rect 497 14874 549 14884
rect 688 14874 740 14884
rect 880 14874 932 14884
rect 1072 14874 1124 14884
rect 1264 14874 1316 14884
rect 1522 14867 1578 14877
rect 1610 14304 1722 15447
rect 1608 14294 1722 14304
rect 1720 14170 1722 14294
rect 1608 14160 1722 14170
rect 304 14129 356 14139
rect 495 14129 547 14139
rect 687 14129 739 14139
rect 879 14129 931 14139
rect 1072 14129 1124 14138
rect 1264 14129 1316 14138
rect 1468 14132 1524 14142
rect 96 14077 304 14129
rect 356 14077 495 14129
rect 547 14077 687 14129
rect 739 14077 879 14129
rect 931 14128 1468 14129
rect 931 14077 1072 14128
rect 304 14067 356 14077
rect 495 14067 547 14077
rect 687 14067 739 14077
rect 879 14067 931 14077
rect 1124 14077 1264 14128
rect 1072 14066 1124 14076
rect 1316 14077 1468 14128
rect 1264 14066 1316 14076
rect 1524 14077 1526 14129
rect 1468 14066 1524 14076
rect 304 13649 356 13659
rect 497 13649 549 13659
rect 688 13649 740 13659
rect 880 13649 932 13659
rect 1072 13649 1124 13659
rect 1264 13649 1316 13659
rect 1522 13650 1578 13660
rect 96 13597 304 13649
rect 356 13597 497 13649
rect 549 13597 688 13649
rect 740 13597 880 13649
rect 932 13597 1072 13649
rect 1124 13597 1264 13649
rect 1316 13597 1522 13649
rect 304 13587 356 13597
rect 497 13587 549 13597
rect 688 13587 740 13597
rect 880 13587 932 13597
rect 1072 13587 1124 13597
rect 1264 13587 1316 13597
rect 1522 13580 1578 13590
rect 1610 13017 1722 14160
rect 1608 13007 1722 13017
rect 1720 12883 1722 13007
rect 1608 12873 1722 12883
rect 304 12842 356 12852
rect 495 12842 547 12852
rect 687 12842 739 12852
rect 879 12842 931 12852
rect 1072 12842 1124 12851
rect 1264 12842 1316 12851
rect 1468 12845 1524 12855
rect 96 12790 304 12842
rect 356 12790 495 12842
rect 547 12790 687 12842
rect 739 12790 879 12842
rect 931 12841 1468 12842
rect 931 12790 1072 12841
rect 304 12780 356 12790
rect 495 12780 547 12790
rect 687 12780 739 12790
rect 879 12780 931 12790
rect 1124 12790 1264 12841
rect 1072 12779 1124 12789
rect 1316 12790 1468 12841
rect 1264 12779 1316 12789
rect 1524 12790 1526 12842
rect 1468 12779 1524 12789
rect 304 12362 356 12372
rect 497 12362 549 12372
rect 688 12362 740 12372
rect 880 12362 932 12372
rect 1072 12362 1124 12372
rect 1264 12362 1316 12372
rect 1522 12363 1578 12373
rect 96 12310 304 12362
rect 356 12310 497 12362
rect 549 12310 688 12362
rect 740 12310 880 12362
rect 932 12310 1072 12362
rect 1124 12310 1264 12362
rect 1316 12310 1522 12362
rect 304 12300 356 12310
rect 497 12300 549 12310
rect 688 12300 740 12310
rect 880 12300 932 12310
rect 1072 12300 1124 12310
rect 1264 12300 1316 12310
rect 1522 12293 1578 12303
rect 1610 11730 1722 12873
rect 1608 11720 1722 11730
rect 1720 11596 1722 11720
rect 1608 11586 1722 11596
rect 304 11555 356 11565
rect 495 11555 547 11565
rect 687 11555 739 11565
rect 879 11555 931 11565
rect 1072 11555 1124 11564
rect 1264 11555 1316 11564
rect 1468 11558 1524 11568
rect 96 11503 304 11555
rect 356 11503 495 11555
rect 547 11503 687 11555
rect 739 11503 879 11555
rect 931 11554 1468 11555
rect 931 11503 1072 11554
rect 304 11493 356 11503
rect 495 11493 547 11503
rect 687 11493 739 11503
rect 879 11493 931 11503
rect 1124 11503 1264 11554
rect 1072 11492 1124 11502
rect 1316 11503 1468 11554
rect 1264 11492 1316 11502
rect 1524 11503 1526 11555
rect 1468 11492 1524 11502
rect 304 11075 356 11085
rect 497 11075 549 11085
rect 688 11075 740 11085
rect 880 11075 932 11085
rect 1072 11075 1124 11085
rect 1264 11075 1316 11085
rect 1522 11076 1578 11086
rect 96 11023 304 11075
rect 356 11023 497 11075
rect 549 11023 688 11075
rect 740 11023 880 11075
rect 932 11023 1072 11075
rect 1124 11023 1264 11075
rect 1316 11023 1522 11075
rect 304 11013 356 11023
rect 497 11013 549 11023
rect 688 11013 740 11023
rect 880 11013 932 11023
rect 1072 11013 1124 11023
rect 1264 11013 1316 11023
rect 1522 11006 1578 11016
rect 1610 10443 1722 11586
rect 1608 10433 1722 10443
rect 1720 10309 1722 10433
rect 1608 10299 1722 10309
rect 304 10268 356 10278
rect 495 10268 547 10278
rect 687 10268 739 10278
rect 879 10268 931 10278
rect 1072 10268 1124 10277
rect 1264 10268 1316 10277
rect 1468 10271 1524 10281
rect 96 10216 304 10268
rect 356 10216 495 10268
rect 547 10216 687 10268
rect 739 10216 879 10268
rect 931 10267 1468 10268
rect 931 10216 1072 10267
rect 304 10206 356 10216
rect 495 10206 547 10216
rect 687 10206 739 10216
rect 879 10206 931 10216
rect 1124 10216 1264 10267
rect 1072 10205 1124 10215
rect 1316 10216 1468 10267
rect 1264 10205 1316 10215
rect 1524 10216 1526 10268
rect 1468 10205 1524 10215
rect 304 9788 356 9798
rect 497 9788 549 9798
rect 688 9788 740 9798
rect 880 9788 932 9798
rect 1072 9788 1124 9798
rect 1264 9788 1316 9798
rect 1522 9789 1578 9799
rect 96 9736 304 9788
rect 356 9736 497 9788
rect 549 9736 688 9788
rect 740 9736 880 9788
rect 932 9736 1072 9788
rect 1124 9736 1264 9788
rect 1316 9736 1522 9788
rect 304 9726 356 9736
rect 497 9726 549 9736
rect 688 9726 740 9736
rect 880 9726 932 9736
rect 1072 9726 1124 9736
rect 1264 9726 1316 9736
rect 1522 9719 1578 9729
rect 1610 9156 1722 10299
rect 1608 9146 1722 9156
rect 1720 9022 1722 9146
rect 1608 9012 1722 9022
rect 304 8981 356 8991
rect 495 8981 547 8991
rect 687 8981 739 8991
rect 879 8981 931 8991
rect 1072 8981 1124 8990
rect 1264 8981 1316 8990
rect 1468 8984 1524 8994
rect 96 8929 304 8981
rect 356 8929 495 8981
rect 547 8929 687 8981
rect 739 8929 879 8981
rect 931 8980 1468 8981
rect 931 8929 1072 8980
rect 304 8919 356 8929
rect 495 8919 547 8929
rect 687 8919 739 8929
rect 879 8919 931 8929
rect 1124 8929 1264 8980
rect 1072 8918 1124 8928
rect 1316 8929 1468 8980
rect 1264 8918 1316 8928
rect 1524 8929 1526 8981
rect 1468 8918 1524 8928
rect 304 8501 356 8511
rect 497 8501 549 8511
rect 688 8501 740 8511
rect 880 8501 932 8511
rect 1072 8501 1124 8511
rect 1264 8501 1316 8511
rect 1522 8502 1578 8512
rect 96 8449 304 8501
rect 356 8449 497 8501
rect 549 8449 688 8501
rect 740 8449 880 8501
rect 932 8449 1072 8501
rect 1124 8449 1264 8501
rect 1316 8449 1522 8501
rect 304 8439 356 8449
rect 497 8439 549 8449
rect 688 8439 740 8449
rect 880 8439 932 8449
rect 1072 8439 1124 8449
rect 1264 8439 1316 8449
rect 1522 8432 1578 8442
rect 1610 7869 1722 9012
rect 1608 7859 1722 7869
rect 1720 7735 1722 7859
rect 1608 7725 1722 7735
rect 304 7694 356 7704
rect 495 7694 547 7704
rect 687 7694 739 7704
rect 879 7694 931 7704
rect 1072 7694 1124 7703
rect 1264 7694 1316 7703
rect 1468 7697 1524 7707
rect 96 7642 304 7694
rect 356 7642 495 7694
rect 547 7642 687 7694
rect 739 7642 879 7694
rect 931 7693 1468 7694
rect 931 7642 1072 7693
rect 304 7632 356 7642
rect 495 7632 547 7642
rect 687 7632 739 7642
rect 879 7632 931 7642
rect 1124 7642 1264 7693
rect 1072 7631 1124 7641
rect 1316 7642 1468 7693
rect 1264 7631 1316 7641
rect 1524 7642 1526 7694
rect 1468 7631 1524 7641
rect 304 7214 356 7224
rect 497 7214 549 7224
rect 688 7214 740 7224
rect 880 7214 932 7224
rect 1072 7214 1124 7224
rect 1264 7214 1316 7224
rect 1522 7215 1578 7225
rect 96 7162 304 7214
rect 356 7162 497 7214
rect 549 7162 688 7214
rect 740 7162 880 7214
rect 932 7162 1072 7214
rect 1124 7162 1264 7214
rect 1316 7162 1522 7214
rect 304 7152 356 7162
rect 497 7152 549 7162
rect 688 7152 740 7162
rect 880 7152 932 7162
rect 1072 7152 1124 7162
rect 1264 7152 1316 7162
rect 1522 7145 1578 7155
rect 1610 6582 1722 7725
rect 1608 6572 1722 6582
rect 1720 6448 1722 6572
rect 1608 6438 1722 6448
rect 304 6407 356 6417
rect 495 6407 547 6417
rect 687 6407 739 6417
rect 879 6407 931 6417
rect 1072 6407 1124 6416
rect 1264 6407 1316 6416
rect 1468 6410 1524 6420
rect 96 6355 304 6407
rect 356 6355 495 6407
rect 547 6355 687 6407
rect 739 6355 879 6407
rect 931 6406 1468 6407
rect 931 6355 1072 6406
rect 304 6345 356 6355
rect 495 6345 547 6355
rect 687 6345 739 6355
rect 879 6345 931 6355
rect 1124 6355 1264 6406
rect 1072 6344 1124 6354
rect 1316 6355 1468 6406
rect 1264 6344 1316 6354
rect 1524 6355 1526 6407
rect 1468 6344 1524 6354
rect 304 5927 356 5937
rect 497 5927 549 5937
rect 688 5927 740 5937
rect 880 5927 932 5937
rect 1072 5927 1124 5937
rect 1264 5927 1316 5937
rect 1522 5928 1578 5938
rect 96 5875 304 5927
rect 356 5875 497 5927
rect 549 5875 688 5927
rect 740 5875 880 5927
rect 932 5875 1072 5927
rect 1124 5875 1264 5927
rect 1316 5875 1522 5927
rect 304 5865 356 5875
rect 497 5865 549 5875
rect 688 5865 740 5875
rect 880 5865 932 5875
rect 1072 5865 1124 5875
rect 1264 5865 1316 5875
rect 1522 5858 1578 5868
rect 1610 5295 1722 6438
rect 1608 5285 1722 5295
rect 1720 5161 1722 5285
rect 1608 5151 1722 5161
rect 304 5120 356 5130
rect 495 5120 547 5130
rect 687 5120 739 5130
rect 879 5120 931 5130
rect 1072 5120 1124 5129
rect 1264 5120 1316 5129
rect 1468 5123 1524 5133
rect 96 5068 304 5120
rect 356 5068 495 5120
rect 547 5068 687 5120
rect 739 5068 879 5120
rect 931 5119 1468 5120
rect 931 5068 1072 5119
rect 304 5058 356 5068
rect 495 5058 547 5068
rect 687 5058 739 5068
rect 879 5058 931 5068
rect 1124 5068 1264 5119
rect 1072 5057 1124 5067
rect 1316 5068 1468 5119
rect 1264 5057 1316 5067
rect 1524 5068 1526 5120
rect 1468 5057 1524 5067
rect 304 4640 356 4650
rect 497 4640 549 4650
rect 688 4640 740 4650
rect 880 4640 932 4650
rect 1072 4640 1124 4650
rect 1264 4640 1316 4650
rect 1522 4641 1578 4651
rect 96 4588 304 4640
rect 356 4588 497 4640
rect 549 4588 688 4640
rect 740 4588 880 4640
rect 932 4588 1072 4640
rect 1124 4588 1264 4640
rect 1316 4588 1522 4640
rect 304 4578 356 4588
rect 497 4578 549 4588
rect 688 4578 740 4588
rect 880 4578 932 4588
rect 1072 4578 1124 4588
rect 1264 4578 1316 4588
rect 1522 4571 1578 4581
rect 1610 4008 1722 5151
rect 1608 3998 1722 4008
rect 1720 3874 1722 3998
rect 1608 3864 1722 3874
rect 304 3833 356 3843
rect 495 3833 547 3843
rect 687 3833 739 3843
rect 879 3833 931 3843
rect 1072 3833 1124 3842
rect 1264 3833 1316 3842
rect 1468 3836 1524 3846
rect 96 3781 304 3833
rect 356 3781 495 3833
rect 547 3781 687 3833
rect 739 3781 879 3833
rect 931 3832 1468 3833
rect 931 3781 1072 3832
rect 304 3771 356 3781
rect 495 3771 547 3781
rect 687 3771 739 3781
rect 879 3771 931 3781
rect 1124 3781 1264 3832
rect 1072 3770 1124 3780
rect 1316 3781 1468 3832
rect 1264 3770 1316 3780
rect 1524 3781 1526 3833
rect 1468 3770 1524 3780
rect 304 3353 356 3363
rect 497 3353 549 3363
rect 688 3353 740 3363
rect 880 3353 932 3363
rect 1072 3353 1124 3363
rect 1264 3353 1316 3363
rect 1522 3354 1578 3364
rect 96 3301 304 3353
rect 356 3301 497 3353
rect 549 3301 688 3353
rect 740 3301 880 3353
rect 932 3301 1072 3353
rect 1124 3301 1264 3353
rect 1316 3301 1522 3353
rect 304 3291 356 3301
rect 497 3291 549 3301
rect 688 3291 740 3301
rect 880 3291 932 3301
rect 1072 3291 1124 3301
rect 1264 3291 1316 3301
rect 1522 3284 1578 3294
rect 1610 2721 1722 3864
rect 1608 2711 1722 2721
rect 1720 2587 1722 2711
rect 1608 2577 1722 2587
rect 304 2546 356 2556
rect 495 2546 547 2556
rect 687 2546 739 2556
rect 879 2546 931 2556
rect 1072 2546 1124 2555
rect 1264 2546 1316 2555
rect 1468 2549 1524 2559
rect 96 2494 304 2546
rect 356 2494 495 2546
rect 547 2494 687 2546
rect 739 2494 879 2546
rect 931 2545 1468 2546
rect 931 2494 1072 2545
rect 304 2484 356 2494
rect 495 2484 547 2494
rect 687 2484 739 2494
rect 879 2484 931 2494
rect 1124 2494 1264 2545
rect 1072 2483 1124 2493
rect 1316 2494 1468 2545
rect 1264 2483 1316 2493
rect 1524 2494 1526 2546
rect 1468 2483 1524 2493
rect 304 2066 356 2076
rect 497 2066 549 2076
rect 688 2066 740 2076
rect 880 2066 932 2076
rect 1072 2066 1124 2076
rect 1264 2066 1316 2076
rect 1522 2067 1578 2077
rect 96 2014 304 2066
rect 356 2014 497 2066
rect 549 2014 688 2066
rect 740 2014 880 2066
rect 932 2014 1072 2066
rect 1124 2014 1264 2066
rect 1316 2014 1522 2066
rect 304 2004 356 2014
rect 497 2004 549 2014
rect 688 2004 740 2014
rect 880 2004 932 2014
rect 1072 2004 1124 2014
rect 1264 2004 1316 2014
rect 1522 1997 1578 2007
rect 1610 1434 1722 2577
rect 1608 1424 1722 1434
rect 1720 1300 1722 1424
rect 1608 1290 1722 1300
rect 304 1259 356 1269
rect 495 1259 547 1269
rect 687 1259 739 1269
rect 879 1259 931 1269
rect 1072 1259 1124 1268
rect 1264 1259 1316 1268
rect 1468 1262 1524 1272
rect 96 1207 304 1259
rect 356 1207 495 1259
rect 547 1207 687 1259
rect 739 1207 879 1259
rect 931 1258 1468 1259
rect 931 1207 1072 1258
rect 304 1197 356 1207
rect 495 1197 547 1207
rect 687 1197 739 1207
rect 879 1197 931 1207
rect 1124 1207 1264 1258
rect 1072 1196 1124 1206
rect 1316 1207 1468 1258
rect 1264 1196 1316 1206
rect 1524 1207 1526 1259
rect 1468 1196 1524 1206
rect 1610 1202 1722 1290
rect 1792 41964 1852 42267
rect 1792 40677 1852 41904
rect 1792 39390 1852 40617
rect 1792 38103 1852 39330
rect 1792 36816 1852 38043
rect 1792 35529 1852 36756
rect 1792 34242 1852 35469
rect 1792 32955 1852 34182
rect 1792 31668 1852 32895
rect 1792 30381 1852 31608
rect 1792 29094 1852 30321
rect 1792 27807 1852 29034
rect 1792 26520 1852 27747
rect 1792 25233 1852 26460
rect 1792 23946 1852 25173
rect 1792 22659 1852 23886
rect 1792 21372 1852 22599
rect 1792 20085 1852 21312
rect 1792 18798 1852 20025
rect 1792 17511 1852 18738
rect 1792 16224 1852 17451
rect 1792 14937 1852 16164
rect 1792 13650 1852 14877
rect 1792 12363 1852 13590
rect 1792 11076 1852 12303
rect 1792 9789 1852 11016
rect 1792 8502 1852 9729
rect 1792 7215 1852 8442
rect 1792 5928 1852 7155
rect 1792 4641 1852 5868
rect 1792 3354 1852 4581
rect 1792 2067 1852 3294
rect 1792 1202 1852 2007
rect 1930 41161 1986 42267
rect 2054 41665 2192 42212
rect 2457 41967 2509 41977
rect 2650 41967 2702 41977
rect 2841 41967 2893 41977
rect 3033 41967 3085 41977
rect 3225 41967 3277 41977
rect 3417 41967 3469 41977
rect 3978 41967 4030 41977
rect 4171 41967 4223 41977
rect 4362 41967 4414 41977
rect 4554 41967 4606 41977
rect 4746 41967 4798 41977
rect 4938 41967 4990 41977
rect 2233 41915 2457 41967
rect 2509 41915 2650 41967
rect 2702 41915 2841 41967
rect 2893 41915 3033 41967
rect 3085 41915 3225 41967
rect 3277 41915 3417 41967
rect 3469 41915 3978 41967
rect 4030 41915 4171 41967
rect 4223 41915 4362 41967
rect 4414 41915 4554 41967
rect 4606 41915 4746 41967
rect 4798 41915 4938 41967
rect 4990 41915 5846 41967
rect 2457 41905 2509 41915
rect 2650 41905 2702 41915
rect 2841 41905 2893 41915
rect 3033 41905 3085 41915
rect 3225 41905 3277 41915
rect 3417 41905 3469 41915
rect 2054 41557 2056 41665
rect 2190 41557 2192 41665
rect 2054 41554 2192 41557
rect 1930 39874 1986 41105
rect 1930 38587 1986 39818
rect 1930 37300 1986 38531
rect 1930 36013 1986 37244
rect 1930 34726 1986 35957
rect 1930 33439 1986 34670
rect 1930 32152 1986 33383
rect 1930 30865 1986 32096
rect 1930 29578 1986 30809
rect 1930 28291 1986 29522
rect 1930 27004 1986 28235
rect 1930 25717 1986 26948
rect 1930 24430 1986 25661
rect 1930 23143 1986 24374
rect 1930 21856 1986 23087
rect 1930 20569 1986 21800
rect 1930 19282 1986 20513
rect 1930 17995 1986 19226
rect 1930 16708 1986 17939
rect 1930 15421 1986 16652
rect 1930 14134 1986 15365
rect 1930 12847 1986 14078
rect 1930 11560 1986 12791
rect 1930 10273 1986 11504
rect 1930 8986 1986 10217
rect 1930 7699 1986 8930
rect 1930 6412 1986 7643
rect 1930 5125 1986 6356
rect 1930 3838 1986 5069
rect 1930 2551 1986 3782
rect 1930 1264 1986 2495
rect 2056 41427 2190 41554
rect 2056 40388 2186 41427
rect 3681 41390 3733 41915
rect 3978 41905 4030 41915
rect 4171 41905 4223 41915
rect 4362 41905 4414 41915
rect 4554 41905 4606 41915
rect 4746 41905 4798 41915
rect 4938 41905 4990 41915
rect 5336 41422 5390 41433
rect 5336 41415 5337 41422
rect 3681 41328 3733 41338
rect 5178 41370 5337 41415
rect 5389 41370 5390 41422
rect 5178 41363 5390 41370
rect 2457 41160 2509 41170
rect 2648 41160 2700 41170
rect 2840 41160 2892 41170
rect 3032 41160 3084 41170
rect 3225 41160 3277 41169
rect 3417 41160 3469 41169
rect 3978 41160 4030 41170
rect 4169 41160 4221 41170
rect 4361 41160 4413 41170
rect 4553 41160 4605 41170
rect 4746 41160 4798 41169
rect 4938 41160 4990 41169
rect 5178 41160 5230 41363
rect 5336 41359 5390 41363
rect 5448 41431 5502 41435
rect 5608 41431 5660 41915
rect 5448 41424 5660 41431
rect 5448 41372 5449 41424
rect 5501 41379 5660 41424
rect 5501 41372 5502 41379
rect 5448 41361 5502 41372
rect 2229 41108 2457 41160
rect 2509 41108 2648 41160
rect 2700 41108 2840 41160
rect 2892 41108 3032 41160
rect 3084 41159 3978 41160
rect 3084 41108 3225 41159
rect 2457 41098 2509 41108
rect 2648 41098 2700 41108
rect 2840 41098 2892 41108
rect 3032 41098 3084 41108
rect 3277 41108 3417 41159
rect 3225 41097 3277 41107
rect 3469 41108 3978 41159
rect 4030 41108 4169 41160
rect 4221 41108 4361 41160
rect 4413 41108 4553 41160
rect 4605 41159 5230 41160
rect 4605 41108 4746 41159
rect 3417 41097 3469 41107
rect 3978 41098 4030 41108
rect 4169 41098 4221 41108
rect 4361 41098 4413 41108
rect 4553 41098 4605 41108
rect 4798 41108 4938 41159
rect 4746 41097 4798 41107
rect 4990 41108 5230 41159
rect 4938 41097 4990 41107
rect 2457 40680 2509 40690
rect 2650 40680 2702 40690
rect 2841 40680 2893 40690
rect 3033 40680 3085 40690
rect 3225 40680 3277 40690
rect 3417 40680 3469 40690
rect 3978 40680 4030 40690
rect 4171 40680 4223 40690
rect 4362 40680 4414 40690
rect 4554 40680 4606 40690
rect 4746 40680 4798 40690
rect 4938 40680 4990 40690
rect 2233 40628 2457 40680
rect 2509 40628 2650 40680
rect 2702 40628 2841 40680
rect 2893 40628 3033 40680
rect 3085 40628 3225 40680
rect 3277 40628 3417 40680
rect 3469 40628 3978 40680
rect 4030 40628 4171 40680
rect 4223 40628 4362 40680
rect 4414 40628 4554 40680
rect 4606 40628 4746 40680
rect 4798 40628 4938 40680
rect 4990 40628 5846 40680
rect 2457 40618 2509 40628
rect 2650 40618 2702 40628
rect 2841 40618 2893 40628
rect 3033 40618 3085 40628
rect 3225 40618 3277 40628
rect 3417 40618 3469 40628
rect 2056 40378 2190 40388
rect 2056 40140 2190 40270
rect 2056 39101 2186 40140
rect 3681 40103 3733 40628
rect 3978 40618 4030 40628
rect 4171 40618 4223 40628
rect 4362 40618 4414 40628
rect 4554 40618 4606 40628
rect 4746 40618 4798 40628
rect 4938 40618 4990 40628
rect 5336 40135 5390 40146
rect 5336 40128 5337 40135
rect 3681 40041 3733 40051
rect 5178 40083 5337 40128
rect 5389 40083 5390 40135
rect 5178 40076 5390 40083
rect 2457 39873 2509 39883
rect 2648 39873 2700 39883
rect 2840 39873 2892 39883
rect 3032 39873 3084 39883
rect 3225 39873 3277 39882
rect 3417 39873 3469 39882
rect 3978 39873 4030 39883
rect 4169 39873 4221 39883
rect 4361 39873 4413 39883
rect 4553 39873 4605 39883
rect 4746 39873 4798 39882
rect 4938 39873 4990 39882
rect 5178 39873 5230 40076
rect 5336 40072 5390 40076
rect 5448 40144 5502 40148
rect 5608 40144 5660 40628
rect 5448 40137 5660 40144
rect 5448 40085 5449 40137
rect 5501 40092 5660 40137
rect 5501 40085 5502 40092
rect 5448 40074 5502 40085
rect 2229 39821 2457 39873
rect 2509 39821 2648 39873
rect 2700 39821 2840 39873
rect 2892 39821 3032 39873
rect 3084 39872 3978 39873
rect 3084 39821 3225 39872
rect 2457 39811 2509 39821
rect 2648 39811 2700 39821
rect 2840 39811 2892 39821
rect 3032 39811 3084 39821
rect 3277 39821 3417 39872
rect 3225 39810 3277 39820
rect 3469 39821 3978 39872
rect 4030 39821 4169 39873
rect 4221 39821 4361 39873
rect 4413 39821 4553 39873
rect 4605 39872 5230 39873
rect 4605 39821 4746 39872
rect 3417 39810 3469 39820
rect 3978 39811 4030 39821
rect 4169 39811 4221 39821
rect 4361 39811 4413 39821
rect 4553 39811 4605 39821
rect 4798 39821 4938 39872
rect 4746 39810 4798 39820
rect 4990 39821 5230 39872
rect 4938 39810 4990 39820
rect 2457 39393 2509 39403
rect 2650 39393 2702 39403
rect 2841 39393 2893 39403
rect 3033 39393 3085 39403
rect 3225 39393 3277 39403
rect 3417 39393 3469 39403
rect 3978 39393 4030 39403
rect 4171 39393 4223 39403
rect 4362 39393 4414 39403
rect 4554 39393 4606 39403
rect 4746 39393 4798 39403
rect 4938 39393 4990 39403
rect 2233 39341 2457 39393
rect 2509 39341 2650 39393
rect 2702 39341 2841 39393
rect 2893 39341 3033 39393
rect 3085 39341 3225 39393
rect 3277 39341 3417 39393
rect 3469 39341 3978 39393
rect 4030 39341 4171 39393
rect 4223 39341 4362 39393
rect 4414 39341 4554 39393
rect 4606 39341 4746 39393
rect 4798 39341 4938 39393
rect 4990 39341 5846 39393
rect 2457 39331 2509 39341
rect 2650 39331 2702 39341
rect 2841 39331 2893 39341
rect 3033 39331 3085 39341
rect 3225 39331 3277 39341
rect 3417 39331 3469 39341
rect 2056 39091 2190 39101
rect 2056 38853 2190 38983
rect 2056 37814 2186 38853
rect 3681 38816 3733 39341
rect 3978 39331 4030 39341
rect 4171 39331 4223 39341
rect 4362 39331 4414 39341
rect 4554 39331 4606 39341
rect 4746 39331 4798 39341
rect 4938 39331 4990 39341
rect 5336 38848 5390 38859
rect 5336 38841 5337 38848
rect 3681 38754 3733 38764
rect 5178 38796 5337 38841
rect 5389 38796 5390 38848
rect 5178 38789 5390 38796
rect 2457 38586 2509 38596
rect 2648 38586 2700 38596
rect 2840 38586 2892 38596
rect 3032 38586 3084 38596
rect 3225 38586 3277 38595
rect 3417 38586 3469 38595
rect 3978 38586 4030 38596
rect 4169 38586 4221 38596
rect 4361 38586 4413 38596
rect 4553 38586 4605 38596
rect 4746 38586 4798 38595
rect 4938 38586 4990 38595
rect 5178 38586 5230 38789
rect 5336 38785 5390 38789
rect 5448 38857 5502 38861
rect 5608 38857 5660 39341
rect 5448 38850 5660 38857
rect 5448 38798 5449 38850
rect 5501 38805 5660 38850
rect 5501 38798 5502 38805
rect 5448 38787 5502 38798
rect 2229 38534 2457 38586
rect 2509 38534 2648 38586
rect 2700 38534 2840 38586
rect 2892 38534 3032 38586
rect 3084 38585 3978 38586
rect 3084 38534 3225 38585
rect 2457 38524 2509 38534
rect 2648 38524 2700 38534
rect 2840 38524 2892 38534
rect 3032 38524 3084 38534
rect 3277 38534 3417 38585
rect 3225 38523 3277 38533
rect 3469 38534 3978 38585
rect 4030 38534 4169 38586
rect 4221 38534 4361 38586
rect 4413 38534 4553 38586
rect 4605 38585 5230 38586
rect 4605 38534 4746 38585
rect 3417 38523 3469 38533
rect 3978 38524 4030 38534
rect 4169 38524 4221 38534
rect 4361 38524 4413 38534
rect 4553 38524 4605 38534
rect 4798 38534 4938 38585
rect 4746 38523 4798 38533
rect 4990 38534 5230 38585
rect 4938 38523 4990 38533
rect 2457 38106 2509 38116
rect 2650 38106 2702 38116
rect 2841 38106 2893 38116
rect 3033 38106 3085 38116
rect 3225 38106 3277 38116
rect 3417 38106 3469 38116
rect 3978 38106 4030 38116
rect 4171 38106 4223 38116
rect 4362 38106 4414 38116
rect 4554 38106 4606 38116
rect 4746 38106 4798 38116
rect 4938 38106 4990 38116
rect 2233 38054 2457 38106
rect 2509 38054 2650 38106
rect 2702 38054 2841 38106
rect 2893 38054 3033 38106
rect 3085 38054 3225 38106
rect 3277 38054 3417 38106
rect 3469 38054 3978 38106
rect 4030 38054 4171 38106
rect 4223 38054 4362 38106
rect 4414 38054 4554 38106
rect 4606 38054 4746 38106
rect 4798 38054 4938 38106
rect 4990 38054 5846 38106
rect 2457 38044 2509 38054
rect 2650 38044 2702 38054
rect 2841 38044 2893 38054
rect 3033 38044 3085 38054
rect 3225 38044 3277 38054
rect 3417 38044 3469 38054
rect 2056 37804 2190 37814
rect 2056 37566 2190 37696
rect 2056 36527 2186 37566
rect 3681 37529 3733 38054
rect 3978 38044 4030 38054
rect 4171 38044 4223 38054
rect 4362 38044 4414 38054
rect 4554 38044 4606 38054
rect 4746 38044 4798 38054
rect 4938 38044 4990 38054
rect 5336 37561 5390 37572
rect 5336 37554 5337 37561
rect 3681 37467 3733 37477
rect 5178 37509 5337 37554
rect 5389 37509 5390 37561
rect 5178 37502 5390 37509
rect 2457 37299 2509 37309
rect 2648 37299 2700 37309
rect 2840 37299 2892 37309
rect 3032 37299 3084 37309
rect 3225 37299 3277 37308
rect 3417 37299 3469 37308
rect 3978 37299 4030 37309
rect 4169 37299 4221 37309
rect 4361 37299 4413 37309
rect 4553 37299 4605 37309
rect 4746 37299 4798 37308
rect 4938 37299 4990 37308
rect 5178 37299 5230 37502
rect 5336 37498 5390 37502
rect 5448 37570 5502 37574
rect 5608 37570 5660 38054
rect 5448 37563 5660 37570
rect 5448 37511 5449 37563
rect 5501 37518 5660 37563
rect 5501 37511 5502 37518
rect 5448 37500 5502 37511
rect 2229 37247 2457 37299
rect 2509 37247 2648 37299
rect 2700 37247 2840 37299
rect 2892 37247 3032 37299
rect 3084 37298 3978 37299
rect 3084 37247 3225 37298
rect 2457 37237 2509 37247
rect 2648 37237 2700 37247
rect 2840 37237 2892 37247
rect 3032 37237 3084 37247
rect 3277 37247 3417 37298
rect 3225 37236 3277 37246
rect 3469 37247 3978 37298
rect 4030 37247 4169 37299
rect 4221 37247 4361 37299
rect 4413 37247 4553 37299
rect 4605 37298 5230 37299
rect 4605 37247 4746 37298
rect 3417 37236 3469 37246
rect 3978 37237 4030 37247
rect 4169 37237 4221 37247
rect 4361 37237 4413 37247
rect 4553 37237 4605 37247
rect 4798 37247 4938 37298
rect 4746 37236 4798 37246
rect 4990 37247 5230 37298
rect 4938 37236 4990 37246
rect 2457 36819 2509 36829
rect 2650 36819 2702 36829
rect 2841 36819 2893 36829
rect 3033 36819 3085 36829
rect 3225 36819 3277 36829
rect 3417 36819 3469 36829
rect 3978 36819 4030 36829
rect 4171 36819 4223 36829
rect 4362 36819 4414 36829
rect 4554 36819 4606 36829
rect 4746 36819 4798 36829
rect 4938 36819 4990 36829
rect 2233 36767 2457 36819
rect 2509 36767 2650 36819
rect 2702 36767 2841 36819
rect 2893 36767 3033 36819
rect 3085 36767 3225 36819
rect 3277 36767 3417 36819
rect 3469 36767 3978 36819
rect 4030 36767 4171 36819
rect 4223 36767 4362 36819
rect 4414 36767 4554 36819
rect 4606 36767 4746 36819
rect 4798 36767 4938 36819
rect 4990 36767 5846 36819
rect 2457 36757 2509 36767
rect 2650 36757 2702 36767
rect 2841 36757 2893 36767
rect 3033 36757 3085 36767
rect 3225 36757 3277 36767
rect 3417 36757 3469 36767
rect 2056 36517 2190 36527
rect 2056 36279 2190 36409
rect 2056 35240 2186 36279
rect 3681 36242 3733 36767
rect 3978 36757 4030 36767
rect 4171 36757 4223 36767
rect 4362 36757 4414 36767
rect 4554 36757 4606 36767
rect 4746 36757 4798 36767
rect 4938 36757 4990 36767
rect 5336 36274 5390 36285
rect 5336 36267 5337 36274
rect 3681 36180 3733 36190
rect 5178 36222 5337 36267
rect 5389 36222 5390 36274
rect 5178 36215 5390 36222
rect 2457 36012 2509 36022
rect 2648 36012 2700 36022
rect 2840 36012 2892 36022
rect 3032 36012 3084 36022
rect 3225 36012 3277 36021
rect 3417 36012 3469 36021
rect 3978 36012 4030 36022
rect 4169 36012 4221 36022
rect 4361 36012 4413 36022
rect 4553 36012 4605 36022
rect 4746 36012 4798 36021
rect 4938 36012 4990 36021
rect 5178 36012 5230 36215
rect 5336 36211 5390 36215
rect 5448 36283 5502 36287
rect 5608 36283 5660 36767
rect 5448 36276 5660 36283
rect 5448 36224 5449 36276
rect 5501 36231 5660 36276
rect 5501 36224 5502 36231
rect 5448 36213 5502 36224
rect 2229 35960 2457 36012
rect 2509 35960 2648 36012
rect 2700 35960 2840 36012
rect 2892 35960 3032 36012
rect 3084 36011 3978 36012
rect 3084 35960 3225 36011
rect 2457 35950 2509 35960
rect 2648 35950 2700 35960
rect 2840 35950 2892 35960
rect 3032 35950 3084 35960
rect 3277 35960 3417 36011
rect 3225 35949 3277 35959
rect 3469 35960 3978 36011
rect 4030 35960 4169 36012
rect 4221 35960 4361 36012
rect 4413 35960 4553 36012
rect 4605 36011 5230 36012
rect 4605 35960 4746 36011
rect 3417 35949 3469 35959
rect 3978 35950 4030 35960
rect 4169 35950 4221 35960
rect 4361 35950 4413 35960
rect 4553 35950 4605 35960
rect 4798 35960 4938 36011
rect 4746 35949 4798 35959
rect 4990 35960 5230 36011
rect 4938 35949 4990 35959
rect 2457 35532 2509 35542
rect 2650 35532 2702 35542
rect 2841 35532 2893 35542
rect 3033 35532 3085 35542
rect 3225 35532 3277 35542
rect 3417 35532 3469 35542
rect 3978 35532 4030 35542
rect 4171 35532 4223 35542
rect 4362 35532 4414 35542
rect 4554 35532 4606 35542
rect 4746 35532 4798 35542
rect 4938 35532 4990 35542
rect 2233 35480 2457 35532
rect 2509 35480 2650 35532
rect 2702 35480 2841 35532
rect 2893 35480 3033 35532
rect 3085 35480 3225 35532
rect 3277 35480 3417 35532
rect 3469 35480 3978 35532
rect 4030 35480 4171 35532
rect 4223 35480 4362 35532
rect 4414 35480 4554 35532
rect 4606 35480 4746 35532
rect 4798 35480 4938 35532
rect 4990 35480 5846 35532
rect 2457 35470 2509 35480
rect 2650 35470 2702 35480
rect 2841 35470 2893 35480
rect 3033 35470 3085 35480
rect 3225 35470 3277 35480
rect 3417 35470 3469 35480
rect 2056 35230 2190 35240
rect 2056 34992 2190 35122
rect 2056 33953 2186 34992
rect 3681 34955 3733 35480
rect 3978 35470 4030 35480
rect 4171 35470 4223 35480
rect 4362 35470 4414 35480
rect 4554 35470 4606 35480
rect 4746 35470 4798 35480
rect 4938 35470 4990 35480
rect 5336 34987 5390 34998
rect 5336 34980 5337 34987
rect 3681 34893 3733 34903
rect 5178 34935 5337 34980
rect 5389 34935 5390 34987
rect 5178 34928 5390 34935
rect 2457 34725 2509 34735
rect 2648 34725 2700 34735
rect 2840 34725 2892 34735
rect 3032 34725 3084 34735
rect 3225 34725 3277 34734
rect 3417 34725 3469 34734
rect 3978 34725 4030 34735
rect 4169 34725 4221 34735
rect 4361 34725 4413 34735
rect 4553 34725 4605 34735
rect 4746 34725 4798 34734
rect 4938 34725 4990 34734
rect 5178 34725 5230 34928
rect 5336 34924 5390 34928
rect 5448 34996 5502 35000
rect 5608 34996 5660 35480
rect 5448 34989 5660 34996
rect 5448 34937 5449 34989
rect 5501 34944 5660 34989
rect 5501 34937 5502 34944
rect 5448 34926 5502 34937
rect 2229 34673 2457 34725
rect 2509 34673 2648 34725
rect 2700 34673 2840 34725
rect 2892 34673 3032 34725
rect 3084 34724 3978 34725
rect 3084 34673 3225 34724
rect 2457 34663 2509 34673
rect 2648 34663 2700 34673
rect 2840 34663 2892 34673
rect 3032 34663 3084 34673
rect 3277 34673 3417 34724
rect 3225 34662 3277 34672
rect 3469 34673 3978 34724
rect 4030 34673 4169 34725
rect 4221 34673 4361 34725
rect 4413 34673 4553 34725
rect 4605 34724 5230 34725
rect 4605 34673 4746 34724
rect 3417 34662 3469 34672
rect 3978 34663 4030 34673
rect 4169 34663 4221 34673
rect 4361 34663 4413 34673
rect 4553 34663 4605 34673
rect 4798 34673 4938 34724
rect 4746 34662 4798 34672
rect 4990 34673 5230 34724
rect 4938 34662 4990 34672
rect 2457 34245 2509 34255
rect 2650 34245 2702 34255
rect 2841 34245 2893 34255
rect 3033 34245 3085 34255
rect 3225 34245 3277 34255
rect 3417 34245 3469 34255
rect 3978 34245 4030 34255
rect 4171 34245 4223 34255
rect 4362 34245 4414 34255
rect 4554 34245 4606 34255
rect 4746 34245 4798 34255
rect 4938 34245 4990 34255
rect 2233 34193 2457 34245
rect 2509 34193 2650 34245
rect 2702 34193 2841 34245
rect 2893 34193 3033 34245
rect 3085 34193 3225 34245
rect 3277 34193 3417 34245
rect 3469 34193 3978 34245
rect 4030 34193 4171 34245
rect 4223 34193 4362 34245
rect 4414 34193 4554 34245
rect 4606 34193 4746 34245
rect 4798 34193 4938 34245
rect 4990 34193 5846 34245
rect 2457 34183 2509 34193
rect 2650 34183 2702 34193
rect 2841 34183 2893 34193
rect 3033 34183 3085 34193
rect 3225 34183 3277 34193
rect 3417 34183 3469 34193
rect 2056 33943 2190 33953
rect 2056 33705 2190 33835
rect 2056 32666 2186 33705
rect 3681 33668 3733 34193
rect 3978 34183 4030 34193
rect 4171 34183 4223 34193
rect 4362 34183 4414 34193
rect 4554 34183 4606 34193
rect 4746 34183 4798 34193
rect 4938 34183 4990 34193
rect 5336 33700 5390 33711
rect 5336 33693 5337 33700
rect 3681 33606 3733 33616
rect 5178 33648 5337 33693
rect 5389 33648 5390 33700
rect 5178 33641 5390 33648
rect 2457 33438 2509 33448
rect 2648 33438 2700 33448
rect 2840 33438 2892 33448
rect 3032 33438 3084 33448
rect 3225 33438 3277 33447
rect 3417 33438 3469 33447
rect 3978 33438 4030 33448
rect 4169 33438 4221 33448
rect 4361 33438 4413 33448
rect 4553 33438 4605 33448
rect 4746 33438 4798 33447
rect 4938 33438 4990 33447
rect 5178 33438 5230 33641
rect 5336 33637 5390 33641
rect 5448 33709 5502 33713
rect 5608 33709 5660 34193
rect 5448 33702 5660 33709
rect 5448 33650 5449 33702
rect 5501 33657 5660 33702
rect 5501 33650 5502 33657
rect 5448 33639 5502 33650
rect 2229 33386 2457 33438
rect 2509 33386 2648 33438
rect 2700 33386 2840 33438
rect 2892 33386 3032 33438
rect 3084 33437 3978 33438
rect 3084 33386 3225 33437
rect 2457 33376 2509 33386
rect 2648 33376 2700 33386
rect 2840 33376 2892 33386
rect 3032 33376 3084 33386
rect 3277 33386 3417 33437
rect 3225 33375 3277 33385
rect 3469 33386 3978 33437
rect 4030 33386 4169 33438
rect 4221 33386 4361 33438
rect 4413 33386 4553 33438
rect 4605 33437 5230 33438
rect 4605 33386 4746 33437
rect 3417 33375 3469 33385
rect 3978 33376 4030 33386
rect 4169 33376 4221 33386
rect 4361 33376 4413 33386
rect 4553 33376 4605 33386
rect 4798 33386 4938 33437
rect 4746 33375 4798 33385
rect 4990 33386 5230 33437
rect 4938 33375 4990 33385
rect 2457 32958 2509 32968
rect 2650 32958 2702 32968
rect 2841 32958 2893 32968
rect 3033 32958 3085 32968
rect 3225 32958 3277 32968
rect 3417 32958 3469 32968
rect 3978 32958 4030 32968
rect 4171 32958 4223 32968
rect 4362 32958 4414 32968
rect 4554 32958 4606 32968
rect 4746 32958 4798 32968
rect 4938 32958 4990 32968
rect 2233 32906 2457 32958
rect 2509 32906 2650 32958
rect 2702 32906 2841 32958
rect 2893 32906 3033 32958
rect 3085 32906 3225 32958
rect 3277 32906 3417 32958
rect 3469 32906 3978 32958
rect 4030 32906 4171 32958
rect 4223 32906 4362 32958
rect 4414 32906 4554 32958
rect 4606 32906 4746 32958
rect 4798 32906 4938 32958
rect 4990 32906 5846 32958
rect 2457 32896 2509 32906
rect 2650 32896 2702 32906
rect 2841 32896 2893 32906
rect 3033 32896 3085 32906
rect 3225 32896 3277 32906
rect 3417 32896 3469 32906
rect 2056 32656 2190 32666
rect 2056 32418 2190 32548
rect 2056 31379 2186 32418
rect 3681 32381 3733 32906
rect 3978 32896 4030 32906
rect 4171 32896 4223 32906
rect 4362 32896 4414 32906
rect 4554 32896 4606 32906
rect 4746 32896 4798 32906
rect 4938 32896 4990 32906
rect 5336 32413 5390 32424
rect 5336 32406 5337 32413
rect 3681 32319 3733 32329
rect 5178 32361 5337 32406
rect 5389 32361 5390 32413
rect 5178 32354 5390 32361
rect 2457 32151 2509 32161
rect 2648 32151 2700 32161
rect 2840 32151 2892 32161
rect 3032 32151 3084 32161
rect 3225 32151 3277 32160
rect 3417 32151 3469 32160
rect 3978 32151 4030 32161
rect 4169 32151 4221 32161
rect 4361 32151 4413 32161
rect 4553 32151 4605 32161
rect 4746 32151 4798 32160
rect 4938 32151 4990 32160
rect 5178 32151 5230 32354
rect 5336 32350 5390 32354
rect 5448 32422 5502 32426
rect 5608 32422 5660 32906
rect 5448 32415 5660 32422
rect 5448 32363 5449 32415
rect 5501 32370 5660 32415
rect 5501 32363 5502 32370
rect 5448 32352 5502 32363
rect 2229 32099 2457 32151
rect 2509 32099 2648 32151
rect 2700 32099 2840 32151
rect 2892 32099 3032 32151
rect 3084 32150 3978 32151
rect 3084 32099 3225 32150
rect 2457 32089 2509 32099
rect 2648 32089 2700 32099
rect 2840 32089 2892 32099
rect 3032 32089 3084 32099
rect 3277 32099 3417 32150
rect 3225 32088 3277 32098
rect 3469 32099 3978 32150
rect 4030 32099 4169 32151
rect 4221 32099 4361 32151
rect 4413 32099 4553 32151
rect 4605 32150 5230 32151
rect 4605 32099 4746 32150
rect 3417 32088 3469 32098
rect 3978 32089 4030 32099
rect 4169 32089 4221 32099
rect 4361 32089 4413 32099
rect 4553 32089 4605 32099
rect 4798 32099 4938 32150
rect 4746 32088 4798 32098
rect 4990 32099 5230 32150
rect 4938 32088 4990 32098
rect 2457 31671 2509 31681
rect 2650 31671 2702 31681
rect 2841 31671 2893 31681
rect 3033 31671 3085 31681
rect 3225 31671 3277 31681
rect 3417 31671 3469 31681
rect 3978 31671 4030 31681
rect 4171 31671 4223 31681
rect 4362 31671 4414 31681
rect 4554 31671 4606 31681
rect 4746 31671 4798 31681
rect 4938 31671 4990 31681
rect 2233 31619 2457 31671
rect 2509 31619 2650 31671
rect 2702 31619 2841 31671
rect 2893 31619 3033 31671
rect 3085 31619 3225 31671
rect 3277 31619 3417 31671
rect 3469 31619 3978 31671
rect 4030 31619 4171 31671
rect 4223 31619 4362 31671
rect 4414 31619 4554 31671
rect 4606 31619 4746 31671
rect 4798 31619 4938 31671
rect 4990 31619 5846 31671
rect 2457 31609 2509 31619
rect 2650 31609 2702 31619
rect 2841 31609 2893 31619
rect 3033 31609 3085 31619
rect 3225 31609 3277 31619
rect 3417 31609 3469 31619
rect 2056 31369 2190 31379
rect 2056 31131 2190 31261
rect 2056 30092 2186 31131
rect 3681 31094 3733 31619
rect 3978 31609 4030 31619
rect 4171 31609 4223 31619
rect 4362 31609 4414 31619
rect 4554 31609 4606 31619
rect 4746 31609 4798 31619
rect 4938 31609 4990 31619
rect 5336 31126 5390 31137
rect 5336 31119 5337 31126
rect 3681 31032 3733 31042
rect 5178 31074 5337 31119
rect 5389 31074 5390 31126
rect 5178 31067 5390 31074
rect 2457 30864 2509 30874
rect 2648 30864 2700 30874
rect 2840 30864 2892 30874
rect 3032 30864 3084 30874
rect 3225 30864 3277 30873
rect 3417 30864 3469 30873
rect 3978 30864 4030 30874
rect 4169 30864 4221 30874
rect 4361 30864 4413 30874
rect 4553 30864 4605 30874
rect 4746 30864 4798 30873
rect 4938 30864 4990 30873
rect 5178 30864 5230 31067
rect 5336 31063 5390 31067
rect 5448 31135 5502 31139
rect 5608 31135 5660 31619
rect 5448 31128 5660 31135
rect 5448 31076 5449 31128
rect 5501 31083 5660 31128
rect 5501 31076 5502 31083
rect 5448 31065 5502 31076
rect 2229 30812 2457 30864
rect 2509 30812 2648 30864
rect 2700 30812 2840 30864
rect 2892 30812 3032 30864
rect 3084 30863 3978 30864
rect 3084 30812 3225 30863
rect 2457 30802 2509 30812
rect 2648 30802 2700 30812
rect 2840 30802 2892 30812
rect 3032 30802 3084 30812
rect 3277 30812 3417 30863
rect 3225 30801 3277 30811
rect 3469 30812 3978 30863
rect 4030 30812 4169 30864
rect 4221 30812 4361 30864
rect 4413 30812 4553 30864
rect 4605 30863 5230 30864
rect 4605 30812 4746 30863
rect 3417 30801 3469 30811
rect 3978 30802 4030 30812
rect 4169 30802 4221 30812
rect 4361 30802 4413 30812
rect 4553 30802 4605 30812
rect 4798 30812 4938 30863
rect 4746 30801 4798 30811
rect 4990 30812 5230 30863
rect 4938 30801 4990 30811
rect 2457 30384 2509 30394
rect 2650 30384 2702 30394
rect 2841 30384 2893 30394
rect 3033 30384 3085 30394
rect 3225 30384 3277 30394
rect 3417 30384 3469 30394
rect 3978 30384 4030 30394
rect 4171 30384 4223 30394
rect 4362 30384 4414 30394
rect 4554 30384 4606 30394
rect 4746 30384 4798 30394
rect 4938 30384 4990 30394
rect 2233 30332 2457 30384
rect 2509 30332 2650 30384
rect 2702 30332 2841 30384
rect 2893 30332 3033 30384
rect 3085 30332 3225 30384
rect 3277 30332 3417 30384
rect 3469 30332 3978 30384
rect 4030 30332 4171 30384
rect 4223 30332 4362 30384
rect 4414 30332 4554 30384
rect 4606 30332 4746 30384
rect 4798 30332 4938 30384
rect 4990 30332 5846 30384
rect 2457 30322 2509 30332
rect 2650 30322 2702 30332
rect 2841 30322 2893 30332
rect 3033 30322 3085 30332
rect 3225 30322 3277 30332
rect 3417 30322 3469 30332
rect 2056 30082 2190 30092
rect 2056 29844 2190 29974
rect 2056 28805 2186 29844
rect 3681 29807 3733 30332
rect 3978 30322 4030 30332
rect 4171 30322 4223 30332
rect 4362 30322 4414 30332
rect 4554 30322 4606 30332
rect 4746 30322 4798 30332
rect 4938 30322 4990 30332
rect 5336 29839 5390 29850
rect 5336 29832 5337 29839
rect 3681 29745 3733 29755
rect 5178 29787 5337 29832
rect 5389 29787 5390 29839
rect 5178 29780 5390 29787
rect 2457 29577 2509 29587
rect 2648 29577 2700 29587
rect 2840 29577 2892 29587
rect 3032 29577 3084 29587
rect 3225 29577 3277 29586
rect 3417 29577 3469 29586
rect 3978 29577 4030 29587
rect 4169 29577 4221 29587
rect 4361 29577 4413 29587
rect 4553 29577 4605 29587
rect 4746 29577 4798 29586
rect 4938 29577 4990 29586
rect 5178 29577 5230 29780
rect 5336 29776 5390 29780
rect 5448 29848 5502 29852
rect 5608 29848 5660 30332
rect 5448 29841 5660 29848
rect 5448 29789 5449 29841
rect 5501 29796 5660 29841
rect 5501 29789 5502 29796
rect 5448 29778 5502 29789
rect 2229 29525 2457 29577
rect 2509 29525 2648 29577
rect 2700 29525 2840 29577
rect 2892 29525 3032 29577
rect 3084 29576 3978 29577
rect 3084 29525 3225 29576
rect 2457 29515 2509 29525
rect 2648 29515 2700 29525
rect 2840 29515 2892 29525
rect 3032 29515 3084 29525
rect 3277 29525 3417 29576
rect 3225 29514 3277 29524
rect 3469 29525 3978 29576
rect 4030 29525 4169 29577
rect 4221 29525 4361 29577
rect 4413 29525 4553 29577
rect 4605 29576 5230 29577
rect 4605 29525 4746 29576
rect 3417 29514 3469 29524
rect 3978 29515 4030 29525
rect 4169 29515 4221 29525
rect 4361 29515 4413 29525
rect 4553 29515 4605 29525
rect 4798 29525 4938 29576
rect 4746 29514 4798 29524
rect 4990 29525 5230 29576
rect 4938 29514 4990 29524
rect 2457 29097 2509 29107
rect 2650 29097 2702 29107
rect 2841 29097 2893 29107
rect 3033 29097 3085 29107
rect 3225 29097 3277 29107
rect 3417 29097 3469 29107
rect 3978 29097 4030 29107
rect 4171 29097 4223 29107
rect 4362 29097 4414 29107
rect 4554 29097 4606 29107
rect 4746 29097 4798 29107
rect 4938 29097 4990 29107
rect 2233 29045 2457 29097
rect 2509 29045 2650 29097
rect 2702 29045 2841 29097
rect 2893 29045 3033 29097
rect 3085 29045 3225 29097
rect 3277 29045 3417 29097
rect 3469 29045 3978 29097
rect 4030 29045 4171 29097
rect 4223 29045 4362 29097
rect 4414 29045 4554 29097
rect 4606 29045 4746 29097
rect 4798 29045 4938 29097
rect 4990 29045 5846 29097
rect 2457 29035 2509 29045
rect 2650 29035 2702 29045
rect 2841 29035 2893 29045
rect 3033 29035 3085 29045
rect 3225 29035 3277 29045
rect 3417 29035 3469 29045
rect 2056 28795 2190 28805
rect 2056 28557 2190 28687
rect 2056 27518 2186 28557
rect 3681 28520 3733 29045
rect 3978 29035 4030 29045
rect 4171 29035 4223 29045
rect 4362 29035 4414 29045
rect 4554 29035 4606 29045
rect 4746 29035 4798 29045
rect 4938 29035 4990 29045
rect 5336 28552 5390 28563
rect 5336 28545 5337 28552
rect 3681 28458 3733 28468
rect 5178 28500 5337 28545
rect 5389 28500 5390 28552
rect 5178 28493 5390 28500
rect 2457 28290 2509 28300
rect 2648 28290 2700 28300
rect 2840 28290 2892 28300
rect 3032 28290 3084 28300
rect 3225 28290 3277 28299
rect 3417 28290 3469 28299
rect 3978 28290 4030 28300
rect 4169 28290 4221 28300
rect 4361 28290 4413 28300
rect 4553 28290 4605 28300
rect 4746 28290 4798 28299
rect 4938 28290 4990 28299
rect 5178 28290 5230 28493
rect 5336 28489 5390 28493
rect 5448 28561 5502 28565
rect 5608 28561 5660 29045
rect 5448 28554 5660 28561
rect 5448 28502 5449 28554
rect 5501 28509 5660 28554
rect 5501 28502 5502 28509
rect 5448 28491 5502 28502
rect 2229 28238 2457 28290
rect 2509 28238 2648 28290
rect 2700 28238 2840 28290
rect 2892 28238 3032 28290
rect 3084 28289 3978 28290
rect 3084 28238 3225 28289
rect 2457 28228 2509 28238
rect 2648 28228 2700 28238
rect 2840 28228 2892 28238
rect 3032 28228 3084 28238
rect 3277 28238 3417 28289
rect 3225 28227 3277 28237
rect 3469 28238 3978 28289
rect 4030 28238 4169 28290
rect 4221 28238 4361 28290
rect 4413 28238 4553 28290
rect 4605 28289 5230 28290
rect 4605 28238 4746 28289
rect 3417 28227 3469 28237
rect 3978 28228 4030 28238
rect 4169 28228 4221 28238
rect 4361 28228 4413 28238
rect 4553 28228 4605 28238
rect 4798 28238 4938 28289
rect 4746 28227 4798 28237
rect 4990 28238 5230 28289
rect 4938 28227 4990 28237
rect 2457 27810 2509 27820
rect 2650 27810 2702 27820
rect 2841 27810 2893 27820
rect 3033 27810 3085 27820
rect 3225 27810 3277 27820
rect 3417 27810 3469 27820
rect 3978 27810 4030 27820
rect 4171 27810 4223 27820
rect 4362 27810 4414 27820
rect 4554 27810 4606 27820
rect 4746 27810 4798 27820
rect 4938 27810 4990 27820
rect 2233 27758 2457 27810
rect 2509 27758 2650 27810
rect 2702 27758 2841 27810
rect 2893 27758 3033 27810
rect 3085 27758 3225 27810
rect 3277 27758 3417 27810
rect 3469 27758 3978 27810
rect 4030 27758 4171 27810
rect 4223 27758 4362 27810
rect 4414 27758 4554 27810
rect 4606 27758 4746 27810
rect 4798 27758 4938 27810
rect 4990 27758 5846 27810
rect 2457 27748 2509 27758
rect 2650 27748 2702 27758
rect 2841 27748 2893 27758
rect 3033 27748 3085 27758
rect 3225 27748 3277 27758
rect 3417 27748 3469 27758
rect 2056 27508 2190 27518
rect 2056 27270 2190 27400
rect 2056 26231 2186 27270
rect 3681 27233 3733 27758
rect 3978 27748 4030 27758
rect 4171 27748 4223 27758
rect 4362 27748 4414 27758
rect 4554 27748 4606 27758
rect 4746 27748 4798 27758
rect 4938 27748 4990 27758
rect 5336 27265 5390 27276
rect 5336 27258 5337 27265
rect 3681 27171 3733 27181
rect 5178 27213 5337 27258
rect 5389 27213 5390 27265
rect 5178 27206 5390 27213
rect 2457 27003 2509 27013
rect 2648 27003 2700 27013
rect 2840 27003 2892 27013
rect 3032 27003 3084 27013
rect 3225 27003 3277 27012
rect 3417 27003 3469 27012
rect 3978 27003 4030 27013
rect 4169 27003 4221 27013
rect 4361 27003 4413 27013
rect 4553 27003 4605 27013
rect 4746 27003 4798 27012
rect 4938 27003 4990 27012
rect 5178 27003 5230 27206
rect 5336 27202 5390 27206
rect 5448 27274 5502 27278
rect 5608 27274 5660 27758
rect 5448 27267 5660 27274
rect 5448 27215 5449 27267
rect 5501 27222 5660 27267
rect 5501 27215 5502 27222
rect 5448 27204 5502 27215
rect 2229 26951 2457 27003
rect 2509 26951 2648 27003
rect 2700 26951 2840 27003
rect 2892 26951 3032 27003
rect 3084 27002 3978 27003
rect 3084 26951 3225 27002
rect 2457 26941 2509 26951
rect 2648 26941 2700 26951
rect 2840 26941 2892 26951
rect 3032 26941 3084 26951
rect 3277 26951 3417 27002
rect 3225 26940 3277 26950
rect 3469 26951 3978 27002
rect 4030 26951 4169 27003
rect 4221 26951 4361 27003
rect 4413 26951 4553 27003
rect 4605 27002 5230 27003
rect 4605 26951 4746 27002
rect 3417 26940 3469 26950
rect 3978 26941 4030 26951
rect 4169 26941 4221 26951
rect 4361 26941 4413 26951
rect 4553 26941 4605 26951
rect 4798 26951 4938 27002
rect 4746 26940 4798 26950
rect 4990 26951 5230 27002
rect 4938 26940 4990 26950
rect 2457 26523 2509 26533
rect 2650 26523 2702 26533
rect 2841 26523 2893 26533
rect 3033 26523 3085 26533
rect 3225 26523 3277 26533
rect 3417 26523 3469 26533
rect 3978 26523 4030 26533
rect 4171 26523 4223 26533
rect 4362 26523 4414 26533
rect 4554 26523 4606 26533
rect 4746 26523 4798 26533
rect 4938 26523 4990 26533
rect 2233 26471 2457 26523
rect 2509 26471 2650 26523
rect 2702 26471 2841 26523
rect 2893 26471 3033 26523
rect 3085 26471 3225 26523
rect 3277 26471 3417 26523
rect 3469 26471 3978 26523
rect 4030 26471 4171 26523
rect 4223 26471 4362 26523
rect 4414 26471 4554 26523
rect 4606 26471 4746 26523
rect 4798 26471 4938 26523
rect 4990 26471 5846 26523
rect 2457 26461 2509 26471
rect 2650 26461 2702 26471
rect 2841 26461 2893 26471
rect 3033 26461 3085 26471
rect 3225 26461 3277 26471
rect 3417 26461 3469 26471
rect 2056 26221 2190 26231
rect 2056 25983 2190 26113
rect 2056 24944 2186 25983
rect 3681 25946 3733 26471
rect 3978 26461 4030 26471
rect 4171 26461 4223 26471
rect 4362 26461 4414 26471
rect 4554 26461 4606 26471
rect 4746 26461 4798 26471
rect 4938 26461 4990 26471
rect 5336 25978 5390 25989
rect 5336 25971 5337 25978
rect 3681 25884 3733 25894
rect 5178 25926 5337 25971
rect 5389 25926 5390 25978
rect 5178 25919 5390 25926
rect 2457 25716 2509 25726
rect 2648 25716 2700 25726
rect 2840 25716 2892 25726
rect 3032 25716 3084 25726
rect 3225 25716 3277 25725
rect 3417 25716 3469 25725
rect 3978 25716 4030 25726
rect 4169 25716 4221 25726
rect 4361 25716 4413 25726
rect 4553 25716 4605 25726
rect 4746 25716 4798 25725
rect 4938 25716 4990 25725
rect 5178 25716 5230 25919
rect 5336 25915 5390 25919
rect 5448 25987 5502 25991
rect 5608 25987 5660 26471
rect 5448 25980 5660 25987
rect 5448 25928 5449 25980
rect 5501 25935 5660 25980
rect 5501 25928 5502 25935
rect 5448 25917 5502 25928
rect 2229 25664 2457 25716
rect 2509 25664 2648 25716
rect 2700 25664 2840 25716
rect 2892 25664 3032 25716
rect 3084 25715 3978 25716
rect 3084 25664 3225 25715
rect 2457 25654 2509 25664
rect 2648 25654 2700 25664
rect 2840 25654 2892 25664
rect 3032 25654 3084 25664
rect 3277 25664 3417 25715
rect 3225 25653 3277 25663
rect 3469 25664 3978 25715
rect 4030 25664 4169 25716
rect 4221 25664 4361 25716
rect 4413 25664 4553 25716
rect 4605 25715 5230 25716
rect 4605 25664 4746 25715
rect 3417 25653 3469 25663
rect 3978 25654 4030 25664
rect 4169 25654 4221 25664
rect 4361 25654 4413 25664
rect 4553 25654 4605 25664
rect 4798 25664 4938 25715
rect 4746 25653 4798 25663
rect 4990 25664 5230 25715
rect 4938 25653 4990 25663
rect 2457 25236 2509 25246
rect 2650 25236 2702 25246
rect 2841 25236 2893 25246
rect 3033 25236 3085 25246
rect 3225 25236 3277 25246
rect 3417 25236 3469 25246
rect 3978 25236 4030 25246
rect 4171 25236 4223 25246
rect 4362 25236 4414 25246
rect 4554 25236 4606 25246
rect 4746 25236 4798 25246
rect 4938 25236 4990 25246
rect 2233 25184 2457 25236
rect 2509 25184 2650 25236
rect 2702 25184 2841 25236
rect 2893 25184 3033 25236
rect 3085 25184 3225 25236
rect 3277 25184 3417 25236
rect 3469 25184 3978 25236
rect 4030 25184 4171 25236
rect 4223 25184 4362 25236
rect 4414 25184 4554 25236
rect 4606 25184 4746 25236
rect 4798 25184 4938 25236
rect 4990 25184 5846 25236
rect 2457 25174 2509 25184
rect 2650 25174 2702 25184
rect 2841 25174 2893 25184
rect 3033 25174 3085 25184
rect 3225 25174 3277 25184
rect 3417 25174 3469 25184
rect 2056 24934 2190 24944
rect 2056 24696 2190 24826
rect 2056 23657 2186 24696
rect 3681 24659 3733 25184
rect 3978 25174 4030 25184
rect 4171 25174 4223 25184
rect 4362 25174 4414 25184
rect 4554 25174 4606 25184
rect 4746 25174 4798 25184
rect 4938 25174 4990 25184
rect 5336 24691 5390 24702
rect 5336 24684 5337 24691
rect 3681 24597 3733 24607
rect 5178 24639 5337 24684
rect 5389 24639 5390 24691
rect 5178 24632 5390 24639
rect 2457 24429 2509 24439
rect 2648 24429 2700 24439
rect 2840 24429 2892 24439
rect 3032 24429 3084 24439
rect 3225 24429 3277 24438
rect 3417 24429 3469 24438
rect 3978 24429 4030 24439
rect 4169 24429 4221 24439
rect 4361 24429 4413 24439
rect 4553 24429 4605 24439
rect 4746 24429 4798 24438
rect 4938 24429 4990 24438
rect 5178 24429 5230 24632
rect 5336 24628 5390 24632
rect 5448 24700 5502 24704
rect 5608 24700 5660 25184
rect 5448 24693 5660 24700
rect 5448 24641 5449 24693
rect 5501 24648 5660 24693
rect 5501 24641 5502 24648
rect 5448 24630 5502 24641
rect 2229 24377 2457 24429
rect 2509 24377 2648 24429
rect 2700 24377 2840 24429
rect 2892 24377 3032 24429
rect 3084 24428 3978 24429
rect 3084 24377 3225 24428
rect 2457 24367 2509 24377
rect 2648 24367 2700 24377
rect 2840 24367 2892 24377
rect 3032 24367 3084 24377
rect 3277 24377 3417 24428
rect 3225 24366 3277 24376
rect 3469 24377 3978 24428
rect 4030 24377 4169 24429
rect 4221 24377 4361 24429
rect 4413 24377 4553 24429
rect 4605 24428 5230 24429
rect 4605 24377 4746 24428
rect 3417 24366 3469 24376
rect 3978 24367 4030 24377
rect 4169 24367 4221 24377
rect 4361 24367 4413 24377
rect 4553 24367 4605 24377
rect 4798 24377 4938 24428
rect 4746 24366 4798 24376
rect 4990 24377 5230 24428
rect 4938 24366 4990 24376
rect 2457 23949 2509 23959
rect 2650 23949 2702 23959
rect 2841 23949 2893 23959
rect 3033 23949 3085 23959
rect 3225 23949 3277 23959
rect 3417 23949 3469 23959
rect 3978 23949 4030 23959
rect 4171 23949 4223 23959
rect 4362 23949 4414 23959
rect 4554 23949 4606 23959
rect 4746 23949 4798 23959
rect 4938 23949 4990 23959
rect 2233 23897 2457 23949
rect 2509 23897 2650 23949
rect 2702 23897 2841 23949
rect 2893 23897 3033 23949
rect 3085 23897 3225 23949
rect 3277 23897 3417 23949
rect 3469 23897 3978 23949
rect 4030 23897 4171 23949
rect 4223 23897 4362 23949
rect 4414 23897 4554 23949
rect 4606 23897 4746 23949
rect 4798 23897 4938 23949
rect 4990 23897 5846 23949
rect 2457 23887 2509 23897
rect 2650 23887 2702 23897
rect 2841 23887 2893 23897
rect 3033 23887 3085 23897
rect 3225 23887 3277 23897
rect 3417 23887 3469 23897
rect 2056 23647 2190 23657
rect 2056 23409 2190 23539
rect 2056 22370 2186 23409
rect 3681 23372 3733 23897
rect 3978 23887 4030 23897
rect 4171 23887 4223 23897
rect 4362 23887 4414 23897
rect 4554 23887 4606 23897
rect 4746 23887 4798 23897
rect 4938 23887 4990 23897
rect 5336 23404 5390 23415
rect 5336 23397 5337 23404
rect 3681 23310 3733 23320
rect 5178 23352 5337 23397
rect 5389 23352 5390 23404
rect 5178 23345 5390 23352
rect 2457 23142 2509 23152
rect 2648 23142 2700 23152
rect 2840 23142 2892 23152
rect 3032 23142 3084 23152
rect 3225 23142 3277 23151
rect 3417 23142 3469 23151
rect 3978 23142 4030 23152
rect 4169 23142 4221 23152
rect 4361 23142 4413 23152
rect 4553 23142 4605 23152
rect 4746 23142 4798 23151
rect 4938 23142 4990 23151
rect 5178 23142 5230 23345
rect 5336 23341 5390 23345
rect 5448 23413 5502 23417
rect 5608 23413 5660 23897
rect 5448 23406 5660 23413
rect 5448 23354 5449 23406
rect 5501 23361 5660 23406
rect 5501 23354 5502 23361
rect 5448 23343 5502 23354
rect 2229 23090 2457 23142
rect 2509 23090 2648 23142
rect 2700 23090 2840 23142
rect 2892 23090 3032 23142
rect 3084 23141 3978 23142
rect 3084 23090 3225 23141
rect 2457 23080 2509 23090
rect 2648 23080 2700 23090
rect 2840 23080 2892 23090
rect 3032 23080 3084 23090
rect 3277 23090 3417 23141
rect 3225 23079 3277 23089
rect 3469 23090 3978 23141
rect 4030 23090 4169 23142
rect 4221 23090 4361 23142
rect 4413 23090 4553 23142
rect 4605 23141 5230 23142
rect 4605 23090 4746 23141
rect 3417 23079 3469 23089
rect 3978 23080 4030 23090
rect 4169 23080 4221 23090
rect 4361 23080 4413 23090
rect 4553 23080 4605 23090
rect 4798 23090 4938 23141
rect 4746 23079 4798 23089
rect 4990 23090 5230 23141
rect 4938 23079 4990 23089
rect 2457 22662 2509 22672
rect 2650 22662 2702 22672
rect 2841 22662 2893 22672
rect 3033 22662 3085 22672
rect 3225 22662 3277 22672
rect 3417 22662 3469 22672
rect 3978 22662 4030 22672
rect 4171 22662 4223 22672
rect 4362 22662 4414 22672
rect 4554 22662 4606 22672
rect 4746 22662 4798 22672
rect 4938 22662 4990 22672
rect 2233 22610 2457 22662
rect 2509 22610 2650 22662
rect 2702 22610 2841 22662
rect 2893 22610 3033 22662
rect 3085 22610 3225 22662
rect 3277 22610 3417 22662
rect 3469 22610 3978 22662
rect 4030 22610 4171 22662
rect 4223 22610 4362 22662
rect 4414 22610 4554 22662
rect 4606 22610 4746 22662
rect 4798 22610 4938 22662
rect 4990 22610 5846 22662
rect 2457 22600 2509 22610
rect 2650 22600 2702 22610
rect 2841 22600 2893 22610
rect 3033 22600 3085 22610
rect 3225 22600 3277 22610
rect 3417 22600 3469 22610
rect 2056 22360 2190 22370
rect 2056 22122 2190 22252
rect 2056 21083 2186 22122
rect 3681 22085 3733 22610
rect 3978 22600 4030 22610
rect 4171 22600 4223 22610
rect 4362 22600 4414 22610
rect 4554 22600 4606 22610
rect 4746 22600 4798 22610
rect 4938 22600 4990 22610
rect 5336 22117 5390 22128
rect 5336 22110 5337 22117
rect 3681 22023 3733 22033
rect 5178 22065 5337 22110
rect 5389 22065 5390 22117
rect 5178 22058 5390 22065
rect 2457 21855 2509 21865
rect 2648 21855 2700 21865
rect 2840 21855 2892 21865
rect 3032 21855 3084 21865
rect 3225 21855 3277 21864
rect 3417 21855 3469 21864
rect 3978 21855 4030 21865
rect 4169 21855 4221 21865
rect 4361 21855 4413 21865
rect 4553 21855 4605 21865
rect 4746 21855 4798 21864
rect 4938 21855 4990 21864
rect 5178 21855 5230 22058
rect 5336 22054 5390 22058
rect 5448 22126 5502 22130
rect 5608 22126 5660 22610
rect 5448 22119 5660 22126
rect 5448 22067 5449 22119
rect 5501 22074 5660 22119
rect 5501 22067 5502 22074
rect 5448 22056 5502 22067
rect 2229 21803 2457 21855
rect 2509 21803 2648 21855
rect 2700 21803 2840 21855
rect 2892 21803 3032 21855
rect 3084 21854 3978 21855
rect 3084 21803 3225 21854
rect 2457 21793 2509 21803
rect 2648 21793 2700 21803
rect 2840 21793 2892 21803
rect 3032 21793 3084 21803
rect 3277 21803 3417 21854
rect 3225 21792 3277 21802
rect 3469 21803 3978 21854
rect 4030 21803 4169 21855
rect 4221 21803 4361 21855
rect 4413 21803 4553 21855
rect 4605 21854 5230 21855
rect 4605 21803 4746 21854
rect 3417 21792 3469 21802
rect 3978 21793 4030 21803
rect 4169 21793 4221 21803
rect 4361 21793 4413 21803
rect 4553 21793 4605 21803
rect 4798 21803 4938 21854
rect 4746 21792 4798 21802
rect 4990 21803 5230 21854
rect 4938 21792 4990 21802
rect 2457 21375 2509 21385
rect 2650 21375 2702 21385
rect 2841 21375 2893 21385
rect 3033 21375 3085 21385
rect 3225 21375 3277 21385
rect 3417 21375 3469 21385
rect 3978 21375 4030 21385
rect 4171 21375 4223 21385
rect 4362 21375 4414 21385
rect 4554 21375 4606 21385
rect 4746 21375 4798 21385
rect 4938 21375 4990 21385
rect 2233 21323 2457 21375
rect 2509 21323 2650 21375
rect 2702 21323 2841 21375
rect 2893 21323 3033 21375
rect 3085 21323 3225 21375
rect 3277 21323 3417 21375
rect 3469 21323 3978 21375
rect 4030 21323 4171 21375
rect 4223 21323 4362 21375
rect 4414 21323 4554 21375
rect 4606 21323 4746 21375
rect 4798 21323 4938 21375
rect 4990 21323 5846 21375
rect 2457 21313 2509 21323
rect 2650 21313 2702 21323
rect 2841 21313 2893 21323
rect 3033 21313 3085 21323
rect 3225 21313 3277 21323
rect 3417 21313 3469 21323
rect 2056 21073 2190 21083
rect 2056 20835 2190 20965
rect 2056 19796 2186 20835
rect 3681 20798 3733 21323
rect 3978 21313 4030 21323
rect 4171 21313 4223 21323
rect 4362 21313 4414 21323
rect 4554 21313 4606 21323
rect 4746 21313 4798 21323
rect 4938 21313 4990 21323
rect 5336 20830 5390 20841
rect 5336 20823 5337 20830
rect 3681 20736 3733 20746
rect 5178 20778 5337 20823
rect 5389 20778 5390 20830
rect 5178 20771 5390 20778
rect 2457 20568 2509 20578
rect 2648 20568 2700 20578
rect 2840 20568 2892 20578
rect 3032 20568 3084 20578
rect 3225 20568 3277 20577
rect 3417 20568 3469 20577
rect 3978 20568 4030 20578
rect 4169 20568 4221 20578
rect 4361 20568 4413 20578
rect 4553 20568 4605 20578
rect 4746 20568 4798 20577
rect 4938 20568 4990 20577
rect 5178 20568 5230 20771
rect 5336 20767 5390 20771
rect 5448 20839 5502 20843
rect 5608 20839 5660 21323
rect 5448 20832 5660 20839
rect 5448 20780 5449 20832
rect 5501 20787 5660 20832
rect 5501 20780 5502 20787
rect 5448 20769 5502 20780
rect 2229 20516 2457 20568
rect 2509 20516 2648 20568
rect 2700 20516 2840 20568
rect 2892 20516 3032 20568
rect 3084 20567 3978 20568
rect 3084 20516 3225 20567
rect 2457 20506 2509 20516
rect 2648 20506 2700 20516
rect 2840 20506 2892 20516
rect 3032 20506 3084 20516
rect 3277 20516 3417 20567
rect 3225 20505 3277 20515
rect 3469 20516 3978 20567
rect 4030 20516 4169 20568
rect 4221 20516 4361 20568
rect 4413 20516 4553 20568
rect 4605 20567 5230 20568
rect 4605 20516 4746 20567
rect 3417 20505 3469 20515
rect 3978 20506 4030 20516
rect 4169 20506 4221 20516
rect 4361 20506 4413 20516
rect 4553 20506 4605 20516
rect 4798 20516 4938 20567
rect 4746 20505 4798 20515
rect 4990 20516 5230 20567
rect 4938 20505 4990 20515
rect 2457 20088 2509 20098
rect 2650 20088 2702 20098
rect 2841 20088 2893 20098
rect 3033 20088 3085 20098
rect 3225 20088 3277 20098
rect 3417 20088 3469 20098
rect 3978 20088 4030 20098
rect 4171 20088 4223 20098
rect 4362 20088 4414 20098
rect 4554 20088 4606 20098
rect 4746 20088 4798 20098
rect 4938 20088 4990 20098
rect 2233 20036 2457 20088
rect 2509 20036 2650 20088
rect 2702 20036 2841 20088
rect 2893 20036 3033 20088
rect 3085 20036 3225 20088
rect 3277 20036 3417 20088
rect 3469 20036 3978 20088
rect 4030 20036 4171 20088
rect 4223 20036 4362 20088
rect 4414 20036 4554 20088
rect 4606 20036 4746 20088
rect 4798 20036 4938 20088
rect 4990 20036 5846 20088
rect 2457 20026 2509 20036
rect 2650 20026 2702 20036
rect 2841 20026 2893 20036
rect 3033 20026 3085 20036
rect 3225 20026 3277 20036
rect 3417 20026 3469 20036
rect 2056 19786 2190 19796
rect 2056 19548 2190 19678
rect 2056 18509 2186 19548
rect 3681 19511 3733 20036
rect 3978 20026 4030 20036
rect 4171 20026 4223 20036
rect 4362 20026 4414 20036
rect 4554 20026 4606 20036
rect 4746 20026 4798 20036
rect 4938 20026 4990 20036
rect 5336 19543 5390 19554
rect 5336 19536 5337 19543
rect 3681 19449 3733 19459
rect 5178 19491 5337 19536
rect 5389 19491 5390 19543
rect 5178 19484 5390 19491
rect 2457 19281 2509 19291
rect 2648 19281 2700 19291
rect 2840 19281 2892 19291
rect 3032 19281 3084 19291
rect 3225 19281 3277 19290
rect 3417 19281 3469 19290
rect 3978 19281 4030 19291
rect 4169 19281 4221 19291
rect 4361 19281 4413 19291
rect 4553 19281 4605 19291
rect 4746 19281 4798 19290
rect 4938 19281 4990 19290
rect 5178 19281 5230 19484
rect 5336 19480 5390 19484
rect 5448 19552 5502 19556
rect 5608 19552 5660 20036
rect 5448 19545 5660 19552
rect 5448 19493 5449 19545
rect 5501 19500 5660 19545
rect 5501 19493 5502 19500
rect 5448 19482 5502 19493
rect 2229 19229 2457 19281
rect 2509 19229 2648 19281
rect 2700 19229 2840 19281
rect 2892 19229 3032 19281
rect 3084 19280 3978 19281
rect 3084 19229 3225 19280
rect 2457 19219 2509 19229
rect 2648 19219 2700 19229
rect 2840 19219 2892 19229
rect 3032 19219 3084 19229
rect 3277 19229 3417 19280
rect 3225 19218 3277 19228
rect 3469 19229 3978 19280
rect 4030 19229 4169 19281
rect 4221 19229 4361 19281
rect 4413 19229 4553 19281
rect 4605 19280 5230 19281
rect 4605 19229 4746 19280
rect 3417 19218 3469 19228
rect 3978 19219 4030 19229
rect 4169 19219 4221 19229
rect 4361 19219 4413 19229
rect 4553 19219 4605 19229
rect 4798 19229 4938 19280
rect 4746 19218 4798 19228
rect 4990 19229 5230 19280
rect 4938 19218 4990 19228
rect 2457 18801 2509 18811
rect 2650 18801 2702 18811
rect 2841 18801 2893 18811
rect 3033 18801 3085 18811
rect 3225 18801 3277 18811
rect 3417 18801 3469 18811
rect 3978 18801 4030 18811
rect 4171 18801 4223 18811
rect 4362 18801 4414 18811
rect 4554 18801 4606 18811
rect 4746 18801 4798 18811
rect 4938 18801 4990 18811
rect 2233 18749 2457 18801
rect 2509 18749 2650 18801
rect 2702 18749 2841 18801
rect 2893 18749 3033 18801
rect 3085 18749 3225 18801
rect 3277 18749 3417 18801
rect 3469 18749 3978 18801
rect 4030 18749 4171 18801
rect 4223 18749 4362 18801
rect 4414 18749 4554 18801
rect 4606 18749 4746 18801
rect 4798 18749 4938 18801
rect 4990 18749 5846 18801
rect 2457 18739 2509 18749
rect 2650 18739 2702 18749
rect 2841 18739 2893 18749
rect 3033 18739 3085 18749
rect 3225 18739 3277 18749
rect 3417 18739 3469 18749
rect 2056 18499 2190 18509
rect 2056 18261 2190 18391
rect 2056 17222 2186 18261
rect 3681 18224 3733 18749
rect 3978 18739 4030 18749
rect 4171 18739 4223 18749
rect 4362 18739 4414 18749
rect 4554 18739 4606 18749
rect 4746 18739 4798 18749
rect 4938 18739 4990 18749
rect 5336 18256 5390 18267
rect 5336 18249 5337 18256
rect 3681 18162 3733 18172
rect 5178 18204 5337 18249
rect 5389 18204 5390 18256
rect 5178 18197 5390 18204
rect 2457 17994 2509 18004
rect 2648 17994 2700 18004
rect 2840 17994 2892 18004
rect 3032 17994 3084 18004
rect 3225 17994 3277 18003
rect 3417 17994 3469 18003
rect 3978 17994 4030 18004
rect 4169 17994 4221 18004
rect 4361 17994 4413 18004
rect 4553 17994 4605 18004
rect 4746 17994 4798 18003
rect 4938 17994 4990 18003
rect 5178 17994 5230 18197
rect 5336 18193 5390 18197
rect 5448 18265 5502 18269
rect 5608 18265 5660 18749
rect 5448 18258 5660 18265
rect 5448 18206 5449 18258
rect 5501 18213 5660 18258
rect 5501 18206 5502 18213
rect 5448 18195 5502 18206
rect 2229 17942 2457 17994
rect 2509 17942 2648 17994
rect 2700 17942 2840 17994
rect 2892 17942 3032 17994
rect 3084 17993 3978 17994
rect 3084 17942 3225 17993
rect 2457 17932 2509 17942
rect 2648 17932 2700 17942
rect 2840 17932 2892 17942
rect 3032 17932 3084 17942
rect 3277 17942 3417 17993
rect 3225 17931 3277 17941
rect 3469 17942 3978 17993
rect 4030 17942 4169 17994
rect 4221 17942 4361 17994
rect 4413 17942 4553 17994
rect 4605 17993 5230 17994
rect 4605 17942 4746 17993
rect 3417 17931 3469 17941
rect 3978 17932 4030 17942
rect 4169 17932 4221 17942
rect 4361 17932 4413 17942
rect 4553 17932 4605 17942
rect 4798 17942 4938 17993
rect 4746 17931 4798 17941
rect 4990 17942 5230 17993
rect 4938 17931 4990 17941
rect 2457 17514 2509 17524
rect 2650 17514 2702 17524
rect 2841 17514 2893 17524
rect 3033 17514 3085 17524
rect 3225 17514 3277 17524
rect 3417 17514 3469 17524
rect 3978 17514 4030 17524
rect 4171 17514 4223 17524
rect 4362 17514 4414 17524
rect 4554 17514 4606 17524
rect 4746 17514 4798 17524
rect 4938 17514 4990 17524
rect 2233 17462 2457 17514
rect 2509 17462 2650 17514
rect 2702 17462 2841 17514
rect 2893 17462 3033 17514
rect 3085 17462 3225 17514
rect 3277 17462 3417 17514
rect 3469 17462 3978 17514
rect 4030 17462 4171 17514
rect 4223 17462 4362 17514
rect 4414 17462 4554 17514
rect 4606 17462 4746 17514
rect 4798 17462 4938 17514
rect 4990 17462 5846 17514
rect 2457 17452 2509 17462
rect 2650 17452 2702 17462
rect 2841 17452 2893 17462
rect 3033 17452 3085 17462
rect 3225 17452 3277 17462
rect 3417 17452 3469 17462
rect 2056 17212 2190 17222
rect 2056 16974 2190 17104
rect 2056 15935 2186 16974
rect 3681 16937 3733 17462
rect 3978 17452 4030 17462
rect 4171 17452 4223 17462
rect 4362 17452 4414 17462
rect 4554 17452 4606 17462
rect 4746 17452 4798 17462
rect 4938 17452 4990 17462
rect 5336 16969 5390 16980
rect 5336 16962 5337 16969
rect 3681 16875 3733 16885
rect 5178 16917 5337 16962
rect 5389 16917 5390 16969
rect 5178 16910 5390 16917
rect 2457 16707 2509 16717
rect 2648 16707 2700 16717
rect 2840 16707 2892 16717
rect 3032 16707 3084 16717
rect 3225 16707 3277 16716
rect 3417 16707 3469 16716
rect 3978 16707 4030 16717
rect 4169 16707 4221 16717
rect 4361 16707 4413 16717
rect 4553 16707 4605 16717
rect 4746 16707 4798 16716
rect 4938 16707 4990 16716
rect 5178 16707 5230 16910
rect 5336 16906 5390 16910
rect 5448 16978 5502 16982
rect 5608 16978 5660 17462
rect 5448 16971 5660 16978
rect 5448 16919 5449 16971
rect 5501 16926 5660 16971
rect 5501 16919 5502 16926
rect 5448 16908 5502 16919
rect 2229 16655 2457 16707
rect 2509 16655 2648 16707
rect 2700 16655 2840 16707
rect 2892 16655 3032 16707
rect 3084 16706 3978 16707
rect 3084 16655 3225 16706
rect 2457 16645 2509 16655
rect 2648 16645 2700 16655
rect 2840 16645 2892 16655
rect 3032 16645 3084 16655
rect 3277 16655 3417 16706
rect 3225 16644 3277 16654
rect 3469 16655 3978 16706
rect 4030 16655 4169 16707
rect 4221 16655 4361 16707
rect 4413 16655 4553 16707
rect 4605 16706 5230 16707
rect 4605 16655 4746 16706
rect 3417 16644 3469 16654
rect 3978 16645 4030 16655
rect 4169 16645 4221 16655
rect 4361 16645 4413 16655
rect 4553 16645 4605 16655
rect 4798 16655 4938 16706
rect 4746 16644 4798 16654
rect 4990 16655 5230 16706
rect 4938 16644 4990 16654
rect 2457 16227 2509 16237
rect 2650 16227 2702 16237
rect 2841 16227 2893 16237
rect 3033 16227 3085 16237
rect 3225 16227 3277 16237
rect 3417 16227 3469 16237
rect 3978 16227 4030 16237
rect 4171 16227 4223 16237
rect 4362 16227 4414 16237
rect 4554 16227 4606 16237
rect 4746 16227 4798 16237
rect 4938 16227 4990 16237
rect 2233 16175 2457 16227
rect 2509 16175 2650 16227
rect 2702 16175 2841 16227
rect 2893 16175 3033 16227
rect 3085 16175 3225 16227
rect 3277 16175 3417 16227
rect 3469 16175 3978 16227
rect 4030 16175 4171 16227
rect 4223 16175 4362 16227
rect 4414 16175 4554 16227
rect 4606 16175 4746 16227
rect 4798 16175 4938 16227
rect 4990 16175 5846 16227
rect 2457 16165 2509 16175
rect 2650 16165 2702 16175
rect 2841 16165 2893 16175
rect 3033 16165 3085 16175
rect 3225 16165 3277 16175
rect 3417 16165 3469 16175
rect 2056 15925 2190 15935
rect 2056 15687 2190 15817
rect 2056 14648 2186 15687
rect 3681 15650 3733 16175
rect 3978 16165 4030 16175
rect 4171 16165 4223 16175
rect 4362 16165 4414 16175
rect 4554 16165 4606 16175
rect 4746 16165 4798 16175
rect 4938 16165 4990 16175
rect 5336 15682 5390 15693
rect 5336 15675 5337 15682
rect 3681 15588 3733 15598
rect 5178 15630 5337 15675
rect 5389 15630 5390 15682
rect 5178 15623 5390 15630
rect 2457 15420 2509 15430
rect 2648 15420 2700 15430
rect 2840 15420 2892 15430
rect 3032 15420 3084 15430
rect 3225 15420 3277 15429
rect 3417 15420 3469 15429
rect 3978 15420 4030 15430
rect 4169 15420 4221 15430
rect 4361 15420 4413 15430
rect 4553 15420 4605 15430
rect 4746 15420 4798 15429
rect 4938 15420 4990 15429
rect 5178 15420 5230 15623
rect 5336 15619 5390 15623
rect 5448 15691 5502 15695
rect 5608 15691 5660 16175
rect 5448 15684 5660 15691
rect 5448 15632 5449 15684
rect 5501 15639 5660 15684
rect 5501 15632 5502 15639
rect 5448 15621 5502 15632
rect 2229 15368 2457 15420
rect 2509 15368 2648 15420
rect 2700 15368 2840 15420
rect 2892 15368 3032 15420
rect 3084 15419 3978 15420
rect 3084 15368 3225 15419
rect 2457 15358 2509 15368
rect 2648 15358 2700 15368
rect 2840 15358 2892 15368
rect 3032 15358 3084 15368
rect 3277 15368 3417 15419
rect 3225 15357 3277 15367
rect 3469 15368 3978 15419
rect 4030 15368 4169 15420
rect 4221 15368 4361 15420
rect 4413 15368 4553 15420
rect 4605 15419 5230 15420
rect 4605 15368 4746 15419
rect 3417 15357 3469 15367
rect 3978 15358 4030 15368
rect 4169 15358 4221 15368
rect 4361 15358 4413 15368
rect 4553 15358 4605 15368
rect 4798 15368 4938 15419
rect 4746 15357 4798 15367
rect 4990 15368 5230 15419
rect 4938 15357 4990 15367
rect 2457 14940 2509 14950
rect 2650 14940 2702 14950
rect 2841 14940 2893 14950
rect 3033 14940 3085 14950
rect 3225 14940 3277 14950
rect 3417 14940 3469 14950
rect 3978 14940 4030 14950
rect 4171 14940 4223 14950
rect 4362 14940 4414 14950
rect 4554 14940 4606 14950
rect 4746 14940 4798 14950
rect 4938 14940 4990 14950
rect 2233 14888 2457 14940
rect 2509 14888 2650 14940
rect 2702 14888 2841 14940
rect 2893 14888 3033 14940
rect 3085 14888 3225 14940
rect 3277 14888 3417 14940
rect 3469 14888 3978 14940
rect 4030 14888 4171 14940
rect 4223 14888 4362 14940
rect 4414 14888 4554 14940
rect 4606 14888 4746 14940
rect 4798 14888 4938 14940
rect 4990 14888 5846 14940
rect 2457 14878 2509 14888
rect 2650 14878 2702 14888
rect 2841 14878 2893 14888
rect 3033 14878 3085 14888
rect 3225 14878 3277 14888
rect 3417 14878 3469 14888
rect 2056 14638 2190 14648
rect 2056 14400 2190 14530
rect 2056 13361 2186 14400
rect 3681 14363 3733 14888
rect 3978 14878 4030 14888
rect 4171 14878 4223 14888
rect 4362 14878 4414 14888
rect 4554 14878 4606 14888
rect 4746 14878 4798 14888
rect 4938 14878 4990 14888
rect 5336 14395 5390 14406
rect 5336 14388 5337 14395
rect 3681 14301 3733 14311
rect 5178 14343 5337 14388
rect 5389 14343 5390 14395
rect 5178 14336 5390 14343
rect 2457 14133 2509 14143
rect 2648 14133 2700 14143
rect 2840 14133 2892 14143
rect 3032 14133 3084 14143
rect 3225 14133 3277 14142
rect 3417 14133 3469 14142
rect 3978 14133 4030 14143
rect 4169 14133 4221 14143
rect 4361 14133 4413 14143
rect 4553 14133 4605 14143
rect 4746 14133 4798 14142
rect 4938 14133 4990 14142
rect 5178 14133 5230 14336
rect 5336 14332 5390 14336
rect 5448 14404 5502 14408
rect 5608 14404 5660 14888
rect 5448 14397 5660 14404
rect 5448 14345 5449 14397
rect 5501 14352 5660 14397
rect 5501 14345 5502 14352
rect 5448 14334 5502 14345
rect 2229 14081 2457 14133
rect 2509 14081 2648 14133
rect 2700 14081 2840 14133
rect 2892 14081 3032 14133
rect 3084 14132 3978 14133
rect 3084 14081 3225 14132
rect 2457 14071 2509 14081
rect 2648 14071 2700 14081
rect 2840 14071 2892 14081
rect 3032 14071 3084 14081
rect 3277 14081 3417 14132
rect 3225 14070 3277 14080
rect 3469 14081 3978 14132
rect 4030 14081 4169 14133
rect 4221 14081 4361 14133
rect 4413 14081 4553 14133
rect 4605 14132 5230 14133
rect 4605 14081 4746 14132
rect 3417 14070 3469 14080
rect 3978 14071 4030 14081
rect 4169 14071 4221 14081
rect 4361 14071 4413 14081
rect 4553 14071 4605 14081
rect 4798 14081 4938 14132
rect 4746 14070 4798 14080
rect 4990 14081 5230 14132
rect 4938 14070 4990 14080
rect 2457 13653 2509 13663
rect 2650 13653 2702 13663
rect 2841 13653 2893 13663
rect 3033 13653 3085 13663
rect 3225 13653 3277 13663
rect 3417 13653 3469 13663
rect 3978 13653 4030 13663
rect 4171 13653 4223 13663
rect 4362 13653 4414 13663
rect 4554 13653 4606 13663
rect 4746 13653 4798 13663
rect 4938 13653 4990 13663
rect 2233 13601 2457 13653
rect 2509 13601 2650 13653
rect 2702 13601 2841 13653
rect 2893 13601 3033 13653
rect 3085 13601 3225 13653
rect 3277 13601 3417 13653
rect 3469 13601 3978 13653
rect 4030 13601 4171 13653
rect 4223 13601 4362 13653
rect 4414 13601 4554 13653
rect 4606 13601 4746 13653
rect 4798 13601 4938 13653
rect 4990 13601 5846 13653
rect 2457 13591 2509 13601
rect 2650 13591 2702 13601
rect 2841 13591 2893 13601
rect 3033 13591 3085 13601
rect 3225 13591 3277 13601
rect 3417 13591 3469 13601
rect 2056 13351 2190 13361
rect 2056 13113 2190 13243
rect 2056 12074 2186 13113
rect 3681 13076 3733 13601
rect 3978 13591 4030 13601
rect 4171 13591 4223 13601
rect 4362 13591 4414 13601
rect 4554 13591 4606 13601
rect 4746 13591 4798 13601
rect 4938 13591 4990 13601
rect 5336 13108 5390 13119
rect 5336 13101 5337 13108
rect 3681 13014 3733 13024
rect 5178 13056 5337 13101
rect 5389 13056 5390 13108
rect 5178 13049 5390 13056
rect 2457 12846 2509 12856
rect 2648 12846 2700 12856
rect 2840 12846 2892 12856
rect 3032 12846 3084 12856
rect 3225 12846 3277 12855
rect 3417 12846 3469 12855
rect 3978 12846 4030 12856
rect 4169 12846 4221 12856
rect 4361 12846 4413 12856
rect 4553 12846 4605 12856
rect 4746 12846 4798 12855
rect 4938 12846 4990 12855
rect 5178 12846 5230 13049
rect 5336 13045 5390 13049
rect 5448 13117 5502 13121
rect 5608 13117 5660 13601
rect 5448 13110 5660 13117
rect 5448 13058 5449 13110
rect 5501 13065 5660 13110
rect 5501 13058 5502 13065
rect 5448 13047 5502 13058
rect 2229 12794 2457 12846
rect 2509 12794 2648 12846
rect 2700 12794 2840 12846
rect 2892 12794 3032 12846
rect 3084 12845 3978 12846
rect 3084 12794 3225 12845
rect 2457 12784 2509 12794
rect 2648 12784 2700 12794
rect 2840 12784 2892 12794
rect 3032 12784 3084 12794
rect 3277 12794 3417 12845
rect 3225 12783 3277 12793
rect 3469 12794 3978 12845
rect 4030 12794 4169 12846
rect 4221 12794 4361 12846
rect 4413 12794 4553 12846
rect 4605 12845 5230 12846
rect 4605 12794 4746 12845
rect 3417 12783 3469 12793
rect 3978 12784 4030 12794
rect 4169 12784 4221 12794
rect 4361 12784 4413 12794
rect 4553 12784 4605 12794
rect 4798 12794 4938 12845
rect 4746 12783 4798 12793
rect 4990 12794 5230 12845
rect 4938 12783 4990 12793
rect 2457 12366 2509 12376
rect 2650 12366 2702 12376
rect 2841 12366 2893 12376
rect 3033 12366 3085 12376
rect 3225 12366 3277 12376
rect 3417 12366 3469 12376
rect 3978 12366 4030 12376
rect 4171 12366 4223 12376
rect 4362 12366 4414 12376
rect 4554 12366 4606 12376
rect 4746 12366 4798 12376
rect 4938 12366 4990 12376
rect 2233 12314 2457 12366
rect 2509 12314 2650 12366
rect 2702 12314 2841 12366
rect 2893 12314 3033 12366
rect 3085 12314 3225 12366
rect 3277 12314 3417 12366
rect 3469 12314 3978 12366
rect 4030 12314 4171 12366
rect 4223 12314 4362 12366
rect 4414 12314 4554 12366
rect 4606 12314 4746 12366
rect 4798 12314 4938 12366
rect 4990 12314 5846 12366
rect 2457 12304 2509 12314
rect 2650 12304 2702 12314
rect 2841 12304 2893 12314
rect 3033 12304 3085 12314
rect 3225 12304 3277 12314
rect 3417 12304 3469 12314
rect 2056 12064 2190 12074
rect 2056 11826 2190 11956
rect 2056 10787 2186 11826
rect 3681 11789 3733 12314
rect 3978 12304 4030 12314
rect 4171 12304 4223 12314
rect 4362 12304 4414 12314
rect 4554 12304 4606 12314
rect 4746 12304 4798 12314
rect 4938 12304 4990 12314
rect 5336 11821 5390 11832
rect 5336 11814 5337 11821
rect 3681 11727 3733 11737
rect 5178 11769 5337 11814
rect 5389 11769 5390 11821
rect 5178 11762 5390 11769
rect 2457 11559 2509 11569
rect 2648 11559 2700 11569
rect 2840 11559 2892 11569
rect 3032 11559 3084 11569
rect 3225 11559 3277 11568
rect 3417 11559 3469 11568
rect 3978 11559 4030 11569
rect 4169 11559 4221 11569
rect 4361 11559 4413 11569
rect 4553 11559 4605 11569
rect 4746 11559 4798 11568
rect 4938 11559 4990 11568
rect 5178 11559 5230 11762
rect 5336 11758 5390 11762
rect 5448 11830 5502 11834
rect 5608 11830 5660 12314
rect 5448 11823 5660 11830
rect 5448 11771 5449 11823
rect 5501 11778 5660 11823
rect 5501 11771 5502 11778
rect 5448 11760 5502 11771
rect 2229 11507 2457 11559
rect 2509 11507 2648 11559
rect 2700 11507 2840 11559
rect 2892 11507 3032 11559
rect 3084 11558 3978 11559
rect 3084 11507 3225 11558
rect 2457 11497 2509 11507
rect 2648 11497 2700 11507
rect 2840 11497 2892 11507
rect 3032 11497 3084 11507
rect 3277 11507 3417 11558
rect 3225 11496 3277 11506
rect 3469 11507 3978 11558
rect 4030 11507 4169 11559
rect 4221 11507 4361 11559
rect 4413 11507 4553 11559
rect 4605 11558 5230 11559
rect 4605 11507 4746 11558
rect 3417 11496 3469 11506
rect 3978 11497 4030 11507
rect 4169 11497 4221 11507
rect 4361 11497 4413 11507
rect 4553 11497 4605 11507
rect 4798 11507 4938 11558
rect 4746 11496 4798 11506
rect 4990 11507 5230 11558
rect 4938 11496 4990 11506
rect 2457 11079 2509 11089
rect 2650 11079 2702 11089
rect 2841 11079 2893 11089
rect 3033 11079 3085 11089
rect 3225 11079 3277 11089
rect 3417 11079 3469 11089
rect 3978 11079 4030 11089
rect 4171 11079 4223 11089
rect 4362 11079 4414 11089
rect 4554 11079 4606 11089
rect 4746 11079 4798 11089
rect 4938 11079 4990 11089
rect 2233 11027 2457 11079
rect 2509 11027 2650 11079
rect 2702 11027 2841 11079
rect 2893 11027 3033 11079
rect 3085 11027 3225 11079
rect 3277 11027 3417 11079
rect 3469 11027 3978 11079
rect 4030 11027 4171 11079
rect 4223 11027 4362 11079
rect 4414 11027 4554 11079
rect 4606 11027 4746 11079
rect 4798 11027 4938 11079
rect 4990 11027 5846 11079
rect 2457 11017 2509 11027
rect 2650 11017 2702 11027
rect 2841 11017 2893 11027
rect 3033 11017 3085 11027
rect 3225 11017 3277 11027
rect 3417 11017 3469 11027
rect 2056 10777 2190 10787
rect 2056 10539 2190 10669
rect 2056 9500 2186 10539
rect 3681 10502 3733 11027
rect 3978 11017 4030 11027
rect 4171 11017 4223 11027
rect 4362 11017 4414 11027
rect 4554 11017 4606 11027
rect 4746 11017 4798 11027
rect 4938 11017 4990 11027
rect 5336 10534 5390 10545
rect 5336 10527 5337 10534
rect 3681 10440 3733 10450
rect 5178 10482 5337 10527
rect 5389 10482 5390 10534
rect 5178 10475 5390 10482
rect 2457 10272 2509 10282
rect 2648 10272 2700 10282
rect 2840 10272 2892 10282
rect 3032 10272 3084 10282
rect 3225 10272 3277 10281
rect 3417 10272 3469 10281
rect 3978 10272 4030 10282
rect 4169 10272 4221 10282
rect 4361 10272 4413 10282
rect 4553 10272 4605 10282
rect 4746 10272 4798 10281
rect 4938 10272 4990 10281
rect 5178 10272 5230 10475
rect 5336 10471 5390 10475
rect 5448 10543 5502 10547
rect 5608 10543 5660 11027
rect 5448 10536 5660 10543
rect 5448 10484 5449 10536
rect 5501 10491 5660 10536
rect 5501 10484 5502 10491
rect 5448 10473 5502 10484
rect 2229 10220 2457 10272
rect 2509 10220 2648 10272
rect 2700 10220 2840 10272
rect 2892 10220 3032 10272
rect 3084 10271 3978 10272
rect 3084 10220 3225 10271
rect 2457 10210 2509 10220
rect 2648 10210 2700 10220
rect 2840 10210 2892 10220
rect 3032 10210 3084 10220
rect 3277 10220 3417 10271
rect 3225 10209 3277 10219
rect 3469 10220 3978 10271
rect 4030 10220 4169 10272
rect 4221 10220 4361 10272
rect 4413 10220 4553 10272
rect 4605 10271 5230 10272
rect 4605 10220 4746 10271
rect 3417 10209 3469 10219
rect 3978 10210 4030 10220
rect 4169 10210 4221 10220
rect 4361 10210 4413 10220
rect 4553 10210 4605 10220
rect 4798 10220 4938 10271
rect 4746 10209 4798 10219
rect 4990 10220 5230 10271
rect 4938 10209 4990 10219
rect 2457 9792 2509 9802
rect 2650 9792 2702 9802
rect 2841 9792 2893 9802
rect 3033 9792 3085 9802
rect 3225 9792 3277 9802
rect 3417 9792 3469 9802
rect 3978 9792 4030 9802
rect 4171 9792 4223 9802
rect 4362 9792 4414 9802
rect 4554 9792 4606 9802
rect 4746 9792 4798 9802
rect 4938 9792 4990 9802
rect 2233 9740 2457 9792
rect 2509 9740 2650 9792
rect 2702 9740 2841 9792
rect 2893 9740 3033 9792
rect 3085 9740 3225 9792
rect 3277 9740 3417 9792
rect 3469 9740 3978 9792
rect 4030 9740 4171 9792
rect 4223 9740 4362 9792
rect 4414 9740 4554 9792
rect 4606 9740 4746 9792
rect 4798 9740 4938 9792
rect 4990 9740 5846 9792
rect 2457 9730 2509 9740
rect 2650 9730 2702 9740
rect 2841 9730 2893 9740
rect 3033 9730 3085 9740
rect 3225 9730 3277 9740
rect 3417 9730 3469 9740
rect 2056 9490 2190 9500
rect 2056 9252 2190 9382
rect 2056 8213 2186 9252
rect 3681 9215 3733 9740
rect 3978 9730 4030 9740
rect 4171 9730 4223 9740
rect 4362 9730 4414 9740
rect 4554 9730 4606 9740
rect 4746 9730 4798 9740
rect 4938 9730 4990 9740
rect 5336 9247 5390 9258
rect 5336 9240 5337 9247
rect 3681 9153 3733 9163
rect 5178 9195 5337 9240
rect 5389 9195 5390 9247
rect 5178 9188 5390 9195
rect 2457 8985 2509 8995
rect 2648 8985 2700 8995
rect 2840 8985 2892 8995
rect 3032 8985 3084 8995
rect 3225 8985 3277 8994
rect 3417 8985 3469 8994
rect 3978 8985 4030 8995
rect 4169 8985 4221 8995
rect 4361 8985 4413 8995
rect 4553 8985 4605 8995
rect 4746 8985 4798 8994
rect 4938 8985 4990 8994
rect 5178 8985 5230 9188
rect 5336 9184 5390 9188
rect 5448 9256 5502 9260
rect 5608 9256 5660 9740
rect 5448 9249 5660 9256
rect 5448 9197 5449 9249
rect 5501 9204 5660 9249
rect 5501 9197 5502 9204
rect 5448 9186 5502 9197
rect 2229 8933 2457 8985
rect 2509 8933 2648 8985
rect 2700 8933 2840 8985
rect 2892 8933 3032 8985
rect 3084 8984 3978 8985
rect 3084 8933 3225 8984
rect 2457 8923 2509 8933
rect 2648 8923 2700 8933
rect 2840 8923 2892 8933
rect 3032 8923 3084 8933
rect 3277 8933 3417 8984
rect 3225 8922 3277 8932
rect 3469 8933 3978 8984
rect 4030 8933 4169 8985
rect 4221 8933 4361 8985
rect 4413 8933 4553 8985
rect 4605 8984 5230 8985
rect 4605 8933 4746 8984
rect 3417 8922 3469 8932
rect 3978 8923 4030 8933
rect 4169 8923 4221 8933
rect 4361 8923 4413 8933
rect 4553 8923 4605 8933
rect 4798 8933 4938 8984
rect 4746 8922 4798 8932
rect 4990 8933 5230 8984
rect 4938 8922 4990 8932
rect 2457 8505 2509 8515
rect 2650 8505 2702 8515
rect 2841 8505 2893 8515
rect 3033 8505 3085 8515
rect 3225 8505 3277 8515
rect 3417 8505 3469 8515
rect 3978 8505 4030 8515
rect 4171 8505 4223 8515
rect 4362 8505 4414 8515
rect 4554 8505 4606 8515
rect 4746 8505 4798 8515
rect 4938 8505 4990 8515
rect 2233 8453 2457 8505
rect 2509 8453 2650 8505
rect 2702 8453 2841 8505
rect 2893 8453 3033 8505
rect 3085 8453 3225 8505
rect 3277 8453 3417 8505
rect 3469 8453 3978 8505
rect 4030 8453 4171 8505
rect 4223 8453 4362 8505
rect 4414 8453 4554 8505
rect 4606 8453 4746 8505
rect 4798 8453 4938 8505
rect 4990 8453 5846 8505
rect 2457 8443 2509 8453
rect 2650 8443 2702 8453
rect 2841 8443 2893 8453
rect 3033 8443 3085 8453
rect 3225 8443 3277 8453
rect 3417 8443 3469 8453
rect 2056 8203 2190 8213
rect 2056 7965 2190 8095
rect 2056 6926 2186 7965
rect 3681 7928 3733 8453
rect 3978 8443 4030 8453
rect 4171 8443 4223 8453
rect 4362 8443 4414 8453
rect 4554 8443 4606 8453
rect 4746 8443 4798 8453
rect 4938 8443 4990 8453
rect 5336 7960 5390 7971
rect 5336 7953 5337 7960
rect 3681 7866 3733 7876
rect 5178 7908 5337 7953
rect 5389 7908 5390 7960
rect 5178 7901 5390 7908
rect 2457 7698 2509 7708
rect 2648 7698 2700 7708
rect 2840 7698 2892 7708
rect 3032 7698 3084 7708
rect 3225 7698 3277 7707
rect 3417 7698 3469 7707
rect 3978 7698 4030 7708
rect 4169 7698 4221 7708
rect 4361 7698 4413 7708
rect 4553 7698 4605 7708
rect 4746 7698 4798 7707
rect 4938 7698 4990 7707
rect 5178 7698 5230 7901
rect 5336 7897 5390 7901
rect 5448 7969 5502 7973
rect 5608 7969 5660 8453
rect 5448 7962 5660 7969
rect 5448 7910 5449 7962
rect 5501 7917 5660 7962
rect 5501 7910 5502 7917
rect 5448 7899 5502 7910
rect 2229 7646 2457 7698
rect 2509 7646 2648 7698
rect 2700 7646 2840 7698
rect 2892 7646 3032 7698
rect 3084 7697 3978 7698
rect 3084 7646 3225 7697
rect 2457 7636 2509 7646
rect 2648 7636 2700 7646
rect 2840 7636 2892 7646
rect 3032 7636 3084 7646
rect 3277 7646 3417 7697
rect 3225 7635 3277 7645
rect 3469 7646 3978 7697
rect 4030 7646 4169 7698
rect 4221 7646 4361 7698
rect 4413 7646 4553 7698
rect 4605 7697 5230 7698
rect 4605 7646 4746 7697
rect 3417 7635 3469 7645
rect 3978 7636 4030 7646
rect 4169 7636 4221 7646
rect 4361 7636 4413 7646
rect 4553 7636 4605 7646
rect 4798 7646 4938 7697
rect 4746 7635 4798 7645
rect 4990 7646 5230 7697
rect 4938 7635 4990 7645
rect 2457 7218 2509 7228
rect 2650 7218 2702 7228
rect 2841 7218 2893 7228
rect 3033 7218 3085 7228
rect 3225 7218 3277 7228
rect 3417 7218 3469 7228
rect 3978 7218 4030 7228
rect 4171 7218 4223 7228
rect 4362 7218 4414 7228
rect 4554 7218 4606 7228
rect 4746 7218 4798 7228
rect 4938 7218 4990 7228
rect 2233 7166 2457 7218
rect 2509 7166 2650 7218
rect 2702 7166 2841 7218
rect 2893 7166 3033 7218
rect 3085 7166 3225 7218
rect 3277 7166 3417 7218
rect 3469 7166 3978 7218
rect 4030 7166 4171 7218
rect 4223 7166 4362 7218
rect 4414 7166 4554 7218
rect 4606 7166 4746 7218
rect 4798 7166 4938 7218
rect 4990 7166 5846 7218
rect 2457 7156 2509 7166
rect 2650 7156 2702 7166
rect 2841 7156 2893 7166
rect 3033 7156 3085 7166
rect 3225 7156 3277 7166
rect 3417 7156 3469 7166
rect 2056 6916 2190 6926
rect 2056 6678 2190 6808
rect 2056 5639 2186 6678
rect 3681 6641 3733 7166
rect 3978 7156 4030 7166
rect 4171 7156 4223 7166
rect 4362 7156 4414 7166
rect 4554 7156 4606 7166
rect 4746 7156 4798 7166
rect 4938 7156 4990 7166
rect 5336 6673 5390 6684
rect 5336 6666 5337 6673
rect 3681 6579 3733 6589
rect 5178 6621 5337 6666
rect 5389 6621 5390 6673
rect 5178 6614 5390 6621
rect 2457 6411 2509 6421
rect 2648 6411 2700 6421
rect 2840 6411 2892 6421
rect 3032 6411 3084 6421
rect 3225 6411 3277 6420
rect 3417 6411 3469 6420
rect 3978 6411 4030 6421
rect 4169 6411 4221 6421
rect 4361 6411 4413 6421
rect 4553 6411 4605 6421
rect 4746 6411 4798 6420
rect 4938 6411 4990 6420
rect 5178 6411 5230 6614
rect 5336 6610 5390 6614
rect 5448 6682 5502 6686
rect 5608 6682 5660 7166
rect 5448 6675 5660 6682
rect 5448 6623 5449 6675
rect 5501 6630 5660 6675
rect 5501 6623 5502 6630
rect 5448 6612 5502 6623
rect 2229 6359 2457 6411
rect 2509 6359 2648 6411
rect 2700 6359 2840 6411
rect 2892 6359 3032 6411
rect 3084 6410 3978 6411
rect 3084 6359 3225 6410
rect 2457 6349 2509 6359
rect 2648 6349 2700 6359
rect 2840 6349 2892 6359
rect 3032 6349 3084 6359
rect 3277 6359 3417 6410
rect 3225 6348 3277 6358
rect 3469 6359 3978 6410
rect 4030 6359 4169 6411
rect 4221 6359 4361 6411
rect 4413 6359 4553 6411
rect 4605 6410 5230 6411
rect 4605 6359 4746 6410
rect 3417 6348 3469 6358
rect 3978 6349 4030 6359
rect 4169 6349 4221 6359
rect 4361 6349 4413 6359
rect 4553 6349 4605 6359
rect 4798 6359 4938 6410
rect 4746 6348 4798 6358
rect 4990 6359 5230 6410
rect 4938 6348 4990 6358
rect 2457 5931 2509 5941
rect 2650 5931 2702 5941
rect 2841 5931 2893 5941
rect 3033 5931 3085 5941
rect 3225 5931 3277 5941
rect 3417 5931 3469 5941
rect 3978 5931 4030 5941
rect 4171 5931 4223 5941
rect 4362 5931 4414 5941
rect 4554 5931 4606 5941
rect 4746 5931 4798 5941
rect 4938 5931 4990 5941
rect 2233 5879 2457 5931
rect 2509 5879 2650 5931
rect 2702 5879 2841 5931
rect 2893 5879 3033 5931
rect 3085 5879 3225 5931
rect 3277 5879 3417 5931
rect 3469 5879 3978 5931
rect 4030 5879 4171 5931
rect 4223 5879 4362 5931
rect 4414 5879 4554 5931
rect 4606 5879 4746 5931
rect 4798 5879 4938 5931
rect 4990 5879 5846 5931
rect 2457 5869 2509 5879
rect 2650 5869 2702 5879
rect 2841 5869 2893 5879
rect 3033 5869 3085 5879
rect 3225 5869 3277 5879
rect 3417 5869 3469 5879
rect 2056 5629 2190 5639
rect 2056 5391 2190 5521
rect 2056 4352 2186 5391
rect 3681 5354 3733 5879
rect 3978 5869 4030 5879
rect 4171 5869 4223 5879
rect 4362 5869 4414 5879
rect 4554 5869 4606 5879
rect 4746 5869 4798 5879
rect 4938 5869 4990 5879
rect 5336 5386 5390 5397
rect 5336 5379 5337 5386
rect 3681 5292 3733 5302
rect 5178 5334 5337 5379
rect 5389 5334 5390 5386
rect 5178 5327 5390 5334
rect 2457 5124 2509 5134
rect 2648 5124 2700 5134
rect 2840 5124 2892 5134
rect 3032 5124 3084 5134
rect 3225 5124 3277 5133
rect 3417 5124 3469 5133
rect 3978 5124 4030 5134
rect 4169 5124 4221 5134
rect 4361 5124 4413 5134
rect 4553 5124 4605 5134
rect 4746 5124 4798 5133
rect 4938 5124 4990 5133
rect 5178 5124 5230 5327
rect 5336 5323 5390 5327
rect 5448 5395 5502 5399
rect 5608 5395 5660 5879
rect 5448 5388 5660 5395
rect 5448 5336 5449 5388
rect 5501 5343 5660 5388
rect 5501 5336 5502 5343
rect 5448 5325 5502 5336
rect 2229 5072 2457 5124
rect 2509 5072 2648 5124
rect 2700 5072 2840 5124
rect 2892 5072 3032 5124
rect 3084 5123 3978 5124
rect 3084 5072 3225 5123
rect 2457 5062 2509 5072
rect 2648 5062 2700 5072
rect 2840 5062 2892 5072
rect 3032 5062 3084 5072
rect 3277 5072 3417 5123
rect 3225 5061 3277 5071
rect 3469 5072 3978 5123
rect 4030 5072 4169 5124
rect 4221 5072 4361 5124
rect 4413 5072 4553 5124
rect 4605 5123 5230 5124
rect 4605 5072 4746 5123
rect 3417 5061 3469 5071
rect 3978 5062 4030 5072
rect 4169 5062 4221 5072
rect 4361 5062 4413 5072
rect 4553 5062 4605 5072
rect 4798 5072 4938 5123
rect 4746 5061 4798 5071
rect 4990 5072 5230 5123
rect 4938 5061 4990 5071
rect 2457 4644 2509 4654
rect 2650 4644 2702 4654
rect 2841 4644 2893 4654
rect 3033 4644 3085 4654
rect 3225 4644 3277 4654
rect 3417 4644 3469 4654
rect 3978 4644 4030 4654
rect 4171 4644 4223 4654
rect 4362 4644 4414 4654
rect 4554 4644 4606 4654
rect 4746 4644 4798 4654
rect 4938 4644 4990 4654
rect 2233 4592 2457 4644
rect 2509 4592 2650 4644
rect 2702 4592 2841 4644
rect 2893 4592 3033 4644
rect 3085 4592 3225 4644
rect 3277 4592 3417 4644
rect 3469 4592 3978 4644
rect 4030 4592 4171 4644
rect 4223 4592 4362 4644
rect 4414 4592 4554 4644
rect 4606 4592 4746 4644
rect 4798 4592 4938 4644
rect 4990 4592 5846 4644
rect 2457 4582 2509 4592
rect 2650 4582 2702 4592
rect 2841 4582 2893 4592
rect 3033 4582 3085 4592
rect 3225 4582 3277 4592
rect 3417 4582 3469 4592
rect 2056 4342 2190 4352
rect 2056 4104 2190 4234
rect 2056 3065 2186 4104
rect 3681 4067 3733 4592
rect 3978 4582 4030 4592
rect 4171 4582 4223 4592
rect 4362 4582 4414 4592
rect 4554 4582 4606 4592
rect 4746 4582 4798 4592
rect 4938 4582 4990 4592
rect 5336 4099 5390 4110
rect 5336 4092 5337 4099
rect 3681 4005 3733 4015
rect 5178 4047 5337 4092
rect 5389 4047 5390 4099
rect 5178 4040 5390 4047
rect 2457 3837 2509 3847
rect 2648 3837 2700 3847
rect 2840 3837 2892 3847
rect 3032 3837 3084 3847
rect 3225 3837 3277 3846
rect 3417 3837 3469 3846
rect 3978 3837 4030 3847
rect 4169 3837 4221 3847
rect 4361 3837 4413 3847
rect 4553 3837 4605 3847
rect 4746 3837 4798 3846
rect 4938 3837 4990 3846
rect 5178 3837 5230 4040
rect 5336 4036 5390 4040
rect 5448 4108 5502 4112
rect 5608 4108 5660 4592
rect 5448 4101 5660 4108
rect 5448 4049 5449 4101
rect 5501 4056 5660 4101
rect 5501 4049 5502 4056
rect 5448 4038 5502 4049
rect 2229 3785 2457 3837
rect 2509 3785 2648 3837
rect 2700 3785 2840 3837
rect 2892 3785 3032 3837
rect 3084 3836 3978 3837
rect 3084 3785 3225 3836
rect 2457 3775 2509 3785
rect 2648 3775 2700 3785
rect 2840 3775 2892 3785
rect 3032 3775 3084 3785
rect 3277 3785 3417 3836
rect 3225 3774 3277 3784
rect 3469 3785 3978 3836
rect 4030 3785 4169 3837
rect 4221 3785 4361 3837
rect 4413 3785 4553 3837
rect 4605 3836 5230 3837
rect 4605 3785 4746 3836
rect 3417 3774 3469 3784
rect 3978 3775 4030 3785
rect 4169 3775 4221 3785
rect 4361 3775 4413 3785
rect 4553 3775 4605 3785
rect 4798 3785 4938 3836
rect 4746 3774 4798 3784
rect 4990 3785 5230 3836
rect 4938 3774 4990 3784
rect 2457 3357 2509 3367
rect 2650 3357 2702 3367
rect 2841 3357 2893 3367
rect 3033 3357 3085 3367
rect 3225 3357 3277 3367
rect 3417 3357 3469 3367
rect 3978 3357 4030 3367
rect 4171 3357 4223 3367
rect 4362 3357 4414 3367
rect 4554 3357 4606 3367
rect 4746 3357 4798 3367
rect 4938 3357 4990 3367
rect 2233 3305 2457 3357
rect 2509 3305 2650 3357
rect 2702 3305 2841 3357
rect 2893 3305 3033 3357
rect 3085 3305 3225 3357
rect 3277 3305 3417 3357
rect 3469 3305 3978 3357
rect 4030 3305 4171 3357
rect 4223 3305 4362 3357
rect 4414 3305 4554 3357
rect 4606 3305 4746 3357
rect 4798 3305 4938 3357
rect 4990 3305 5846 3357
rect 2457 3295 2509 3305
rect 2650 3295 2702 3305
rect 2841 3295 2893 3305
rect 3033 3295 3085 3305
rect 3225 3295 3277 3305
rect 3417 3295 3469 3305
rect 2056 3055 2190 3065
rect 2056 2817 2190 2947
rect 2056 1778 2186 2817
rect 3681 2780 3733 3305
rect 3978 3295 4030 3305
rect 4171 3295 4223 3305
rect 4362 3295 4414 3305
rect 4554 3295 4606 3305
rect 4746 3295 4798 3305
rect 4938 3295 4990 3305
rect 5336 2812 5390 2823
rect 5336 2805 5337 2812
rect 3681 2718 3733 2728
rect 5178 2760 5337 2805
rect 5389 2760 5390 2812
rect 5178 2753 5390 2760
rect 2457 2550 2509 2560
rect 2648 2550 2700 2560
rect 2840 2550 2892 2560
rect 3032 2550 3084 2560
rect 3225 2550 3277 2559
rect 3417 2550 3469 2559
rect 3978 2550 4030 2560
rect 4169 2550 4221 2560
rect 4361 2550 4413 2560
rect 4553 2550 4605 2560
rect 4746 2550 4798 2559
rect 4938 2550 4990 2559
rect 5178 2550 5230 2753
rect 5336 2749 5390 2753
rect 5448 2821 5502 2825
rect 5608 2821 5660 3305
rect 5448 2814 5660 2821
rect 5448 2762 5449 2814
rect 5501 2769 5660 2814
rect 5501 2762 5502 2769
rect 5448 2751 5502 2762
rect 2229 2498 2457 2550
rect 2509 2498 2648 2550
rect 2700 2498 2840 2550
rect 2892 2498 3032 2550
rect 3084 2549 3978 2550
rect 3084 2498 3225 2549
rect 2457 2488 2509 2498
rect 2648 2488 2700 2498
rect 2840 2488 2892 2498
rect 3032 2488 3084 2498
rect 3277 2498 3417 2549
rect 3225 2487 3277 2497
rect 3469 2498 3978 2549
rect 4030 2498 4169 2550
rect 4221 2498 4361 2550
rect 4413 2498 4553 2550
rect 4605 2549 5230 2550
rect 4605 2498 4746 2549
rect 3417 2487 3469 2497
rect 3978 2488 4030 2498
rect 4169 2488 4221 2498
rect 4361 2488 4413 2498
rect 4553 2488 4605 2498
rect 4798 2498 4938 2549
rect 4746 2487 4798 2497
rect 4990 2498 5230 2549
rect 4938 2487 4990 2497
rect 2457 2070 2509 2080
rect 2650 2070 2702 2080
rect 2841 2070 2893 2080
rect 3033 2070 3085 2080
rect 3225 2070 3277 2080
rect 3417 2070 3469 2080
rect 3978 2070 4030 2080
rect 4171 2070 4223 2080
rect 4362 2070 4414 2080
rect 4554 2070 4606 2080
rect 4746 2070 4798 2080
rect 4938 2070 4990 2080
rect 2233 2018 2457 2070
rect 2509 2018 2650 2070
rect 2702 2018 2841 2070
rect 2893 2018 3033 2070
rect 3085 2018 3225 2070
rect 3277 2018 3417 2070
rect 3469 2018 3978 2070
rect 4030 2018 4171 2070
rect 4223 2018 4362 2070
rect 4414 2018 4554 2070
rect 4606 2018 4746 2070
rect 4798 2018 4938 2070
rect 4990 2018 5846 2070
rect 2457 2008 2509 2018
rect 2650 2008 2702 2018
rect 2841 2008 2893 2018
rect 3033 2008 3085 2018
rect 3225 2008 3277 2018
rect 3417 2008 3469 2018
rect 2056 1768 2190 1778
rect 2056 1618 2190 1660
rect 3681 1493 3733 2018
rect 3978 2008 4030 2018
rect 4171 2008 4223 2018
rect 4362 2008 4414 2018
rect 4554 2008 4606 2018
rect 4746 2008 4798 2018
rect 4938 2008 4990 2018
rect 5336 1525 5390 1536
rect 5336 1518 5337 1525
rect 3681 1431 3733 1441
rect 5178 1473 5337 1518
rect 5389 1473 5390 1525
rect 5178 1466 5390 1473
rect 2457 1263 2509 1273
rect 2648 1263 2700 1273
rect 2840 1263 2892 1273
rect 3032 1263 3084 1273
rect 3225 1263 3277 1272
rect 3417 1263 3469 1272
rect 3978 1263 4030 1273
rect 4169 1263 4221 1273
rect 4361 1263 4413 1273
rect 4553 1263 4605 1273
rect 4746 1263 4798 1272
rect 4938 1263 4990 1272
rect 5178 1263 5230 1466
rect 5336 1462 5390 1466
rect 5448 1534 5502 1538
rect 5608 1534 5660 2018
rect 5448 1527 5660 1534
rect 5448 1475 5449 1527
rect 5501 1482 5660 1527
rect 5501 1475 5502 1482
rect 5448 1464 5502 1475
rect 2270 1211 2457 1263
rect 2509 1211 2648 1263
rect 2700 1211 2840 1263
rect 2892 1211 3032 1263
rect 3084 1262 3978 1263
rect 3084 1211 3225 1262
rect 1930 1202 1986 1208
rect 2457 1201 2509 1211
rect 2648 1201 2700 1211
rect 2840 1201 2892 1211
rect 3032 1201 3084 1211
rect 3277 1211 3417 1262
rect 3225 1200 3277 1210
rect 3469 1211 3978 1262
rect 4030 1211 4169 1263
rect 4221 1211 4361 1263
rect 4413 1211 4553 1263
rect 4605 1262 5230 1263
rect 4605 1211 4746 1262
rect 3417 1200 3469 1210
rect 3978 1201 4030 1211
rect 4169 1201 4221 1211
rect 4361 1201 4413 1211
rect 4553 1201 4605 1211
rect 4798 1211 4938 1262
rect 4746 1200 4798 1210
rect 4990 1211 5230 1262
rect 4938 1200 4990 1210
<< labels >>
flabel metal1 5724 41380 5882 41516 1 FreeSans 480 0 0 0 out
port 1 n signal bidirectional
flabel metal2 5794 2018 5846 2070 1 FreeSans 480 0 0 0 en31_b
port 2 n signal bidirectional
flabel metal1 0 1527 34 1561 1 FreeSans 480 0 0 0 in_31
port 3 n signal bidirectional
flabel metal2 5794 3305 5846 3357 1 FreeSans 480 0 0 0 en30_b
port 4 n signal bidirectional
flabel metal1 0 2814 34 2848 1 FreeSans 480 0 0 0 in_30
port 5 n signal bidirectional
flabel metal2 5794 4592 5846 4644 1 FreeSans 480 0 0 0 en29_b
port 6 n signal bidirectional
flabel metal1 0 4101 34 4135 1 FreeSans 480 0 0 0 in_29
port 7 n signal bidirectional
flabel metal2 5794 5879 5846 5931 1 FreeSans 480 0 0 0 en28_b
port 8 n signal bidirectional
flabel metal1 0 5388 34 5422 1 FreeSans 480 0 0 0 in_28
port 9 n signal bidirectional
flabel metal2 5794 7166 5846 7218 1 FreeSans 480 0 0 0 en27_b
port 10 n signal bidirectional
flabel metal1 0 6675 34 6709 1 FreeSans 480 0 0 0 in_27
port 11 n signal bidirectional
flabel metal2 5794 8453 5846 8505 1 FreeSans 480 0 0 0 en26_b
port 12 n signal bidirectional
flabel metal1 0 7962 34 7996 1 FreeSans 480 0 0 0 in_26
port 13 n signal bidirectional
flabel metal2 5794 9740 5846 9792 1 FreeSans 480 0 0 0 en25_b
port 14 n signal bidirectional
flabel metal1 0 9249 34 9283 1 FreeSans 480 0 0 0 in_25
port 15 n signal bidirectional
flabel metal2 5794 11027 5846 11079 1 FreeSans 480 0 0 0 en24_b
port 16 n signal bidirectional
flabel metal1 0 10536 34 10570 1 FreeSans 480 0 0 0 in_24
port 17 n signal bidirectional
flabel metal2 5794 12314 5846 12366 1 FreeSans 480 0 0 0 en23_b
port 18 n signal bidirectional
flabel metal1 0 11823 34 11857 1 FreeSans 480 0 0 0 in_23
port 19 n signal bidirectional
flabel metal2 5794 13601 5846 13653 1 FreeSans 480 0 0 0 en22_b
port 20 n signal bidirectional
flabel metal1 0 13110 34 13144 1 FreeSans 480 0 0 0 in_22
port 21 n signal bidirectional
flabel metal2 5794 14888 5846 14940 1 FreeSans 480 0 0 0 en21_b
port 22 n signal bidirectional
flabel metal1 0 14397 34 14431 1 FreeSans 480 0 0 0 in_21
port 23 n signal bidirectional
flabel metal2 5794 16175 5846 16227 1 FreeSans 480 0 0 0 en20_b
port 24 n signal bidirectional
flabel metal1 0 15684 34 15718 1 FreeSans 480 0 0 0 in_20
port 25 n signal bidirectional
flabel metal2 5794 17462 5846 17514 1 FreeSans 480 0 0 0 en19_b
port 26 n signal bidirectional
flabel metal1 0 16971 34 17005 1 FreeSans 480 0 0 0 in_19
port 27 n signal bidirectional
flabel metal2 5794 18749 5846 18801 1 FreeSans 480 0 0 0 en18_b
port 28 n signal bidirectional
flabel metal1 0 18258 34 18292 1 FreeSans 480 0 0 0 in_18
port 29 n signal bidirectional
flabel metal2 5794 20036 5846 20088 1 FreeSans 480 0 0 0 en17_b
port 30 n signal bidirectional
flabel metal1 0 19545 34 19579 1 FreeSans 480 0 0 0 in_17
port 31 n signal bidirectional
flabel metal2 5794 21323 5846 21375 1 FreeSans 480 0 0 0 en16_b
port 32 n signal bidirectional
flabel metal1 0 20832 34 20866 1 FreeSans 480 0 0 0 in_16
port 33 n signal bidirectional
flabel metal2 5794 22610 5846 22662 1 FreeSans 480 0 0 0 en15_b
port 34 n signal bidirectional
flabel metal1 0 22119 34 22153 1 FreeSans 480 0 0 0 in_15
port 35 n signal bidirectional
flabel metal2 5794 23897 5846 23949 1 FreeSans 480 0 0 0 en14_b
port 36 n signal bidirectional
flabel metal1 0 23406 34 23440 1 FreeSans 480 0 0 0 in_14
port 37 n signal bidirectional
flabel metal2 5794 25184 5846 25236 1 FreeSans 480 0 0 0 en13_b
port 38 n signal bidirectional
flabel metal1 0 24693 34 24727 1 FreeSans 480 0 0 0 in_13
port 39 n signal bidirectional
flabel metal2 5794 26471 5846 26523 1 FreeSans 480 0 0 0 en12_b
port 40 n signal bidirectional
flabel metal1 0 25980 34 26014 1 FreeSans 480 0 0 0 in_12
port 41 n signal bidirectional
flabel metal2 5794 27758 5846 27810 1 FreeSans 480 0 0 0 en11_b
port 42 n signal bidirectional
flabel metal1 0 27267 34 27301 1 FreeSans 480 0 0 0 in_11
port 43 n signal bidirectional
flabel metal2 5794 29045 5846 29097 1 FreeSans 480 0 0 0 en10_b
port 44 n signal bidirectional
flabel metal1 0 28554 34 28588 1 FreeSans 480 0 0 0 in_10
port 45 n signal bidirectional
flabel metal2 5794 30332 5846 30384 1 FreeSans 480 0 0 0 en9_b
port 46 n signal bidirectional
flabel metal1 0 29841 34 29875 1 FreeSans 480 0 0 0 in_9
port 47 n signal bidirectional
flabel metal2 5794 31619 5846 31671 1 FreeSans 480 0 0 0 en8_b
port 48 n signal bidirectional
flabel metal1 0 31128 34 31162 1 FreeSans 480 0 0 0 in_8
port 49 n signal bidirectional
flabel metal2 5794 32906 5846 32958 1 FreeSans 480 0 0 0 en7_b
port 50 n signal bidirectional
flabel metal1 0 32415 34 32449 1 FreeSans 480 0 0 0 in_7
port 51 n signal bidirectional
flabel metal2 5794 34193 5846 34245 1 FreeSans 480 0 0 0 en6_b
port 52 n signal bidirectional
flabel metal1 0 33702 34 33736 1 FreeSans 480 0 0 0 in_6
port 53 n signal bidirectional
flabel metal2 5794 35480 5846 35532 1 FreeSans 480 0 0 0 en5_b
port 54 n signal bidirectional
flabel metal1 0 34989 34 35023 1 FreeSans 480 0 0 0 in_5
port 55 n signal bidirectional
flabel metal2 5794 36767 5846 36819 1 FreeSans 480 0 0 0 en4_b
port 56 n signal bidirectional
flabel metal1 0 36276 34 36310 1 FreeSans 480 0 0 0 in_4
port 57 n signal bidirectional
flabel metal2 5794 38054 5846 38106 1 FreeSans 480 0 0 0 en3_b
port 58 n signal bidirectional
flabel metal1 0 37563 34 37597 1 FreeSans 480 0 0 0 in_3
port 59 n signal bidirectional
flabel metal2 5794 39341 5846 39393 1 FreeSans 480 0 0 0 en2_b
port 60 n signal bidirectional
flabel metal1 0 38850 34 38884 1 FreeSans 480 0 0 0 in_2
port 61 n signal bidirectional
flabel metal2 5794 40628 5846 40680 1 FreeSans 480 0 0 0 en1_b
port 62 n signal bidirectional
flabel metal1 0 40137 34 40171 1 FreeSans 480 0 0 0 in_1
port 63 n signal bidirectional
flabel metal2 5794 41915 5846 41967 1 FreeSans 480 0 0 0 en0_b
port 64 n signal bidirectional
flabel metal1 0 41424 34 41458 1 FreeSans 480 0 0 0 in_0
port 65 n signal bidirectional
flabel metal2 1792 42206 1852 42260 1 FreeSans 480 0 0 0 en_b
port 66 n signal bidirectional
flabel metal2 1930 42206 1986 42260 1 FreeSans 480 0 0 0 en
port 67 n signal bidirectional
flabel metal2 1610 42114 1722 42188 1 FreeSans 480 0 0 0 VGND
port 68 n ground bidirectional
flabel metal2 2058 42114 2186 42188 1 FreeSans 480 0 0 0 VPWR
port 69 n power bidirectional
<< end >>
