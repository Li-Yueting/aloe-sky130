magic
tech sky130A
magscale 1 2
timestamp 1654309566
<< pwell >>
rect -636 -252 638 190
<< nmos >>
rect -446 -52 -416 52
rect -350 -52 -320 52
rect -254 -52 -224 52
rect -158 -52 -128 52
rect -62 -52 -32 52
rect 34 -52 64 52
rect 130 -52 160 52
rect 226 -52 256 52
rect 322 -52 352 52
rect 418 -52 448 52
<< ndiff >>
rect -508 17 -446 52
rect -508 -17 -496 17
rect -462 -17 -446 17
rect -508 -52 -446 -17
rect -416 17 -350 52
rect -416 -17 -400 17
rect -366 -17 -350 17
rect -416 -52 -350 -17
rect -320 17 -254 52
rect -320 -17 -304 17
rect -270 -17 -254 17
rect -320 -52 -254 -17
rect -224 17 -158 52
rect -224 -17 -208 17
rect -174 -17 -158 17
rect -224 -52 -158 -17
rect -128 17 -62 52
rect -128 -17 -112 17
rect -78 -17 -62 17
rect -128 -52 -62 -17
rect -32 17 34 52
rect -32 -17 -16 17
rect 18 -17 34 17
rect -32 -52 34 -17
rect 64 17 130 52
rect 64 -17 80 17
rect 114 -17 130 17
rect 64 -52 130 -17
rect 160 17 226 52
rect 160 -17 176 17
rect 210 -17 226 17
rect 160 -52 226 -17
rect 256 17 322 52
rect 256 -17 272 17
rect 306 -17 322 17
rect 256 -52 322 -17
rect 352 17 418 52
rect 352 -17 368 17
rect 402 -17 418 17
rect 352 -52 418 -17
rect 448 17 510 52
rect 448 -17 464 17
rect 498 -17 510 17
rect 448 -52 510 -17
<< ndiffc >>
rect -496 -17 -462 17
rect -400 -17 -366 17
rect -304 -17 -270 17
rect -208 -17 -174 17
rect -112 -17 -78 17
rect -16 -17 18 17
rect 80 -17 114 17
rect 176 -17 210 17
rect 272 -17 306 17
rect 368 -17 402 17
rect 464 -17 498 17
<< psubdiff >>
rect -610 130 -492 164
rect -458 130 -424 164
rect -390 130 -356 164
rect -322 130 -288 164
rect -254 130 -220 164
rect -186 130 -152 164
rect -118 130 -84 164
rect -50 130 -16 164
rect 18 130 52 164
rect 86 130 120 164
rect 154 130 188 164
rect 222 130 256 164
rect 290 130 324 164
rect 358 130 392 164
rect 426 130 460 164
rect 494 130 612 164
rect -610 54 -576 130
rect 578 54 612 130
rect -610 -14 -576 20
rect -610 -82 -576 -48
rect 578 -14 612 20
rect -610 -192 -576 -116
rect 578 -82 612 -48
rect 578 -192 612 -116
rect -610 -226 -492 -192
rect -458 -226 -424 -192
rect -390 -226 -356 -192
rect -322 -226 -288 -192
rect -254 -226 -220 -192
rect -186 -226 -152 -192
rect -118 -226 -84 -192
rect -50 -226 -16 -192
rect 18 -226 52 -192
rect 86 -226 120 -192
rect 154 -226 188 -192
rect 222 -226 256 -192
rect 290 -226 324 -192
rect 358 -226 392 -192
rect 426 -226 460 -192
rect 494 -226 612 -192
<< psubdiffcont >>
rect -492 130 -458 164
rect -424 130 -390 164
rect -356 130 -322 164
rect -288 130 -254 164
rect -220 130 -186 164
rect -152 130 -118 164
rect -84 130 -50 164
rect -16 130 18 164
rect 52 130 86 164
rect 120 130 154 164
rect 188 130 222 164
rect 256 130 290 164
rect 324 130 358 164
rect 392 130 426 164
rect 460 130 494 164
rect -610 20 -576 54
rect -610 -48 -576 -14
rect 578 20 612 54
rect 578 -48 612 -14
rect -610 -116 -576 -82
rect 578 -116 612 -82
rect -492 -226 -458 -192
rect -424 -226 -390 -192
rect -356 -226 -322 -192
rect -288 -226 -254 -192
rect -220 -226 -186 -192
rect -152 -226 -118 -192
rect -84 -226 -50 -192
rect -16 -226 18 -192
rect 52 -226 86 -192
rect 120 -226 154 -192
rect 188 -226 222 -192
rect 256 -226 290 -192
rect 324 -226 358 -192
rect 392 -226 426 -192
rect 460 -226 494 -192
<< poly >>
rect -446 52 -416 78
rect -350 52 -320 78
rect -254 52 -224 78
rect -158 52 -128 78
rect -62 52 -32 78
rect 34 52 64 78
rect 130 52 160 78
rect 226 52 256 78
rect 322 52 352 78
rect 418 52 448 78
rect -446 -74 -416 -52
rect -350 -74 -320 -52
rect -254 -74 -224 -52
rect -158 -74 -128 -52
rect -62 -74 -32 -52
rect 34 -74 64 -52
rect 130 -74 160 -52
rect 226 -74 256 -52
rect 322 -74 352 -52
rect 418 -74 448 -52
rect -512 -94 514 -74
rect -512 -128 -496 -94
rect -462 -128 -304 -94
rect -270 -128 -112 -94
rect -78 -128 80 -94
rect 114 -128 272 -94
rect 306 -128 464 -94
rect 498 -128 514 -94
rect -512 -140 514 -128
<< polycont >>
rect -496 -128 -462 -94
rect -304 -128 -270 -94
rect -112 -128 -78 -94
rect 80 -128 114 -94
rect 272 -128 306 -94
rect 464 -128 498 -94
<< locali >>
rect -610 130 -492 164
rect -458 130 -424 164
rect -390 130 -356 164
rect -322 130 -288 164
rect -254 130 -220 164
rect -186 130 -152 164
rect -118 130 -84 164
rect -50 130 -16 164
rect 18 130 52 164
rect 86 130 120 164
rect 154 130 188 164
rect 222 130 256 164
rect 290 130 324 164
rect 358 130 392 164
rect 426 130 460 164
rect 494 130 612 164
rect -610 54 -576 130
rect -610 -14 -576 20
rect -610 -82 -576 -48
rect -496 17 -462 56
rect -496 -56 -462 -17
rect -400 17 -366 56
rect -400 -56 -366 -17
rect -304 17 -270 56
rect -304 -56 -270 -17
rect -208 17 -174 56
rect -208 -56 -174 -17
rect -112 17 -78 56
rect -112 -56 -78 -17
rect -16 17 18 56
rect -16 -56 18 -17
rect 80 17 114 56
rect 80 -56 114 -17
rect 176 17 210 56
rect 176 -56 210 -17
rect 272 17 306 56
rect 272 -56 306 -17
rect 368 17 402 56
rect 368 -56 402 -17
rect 464 17 498 56
rect 464 -56 498 -17
rect 578 54 612 130
rect 578 -14 612 20
rect 578 -82 612 -48
rect -610 -192 -576 -116
rect -512 -128 -496 -94
rect -462 -128 -446 -94
rect -320 -128 -304 -94
rect -270 -128 -254 -94
rect -128 -128 -112 -94
rect -78 -128 -62 -94
rect 64 -128 80 -94
rect 114 -128 130 -94
rect 256 -128 272 -94
rect 306 -128 322 -94
rect 448 -128 464 -94
rect 498 -128 514 -94
rect 578 -192 612 -116
rect -610 -226 -492 -192
rect -458 -226 -424 -192
rect -390 -226 -356 -192
rect -322 -226 -288 -192
rect -254 -226 -220 -192
rect -186 -226 -152 -192
rect -118 -226 -84 -192
rect -50 -226 -16 -192
rect 18 -226 52 -192
rect 86 -226 120 -192
rect 154 -226 188 -192
rect 222 -226 256 -192
rect 290 -226 324 -192
rect 358 -226 392 -192
rect 426 -226 460 -192
rect 494 -226 612 -192
<< viali >>
rect -496 -17 -462 17
rect -400 -17 -366 17
rect -304 -17 -270 17
rect -208 -17 -174 17
rect -112 -17 -78 17
rect -16 -17 18 17
rect 80 -17 114 17
rect 176 -17 210 17
rect 272 -17 306 17
rect 368 -17 402 17
rect 464 -17 498 17
rect -496 -128 -462 -94
rect -304 -128 -270 -94
rect -112 -128 -78 -94
rect 80 -128 114 -94
rect 272 -128 306 -94
rect 464 -128 498 -94
<< metal1 >>
rect -502 17 -456 52
rect -502 -17 -496 17
rect -462 -17 -456 17
rect -502 -52 -456 -17
rect -406 17 -360 52
rect -406 -17 -400 17
rect -366 -17 -360 17
rect -406 -52 -360 -17
rect -310 17 -264 52
rect -310 -17 -304 17
rect -270 -17 -264 17
rect -310 -52 -264 -17
rect -214 17 -168 52
rect -214 -17 -208 17
rect -174 -17 -168 17
rect -214 -52 -168 -17
rect -118 17 -72 52
rect -118 -17 -112 17
rect -78 -17 -72 17
rect -118 -52 -72 -17
rect -22 17 24 52
rect -22 -17 -16 17
rect 18 -17 24 17
rect -22 -52 24 -17
rect 74 17 120 52
rect 74 -17 80 17
rect 114 -17 120 17
rect 74 -52 120 -17
rect 170 17 216 52
rect 170 -17 176 17
rect 210 -17 216 17
rect 170 -52 216 -17
rect 266 17 312 52
rect 266 -17 272 17
rect 306 -17 312 17
rect 266 -52 312 -17
rect 362 17 408 52
rect 362 -17 368 17
rect 402 -17 408 17
rect 362 -52 408 -17
rect 458 17 504 52
rect 458 -17 464 17
rect 498 -17 504 17
rect 458 -52 504 -17
rect -512 -94 -446 -80
rect -512 -128 -496 -94
rect -462 -128 -446 -94
rect -512 -140 -446 -128
rect -320 -94 -254 -80
rect -320 -128 -304 -94
rect -270 -128 -254 -94
rect -320 -140 -254 -128
rect -128 -94 -62 -80
rect -128 -128 -112 -94
rect -78 -128 -62 -94
rect -128 -140 -62 -128
rect 64 -94 130 -80
rect 64 -128 80 -94
rect 114 -128 130 -94
rect 64 -140 130 -128
rect 256 -94 322 -80
rect 256 -128 272 -94
rect 306 -128 322 -94
rect 256 -140 322 -128
rect 448 -94 514 -80
rect 448 -128 464 -94
rect 498 -128 514 -94
rect 448 -140 514 -128
<< properties >>
string FIXED_BBOX -594 -210 594 210
<< end >>
