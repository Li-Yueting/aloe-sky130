magic
tech sky130A
magscale 1 2
timestamp 1654747315
<< nwell >>
rect -2742 562 2644 940
rect -2742 -562 2645 562
<< pmoslvt >>
rect -2551 -500 -2351 500
rect -2293 -500 -2093 500
rect -2035 -500 -1835 500
rect -1777 -500 -1577 500
rect -1519 -500 -1319 500
rect -1261 -500 -1061 500
rect -1003 -500 -803 500
rect -745 -500 -545 500
rect -487 -500 -287 500
rect -229 -500 -29 500
rect 29 -500 229 500
rect 287 -500 487 500
rect 545 -500 745 500
rect 803 -500 1003 500
rect 1061 -500 1261 500
rect 1319 -500 1519 500
rect 1577 -500 1777 500
rect 1835 -500 2035 500
rect 2093 -500 2293 500
rect 2351 -500 2551 500
<< pdiff >>
rect -2609 488 -2551 500
rect -2609 -488 -2597 488
rect -2563 -488 -2551 488
rect -2609 -500 -2551 -488
rect -2351 488 -2293 500
rect -2351 -488 -2339 488
rect -2305 -488 -2293 488
rect -2351 -500 -2293 -488
rect -2093 488 -2035 500
rect -2093 -488 -2081 488
rect -2047 -488 -2035 488
rect -2093 -500 -2035 -488
rect -1835 488 -1777 500
rect -1835 -488 -1823 488
rect -1789 -488 -1777 488
rect -1835 -500 -1777 -488
rect -1577 488 -1519 500
rect -1577 -488 -1565 488
rect -1531 -488 -1519 488
rect -1577 -500 -1519 -488
rect -1319 488 -1261 500
rect -1319 -488 -1307 488
rect -1273 -488 -1261 488
rect -1319 -500 -1261 -488
rect -1061 488 -1003 500
rect -1061 -488 -1049 488
rect -1015 -488 -1003 488
rect -1061 -500 -1003 -488
rect -803 488 -745 500
rect -803 -488 -791 488
rect -757 -488 -745 488
rect -803 -500 -745 -488
rect -545 488 -487 500
rect -545 -488 -533 488
rect -499 -488 -487 488
rect -545 -500 -487 -488
rect -287 488 -229 500
rect -287 -488 -275 488
rect -241 -488 -229 488
rect -287 -500 -229 -488
rect -29 488 29 500
rect -29 -488 -17 488
rect 17 -488 29 488
rect -29 -500 29 -488
rect 229 488 287 500
rect 229 -488 241 488
rect 275 -488 287 488
rect 229 -500 287 -488
rect 487 488 545 500
rect 487 -488 499 488
rect 533 -488 545 488
rect 487 -500 545 -488
rect 745 488 803 500
rect 745 -488 757 488
rect 791 -488 803 488
rect 745 -500 803 -488
rect 1003 488 1061 500
rect 1003 -488 1015 488
rect 1049 -488 1061 488
rect 1003 -500 1061 -488
rect 1261 488 1319 500
rect 1261 -488 1273 488
rect 1307 -488 1319 488
rect 1261 -500 1319 -488
rect 1519 488 1577 500
rect 1519 -488 1531 488
rect 1565 -488 1577 488
rect 1519 -500 1577 -488
rect 1777 488 1835 500
rect 1777 -488 1789 488
rect 1823 -488 1835 488
rect 1777 -500 1835 -488
rect 2035 488 2093 500
rect 2035 -488 2047 488
rect 2081 -488 2093 488
rect 2035 -500 2093 -488
rect 2293 488 2351 500
rect 2293 -488 2305 488
rect 2339 -488 2351 488
rect 2293 -500 2351 -488
rect 2551 488 2609 500
rect 2551 -488 2563 488
rect 2597 -488 2609 488
rect 2551 -500 2609 -488
<< pdiffc >>
rect -2597 -488 -2563 488
rect -2339 -488 -2305 488
rect -2081 -488 -2047 488
rect -1823 -488 -1789 488
rect -1565 -488 -1531 488
rect -1307 -488 -1273 488
rect -1049 -488 -1015 488
rect -791 -488 -757 488
rect -533 -488 -499 488
rect -275 -488 -241 488
rect -17 -488 17 488
rect 241 -488 275 488
rect 499 -488 533 488
rect 757 -488 791 488
rect 1015 -488 1049 488
rect 1273 -488 1307 488
rect 1531 -488 1565 488
rect 1789 -488 1823 488
rect 2047 -488 2081 488
rect 2305 -488 2339 488
rect 2563 -488 2597 488
<< nsubdiff >>
rect -1646 808 -1526 810
rect -2704 760 -2664 800
rect -1646 772 -1606 808
rect -1562 772 -1526 808
rect -1646 770 -1526 772
rect -346 808 -226 810
rect -346 772 -306 808
rect -262 772 -226 808
rect -346 770 -226 772
rect 954 808 1074 810
rect 954 772 994 808
rect 1038 772 1074 808
rect 954 770 1074 772
rect -2704 680 -2664 720
<< nsubdiffcont >>
rect -1606 772 -1562 808
rect -306 772 -262 808
rect 994 772 1038 808
rect -2704 720 -2664 760
<< poly >>
rect -2551 500 -2351 526
rect -2293 500 -2093 526
rect -2035 500 -1835 526
rect -1777 500 -1577 526
rect -1519 500 -1319 526
rect -1261 500 -1061 526
rect -1003 500 -803 526
rect -745 500 -545 526
rect -487 500 -287 526
rect -229 500 -29 526
rect 29 500 229 526
rect 287 500 487 526
rect 545 500 745 526
rect 803 500 1003 526
rect 1061 500 1261 526
rect 1319 500 1519 526
rect 1577 500 1777 526
rect 1835 500 2035 526
rect 2093 500 2293 526
rect 2351 500 2551 526
rect -2551 -526 -2351 -500
rect -2293 -526 -2093 -500
rect -2035 -526 -1835 -500
rect -1777 -526 -1577 -500
rect -1519 -526 -1319 -500
rect -1261 -526 -1061 -500
rect -1003 -526 -803 -500
rect -745 -526 -545 -500
rect -487 -526 -287 -500
rect -229 -526 -29 -500
rect 29 -526 229 -500
rect 287 -526 487 -500
rect 545 -526 745 -500
rect 803 -526 1003 -500
rect 1061 -526 1261 -500
rect 1319 -526 1519 -500
rect 1577 -526 1777 -500
rect 1835 -526 2035 -500
rect 2093 -526 2293 -500
rect 2351 -526 2551 -500
rect -2518 -672 -2398 -526
rect -2259 -672 -2139 -526
rect -2000 -672 -1880 -526
rect -1741 -672 -1621 -526
rect -1482 -672 -1362 -526
rect -1223 -672 -1103 -526
rect -964 -672 -844 -526
rect -705 -672 -585 -526
rect -446 -672 -326 -526
rect -187 -672 -67 -526
rect 72 -672 192 -526
rect 331 -672 451 -526
rect 590 -672 710 -526
rect 849 -672 969 -526
rect 1108 -672 1228 -526
rect 1367 -672 1487 -526
rect 1626 -672 1746 -526
rect 1885 -672 2005 -526
rect 2144 -672 2264 -526
rect 2403 -672 2523 -526
rect -2644 -692 2644 -672
rect -2644 -752 -2474 -692
rect -2414 -752 -2274 -692
rect -2214 -752 -2074 -692
rect -2014 -752 -1874 -692
rect -1814 -752 -1674 -692
rect -1614 -752 -1474 -692
rect -1414 -752 -1274 -692
rect -1214 -752 -1074 -692
rect -1014 -752 -874 -692
rect -814 -752 -674 -692
rect -614 -752 -474 -692
rect -414 -752 -274 -692
rect -214 -752 -74 -692
rect -14 -752 126 -692
rect 186 -752 326 -692
rect 386 -752 526 -692
rect 586 -752 726 -692
rect 786 -752 926 -692
rect 986 -752 1126 -692
rect 1186 -752 1326 -692
rect 1386 -752 1526 -692
rect 1586 -752 1726 -692
rect 1786 -752 1926 -692
rect 1986 -752 2126 -692
rect 2186 -752 2326 -692
rect 2386 -752 2526 -692
rect 2586 -752 2644 -692
rect -2644 -772 2644 -752
<< polycont >>
rect -2474 -752 -2414 -692
rect -2274 -752 -2214 -692
rect -2074 -752 -2014 -692
rect -1874 -752 -1814 -692
rect -1674 -752 -1614 -692
rect -1474 -752 -1414 -692
rect -1274 -752 -1214 -692
rect -1074 -752 -1014 -692
rect -874 -752 -814 -692
rect -674 -752 -614 -692
rect -474 -752 -414 -692
rect -274 -752 -214 -692
rect -74 -752 -14 -692
rect 126 -752 186 -692
rect 326 -752 386 -692
rect 526 -752 586 -692
rect 726 -752 786 -692
rect 926 -752 986 -692
rect 1126 -752 1186 -692
rect 1326 -752 1386 -692
rect 1526 -752 1586 -692
rect 1726 -752 1786 -692
rect 1926 -752 1986 -692
rect 2126 -752 2186 -692
rect 2326 -752 2386 -692
rect 2526 -752 2586 -692
<< locali >>
rect -2742 850 -2474 910
rect -2414 850 -2274 910
rect -2214 850 -2074 910
rect -2014 850 -1874 910
rect -1814 850 -1674 910
rect -1614 850 -1474 910
rect -1414 850 -1274 910
rect -1214 850 -1074 910
rect -1014 850 -874 910
rect -814 850 -674 910
rect -614 850 -474 910
rect -414 850 -274 910
rect -214 850 -74 910
rect -14 850 126 910
rect 186 850 326 910
rect 386 850 526 910
rect 586 850 726 910
rect 786 850 926 910
rect 986 850 1126 910
rect 1186 850 1326 910
rect 1386 850 1526 910
rect 1586 850 1726 910
rect 1786 850 1926 910
rect 1986 850 2126 910
rect 2186 850 2326 910
rect 2386 850 2526 910
rect 2586 850 2644 910
rect -2714 760 -2654 850
rect -1666 808 -1506 850
rect -1666 772 -1606 808
rect -1562 772 -1506 808
rect -1666 770 -1506 772
rect -366 808 -206 850
rect -366 772 -306 808
rect -262 772 -206 808
rect -366 770 -206 772
rect 934 808 1094 850
rect 934 772 994 808
rect 1038 772 1094 808
rect 934 770 1094 772
rect -2714 720 -2704 760
rect -2664 720 -2654 760
rect -2714 640 -2654 720
rect -2584 690 2644 730
rect -2597 488 -2563 504
rect -2597 -692 -2563 -488
rect -2339 488 -2305 690
rect -2339 -504 -2305 -488
rect -2081 488 -2047 504
rect -2081 -692 -2047 -488
rect -1823 488 -1789 690
rect -1823 -504 -1789 -488
rect -1565 488 -1531 504
rect -1565 -692 -1531 -488
rect -1307 488 -1273 690
rect -1307 -504 -1273 -488
rect -1049 488 -1015 504
rect -1049 -692 -1015 -488
rect -791 488 -757 690
rect -791 -504 -757 -488
rect -533 488 -499 504
rect -533 -692 -499 -488
rect -275 488 -241 690
rect -275 -504 -241 -488
rect -17 488 17 504
rect -17 -692 17 -488
rect 241 488 275 690
rect 241 -504 275 -488
rect 499 488 533 504
rect 499 -692 533 -488
rect 757 488 791 690
rect 757 -504 791 -488
rect 1015 488 1049 504
rect 1015 -692 1049 -488
rect 1273 488 1307 690
rect 1273 -504 1307 -488
rect 1531 488 1565 504
rect 1531 -692 1565 -488
rect 1789 488 1823 690
rect 1789 -504 1823 -488
rect 2047 488 2081 504
rect 2047 -692 2081 -488
rect 2305 488 2339 690
rect 2305 -504 2339 -488
rect 2563 488 2597 504
rect 2563 -692 2597 -488
rect -2644 -752 -2474 -692
rect -2414 -752 -2274 -692
rect -2214 -752 -2074 -692
rect -2014 -752 -1874 -692
rect -1814 -752 -1674 -692
rect -1614 -752 -1474 -692
rect -1414 -752 -1274 -692
rect -1214 -752 -1074 -692
rect -1014 -752 -874 -692
rect -814 -752 -674 -692
rect -614 -752 -474 -692
rect -414 -752 -274 -692
rect -214 -752 -74 -692
rect -14 -752 126 -692
rect 186 -752 326 -692
rect 386 -752 526 -692
rect 586 -752 726 -692
rect 786 -752 926 -692
rect 986 -752 1126 -692
rect 1186 -752 1326 -692
rect 1386 -752 1526 -692
rect 1586 -752 1726 -692
rect 1786 -752 1926 -692
rect 1986 -752 2126 -692
rect 2186 -752 2326 -692
rect 2386 -752 2526 -692
rect 2586 -752 2644 -692
rect -2644 -790 2644 -752
rect -2742 -1030 -2474 -970
rect -2414 -1030 -2274 -970
rect -2214 -1030 -2074 -970
rect -2014 -1030 -1874 -970
rect -1814 -1030 -1674 -970
rect -1614 -1030 -1474 -970
rect -1414 -1030 -1274 -970
rect -1214 -1030 -1074 -970
rect -1014 -1030 -874 -970
rect -814 -1030 -674 -970
rect -614 -1030 -474 -970
rect -414 -1030 -274 -970
rect -214 -1030 -74 -970
rect -14 -1030 126 -970
rect 186 -1030 326 -970
rect 386 -1030 526 -970
rect 586 -1030 726 -970
rect 786 -1030 926 -970
rect 986 -1030 1126 -970
rect 1186 -1030 1326 -970
rect 1386 -1030 1526 -970
rect 1586 -1030 1726 -970
rect 1786 -1030 1926 -970
rect 1986 -1030 2126 -970
rect 2186 -1030 2326 -970
rect 2386 -1030 2526 -970
rect 2586 -1030 2644 -970
<< viali >>
rect -2474 850 -2414 910
rect -2274 850 -2214 910
rect -2074 850 -2014 910
rect -1874 850 -1814 910
rect -1674 850 -1614 910
rect -1474 850 -1414 910
rect -1274 850 -1214 910
rect -1074 850 -1014 910
rect -874 850 -814 910
rect -674 850 -614 910
rect -474 850 -414 910
rect -274 850 -214 910
rect -74 850 -14 910
rect 126 850 186 910
rect 326 850 386 910
rect 526 850 586 910
rect 726 850 786 910
rect 926 850 986 910
rect 1126 850 1186 910
rect 1326 850 1386 910
rect 1526 850 1586 910
rect 1726 850 1786 910
rect 1926 850 1986 910
rect 2126 850 2186 910
rect 2326 850 2386 910
rect 2526 850 2586 910
rect -2597 -488 -2563 488
rect -2339 -488 -2305 488
rect -2081 -488 -2047 488
rect -1823 -488 -1789 488
rect -1565 -488 -1531 488
rect -1307 -488 -1273 488
rect -1049 -488 -1015 488
rect -791 -488 -757 488
rect -533 -488 -499 488
rect -275 -488 -241 488
rect -17 -488 17 488
rect 241 -488 275 488
rect 499 -488 533 488
rect 757 -488 791 488
rect 1015 -488 1049 488
rect 1273 -488 1307 488
rect 1531 -488 1565 488
rect 1789 -488 1823 488
rect 2047 -488 2081 488
rect 2305 -488 2339 488
rect 2563 -488 2597 488
rect -2474 -1030 -2414 -970
rect -2274 -1030 -2214 -970
rect -2074 -1030 -2014 -970
rect -1874 -1030 -1814 -970
rect -1674 -1030 -1614 -970
rect -1474 -1030 -1414 -970
rect -1274 -1030 -1214 -970
rect -1074 -1030 -1014 -970
rect -874 -1030 -814 -970
rect -674 -1030 -614 -970
rect -474 -1030 -414 -970
rect -274 -1030 -214 -970
rect -74 -1030 -14 -970
rect 126 -1030 186 -970
rect 326 -1030 386 -970
rect 526 -1030 586 -970
rect 726 -1030 786 -970
rect 926 -1030 986 -970
rect 1126 -1030 1186 -970
rect 1326 -1030 1386 -970
rect 1526 -1030 1586 -970
rect 1726 -1030 1786 -970
rect 1926 -1030 1986 -970
rect 2126 -1030 2186 -970
rect 2326 -1030 2386 -970
rect 2526 -1030 2586 -970
<< metal1 >>
rect -2742 910 2644 940
rect -2742 850 -2474 910
rect -2414 850 -2274 910
rect -2214 850 -2074 910
rect -2014 850 -1874 910
rect -1814 850 -1674 910
rect -1614 850 -1474 910
rect -1414 850 -1274 910
rect -1214 850 -1074 910
rect -1014 850 -874 910
rect -814 850 -674 910
rect -614 850 -474 910
rect -414 850 -274 910
rect -214 850 -74 910
rect -14 850 126 910
rect 186 850 326 910
rect 386 850 526 910
rect 586 850 726 910
rect 786 850 926 910
rect 986 850 1126 910
rect 1186 850 1326 910
rect 1386 850 1526 910
rect 1586 850 1726 910
rect 1786 850 1926 910
rect 1986 850 2126 910
rect 2186 850 2326 910
rect 2386 850 2526 910
rect 2586 850 2644 910
rect -2742 820 2644 850
rect -2603 488 -2557 500
rect -2603 -488 -2597 488
rect -2563 -488 -2557 488
rect -2603 -500 -2557 -488
rect -2345 488 -2299 500
rect -2345 -488 -2339 488
rect -2305 -488 -2299 488
rect -2345 -500 -2299 -488
rect -2087 488 -2041 500
rect -2087 -488 -2081 488
rect -2047 -488 -2041 488
rect -2087 -500 -2041 -488
rect -1829 488 -1783 500
rect -1829 -488 -1823 488
rect -1789 -488 -1783 488
rect -1829 -500 -1783 -488
rect -1571 488 -1525 500
rect -1571 -488 -1565 488
rect -1531 -488 -1525 488
rect -1571 -500 -1525 -488
rect -1313 488 -1267 500
rect -1313 -488 -1307 488
rect -1273 -488 -1267 488
rect -1313 -500 -1267 -488
rect -1055 488 -1009 500
rect -1055 -488 -1049 488
rect -1015 -488 -1009 488
rect -1055 -500 -1009 -488
rect -797 488 -751 500
rect -797 -488 -791 488
rect -757 -488 -751 488
rect -797 -500 -751 -488
rect -539 488 -493 500
rect -539 -488 -533 488
rect -499 -488 -493 488
rect -539 -500 -493 -488
rect -281 488 -235 500
rect -281 -488 -275 488
rect -241 -488 -235 488
rect -281 -500 -235 -488
rect -23 488 23 500
rect -23 -488 -17 488
rect 17 -488 23 488
rect -23 -500 23 -488
rect 235 488 281 500
rect 235 -488 241 488
rect 275 -488 281 488
rect 235 -500 281 -488
rect 493 488 539 500
rect 493 -488 499 488
rect 533 -488 539 488
rect 493 -500 539 -488
rect 751 488 797 500
rect 751 -488 757 488
rect 791 -488 797 488
rect 751 -500 797 -488
rect 1009 488 1055 500
rect 1009 -488 1015 488
rect 1049 -488 1055 488
rect 1009 -500 1055 -488
rect 1267 488 1313 500
rect 1267 -488 1273 488
rect 1307 -488 1313 488
rect 1267 -500 1313 -488
rect 1525 488 1571 500
rect 1525 -488 1531 488
rect 1565 -488 1571 488
rect 1525 -500 1571 -488
rect 1783 488 1829 500
rect 1783 -488 1789 488
rect 1823 -488 1829 488
rect 1783 -500 1829 -488
rect 2041 488 2087 500
rect 2041 -488 2047 488
rect 2081 -488 2087 488
rect 2041 -500 2087 -488
rect 2299 488 2345 500
rect 2299 -488 2305 488
rect 2339 -488 2345 488
rect 2299 -500 2345 -488
rect 2557 488 2603 500
rect 2557 -488 2563 488
rect 2597 -488 2603 488
rect 2557 -500 2603 -488
rect -2742 -970 2644 -940
rect -2742 -1030 -2474 -970
rect -2414 -1030 -2274 -970
rect -2214 -1030 -2074 -970
rect -2014 -1030 -1874 -970
rect -1814 -1030 -1674 -970
rect -1614 -1030 -1474 -970
rect -1414 -1030 -1274 -970
rect -1214 -1030 -1074 -970
rect -1014 -1030 -874 -970
rect -814 -1030 -674 -970
rect -614 -1030 -474 -970
rect -414 -1030 -274 -970
rect -214 -1030 -74 -970
rect -14 -1030 126 -970
rect 186 -1030 326 -970
rect 386 -1030 526 -970
rect 586 -1030 726 -970
rect 786 -1030 926 -970
rect 986 -1030 1126 -970
rect 1186 -1030 1326 -970
rect 1386 -1030 1526 -970
rect 1586 -1030 1726 -970
rect 1786 -1030 1926 -970
rect 1986 -1030 2126 -970
rect 2186 -1030 2326 -970
rect 2386 -1030 2526 -970
rect 2586 -1030 2644 -970
rect -2742 -1060 2644 -1030
<< labels >>
flabel nwell -2742 850 -2682 910 1 FreeSans 800 0 0 0 VPWR
flabel metal1 -2742 -1030 -2584 -970 1 FreeSans 800 0 0 0 VGND
flabel locali 2584 690 2644 730 1 FreeSans 800 0 0 0 SOURCE
flabel locali 2584 -790 2644 -730 1 FreeSans 800 0 0 0 DRAIN
flabel locali 2584 -752 2644 -692 1 FreeSans 800 0 0 0 GATE
<< end >>
