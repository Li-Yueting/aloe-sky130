VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO decoder5x32
  CLASS BLOCK ;
  FOREIGN decoder5x32 ;
  ORIGIN 0.000 0.000 ;
  SIZE 41.400 BY 36.040 ;
  PIN a[4]
    ANTENNAGATEAREA 0.373500 ;
    PORT
      LAYER li1 ;
        RECT 16.120 11.135 16.455 11.185 ;
        RECT 18.030 11.135 18.380 11.175 ;
        RECT 16.120 10.965 18.380 11.135 ;
        RECT 16.120 10.935 16.455 10.965 ;
        RECT 18.030 10.935 18.380 10.965 ;
      LAYER mcon ;
        RECT 18.085 10.965 18.255 11.135 ;
      LAYER met1 ;
        RECT 18.010 11.120 18.330 11.180 ;
        RECT 17.735 10.980 18.330 11.120 ;
        RECT 18.010 10.920 18.330 10.980 ;
      LAYER via ;
        RECT 18.040 10.920 18.300 11.180 ;
      LAYER met2 ;
        RECT 18.040 10.890 18.300 11.210 ;
        RECT 18.100 1.065 18.240 10.890 ;
        RECT 18.030 0.695 18.310 1.065 ;
      LAYER via2 ;
        RECT 18.030 0.740 18.310 1.020 ;
      LAYER met3 ;
        RECT 18.005 1.030 18.335 1.045 ;
        RECT 0.000 0.730 18.335 1.030 ;
        RECT 18.005 0.715 18.335 0.730 ;
    END
  END a[4]
  PIN a[3]
    ANTENNAGATEAREA 0.810000 ;
    PORT
      LAYER li1 ;
        RECT 15.265 13.975 15.615 14.225 ;
        RECT 17.565 13.975 17.805 14.925 ;
        RECT 18.945 13.975 19.295 14.225 ;
      LAYER mcon ;
        RECT 15.325 14.025 15.495 14.195 ;
        RECT 17.625 14.025 17.795 14.195 ;
        RECT 19.005 14.025 19.175 14.195 ;
      LAYER met1 ;
        RECT 15.265 13.995 15.555 14.225 ;
        RECT 17.090 14.180 17.410 14.240 ;
        RECT 17.565 14.180 17.855 14.225 ;
        RECT 18.945 14.180 19.235 14.225 ;
        RECT 16.720 14.040 19.235 14.180 ;
        RECT 15.340 13.840 15.480 13.995 ;
        RECT 16.720 13.840 16.860 14.040 ;
        RECT 17.090 13.980 17.410 14.040 ;
        RECT 17.565 13.995 17.855 14.040 ;
        RECT 18.945 13.995 19.235 14.040 ;
        RECT 15.340 13.700 16.860 13.840 ;
      LAYER via ;
        RECT 17.120 13.980 17.380 14.240 ;
      LAYER met2 ;
        RECT 17.120 13.950 17.380 14.270 ;
        RECT 17.180 11.120 17.320 13.950 ;
        RECT 16.720 10.980 17.320 11.120 ;
        RECT 16.720 3.640 16.860 10.980 ;
        RECT 16.720 3.500 17.320 3.640 ;
        RECT 17.180 2.895 17.320 3.500 ;
        RECT 17.110 2.525 17.390 2.895 ;
      LAYER via2 ;
        RECT 17.110 2.570 17.390 2.850 ;
      LAYER met3 ;
        RECT 17.085 2.860 17.415 2.875 ;
        RECT 0.000 2.560 17.415 2.860 ;
        RECT 17.085 2.545 17.415 2.560 ;
    END
  END a[3]
  PIN a[2]
    ANTENNAGATEAREA 4.950000 ;
    PORT
      LAYER li1 ;
        RECT 14.325 25.075 14.610 25.185 ;
        RECT 14.830 25.075 15.050 25.435 ;
        RECT 14.325 24.905 15.050 25.075 ;
        RECT 14.325 24.855 14.610 24.905 ;
        RECT 14.830 24.855 15.050 24.905 ;
        RECT 26.285 24.855 26.570 25.185 ;
        RECT 27.740 24.855 28.115 25.415 ;
        RECT 16.240 21.505 16.615 22.065 ;
        RECT 25.435 21.735 25.815 22.065 ;
        RECT 25.435 21.040 25.650 21.735 ;
        RECT 29.090 21.485 29.310 22.065 ;
        RECT 18.510 19.745 18.725 20.440 ;
        RECT 18.345 19.415 18.725 19.745 ;
        RECT 21.660 19.415 22.025 19.675 ;
        RECT 13.450 16.045 13.670 16.625 ;
        RECT 16.155 16.365 16.520 16.625 ;
        RECT 24.420 16.365 24.785 16.625 ;
        RECT 27.665 16.295 27.950 16.625 ;
        RECT 28.660 16.065 29.035 16.625 ;
        RECT 11.175 14.305 11.390 15.000 ;
        RECT 11.175 13.975 11.555 14.305 ;
        RECT 14.205 13.975 14.580 14.535 ;
        RECT 25.410 14.305 25.625 15.000 ;
        RECT 21.200 13.975 21.565 14.235 ;
        RECT 25.245 13.975 25.625 14.305 ;
        RECT 10.690 10.855 10.975 11.185 ;
        RECT 25.430 10.605 25.650 11.185 ;
      LAYER mcon ;
        RECT 14.405 24.905 14.575 25.075 ;
        RECT 26.365 24.905 26.535 25.075 ;
        RECT 27.745 24.905 27.915 25.075 ;
        RECT 16.245 21.845 16.415 22.015 ;
        RECT 29.125 21.845 29.295 22.015 ;
        RECT 25.445 21.505 25.615 21.675 ;
        RECT 18.545 19.465 18.715 19.635 ;
        RECT 21.765 19.465 21.935 19.635 ;
        RECT 16.245 16.405 16.415 16.575 ;
        RECT 24.525 16.405 24.695 16.575 ;
        RECT 27.745 16.405 27.915 16.575 ;
        RECT 28.665 16.405 28.835 16.575 ;
        RECT 13.485 16.065 13.655 16.235 ;
        RECT 14.405 14.365 14.575 14.535 ;
        RECT 11.185 14.025 11.355 14.195 ;
        RECT 25.445 14.365 25.615 14.535 ;
        RECT 21.305 14.025 21.475 14.195 ;
        RECT 10.725 10.965 10.895 11.135 ;
        RECT 25.445 10.965 25.615 11.135 ;
      LAYER met1 ;
        RECT 14.330 25.060 14.650 25.120 ;
        RECT 14.055 24.920 14.650 25.060 ;
        RECT 14.330 24.860 14.650 24.920 ;
        RECT 26.305 25.060 26.595 25.105 ;
        RECT 27.685 25.060 27.975 25.105 ;
        RECT 26.305 24.920 27.975 25.060 ;
        RECT 26.305 24.875 26.595 24.920 ;
        RECT 27.685 24.875 27.975 24.920 ;
        RECT 27.760 24.720 27.900 24.875 ;
        RECT 29.050 24.720 29.370 24.780 ;
        RECT 27.760 24.580 29.370 24.720 ;
        RECT 29.050 24.520 29.370 24.580 ;
        RECT 14.790 22.680 15.110 22.740 ;
        RECT 14.790 22.540 15.940 22.680 ;
        RECT 14.790 22.480 15.110 22.540 ;
        RECT 15.800 22.000 15.940 22.540 ;
        RECT 16.185 22.000 16.475 22.045 ;
        RECT 18.010 22.000 18.330 22.060 ;
        RECT 29.050 22.000 29.370 22.060 ;
        RECT 15.800 21.860 18.330 22.000 ;
        RECT 28.775 21.860 29.370 22.000 ;
        RECT 16.185 21.815 16.475 21.860 ;
        RECT 18.010 21.800 18.330 21.860 ;
        RECT 29.050 21.800 29.370 21.860 ;
        RECT 25.370 21.660 25.690 21.720 ;
        RECT 25.095 21.520 25.690 21.660 ;
        RECT 25.370 21.460 25.690 21.520 ;
        RECT 18.010 19.620 18.330 19.680 ;
        RECT 18.485 19.620 18.775 19.665 ;
        RECT 21.690 19.620 22.010 19.680 ;
        RECT 18.010 19.480 18.775 19.620 ;
        RECT 21.415 19.480 22.010 19.620 ;
        RECT 18.010 19.420 18.330 19.480 ;
        RECT 18.485 19.435 18.775 19.480 ;
        RECT 21.690 19.420 22.010 19.480 ;
        RECT 18.010 16.900 18.330 16.960 ;
        RECT 21.230 16.900 21.550 16.960 ;
        RECT 13.500 16.760 21.550 16.900 ;
        RECT 10.650 16.220 10.970 16.280 ;
        RECT 13.500 16.265 13.640 16.760 ;
        RECT 16.260 16.605 16.400 16.760 ;
        RECT 18.010 16.700 18.330 16.760 ;
        RECT 21.230 16.700 21.550 16.760 ;
        RECT 16.185 16.560 16.475 16.605 ;
        RECT 16.630 16.560 16.950 16.620 ;
        RECT 24.450 16.560 24.770 16.620 ;
        RECT 27.670 16.560 27.990 16.620 ;
        RECT 16.185 16.420 16.950 16.560 ;
        RECT 16.185 16.375 16.475 16.420 ;
        RECT 16.630 16.360 16.950 16.420 ;
        RECT 24.080 16.420 24.770 16.560 ;
        RECT 27.395 16.420 27.990 16.560 ;
        RECT 13.425 16.220 13.715 16.265 ;
        RECT 10.650 16.080 13.715 16.220 ;
        RECT 10.650 16.020 10.970 16.080 ;
        RECT 13.425 16.035 13.715 16.080 ;
        RECT 21.230 16.220 21.550 16.280 ;
        RECT 24.080 16.220 24.220 16.420 ;
        RECT 24.450 16.360 24.770 16.420 ;
        RECT 27.670 16.360 27.990 16.420 ;
        RECT 28.590 16.560 28.910 16.620 ;
        RECT 28.590 16.420 29.185 16.560 ;
        RECT 28.590 16.360 28.910 16.420 ;
        RECT 21.230 16.080 24.220 16.220 ;
        RECT 21.230 16.020 21.550 16.080 ;
        RECT 14.345 14.520 14.635 14.565 ;
        RECT 16.630 14.520 16.950 14.580 ;
        RECT 23.070 14.520 23.390 14.580 ;
        RECT 25.385 14.520 25.675 14.565 ;
        RECT 14.345 14.380 16.950 14.520 ;
        RECT 14.345 14.335 14.635 14.380 ;
        RECT 16.630 14.320 16.950 14.380 ;
        RECT 21.780 14.380 25.675 14.520 ;
        RECT 10.650 14.180 10.970 14.240 ;
        RECT 11.125 14.180 11.415 14.225 ;
        RECT 10.650 14.040 11.415 14.180 ;
        RECT 10.650 13.980 10.970 14.040 ;
        RECT 11.125 13.995 11.415 14.040 ;
        RECT 21.230 14.180 21.550 14.240 ;
        RECT 21.780 14.180 21.920 14.380 ;
        RECT 23.070 14.320 23.390 14.380 ;
        RECT 25.385 14.335 25.675 14.380 ;
        RECT 21.230 14.040 21.920 14.180 ;
        RECT 21.230 13.980 21.550 14.040 ;
        RECT 23.530 11.800 23.850 11.860 ;
        RECT 23.530 11.660 25.600 11.800 ;
        RECT 23.530 11.600 23.850 11.660 ;
        RECT 4.210 11.120 4.530 11.180 ;
        RECT 10.650 11.120 10.970 11.180 ;
        RECT 25.460 11.165 25.600 11.660 ;
        RECT 4.210 10.980 10.970 11.120 ;
        RECT 4.210 10.920 4.530 10.980 ;
        RECT 10.650 10.920 10.970 10.980 ;
        RECT 25.385 10.935 25.675 11.165 ;
      LAYER via ;
        RECT 14.360 24.860 14.620 25.120 ;
        RECT 29.080 24.520 29.340 24.780 ;
        RECT 14.820 22.480 15.080 22.740 ;
        RECT 18.040 21.800 18.300 22.060 ;
        RECT 29.080 21.800 29.340 22.060 ;
        RECT 25.400 21.460 25.660 21.720 ;
        RECT 18.040 19.420 18.300 19.680 ;
        RECT 21.720 19.420 21.980 19.680 ;
        RECT 10.680 16.020 10.940 16.280 ;
        RECT 18.040 16.700 18.300 16.960 ;
        RECT 21.260 16.700 21.520 16.960 ;
        RECT 16.660 16.360 16.920 16.620 ;
        RECT 21.260 16.020 21.520 16.280 ;
        RECT 24.480 16.360 24.740 16.620 ;
        RECT 27.700 16.360 27.960 16.620 ;
        RECT 28.620 16.360 28.880 16.620 ;
        RECT 16.660 14.320 16.920 14.580 ;
        RECT 10.680 13.980 10.940 14.240 ;
        RECT 21.260 13.980 21.520 14.240 ;
        RECT 23.100 14.320 23.360 14.580 ;
        RECT 23.560 11.600 23.820 11.860 ;
        RECT 4.240 10.920 4.500 11.180 ;
        RECT 10.680 10.920 10.940 11.180 ;
      LAYER met2 ;
        RECT 14.360 24.830 14.620 25.150 ;
        RECT 14.420 22.680 14.560 24.830 ;
        RECT 29.080 24.490 29.340 24.810 ;
        RECT 29.140 23.025 29.280 24.490 ;
        RECT 14.820 22.680 15.080 22.770 ;
        RECT 14.420 22.540 15.080 22.680 ;
        RECT 29.070 22.655 29.350 23.025 ;
        RECT 14.820 22.450 15.080 22.540 ;
        RECT 29.140 22.090 29.280 22.655 ;
        RECT 18.040 21.770 18.300 22.090 ;
        RECT 29.080 21.770 29.340 22.090 ;
        RECT 18.100 19.975 18.240 21.770 ;
        RECT 25.400 21.430 25.660 21.750 ;
        RECT 25.460 21.195 25.600 21.430 ;
        RECT 25.390 20.825 25.670 21.195 ;
        RECT 18.030 19.605 18.310 19.975 ;
        RECT 21.710 19.605 21.990 19.975 ;
        RECT 18.040 19.390 18.300 19.605 ;
        RECT 21.720 19.390 21.980 19.605 ;
        RECT 18.100 16.990 18.240 19.390 ;
        RECT 18.040 16.670 18.300 16.990 ;
        RECT 21.260 16.670 21.520 16.990 ;
        RECT 16.660 16.330 16.920 16.650 ;
        RECT 10.680 15.990 10.940 16.310 ;
        RECT 10.740 14.270 10.880 15.990 ;
        RECT 16.720 14.610 16.860 16.330 ;
        RECT 21.320 16.310 21.460 16.670 ;
        RECT 24.470 16.555 24.750 16.925 ;
        RECT 27.690 16.560 27.970 16.925 ;
        RECT 28.620 16.560 28.880 16.650 ;
        RECT 27.690 16.555 28.880 16.560 ;
        RECT 24.480 16.330 24.740 16.555 ;
        RECT 27.700 16.420 28.880 16.555 ;
        RECT 27.700 16.330 27.960 16.420 ;
        RECT 28.620 16.330 28.880 16.420 ;
        RECT 21.260 15.990 21.520 16.310 ;
        RECT 16.660 14.290 16.920 14.610 ;
        RECT 21.320 14.270 21.460 15.990 ;
        RECT 23.100 14.290 23.360 14.610 ;
        RECT 10.680 13.950 10.940 14.270 ;
        RECT 21.260 13.950 21.520 14.270 ;
        RECT 10.740 11.210 10.880 13.950 ;
        RECT 23.160 13.840 23.300 14.290 ;
        RECT 23.160 13.700 23.760 13.840 ;
        RECT 23.620 11.890 23.760 13.700 ;
        RECT 23.560 11.570 23.820 11.890 ;
        RECT 4.240 10.890 4.500 11.210 ;
        RECT 10.680 10.890 10.940 11.210 ;
        RECT 4.300 4.725 4.440 10.890 ;
        RECT 4.230 4.355 4.510 4.725 ;
      LAYER via2 ;
        RECT 29.070 22.700 29.350 22.980 ;
        RECT 25.390 20.870 25.670 21.150 ;
        RECT 18.030 19.650 18.310 19.930 ;
        RECT 21.710 19.650 21.990 19.930 ;
        RECT 24.470 16.600 24.750 16.880 ;
        RECT 27.690 16.600 27.970 16.880 ;
        RECT 4.230 4.400 4.510 4.680 ;
      LAYER met3 ;
        RECT 29.045 22.990 29.375 23.005 ;
        RECT 24.000 22.690 29.375 22.990 ;
        RECT 24.000 21.160 24.300 22.690 ;
        RECT 29.045 22.675 29.375 22.690 ;
        RECT 25.365 21.160 25.695 21.175 ;
        RECT 24.000 20.860 25.695 21.160 ;
        RECT 18.005 19.940 18.335 19.955 ;
        RECT 21.685 19.940 22.015 19.955 ;
        RECT 24.000 19.940 24.300 20.860 ;
        RECT 25.365 20.845 25.695 20.860 ;
        RECT 18.005 19.640 24.300 19.940 ;
        RECT 18.005 19.625 18.335 19.640 ;
        RECT 21.685 19.625 22.015 19.640 ;
        RECT 24.445 16.890 24.775 16.905 ;
        RECT 27.665 16.890 27.995 16.905 ;
        RECT 24.445 16.590 27.995 16.890 ;
        RECT 24.445 16.575 24.775 16.590 ;
        RECT 27.665 16.575 27.995 16.590 ;
        RECT 4.205 4.690 4.535 4.705 ;
        RECT 0.000 4.390 4.535 4.690 ;
        RECT 4.205 4.375 4.535 4.390 ;
    END
  END a[2]
  PIN a[1]
    ANTENNAGATEAREA 4.230000 ;
    PORT
      LAYER li1 ;
        RECT 10.665 24.855 10.975 25.185 ;
        RECT 12.505 24.515 12.745 25.185 ;
        RECT 19.805 24.855 20.155 25.105 ;
        RECT 24.465 24.515 24.705 25.185 ;
        RECT 27.225 21.735 27.535 22.065 ;
        RECT 11.175 19.415 11.415 20.365 ;
        RECT 12.945 19.415 13.255 19.745 ;
        RECT 15.205 19.415 15.555 19.665 ;
        RECT 19.405 19.415 19.645 20.365 ;
        RECT 23.085 19.415 23.325 20.365 ;
        RECT 26.765 19.415 27.115 19.665 ;
        RECT 25.845 16.295 26.085 16.965 ;
        RECT 22.625 13.975 22.865 14.925 ;
        RECT 12.555 10.855 12.795 11.525 ;
        RECT 20.325 10.935 20.675 11.185 ;
        RECT 27.685 10.855 27.995 11.185 ;
      LAYER mcon ;
        RECT 10.725 24.905 10.895 25.075 ;
        RECT 19.925 24.905 20.095 25.075 ;
        RECT 24.525 24.905 24.695 25.075 ;
        RECT 12.565 24.565 12.735 24.735 ;
        RECT 27.285 21.845 27.455 22.015 ;
        RECT 11.185 20.145 11.355 20.315 ;
        RECT 19.465 19.805 19.635 19.975 ;
        RECT 13.025 19.465 13.195 19.635 ;
        RECT 15.325 19.465 15.495 19.635 ;
        RECT 23.145 19.465 23.315 19.635 ;
        RECT 26.825 19.465 26.995 19.635 ;
        RECT 25.905 16.405 26.075 16.575 ;
        RECT 22.685 14.025 22.855 14.195 ;
        RECT 12.565 10.965 12.735 11.135 ;
        RECT 20.385 10.965 20.555 11.135 ;
        RECT 27.745 10.965 27.915 11.135 ;
      LAYER met1 ;
        RECT 10.665 24.875 10.955 25.105 ;
        RECT 19.850 25.060 20.170 25.120 ;
        RECT 24.465 25.060 24.755 25.105 ;
        RECT 19.850 24.920 24.755 25.060 ;
        RECT 9.730 24.720 10.050 24.780 ;
        RECT 10.740 24.720 10.880 24.875 ;
        RECT 19.850 24.860 20.170 24.920 ;
        RECT 24.465 24.875 24.755 24.920 ;
        RECT 12.505 24.720 12.795 24.765 ;
        RECT 9.730 24.580 12.795 24.720 ;
        RECT 9.730 24.520 10.050 24.580 ;
        RECT 12.505 24.535 12.795 24.580 ;
        RECT 27.210 22.000 27.530 22.060 ;
        RECT 27.210 21.860 27.805 22.000 ;
        RECT 27.210 21.800 27.530 21.860 ;
        RECT 9.730 20.300 10.050 20.360 ;
        RECT 11.125 20.300 11.415 20.345 ;
        RECT 27.210 20.300 27.530 20.360 ;
        RECT 9.730 20.160 11.415 20.300 ;
        RECT 9.730 20.100 10.050 20.160 ;
        RECT 10.280 19.280 10.420 20.160 ;
        RECT 11.125 20.115 11.415 20.160 ;
        RECT 25.000 20.160 27.530 20.300 ;
        RECT 19.390 19.960 19.710 20.020 ;
        RECT 19.115 19.820 19.710 19.960 ;
        RECT 19.390 19.760 19.710 19.820 ;
        RECT 12.965 19.620 13.255 19.665 ;
        RECT 15.265 19.620 15.555 19.665 ;
        RECT 23.085 19.620 23.375 19.665 ;
        RECT 25.000 19.620 25.140 20.160 ;
        RECT 26.840 19.665 26.980 20.160 ;
        RECT 27.210 20.100 27.530 20.160 ;
        RECT 12.965 19.480 17.320 19.620 ;
        RECT 12.965 19.435 13.255 19.480 ;
        RECT 15.265 19.435 15.555 19.480 ;
        RECT 13.040 19.280 13.180 19.435 ;
        RECT 10.280 19.140 13.180 19.280 ;
        RECT 17.180 19.280 17.320 19.480 ;
        RECT 22.240 19.480 25.140 19.620 ;
        RECT 19.390 19.280 19.710 19.340 ;
        RECT 22.240 19.280 22.380 19.480 ;
        RECT 23.085 19.435 23.375 19.480 ;
        RECT 26.765 19.435 27.055 19.665 ;
        RECT 17.180 19.140 22.380 19.280 ;
        RECT 19.390 19.080 19.710 19.140 ;
        RECT 22.240 19.000 22.380 19.140 ;
        RECT 22.150 18.740 22.470 19.000 ;
        RECT 22.150 16.900 22.470 16.960 ;
        RECT 22.150 16.760 25.140 16.900 ;
        RECT 22.150 16.700 22.470 16.760 ;
        RECT 25.000 16.560 25.140 16.760 ;
        RECT 25.845 16.560 26.135 16.605 ;
        RECT 25.000 16.420 26.135 16.560 ;
        RECT 25.845 16.375 26.135 16.420 ;
        RECT 22.625 13.995 22.915 14.225 ;
        RECT 20.770 13.840 21.090 13.900 ;
        RECT 22.150 13.840 22.470 13.900 ;
        RECT 22.700 13.840 22.840 13.995 ;
        RECT 20.770 13.700 22.840 13.840 ;
        RECT 20.770 13.640 21.090 13.700 ;
        RECT 22.150 13.640 22.470 13.700 ;
        RECT 27.670 11.940 27.990 12.200 ;
        RECT 13.960 11.490 18.700 11.630 ;
        RECT 13.960 11.460 14.100 11.490 ;
        RECT 13.040 11.320 14.100 11.460 ;
        RECT 18.560 11.460 18.700 11.490 ;
        RECT 20.770 11.460 21.090 11.520 ;
        RECT 18.560 11.320 21.090 11.460 ;
        RECT 12.030 11.120 12.350 11.180 ;
        RECT 12.505 11.120 12.795 11.165 ;
        RECT 13.040 11.120 13.180 11.320 ;
        RECT 12.030 10.980 13.180 11.120 ;
        RECT 19.480 11.120 19.620 11.320 ;
        RECT 20.770 11.260 21.090 11.320 ;
        RECT 27.760 11.165 27.900 11.940 ;
        RECT 20.325 11.120 20.615 11.165 ;
        RECT 19.480 10.980 20.615 11.120 ;
        RECT 12.030 10.920 12.350 10.980 ;
        RECT 12.505 10.935 12.795 10.980 ;
        RECT 20.325 10.935 20.615 10.980 ;
        RECT 27.685 10.935 27.975 11.165 ;
      LAYER via ;
        RECT 9.760 24.520 10.020 24.780 ;
        RECT 19.880 24.860 20.140 25.120 ;
        RECT 27.240 21.800 27.500 22.060 ;
        RECT 9.760 20.100 10.020 20.360 ;
        RECT 19.420 19.760 19.680 20.020 ;
        RECT 27.240 20.100 27.500 20.360 ;
        RECT 19.420 19.080 19.680 19.340 ;
        RECT 22.180 18.740 22.440 19.000 ;
        RECT 22.180 16.700 22.440 16.960 ;
        RECT 20.800 13.640 21.060 13.900 ;
        RECT 22.180 13.640 22.440 13.900 ;
        RECT 27.700 11.940 27.960 12.200 ;
        RECT 12.060 10.920 12.320 11.180 ;
        RECT 20.800 11.260 21.060 11.520 ;
      LAYER met2 ;
        RECT 19.880 24.830 20.140 25.150 ;
        RECT 9.760 24.490 10.020 24.810 ;
        RECT 9.820 20.390 9.960 24.490 ;
        RECT 19.940 24.040 20.080 24.830 ;
        RECT 19.020 23.900 20.080 24.040 ;
        RECT 19.020 20.980 19.160 23.900 ;
        RECT 27.240 21.770 27.500 22.090 ;
        RECT 19.020 20.840 19.620 20.980 ;
        RECT 9.760 20.070 10.020 20.390 ;
        RECT 19.480 20.050 19.620 20.840 ;
        RECT 27.300 20.390 27.440 21.770 ;
        RECT 27.240 20.070 27.500 20.390 ;
        RECT 19.420 19.730 19.680 20.050 ;
        RECT 19.480 19.370 19.620 19.730 ;
        RECT 19.420 19.050 19.680 19.370 ;
        RECT 22.180 18.710 22.440 19.030 ;
        RECT 22.240 16.990 22.380 18.710 ;
        RECT 22.180 16.670 22.440 16.990 ;
        RECT 22.240 15.095 22.380 16.670 ;
        RECT 22.170 14.725 22.450 15.095 ;
        RECT 27.690 14.725 27.970 15.095 ;
        RECT 22.240 13.930 22.380 14.725 ;
        RECT 20.800 13.610 21.060 13.930 ;
        RECT 22.180 13.610 22.440 13.930 ;
        RECT 20.860 11.520 21.000 13.610 ;
        RECT 27.760 12.230 27.900 14.725 ;
        RECT 27.700 11.910 27.960 12.230 ;
        RECT 20.770 11.260 21.090 11.520 ;
        RECT 12.060 10.890 12.320 11.210 ;
        RECT 12.120 6.555 12.260 10.890 ;
        RECT 12.050 6.185 12.330 6.555 ;
      LAYER via2 ;
        RECT 22.170 14.770 22.450 15.050 ;
        RECT 27.690 14.770 27.970 15.050 ;
        RECT 12.050 6.230 12.330 6.510 ;
      LAYER met3 ;
        RECT 22.145 15.060 22.475 15.075 ;
        RECT 27.665 15.060 27.995 15.075 ;
        RECT 22.145 14.760 27.995 15.060 ;
        RECT 22.145 14.745 22.475 14.760 ;
        RECT 27.665 14.745 27.995 14.760 ;
        RECT 12.025 6.520 12.355 6.535 ;
        RECT 0.000 6.220 12.355 6.520 ;
        RECT 12.025 6.205 12.355 6.220 ;
    END
  END a[1]
  PIN a[0]
    ANTENNAGATEAREA 5.940000 ;
    PORT
      LAYER li1 ;
        RECT 11.180 24.855 11.555 25.415 ;
        RECT 13.370 25.355 13.720 25.880 ;
        RECT 25.330 25.355 25.680 25.880 ;
        RECT 13.370 25.185 13.575 25.355 ;
        RECT 25.330 25.185 25.535 25.355 ;
        RECT 13.265 24.855 13.575 25.185 ;
        RECT 18.945 24.855 19.295 25.105 ;
        RECT 25.225 24.855 25.535 25.185 ;
        RECT 12.025 21.735 12.335 22.065 ;
        RECT 18.085 22.015 18.255 23.035 ;
        RECT 18.485 22.015 18.835 22.065 ;
        RECT 18.085 21.845 18.835 22.015 ;
        RECT 18.485 21.815 18.835 21.845 ;
        RECT 21.225 21.735 21.535 22.065 ;
        RECT 23.545 21.815 23.895 22.065 ;
        RECT 26.815 21.735 27.055 22.405 ;
        RECT 27.740 21.505 28.115 22.065 ;
        RECT 12.365 19.415 12.740 19.975 ;
        RECT 13.945 19.635 14.115 19.975 ;
        RECT 14.345 19.635 14.695 19.665 ;
        RECT 13.945 19.465 14.695 19.635 ;
        RECT 16.245 19.635 16.415 19.975 ;
        RECT 17.105 19.635 17.345 19.745 ;
        RECT 16.245 19.465 17.345 19.635 ;
        RECT 14.345 19.415 14.695 19.465 ;
        RECT 17.105 19.075 17.345 19.465 ;
        RECT 26.285 19.415 26.595 19.745 ;
        RECT 27.625 19.415 27.975 19.665 ;
        RECT 12.905 16.375 13.255 16.625 ;
        RECT 26.605 16.295 26.915 16.625 ;
        RECT 26.710 16.125 26.915 16.295 ;
        RECT 26.710 15.600 27.060 16.125 ;
        RECT 12.555 13.635 12.795 14.305 ;
        RECT 24.005 13.635 24.245 14.305 ;
        RECT 26.765 14.195 27.115 14.225 ;
        RECT 26.365 14.025 27.115 14.195 ;
        RECT 26.365 13.345 26.535 14.025 ;
        RECT 26.765 13.975 27.115 14.025 ;
        RECT 11.725 10.855 12.035 11.185 ;
        RECT 21.185 10.935 21.535 11.185 ;
        RECT 25.845 10.855 26.155 11.185 ;
        RECT 11.725 10.685 11.930 10.855 ;
        RECT 11.580 10.160 11.930 10.685 ;
        RECT 28.200 10.625 28.575 11.185 ;
      LAYER mcon ;
        RECT 13.485 25.585 13.655 25.755 ;
        RECT 25.445 25.585 25.615 25.755 ;
        RECT 11.185 24.905 11.355 25.075 ;
        RECT 19.005 24.905 19.175 25.075 ;
        RECT 18.085 22.865 18.255 23.035 ;
        RECT 12.105 21.845 12.275 22.015 ;
        RECT 26.825 22.185 26.995 22.355 ;
        RECT 21.305 21.845 21.475 22.015 ;
        RECT 23.605 21.845 23.775 22.015 ;
        RECT 27.745 21.505 27.915 21.675 ;
        RECT 12.565 19.465 12.735 19.635 ;
        RECT 13.945 19.805 14.115 19.975 ;
        RECT 16.245 19.805 16.415 19.975 ;
        RECT 26.365 19.465 26.535 19.635 ;
        RECT 27.745 19.465 27.915 19.635 ;
        RECT 13.025 16.405 13.195 16.575 ;
        RECT 26.825 15.725 26.995 15.895 ;
        RECT 12.565 13.685 12.735 13.855 ;
        RECT 24.065 13.685 24.235 13.855 ;
        RECT 21.305 10.965 21.475 11.135 ;
        RECT 25.905 10.965 26.075 11.135 ;
        RECT 28.205 10.965 28.375 11.135 ;
        RECT 11.645 10.285 11.815 10.455 ;
      LAYER met1 ;
        RECT 13.425 25.740 13.715 25.785 ;
        RECT 13.040 25.600 13.715 25.740 ;
        RECT 13.040 25.400 13.180 25.600 ;
        RECT 13.425 25.555 13.715 25.600 ;
        RECT 23.990 25.740 24.310 25.800 ;
        RECT 25.385 25.740 25.675 25.785 ;
        RECT 23.990 25.600 25.675 25.740 ;
        RECT 23.990 25.540 24.310 25.600 ;
        RECT 25.385 25.555 25.675 25.600 ;
        RECT 11.200 25.260 16.400 25.400 ;
        RECT 11.200 25.120 11.340 25.260 ;
        RECT 11.110 25.060 11.430 25.120 ;
        RECT 16.260 25.060 16.400 25.260 ;
        RECT 18.010 25.060 18.330 25.120 ;
        RECT 18.945 25.060 19.235 25.105 ;
        RECT 11.110 24.920 11.705 25.060 ;
        RECT 16.260 24.920 19.235 25.060 ;
        RECT 11.110 24.860 11.430 24.920 ;
        RECT 18.010 24.860 18.330 24.920 ;
        RECT 18.945 24.875 19.235 24.920 ;
        RECT 18.010 23.020 18.330 23.080 ;
        RECT 20.310 23.020 20.630 23.080 ;
        RECT 17.735 22.880 20.630 23.020 ;
        RECT 18.010 22.820 18.330 22.880 ;
        RECT 20.310 22.820 20.630 22.880 ;
        RECT 23.990 22.340 24.310 22.400 ;
        RECT 26.765 22.340 27.055 22.385 ;
        RECT 23.620 22.200 27.055 22.340 ;
        RECT 11.110 22.000 11.430 22.060 ;
        RECT 12.045 22.000 12.335 22.045 ;
        RECT 11.110 21.860 12.335 22.000 ;
        RECT 11.110 21.800 11.430 21.860 ;
        RECT 12.045 21.815 12.335 21.860 ;
        RECT 20.310 22.000 20.630 22.060 ;
        RECT 23.620 22.045 23.760 22.200 ;
        RECT 23.990 22.140 24.310 22.200 ;
        RECT 26.765 22.155 27.055 22.200 ;
        RECT 21.245 22.000 21.535 22.045 ;
        RECT 23.545 22.000 23.835 22.045 ;
        RECT 20.310 21.860 21.535 22.000 ;
        RECT 20.310 21.800 20.630 21.860 ;
        RECT 21.245 21.815 21.535 21.860 ;
        RECT 23.160 21.860 23.835 22.000 ;
        RECT 20.400 21.320 20.540 21.800 ;
        RECT 23.160 21.320 23.300 21.860 ;
        RECT 23.545 21.815 23.835 21.860 ;
        RECT 26.840 21.660 26.980 22.155 ;
        RECT 27.670 21.660 27.990 21.720 ;
        RECT 26.840 21.520 27.990 21.660 ;
        RECT 27.670 21.460 27.990 21.520 ;
        RECT 20.400 21.180 23.300 21.320 ;
        RECT 13.410 19.960 13.730 20.020 ;
        RECT 13.885 19.960 14.175 20.005 ;
        RECT 16.185 19.960 16.475 20.005 ;
        RECT 12.580 19.820 16.475 19.960 ;
        RECT 10.650 19.620 10.970 19.680 ;
        RECT 12.580 19.665 12.720 19.820 ;
        RECT 13.410 19.760 13.730 19.820 ;
        RECT 13.885 19.775 14.175 19.820 ;
        RECT 16.185 19.775 16.475 19.820 ;
        RECT 12.505 19.620 12.795 19.665 ;
        RECT 10.650 19.480 12.795 19.620 ;
        RECT 10.650 19.420 10.970 19.480 ;
        RECT 12.505 19.435 12.795 19.480 ;
        RECT 26.305 19.435 26.595 19.665 ;
        RECT 27.670 19.620 27.990 19.680 ;
        RECT 27.300 19.480 27.990 19.620 ;
        RECT 26.380 19.280 26.520 19.435 ;
        RECT 27.300 19.280 27.440 19.480 ;
        RECT 27.670 19.420 27.990 19.480 ;
        RECT 26.380 19.140 27.440 19.280 ;
        RECT 12.950 16.560 13.270 16.620 ;
        RECT 12.675 16.420 13.270 16.560 ;
        RECT 12.950 16.360 13.270 16.420 ;
        RECT 25.830 15.880 26.150 15.940 ;
        RECT 26.765 15.880 27.055 15.925 ;
        RECT 25.830 15.740 27.055 15.880 ;
        RECT 25.830 15.680 26.150 15.740 ;
        RECT 26.765 15.695 27.055 15.740 ;
        RECT 12.490 13.840 12.810 13.900 ;
        RECT 12.215 13.700 12.810 13.840 ;
        RECT 12.490 13.640 12.810 13.700 ;
        RECT 24.005 13.655 24.295 13.885 ;
        RECT 24.080 13.500 24.220 13.655 ;
        RECT 25.830 13.500 26.150 13.560 ;
        RECT 26.305 13.500 26.595 13.545 ;
        RECT 24.080 13.360 26.595 13.500 ;
        RECT 25.830 13.300 26.150 13.360 ;
        RECT 26.305 13.315 26.595 13.360 ;
        RECT 21.230 11.120 21.550 11.180 ;
        RECT 20.955 10.980 21.550 11.120 ;
        RECT 21.230 10.920 21.550 10.980 ;
        RECT 25.830 11.120 26.150 11.180 ;
        RECT 28.130 11.120 28.450 11.180 ;
        RECT 25.830 10.980 26.425 11.120 ;
        RECT 28.130 10.980 28.725 11.120 ;
        RECT 25.830 10.920 26.150 10.980 ;
        RECT 28.130 10.920 28.450 10.980 ;
        RECT 1.450 10.440 1.770 10.500 ;
        RECT 2.460 10.470 10.880 10.610 ;
        RECT 2.460 10.440 2.600 10.470 ;
        RECT 1.450 10.300 2.600 10.440 ;
        RECT 10.740 10.440 10.880 10.470 ;
        RECT 11.585 10.440 11.875 10.485 ;
        RECT 12.490 10.440 12.810 10.500 ;
        RECT 20.310 10.440 20.630 10.500 ;
        RECT 10.740 10.300 20.630 10.440 ;
        RECT 1.450 10.240 1.770 10.300 ;
        RECT 11.585 10.255 11.875 10.300 ;
        RECT 12.490 10.240 12.810 10.300 ;
        RECT 20.310 10.240 20.630 10.300 ;
      LAYER via ;
        RECT 24.020 25.540 24.280 25.800 ;
        RECT 11.140 24.860 11.400 25.120 ;
        RECT 18.040 24.860 18.300 25.120 ;
        RECT 18.040 22.820 18.300 23.080 ;
        RECT 20.340 22.820 20.600 23.080 ;
        RECT 11.140 21.800 11.400 22.060 ;
        RECT 20.340 21.800 20.600 22.060 ;
        RECT 24.020 22.140 24.280 22.400 ;
        RECT 27.700 21.460 27.960 21.720 ;
        RECT 10.680 19.420 10.940 19.680 ;
        RECT 13.440 19.760 13.700 20.020 ;
        RECT 27.700 19.420 27.960 19.680 ;
        RECT 12.980 16.360 13.240 16.620 ;
        RECT 25.860 15.680 26.120 15.940 ;
        RECT 12.520 13.640 12.780 13.900 ;
        RECT 25.860 13.300 26.120 13.560 ;
        RECT 21.260 10.920 21.520 11.180 ;
        RECT 25.860 10.920 26.120 11.180 ;
        RECT 28.160 10.920 28.420 11.180 ;
        RECT 1.480 10.240 1.740 10.500 ;
        RECT 12.520 10.240 12.780 10.500 ;
        RECT 20.340 10.240 20.600 10.500 ;
      LAYER met2 ;
        RECT 24.020 25.510 24.280 25.830 ;
        RECT 11.140 24.830 11.400 25.150 ;
        RECT 18.040 24.830 18.300 25.150 ;
        RECT 11.200 22.090 11.340 24.830 ;
        RECT 18.100 23.110 18.240 24.830 ;
        RECT 18.040 22.790 18.300 23.110 ;
        RECT 20.340 22.790 20.600 23.110 ;
        RECT 20.400 22.090 20.540 22.790 ;
        RECT 24.080 22.430 24.220 25.510 ;
        RECT 24.020 22.110 24.280 22.430 ;
        RECT 11.140 22.000 11.400 22.090 ;
        RECT 10.740 21.860 11.400 22.000 ;
        RECT 10.740 19.710 10.880 21.860 ;
        RECT 11.140 21.770 11.400 21.860 ;
        RECT 20.340 21.770 20.600 22.090 ;
        RECT 27.700 21.430 27.960 21.750 ;
        RECT 13.440 19.730 13.700 20.050 ;
        RECT 10.680 19.390 10.940 19.710 ;
        RECT 13.500 17.920 13.640 19.730 ;
        RECT 27.760 19.710 27.900 21.430 ;
        RECT 27.700 19.390 27.960 19.710 ;
        RECT 13.040 17.780 13.640 17.920 ;
        RECT 13.040 16.650 13.180 17.780 ;
        RECT 12.980 16.330 13.240 16.650 ;
        RECT 12.520 13.840 12.780 13.930 ;
        RECT 13.040 13.840 13.180 16.330 ;
        RECT 25.860 15.650 26.120 15.970 ;
        RECT 12.520 13.700 13.180 13.840 ;
        RECT 12.520 13.610 12.780 13.700 ;
        RECT 12.580 10.530 12.720 13.610 ;
        RECT 25.920 13.590 26.060 15.650 ;
        RECT 25.860 13.270 26.120 13.590 ;
        RECT 25.920 12.045 26.060 13.270 ;
        RECT 21.250 11.675 21.530 12.045 ;
        RECT 25.850 11.675 26.130 12.045 ;
        RECT 28.150 11.675 28.430 12.045 ;
        RECT 21.320 11.210 21.460 11.675 ;
        RECT 25.920 11.210 26.060 11.675 ;
        RECT 28.220 11.210 28.360 11.675 ;
        RECT 21.260 11.120 21.520 11.210 ;
        RECT 20.400 10.980 21.520 11.120 ;
        RECT 20.400 10.530 20.540 10.980 ;
        RECT 21.260 10.890 21.520 10.980 ;
        RECT 25.860 10.890 26.120 11.210 ;
        RECT 28.160 10.890 28.420 11.210 ;
        RECT 1.480 10.210 1.740 10.530 ;
        RECT 12.520 10.210 12.780 10.530 ;
        RECT 20.340 10.210 20.600 10.530 ;
        RECT 1.540 8.385 1.680 10.210 ;
        RECT 1.470 8.015 1.750 8.385 ;
      LAYER via2 ;
        RECT 21.250 11.720 21.530 12.000 ;
        RECT 25.850 11.720 26.130 12.000 ;
        RECT 28.150 11.720 28.430 12.000 ;
        RECT 1.470 8.060 1.750 8.340 ;
      LAYER met3 ;
        RECT 21.225 12.010 21.555 12.025 ;
        RECT 25.825 12.010 26.155 12.025 ;
        RECT 28.125 12.010 28.455 12.025 ;
        RECT 21.225 11.710 28.455 12.010 ;
        RECT 21.225 11.695 21.555 11.710 ;
        RECT 25.825 11.695 26.155 11.710 ;
        RECT 28.125 11.695 28.455 11.710 ;
        RECT 1.445 8.350 1.775 8.365 ;
        RECT 0.000 8.050 1.775 8.350 ;
        RECT 1.445 8.035 1.775 8.050 ;
    END
  END a[0]
  PIN en
    ANTENNAGATEAREA 0.495000 ;
    PORT
      LAYER li1 ;
        RECT 15.275 11.135 15.610 11.185 ;
        RECT 14.865 10.965 15.610 11.135 ;
        RECT 15.275 10.915 15.610 10.965 ;
        RECT 18.550 10.935 19.025 11.175 ;
      LAYER mcon ;
        RECT 18.775 10.965 18.945 11.135 ;
      LAYER met1 ;
        RECT 13.410 11.120 13.730 11.180 ;
        RECT 14.805 11.120 15.095 11.165 ;
        RECT 13.410 10.980 17.320 11.120 ;
        RECT 13.410 10.920 13.730 10.980 ;
        RECT 14.805 10.935 15.095 10.980 ;
        RECT 17.180 10.780 17.320 10.980 ;
        RECT 18.715 10.935 19.005 11.165 ;
        RECT 18.790 10.780 18.930 10.935 ;
        RECT 17.180 10.640 18.930 10.780 ;
      LAYER via ;
        RECT 13.440 10.920 13.700 11.180 ;
      LAYER met2 ;
        RECT 13.430 10.455 13.710 11.210 ;
      LAYER via2 ;
        RECT 13.430 10.500 13.710 10.780 ;
      LAYER met3 ;
        RECT 13.405 10.790 13.735 10.805 ;
        RECT 1.000 10.490 13.735 10.790 ;
        RECT 1.000 10.180 1.300 10.490 ;
        RECT 13.405 10.475 13.735 10.490 ;
        RECT 0.000 9.880 1.300 10.180 ;
    END
  END en
  PIN y[31]
    ANTENNADIFFAREA 0.795000 ;
    PORT
      LAYER li1 ;
        RECT 11.095 11.525 11.425 12.325 ;
        RECT 11.965 11.525 12.295 12.325 ;
        RECT 11.095 11.355 12.375 11.525 ;
        RECT 12.205 10.685 12.375 11.355 ;
        RECT 12.100 10.115 12.795 10.685 ;
      LAYER mcon ;
        RECT 11.185 11.985 11.355 12.155 ;
      LAYER met1 ;
        RECT 0.990 12.140 1.310 12.200 ;
        RECT 11.125 12.140 11.415 12.185 ;
        RECT 0.990 12.000 5.820 12.140 ;
        RECT 0.990 11.940 1.310 12.000 ;
        RECT 5.680 11.800 5.820 12.000 ;
        RECT 10.280 12.000 11.415 12.140 ;
        RECT 10.280 11.800 10.420 12.000 ;
        RECT 11.125 11.955 11.415 12.000 ;
        RECT 5.680 11.660 10.420 11.800 ;
      LAYER via ;
        RECT 1.020 11.940 1.280 12.200 ;
      LAYER met2 ;
        RECT 1.010 11.910 1.290 12.655 ;
      LAYER via2 ;
        RECT 1.010 12.330 1.290 12.610 ;
      LAYER met3 ;
        RECT 0.985 12.620 1.315 12.635 ;
        RECT 0.000 12.320 1.315 12.620 ;
        RECT 0.985 12.305 1.315 12.320 ;
    END
  END y[31]
  PIN y[30]
    ANTENNADIFFAREA 0.699000 ;
    PORT
      LAYER li1 ;
        RECT 13.855 14.705 15.085 15.045 ;
        RECT 13.855 13.805 14.035 14.705 ;
        RECT 14.755 14.475 15.085 14.705 ;
        RECT 13.855 13.635 15.085 13.805 ;
        RECT 13.855 12.835 14.185 13.635 ;
        RECT 14.755 12.835 15.085 13.635 ;
      LAYER mcon ;
        RECT 13.945 14.705 14.115 14.875 ;
      LAYER met1 ;
        RECT 12.490 14.860 12.810 14.920 ;
        RECT 13.885 14.860 14.175 14.905 ;
        RECT 12.490 14.720 14.175 14.860 ;
        RECT 12.490 14.660 12.810 14.720 ;
        RECT 13.885 14.675 14.175 14.720 ;
      LAYER via ;
        RECT 12.520 14.660 12.780 14.920 ;
      LAYER met2 ;
        RECT 12.520 14.630 12.780 14.950 ;
        RECT 12.580 14.485 12.720 14.630 ;
        RECT 12.510 14.115 12.790 14.485 ;
      LAYER via2 ;
        RECT 12.510 14.160 12.790 14.440 ;
      LAYER met3 ;
        RECT 12.485 14.450 12.815 14.465 ;
        RECT 0.000 14.150 12.815 14.450 ;
        RECT 12.485 14.135 12.815 14.150 ;
    END
  END y[30]
  PIN y[29]
    ANTENNADIFFAREA 0.795000 ;
    PORT
      LAYER li1 ;
        RECT 12.100 14.475 12.795 15.045 ;
        RECT 12.205 13.805 12.375 14.475 ;
        RECT 11.095 13.635 12.375 13.805 ;
        RECT 11.095 12.835 11.425 13.635 ;
        RECT 11.965 12.835 12.295 13.635 ;
      LAYER mcon ;
        RECT 11.185 13.345 11.355 13.515 ;
      LAYER met1 ;
        RECT 7.060 13.700 9.960 13.840 ;
        RECT 6.050 13.500 6.370 13.560 ;
        RECT 7.060 13.500 7.200 13.700 ;
        RECT 6.050 13.360 7.200 13.500 ;
        RECT 9.820 13.500 9.960 13.700 ;
        RECT 11.125 13.500 11.415 13.545 ;
        RECT 9.820 13.360 11.415 13.500 ;
        RECT 6.050 13.300 6.370 13.360 ;
        RECT 11.125 13.315 11.415 13.360 ;
      LAYER via ;
        RECT 6.080 13.300 6.340 13.560 ;
      LAYER met2 ;
        RECT 6.070 15.945 6.350 16.315 ;
        RECT 6.140 13.590 6.280 15.945 ;
        RECT 6.080 13.270 6.340 13.590 ;
      LAYER via2 ;
        RECT 6.070 15.990 6.350 16.270 ;
      LAYER met3 ;
        RECT 6.045 16.280 6.375 16.295 ;
        RECT 0.000 15.980 6.375 16.280 ;
        RECT 6.045 15.965 6.375 15.980 ;
    END
  END y[29]
  PIN y[28]
    ANTENNADIFFAREA 0.699000 ;
    PORT
      LAYER li1 ;
        RECT 13.855 16.965 14.185 17.765 ;
        RECT 14.755 16.965 15.085 17.765 ;
        RECT 13.855 16.795 15.085 16.965 ;
        RECT 13.855 15.895 14.035 16.795 ;
        RECT 14.755 15.895 15.085 16.125 ;
        RECT 13.855 15.555 15.085 15.895 ;
      LAYER mcon ;
        RECT 13.945 17.085 14.115 17.255 ;
      LAYER met1 ;
        RECT 0.990 17.240 1.310 17.300 ;
        RECT 13.885 17.240 14.175 17.285 ;
        RECT 0.990 17.100 5.820 17.240 ;
        RECT 0.990 17.040 1.310 17.100 ;
        RECT 5.680 16.900 5.820 17.100 ;
        RECT 12.580 17.100 14.175 17.240 ;
        RECT 12.580 17.070 12.720 17.100 ;
        RECT 9.820 16.930 12.720 17.070 ;
        RECT 13.885 17.055 14.175 17.100 ;
        RECT 9.820 16.900 9.960 16.930 ;
        RECT 5.680 16.760 9.960 16.900 ;
      LAYER via ;
        RECT 1.020 17.040 1.280 17.300 ;
      LAYER met2 ;
        RECT 1.010 17.775 1.290 18.145 ;
        RECT 1.080 17.330 1.220 17.775 ;
        RECT 1.020 17.010 1.280 17.330 ;
      LAYER via2 ;
        RECT 1.010 17.820 1.290 18.100 ;
      LAYER met3 ;
        RECT 0.985 18.110 1.315 18.125 ;
        RECT 0.000 17.810 1.315 18.110 ;
        RECT 0.985 17.795 1.315 17.810 ;
    END
  END y[28]
  PIN y[27]
    ANTENNADIFFAREA 0.699000 ;
    PORT
      LAYER li1 ;
        RECT 12.015 20.145 13.245 20.485 ;
        RECT 12.015 19.245 12.195 20.145 ;
        RECT 12.915 19.915 13.245 20.145 ;
        RECT 12.015 19.075 13.245 19.245 ;
        RECT 12.015 18.275 12.345 19.075 ;
        RECT 12.915 18.275 13.245 19.075 ;
      LAYER mcon ;
        RECT 13.025 20.145 13.195 20.315 ;
      LAYER met1 ;
        RECT 12.950 20.300 13.270 20.360 ;
        RECT 12.675 20.160 13.270 20.300 ;
        RECT 12.950 20.100 13.270 20.160 ;
      LAYER via ;
        RECT 12.980 20.100 13.240 20.360 ;
      LAYER met2 ;
        RECT 12.970 19.605 13.250 20.390 ;
      LAYER via2 ;
        RECT 12.970 19.650 13.250 19.930 ;
      LAYER met3 ;
        RECT 12.945 19.940 13.275 19.955 ;
        RECT 0.000 19.640 13.275 19.940 ;
        RECT 12.945 19.625 13.275 19.640 ;
    END
  END y[27]
  PIN y[26]
    ANTENNADIFFAREA 0.439000 ;
    PORT
      LAYER li1 ;
        RECT 12.955 22.225 13.285 23.205 ;
        RECT 13.020 22.185 13.195 22.225 ;
        RECT 13.020 21.625 13.190 22.185 ;
        RECT 13.020 20.995 13.715 21.625 ;
      LAYER mcon ;
        RECT 13.025 22.185 13.195 22.355 ;
      LAYER met1 ;
        RECT 2.370 22.340 2.690 22.400 ;
        RECT 12.965 22.340 13.255 22.385 ;
        RECT 2.370 22.200 4.440 22.340 ;
        RECT 2.370 22.140 2.690 22.200 ;
        RECT 4.300 22.000 4.440 22.200 ;
        RECT 10.280 22.200 13.255 22.340 ;
        RECT 10.280 22.000 10.420 22.200 ;
        RECT 12.965 22.155 13.255 22.200 ;
        RECT 4.300 21.860 10.420 22.000 ;
      LAYER via ;
        RECT 2.400 22.140 2.660 22.400 ;
      LAYER met2 ;
        RECT 2.400 22.110 2.660 22.430 ;
        RECT 2.460 21.805 2.600 22.110 ;
        RECT 2.390 21.435 2.670 21.805 ;
      LAYER via2 ;
        RECT 2.390 21.480 2.670 21.760 ;
      LAYER met3 ;
        RECT 2.365 21.770 2.695 21.785 ;
        RECT 0.000 21.470 2.695 21.770 ;
        RECT 2.365 21.455 2.695 21.470 ;
    END
  END y[26]
  PIN y[25]
    ANTENNADIFFAREA 0.699000 ;
    PORT
      LAYER li1 ;
        RECT 11.095 22.405 11.425 23.205 ;
        RECT 11.995 22.405 12.325 23.205 ;
        RECT 11.095 22.235 12.325 22.405 ;
        RECT 11.095 21.335 11.275 22.235 ;
        RECT 11.995 21.335 12.325 21.565 ;
        RECT 11.095 20.995 12.325 21.335 ;
      LAYER mcon ;
        RECT 11.185 22.865 11.355 23.035 ;
      LAYER met1 ;
        RECT 4.670 23.020 4.990 23.080 ;
        RECT 11.125 23.020 11.415 23.065 ;
        RECT 4.670 22.880 5.820 23.020 ;
        RECT 4.670 22.820 4.990 22.880 ;
        RECT 5.680 22.680 5.820 22.880 ;
        RECT 9.360 22.880 11.415 23.020 ;
        RECT 9.360 22.680 9.500 22.880 ;
        RECT 11.125 22.835 11.415 22.880 ;
        RECT 5.680 22.540 9.500 22.680 ;
      LAYER via ;
        RECT 4.700 22.820 4.960 23.080 ;
      LAYER met2 ;
        RECT 4.690 23.875 4.970 24.245 ;
        RECT 4.760 23.110 4.900 23.875 ;
        RECT 4.700 22.790 4.960 23.110 ;
      LAYER via2 ;
        RECT 4.690 23.920 4.970 24.200 ;
      LAYER met3 ;
        RECT 4.665 24.210 4.995 24.225 ;
        RECT 0.000 23.910 4.995 24.210 ;
        RECT 4.665 23.895 4.995 23.910 ;
    END
  END y[25]
  PIN y[24]
    ANTENNADIFFAREA 0.439000 ;
    PORT
      LAYER li1 ;
        RECT 14.335 22.225 14.665 23.205 ;
        RECT 14.400 21.625 14.570 22.225 ;
        RECT 14.400 20.995 15.095 21.625 ;
      LAYER mcon ;
        RECT 14.405 22.865 14.575 23.035 ;
      LAYER met1 ;
        RECT 14.345 23.020 14.635 23.065 ;
        RECT 16.170 23.020 16.490 23.080 ;
        RECT 14.345 22.880 16.490 23.020 ;
        RECT 14.345 22.835 14.635 22.880 ;
        RECT 16.170 22.820 16.490 22.880 ;
      LAYER via ;
        RECT 16.200 22.820 16.460 23.080 ;
      LAYER met2 ;
        RECT 16.190 25.095 16.470 25.465 ;
        RECT 16.260 23.110 16.400 25.095 ;
        RECT 16.200 22.790 16.460 23.110 ;
      LAYER via2 ;
        RECT 16.190 25.140 16.470 25.420 ;
      LAYER met3 ;
        RECT 0.000 25.740 1.300 26.040 ;
        RECT 1.000 25.430 1.300 25.740 ;
        RECT 16.165 25.430 16.495 25.445 ;
        RECT 1.000 25.130 16.495 25.430 ;
        RECT 16.165 25.115 16.495 25.130 ;
    END
  END y[24]
  PIN y[23]
    ANTENNADIFFAREA 0.795000 ;
    PORT
      LAYER li1 ;
        RECT 12.505 25.355 13.200 25.925 ;
        RECT 12.925 24.685 13.095 25.355 ;
        RECT 12.925 24.515 14.205 24.685 ;
        RECT 13.005 23.715 13.335 24.515 ;
        RECT 13.875 23.715 14.205 24.515 ;
      LAYER mcon ;
        RECT 12.565 25.585 12.735 25.755 ;
      LAYER met1 ;
        RECT 12.030 25.740 12.350 25.800 ;
        RECT 12.505 25.740 12.795 25.785 ;
        RECT 12.030 25.600 12.795 25.740 ;
        RECT 12.030 25.540 12.350 25.600 ;
        RECT 12.505 25.555 12.795 25.600 ;
      LAYER via ;
        RECT 12.060 25.540 12.320 25.800 ;
      LAYER met2 ;
        RECT 12.050 26.315 12.330 26.685 ;
        RECT 12.120 25.830 12.260 26.315 ;
        RECT 12.060 25.510 12.320 25.830 ;
      LAYER via2 ;
        RECT 12.050 26.360 12.330 26.640 ;
      LAYER met3 ;
        RECT 0.000 27.570 12.340 27.870 ;
        RECT 12.040 26.665 12.340 27.570 ;
        RECT 12.025 26.335 12.355 26.665 ;
    END
  END y[23]
  PIN y[22]
    ANTENNADIFFAREA 0.699000 ;
    PORT
      LAYER li1 ;
        RECT 15.735 22.405 16.065 23.205 ;
        RECT 16.635 22.405 16.965 23.205 ;
        RECT 15.735 22.235 16.965 22.405 ;
        RECT 15.735 21.335 16.065 21.565 ;
        RECT 16.785 21.335 16.965 22.235 ;
        RECT 15.735 20.995 16.965 21.335 ;
      LAYER mcon ;
        RECT 16.705 22.865 16.875 23.035 ;
      LAYER met1 ;
        RECT 16.645 23.020 16.935 23.065 ;
        RECT 17.090 23.020 17.410 23.080 ;
        RECT 16.645 22.880 17.410 23.020 ;
        RECT 16.645 22.835 16.935 22.880 ;
        RECT 17.090 22.820 17.410 22.880 ;
      LAYER via ;
        RECT 17.120 22.820 17.380 23.080 ;
      LAYER met2 ;
        RECT 17.110 29.365 17.390 29.735 ;
        RECT 17.180 23.110 17.320 29.365 ;
        RECT 17.120 22.790 17.380 23.110 ;
      LAYER via2 ;
        RECT 17.110 29.410 17.390 29.690 ;
      LAYER met3 ;
        RECT 17.085 29.700 17.415 29.715 ;
        RECT 0.000 29.400 17.415 29.700 ;
        RECT 17.085 29.385 17.415 29.400 ;
    END
  END y[22]
  PIN y[21]
    ANTENNADIFFAREA 0.795000 ;
    PORT
      LAYER li1 ;
        RECT 17.105 19.915 17.800 20.485 ;
        RECT 17.525 19.245 17.695 19.915 ;
        RECT 17.525 19.075 18.805 19.245 ;
        RECT 17.605 18.275 17.935 19.075 ;
        RECT 18.475 18.275 18.805 19.075 ;
      LAYER mcon ;
        RECT 17.625 18.785 17.795 18.955 ;
      LAYER met1 ;
        RECT 6.600 19.140 9.500 19.280 ;
        RECT 5.590 18.940 5.910 19.000 ;
        RECT 6.600 18.940 6.740 19.140 ;
        RECT 5.590 18.800 6.740 18.940 ;
        RECT 9.360 18.940 9.500 19.140 ;
        RECT 17.565 18.940 17.855 18.985 ;
        RECT 9.360 18.800 10.420 18.940 ;
        RECT 5.590 18.740 5.910 18.800 ;
        RECT 10.280 18.770 10.420 18.800 ;
        RECT 13.500 18.800 17.855 18.940 ;
        RECT 13.500 18.770 13.640 18.800 ;
        RECT 10.280 18.630 13.640 18.770 ;
        RECT 17.565 18.755 17.855 18.800 ;
      LAYER via ;
        RECT 5.620 18.740 5.880 19.000 ;
      LAYER met2 ;
        RECT 5.610 31.195 5.890 31.565 ;
        RECT 5.680 19.030 5.820 31.195 ;
        RECT 5.620 18.710 5.880 19.030 ;
      LAYER via2 ;
        RECT 5.610 31.240 5.890 31.520 ;
      LAYER met3 ;
        RECT 5.585 31.530 5.915 31.545 ;
        RECT 0.000 31.230 5.915 31.530 ;
        RECT 5.585 31.215 5.915 31.230 ;
    END
  END y[21]
  PIN y[20]
    ANTENNADIFFAREA 0.699000 ;
    PORT
      LAYER li1 ;
        RECT 15.235 25.585 16.465 25.925 ;
        RECT 15.235 24.685 15.415 25.585 ;
        RECT 16.135 25.355 16.465 25.585 ;
        RECT 15.235 24.515 16.465 24.685 ;
        RECT 15.235 23.715 15.565 24.515 ;
        RECT 16.135 23.715 16.465 24.515 ;
      LAYER mcon ;
        RECT 15.325 25.585 15.495 25.755 ;
      LAYER met1 ;
        RECT 15.250 25.740 15.570 25.800 ;
        RECT 14.975 25.600 15.570 25.740 ;
        RECT 15.250 25.540 15.570 25.600 ;
      LAYER via ;
        RECT 15.280 25.540 15.540 25.800 ;
      LAYER met2 ;
        RECT 15.270 33.025 15.550 33.395 ;
        RECT 15.340 25.830 15.480 33.025 ;
        RECT 15.280 25.510 15.540 25.830 ;
      LAYER via2 ;
        RECT 15.270 33.070 15.550 33.350 ;
      LAYER met3 ;
        RECT 15.245 33.360 15.575 33.375 ;
        RECT 0.000 33.060 15.575 33.360 ;
        RECT 15.245 33.045 15.575 33.060 ;
    END
  END y[20]
  PIN y[19]
    ANTENNADIFFAREA 0.699000 ;
    PORT
      LAYER li1 ;
        RECT 10.675 25.585 11.905 25.925 ;
        RECT 10.675 25.355 11.005 25.585 ;
        RECT 11.725 24.685 11.905 25.585 ;
        RECT 10.675 24.515 11.905 24.685 ;
        RECT 10.675 23.715 11.005 24.515 ;
        RECT 11.575 23.715 11.905 24.515 ;
      LAYER mcon ;
        RECT 10.725 25.585 10.895 25.755 ;
      LAYER met1 ;
        RECT 10.650 25.740 10.970 25.800 ;
        RECT 10.375 25.600 10.970 25.740 ;
        RECT 10.650 25.540 10.970 25.600 ;
      LAYER via ;
        RECT 10.680 25.540 10.940 25.800 ;
      LAYER met2 ;
        RECT 10.670 34.855 10.950 35.225 ;
        RECT 10.740 25.830 10.880 34.855 ;
        RECT 10.680 25.510 10.940 25.830 ;
      LAYER via2 ;
        RECT 10.670 34.900 10.950 35.180 ;
      LAYER met3 ;
        RECT 10.645 35.190 10.975 35.205 ;
        RECT 0.000 34.890 10.975 35.190 ;
        RECT 10.645 34.875 10.975 34.890 ;
    END
  END y[19]
  PIN y[18]
    ANTENNADIFFAREA 0.439000 ;
    PORT
      LAYER li1 ;
        RECT 22.155 22.225 22.485 23.205 ;
        RECT 22.220 21.625 22.390 22.225 ;
        RECT 22.220 20.995 22.915 21.625 ;
      LAYER mcon ;
        RECT 22.225 22.865 22.395 23.035 ;
      LAYER met1 ;
        RECT 22.165 23.020 22.455 23.065 ;
        RECT 25.370 23.020 25.690 23.080 ;
        RECT 22.165 22.880 25.690 23.020 ;
        RECT 22.165 22.835 22.455 22.880 ;
        RECT 25.370 22.820 25.690 22.880 ;
      LAYER via ;
        RECT 25.400 22.820 25.660 23.080 ;
      LAYER met2 ;
        RECT 25.390 35.465 25.670 35.835 ;
        RECT 25.460 23.110 25.600 35.465 ;
        RECT 25.400 22.790 25.660 23.110 ;
      LAYER via2 ;
        RECT 25.390 35.510 25.670 35.790 ;
      LAYER met3 ;
        RECT 25.365 35.800 25.695 35.815 ;
        RECT 25.365 35.500 41.400 35.800 ;
        RECT 25.365 35.485 25.695 35.500 ;
    END
  END y[18]
  PIN y[17]
    ANTENNADIFFAREA 0.699000 ;
    PORT
      LAYER li1 ;
        RECT 20.295 22.405 20.625 23.205 ;
        RECT 21.195 22.405 21.525 23.205 ;
        RECT 20.295 22.235 21.525 22.405 ;
        RECT 20.295 21.335 20.475 22.235 ;
        RECT 21.195 21.335 21.525 21.565 ;
        RECT 20.295 20.995 21.525 21.335 ;
      LAYER mcon ;
        RECT 21.305 22.865 21.475 23.035 ;
      LAYER met1 ;
        RECT 21.245 23.020 21.535 23.065 ;
        RECT 21.690 23.020 22.010 23.080 ;
        RECT 21.245 22.880 22.010 23.020 ;
        RECT 21.245 22.835 21.535 22.880 ;
        RECT 21.690 22.820 22.010 22.880 ;
      LAYER via ;
        RECT 21.720 22.820 21.980 23.080 ;
      LAYER met2 ;
        RECT 21.710 33.635 21.990 34.005 ;
        RECT 21.780 23.110 21.920 33.635 ;
        RECT 21.720 22.790 21.980 23.110 ;
      LAYER via2 ;
        RECT 21.710 33.680 21.990 33.960 ;
      LAYER met3 ;
        RECT 21.685 33.970 22.015 33.985 ;
        RECT 21.685 33.670 41.400 33.970 ;
        RECT 21.685 33.655 22.015 33.670 ;
    END
  END y[17]
  PIN y[16]
    ANTENNADIFFAREA 0.439000 ;
    PORT
      LAYER li1 ;
        RECT 21.245 25.295 21.940 25.925 ;
        RECT 21.770 24.695 21.940 25.295 ;
        RECT 21.675 23.715 22.005 24.695 ;
      LAYER mcon ;
        RECT 21.765 25.585 21.935 25.755 ;
      LAYER met1 ;
        RECT 21.705 25.740 21.995 25.785 ;
        RECT 23.530 25.740 23.850 25.800 ;
        RECT 21.705 25.600 23.850 25.740 ;
        RECT 21.705 25.555 21.995 25.600 ;
        RECT 23.530 25.540 23.850 25.600 ;
      LAYER via ;
        RECT 23.560 25.540 23.820 25.800 ;
      LAYER met2 ;
        RECT 23.550 31.805 23.830 32.175 ;
        RECT 23.620 25.830 23.760 31.805 ;
        RECT 23.560 25.510 23.820 25.830 ;
      LAYER via2 ;
        RECT 23.550 31.850 23.830 32.130 ;
      LAYER met3 ;
        RECT 23.525 32.140 23.855 32.155 ;
        RECT 23.525 31.840 41.400 32.140 ;
        RECT 23.525 31.825 23.855 31.840 ;
    END
  END y[16]
  PIN y[15]
    ANTENNADIFFAREA 0.795000 ;
    PORT
      LAYER li1 ;
        RECT 24.465 25.355 25.160 25.925 ;
        RECT 24.885 24.685 25.055 25.355 ;
        RECT 24.885 24.515 26.165 24.685 ;
        RECT 24.965 23.715 25.295 24.515 ;
        RECT 25.835 23.715 26.165 24.515 ;
      LAYER mcon ;
        RECT 25.905 24.225 26.075 24.395 ;
      LAYER met1 ;
        RECT 30.980 24.580 34.340 24.720 ;
        RECT 25.845 24.380 26.135 24.425 ;
        RECT 30.980 24.380 31.120 24.580 ;
        RECT 25.845 24.240 26.980 24.380 ;
        RECT 25.845 24.195 26.135 24.240 ;
        RECT 26.840 24.210 26.980 24.240 ;
        RECT 30.060 24.240 31.120 24.380 ;
        RECT 34.200 24.380 34.340 24.580 ;
        RECT 35.030 24.380 35.350 24.440 ;
        RECT 34.200 24.240 35.350 24.380 ;
        RECT 30.060 24.210 30.200 24.240 ;
        RECT 26.840 24.070 30.200 24.210 ;
        RECT 35.030 24.180 35.350 24.240 ;
      LAYER via ;
        RECT 35.060 24.180 35.320 24.440 ;
      LAYER met2 ;
        RECT 35.050 29.975 35.330 30.345 ;
        RECT 35.120 24.470 35.260 29.975 ;
        RECT 35.060 24.150 35.320 24.470 ;
      LAYER via2 ;
        RECT 35.050 30.020 35.330 30.300 ;
      LAYER met3 ;
        RECT 35.025 30.310 35.355 30.325 ;
        RECT 35.025 30.010 41.400 30.310 ;
        RECT 35.025 29.995 35.355 30.010 ;
    END
  END y[15]
  PIN y[14]
    ANTENNADIFFAREA 0.699000 ;
    PORT
      LAYER li1 ;
        RECT 27.235 25.585 28.465 25.925 ;
        RECT 27.235 25.355 27.565 25.585 ;
        RECT 28.285 24.685 28.465 25.585 ;
        RECT 27.235 24.515 28.465 24.685 ;
        RECT 27.235 23.715 27.565 24.515 ;
        RECT 28.135 23.715 28.465 24.515 ;
      LAYER mcon ;
        RECT 28.205 25.585 28.375 25.755 ;
      LAYER met1 ;
        RECT 28.130 25.740 28.450 25.800 ;
        RECT 27.855 25.600 28.450 25.740 ;
        RECT 28.130 25.540 28.450 25.600 ;
      LAYER via ;
        RECT 28.160 25.540 28.420 25.800 ;
      LAYER met2 ;
        RECT 28.150 28.145 28.430 28.515 ;
        RECT 28.220 25.830 28.360 28.145 ;
        RECT 28.160 25.510 28.420 25.830 ;
      LAYER via2 ;
        RECT 28.150 28.190 28.430 28.470 ;
      LAYER met3 ;
        RECT 28.125 28.480 28.455 28.495 ;
        RECT 28.125 28.180 41.400 28.480 ;
        RECT 28.125 28.165 28.455 28.180 ;
    END
  END y[14]
  PIN y[13]
    ANTENNADIFFAREA 0.795000 ;
    PORT
      LAYER li1 ;
        RECT 25.355 22.405 25.685 23.205 ;
        RECT 26.225 22.405 26.555 23.205 ;
        RECT 25.355 22.235 26.635 22.405 ;
        RECT 26.465 21.565 26.635 22.235 ;
        RECT 26.360 20.995 27.055 21.565 ;
      LAYER mcon ;
        RECT 26.365 22.865 26.535 23.035 ;
      LAYER met1 ;
        RECT 26.290 23.020 26.610 23.080 ;
        RECT 26.015 22.880 26.610 23.020 ;
        RECT 26.290 22.820 26.610 22.880 ;
      LAYER via ;
        RECT 26.320 22.820 26.580 23.080 ;
      LAYER met2 ;
        RECT 26.310 25.095 26.590 25.465 ;
        RECT 26.380 23.110 26.520 25.095 ;
        RECT 26.320 22.790 26.580 23.110 ;
      LAYER via2 ;
        RECT 26.310 25.140 26.590 25.420 ;
      LAYER met3 ;
        RECT 39.640 26.350 41.400 26.650 ;
        RECT 26.285 25.430 26.615 25.445 ;
        RECT 39.640 25.430 39.940 26.350 ;
        RECT 26.285 25.130 39.940 25.430 ;
        RECT 26.285 25.115 26.615 25.130 ;
    END
  END y[13]
  PIN y[12]
    ANTENNADIFFAREA 0.699000 ;
    PORT
      LAYER li1 ;
        RECT 29.495 22.405 29.825 23.205 ;
        RECT 30.395 22.405 30.725 23.205 ;
        RECT 29.495 22.235 30.725 22.405 ;
        RECT 29.495 21.335 29.675 22.235 ;
        RECT 30.395 21.335 30.725 21.565 ;
        RECT 29.495 20.995 30.725 21.335 ;
      LAYER mcon ;
        RECT 30.505 22.865 30.675 23.035 ;
      LAYER met1 ;
        RECT 30.445 23.020 30.735 23.065 ;
        RECT 35.950 23.020 36.270 23.080 ;
        RECT 30.445 22.880 31.580 23.020 ;
        RECT 30.445 22.835 30.735 22.880 ;
        RECT 31.440 22.680 31.580 22.880 ;
        RECT 35.120 22.880 36.270 23.020 ;
        RECT 35.120 22.680 35.260 22.880 ;
        RECT 35.950 22.820 36.270 22.880 ;
        RECT 31.440 22.540 35.260 22.680 ;
      LAYER via ;
        RECT 35.980 22.820 36.240 23.080 ;
      LAYER met2 ;
        RECT 35.970 23.875 36.250 24.245 ;
        RECT 36.040 23.110 36.180 23.875 ;
        RECT 35.980 22.790 36.240 23.110 ;
      LAYER via2 ;
        RECT 35.970 23.920 36.250 24.200 ;
      LAYER met3 ;
        RECT 35.945 24.210 36.275 24.225 ;
        RECT 35.945 23.910 41.400 24.210 ;
        RECT 35.945 23.895 36.275 23.910 ;
    END
  END y[12]
  PIN y[11]
    ANTENNADIFFAREA 0.699000 ;
    PORT
      LAYER li1 ;
        RECT 27.235 22.405 27.565 23.205 ;
        RECT 28.135 22.405 28.465 23.205 ;
        RECT 27.235 22.235 28.465 22.405 ;
        RECT 27.235 21.335 27.565 21.565 ;
        RECT 28.285 21.335 28.465 22.235 ;
        RECT 27.235 20.995 28.465 21.335 ;
      LAYER mcon ;
        RECT 28.205 21.165 28.375 21.335 ;
      LAYER met1 ;
        RECT 30.980 21.860 39.400 22.000 ;
        RECT 28.145 21.320 28.435 21.365 ;
        RECT 30.980 21.320 31.120 21.860 ;
        RECT 28.145 21.180 31.120 21.320 ;
        RECT 39.260 21.320 39.400 21.860 ;
        RECT 40.090 21.320 40.410 21.380 ;
        RECT 39.260 21.180 40.410 21.320 ;
        RECT 28.145 21.135 28.435 21.180 ;
        RECT 40.090 21.120 40.410 21.180 ;
      LAYER via ;
        RECT 40.120 21.120 40.380 21.380 ;
      LAYER met2 ;
        RECT 40.110 22.045 40.390 22.415 ;
        RECT 40.180 21.410 40.320 22.045 ;
        RECT 40.120 21.090 40.380 21.410 ;
      LAYER via2 ;
        RECT 40.110 22.090 40.390 22.370 ;
      LAYER met3 ;
        RECT 40.085 22.380 40.415 22.395 ;
        RECT 40.085 22.080 41.400 22.380 ;
        RECT 40.085 22.065 40.415 22.080 ;
    END
  END y[11]
  PIN y[10]
    ANTENNADIFFAREA 0.439000 ;
    PORT
      LAYER li1 ;
        RECT 28.660 19.855 29.355 20.485 ;
        RECT 28.660 19.255 28.830 19.855 ;
        RECT 28.595 18.275 28.925 19.255 ;
      LAYER mcon ;
        RECT 29.125 20.145 29.295 20.315 ;
      LAYER met1 ;
        RECT 29.065 20.300 29.355 20.345 ;
        RECT 39.630 20.300 39.950 20.360 ;
        RECT 29.065 20.160 30.200 20.300 ;
        RECT 29.065 20.115 29.355 20.160 ;
        RECT 30.060 19.960 30.200 20.160 ;
        RECT 38.800 20.160 39.950 20.300 ;
        RECT 38.800 19.960 38.940 20.160 ;
        RECT 39.630 20.100 39.950 20.160 ;
        RECT 30.060 19.820 38.940 19.960 ;
      LAYER via ;
        RECT 39.660 20.100 39.920 20.360 ;
      LAYER met2 ;
        RECT 39.650 20.215 39.930 20.585 ;
        RECT 39.660 20.070 39.920 20.215 ;
      LAYER via2 ;
        RECT 39.650 20.260 39.930 20.540 ;
      LAYER met3 ;
        RECT 39.625 20.550 39.955 20.565 ;
        RECT 39.625 20.250 41.400 20.550 ;
        RECT 39.625 20.235 39.955 20.250 ;
    END
  END y[10]
  PIN y[9]
    ANTENNADIFFAREA 0.699000 ;
    PORT
      LAYER li1 ;
        RECT 25.355 20.145 26.585 20.485 ;
        RECT 25.355 19.245 25.535 20.145 ;
        RECT 26.255 19.915 26.585 20.145 ;
        RECT 25.355 19.075 26.585 19.245 ;
        RECT 25.355 18.275 25.685 19.075 ;
        RECT 26.255 18.275 26.585 19.075 ;
      LAYER mcon ;
        RECT 26.365 18.785 26.535 18.955 ;
      LAYER met1 ;
        RECT 30.060 19.140 35.720 19.280 ;
        RECT 26.305 18.940 26.595 18.985 ;
        RECT 30.060 18.940 30.200 19.140 ;
        RECT 26.305 18.800 30.200 18.940 ;
        RECT 35.580 18.940 35.720 19.140 ;
        RECT 36.410 18.940 36.730 19.000 ;
        RECT 35.580 18.800 36.730 18.940 ;
        RECT 26.305 18.755 26.595 18.800 ;
        RECT 36.410 18.740 36.730 18.800 ;
      LAYER via ;
        RECT 36.440 18.740 36.700 19.000 ;
      LAYER met2 ;
        RECT 36.440 18.755 36.700 19.030 ;
        RECT 36.430 18.385 36.710 18.755 ;
      LAYER via2 ;
        RECT 36.430 18.430 36.710 18.710 ;
      LAYER met3 ;
        RECT 36.405 18.720 36.735 18.735 ;
        RECT 36.405 18.420 41.400 18.720 ;
        RECT 36.405 18.405 36.735 18.420 ;
    END
  END y[9]
  PIN y[8]
    ANTENNADIFFAREA 0.439000 ;
    PORT
      LAYER li1 ;
        RECT 30.435 16.785 30.765 17.765 ;
        RECT 30.500 16.745 30.675 16.785 ;
        RECT 30.500 16.185 30.670 16.745 ;
        RECT 30.500 15.555 31.195 16.185 ;
      LAYER mcon ;
        RECT 30.505 16.745 30.675 16.915 ;
      LAYER met1 ;
        RECT 30.445 16.900 30.735 16.945 ;
        RECT 35.490 16.900 35.810 16.960 ;
        RECT 30.445 16.760 35.810 16.900 ;
        RECT 30.445 16.715 30.735 16.760 ;
        RECT 35.490 16.700 35.810 16.760 ;
      LAYER via ;
        RECT 35.520 16.700 35.780 16.960 ;
      LAYER met2 ;
        RECT 35.520 16.925 35.780 16.990 ;
        RECT 35.510 16.555 35.790 16.925 ;
        RECT 35.580 16.505 35.720 16.555 ;
      LAYER via2 ;
        RECT 35.510 16.600 35.790 16.880 ;
      LAYER met3 ;
        RECT 35.485 16.890 35.815 16.905 ;
        RECT 35.485 16.590 41.400 16.890 ;
        RECT 35.485 16.575 35.815 16.590 ;
    END
  END y[8]
  PIN y[7]
    ANTENNADIFFAREA 0.795000 ;
    PORT
      LAYER li1 ;
        RECT 26.345 16.965 26.675 17.765 ;
        RECT 27.215 16.965 27.545 17.765 ;
        RECT 26.265 16.795 27.545 16.965 ;
        RECT 26.265 16.125 26.435 16.795 ;
        RECT 25.845 15.555 26.540 16.125 ;
      LAYER mcon ;
        RECT 27.285 17.425 27.455 17.595 ;
      LAYER met1 ;
        RECT 27.225 17.580 27.515 17.625 ;
        RECT 40.090 17.580 40.410 17.640 ;
        RECT 27.225 17.440 28.360 17.580 ;
        RECT 27.225 17.395 27.515 17.440 ;
        RECT 28.220 17.410 28.360 17.440 ;
        RECT 35.580 17.440 40.410 17.580 ;
        RECT 35.580 17.410 35.720 17.440 ;
        RECT 28.220 17.270 35.720 17.410 ;
        RECT 40.090 17.380 40.410 17.440 ;
      LAYER via ;
        RECT 40.120 17.380 40.380 17.640 ;
      LAYER met2 ;
        RECT 40.120 17.350 40.380 17.670 ;
        RECT 40.180 15.095 40.320 17.350 ;
        RECT 40.110 14.725 40.390 15.095 ;
      LAYER via2 ;
        RECT 40.110 14.770 40.390 15.050 ;
      LAYER met3 ;
        RECT 40.085 15.060 40.415 15.075 ;
        RECT 40.085 14.760 41.400 15.060 ;
        RECT 40.085 14.745 40.415 14.760 ;
    END
  END y[7]
  PIN y[6]
    ANTENNADIFFAREA 0.699000 ;
    PORT
      LAYER li1 ;
        RECT 28.155 16.965 28.485 17.765 ;
        RECT 29.055 16.965 29.385 17.765 ;
        RECT 28.155 16.795 29.385 16.965 ;
        RECT 28.155 15.895 28.485 16.125 ;
        RECT 29.205 15.895 29.385 16.795 ;
        RECT 28.155 15.555 29.385 15.895 ;
      LAYER mcon ;
        RECT 28.205 15.725 28.375 15.895 ;
      LAYER met1 ;
        RECT 30.980 16.080 35.260 16.220 ;
        RECT 28.145 15.880 28.435 15.925 ;
        RECT 30.980 15.880 31.120 16.080 ;
        RECT 28.145 15.740 31.120 15.880 ;
        RECT 35.120 15.880 35.260 16.080 ;
        RECT 35.950 15.880 36.270 15.940 ;
        RECT 35.120 15.740 36.270 15.880 ;
        RECT 28.145 15.695 28.435 15.740 ;
        RECT 35.950 15.680 36.270 15.740 ;
      LAYER via ;
        RECT 35.980 15.680 36.240 15.940 ;
      LAYER met2 ;
        RECT 35.980 15.650 36.240 15.970 ;
        RECT 36.040 12.655 36.180 15.650 ;
        RECT 35.970 12.285 36.250 12.655 ;
      LAYER via2 ;
        RECT 35.970 12.330 36.250 12.610 ;
      LAYER met3 ;
        RECT 35.945 12.620 36.275 12.635 ;
        RECT 35.945 12.320 41.400 12.620 ;
        RECT 35.945 12.305 36.275 12.320 ;
    END
  END y[6]
  PIN y[5]
    ANTENNADIFFAREA 0.795000 ;
    PORT
      LAYER li1 ;
        RECT 24.005 14.475 24.700 15.045 ;
        RECT 24.425 13.805 24.595 14.475 ;
        RECT 24.425 13.635 25.705 13.805 ;
        RECT 24.505 12.835 24.835 13.635 ;
        RECT 25.375 12.835 25.705 13.635 ;
      LAYER mcon ;
        RECT 25.445 13.005 25.615 13.175 ;
      LAYER met1 ;
        RECT 25.370 13.160 25.690 13.220 ;
        RECT 25.095 13.020 25.690 13.160 ;
        RECT 25.370 12.960 25.690 13.020 ;
      LAYER via ;
        RECT 25.400 12.960 25.660 13.220 ;
      LAYER met2 ;
        RECT 25.400 12.930 25.660 13.250 ;
        RECT 25.460 10.825 25.600 12.930 ;
        RECT 25.390 10.455 25.670 10.825 ;
      LAYER via2 ;
        RECT 25.390 10.500 25.670 10.780 ;
      LAYER met3 ;
        RECT 25.365 10.790 25.695 10.805 ;
        RECT 25.365 10.490 41.400 10.790 ;
        RECT 25.365 10.475 25.695 10.490 ;
    END
  END y[5]
  PIN y[4]
    ANTENNADIFFAREA 0.699000 ;
    PORT
      LAYER li1 ;
        RECT 24.015 11.525 24.345 12.325 ;
        RECT 24.915 11.525 25.245 12.325 ;
        RECT 24.015 11.355 25.245 11.525 ;
        RECT 24.015 10.455 24.345 10.685 ;
        RECT 25.065 10.455 25.245 11.355 ;
        RECT 24.015 10.115 25.245 10.455 ;
      LAYER mcon ;
        RECT 24.065 10.285 24.235 10.455 ;
      LAYER met1 ;
        RECT 23.990 10.440 24.310 10.500 ;
        RECT 23.715 10.300 24.310 10.440 ;
        RECT 23.990 10.240 24.310 10.300 ;
      LAYER via ;
        RECT 24.020 10.240 24.280 10.500 ;
      LAYER met2 ;
        RECT 24.020 10.210 24.280 10.530 ;
        RECT 24.080 9.760 24.220 10.210 ;
        RECT 24.080 9.620 24.680 9.760 ;
        RECT 24.540 8.995 24.680 9.620 ;
        RECT 24.470 8.625 24.750 8.995 ;
      LAYER via2 ;
        RECT 24.470 8.670 24.750 8.950 ;
      LAYER met3 ;
        RECT 24.445 8.960 24.775 8.975 ;
        RECT 24.445 8.660 41.400 8.960 ;
        RECT 24.445 8.645 24.775 8.660 ;
    END
  END y[4]
  PIN y[3]
    ANTENNADIFFAREA 0.699000 ;
    PORT
      LAYER li1 ;
        RECT 27.695 11.525 28.025 12.325 ;
        RECT 28.595 11.525 28.925 12.325 ;
        RECT 27.695 11.355 28.925 11.525 ;
        RECT 27.695 10.455 28.025 10.685 ;
        RECT 28.745 10.455 28.925 11.355 ;
        RECT 27.695 10.115 28.925 10.455 ;
      LAYER mcon ;
        RECT 28.665 10.285 28.835 10.455 ;
      LAYER met1 ;
        RECT 28.590 10.440 28.910 10.500 ;
        RECT 28.315 10.300 28.910 10.440 ;
        RECT 28.590 10.240 28.910 10.300 ;
      LAYER via ;
        RECT 28.620 10.240 28.880 10.500 ;
      LAYER met2 ;
        RECT 28.620 10.210 28.880 10.530 ;
        RECT 28.680 7.165 28.820 10.210 ;
        RECT 28.610 6.795 28.890 7.165 ;
      LAYER via2 ;
        RECT 28.610 6.840 28.890 7.120 ;
      LAYER met3 ;
        RECT 28.585 7.130 28.915 7.145 ;
        RECT 28.585 6.830 41.400 7.130 ;
        RECT 28.585 6.815 28.915 6.830 ;
    END
  END y[3]
  PIN y[2]
    ANTENNADIFFAREA 0.439000 ;
    PORT
      LAYER li1 ;
        RECT 28.660 14.415 29.355 15.045 ;
        RECT 28.660 13.815 28.830 14.415 ;
        RECT 28.595 12.835 28.925 13.815 ;
      LAYER mcon ;
        RECT 28.665 13.005 28.835 13.175 ;
      LAYER met1 ;
        RECT 28.605 13.160 28.895 13.205 ;
        RECT 29.510 13.160 29.830 13.220 ;
        RECT 28.605 13.020 29.830 13.160 ;
        RECT 28.605 12.975 28.895 13.020 ;
        RECT 29.510 12.960 29.830 13.020 ;
      LAYER via ;
        RECT 29.540 12.960 29.800 13.220 ;
      LAYER met2 ;
        RECT 29.540 12.930 29.800 13.250 ;
        RECT 29.600 11.120 29.740 12.930 ;
        RECT 29.600 10.980 30.200 11.120 ;
        RECT 30.060 6.360 30.200 10.980 ;
        RECT 29.600 6.220 30.200 6.360 ;
        RECT 29.600 5.335 29.740 6.220 ;
        RECT 29.530 4.965 29.810 5.335 ;
      LAYER via2 ;
        RECT 29.530 5.010 29.810 5.290 ;
      LAYER met3 ;
        RECT 29.505 5.300 29.835 5.315 ;
        RECT 29.505 5.000 41.400 5.300 ;
        RECT 29.505 4.985 29.835 5.000 ;
    END
  END y[2]
  PIN y[1]
    ANTENNADIFFAREA 0.699000 ;
    PORT
      LAYER li1 ;
        RECT 25.855 11.525 26.185 12.325 ;
        RECT 26.755 11.525 27.085 12.325 ;
        RECT 25.855 11.355 27.085 11.525 ;
        RECT 25.855 10.455 26.185 10.685 ;
        RECT 26.905 10.455 27.085 11.355 ;
        RECT 25.855 10.115 27.085 10.455 ;
      LAYER mcon ;
        RECT 25.905 10.285 26.075 10.455 ;
      LAYER met1 ;
        RECT 25.830 10.440 26.150 10.500 ;
        RECT 25.555 10.300 26.150 10.440 ;
        RECT 25.830 10.240 26.150 10.300 ;
      LAYER via ;
        RECT 25.860 10.240 26.120 10.500 ;
      LAYER met2 ;
        RECT 25.860 10.210 26.120 10.530 ;
        RECT 25.920 3.505 26.060 10.210 ;
        RECT 25.850 3.135 26.130 3.505 ;
      LAYER via2 ;
        RECT 25.850 3.180 26.130 3.460 ;
      LAYER met3 ;
        RECT 25.825 3.470 26.155 3.485 ;
        RECT 25.825 3.170 41.400 3.470 ;
        RECT 25.825 3.155 26.155 3.170 ;
    END
  END y[1]
  PIN y[0]
    ANTENNADIFFAREA 0.439000 ;
    PORT
      LAYER li1 ;
        RECT 22.135 11.345 22.465 12.325 ;
        RECT 22.230 10.745 22.400 11.345 ;
        RECT 21.705 10.115 22.400 10.745 ;
      LAYER mcon ;
        RECT 21.765 10.285 21.935 10.455 ;
      LAYER met1 ;
        RECT 21.690 10.440 22.010 10.500 ;
        RECT 21.415 10.300 22.010 10.440 ;
        RECT 21.690 10.240 22.010 10.300 ;
      LAYER via ;
        RECT 21.720 10.240 21.980 10.500 ;
      LAYER met2 ;
        RECT 21.720 10.210 21.980 10.530 ;
        RECT 21.780 1.675 21.920 10.210 ;
        RECT 21.710 1.305 21.990 1.675 ;
      LAYER via2 ;
        RECT 21.710 1.350 21.990 1.630 ;
      LAYER met3 ;
        RECT 21.685 1.640 22.015 1.655 ;
        RECT 21.685 1.340 41.400 1.640 ;
        RECT 21.685 1.325 22.015 1.340 ;
    END
  END y[0]
  OBS
      LAYER pwell ;
        RECT 12.100 26.075 12.270 26.265 ;
        RECT 14.400 26.075 14.570 26.265 ;
        RECT 14.870 26.075 15.040 26.265 ;
        RECT 17.195 26.120 17.305 26.240 ;
        RECT 19.010 26.075 19.180 26.265 ;
        RECT 20.395 26.120 20.555 26.230 ;
        RECT 22.230 26.075 22.400 26.265 ;
        RECT 22.680 26.125 22.800 26.235 ;
        RECT 23.615 26.120 23.775 26.230 ;
        RECT 26.360 26.075 26.530 26.265 ;
        RECT 26.820 26.125 26.940 26.235 ;
        RECT 28.660 26.075 28.830 26.265 ;
        RECT 29.120 26.125 29.240 26.235 ;
        RECT 30.055 26.120 30.215 26.230 ;
        RECT 30.960 26.125 31.080 26.235 ;
        RECT 10.135 25.205 10.565 25.990 ;
        RECT 10.585 25.165 12.415 26.075 ;
        RECT 12.425 25.165 14.715 26.075 ;
        RECT 14.725 25.165 16.555 26.075 ;
        RECT 16.575 25.205 17.005 25.990 ;
        RECT 18.865 25.165 20.215 26.075 ;
        RECT 21.165 25.165 22.515 26.075 ;
        RECT 23.015 25.205 23.445 25.990 ;
        RECT 24.385 25.165 26.675 26.075 ;
        RECT 27.145 25.165 28.975 26.075 ;
        RECT 29.455 25.205 29.885 25.990 ;
      LAYER nwell ;
        RECT 9.930 22.045 31.470 24.875 ;
      LAYER pwell ;
        RECT 10.135 20.930 10.565 21.715 ;
        RECT 10.585 20.845 12.415 21.755 ;
        RECT 12.445 20.845 13.795 21.755 ;
        RECT 13.825 20.845 15.175 21.755 ;
        RECT 15.645 20.845 17.475 21.755 ;
        RECT 18.425 20.845 19.775 21.755 ;
        RECT 19.785 20.845 21.615 21.755 ;
        RECT 21.645 20.845 22.995 21.755 ;
        RECT 23.015 20.930 23.445 21.715 ;
        RECT 23.485 20.845 24.835 21.755 ;
        RECT 24.845 20.845 27.135 21.755 ;
        RECT 27.145 20.845 28.975 21.755 ;
        RECT 28.985 20.845 30.815 21.755 ;
        RECT 10.730 20.655 10.900 20.845 ;
        RECT 11.185 20.655 11.355 20.825 ;
        RECT 11.650 20.635 11.820 20.825 ;
        RECT 12.560 20.655 12.730 20.845 ;
        RECT 13.495 20.680 13.655 20.790 ;
        RECT 13.940 20.655 14.110 20.845 ;
        RECT 14.410 20.635 14.580 20.825 ;
        RECT 15.320 20.685 15.440 20.795 ;
        RECT 15.795 20.680 15.955 20.790 ;
        RECT 17.160 20.655 17.330 20.845 ;
        RECT 19.460 20.825 19.630 20.845 ;
        RECT 17.635 20.690 17.795 20.800 ;
        RECT 19.000 20.635 19.170 20.825 ;
        RECT 19.460 20.655 19.635 20.825 ;
        RECT 19.930 20.655 20.100 20.845 ;
        RECT 20.845 20.655 21.015 20.825 ;
        RECT 21.760 20.655 21.930 20.845 ;
        RECT 23.145 20.655 23.315 20.825 ;
        RECT 24.520 20.655 24.690 20.845 ;
        RECT 20.940 20.635 21.015 20.655 ;
        RECT 24.990 20.635 25.160 20.845 ;
        RECT 27.740 20.635 27.910 20.825 ;
        RECT 28.200 20.635 28.370 20.825 ;
        RECT 28.660 20.655 28.830 20.845 ;
        RECT 29.130 20.655 29.300 20.845 ;
        RECT 30.055 20.680 30.215 20.790 ;
        RECT 30.960 20.685 31.080 20.795 ;
        RECT 10.125 19.955 11.080 20.635 ;
        RECT 11.505 19.725 13.335 20.635 ;
        RECT 14.265 19.725 15.615 20.635 ;
        RECT 16.575 19.765 17.005 20.550 ;
        RECT 17.025 19.725 19.315 20.635 ;
        RECT 19.740 19.955 20.695 20.635 ;
        RECT 20.940 19.955 22.775 20.635 ;
        RECT 23.420 19.955 24.375 20.635 ;
        RECT 21.425 19.725 22.775 19.955 ;
        RECT 24.845 19.725 26.675 20.635 ;
        RECT 26.705 19.725 28.055 20.635 ;
        RECT 28.085 19.725 29.435 20.635 ;
        RECT 29.455 19.765 29.885 20.550 ;
      LAYER nwell ;
        RECT 9.930 16.605 31.470 19.435 ;
      LAYER pwell ;
        RECT 10.135 15.490 10.565 16.275 ;
        RECT 11.965 15.405 13.315 16.315 ;
        RECT 13.345 15.405 15.175 16.315 ;
        RECT 15.405 16.085 16.755 16.315 ;
        RECT 15.405 15.405 17.240 16.085 ;
        RECT 17.485 15.405 18.835 16.315 ;
        RECT 18.885 15.405 20.235 16.315 ;
        RECT 23.015 15.490 23.445 16.275 ;
        RECT 24.185 16.085 25.535 16.315 ;
        RECT 23.700 15.405 25.535 16.085 ;
        RECT 25.765 15.405 28.055 16.315 ;
        RECT 28.065 15.405 29.895 16.315 ;
        RECT 29.925 15.405 31.275 16.315 ;
        RECT 10.260 15.245 10.380 15.355 ;
        RECT 10.730 15.195 10.900 15.385 ;
        RECT 11.640 15.245 11.760 15.355 ;
        RECT 12.110 15.215 12.280 15.405 ;
        RECT 13.020 15.245 13.140 15.355 ;
        RECT 13.490 15.195 13.660 15.405 ;
        RECT 17.165 15.385 17.240 15.405 ;
        RECT 17.630 15.385 17.800 15.405 ;
        RECT 16.240 15.195 16.410 15.385 ;
        RECT 17.165 15.355 17.335 15.385 ;
        RECT 17.160 15.245 17.335 15.355 ;
        RECT 17.165 15.215 17.335 15.245 ;
        RECT 17.625 15.215 17.800 15.385 ;
        RECT 19.920 15.195 20.090 15.405 ;
        RECT 23.700 15.385 23.775 15.405 ;
        RECT 20.385 15.215 20.555 15.385 ;
        RECT 22.235 15.250 22.395 15.360 ;
        RECT 22.685 15.215 22.855 15.385 ;
        RECT 23.605 15.215 23.775 15.385 ;
        RECT 20.480 15.195 20.555 15.215 ;
        RECT 25.900 15.195 26.070 15.385 ;
        RECT 26.360 15.245 26.480 15.355 ;
        RECT 27.740 15.195 27.910 15.405 ;
        RECT 28.200 15.195 28.370 15.385 ;
        RECT 29.580 15.215 29.750 15.405 ;
        RECT 30.040 15.350 30.210 15.405 ;
        RECT 30.040 15.240 30.215 15.350 ;
        RECT 30.960 15.245 31.080 15.355 ;
        RECT 30.040 15.215 30.210 15.240 ;
        RECT 10.585 14.285 12.875 15.195 ;
        RECT 13.345 14.285 15.175 15.195 ;
        RECT 15.205 14.285 16.555 15.195 ;
        RECT 16.575 14.325 17.005 15.110 ;
        RECT 17.900 14.515 18.855 15.195 ;
        RECT 18.885 14.285 20.235 15.195 ;
        RECT 20.480 14.515 22.315 15.195 ;
        RECT 22.960 14.515 23.915 15.195 ;
        RECT 20.965 14.285 22.315 14.515 ;
        RECT 23.925 14.285 26.215 15.195 ;
        RECT 26.705 14.285 28.055 15.195 ;
        RECT 28.085 14.285 29.435 15.195 ;
        RECT 29.455 14.325 29.885 15.110 ;
      LAYER nwell ;
        RECT 9.930 11.165 31.470 13.995 ;
      LAYER pwell ;
        RECT 10.135 10.050 10.565 10.835 ;
        RECT 10.585 9.965 12.875 10.875 ;
        RECT 15.205 9.965 16.555 10.875 ;
        RECT 16.575 10.050 17.005 10.835 ;
        RECT 17.945 10.195 19.780 10.875 ;
        RECT 18.090 9.965 19.780 10.195 ;
        RECT 20.265 9.965 21.615 10.875 ;
        RECT 21.625 9.965 22.975 10.875 ;
        RECT 23.015 10.050 23.445 10.835 ;
        RECT 23.925 9.965 25.755 10.875 ;
        RECT 25.765 9.965 27.595 10.875 ;
        RECT 27.605 9.965 29.435 10.875 ;
        RECT 29.455 10.050 29.885 10.835 ;
        RECT 10.730 9.775 10.900 9.965 ;
        RECT 13.055 9.800 13.165 9.920 ;
        RECT 14.860 9.805 14.980 9.915 ;
        RECT 15.320 9.775 15.490 9.965 ;
        RECT 17.175 9.810 17.335 9.920 ;
        RECT 18.090 9.775 18.260 9.965 ;
        RECT 21.300 9.775 21.470 9.965 ;
        RECT 22.690 9.775 22.860 9.965 ;
        RECT 23.600 9.805 23.720 9.915 ;
        RECT 25.440 9.775 25.610 9.965 ;
        RECT 27.280 9.775 27.450 9.965 ;
        RECT 29.120 9.775 29.290 9.965 ;
        RECT 30.055 9.810 30.215 9.920 ;
        RECT 30.960 9.805 31.080 9.915 ;
      LAYER li1 ;
        RECT 10.120 26.095 31.280 26.265 ;
        RECT 10.205 25.370 10.495 26.095 ;
        RECT 12.075 25.605 12.330 26.095 ;
        RECT 12.090 24.855 12.310 25.435 ;
        RECT 13.910 25.185 14.125 25.880 ;
        RECT 14.295 25.355 14.630 26.095 ;
        RECT 14.810 25.605 15.065 26.095 ;
        RECT 13.745 24.855 14.125 25.185 ;
        RECT 15.585 24.855 15.960 25.415 ;
        RECT 16.645 25.370 16.935 26.095 ;
        RECT 18.965 25.285 19.205 26.095 ;
        RECT 19.375 25.285 19.705 25.925 ;
        RECT 19.875 25.285 20.145 26.095 ;
        RECT 22.145 25.295 22.455 26.095 ;
        RECT 23.085 25.370 23.375 26.095 ;
        RECT 16.165 25.075 16.475 25.185 ;
        RECT 16.165 24.905 18.715 25.075 ;
        RECT 16.165 24.855 16.475 24.905 ;
        RECT 10.205 23.545 10.495 24.710 ;
        RECT 11.175 23.545 11.405 24.345 ;
        RECT 12.075 23.545 12.330 24.685 ;
        RECT 12.525 23.545 12.805 24.345 ;
        RECT 13.535 23.545 13.705 24.345 ;
        RECT 14.375 23.545 14.635 24.685 ;
        RECT 14.810 23.545 15.065 24.685 ;
        RECT 15.735 23.545 15.965 24.345 ;
        RECT 16.645 23.545 16.935 24.710 ;
        RECT 18.545 24.395 18.715 24.905 ;
        RECT 19.465 24.685 19.635 25.285 ;
        RECT 25.870 25.185 26.085 25.880 ;
        RECT 26.255 25.355 26.590 26.095 ;
        RECT 28.635 25.605 28.890 26.095 ;
        RECT 21.265 25.075 21.600 25.105 ;
        RECT 20.845 24.905 21.600 25.075 ;
        RECT 18.955 24.515 19.635 24.685 ;
        RECT 18.955 24.395 19.285 24.515 ;
        RECT 18.545 24.225 19.285 24.395 ;
        RECT 18.955 23.730 19.285 24.225 ;
        RECT 19.815 23.545 20.145 24.685 ;
        RECT 20.845 24.565 21.015 24.905 ;
        RECT 21.265 24.855 21.600 24.905 ;
        RECT 22.110 25.075 22.445 25.125 ;
        RECT 22.110 24.905 22.855 25.075 ;
        RECT 22.110 24.855 22.445 24.905 ;
        RECT 21.245 23.545 21.505 24.685 ;
        RECT 22.175 23.545 22.455 24.685 ;
        RECT 22.685 24.225 22.855 24.905 ;
        RECT 25.705 24.855 26.085 25.185 ;
        RECT 26.825 25.075 26.995 25.415 ;
        RECT 27.225 25.075 27.535 25.185 ;
        RECT 26.825 24.905 27.535 25.075 ;
        RECT 27.225 24.855 27.535 24.905 ;
        RECT 28.650 24.855 28.870 25.435 ;
        RECT 29.525 25.370 29.815 26.095 ;
        RECT 23.085 23.545 23.375 24.710 ;
        RECT 24.485 23.545 24.765 24.345 ;
        RECT 25.495 23.545 25.665 24.345 ;
        RECT 26.335 23.545 26.595 24.685 ;
        RECT 27.735 23.545 27.965 24.345 ;
        RECT 28.635 23.545 28.890 24.685 ;
        RECT 29.525 23.545 29.815 24.710 ;
        RECT 10.120 23.375 31.280 23.545 ;
        RECT 10.205 22.210 10.495 23.375 ;
        RECT 10.670 22.235 10.925 23.375 ;
        RECT 11.595 22.575 11.825 23.375 ;
        RECT 12.505 22.235 12.785 23.375 ;
        RECT 13.455 22.235 13.715 23.375 ;
        RECT 13.885 22.235 14.165 23.375 ;
        RECT 14.835 22.235 15.095 23.375 ;
        RECT 16.235 22.575 16.465 23.375 ;
        RECT 10.690 22.015 10.910 22.065 ;
        RECT 9.345 21.845 10.910 22.015 ;
        RECT 9.345 19.975 9.515 21.845 ;
        RECT 10.205 20.825 10.495 21.550 ;
        RECT 10.690 21.485 10.910 21.845 ;
        RECT 11.445 21.505 11.820 22.065 ;
        RECT 12.515 21.795 12.850 22.065 ;
        RECT 13.360 22.015 13.695 22.065 ;
        RECT 13.895 22.015 14.230 22.065 ;
        RECT 13.360 21.845 14.230 22.015 ;
        RECT 13.360 21.815 13.695 21.845 ;
        RECT 13.895 21.795 14.230 21.845 ;
        RECT 14.740 21.815 15.075 22.065 ;
        RECT 15.325 22.015 15.495 22.355 ;
        RECT 17.135 22.235 17.390 23.375 ;
        RECT 18.495 22.235 18.825 23.375 ;
        RECT 19.355 22.405 19.685 23.190 ;
        RECT 19.005 22.235 19.685 22.405 ;
        RECT 19.870 22.235 20.125 23.375 ;
        RECT 20.795 22.575 21.025 23.375 ;
        RECT 21.705 22.235 21.985 23.375 ;
        RECT 22.655 22.235 22.915 23.375 ;
        RECT 15.725 22.015 16.035 22.065 ;
        RECT 15.325 21.845 16.035 22.015 ;
        RECT 15.725 21.735 16.035 21.845 ;
        RECT 10.670 20.825 10.925 21.315 ;
        RECT 12.505 20.825 12.815 21.625 ;
        RECT 13.885 20.825 14.195 21.625 ;
        RECT 17.150 21.485 17.370 22.065 ;
        RECT 19.005 21.635 19.175 22.235 ;
        RECT 23.085 22.210 23.375 23.375 ;
        RECT 23.555 22.235 23.885 23.375 ;
        RECT 24.415 22.405 24.745 23.190 ;
        RECT 24.065 22.235 24.745 22.405 ;
        RECT 24.925 22.235 25.185 23.375 ;
        RECT 25.855 22.575 26.025 23.375 ;
        RECT 26.755 22.575 27.035 23.375 ;
        RECT 27.735 22.575 27.965 23.375 ;
        RECT 28.635 22.235 28.890 23.375 ;
        RECT 29.070 22.235 29.325 23.375 ;
        RECT 29.995 22.575 30.225 23.375 ;
        RECT 19.345 22.015 19.695 22.065 ;
        RECT 19.890 22.015 20.110 22.065 ;
        RECT 19.345 21.845 20.110 22.015 ;
        RECT 19.345 21.815 19.695 21.845 ;
        RECT 17.135 20.825 17.390 21.315 ;
        RECT 18.495 20.825 18.765 21.635 ;
        RECT 18.935 20.995 19.265 21.635 ;
        RECT 19.435 20.825 19.675 21.635 ;
        RECT 19.890 21.485 20.110 21.845 ;
        RECT 20.645 21.505 21.020 22.065 ;
        RECT 21.715 21.795 22.050 22.065 ;
        RECT 22.560 21.815 22.895 22.065 ;
        RECT 24.065 21.635 24.235 22.235 ;
        RECT 24.405 22.015 24.755 22.065 ;
        RECT 24.950 22.015 25.235 22.065 ;
        RECT 24.405 21.845 25.235 22.015 ;
        RECT 24.405 21.815 24.755 21.845 ;
        RECT 24.950 21.735 25.235 21.845 ;
        RECT 25.985 21.735 26.295 22.065 ;
        RECT 19.870 20.825 20.125 21.315 ;
        RECT 21.705 20.825 22.015 21.625 ;
        RECT 23.085 20.825 23.375 21.550 ;
        RECT 23.555 20.825 23.825 21.635 ;
        RECT 23.995 20.995 24.325 21.635 ;
        RECT 24.495 20.825 24.735 21.635 ;
        RECT 25.985 21.565 26.190 21.735 ;
        RECT 24.930 20.825 25.265 21.565 ;
        RECT 25.840 21.040 26.190 21.565 ;
        RECT 28.650 21.485 28.870 22.065 ;
        RECT 29.845 21.505 30.220 22.065 ;
        RECT 30.425 22.015 30.735 22.065 ;
        RECT 30.425 21.845 32.055 22.015 ;
        RECT 30.425 21.735 30.735 21.845 ;
        RECT 28.635 20.825 28.890 21.315 ;
        RECT 29.070 20.825 29.325 21.315 ;
        RECT 10.120 20.655 31.280 20.825 ;
        RECT 10.205 20.150 10.490 20.655 ;
        RECT 10.660 19.980 10.985 20.485 ;
        RECT 11.590 20.165 11.845 20.655 ;
        RECT 10.205 19.975 10.985 19.980 ;
        RECT 9.345 19.805 10.985 19.975 ;
        RECT 9.345 16.575 9.515 19.805 ;
        RECT 10.205 19.450 10.985 19.805 ;
        RECT 10.205 18.105 10.485 19.075 ;
        RECT 10.655 18.275 10.985 19.450 ;
        RECT 11.610 19.415 11.830 19.995 ;
        RECT 14.365 19.845 14.605 20.655 ;
        RECT 14.775 19.845 15.105 20.485 ;
        RECT 15.275 19.845 15.545 20.655 ;
        RECT 16.645 19.930 16.935 20.655 ;
        RECT 17.970 19.915 18.320 20.440 ;
        RECT 18.895 19.915 19.230 20.655 ;
        RECT 19.835 19.980 20.160 20.485 ;
        RECT 20.330 20.150 20.615 20.655 ;
        RECT 21.030 20.195 21.375 20.370 ;
        RECT 14.865 19.245 15.035 19.845 ;
        RECT 17.970 19.745 18.175 19.915 ;
        RECT 17.865 19.415 18.175 19.745 ;
        RECT 18.925 19.415 19.210 19.745 ;
        RECT 19.835 19.450 20.615 19.980 ;
        RECT 11.155 18.105 11.415 19.075 ;
        RECT 11.590 18.105 11.845 19.245 ;
        RECT 14.355 19.075 15.035 19.245 ;
        RECT 12.515 18.105 12.745 18.905 ;
        RECT 14.355 18.290 14.685 19.075 ;
        RECT 15.215 18.105 15.545 19.245 ;
        RECT 16.645 18.105 16.935 19.270 ;
        RECT 17.125 18.105 17.405 18.905 ;
        RECT 18.135 18.105 18.305 18.905 ;
        RECT 18.975 18.105 19.235 19.245 ;
        RECT 19.405 18.105 19.665 19.075 ;
        RECT 19.835 18.275 20.165 19.450 ;
        RECT 20.800 19.415 21.025 20.015 ;
        RECT 21.195 19.230 21.375 20.195 ;
        RECT 21.555 19.845 21.765 20.655 ;
        RECT 21.935 20.015 22.265 20.485 ;
        RECT 22.435 20.185 22.820 20.655 ;
        RECT 21.935 19.845 22.915 20.015 ;
        RECT 22.235 19.495 22.565 19.665 ;
        RECT 22.235 19.230 22.405 19.495 ;
        RECT 22.735 19.295 22.915 19.845 ;
        RECT 20.335 18.105 20.615 19.075 ;
        RECT 21.115 19.060 22.405 19.230 ;
        RECT 22.685 19.125 22.915 19.295 ;
        RECT 21.115 18.835 21.375 19.060 ;
        RECT 22.735 18.890 22.915 19.125 ;
        RECT 23.515 19.980 23.840 20.485 ;
        RECT 24.010 20.150 24.295 20.655 ;
        RECT 23.515 19.975 24.295 19.980 ;
        RECT 24.525 19.975 24.695 20.315 ;
        RECT 24.930 20.165 25.185 20.655 ;
        RECT 24.950 19.975 25.170 19.995 ;
        RECT 23.515 19.805 25.170 19.975 ;
        RECT 23.515 19.450 24.295 19.805 ;
        RECT 21.575 18.105 21.905 18.885 ;
        RECT 22.355 18.275 22.915 18.890 ;
        RECT 23.085 18.105 23.345 19.075 ;
        RECT 23.515 18.275 23.845 19.450 ;
        RECT 24.950 19.415 25.170 19.805 ;
        RECT 25.705 19.415 26.080 19.975 ;
        RECT 26.775 19.845 27.045 20.655 ;
        RECT 27.215 19.845 27.545 20.485 ;
        RECT 27.715 19.845 27.955 20.655 ;
        RECT 28.145 19.855 28.455 20.655 ;
        RECT 29.525 19.930 29.815 20.655 ;
        RECT 27.285 19.245 27.455 19.845 ;
        RECT 28.155 19.415 28.490 19.685 ;
        RECT 29.000 19.415 29.335 19.665 ;
        RECT 24.015 18.105 24.295 19.075 ;
        RECT 24.930 18.105 25.185 19.245 ;
        RECT 25.855 18.105 26.085 18.905 ;
        RECT 26.775 18.105 27.105 19.245 ;
        RECT 27.285 19.075 27.965 19.245 ;
        RECT 27.635 18.290 27.965 19.075 ;
        RECT 28.145 18.105 28.425 19.245 ;
        RECT 29.095 18.105 29.355 19.245 ;
        RECT 29.525 18.105 29.815 19.270 ;
        RECT 10.120 17.935 31.280 18.105 ;
        RECT 10.205 16.770 10.495 17.935 ;
        RECT 12.055 16.965 12.385 17.750 ;
        RECT 12.055 16.795 12.735 16.965 ;
        RECT 12.915 16.795 13.245 17.935 ;
        RECT 13.430 16.795 13.685 17.935 ;
        RECT 14.355 17.135 14.585 17.935 ;
        RECT 15.265 17.150 15.825 17.765 ;
        RECT 16.275 17.155 16.605 17.935 ;
        RECT 12.045 16.575 12.395 16.625 ;
        RECT 9.345 16.405 12.395 16.575 ;
        RECT 9.345 14.195 9.515 16.405 ;
        RECT 12.045 16.375 12.395 16.405 ;
        RECT 12.565 16.195 12.735 16.795 ;
        RECT 10.205 15.385 10.495 16.110 ;
        RECT 12.065 15.385 12.305 16.195 ;
        RECT 12.475 15.555 12.805 16.195 ;
        RECT 12.975 15.385 13.245 16.195 ;
        RECT 14.205 16.065 14.580 16.625 ;
        RECT 14.785 16.295 15.095 16.625 ;
        RECT 15.265 16.195 15.445 17.150 ;
        RECT 16.805 16.980 17.065 17.205 ;
        RECT 15.775 16.810 17.065 16.980 ;
        RECT 17.575 16.965 17.905 17.750 ;
        RECT 15.775 16.545 15.945 16.810 ;
        RECT 15.615 16.375 15.945 16.545 ;
        RECT 15.265 16.025 16.245 16.195 ;
        RECT 13.430 15.385 13.685 15.875 ;
        RECT 15.360 15.385 15.745 15.855 ;
        RECT 15.915 15.555 16.245 16.025 ;
        RECT 16.415 15.385 16.625 16.195 ;
        RECT 16.805 15.845 16.985 16.810 ;
        RECT 17.575 16.795 18.255 16.965 ;
        RECT 18.435 16.795 18.765 17.935 ;
        RECT 18.955 16.795 19.285 17.935 ;
        RECT 19.815 17.255 20.145 17.750 ;
        RECT 19.815 17.085 20.555 17.255 ;
        RECT 19.815 16.965 20.145 17.085 ;
        RECT 19.465 16.795 20.145 16.965 ;
        RECT 17.155 16.025 17.380 16.625 ;
        RECT 17.565 16.375 17.915 16.625 ;
        RECT 18.085 16.195 18.255 16.795 ;
        RECT 18.425 16.575 18.775 16.625 ;
        RECT 18.945 16.575 19.295 16.625 ;
        RECT 18.425 16.405 19.295 16.575 ;
        RECT 18.425 16.375 18.775 16.405 ;
        RECT 18.945 16.375 19.295 16.405 ;
        RECT 19.465 16.195 19.635 16.795 ;
        RECT 19.805 16.375 20.155 16.625 ;
        RECT 20.385 16.575 20.555 17.085 ;
        RECT 23.085 16.770 23.375 17.935 ;
        RECT 23.875 16.980 24.135 17.205 ;
        RECT 24.335 17.155 24.665 17.935 ;
        RECT 25.115 17.150 25.675 17.765 ;
        RECT 23.875 16.810 25.165 16.980 ;
        RECT 25.495 16.915 25.675 17.150 ;
        RECT 25.865 17.135 26.145 17.935 ;
        RECT 26.875 17.135 27.045 17.935 ;
        RECT 23.560 16.575 23.785 16.625 ;
        RECT 20.385 16.405 23.785 16.575 ;
        RECT 16.805 15.670 17.150 15.845 ;
        RECT 17.585 15.385 17.825 16.195 ;
        RECT 17.995 15.555 18.325 16.195 ;
        RECT 18.495 15.385 18.765 16.195 ;
        RECT 18.955 15.385 19.225 16.195 ;
        RECT 19.395 15.555 19.725 16.195 ;
        RECT 19.895 15.385 20.135 16.195 ;
        RECT 23.085 15.385 23.375 16.110 ;
        RECT 23.560 16.025 23.785 16.405 ;
        RECT 23.955 15.845 24.135 16.810 ;
        RECT 24.995 16.545 25.165 16.810 ;
        RECT 25.445 16.745 25.675 16.915 ;
        RECT 27.715 16.795 27.975 17.935 ;
        RECT 28.655 17.135 28.885 17.935 ;
        RECT 29.555 16.795 29.810 17.935 ;
        RECT 29.985 16.795 30.265 17.935 ;
        RECT 30.935 16.795 31.195 17.935 ;
        RECT 24.995 16.375 25.325 16.545 ;
        RECT 25.495 16.195 25.675 16.745 ;
        RECT 27.085 16.295 27.465 16.625 ;
        RECT 28.145 16.295 28.455 16.625 ;
        RECT 23.790 15.670 24.135 15.845 ;
        RECT 24.315 15.385 24.525 16.195 ;
        RECT 24.695 16.025 25.675 16.195 ;
        RECT 24.695 15.555 25.025 16.025 ;
        RECT 25.195 15.385 25.580 15.855 ;
        RECT 27.250 15.600 27.465 16.295 ;
        RECT 27.635 15.385 27.970 16.125 ;
        RECT 29.570 16.045 29.790 16.625 ;
        RECT 29.995 16.355 30.330 16.625 ;
        RECT 30.840 16.575 31.175 16.625 ;
        RECT 31.885 16.575 32.055 21.845 ;
        RECT 30.840 16.405 32.055 16.575 ;
        RECT 30.840 16.375 31.175 16.405 ;
        RECT 29.555 15.385 29.810 15.875 ;
        RECT 29.985 15.385 30.295 16.185 ;
        RECT 10.120 15.215 31.280 15.385 ;
        RECT 10.670 14.475 11.005 15.215 ;
        RECT 11.580 14.475 11.930 15.000 ;
        RECT 13.430 14.725 13.685 15.215 ;
        RECT 11.725 14.305 11.930 14.475 ;
        RECT 10.690 14.195 10.975 14.305 ;
        RECT 9.345 14.025 10.975 14.195 ;
        RECT 10.690 13.975 10.975 14.025 ;
        RECT 11.725 13.975 12.035 14.305 ;
        RECT 13.450 13.975 13.670 14.555 ;
        RECT 15.275 14.405 15.545 15.215 ;
        RECT 15.715 14.405 16.045 15.045 ;
        RECT 16.215 14.405 16.455 15.215 ;
        RECT 16.645 14.490 16.935 15.215 ;
        RECT 17.995 14.540 18.320 15.045 ;
        RECT 18.490 14.710 18.775 15.215 ;
        RECT 14.785 13.975 15.095 14.305 ;
        RECT 15.785 13.805 15.955 14.405 ;
        RECT 16.125 13.975 16.475 14.225 ;
        RECT 17.995 14.010 18.775 14.540 ;
        RECT 18.955 14.405 19.225 15.215 ;
        RECT 19.395 14.405 19.725 15.045 ;
        RECT 19.895 14.405 20.135 15.215 ;
        RECT 20.570 14.755 20.915 14.930 ;
        RECT 10.665 12.665 10.925 13.805 ;
        RECT 11.595 12.665 11.765 13.465 ;
        RECT 12.495 12.665 12.775 13.465 ;
        RECT 13.430 12.665 13.685 13.805 ;
        RECT 14.355 12.665 14.585 13.465 ;
        RECT 15.275 12.665 15.605 13.805 ;
        RECT 15.785 13.635 16.465 13.805 ;
        RECT 16.135 12.850 16.465 13.635 ;
        RECT 16.645 12.665 16.935 13.830 ;
        RECT 17.565 12.665 17.825 13.635 ;
        RECT 17.995 12.835 18.325 14.010 ;
        RECT 19.465 13.805 19.635 14.405 ;
        RECT 19.805 13.975 20.155 14.225 ;
        RECT 20.340 13.975 20.565 14.575 ;
        RECT 18.495 12.665 18.775 13.635 ;
        RECT 18.955 12.665 19.285 13.805 ;
        RECT 19.465 13.635 20.145 13.805 ;
        RECT 20.735 13.790 20.915 14.755 ;
        RECT 21.095 14.405 21.305 15.215 ;
        RECT 21.475 14.575 21.805 15.045 ;
        RECT 21.975 14.745 22.360 15.215 ;
        RECT 21.475 14.405 22.455 14.575 ;
        RECT 21.775 14.055 22.105 14.225 ;
        RECT 21.775 13.790 21.945 14.055 ;
        RECT 19.815 12.850 20.145 13.635 ;
        RECT 20.655 13.620 21.945 13.790 ;
        RECT 20.655 13.395 20.915 13.620 ;
        RECT 22.275 13.450 22.455 14.405 ;
        RECT 23.055 14.540 23.380 15.045 ;
        RECT 23.550 14.710 23.835 15.215 ;
        RECT 23.055 14.010 23.835 14.540 ;
        RECT 24.870 14.475 25.220 15.000 ;
        RECT 25.795 14.475 26.130 15.215 ;
        RECT 24.870 14.305 25.075 14.475 ;
        RECT 26.775 14.405 27.045 15.215 ;
        RECT 27.215 14.405 27.545 15.045 ;
        RECT 27.715 14.405 27.955 15.215 ;
        RECT 28.145 14.415 28.455 15.215 ;
        RECT 29.525 14.490 29.815 15.215 ;
        RECT 21.115 12.665 21.445 13.445 ;
        RECT 21.895 12.835 22.455 13.450 ;
        RECT 22.625 12.665 22.885 13.635 ;
        RECT 23.055 12.835 23.385 14.010 ;
        RECT 24.765 13.975 25.075 14.305 ;
        RECT 25.825 13.975 26.110 14.305 ;
        RECT 27.285 13.805 27.455 14.405 ;
        RECT 27.625 13.975 27.975 14.225 ;
        RECT 28.155 13.975 28.490 14.245 ;
        RECT 29.000 13.975 29.335 14.225 ;
        RECT 23.555 12.665 23.835 13.635 ;
        RECT 24.025 12.665 24.305 13.465 ;
        RECT 25.035 12.665 25.205 13.465 ;
        RECT 25.875 12.665 26.135 13.805 ;
        RECT 26.775 12.665 27.105 13.805 ;
        RECT 27.285 13.635 27.965 13.805 ;
        RECT 27.635 12.850 27.965 13.635 ;
        RECT 28.145 12.665 28.425 13.805 ;
        RECT 29.095 12.665 29.355 13.805 ;
        RECT 29.525 12.665 29.815 13.830 ;
        RECT 10.120 12.495 31.280 12.665 ;
        RECT 10.205 11.330 10.495 12.495 ;
        RECT 10.665 11.355 10.925 12.495 ;
        RECT 11.595 11.695 11.765 12.495 ;
        RECT 12.495 11.695 12.775 12.495 ;
        RECT 15.265 11.355 15.545 12.495 ;
        RECT 15.715 11.345 16.045 12.325 ;
        RECT 16.215 11.355 16.475 12.495 ;
        RECT 11.175 10.855 11.555 11.185 ;
        RECT 10.205 9.945 10.495 10.670 ;
        RECT 10.670 9.945 11.005 10.685 ;
        RECT 11.175 10.160 11.390 10.855 ;
        RECT 15.780 10.745 15.950 11.345 ;
        RECT 16.645 11.330 16.935 12.495 ;
        RECT 18.520 11.695 18.770 12.495 ;
        RECT 18.940 11.865 19.270 12.325 ;
        RECT 19.440 12.035 19.655 12.495 ;
        RECT 18.940 11.695 20.110 11.865 ;
        RECT 18.030 11.525 18.310 11.685 ;
        RECT 18.030 11.355 19.365 11.525 ;
        RECT 19.195 11.185 19.365 11.355 ;
        RECT 19.195 10.935 19.570 11.185 ;
        RECT 19.195 10.765 19.365 10.935 ;
        RECT 15.265 9.945 15.575 10.745 ;
        RECT 15.780 10.115 16.475 10.745 ;
        RECT 16.645 9.945 16.935 10.670 ;
        RECT 18.030 10.595 19.365 10.765 ;
        RECT 18.030 10.385 18.300 10.595 ;
        RECT 19.740 10.405 20.110 11.695 ;
        RECT 20.335 11.355 20.665 12.495 ;
        RECT 21.195 11.525 21.525 12.310 ;
        RECT 20.845 11.355 21.525 11.525 ;
        RECT 21.705 11.355 21.965 12.495 ;
        RECT 22.635 11.355 22.915 12.495 ;
        RECT 20.845 10.755 21.015 11.355 ;
        RECT 23.085 11.330 23.375 12.495 ;
        RECT 24.515 11.695 24.745 12.495 ;
        RECT 25.415 11.355 25.670 12.495 ;
        RECT 26.355 11.695 26.585 12.495 ;
        RECT 27.255 11.355 27.510 12.495 ;
        RECT 28.195 11.695 28.425 12.495 ;
        RECT 29.095 11.355 29.350 12.495 ;
        RECT 29.525 11.330 29.815 12.495 ;
        RECT 21.725 10.935 22.060 11.185 ;
        RECT 22.570 10.915 22.905 11.185 ;
        RECT 24.005 11.135 24.315 11.185 ;
        RECT 23.605 10.965 24.315 11.135 ;
        RECT 18.520 9.945 18.850 10.405 ;
        RECT 19.360 10.115 20.110 10.405 ;
        RECT 20.335 9.945 20.605 10.755 ;
        RECT 20.775 10.115 21.105 10.755 ;
        RECT 21.275 9.945 21.515 10.755 ;
        RECT 22.605 9.945 22.915 10.745 ;
        RECT 23.085 9.945 23.375 10.670 ;
        RECT 23.605 10.625 23.775 10.965 ;
        RECT 24.005 10.855 24.315 10.965 ;
        RECT 24.520 10.625 24.895 11.185 ;
        RECT 26.360 10.625 26.735 11.185 ;
        RECT 27.270 10.605 27.490 11.185 ;
        RECT 29.110 10.605 29.330 11.185 ;
        RECT 25.415 9.945 25.670 10.435 ;
        RECT 27.255 9.945 27.510 10.435 ;
        RECT 29.095 9.945 29.350 10.435 ;
        RECT 29.525 9.945 29.815 10.670 ;
        RECT 10.120 9.775 31.280 9.945 ;
      LAYER mcon ;
        RECT 10.265 26.095 10.435 26.265 ;
        RECT 10.725 26.095 10.895 26.265 ;
        RECT 11.185 26.095 11.355 26.265 ;
        RECT 11.645 26.095 11.815 26.265 ;
        RECT 12.105 26.095 12.275 26.265 ;
        RECT 12.565 26.095 12.735 26.265 ;
        RECT 13.025 26.095 13.195 26.265 ;
        RECT 13.485 26.095 13.655 26.265 ;
        RECT 13.945 26.095 14.115 26.265 ;
        RECT 14.405 26.095 14.575 26.265 ;
        RECT 14.865 26.095 15.035 26.265 ;
        RECT 15.325 26.095 15.495 26.265 ;
        RECT 15.785 26.095 15.955 26.265 ;
        RECT 16.245 26.095 16.415 26.265 ;
        RECT 16.705 26.095 16.875 26.265 ;
        RECT 17.165 26.095 17.335 26.265 ;
        RECT 17.625 26.095 17.795 26.265 ;
        RECT 18.085 26.095 18.255 26.265 ;
        RECT 18.545 26.095 18.715 26.265 ;
        RECT 19.005 26.095 19.175 26.265 ;
        RECT 19.465 26.095 19.635 26.265 ;
        RECT 19.925 26.095 20.095 26.265 ;
        RECT 20.385 26.095 20.555 26.265 ;
        RECT 20.845 26.095 21.015 26.265 ;
        RECT 21.305 26.095 21.475 26.265 ;
        RECT 21.765 26.095 21.935 26.265 ;
        RECT 22.225 26.095 22.395 26.265 ;
        RECT 22.685 26.095 22.855 26.265 ;
        RECT 23.145 26.095 23.315 26.265 ;
        RECT 23.605 26.095 23.775 26.265 ;
        RECT 24.065 26.095 24.235 26.265 ;
        RECT 24.525 26.095 24.695 26.265 ;
        RECT 24.985 26.095 25.155 26.265 ;
        RECT 25.445 26.095 25.615 26.265 ;
        RECT 25.905 26.095 26.075 26.265 ;
        RECT 26.365 26.095 26.535 26.265 ;
        RECT 26.825 26.095 26.995 26.265 ;
        RECT 27.285 26.095 27.455 26.265 ;
        RECT 27.745 26.095 27.915 26.265 ;
        RECT 28.205 26.095 28.375 26.265 ;
        RECT 28.665 26.095 28.835 26.265 ;
        RECT 29.125 26.095 29.295 26.265 ;
        RECT 29.585 26.095 29.755 26.265 ;
        RECT 30.045 26.095 30.215 26.265 ;
        RECT 30.505 26.095 30.675 26.265 ;
        RECT 30.965 26.095 31.135 26.265 ;
        RECT 13.945 25.585 14.115 25.755 ;
        RECT 12.105 24.905 12.275 25.075 ;
        RECT 15.785 24.905 15.955 25.075 ;
        RECT 25.905 25.245 26.075 25.415 ;
        RECT 19.465 24.565 19.635 24.735 ;
        RECT 26.825 25.245 26.995 25.415 ;
        RECT 28.665 24.905 28.835 25.075 ;
        RECT 10.265 23.375 10.435 23.545 ;
        RECT 10.725 23.375 10.895 23.545 ;
        RECT 11.185 23.375 11.355 23.545 ;
        RECT 11.645 23.375 11.815 23.545 ;
        RECT 12.105 23.375 12.275 23.545 ;
        RECT 12.565 23.375 12.735 23.545 ;
        RECT 13.025 23.375 13.195 23.545 ;
        RECT 13.485 23.375 13.655 23.545 ;
        RECT 13.945 23.375 14.115 23.545 ;
        RECT 14.405 23.375 14.575 23.545 ;
        RECT 14.865 23.375 15.035 23.545 ;
        RECT 15.325 23.375 15.495 23.545 ;
        RECT 15.785 23.375 15.955 23.545 ;
        RECT 16.245 23.375 16.415 23.545 ;
        RECT 16.705 23.375 16.875 23.545 ;
        RECT 17.165 23.375 17.335 23.545 ;
        RECT 17.625 23.375 17.795 23.545 ;
        RECT 18.085 23.375 18.255 23.545 ;
        RECT 18.545 23.375 18.715 23.545 ;
        RECT 19.005 23.375 19.175 23.545 ;
        RECT 19.465 23.375 19.635 23.545 ;
        RECT 19.925 23.375 20.095 23.545 ;
        RECT 20.385 23.375 20.555 23.545 ;
        RECT 20.845 23.375 21.015 23.545 ;
        RECT 21.305 23.375 21.475 23.545 ;
        RECT 21.765 23.375 21.935 23.545 ;
        RECT 22.225 23.375 22.395 23.545 ;
        RECT 22.685 23.375 22.855 23.545 ;
        RECT 23.145 23.375 23.315 23.545 ;
        RECT 23.605 23.375 23.775 23.545 ;
        RECT 24.065 23.375 24.235 23.545 ;
        RECT 24.525 23.375 24.695 23.545 ;
        RECT 24.985 23.375 25.155 23.545 ;
        RECT 25.445 23.375 25.615 23.545 ;
        RECT 25.905 23.375 26.075 23.545 ;
        RECT 26.365 23.375 26.535 23.545 ;
        RECT 26.825 23.375 26.995 23.545 ;
        RECT 27.285 23.375 27.455 23.545 ;
        RECT 27.745 23.375 27.915 23.545 ;
        RECT 28.205 23.375 28.375 23.545 ;
        RECT 28.665 23.375 28.835 23.545 ;
        RECT 29.125 23.375 29.295 23.545 ;
        RECT 29.585 23.375 29.755 23.545 ;
        RECT 30.045 23.375 30.215 23.545 ;
        RECT 30.505 23.375 30.675 23.545 ;
        RECT 30.965 23.375 31.135 23.545 ;
        RECT 15.325 22.185 15.495 22.355 ;
        RECT 12.565 21.845 12.735 22.015 ;
        RECT 13.485 21.845 13.655 22.015 ;
        RECT 14.865 21.845 15.035 22.015 ;
        RECT 11.645 21.505 11.815 21.675 ;
        RECT 17.165 21.505 17.335 21.675 ;
        RECT 24.525 22.525 24.695 22.695 ;
        RECT 19.005 21.505 19.175 21.675 ;
        RECT 19.925 21.505 20.095 21.675 ;
        RECT 21.765 21.845 21.935 22.015 ;
        RECT 22.685 21.845 22.855 22.015 ;
        RECT 20.845 21.505 21.015 21.675 ;
        RECT 24.525 21.845 24.695 22.015 ;
        RECT 28.665 21.505 28.835 21.675 ;
        RECT 30.045 21.845 30.215 22.015 ;
        RECT 25.905 21.165 26.075 21.335 ;
        RECT 10.265 20.655 10.435 20.825 ;
        RECT 10.725 20.655 10.895 20.825 ;
        RECT 11.185 20.655 11.355 20.825 ;
        RECT 11.645 20.655 11.815 20.825 ;
        RECT 12.105 20.655 12.275 20.825 ;
        RECT 12.565 20.655 12.735 20.825 ;
        RECT 13.025 20.655 13.195 20.825 ;
        RECT 13.485 20.655 13.655 20.825 ;
        RECT 13.945 20.655 14.115 20.825 ;
        RECT 14.405 20.655 14.575 20.825 ;
        RECT 14.865 20.655 15.035 20.825 ;
        RECT 15.325 20.655 15.495 20.825 ;
        RECT 15.785 20.655 15.955 20.825 ;
        RECT 16.245 20.655 16.415 20.825 ;
        RECT 16.705 20.655 16.875 20.825 ;
        RECT 17.165 20.655 17.335 20.825 ;
        RECT 17.625 20.655 17.795 20.825 ;
        RECT 18.085 20.655 18.255 20.825 ;
        RECT 18.545 20.655 18.715 20.825 ;
        RECT 19.005 20.655 19.175 20.825 ;
        RECT 19.465 20.655 19.635 20.825 ;
        RECT 19.925 20.655 20.095 20.825 ;
        RECT 20.385 20.655 20.555 20.825 ;
        RECT 20.845 20.655 21.015 20.825 ;
        RECT 21.305 20.655 21.475 20.825 ;
        RECT 21.765 20.655 21.935 20.825 ;
        RECT 22.225 20.655 22.395 20.825 ;
        RECT 22.685 20.655 22.855 20.825 ;
        RECT 23.145 20.655 23.315 20.825 ;
        RECT 23.605 20.655 23.775 20.825 ;
        RECT 24.065 20.655 24.235 20.825 ;
        RECT 24.525 20.655 24.695 20.825 ;
        RECT 24.985 20.655 25.155 20.825 ;
        RECT 25.445 20.655 25.615 20.825 ;
        RECT 25.905 20.655 26.075 20.825 ;
        RECT 26.365 20.655 26.535 20.825 ;
        RECT 26.825 20.655 26.995 20.825 ;
        RECT 27.285 20.655 27.455 20.825 ;
        RECT 27.745 20.655 27.915 20.825 ;
        RECT 28.205 20.655 28.375 20.825 ;
        RECT 28.665 20.655 28.835 20.825 ;
        RECT 29.125 20.655 29.295 20.825 ;
        RECT 29.585 20.655 29.755 20.825 ;
        RECT 30.045 20.655 30.215 20.825 ;
        RECT 30.505 20.655 30.675 20.825 ;
        RECT 30.965 20.655 31.135 20.825 ;
        RECT 11.645 19.805 11.815 19.975 ;
        RECT 14.865 20.145 15.035 20.315 ;
        RECT 18.085 20.145 18.255 20.315 ;
        RECT 19.005 19.465 19.175 19.635 ;
        RECT 19.925 19.465 20.095 19.635 ;
        RECT 20.845 19.805 21.015 19.975 ;
        RECT 24.525 20.145 24.695 20.315 ;
        RECT 25.905 19.805 26.075 19.975 ;
        RECT 28.205 19.465 28.375 19.635 ;
        RECT 29.125 19.465 29.295 19.635 ;
        RECT 27.745 18.445 27.915 18.615 ;
        RECT 31.885 18.445 32.055 18.615 ;
        RECT 10.265 17.935 10.435 18.105 ;
        RECT 10.725 17.935 10.895 18.105 ;
        RECT 11.185 17.935 11.355 18.105 ;
        RECT 11.645 17.935 11.815 18.105 ;
        RECT 12.105 17.935 12.275 18.105 ;
        RECT 12.565 17.935 12.735 18.105 ;
        RECT 13.025 17.935 13.195 18.105 ;
        RECT 13.485 17.935 13.655 18.105 ;
        RECT 13.945 17.935 14.115 18.105 ;
        RECT 14.405 17.935 14.575 18.105 ;
        RECT 14.865 17.935 15.035 18.105 ;
        RECT 15.325 17.935 15.495 18.105 ;
        RECT 15.785 17.935 15.955 18.105 ;
        RECT 16.245 17.935 16.415 18.105 ;
        RECT 16.705 17.935 16.875 18.105 ;
        RECT 17.165 17.935 17.335 18.105 ;
        RECT 17.625 17.935 17.795 18.105 ;
        RECT 18.085 17.935 18.255 18.105 ;
        RECT 18.545 17.935 18.715 18.105 ;
        RECT 19.005 17.935 19.175 18.105 ;
        RECT 19.465 17.935 19.635 18.105 ;
        RECT 19.925 17.935 20.095 18.105 ;
        RECT 20.385 17.935 20.555 18.105 ;
        RECT 20.845 17.935 21.015 18.105 ;
        RECT 21.305 17.935 21.475 18.105 ;
        RECT 21.765 17.935 21.935 18.105 ;
        RECT 22.225 17.935 22.395 18.105 ;
        RECT 22.685 17.935 22.855 18.105 ;
        RECT 23.145 17.935 23.315 18.105 ;
        RECT 23.605 17.935 23.775 18.105 ;
        RECT 24.065 17.935 24.235 18.105 ;
        RECT 24.525 17.935 24.695 18.105 ;
        RECT 24.985 17.935 25.155 18.105 ;
        RECT 25.445 17.935 25.615 18.105 ;
        RECT 25.905 17.935 26.075 18.105 ;
        RECT 26.365 17.935 26.535 18.105 ;
        RECT 26.825 17.935 26.995 18.105 ;
        RECT 27.285 17.935 27.455 18.105 ;
        RECT 27.745 17.935 27.915 18.105 ;
        RECT 28.205 17.935 28.375 18.105 ;
        RECT 28.665 17.935 28.835 18.105 ;
        RECT 29.125 17.935 29.295 18.105 ;
        RECT 29.585 17.935 29.755 18.105 ;
        RECT 30.045 17.935 30.215 18.105 ;
        RECT 30.505 17.935 30.675 18.105 ;
        RECT 30.965 17.935 31.135 18.105 ;
        RECT 15.325 17.425 15.495 17.595 ;
        RECT 14.865 16.405 15.035 16.575 ;
        RECT 12.565 15.725 12.735 15.895 ;
        RECT 14.405 16.065 14.575 16.235 ;
        RECT 17.625 16.405 17.795 16.575 ;
        RECT 17.165 16.065 17.335 16.235 ;
        RECT 18.545 16.405 18.715 16.575 ;
        RECT 18.085 16.065 18.255 16.235 ;
        RECT 19.925 16.405 20.095 16.575 ;
        RECT 23.605 16.405 23.775 16.575 ;
        RECT 28.205 16.405 28.375 16.575 ;
        RECT 27.285 16.065 27.455 16.235 ;
        RECT 30.045 16.405 30.215 16.575 ;
        RECT 29.585 16.065 29.755 16.235 ;
        RECT 10.265 15.215 10.435 15.385 ;
        RECT 10.725 15.215 10.895 15.385 ;
        RECT 11.185 15.215 11.355 15.385 ;
        RECT 11.645 15.215 11.815 15.385 ;
        RECT 12.105 15.215 12.275 15.385 ;
        RECT 12.565 15.215 12.735 15.385 ;
        RECT 13.025 15.215 13.195 15.385 ;
        RECT 13.485 15.215 13.655 15.385 ;
        RECT 13.945 15.215 14.115 15.385 ;
        RECT 14.405 15.215 14.575 15.385 ;
        RECT 14.865 15.215 15.035 15.385 ;
        RECT 15.325 15.215 15.495 15.385 ;
        RECT 15.785 15.215 15.955 15.385 ;
        RECT 16.245 15.215 16.415 15.385 ;
        RECT 16.705 15.215 16.875 15.385 ;
        RECT 17.165 15.215 17.335 15.385 ;
        RECT 17.625 15.215 17.795 15.385 ;
        RECT 18.085 15.215 18.255 15.385 ;
        RECT 18.545 15.215 18.715 15.385 ;
        RECT 19.005 15.215 19.175 15.385 ;
        RECT 19.465 15.215 19.635 15.385 ;
        RECT 19.925 15.215 20.095 15.385 ;
        RECT 20.385 15.215 20.555 15.385 ;
        RECT 20.845 15.215 21.015 15.385 ;
        RECT 21.305 15.215 21.475 15.385 ;
        RECT 21.765 15.215 21.935 15.385 ;
        RECT 22.225 15.215 22.395 15.385 ;
        RECT 22.685 15.215 22.855 15.385 ;
        RECT 23.145 15.215 23.315 15.385 ;
        RECT 23.605 15.215 23.775 15.385 ;
        RECT 24.065 15.215 24.235 15.385 ;
        RECT 24.525 15.215 24.695 15.385 ;
        RECT 24.985 15.215 25.155 15.385 ;
        RECT 25.445 15.215 25.615 15.385 ;
        RECT 25.905 15.215 26.075 15.385 ;
        RECT 26.365 15.215 26.535 15.385 ;
        RECT 26.825 15.215 26.995 15.385 ;
        RECT 27.285 15.215 27.455 15.385 ;
        RECT 27.745 15.215 27.915 15.385 ;
        RECT 28.205 15.215 28.375 15.385 ;
        RECT 28.665 15.215 28.835 15.385 ;
        RECT 29.125 15.215 29.295 15.385 ;
        RECT 29.585 15.215 29.755 15.385 ;
        RECT 30.045 15.215 30.215 15.385 ;
        RECT 30.505 15.215 30.675 15.385 ;
        RECT 30.965 15.215 31.135 15.385 ;
        RECT 11.645 14.705 11.815 14.875 ;
        RECT 13.485 14.365 13.655 14.535 ;
        RECT 15.785 14.705 15.955 14.875 ;
        RECT 18.085 14.705 18.255 14.875 ;
        RECT 14.865 14.025 15.035 14.195 ;
        RECT 16.245 14.025 16.415 14.195 ;
        RECT 19.465 14.705 19.635 14.875 ;
        RECT 20.385 14.365 20.555 14.535 ;
        RECT 19.925 14.025 20.095 14.195 ;
        RECT 24.985 14.705 25.155 14.875 ;
        RECT 27.285 14.365 27.455 14.535 ;
        RECT 23.605 14.025 23.775 14.195 ;
        RECT 22.225 13.005 22.395 13.175 ;
        RECT 25.905 14.025 26.075 14.195 ;
        RECT 27.745 14.025 27.915 14.195 ;
        RECT 28.205 14.025 28.375 14.195 ;
        RECT 29.125 14.025 29.295 14.195 ;
        RECT 10.265 12.495 10.435 12.665 ;
        RECT 10.725 12.495 10.895 12.665 ;
        RECT 11.185 12.495 11.355 12.665 ;
        RECT 11.645 12.495 11.815 12.665 ;
        RECT 12.105 12.495 12.275 12.665 ;
        RECT 12.565 12.495 12.735 12.665 ;
        RECT 13.025 12.495 13.195 12.665 ;
        RECT 13.485 12.495 13.655 12.665 ;
        RECT 13.945 12.495 14.115 12.665 ;
        RECT 14.405 12.495 14.575 12.665 ;
        RECT 14.865 12.495 15.035 12.665 ;
        RECT 15.325 12.495 15.495 12.665 ;
        RECT 15.785 12.495 15.955 12.665 ;
        RECT 16.245 12.495 16.415 12.665 ;
        RECT 16.705 12.495 16.875 12.665 ;
        RECT 17.165 12.495 17.335 12.665 ;
        RECT 17.625 12.495 17.795 12.665 ;
        RECT 18.085 12.495 18.255 12.665 ;
        RECT 18.545 12.495 18.715 12.665 ;
        RECT 19.005 12.495 19.175 12.665 ;
        RECT 19.465 12.495 19.635 12.665 ;
        RECT 19.925 12.495 20.095 12.665 ;
        RECT 20.385 12.495 20.555 12.665 ;
        RECT 20.845 12.495 21.015 12.665 ;
        RECT 21.305 12.495 21.475 12.665 ;
        RECT 21.765 12.495 21.935 12.665 ;
        RECT 22.225 12.495 22.395 12.665 ;
        RECT 22.685 12.495 22.855 12.665 ;
        RECT 23.145 12.495 23.315 12.665 ;
        RECT 23.605 12.495 23.775 12.665 ;
        RECT 24.065 12.495 24.235 12.665 ;
        RECT 24.525 12.495 24.695 12.665 ;
        RECT 24.985 12.495 25.155 12.665 ;
        RECT 25.445 12.495 25.615 12.665 ;
        RECT 25.905 12.495 26.075 12.665 ;
        RECT 26.365 12.495 26.535 12.665 ;
        RECT 26.825 12.495 26.995 12.665 ;
        RECT 27.285 12.495 27.455 12.665 ;
        RECT 27.745 12.495 27.915 12.665 ;
        RECT 28.205 12.495 28.375 12.665 ;
        RECT 28.665 12.495 28.835 12.665 ;
        RECT 29.125 12.495 29.295 12.665 ;
        RECT 29.585 12.495 29.755 12.665 ;
        RECT 30.045 12.495 30.215 12.665 ;
        RECT 30.505 12.495 30.675 12.665 ;
        RECT 30.965 12.495 31.135 12.665 ;
        RECT 15.785 11.985 15.955 12.155 ;
        RECT 11.185 10.965 11.355 11.135 ;
        RECT 19.005 11.985 19.175 12.155 ;
        RECT 21.765 10.965 21.935 11.135 ;
        RECT 22.685 10.965 22.855 11.135 ;
        RECT 20.845 10.625 21.015 10.795 ;
        RECT 24.525 10.625 24.695 10.795 ;
        RECT 26.365 10.625 26.535 10.795 ;
        RECT 27.285 10.965 27.455 11.135 ;
        RECT 29.125 10.625 29.295 10.795 ;
        RECT 10.265 9.775 10.435 9.945 ;
        RECT 10.725 9.775 10.895 9.945 ;
        RECT 11.185 9.775 11.355 9.945 ;
        RECT 11.645 9.775 11.815 9.945 ;
        RECT 12.105 9.775 12.275 9.945 ;
        RECT 12.565 9.775 12.735 9.945 ;
        RECT 13.025 9.775 13.195 9.945 ;
        RECT 13.485 9.775 13.655 9.945 ;
        RECT 13.945 9.775 14.115 9.945 ;
        RECT 14.405 9.775 14.575 9.945 ;
        RECT 14.865 9.775 15.035 9.945 ;
        RECT 15.325 9.775 15.495 9.945 ;
        RECT 15.785 9.775 15.955 9.945 ;
        RECT 16.245 9.775 16.415 9.945 ;
        RECT 16.705 9.775 16.875 9.945 ;
        RECT 17.165 9.775 17.335 9.945 ;
        RECT 17.625 9.775 17.795 9.945 ;
        RECT 18.085 9.775 18.255 9.945 ;
        RECT 18.545 9.775 18.715 9.945 ;
        RECT 19.005 9.775 19.175 9.945 ;
        RECT 19.465 9.775 19.635 9.945 ;
        RECT 19.925 9.775 20.095 9.945 ;
        RECT 20.385 9.775 20.555 9.945 ;
        RECT 20.845 9.775 21.015 9.945 ;
        RECT 21.305 9.775 21.475 9.945 ;
        RECT 21.765 9.775 21.935 9.945 ;
        RECT 22.225 9.775 22.395 9.945 ;
        RECT 22.685 9.775 22.855 9.945 ;
        RECT 23.145 9.775 23.315 9.945 ;
        RECT 23.605 9.775 23.775 9.945 ;
        RECT 24.065 9.775 24.235 9.945 ;
        RECT 24.525 9.775 24.695 9.945 ;
        RECT 24.985 9.775 25.155 9.945 ;
        RECT 25.445 9.775 25.615 9.945 ;
        RECT 25.905 9.775 26.075 9.945 ;
        RECT 26.365 9.775 26.535 9.945 ;
        RECT 26.825 9.775 26.995 9.945 ;
        RECT 27.285 9.775 27.455 9.945 ;
        RECT 27.745 9.775 27.915 9.945 ;
        RECT 28.205 9.775 28.375 9.945 ;
        RECT 28.665 9.775 28.835 9.945 ;
        RECT 29.125 9.775 29.295 9.945 ;
        RECT 29.585 9.775 29.755 9.945 ;
        RECT 30.045 9.775 30.215 9.945 ;
        RECT 30.505 9.775 30.675 9.945 ;
        RECT 30.965 9.775 31.135 9.945 ;
      LAYER met1 ;
        RECT 2.120 25.940 39.280 26.420 ;
        RECT 13.870 25.540 14.190 25.800 ;
        RECT 25.845 25.400 26.135 25.445 ;
        RECT 26.765 25.400 27.055 25.445 ;
        RECT 25.845 25.260 30.200 25.400 ;
        RECT 25.845 25.215 26.135 25.260 ;
        RECT 26.765 25.215 27.055 25.260 ;
        RECT 30.060 25.120 30.200 25.260 ;
        RECT 12.045 25.060 12.335 25.105 ;
        RECT 15.725 25.060 16.015 25.105 ;
        RECT 12.045 24.920 13.180 25.060 ;
        RECT 12.045 24.875 12.335 24.920 ;
        RECT 13.040 24.380 13.180 24.920 ;
        RECT 14.880 24.920 16.015 25.060 ;
        RECT 13.870 24.720 14.190 24.780 ;
        RECT 14.880 24.720 15.020 24.920 ;
        RECT 15.725 24.875 16.015 24.920 ;
        RECT 28.130 25.060 28.450 25.120 ;
        RECT 28.605 25.060 28.895 25.105 ;
        RECT 28.130 24.920 28.895 25.060 ;
        RECT 28.130 24.860 28.450 24.920 ;
        RECT 28.605 24.875 28.895 24.920 ;
        RECT 29.970 24.860 30.290 25.120 ;
        RECT 15.250 24.720 15.570 24.780 ;
        RECT 13.870 24.580 15.570 24.720 ;
        RECT 13.870 24.520 14.190 24.580 ;
        RECT 15.250 24.520 15.570 24.580 ;
        RECT 19.405 24.720 19.695 24.765 ;
        RECT 20.785 24.720 21.075 24.765 ;
        RECT 19.405 24.580 21.075 24.720 ;
        RECT 19.405 24.535 19.695 24.580 ;
        RECT 20.785 24.535 21.075 24.580 ;
        RECT 22.610 24.380 22.930 24.440 ;
        RECT 13.040 24.240 19.160 24.380 ;
        RECT 19.020 24.210 19.160 24.240 ;
        RECT 21.780 24.240 22.930 24.380 ;
        RECT 21.780 24.210 21.920 24.240 ;
        RECT 19.020 24.070 21.920 24.210 ;
        RECT 22.610 24.180 22.930 24.240 ;
        RECT 6.120 23.220 35.280 23.700 ;
        RECT 24.465 22.680 24.755 22.725 ;
        RECT 28.130 22.680 28.450 22.740 ;
        RECT 24.465 22.540 28.450 22.680 ;
        RECT 24.465 22.495 24.755 22.540 ;
        RECT 28.130 22.480 28.450 22.540 ;
        RECT 15.250 22.340 15.570 22.400 ;
        RECT 14.975 22.200 15.570 22.340 ;
        RECT 15.250 22.140 15.570 22.200 ;
        RECT 19.020 22.200 21.920 22.340 ;
        RECT 12.490 22.000 12.810 22.060 ;
        RECT 12.490 21.860 13.085 22.000 ;
        RECT 12.490 21.800 12.810 21.860 ;
        RECT 13.425 21.815 13.715 22.045 ;
        RECT 14.330 22.000 14.650 22.060 ;
        RECT 14.805 22.000 15.095 22.045 ;
        RECT 14.330 21.860 15.095 22.000 ;
        RECT 11.570 21.660 11.890 21.720 ;
        RECT 13.500 21.660 13.640 21.815 ;
        RECT 14.330 21.800 14.650 21.860 ;
        RECT 14.805 21.815 15.095 21.860 ;
        RECT 19.020 21.705 19.160 22.200 ;
        RECT 21.780 22.045 21.920 22.200 ;
        RECT 21.705 21.815 21.995 22.045 ;
        RECT 22.610 22.000 22.930 22.060 ;
        RECT 24.450 22.000 24.770 22.060 ;
        RECT 29.970 22.000 30.290 22.060 ;
        RECT 22.240 21.860 22.930 22.000 ;
        RECT 24.175 21.860 24.770 22.000 ;
        RECT 29.695 21.860 30.290 22.000 ;
        RECT 11.570 21.520 13.640 21.660 ;
        RECT 17.105 21.660 17.395 21.705 ;
        RECT 18.945 21.660 19.235 21.705 ;
        RECT 19.850 21.660 20.170 21.720 ;
        RECT 17.105 21.520 19.235 21.660 ;
        RECT 19.575 21.520 20.170 21.660 ;
        RECT 11.570 21.460 11.890 21.520 ;
        RECT 17.105 21.475 17.395 21.520 ;
        RECT 18.945 21.475 19.235 21.520 ;
        RECT 19.850 21.460 20.170 21.520 ;
        RECT 20.785 21.660 21.075 21.705 ;
        RECT 22.240 21.660 22.380 21.860 ;
        RECT 22.610 21.800 22.930 21.860 ;
        RECT 24.450 21.800 24.770 21.860 ;
        RECT 29.970 21.800 30.290 21.860 ;
        RECT 28.590 21.660 28.910 21.720 ;
        RECT 20.785 21.520 22.380 21.660 ;
        RECT 28.315 21.520 28.910 21.660 ;
        RECT 20.785 21.475 21.075 21.520 ;
        RECT 28.590 21.460 28.910 21.520 ;
        RECT 23.530 21.320 23.850 21.380 ;
        RECT 25.830 21.320 26.150 21.380 ;
        RECT 23.530 21.180 26.150 21.320 ;
        RECT 23.530 21.120 23.850 21.180 ;
        RECT 25.830 21.120 26.150 21.180 ;
        RECT 2.120 20.500 39.280 20.980 ;
        RECT 14.330 20.300 14.650 20.360 ;
        RECT 14.805 20.300 15.095 20.345 ;
        RECT 14.330 20.160 15.095 20.300 ;
        RECT 14.330 20.100 14.650 20.160 ;
        RECT 14.805 20.115 15.095 20.160 ;
        RECT 15.250 20.300 15.570 20.360 ;
        RECT 18.025 20.300 18.315 20.345 ;
        RECT 24.450 20.300 24.770 20.360 ;
        RECT 15.250 20.160 20.080 20.300 ;
        RECT 24.175 20.160 24.770 20.300 ;
        RECT 15.250 20.100 15.570 20.160 ;
        RECT 18.025 20.115 18.315 20.160 ;
        RECT 11.570 19.960 11.890 20.020 ;
        RECT 11.295 19.820 11.890 19.960 ;
        RECT 19.940 19.960 20.080 20.160 ;
        RECT 24.450 20.100 24.770 20.160 ;
        RECT 28.130 20.100 28.450 20.360 ;
        RECT 20.785 19.960 21.075 20.005 ;
        RECT 19.940 19.820 21.075 19.960 ;
        RECT 11.570 19.760 11.890 19.820 ;
        RECT 20.785 19.775 21.075 19.820 ;
        RECT 25.370 19.960 25.690 20.020 ;
        RECT 25.845 19.960 26.135 20.005 ;
        RECT 25.370 19.820 26.135 19.960 ;
        RECT 25.370 19.760 25.690 19.820 ;
        RECT 25.845 19.775 26.135 19.820 ;
        RECT 18.945 19.620 19.235 19.665 ;
        RECT 19.850 19.620 20.170 19.680 ;
        RECT 28.220 19.665 28.360 20.100 ;
        RECT 18.945 19.480 20.170 19.620 ;
        RECT 18.945 19.435 19.235 19.480 ;
        RECT 19.850 19.420 20.170 19.480 ;
        RECT 28.145 19.435 28.435 19.665 ;
        RECT 29.050 19.620 29.370 19.680 ;
        RECT 28.775 19.480 29.370 19.620 ;
        RECT 29.050 19.420 29.370 19.480 ;
        RECT 22.610 19.280 22.930 19.340 ;
        RECT 22.610 19.140 23.205 19.280 ;
        RECT 22.610 19.080 22.930 19.140 ;
        RECT 27.685 18.600 27.975 18.645 ;
        RECT 31.825 18.600 32.115 18.645 ;
        RECT 27.685 18.460 32.115 18.600 ;
        RECT 27.685 18.415 27.975 18.460 ;
        RECT 31.825 18.415 32.115 18.460 ;
        RECT 6.120 17.780 35.280 18.260 ;
        RECT 11.570 17.580 11.890 17.640 ;
        RECT 15.265 17.580 15.555 17.625 ;
        RECT 11.570 17.440 15.555 17.580 ;
        RECT 11.570 17.380 11.890 17.440 ;
        RECT 15.265 17.395 15.555 17.440 ;
        RECT 25.370 16.900 25.690 16.960 ;
        RECT 25.370 16.760 30.200 16.900 ;
        RECT 25.370 16.700 25.690 16.760 ;
        RECT 14.790 16.560 15.110 16.620 ;
        RECT 17.550 16.560 17.870 16.620 ;
        RECT 18.470 16.560 18.790 16.620 ;
        RECT 19.850 16.560 20.170 16.620 ;
        RECT 23.530 16.560 23.850 16.620 ;
        RECT 30.060 16.605 30.200 16.760 ;
        RECT 14.515 16.420 15.110 16.560 ;
        RECT 17.275 16.420 17.870 16.560 ;
        RECT 18.195 16.420 18.790 16.560 ;
        RECT 19.575 16.420 20.170 16.560 ;
        RECT 23.255 16.420 23.850 16.560 ;
        RECT 14.790 16.360 15.110 16.420 ;
        RECT 17.550 16.360 17.870 16.420 ;
        RECT 18.470 16.360 18.790 16.420 ;
        RECT 19.850 16.360 20.170 16.420 ;
        RECT 23.530 16.360 23.850 16.420 ;
        RECT 28.145 16.375 28.435 16.605 ;
        RECT 29.985 16.375 30.275 16.605 ;
        RECT 13.870 16.220 14.190 16.280 ;
        RECT 14.345 16.220 14.635 16.265 ;
        RECT 17.105 16.220 17.395 16.265 ;
        RECT 18.025 16.220 18.315 16.265 ;
        RECT 27.225 16.220 27.515 16.265 ;
        RECT 28.220 16.220 28.360 16.375 ;
        RECT 13.870 16.080 18.315 16.220 ;
        RECT 13.870 16.020 14.190 16.080 ;
        RECT 14.345 16.035 14.635 16.080 ;
        RECT 17.105 16.035 17.395 16.080 ;
        RECT 18.025 16.035 18.315 16.080 ;
        RECT 25.460 16.080 28.360 16.220 ;
        RECT 29.050 16.220 29.370 16.280 ;
        RECT 29.525 16.220 29.815 16.265 ;
        RECT 29.050 16.080 29.815 16.220 ;
        RECT 12.030 15.880 12.350 15.940 ;
        RECT 12.505 15.880 12.795 15.925 ;
        RECT 12.030 15.740 12.795 15.880 ;
        RECT 12.030 15.680 12.350 15.740 ;
        RECT 12.505 15.695 12.795 15.740 ;
        RECT 24.450 15.880 24.770 15.940 ;
        RECT 25.460 15.880 25.600 16.080 ;
        RECT 27.225 16.035 27.515 16.080 ;
        RECT 29.050 16.020 29.370 16.080 ;
        RECT 29.525 16.035 29.815 16.080 ;
        RECT 24.450 15.740 25.600 15.880 ;
        RECT 24.450 15.680 24.770 15.740 ;
        RECT 2.120 15.060 39.280 15.540 ;
        RECT 11.570 14.860 11.890 14.920 ;
        RECT 15.710 14.860 16.030 14.920 ;
        RECT 11.295 14.720 11.890 14.860 ;
        RECT 15.435 14.720 16.030 14.860 ;
        RECT 11.570 14.660 11.890 14.720 ;
        RECT 15.710 14.660 16.030 14.720 ;
        RECT 18.025 14.860 18.315 14.905 ;
        RECT 18.470 14.860 18.790 14.920 ;
        RECT 18.025 14.720 18.790 14.860 ;
        RECT 18.025 14.675 18.315 14.720 ;
        RECT 18.470 14.660 18.790 14.720 ;
        RECT 19.405 14.860 19.695 14.905 ;
        RECT 24.450 14.860 24.770 14.920 ;
        RECT 24.925 14.860 25.215 14.905 ;
        RECT 19.405 14.720 25.215 14.860 ;
        RECT 19.405 14.675 19.695 14.720 ;
        RECT 12.030 14.520 12.350 14.580 ;
        RECT 20.400 14.565 20.540 14.720 ;
        RECT 24.450 14.660 24.770 14.720 ;
        RECT 24.925 14.675 25.215 14.720 ;
        RECT 29.050 14.660 29.370 14.920 ;
        RECT 13.425 14.520 13.715 14.565 ;
        RECT 12.030 14.380 13.715 14.520 ;
        RECT 12.030 14.320 12.350 14.380 ;
        RECT 13.425 14.335 13.715 14.380 ;
        RECT 20.325 14.335 20.615 14.565 ;
        RECT 27.225 14.520 27.515 14.565 ;
        RECT 29.140 14.520 29.280 14.660 ;
        RECT 27.225 14.380 29.280 14.520 ;
        RECT 27.225 14.335 27.515 14.380 ;
        RECT 11.570 14.180 11.890 14.240 ;
        RECT 13.870 14.180 14.190 14.240 ;
        RECT 14.805 14.180 15.095 14.225 ;
        RECT 16.170 14.180 16.490 14.240 ;
        RECT 19.850 14.180 20.170 14.240 ;
        RECT 28.220 14.225 28.360 14.380 ;
        RECT 11.570 14.040 15.095 14.180 ;
        RECT 15.895 14.040 16.490 14.180 ;
        RECT 19.575 14.040 20.170 14.180 ;
        RECT 11.570 13.980 11.890 14.040 ;
        RECT 13.870 13.980 14.190 14.040 ;
        RECT 14.805 13.995 15.095 14.040 ;
        RECT 16.170 13.980 16.490 14.040 ;
        RECT 19.850 13.980 20.170 14.040 ;
        RECT 23.545 14.180 23.835 14.225 ;
        RECT 25.845 14.180 26.135 14.225 ;
        RECT 23.545 14.040 26.520 14.180 ;
        RECT 23.545 13.995 23.835 14.040 ;
        RECT 25.845 13.995 26.135 14.040 ;
        RECT 26.380 13.840 26.520 14.040 ;
        RECT 27.685 13.995 27.975 14.225 ;
        RECT 28.145 13.995 28.435 14.225 ;
        RECT 29.050 14.180 29.370 14.240 ;
        RECT 28.775 14.040 29.370 14.180 ;
        RECT 27.210 13.840 27.530 13.900 ;
        RECT 27.760 13.840 27.900 13.995 ;
        RECT 29.050 13.980 29.370 14.040 ;
        RECT 26.380 13.700 27.900 13.840 ;
        RECT 27.210 13.640 27.530 13.700 ;
        RECT 22.165 13.160 22.455 13.205 ;
        RECT 22.610 13.160 22.930 13.220 ;
        RECT 22.165 13.020 22.930 13.160 ;
        RECT 22.165 12.975 22.455 13.020 ;
        RECT 22.610 12.960 22.930 13.020 ;
        RECT 6.120 12.340 35.280 12.820 ;
        RECT 15.725 12.140 16.015 12.185 ;
        RECT 16.170 12.140 16.490 12.200 ;
        RECT 15.725 12.000 16.490 12.140 ;
        RECT 15.725 11.955 16.015 12.000 ;
        RECT 16.170 11.940 16.490 12.000 ;
        RECT 18.945 12.140 19.235 12.185 ;
        RECT 19.850 12.140 20.170 12.200 ;
        RECT 18.945 12.000 20.170 12.140 ;
        RECT 18.945 11.955 19.235 12.000 ;
        RECT 19.850 11.940 20.170 12.000 ;
        RECT 11.125 11.120 11.415 11.165 ;
        RECT 11.570 11.120 11.890 11.180 ;
        RECT 11.125 10.980 11.890 11.120 ;
        RECT 11.125 10.935 11.415 10.980 ;
        RECT 11.570 10.920 11.890 10.980 ;
        RECT 21.705 10.935 21.995 11.165 ;
        RECT 22.610 11.120 22.930 11.180 ;
        RECT 27.210 11.120 27.530 11.180 ;
        RECT 22.335 10.980 25.140 11.120 ;
        RECT 26.935 10.980 27.530 11.120 ;
        RECT 20.785 10.780 21.075 10.825 ;
        RECT 21.780 10.780 21.920 10.935 ;
        RECT 22.610 10.920 22.930 10.980 ;
        RECT 23.545 10.780 23.835 10.825 ;
        RECT 24.450 10.780 24.770 10.840 ;
        RECT 20.785 10.640 23.835 10.780 ;
        RECT 24.175 10.640 24.770 10.780 ;
        RECT 25.000 10.780 25.140 10.980 ;
        RECT 27.210 10.920 27.530 10.980 ;
        RECT 26.305 10.780 26.595 10.825 ;
        RECT 29.065 10.780 29.355 10.825 ;
        RECT 25.000 10.640 29.355 10.780 ;
        RECT 20.785 10.595 21.075 10.640 ;
        RECT 23.545 10.595 23.835 10.640 ;
        RECT 24.450 10.580 24.770 10.640 ;
        RECT 26.305 10.595 26.595 10.640 ;
        RECT 29.065 10.595 29.355 10.640 ;
        RECT 2.120 9.620 39.280 10.100 ;
      LAYER via ;
        RECT 2.190 26.050 2.450 26.310 ;
        RECT 2.510 26.050 2.770 26.310 ;
        RECT 2.830 26.050 3.090 26.310 ;
        RECT 3.150 26.050 3.410 26.310 ;
        RECT 3.470 26.050 3.730 26.310 ;
        RECT 3.790 26.050 4.050 26.310 ;
        RECT 37.350 26.050 37.610 26.310 ;
        RECT 37.670 26.050 37.930 26.310 ;
        RECT 37.990 26.050 38.250 26.310 ;
        RECT 38.310 26.050 38.570 26.310 ;
        RECT 38.630 26.050 38.890 26.310 ;
        RECT 38.950 26.050 39.210 26.310 ;
        RECT 13.900 25.540 14.160 25.800 ;
        RECT 13.900 24.520 14.160 24.780 ;
        RECT 28.160 24.860 28.420 25.120 ;
        RECT 30.000 24.860 30.260 25.120 ;
        RECT 15.280 24.520 15.540 24.780 ;
        RECT 22.640 24.180 22.900 24.440 ;
        RECT 6.190 23.330 6.450 23.590 ;
        RECT 6.510 23.330 6.770 23.590 ;
        RECT 6.830 23.330 7.090 23.590 ;
        RECT 7.150 23.330 7.410 23.590 ;
        RECT 7.470 23.330 7.730 23.590 ;
        RECT 7.790 23.330 8.050 23.590 ;
        RECT 33.350 23.330 33.610 23.590 ;
        RECT 33.670 23.330 33.930 23.590 ;
        RECT 33.990 23.330 34.250 23.590 ;
        RECT 34.310 23.330 34.570 23.590 ;
        RECT 34.630 23.330 34.890 23.590 ;
        RECT 34.950 23.330 35.210 23.590 ;
        RECT 28.160 22.480 28.420 22.740 ;
        RECT 15.280 22.140 15.540 22.400 ;
        RECT 12.520 21.800 12.780 22.060 ;
        RECT 11.600 21.460 11.860 21.720 ;
        RECT 14.360 21.800 14.620 22.060 ;
        RECT 19.880 21.460 20.140 21.720 ;
        RECT 22.640 21.800 22.900 22.060 ;
        RECT 24.480 21.800 24.740 22.060 ;
        RECT 30.000 21.800 30.260 22.060 ;
        RECT 28.620 21.460 28.880 21.720 ;
        RECT 23.560 21.120 23.820 21.380 ;
        RECT 25.860 21.120 26.120 21.380 ;
        RECT 2.190 20.610 2.450 20.870 ;
        RECT 2.510 20.610 2.770 20.870 ;
        RECT 2.830 20.610 3.090 20.870 ;
        RECT 3.150 20.610 3.410 20.870 ;
        RECT 3.470 20.610 3.730 20.870 ;
        RECT 3.790 20.610 4.050 20.870 ;
        RECT 37.350 20.610 37.610 20.870 ;
        RECT 37.670 20.610 37.930 20.870 ;
        RECT 37.990 20.610 38.250 20.870 ;
        RECT 38.310 20.610 38.570 20.870 ;
        RECT 38.630 20.610 38.890 20.870 ;
        RECT 38.950 20.610 39.210 20.870 ;
        RECT 14.360 20.100 14.620 20.360 ;
        RECT 15.280 20.100 15.540 20.360 ;
        RECT 11.600 19.760 11.860 20.020 ;
        RECT 24.480 20.100 24.740 20.360 ;
        RECT 28.160 20.100 28.420 20.360 ;
        RECT 25.400 19.760 25.660 20.020 ;
        RECT 19.880 19.420 20.140 19.680 ;
        RECT 29.080 19.420 29.340 19.680 ;
        RECT 22.640 19.080 22.900 19.340 ;
        RECT 6.190 17.890 6.450 18.150 ;
        RECT 6.510 17.890 6.770 18.150 ;
        RECT 6.830 17.890 7.090 18.150 ;
        RECT 7.150 17.890 7.410 18.150 ;
        RECT 7.470 17.890 7.730 18.150 ;
        RECT 7.790 17.890 8.050 18.150 ;
        RECT 33.350 17.890 33.610 18.150 ;
        RECT 33.670 17.890 33.930 18.150 ;
        RECT 33.990 17.890 34.250 18.150 ;
        RECT 34.310 17.890 34.570 18.150 ;
        RECT 34.630 17.890 34.890 18.150 ;
        RECT 34.950 17.890 35.210 18.150 ;
        RECT 11.600 17.380 11.860 17.640 ;
        RECT 25.400 16.700 25.660 16.960 ;
        RECT 14.820 16.360 15.080 16.620 ;
        RECT 17.580 16.360 17.840 16.620 ;
        RECT 18.500 16.360 18.760 16.620 ;
        RECT 19.880 16.360 20.140 16.620 ;
        RECT 23.560 16.360 23.820 16.620 ;
        RECT 13.900 16.020 14.160 16.280 ;
        RECT 12.060 15.680 12.320 15.940 ;
        RECT 24.480 15.680 24.740 15.940 ;
        RECT 29.080 16.020 29.340 16.280 ;
        RECT 2.190 15.170 2.450 15.430 ;
        RECT 2.510 15.170 2.770 15.430 ;
        RECT 2.830 15.170 3.090 15.430 ;
        RECT 3.150 15.170 3.410 15.430 ;
        RECT 3.470 15.170 3.730 15.430 ;
        RECT 3.790 15.170 4.050 15.430 ;
        RECT 37.350 15.170 37.610 15.430 ;
        RECT 37.670 15.170 37.930 15.430 ;
        RECT 37.990 15.170 38.250 15.430 ;
        RECT 38.310 15.170 38.570 15.430 ;
        RECT 38.630 15.170 38.890 15.430 ;
        RECT 38.950 15.170 39.210 15.430 ;
        RECT 11.600 14.660 11.860 14.920 ;
        RECT 15.740 14.660 16.000 14.920 ;
        RECT 18.500 14.660 18.760 14.920 ;
        RECT 12.060 14.320 12.320 14.580 ;
        RECT 24.480 14.660 24.740 14.920 ;
        RECT 29.080 14.660 29.340 14.920 ;
        RECT 11.600 13.980 11.860 14.240 ;
        RECT 13.900 13.980 14.160 14.240 ;
        RECT 16.200 13.980 16.460 14.240 ;
        RECT 19.880 13.980 20.140 14.240 ;
        RECT 27.240 13.640 27.500 13.900 ;
        RECT 29.080 13.980 29.340 14.240 ;
        RECT 22.640 12.960 22.900 13.220 ;
        RECT 6.190 12.450 6.450 12.710 ;
        RECT 6.510 12.450 6.770 12.710 ;
        RECT 6.830 12.450 7.090 12.710 ;
        RECT 7.150 12.450 7.410 12.710 ;
        RECT 7.470 12.450 7.730 12.710 ;
        RECT 7.790 12.450 8.050 12.710 ;
        RECT 33.350 12.450 33.610 12.710 ;
        RECT 33.670 12.450 33.930 12.710 ;
        RECT 33.990 12.450 34.250 12.710 ;
        RECT 34.310 12.450 34.570 12.710 ;
        RECT 34.630 12.450 34.890 12.710 ;
        RECT 34.950 12.450 35.210 12.710 ;
        RECT 16.200 11.940 16.460 12.200 ;
        RECT 19.880 11.940 20.140 12.200 ;
        RECT 11.600 10.920 11.860 11.180 ;
        RECT 22.640 10.920 22.900 11.180 ;
        RECT 24.480 10.580 24.740 10.840 ;
        RECT 27.240 10.920 27.500 11.180 ;
        RECT 2.190 9.730 2.450 9.990 ;
        RECT 2.510 9.730 2.770 9.990 ;
        RECT 2.830 9.730 3.090 9.990 ;
        RECT 3.150 9.730 3.410 9.990 ;
        RECT 3.470 9.730 3.730 9.990 ;
        RECT 3.790 9.730 4.050 9.990 ;
        RECT 37.350 9.730 37.610 9.990 ;
        RECT 37.670 9.730 37.930 9.990 ;
        RECT 37.990 9.730 38.250 9.990 ;
        RECT 38.310 9.730 38.570 9.990 ;
        RECT 38.630 9.730 38.890 9.990 ;
        RECT 38.950 9.730 39.210 9.990 ;
      LAYER met2 ;
        RECT 2.120 25.940 4.120 26.420 ;
        RECT 37.280 25.940 39.280 26.420 ;
        RECT 13.900 25.510 14.160 25.830 ;
        RECT 13.960 24.810 14.100 25.510 ;
        RECT 28.160 24.830 28.420 25.150 ;
        RECT 30.000 24.830 30.260 25.150 ;
        RECT 13.900 24.490 14.160 24.810 ;
        RECT 15.280 24.490 15.540 24.810 ;
        RECT 6.120 23.220 8.120 23.700 ;
        RECT 15.340 22.430 15.480 24.490 ;
        RECT 22.640 24.150 22.900 24.470 ;
        RECT 15.280 22.110 15.540 22.430 ;
        RECT 12.520 21.770 12.780 22.090 ;
        RECT 14.360 21.770 14.620 22.090 ;
        RECT 11.600 21.430 11.860 21.750 ;
        RECT 2.120 20.500 4.120 20.980 ;
        RECT 11.660 20.050 11.800 21.430 ;
        RECT 12.580 20.640 12.720 21.770 ;
        RECT 12.350 20.500 12.720 20.640 ;
        RECT 11.600 19.730 11.860 20.050 ;
        RECT 6.120 17.780 8.120 18.260 ;
        RECT 11.660 17.670 11.800 19.730 ;
        RECT 11.600 17.350 11.860 17.670 ;
        RECT 12.350 16.900 12.490 20.500 ;
        RECT 14.420 20.390 14.560 21.770 ;
        RECT 15.340 20.390 15.480 22.110 ;
        RECT 22.700 22.090 22.840 24.150 ;
        RECT 28.220 22.770 28.360 24.830 ;
        RECT 28.160 22.450 28.420 22.770 ;
        RECT 22.640 21.770 22.900 22.090 ;
        RECT 24.480 21.770 24.740 22.090 ;
        RECT 19.880 21.430 20.140 21.750 ;
        RECT 14.360 20.070 14.620 20.390 ;
        RECT 15.280 20.070 15.540 20.390 ;
        RECT 14.420 17.240 14.560 20.070 ;
        RECT 14.420 17.100 15.020 17.240 ;
        RECT 12.120 16.760 12.490 16.900 ;
        RECT 12.120 15.970 12.260 16.760 ;
        RECT 14.880 16.650 15.020 17.100 ;
        RECT 14.820 16.330 15.080 16.650 ;
        RECT 15.340 16.560 15.480 20.070 ;
        RECT 19.940 19.710 20.080 21.430 ;
        RECT 19.880 19.390 20.140 19.710 ;
        RECT 22.700 19.370 22.840 21.770 ;
        RECT 23.560 21.090 23.820 21.410 ;
        RECT 22.640 19.050 22.900 19.370 ;
        RECT 23.620 16.650 23.760 21.090 ;
        RECT 24.540 20.390 24.680 21.770 ;
        RECT 25.850 21.090 26.130 21.805 ;
        RECT 28.220 20.390 28.360 22.450 ;
        RECT 30.060 22.090 30.200 24.830 ;
        RECT 33.280 23.220 35.280 23.700 ;
        RECT 30.000 21.805 30.260 22.090 ;
        RECT 28.620 21.430 28.880 21.750 ;
        RECT 29.990 21.435 30.270 21.805 ;
        RECT 28.680 20.640 28.820 21.430 ;
        RECT 28.680 20.500 29.280 20.640 ;
        RECT 37.280 20.500 39.280 20.980 ;
        RECT 24.480 20.070 24.740 20.390 ;
        RECT 28.160 20.070 28.420 20.390 ;
        RECT 25.400 19.975 25.660 20.050 ;
        RECT 29.140 19.975 29.280 20.500 ;
        RECT 25.390 19.605 25.670 19.975 ;
        RECT 29.070 19.605 29.350 19.975 ;
        RECT 25.460 16.990 25.600 19.605 ;
        RECT 29.080 19.390 29.340 19.605 ;
        RECT 33.280 17.780 35.280 18.260 ;
        RECT 25.400 16.670 25.660 16.990 ;
        RECT 15.340 16.420 15.940 16.560 ;
        RECT 13.900 15.990 14.160 16.310 ;
        RECT 12.060 15.650 12.320 15.970 ;
        RECT 2.120 15.060 4.120 15.540 ;
        RECT 11.600 14.630 11.860 14.950 ;
        RECT 11.660 14.270 11.800 14.630 ;
        RECT 12.120 14.610 12.260 15.650 ;
        RECT 12.060 14.290 12.320 14.610 ;
        RECT 13.960 14.270 14.100 15.990 ;
        RECT 15.800 14.950 15.940 16.420 ;
        RECT 17.580 16.330 17.840 16.650 ;
        RECT 18.500 16.330 18.760 16.650 ;
        RECT 19.880 16.330 20.140 16.650 ;
        RECT 23.560 16.330 23.820 16.650 ;
        RECT 15.740 14.630 16.000 14.950 ;
        RECT 17.640 14.485 17.780 16.330 ;
        RECT 18.560 14.950 18.700 16.330 ;
        RECT 18.500 14.630 18.760 14.950 ;
        RECT 11.600 13.950 11.860 14.270 ;
        RECT 13.900 13.950 14.160 14.270 ;
        RECT 16.190 14.115 16.470 14.485 ;
        RECT 17.570 14.115 17.850 14.485 ;
        RECT 19.940 14.270 20.080 16.330 ;
        RECT 29.080 15.990 29.340 16.310 ;
        RECT 24.480 15.650 24.740 15.970 ;
        RECT 24.540 14.950 24.680 15.650 ;
        RECT 29.140 14.950 29.280 15.990 ;
        RECT 37.280 15.060 39.280 15.540 ;
        RECT 24.480 14.630 24.740 14.950 ;
        RECT 29.080 14.630 29.340 14.950 ;
        RECT 16.200 13.950 16.460 14.115 ;
        RECT 19.880 13.950 20.140 14.270 ;
        RECT 6.120 12.340 8.120 12.820 ;
        RECT 11.660 11.210 11.800 13.950 ;
        RECT 16.260 12.230 16.400 13.950 ;
        RECT 19.940 12.230 20.080 13.950 ;
        RECT 22.630 13.505 22.910 13.875 ;
        RECT 22.700 13.250 22.840 13.505 ;
        RECT 22.640 12.930 22.900 13.250 ;
        RECT 16.200 11.910 16.460 12.230 ;
        RECT 19.880 11.910 20.140 12.230 ;
        RECT 22.700 11.210 22.840 12.930 ;
        RECT 11.600 10.890 11.860 11.210 ;
        RECT 22.640 10.890 22.900 11.210 ;
        RECT 24.540 10.870 24.680 14.630 ;
        RECT 27.240 13.610 27.500 13.930 ;
        RECT 27.300 11.210 27.440 13.610 ;
        RECT 29.070 13.505 29.350 14.270 ;
        RECT 33.280 12.340 35.280 12.820 ;
        RECT 27.240 10.890 27.500 11.210 ;
        RECT 24.480 10.550 24.740 10.870 ;
        RECT 2.120 9.620 4.120 10.100 ;
        RECT 37.280 9.620 39.280 10.100 ;
      LAYER via2 ;
        RECT 2.180 26.040 2.460 26.320 ;
        RECT 2.580 26.040 2.860 26.320 ;
        RECT 2.980 26.040 3.260 26.320 ;
        RECT 3.380 26.040 3.660 26.320 ;
        RECT 3.780 26.040 4.060 26.320 ;
        RECT 37.340 26.040 37.620 26.320 ;
        RECT 37.740 26.040 38.020 26.320 ;
        RECT 38.140 26.040 38.420 26.320 ;
        RECT 38.540 26.040 38.820 26.320 ;
        RECT 38.940 26.040 39.220 26.320 ;
        RECT 6.180 23.320 6.460 23.600 ;
        RECT 6.580 23.320 6.860 23.600 ;
        RECT 6.980 23.320 7.260 23.600 ;
        RECT 7.380 23.320 7.660 23.600 ;
        RECT 7.780 23.320 8.060 23.600 ;
        RECT 2.180 20.600 2.460 20.880 ;
        RECT 2.580 20.600 2.860 20.880 ;
        RECT 2.980 20.600 3.260 20.880 ;
        RECT 3.380 20.600 3.660 20.880 ;
        RECT 3.780 20.600 4.060 20.880 ;
        RECT 6.180 17.880 6.460 18.160 ;
        RECT 6.580 17.880 6.860 18.160 ;
        RECT 6.980 17.880 7.260 18.160 ;
        RECT 7.380 17.880 7.660 18.160 ;
        RECT 7.780 17.880 8.060 18.160 ;
        RECT 25.850 21.480 26.130 21.760 ;
        RECT 33.340 23.320 33.620 23.600 ;
        RECT 33.740 23.320 34.020 23.600 ;
        RECT 34.140 23.320 34.420 23.600 ;
        RECT 34.540 23.320 34.820 23.600 ;
        RECT 34.940 23.320 35.220 23.600 ;
        RECT 29.990 21.480 30.270 21.760 ;
        RECT 37.340 20.600 37.620 20.880 ;
        RECT 37.740 20.600 38.020 20.880 ;
        RECT 38.140 20.600 38.420 20.880 ;
        RECT 38.540 20.600 38.820 20.880 ;
        RECT 38.940 20.600 39.220 20.880 ;
        RECT 25.390 19.650 25.670 19.930 ;
        RECT 29.070 19.650 29.350 19.930 ;
        RECT 33.340 17.880 33.620 18.160 ;
        RECT 33.740 17.880 34.020 18.160 ;
        RECT 34.140 17.880 34.420 18.160 ;
        RECT 34.540 17.880 34.820 18.160 ;
        RECT 34.940 17.880 35.220 18.160 ;
        RECT 2.180 15.160 2.460 15.440 ;
        RECT 2.580 15.160 2.860 15.440 ;
        RECT 2.980 15.160 3.260 15.440 ;
        RECT 3.380 15.160 3.660 15.440 ;
        RECT 3.780 15.160 4.060 15.440 ;
        RECT 16.190 14.160 16.470 14.440 ;
        RECT 17.570 14.160 17.850 14.440 ;
        RECT 37.340 15.160 37.620 15.440 ;
        RECT 37.740 15.160 38.020 15.440 ;
        RECT 38.140 15.160 38.420 15.440 ;
        RECT 38.540 15.160 38.820 15.440 ;
        RECT 38.940 15.160 39.220 15.440 ;
        RECT 6.180 12.440 6.460 12.720 ;
        RECT 6.580 12.440 6.860 12.720 ;
        RECT 6.980 12.440 7.260 12.720 ;
        RECT 7.380 12.440 7.660 12.720 ;
        RECT 7.780 12.440 8.060 12.720 ;
        RECT 22.630 13.550 22.910 13.830 ;
        RECT 29.070 13.550 29.350 13.830 ;
        RECT 33.340 12.440 33.620 12.720 ;
        RECT 33.740 12.440 34.020 12.720 ;
        RECT 34.140 12.440 34.420 12.720 ;
        RECT 34.540 12.440 34.820 12.720 ;
        RECT 34.940 12.440 35.220 12.720 ;
        RECT 2.180 9.720 2.460 10.000 ;
        RECT 2.580 9.720 2.860 10.000 ;
        RECT 2.980 9.720 3.260 10.000 ;
        RECT 3.380 9.720 3.660 10.000 ;
        RECT 3.780 9.720 4.060 10.000 ;
        RECT 37.340 9.720 37.620 10.000 ;
        RECT 37.740 9.720 38.020 10.000 ;
        RECT 38.140 9.720 38.420 10.000 ;
        RECT 38.540 9.720 38.820 10.000 ;
        RECT 38.940 9.720 39.220 10.000 ;
      LAYER met3 ;
        RECT 2.120 25.940 4.120 26.420 ;
        RECT 37.280 25.940 39.280 26.420 ;
        RECT 6.120 23.220 8.120 23.700 ;
        RECT 33.280 23.220 35.280 23.700 ;
        RECT 25.825 21.770 26.155 21.785 ;
        RECT 29.965 21.770 30.295 21.785 ;
        RECT 25.825 21.470 30.295 21.770 ;
        RECT 25.825 21.455 26.155 21.470 ;
        RECT 29.965 21.455 30.295 21.470 ;
        RECT 2.120 20.500 4.120 20.980 ;
        RECT 37.280 20.500 39.280 20.980 ;
        RECT 25.365 19.940 25.695 19.955 ;
        RECT 29.045 19.940 29.375 19.955 ;
        RECT 25.365 19.640 29.375 19.940 ;
        RECT 25.365 19.625 25.695 19.640 ;
        RECT 29.045 19.625 29.375 19.640 ;
        RECT 6.120 17.780 8.120 18.260 ;
        RECT 33.280 17.780 35.280 18.260 ;
        RECT 2.120 15.060 4.120 15.540 ;
        RECT 37.280 15.060 39.280 15.540 ;
        RECT 16.165 14.450 16.495 14.465 ;
        RECT 17.545 14.450 17.875 14.465 ;
        RECT 16.165 14.150 17.875 14.450 ;
        RECT 16.165 14.135 16.495 14.150 ;
        RECT 17.545 14.135 17.875 14.150 ;
        RECT 22.605 13.840 22.935 13.855 ;
        RECT 29.045 13.840 29.375 13.855 ;
        RECT 22.605 13.540 29.375 13.840 ;
        RECT 22.605 13.525 22.935 13.540 ;
        RECT 29.045 13.525 29.375 13.540 ;
        RECT 6.120 12.340 8.120 12.820 ;
        RECT 33.280 12.340 35.280 12.820 ;
        RECT 2.120 9.620 4.120 10.100 ;
        RECT 37.280 9.620 39.280 10.100 ;
      LAYER via3 ;
        RECT 2.160 26.020 2.480 26.340 ;
        RECT 2.560 26.020 2.880 26.340 ;
        RECT 2.960 26.020 3.280 26.340 ;
        RECT 3.360 26.020 3.680 26.340 ;
        RECT 3.760 26.020 4.080 26.340 ;
        RECT 37.320 26.020 37.640 26.340 ;
        RECT 37.720 26.020 38.040 26.340 ;
        RECT 38.120 26.020 38.440 26.340 ;
        RECT 38.520 26.020 38.840 26.340 ;
        RECT 38.920 26.020 39.240 26.340 ;
        RECT 6.160 23.300 6.480 23.620 ;
        RECT 6.560 23.300 6.880 23.620 ;
        RECT 6.960 23.300 7.280 23.620 ;
        RECT 7.360 23.300 7.680 23.620 ;
        RECT 7.760 23.300 8.080 23.620 ;
        RECT 33.320 23.300 33.640 23.620 ;
        RECT 33.720 23.300 34.040 23.620 ;
        RECT 34.120 23.300 34.440 23.620 ;
        RECT 34.520 23.300 34.840 23.620 ;
        RECT 34.920 23.300 35.240 23.620 ;
        RECT 2.160 20.580 2.480 20.900 ;
        RECT 2.560 20.580 2.880 20.900 ;
        RECT 2.960 20.580 3.280 20.900 ;
        RECT 3.360 20.580 3.680 20.900 ;
        RECT 3.760 20.580 4.080 20.900 ;
        RECT 37.320 20.580 37.640 20.900 ;
        RECT 37.720 20.580 38.040 20.900 ;
        RECT 38.120 20.580 38.440 20.900 ;
        RECT 38.520 20.580 38.840 20.900 ;
        RECT 38.920 20.580 39.240 20.900 ;
        RECT 6.160 17.860 6.480 18.180 ;
        RECT 6.560 17.860 6.880 18.180 ;
        RECT 6.960 17.860 7.280 18.180 ;
        RECT 7.360 17.860 7.680 18.180 ;
        RECT 7.760 17.860 8.080 18.180 ;
        RECT 33.320 17.860 33.640 18.180 ;
        RECT 33.720 17.860 34.040 18.180 ;
        RECT 34.120 17.860 34.440 18.180 ;
        RECT 34.520 17.860 34.840 18.180 ;
        RECT 34.920 17.860 35.240 18.180 ;
        RECT 2.160 15.140 2.480 15.460 ;
        RECT 2.560 15.140 2.880 15.460 ;
        RECT 2.960 15.140 3.280 15.460 ;
        RECT 3.360 15.140 3.680 15.460 ;
        RECT 3.760 15.140 4.080 15.460 ;
        RECT 37.320 15.140 37.640 15.460 ;
        RECT 37.720 15.140 38.040 15.460 ;
        RECT 38.120 15.140 38.440 15.460 ;
        RECT 38.520 15.140 38.840 15.460 ;
        RECT 38.920 15.140 39.240 15.460 ;
        RECT 6.160 12.420 6.480 12.740 ;
        RECT 6.560 12.420 6.880 12.740 ;
        RECT 6.960 12.420 7.280 12.740 ;
        RECT 7.360 12.420 7.680 12.740 ;
        RECT 7.760 12.420 8.080 12.740 ;
        RECT 33.320 12.420 33.640 12.740 ;
        RECT 33.720 12.420 34.040 12.740 ;
        RECT 34.120 12.420 34.440 12.740 ;
        RECT 34.520 12.420 34.840 12.740 ;
        RECT 34.920 12.420 35.240 12.740 ;
        RECT 2.160 9.700 2.480 10.020 ;
        RECT 2.560 9.700 2.880 10.020 ;
        RECT 2.960 9.700 3.280 10.020 ;
        RECT 3.360 9.700 3.680 10.020 ;
        RECT 3.760 9.700 4.080 10.020 ;
        RECT 37.320 9.700 37.640 10.020 ;
        RECT 37.720 9.700 38.040 10.020 ;
        RECT 38.120 9.700 38.440 10.020 ;
        RECT 38.520 9.700 38.840 10.020 ;
        RECT 38.920 9.700 39.240 10.020 ;
      LAYER met4 ;
        RECT 2.120 0.000 4.120 36.040 ;
        RECT 6.120 0.000 8.120 36.040 ;
        RECT 33.280 0.000 35.280 36.040 ;
        RECT 37.280 0.000 39.280 36.040 ;
      LAYER via4 ;
        RECT 2.530 32.590 3.710 33.770 ;
        RECT 2.530 2.270 3.710 3.450 ;
        RECT 6.530 28.590 7.710 29.770 ;
        RECT 6.530 6.270 7.710 7.450 ;
        RECT 33.690 28.590 34.870 29.770 ;
        RECT 33.690 6.270 34.870 7.450 ;
        RECT 37.690 32.590 38.870 33.770 ;
        RECT 37.690 2.270 38.870 3.450 ;
      LAYER met5 ;
        RECT 0.000 32.180 41.400 34.180 ;
        RECT 0.000 28.180 41.400 30.180 ;
        RECT 0.000 5.860 41.400 7.860 ;
        RECT 0.000 1.860 41.400 3.860 ;
      LAYER li ;
        RECT 2.110 1.890 39.250 34.100 ;
      LAYER m1 ;
        RECT 2.110 1.890 39.250 34.100 ;
      LAYER m2 ;
        RECT 2.110 1.890 39.250 34.100 ;
      LAYER m3 ;
        RECT 2.110 1.890 39.250 34.100 ;
  END
END decoder5x32
END LIBRARY

