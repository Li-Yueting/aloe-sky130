magic
tech sky130A
magscale 1 2
timestamp 1653197205
<< locali >>
rect 92 1850 262 1910
rect 322 1850 662 1910
rect 722 1850 1062 1910
rect 1122 1850 1462 1910
rect 1522 1850 1862 1910
rect 1922 1850 2262 1910
rect 2322 1850 2662 1910
rect 2722 1850 3062 1910
rect 3122 1850 3462 1910
rect 3522 1850 3862 1910
rect 3922 1850 4262 1910
rect 4322 1850 4662 1910
rect 4722 1850 5062 1910
rect 5122 1850 5462 1910
rect 5522 1850 5862 1910
rect 5922 1850 6262 1910
rect 6322 1850 6662 1910
rect 6722 1850 7062 1910
rect 7122 1850 7260 1910
rect 92 -30 262 30
rect 322 -30 662 30
rect 722 -30 1062 30
rect 1122 -30 1462 30
rect 1522 -30 1862 30
rect 1922 -30 2262 30
rect 2322 -30 2662 30
rect 2722 -30 3062 30
rect 3122 -30 3462 30
rect 3522 -30 3862 30
rect 3922 -30 4262 30
rect 4322 -30 4662 30
rect 4722 -30 5062 30
rect 5122 -30 5462 30
rect 5522 -30 5862 30
rect 5922 -30 6262 30
rect 6322 -30 6662 30
rect 6722 -30 7062 30
rect 7122 -30 7260 30
<< viali >>
rect 262 1850 322 1910
rect 662 1850 722 1910
rect 1062 1850 1122 1910
rect 1462 1850 1522 1910
rect 1862 1850 1922 1910
rect 2262 1850 2322 1910
rect 2662 1850 2722 1910
rect 3062 1850 3122 1910
rect 3462 1850 3522 1910
rect 3862 1850 3922 1910
rect 4262 1850 4322 1910
rect 4662 1850 4722 1910
rect 5062 1850 5122 1910
rect 5462 1850 5522 1910
rect 5862 1850 5922 1910
rect 6262 1850 6322 1910
rect 6662 1850 6722 1910
rect 7062 1850 7122 1910
rect 262 -30 322 30
rect 662 -30 722 30
rect 1062 -30 1122 30
rect 1462 -30 1522 30
rect 1862 -30 1922 30
rect 2262 -30 2322 30
rect 2662 -30 2722 30
rect 3062 -30 3122 30
rect 3462 -30 3522 30
rect 3862 -30 3922 30
rect 4262 -30 4322 30
rect 4662 -30 4722 30
rect 5062 -30 5122 30
rect 5462 -30 5522 30
rect 5862 -30 5922 30
rect 6262 -30 6322 30
rect 6662 -30 6722 30
rect 7062 -30 7122 30
<< metal1 >>
rect 92 1910 7260 1940
rect 92 1850 262 1910
rect 322 1850 662 1910
rect 722 1850 1062 1910
rect 1122 1850 1462 1910
rect 1522 1850 1862 1910
rect 1922 1850 2262 1910
rect 2322 1850 2662 1910
rect 2722 1850 3062 1910
rect 3122 1850 3462 1910
rect 3522 1850 3862 1910
rect 3922 1850 4262 1910
rect 4322 1850 4662 1910
rect 4722 1850 5062 1910
rect 5122 1850 5462 1910
rect 5522 1850 5862 1910
rect 5922 1850 6262 1910
rect 6322 1850 6662 1910
rect 6722 1850 7062 1910
rect 7122 1850 7260 1910
rect 92 1820 7260 1850
rect 92 30 7260 60
rect 92 -30 262 30
rect 322 -30 662 30
rect 722 -30 1062 30
rect 1122 -30 1462 30
rect 1522 -30 1862 30
rect 1922 -30 2262 30
rect 2322 -30 2662 30
rect 2722 -30 3062 30
rect 3122 -30 3462 30
rect 3522 -30 3862 30
rect 3922 -30 4262 30
rect 4322 -30 4662 30
rect 4722 -30 5062 30
rect 5122 -30 5462 30
rect 5522 -30 5862 30
rect 5922 -30 6262 30
rect 6322 -30 6662 30
rect 6722 -30 7062 30
rect 7122 -30 7260 30
rect 92 -60 7260 -30
<< metal2 >>
rect 90 1640 290 1650
rect 90 1580 110 1640
rect 270 1580 290 1640
rect 90 1570 290 1580
rect 112 250 272 260
rect 112 170 132 250
rect 252 170 272 250
rect 112 160 272 170
<< via2 >>
rect 110 1580 270 1640
rect 132 170 252 250
<< metal3 >>
rect 90 1640 7262 1650
rect 90 1580 110 1640
rect 270 1622 7262 1640
rect 270 1580 706 1622
rect 90 1078 706 1580
rect 770 1078 1425 1622
rect 1489 1078 2144 1622
rect 2208 1078 2863 1622
rect 2927 1078 3582 1622
rect 3646 1078 4301 1622
rect 4365 1078 5020 1622
rect 5084 1078 5739 1622
rect 5803 1078 6458 1622
rect 6522 1078 7177 1622
rect 7241 1078 7262 1622
rect 90 922 7262 1078
rect 90 378 706 922
rect 770 378 1425 922
rect 1489 378 2144 922
rect 2208 378 2863 922
rect 2927 378 3582 922
rect 3646 378 4301 922
rect 4365 378 5020 922
rect 5084 378 5739 922
rect 5803 378 6458 922
rect 6522 378 7177 922
rect 7241 378 7262 922
rect 90 350 7262 378
rect 92 260 292 270
rect 92 160 112 260
rect 272 160 292 260
rect 92 150 292 160
<< via3 >>
rect 706 1078 770 1622
rect 1425 1078 1489 1622
rect 2144 1078 2208 1622
rect 2863 1078 2927 1622
rect 3582 1078 3646 1622
rect 4301 1078 4365 1622
rect 5020 1078 5084 1622
rect 5739 1078 5803 1622
rect 6458 1078 6522 1622
rect 7177 1078 7241 1622
rect 706 378 770 922
rect 1425 378 1489 922
rect 2144 378 2208 922
rect 2863 378 2927 922
rect 3582 378 3646 922
rect 4301 378 4365 922
rect 5020 378 5084 922
rect 5739 378 5803 922
rect 6458 378 6522 922
rect 7177 378 7241 922
rect 112 250 272 260
rect 112 170 132 250
rect 132 170 252 250
rect 252 170 272 250
rect 112 160 272 170
<< mimcap >>
rect 191 1510 591 1550
rect 191 1190 231 1510
rect 551 1190 591 1510
rect 191 1150 591 1190
rect 910 1510 1310 1550
rect 910 1190 950 1510
rect 1270 1190 1310 1510
rect 910 1150 1310 1190
rect 1629 1510 2029 1550
rect 1629 1190 1669 1510
rect 1989 1190 2029 1510
rect 1629 1150 2029 1190
rect 2348 1510 2748 1550
rect 2348 1190 2388 1510
rect 2708 1190 2748 1510
rect 2348 1150 2748 1190
rect 3067 1510 3467 1550
rect 3067 1190 3107 1510
rect 3427 1190 3467 1510
rect 3067 1150 3467 1190
rect 3786 1510 4186 1550
rect 3786 1190 3826 1510
rect 4146 1190 4186 1510
rect 3786 1150 4186 1190
rect 4505 1510 4905 1550
rect 4505 1190 4545 1510
rect 4865 1190 4905 1510
rect 4505 1150 4905 1190
rect 5224 1510 5624 1550
rect 5224 1190 5264 1510
rect 5584 1190 5624 1510
rect 5224 1150 5624 1190
rect 5943 1510 6343 1550
rect 5943 1190 5983 1510
rect 6303 1190 6343 1510
rect 5943 1150 6343 1190
rect 6662 1510 7062 1550
rect 6662 1190 6702 1510
rect 7022 1190 7062 1510
rect 6662 1150 7062 1190
rect 191 810 591 850
rect 191 490 231 810
rect 551 490 591 810
rect 191 450 591 490
rect 910 810 1310 850
rect 910 490 950 810
rect 1270 490 1310 810
rect 910 450 1310 490
rect 1629 810 2029 850
rect 1629 490 1669 810
rect 1989 490 2029 810
rect 1629 450 2029 490
rect 2348 810 2748 850
rect 2348 490 2388 810
rect 2708 490 2748 810
rect 2348 450 2748 490
rect 3067 810 3467 850
rect 3067 490 3107 810
rect 3427 490 3467 810
rect 3067 450 3467 490
rect 3786 810 4186 850
rect 3786 490 3826 810
rect 4146 490 4186 810
rect 3786 450 4186 490
rect 4505 810 4905 850
rect 4505 490 4545 810
rect 4865 490 4905 810
rect 4505 450 4905 490
rect 5224 810 5624 850
rect 5224 490 5264 810
rect 5584 490 5624 810
rect 5224 450 5624 490
rect 5943 810 6343 850
rect 5943 490 5983 810
rect 6303 490 6343 810
rect 5943 450 6343 490
rect 6662 810 7062 850
rect 6662 490 6702 810
rect 7022 490 7062 810
rect 6662 450 7062 490
<< mimcapcontact >>
rect 231 1190 551 1510
rect 950 1190 1270 1510
rect 1669 1190 1989 1510
rect 2388 1190 2708 1510
rect 3107 1190 3427 1510
rect 3826 1190 4146 1510
rect 4545 1190 4865 1510
rect 5264 1190 5584 1510
rect 5983 1190 6303 1510
rect 6702 1190 7022 1510
rect 231 490 551 810
rect 950 490 1270 810
rect 1669 490 1989 810
rect 2388 490 2708 810
rect 3107 490 3427 810
rect 3826 490 4146 810
rect 4545 490 4865 810
rect 5264 490 5584 810
rect 5983 490 6303 810
rect 6702 490 7022 810
<< metal4 >>
rect 690 1622 786 1638
rect 230 1511 550 1530
rect 230 1510 552 1511
rect 230 1190 231 1510
rect 551 1190 552 1510
rect 230 1189 552 1190
rect 230 811 550 1189
rect 690 1078 706 1622
rect 770 1078 786 1622
rect 1409 1622 1505 1638
rect 950 1511 1270 1530
rect 949 1510 1271 1511
rect 949 1190 950 1510
rect 1270 1190 1271 1510
rect 949 1189 1271 1190
rect 690 1062 786 1078
rect 690 922 786 938
rect 230 810 552 811
rect 230 490 231 810
rect 551 490 552 810
rect 230 489 552 490
rect 230 290 550 489
rect 690 378 706 922
rect 770 378 786 922
rect 950 811 1270 1189
rect 1409 1078 1425 1622
rect 1489 1078 1505 1622
rect 2128 1622 2224 1638
rect 1670 1511 1990 1530
rect 1668 1510 1990 1511
rect 1668 1190 1669 1510
rect 1989 1190 1990 1510
rect 1668 1189 1990 1190
rect 1409 1062 1505 1078
rect 1409 922 1505 938
rect 949 810 1271 811
rect 949 490 950 810
rect 1270 490 1271 810
rect 949 489 1271 490
rect 690 362 786 378
rect 950 290 1270 489
rect 1409 378 1425 922
rect 1489 378 1505 922
rect 1670 811 1990 1189
rect 2128 1078 2144 1622
rect 2208 1078 2224 1622
rect 2847 1622 2943 1638
rect 2390 1511 2710 1530
rect 2387 1510 2710 1511
rect 2387 1190 2388 1510
rect 2708 1190 2710 1510
rect 2387 1189 2710 1190
rect 2128 1062 2224 1078
rect 1668 810 1990 811
rect 1668 490 1669 810
rect 1989 490 1990 810
rect 1668 489 1990 490
rect 1409 362 1505 378
rect 1670 290 1990 489
rect 2128 922 2224 938
rect 2128 378 2144 922
rect 2208 378 2224 922
rect 2390 811 2710 1189
rect 2847 1078 2863 1622
rect 2927 1078 2943 1622
rect 3566 1622 3662 1638
rect 3110 1511 3430 1530
rect 3106 1510 3430 1511
rect 3106 1190 3107 1510
rect 3427 1190 3430 1510
rect 3106 1189 3430 1190
rect 2847 1062 2943 1078
rect 2387 810 2710 811
rect 2387 490 2388 810
rect 2708 490 2710 810
rect 2387 489 2710 490
rect 2128 362 2224 378
rect 2390 290 2710 489
rect 2847 922 2943 938
rect 2847 378 2863 922
rect 2927 378 2943 922
rect 3110 811 3430 1189
rect 3566 1078 3582 1622
rect 3646 1078 3662 1622
rect 4285 1622 4381 1638
rect 3830 1511 4150 1530
rect 3825 1510 4150 1511
rect 3825 1190 3826 1510
rect 4146 1190 4150 1510
rect 3825 1189 4150 1190
rect 3566 1062 3662 1078
rect 3106 810 3430 811
rect 3106 490 3107 810
rect 3427 490 3430 810
rect 3106 489 3430 490
rect 2847 362 2943 378
rect 3110 290 3430 489
rect 3566 922 3662 938
rect 3566 378 3582 922
rect 3646 378 3662 922
rect 3830 811 4150 1189
rect 4285 1078 4301 1622
rect 4365 1078 4381 1622
rect 5004 1622 5100 1638
rect 4550 1511 4870 1530
rect 4544 1510 4870 1511
rect 4544 1190 4545 1510
rect 4865 1190 4870 1510
rect 4544 1189 4870 1190
rect 4285 1062 4381 1078
rect 3825 810 4150 811
rect 3825 490 3826 810
rect 4146 490 4150 810
rect 3825 489 4150 490
rect 3566 362 3662 378
rect 3830 290 4150 489
rect 4285 922 4381 938
rect 4285 378 4301 922
rect 4365 378 4381 922
rect 4550 811 4870 1189
rect 5004 1078 5020 1622
rect 5084 1078 5100 1622
rect 5723 1622 5819 1638
rect 5270 1511 5590 1530
rect 5263 1510 5590 1511
rect 5263 1190 5264 1510
rect 5584 1190 5590 1510
rect 5263 1189 5590 1190
rect 5004 1062 5100 1078
rect 4544 810 4870 811
rect 4544 490 4545 810
rect 4865 490 4870 810
rect 4544 489 4870 490
rect 4285 362 4381 378
rect 4550 290 4870 489
rect 5004 922 5100 938
rect 5004 378 5020 922
rect 5084 378 5100 922
rect 5270 811 5590 1189
rect 5723 1078 5739 1622
rect 5803 1078 5819 1622
rect 6442 1622 6538 1638
rect 5990 1511 6310 1530
rect 5982 1510 6310 1511
rect 5982 1190 5983 1510
rect 6303 1190 6310 1510
rect 5982 1189 6310 1190
rect 5723 1062 5819 1078
rect 5263 810 5590 811
rect 5263 490 5264 810
rect 5584 490 5590 810
rect 5263 489 5590 490
rect 5004 362 5100 378
rect 5270 290 5590 489
rect 5723 922 5819 938
rect 5723 378 5739 922
rect 5803 378 5819 922
rect 5990 811 6310 1189
rect 6442 1078 6458 1622
rect 6522 1078 6538 1622
rect 7161 1622 7257 1638
rect 6710 1511 7030 1530
rect 6701 1510 7030 1511
rect 6701 1190 6702 1510
rect 7022 1190 7030 1510
rect 6701 1189 7030 1190
rect 6442 1062 6538 1078
rect 5982 810 6310 811
rect 5982 490 5983 810
rect 6303 490 6310 810
rect 5982 489 6310 490
rect 5723 362 5819 378
rect 5990 290 6310 489
rect 6442 922 6538 938
rect 6442 378 6458 922
rect 6522 378 6538 922
rect 6710 811 7030 1189
rect 7161 1078 7177 1622
rect 7241 1078 7257 1622
rect 7161 1062 7257 1078
rect 6701 810 7030 811
rect 6701 490 6702 810
rect 7022 490 7030 810
rect 6701 489 7030 490
rect 6442 362 6538 378
rect 6710 290 7030 489
rect 7161 922 7257 938
rect 7161 378 7177 922
rect 7241 378 7257 922
rect 7161 362 7257 378
rect 92 260 7260 290
rect 92 160 112 260
rect 272 160 7260 260
rect 92 150 7260 160
<< labels >>
flabel metal2 90 1570 290 1650 1 FreeSans 800 0 0 0 Cin
port 1 n default bidirectional
flabel metal2 112 160 272 260 1 FreeSans 800 0 0 0 Cout
port 2 n default bidirectional
flabel metal1 92 1850 152 1910 1 FreeSans 800 0 0 0 VPWR
port 3 n power bidirectional
flabel metal1 92 -30 152 30 1 FreeSans 800 0 0 0 VGND
port 4 n ground bidirectional
<< properties >>
string FIXED_BBOX 0 0 7371 1880
string LEFclass CORE
string LEFsite unitasc
<< end >>
