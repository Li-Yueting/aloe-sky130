.subckt sky130_asc_pfet_01v8_lvt_1 GATE SOURCE DRAIN VGND VPWR
X0 SOURCE GATE DRAIN VPWR sky130_fd_pr__pfet_01v8_lvt ad=1.8705e+12p pd=1.348e+07u as=1.8705e+12p ps=1.348e+07u w=6.45e+06u l=2e+06u
.ends


.subckt sky130_asc_nfet_01v8_lvt_1 GATE SOURCE DRAIN VPWR VGND
X0 SOURCE GATE DRAIN VGND sky130_fd_pr__nfet_01v8_lvt ad=1.16e+12p pd=8.58e+06u as=1.16e+12p ps=8.58e+06u w=4e+06u l=2e+06u
.ends


