VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO sky130_asc_pfet_01v8_lvt_1
  CLASS CORE ;
  FOREIGN sky130_asc_pfet_01v8_lvt_1 ;
  ORIGIN 0.000 0.000 ;
  SIZE 2.940 BY 9.400 ;
  SITE unitasc ;
  PIN GATE
    DIRECTION INOUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 12.900000 ;
    PORT
      LAYER li1 ;
        RECT 0.000 0.520 2.940 0.820 ;
    END
  END GATE
  PIN SOURCE
    DIRECTION INOUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.870500 ;
    PORT
      LAYER li1 ;
        RECT 0.000 8.650 2.940 8.950 ;
        RECT 2.525 8.245 2.695 8.650 ;
        RECT 2.525 8.130 2.700 8.245 ;
        RECT 2.530 1.755 2.700 8.130 ;
      LAYER mcon ;
        RECT 2.530 1.835 2.700 8.165 ;
      LAYER met1 ;
        RECT 2.500 1.775 2.730 8.225 ;
    END
  END SOURCE
  PIN DRAIN
    DIRECTION INOUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.870500 ;
    PORT
      LAYER li1 ;
        RECT 0.240 1.870 0.410 8.245 ;
        RECT 0.235 1.755 0.410 1.870 ;
        RECT 0.235 1.350 0.405 1.755 ;
        RECT 0.000 1.050 2.940 1.350 ;
      LAYER mcon ;
        RECT 0.240 1.835 0.410 8.165 ;
      LAYER met1 ;
        RECT 0.210 1.775 0.440 8.225 ;
    END
  END DRAIN
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT 0.000 1.465 2.940 9.700 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER li1 ;
        RECT 0.000 9.250 2.940 9.550 ;
      LAYER mcon ;
        RECT 0.850 9.250 1.150 9.550 ;
      LAYER met1 ;
        RECT 0.000 9.100 2.940 9.700 ;
    END
  END VPWR
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER li1 ;
        RECT 0.000 -0.150 2.940 0.150 ;
      LAYER mcon ;
        RECT 0.850 -0.150 1.150 0.150 ;
      LAYER met1 ;
        RECT 0.000 -0.300 2.940 0.300 ;
    END
  END VGND
END sky130_asc_pfet_01v8_lvt_1

#--------EOF---------

MACRO sky130_asc_nfet_01v8_lvt_1
  CLASS CORE ;
  FOREIGN sky130_asc_nfet_01v8_lvt_1 ;
  ORIGIN 0.000 0.000 ;
  SIZE 2.580 BY 9.400 ;
  SITE unitasc ;
  PIN VNB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER pwell ;
        RECT 0.000 0.150 2.580 5.000 ;
        RECT 0.150 -0.150 0.450 0.150 ;
    END
  END VNB
  PIN GATE
    DIRECTION INOUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 8.000000 ;
    PORT
      LAYER li1 ;
        RECT 0.000 0.720 2.580 1.020 ;
    END
  END GATE
  PIN SOURCE
    DIRECTION INOUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.160000 ;
    PORT
      LAYER li1 ;
        RECT 0.000 8.250 2.580 8.550 ;
        RECT 2.345 7.020 2.515 8.250 ;
        RECT 2.345 6.730 2.520 7.020 ;
        RECT 2.350 2.980 2.520 6.730 ;
      LAYER mcon ;
        RECT 2.350 3.060 2.520 6.940 ;
      LAYER met1 ;
        RECT 2.320 3.000 2.550 7.000 ;
    END
  END SOURCE
  PIN DRAIN
    DIRECTION INOUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.160000 ;
    PORT
      LAYER li1 ;
        RECT 0.060 3.270 0.230 7.020 ;
        RECT 0.055 2.980 0.230 3.270 ;
        RECT 0.055 2.520 0.225 2.980 ;
        RECT 0.000 2.220 2.580 2.520 ;
      LAYER mcon ;
        RECT 0.060 3.060 0.230 6.940 ;
      LAYER met1 ;
        RECT 0.030 3.000 0.260 7.000 ;
    END
  END DRAIN
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER li1 ;
        RECT 0.000 9.250 2.580 9.550 ;
      LAYER mcon ;
        RECT 0.850 9.250 1.150 9.550 ;
      LAYER met1 ;
        RECT 0.000 9.100 2.580 9.700 ;
    END
  END VPWR
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER li1 ;
        RECT 0.000 -0.150 2.580 0.150 ;
      LAYER mcon ;
        RECT 0.850 -0.150 1.150 0.150 ;
      LAYER met1 ;
        RECT 0.000 -0.300 2.580 0.300 ;
    END
  END VGND
END sky130_asc_nfet_01v8_lvt_1

# -------------EOF--------------------

MACRO sky130_fd_sc_hd__inv_2
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__inv_2 ;
  ORIGIN 0.000 0.000 ;
  SIZE 1.380 BY 2.720 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.495000 ;
    PORT
      LAYER li1 ;
        RECT 0.105 1.075 0.435 1.325 ;
    END
  END A
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met1 ;
        RECT 0.000 -0.240 1.380 0.240 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.015 0.105 1.365 1.015 ;
        RECT 0.145 -0.085 0.315 0.105 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190 1.305 1.570 2.910 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met1 ;
        RECT 0.000 2.480 1.380 2.960 ;
    END
  END VPWR
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER li1 ;
        RECT 0.525 1.485 0.855 2.465 ;
        RECT 0.605 0.885 0.855 1.485 ;
        RECT 0.525 0.255 0.855 0.885 ;
    END
  END Y
  OBS
      LAYER li1 ;
        RECT 0.000 2.635 1.380 2.805 ;
        RECT 0.125 1.495 0.355 2.635 ;
        RECT 1.025 1.495 1.235 2.635 ;
        RECT 0.125 0.085 0.355 0.905 ;
        RECT 1.025 0.085 1.235 0.905 ;
        RECT 0.000 -0.085 1.380 0.085 ;
      LAYER mcon ;
        RECT 0.145 2.635 0.315 2.805 ;
        RECT 0.605 2.635 0.775 2.805 ;
        RECT 1.065 2.635 1.235 2.805 ;
        RECT 0.145 -0.085 0.315 0.085 ;
        RECT 0.605 -0.085 0.775 0.085 ;
        RECT 1.065 -0.085 1.235 0.085 ;
  END
END sky130_fd_sc_hd__inv_2

END LIBRARY





