magic
tech sky130A
magscale 1 2
timestamp 1652142558
<< pwell >>
rect 0 -60 2440 1650
<< psubdiff >>
rect 912 940 1528 970
rect 912 820 972 940
rect 1468 820 1528 940
rect 912 790 1528 820
<< psubdiffcont >>
rect 972 820 1468 940
<< xpolycontact >>
rect 0 1075 432 1645
rect 2008 1075 2440 1645
rect 0 115 432 685
rect 2008 115 2440 685
<< xpolyres >>
rect 432 1075 2008 1645
rect 432 115 2008 685
<< locali >>
rect 0 1850 170 1910
rect 230 1850 370 1910
rect 430 1850 570 1910
rect 630 1850 770 1910
rect 830 1850 970 1910
rect 1030 1850 1170 1910
rect 1230 1850 1370 1910
rect 1430 1850 1570 1910
rect 1630 1850 1770 1910
rect 1830 1850 1970 1910
rect 2030 1850 2170 1910
rect 2230 1850 2440 1910
rect 912 940 1528 970
rect 912 820 972 940
rect 1468 820 1528 940
rect 912 30 1528 820
rect 2008 685 2440 1075
rect 0 -30 170 30
rect 230 -30 370 30
rect 430 -30 570 30
rect 630 -30 770 30
rect 830 -30 970 30
rect 1030 -30 1170 30
rect 1230 -30 1370 30
rect 1430 -30 1570 30
rect 1630 -30 1770 30
rect 1830 -30 1970 30
rect 2030 -30 2170 30
rect 2230 -30 2440 30
<< viali >>
rect 170 1850 230 1910
rect 370 1850 430 1910
rect 570 1850 630 1910
rect 770 1850 830 1910
rect 970 1850 1030 1910
rect 1170 1850 1230 1910
rect 1370 1850 1430 1910
rect 1570 1850 1630 1910
rect 1770 1850 1830 1910
rect 1970 1850 2030 1910
rect 2170 1850 2230 1910
rect 18 1091 415 1629
rect 2025 1091 2422 1629
rect 18 131 415 669
rect 2025 131 2422 669
rect 170 -30 230 30
rect 370 -30 430 30
rect 570 -30 630 30
rect 770 -30 830 30
rect 970 -30 1030 30
rect 1170 -30 1230 30
rect 1370 -30 1430 30
rect 1570 -30 1630 30
rect 1770 -30 1830 30
rect 1970 -30 2030 30
rect 2170 -30 2230 30
<< metal1 >>
rect 0 1910 2440 1940
rect 0 1850 170 1910
rect 230 1850 370 1910
rect 430 1850 570 1910
rect 630 1850 770 1910
rect 830 1850 970 1910
rect 1030 1850 1170 1910
rect 1230 1850 1370 1910
rect 1430 1850 1570 1910
rect 1630 1850 1770 1910
rect 1830 1850 1970 1910
rect 2030 1850 2170 1910
rect 2230 1850 2440 1910
rect 0 1820 2440 1850
rect 11 1629 421 1641
rect 11 1091 18 1629
rect 415 1091 421 1629
rect 11 1079 421 1091
rect 2019 1629 2429 1641
rect 2019 1091 2025 1629
rect 2422 1091 2429 1629
rect 2019 1079 2429 1091
rect 11 669 421 681
rect 11 131 18 669
rect 415 131 421 669
rect 11 119 421 131
rect 2008 669 2440 1079
rect 2008 131 2025 669
rect 2422 131 2440 669
rect 2008 115 2440 131
rect 0 30 2440 60
rect 0 -30 170 30
rect 230 -30 370 30
rect 430 -30 570 30
rect 630 -30 770 30
rect 830 -30 970 30
rect 1030 -30 1170 30
rect 1230 -30 1370 30
rect 1430 -30 1570 30
rect 1630 -30 1770 30
rect 1830 -30 1970 30
rect 2030 -30 2170 30
rect 2230 -30 2440 30
rect 0 -60 2440 -30
<< labels >>
flabel metal1 120 1300 240 1420 1 FreeSans 480 0 0 0 Rin
port 1 n default bidirectional
flabel metal1 120 340 240 460 1 FreeSans 480 0 0 0 Rout
port 2 n default bidirectional
flabel metal1 0 1850 60 1910 1 FreeSans 800 0 0 0 VPWR
port 3 n power bidirectional
flabel metal1 0 -30 60 30 1 FreeSans 800 0 0 0 VGND
port 4 n ground bidirectional
<< properties >>
string FIXED_BBOX 0 0 2440 1880
string LEFclass CORE
string LEFsite unitasc
<< end >>
