magic
tech sky130A
magscale 1 2
timestamp 1654738924
<< nwell >>
rect -2742 -562 2644 940
<< nsubdiff >>
rect -1646 808 -1526 810
rect -2704 760 -2664 800
rect -1646 772 -1606 808
rect -1562 772 -1526 808
rect -1646 770 -1526 772
rect -346 808 -226 810
rect -346 772 -306 808
rect -262 772 -226 808
rect -346 770 -226 772
rect 954 808 1074 810
rect 954 772 994 808
rect 1038 772 1074 808
rect 954 770 1074 772
rect -2704 680 -2664 720
<< nsubdiffcont >>
rect -1606 772 -1562 808
rect -306 772 -262 808
rect 994 772 1038 808
rect -2704 720 -2664 760
<< poly >>
rect -2518 -672 -2398 -502
rect -2259 -672 -2139 -502
rect -2000 -672 -1880 -502
rect -1741 -672 -1621 -502
rect -1482 -672 -1362 -502
rect -1223 -672 -1103 -502
rect -964 -672 -844 -502
rect -705 -672 -585 -502
rect -446 -672 -326 -502
rect -187 -672 -67 -502
rect 72 -672 192 -502
rect 331 -672 451 -502
rect 590 -672 710 -502
rect 849 -672 969 -502
rect 1108 -672 1228 -502
rect 1367 -672 1487 -502
rect 1626 -672 1746 -502
rect 1885 -672 2005 -502
rect 2144 -672 2264 -502
rect 2403 -672 2523 -502
rect -2644 -692 2644 -672
rect -2644 -752 -2474 -692
rect -2414 -752 -2274 -692
rect -2214 -752 -2074 -692
rect -2014 -752 -1874 -692
rect -1814 -752 -1674 -692
rect -1614 -752 -1474 -692
rect -1414 -752 -1274 -692
rect -1214 -752 -1074 -692
rect -1014 -752 -874 -692
rect -814 -752 -674 -692
rect -614 -752 -474 -692
rect -414 -752 -274 -692
rect -214 -752 -74 -692
rect -14 -752 126 -692
rect 186 -752 326 -692
rect 386 -752 526 -692
rect 586 -752 726 -692
rect 786 -752 926 -692
rect 986 -752 1126 -692
rect 1186 -752 1326 -692
rect 1386 -752 1526 -692
rect 1586 -752 1726 -692
rect 1786 -752 1926 -692
rect 1986 -752 2126 -692
rect 2186 -752 2326 -692
rect 2386 -752 2526 -692
rect 2586 -752 2644 -692
rect -2644 -772 2644 -752
<< polycont >>
rect -2474 -752 -2414 -692
rect -2274 -752 -2214 -692
rect -2074 -752 -2014 -692
rect -1874 -752 -1814 -692
rect -1674 -752 -1614 -692
rect -1474 -752 -1414 -692
rect -1274 -752 -1214 -692
rect -1074 -752 -1014 -692
rect -874 -752 -814 -692
rect -674 -752 -614 -692
rect -474 -752 -414 -692
rect -274 -752 -214 -692
rect -74 -752 -14 -692
rect 126 -752 186 -692
rect 326 -752 386 -692
rect 526 -752 586 -692
rect 726 -752 786 -692
rect 926 -752 986 -692
rect 1126 -752 1186 -692
rect 1326 -752 1386 -692
rect 1526 -752 1586 -692
rect 1726 -752 1786 -692
rect 1926 -752 1986 -692
rect 2126 -752 2186 -692
rect 2326 -752 2386 -692
rect 2526 -752 2586 -692
<< locali >>
rect -2742 850 -2474 910
rect -2414 850 -2274 910
rect -2214 850 -2074 910
rect -2014 850 -1874 910
rect -1814 850 -1674 910
rect -1614 850 -1474 910
rect -1414 850 -1274 910
rect -1214 850 -1074 910
rect -1014 850 -874 910
rect -814 850 -674 910
rect -614 850 -474 910
rect -414 850 -274 910
rect -214 850 -74 910
rect -14 850 126 910
rect 186 850 326 910
rect 386 850 526 910
rect 586 850 726 910
rect 786 850 926 910
rect 986 850 1126 910
rect 1186 850 1326 910
rect 1386 850 1526 910
rect 1586 850 1726 910
rect 1786 850 1926 910
rect 1986 850 2126 910
rect 2186 850 2326 910
rect 2386 850 2526 910
rect 2586 850 2644 910
rect -2714 760 -2654 850
rect -1666 808 -1506 850
rect -1666 772 -1606 808
rect -1562 772 -1506 808
rect -1666 770 -1506 772
rect -366 808 -206 850
rect -366 772 -306 808
rect -262 772 -206 808
rect -366 770 -206 772
rect 934 808 1094 850
rect 934 772 994 808
rect 1038 772 1094 808
rect 934 770 1094 772
rect -2714 720 -2704 760
rect -2664 720 -2654 760
rect -2714 640 -2654 720
rect -2584 690 2644 730
rect -2339 482 -2305 690
rect -1823 482 -1789 690
rect -1307 482 -1273 690
rect -791 482 -757 690
rect -275 482 -241 690
rect 241 482 275 690
rect 757 482 791 690
rect 1273 482 1307 690
rect 1789 482 1823 690
rect 2305 482 2339 690
rect -2597 -692 -2563 -482
rect -2081 -692 -2047 -482
rect -1565 -692 -1531 -482
rect -1049 -692 -1015 -482
rect -533 -692 -499 -482
rect -17 -692 17 -482
rect 499 -692 533 -482
rect 1015 -692 1049 -482
rect 1531 -692 1565 -482
rect 2047 -692 2081 -482
rect 2563 -692 2597 -482
rect -2644 -752 -2474 -692
rect -2414 -752 -2274 -692
rect -2214 -752 -2074 -692
rect -2014 -752 -1874 -692
rect -1814 -752 -1674 -692
rect -1614 -752 -1474 -692
rect -1414 -752 -1274 -692
rect -1214 -752 -1074 -692
rect -1014 -752 -874 -692
rect -814 -752 -674 -692
rect -614 -752 -474 -692
rect -414 -752 -274 -692
rect -214 -752 -74 -692
rect -14 -752 126 -692
rect 186 -752 326 -692
rect 386 -752 526 -692
rect 586 -752 726 -692
rect 786 -752 926 -692
rect 986 -752 1126 -692
rect 1186 -752 1326 -692
rect 1386 -752 1526 -692
rect 1586 -752 1726 -692
rect 1786 -752 1926 -692
rect 1986 -752 2126 -692
rect 2186 -752 2326 -692
rect 2386 -752 2526 -692
rect 2586 -752 2644 -692
rect -2644 -790 2644 -752
rect -2742 -1030 -2474 -970
rect -2414 -1030 -2274 -970
rect -2214 -1030 -2074 -970
rect -2014 -1030 -1874 -970
rect -1814 -1030 -1674 -970
rect -1614 -1030 -1474 -970
rect -1414 -1030 -1274 -970
rect -1214 -1030 -1074 -970
rect -1014 -1030 -874 -970
rect -814 -1030 -674 -970
rect -614 -1030 -474 -970
rect -414 -1030 -274 -970
rect -214 -1030 -74 -970
rect -14 -1030 126 -970
rect 186 -1030 326 -970
rect 386 -1030 526 -970
rect 586 -1030 726 -970
rect 786 -1030 926 -970
rect 986 -1030 1126 -970
rect 1186 -1030 1326 -970
rect 1386 -1030 1526 -970
rect 1586 -1030 1726 -970
rect 1786 -1030 1926 -970
rect 1986 -1030 2126 -970
rect 2186 -1030 2326 -970
rect 2386 -1030 2526 -970
rect 2586 -1030 2644 -970
<< viali >>
rect -2474 850 -2414 910
rect -2274 850 -2214 910
rect -2074 850 -2014 910
rect -1874 850 -1814 910
rect -1674 850 -1614 910
rect -1474 850 -1414 910
rect -1274 850 -1214 910
rect -1074 850 -1014 910
rect -874 850 -814 910
rect -674 850 -614 910
rect -474 850 -414 910
rect -274 850 -214 910
rect -74 850 -14 910
rect 126 850 186 910
rect 326 850 386 910
rect 526 850 586 910
rect 726 850 786 910
rect 926 850 986 910
rect 1126 850 1186 910
rect 1326 850 1386 910
rect 1526 850 1586 910
rect 1726 850 1786 910
rect 1926 850 1986 910
rect 2126 850 2186 910
rect 2326 850 2386 910
rect 2526 850 2586 910
rect -2474 -1030 -2414 -970
rect -2274 -1030 -2214 -970
rect -2074 -1030 -2014 -970
rect -1874 -1030 -1814 -970
rect -1674 -1030 -1614 -970
rect -1474 -1030 -1414 -970
rect -1274 -1030 -1214 -970
rect -1074 -1030 -1014 -970
rect -874 -1030 -814 -970
rect -674 -1030 -614 -970
rect -474 -1030 -414 -970
rect -274 -1030 -214 -970
rect -74 -1030 -14 -970
rect 126 -1030 186 -970
rect 326 -1030 386 -970
rect 526 -1030 586 -970
rect 726 -1030 786 -970
rect 926 -1030 986 -970
rect 1126 -1030 1186 -970
rect 1326 -1030 1386 -970
rect 1526 -1030 1586 -970
rect 1726 -1030 1786 -970
rect 1926 -1030 1986 -970
rect 2126 -1030 2186 -970
rect 2326 -1030 2386 -970
rect 2526 -1030 2586 -970
<< metal1 >>
rect -2742 910 2644 940
rect -2742 850 -2474 910
rect -2414 850 -2274 910
rect -2214 850 -2074 910
rect -2014 850 -1874 910
rect -1814 850 -1674 910
rect -1614 850 -1474 910
rect -1414 850 -1274 910
rect -1214 850 -1074 910
rect -1014 850 -874 910
rect -814 850 -674 910
rect -614 850 -474 910
rect -414 850 -274 910
rect -214 850 -74 910
rect -14 850 126 910
rect 186 850 326 910
rect 386 850 526 910
rect 586 850 726 910
rect 786 850 926 910
rect 986 850 1126 910
rect 1186 850 1326 910
rect 1386 850 1526 910
rect 1586 850 1726 910
rect 1786 850 1926 910
rect 1986 850 2126 910
rect 2186 850 2326 910
rect 2386 850 2526 910
rect 2586 850 2644 910
rect -2742 820 2644 850
rect -2742 -970 2644 -940
rect -2742 -1030 -2474 -970
rect -2414 -1030 -2274 -970
rect -2214 -1030 -2074 -970
rect -2014 -1030 -1874 -970
rect -1814 -1030 -1674 -970
rect -1614 -1030 -1474 -970
rect -1414 -1030 -1274 -970
rect -1214 -1030 -1074 -970
rect -1014 -1030 -874 -970
rect -814 -1030 -674 -970
rect -614 -1030 -474 -970
rect -414 -1030 -274 -970
rect -214 -1030 -74 -970
rect -14 -1030 126 -970
rect 186 -1030 326 -970
rect 386 -1030 526 -970
rect 586 -1030 726 -970
rect 786 -1030 926 -970
rect 986 -1030 1126 -970
rect 1186 -1030 1326 -970
rect 1386 -1030 1526 -970
rect 1586 -1030 1726 -970
rect 1786 -1030 1926 -970
rect 1986 -1030 2126 -970
rect 2186 -1030 2326 -970
rect 2386 -1030 2526 -970
rect 2586 -1030 2644 -970
rect -2742 -1060 2644 -1030
use sky130_fd_pr__pfet_01v8_lvt_W76TCA  xm0
timestamp 0
transform 1 0 0 0 1 0
box -2645 -562 2645 562
<< labels >>
flabel nwell -2742 850 -2682 910 1 FreeSans 800 0 0 0 VPWR
flabel metal1 -2742 -1030 -2584 -970 1 FreeSans 800 0 0 0 VGND
flabel locali 2584 690 2644 730 1 FreeSans 800 0 0 0 SOURCE
flabel locali 2584 -790 2644 -730 1 FreeSans 800 0 0 0 DRAIN
flabel locali 2584 -752 2644 -692 1 FreeSans 800 0 0 0 GATE
<< end >>
