VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO sky130_asc_nfet_01v8_lvt_9
  CLASS CORE ;
  FOREIGN sky130_asc_nfet_01v8_lvt_9 ;
  ORIGIN 0.000 0.000 ;
  SIZE 22.590 BY 9.400 ;
  SITE unitasc ;
  PIN GATE
    DIRECTION INOUT ;
    ANTENNAGATEAREA 72.000000 ;
    PORT
      LAYER li1 ;
        RECT 0.600 0.570 21.500 0.870 ;
    END
  END GATE
  PIN SOURCE
    DIRECTION INOUT ;
    ANTENNADIFFAREA 5.800000 ;
    PORT
      LAYER li1 ;
        RECT 0.600 5.950 21.500 6.250 ;
        RECT 2.945 5.670 3.115 5.950 ;
        RECT 7.525 5.670 7.695 5.950 ;
        RECT 12.105 5.670 12.275 5.950 ;
        RECT 16.685 5.670 16.855 5.950 ;
        RECT 21.265 5.670 21.435 5.950 ;
        RECT 2.945 5.380 3.120 5.670 ;
        RECT 7.525 5.380 7.700 5.670 ;
        RECT 12.105 5.380 12.280 5.670 ;
        RECT 16.685 5.380 16.860 5.670 ;
        RECT 21.265 5.380 21.440 5.670 ;
        RECT 2.950 1.630 3.120 5.380 ;
        RECT 7.530 1.630 7.700 5.380 ;
        RECT 12.110 1.630 12.280 5.380 ;
        RECT 16.690 1.630 16.860 5.380 ;
        RECT 21.270 1.630 21.440 5.380 ;
      LAYER mcon ;
        RECT 2.950 1.710 3.120 5.590 ;
        RECT 7.530 1.710 7.700 5.590 ;
        RECT 12.110 1.710 12.280 5.590 ;
        RECT 16.690 1.710 16.860 5.590 ;
        RECT 21.270 1.710 21.440 5.590 ;
      LAYER met1 ;
        RECT 2.920 1.650 3.150 5.650 ;
        RECT 7.500 1.650 7.730 5.650 ;
        RECT 12.080 1.650 12.310 5.650 ;
        RECT 16.660 1.650 16.890 5.650 ;
        RECT 21.240 1.650 21.470 5.650 ;
    END
  END SOURCE
  PIN DRAIN
    DIRECTION INOUT ;
    ANTENNADIFFAREA 5.800000 ;
    PORT
      LAYER li1 ;
        RECT 0.660 1.920 0.830 5.670 ;
        RECT 5.240 1.920 5.410 5.670 ;
        RECT 9.820 1.920 9.990 5.670 ;
        RECT 14.400 1.920 14.570 5.670 ;
        RECT 18.980 1.920 19.150 5.670 ;
        RECT 0.655 1.630 0.830 1.920 ;
        RECT 5.235 1.630 5.410 1.920 ;
        RECT 9.815 1.630 9.990 1.920 ;
        RECT 14.395 1.630 14.570 1.920 ;
        RECT 18.975 1.630 19.150 1.920 ;
        RECT 0.655 1.350 0.825 1.630 ;
        RECT 5.235 1.350 5.405 1.630 ;
        RECT 9.815 1.350 9.985 1.630 ;
        RECT 14.395 1.350 14.565 1.630 ;
        RECT 18.975 1.350 19.145 1.630 ;
        RECT 0.600 1.050 21.500 1.350 ;
      LAYER mcon ;
        RECT 0.660 1.710 0.830 5.590 ;
        RECT 5.240 1.710 5.410 5.590 ;
        RECT 9.820 1.710 9.990 5.590 ;
        RECT 14.400 1.710 14.570 5.590 ;
        RECT 18.980 1.710 19.150 5.590 ;
      LAYER met1 ;
        RECT 0.630 1.650 0.860 5.650 ;
        RECT 5.210 1.650 5.440 5.650 ;
        RECT 9.790 1.650 10.020 5.650 ;
        RECT 14.370 1.650 14.600 5.650 ;
        RECT 18.950 1.650 19.180 5.650 ;
    END
  END DRAIN
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER li1 ;
        RECT 0.600 6.550 21.500 6.850 ;
      LAYER mcon ;
        RECT 1.450 6.550 1.750 6.850 ;
        RECT 3.450 6.550 3.750 6.850 ;
        RECT 5.450 6.550 5.750 6.850 ;
        RECT 7.450 6.550 7.750 6.850 ;
        RECT 9.450 6.550 9.750 6.850 ;
        RECT 11.450 6.550 11.750 6.850 ;
        RECT 13.450 6.550 13.750 6.850 ;
        RECT 15.450 6.550 15.750 6.850 ;
        RECT 17.450 6.550 17.750 6.850 ;
        RECT 19.450 6.550 19.750 6.850 ;
      LAYER met1 ;
        RECT 0.600 6.400 21.500 7.000 ;
    END
  END VPWR
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER li1 ;
        RECT 0.600 -0.150 21.500 0.150 ;
      LAYER mcon ;
        RECT 1.450 -0.150 1.750 0.150 ;
        RECT 3.450 -0.150 3.750 0.150 ;
        RECT 5.450 -0.150 5.750 0.150 ;
        RECT 7.450 -0.150 7.750 0.150 ;
        RECT 9.450 -0.150 9.750 0.150 ;
        RECT 11.450 -0.150 11.750 0.150 ;
        RECT 13.450 -0.150 13.750 0.150 ;
        RECT 15.450 -0.150 15.750 0.150 ;
        RECT 17.450 -0.150 17.750 0.150 ;
        RECT 19.450 -0.150 19.750 0.150 ;
      LAYER met1 ;
        RECT 0.600 -0.300 21.500 0.300 ;
    END
  END VGND
  OBS
      LAYER pwell ;
        RECT 0.600 0.150 21.500 3.650 ;
  END
END sky130_asc_nfet_01v8_lvt_9
END LIBRARY

