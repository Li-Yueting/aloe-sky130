magic
tech sky130A
magscale 1 2
timestamp 1658609781
<< pwell >>
rect 120 30 4300 730
<< nmoslvt >>
rect 178 330 578 1130
rect 636 330 1036 1130
rect 1094 330 1494 1130
rect 1552 330 1952 1130
rect 2010 330 2410 1130
rect 2468 330 2868 1130
rect 2926 330 3326 1130
rect 3384 330 3784 1130
rect 3842 330 4242 1130
<< ndiff >>
rect 120 1118 178 1130
rect 120 342 132 1118
rect 166 342 178 1118
rect 120 330 178 342
rect 578 1118 636 1130
rect 578 342 590 1118
rect 624 342 636 1118
rect 578 330 636 342
rect 1036 1118 1094 1130
rect 1036 342 1048 1118
rect 1082 342 1094 1118
rect 1036 330 1094 342
rect 1494 1118 1552 1130
rect 1494 342 1506 1118
rect 1540 342 1552 1118
rect 1494 330 1552 342
rect 1952 1118 2010 1130
rect 1952 342 1964 1118
rect 1998 342 2010 1118
rect 1952 330 2010 342
rect 2410 1118 2468 1130
rect 2410 342 2422 1118
rect 2456 342 2468 1118
rect 2410 330 2468 342
rect 2868 1118 2926 1130
rect 2868 342 2880 1118
rect 2914 342 2926 1118
rect 2868 330 2926 342
rect 3326 1118 3384 1130
rect 3326 342 3338 1118
rect 3372 342 3384 1118
rect 3326 330 3384 342
rect 3784 1118 3842 1130
rect 3784 342 3796 1118
rect 3830 342 3842 1118
rect 3784 330 3842 342
rect 4242 1118 4300 1130
rect 4242 342 4254 1118
rect 4288 342 4300 1118
rect 4242 330 4300 342
<< ndiffc >>
rect 132 342 166 1118
rect 590 342 624 1118
rect 1048 342 1082 1118
rect 1506 342 1540 1118
rect 1964 342 1998 1118
rect 2422 342 2456 1118
rect 2880 342 2914 1118
rect 3338 342 3372 1118
rect 3796 342 3830 1118
rect 4254 342 4288 1118
<< poly >>
rect 178 1130 578 1156
rect 636 1130 1036 1156
rect 1094 1130 1494 1156
rect 1552 1130 1952 1156
rect 2010 1130 2410 1156
rect 2468 1130 2868 1156
rect 2926 1130 3326 1156
rect 3384 1130 3784 1156
rect 3842 1130 4242 1156
rect 178 304 578 330
rect 636 304 1036 330
rect 1094 304 1494 330
rect 1552 304 1952 330
rect 2010 304 2410 330
rect 2468 304 2868 330
rect 2926 304 3326 330
rect 3384 304 3784 330
rect 3842 304 4242 330
rect 326 194 446 304
rect 782 194 902 304
rect 1238 194 1358 304
rect 1694 194 1814 304
rect 2150 194 2270 304
rect 2606 194 2726 304
rect 3062 194 3182 304
rect 3518 194 3638 304
rect 3974 194 4094 304
rect 120 174 4300 194
rect 120 114 290 174
rect 350 114 690 174
rect 750 114 1090 174
rect 1150 114 1490 174
rect 1550 114 1890 174
rect 1950 114 2290 174
rect 2350 114 2690 174
rect 2750 114 3090 174
rect 3150 114 3490 174
rect 3550 114 3890 174
rect 3950 114 4300 174
rect 120 94 4300 114
<< polycont >>
rect 290 114 350 174
rect 690 114 750 174
rect 1090 114 1150 174
rect 1490 114 1550 174
rect 1890 114 1950 174
rect 2290 114 2350 174
rect 2690 114 2750 174
rect 3090 114 3150 174
rect 3490 114 3550 174
rect 3890 114 3950 174
<< locali >>
rect 120 1310 290 1370
rect 350 1310 690 1370
rect 750 1310 1090 1370
rect 1150 1310 1490 1370
rect 1550 1310 1890 1370
rect 1950 1310 2290 1370
rect 2350 1310 2690 1370
rect 2750 1310 3090 1370
rect 3150 1310 3490 1370
rect 3550 1310 3890 1370
rect 3950 1310 4300 1370
rect 120 1190 4300 1250
rect 589 1134 623 1190
rect 1505 1134 1539 1190
rect 2421 1134 2455 1190
rect 3337 1134 3371 1190
rect 4253 1134 4287 1190
rect 132 1118 166 1134
rect 131 342 132 384
rect 589 1118 624 1134
rect 589 1076 590 1118
rect 131 326 166 342
rect 1048 1118 1082 1134
rect 590 326 624 342
rect 1047 342 1048 384
rect 1505 1118 1540 1134
rect 1505 1076 1506 1118
rect 1047 326 1082 342
rect 1964 1118 1998 1134
rect 1506 326 1540 342
rect 1963 342 1964 384
rect 2421 1118 2456 1134
rect 2421 1076 2422 1118
rect 1963 326 1998 342
rect 2880 1118 2914 1134
rect 2422 326 2456 342
rect 2879 342 2880 384
rect 3337 1118 3372 1134
rect 3337 1076 3338 1118
rect 2879 326 2914 342
rect 3796 1118 3830 1134
rect 3338 326 3372 342
rect 3795 342 3796 384
rect 4253 1118 4288 1134
rect 4253 1076 4254 1118
rect 3795 326 3830 342
rect 4254 326 4288 342
rect 131 270 165 326
rect 1047 270 1081 326
rect 1963 270 1997 326
rect 2879 270 2913 326
rect 3795 270 3829 326
rect 120 210 4300 270
rect 120 114 290 174
rect 350 114 690 174
rect 750 114 1090 174
rect 1150 114 1490 174
rect 1550 114 1890 174
rect 1950 114 2290 174
rect 2350 114 2690 174
rect 2750 114 3090 174
rect 3150 114 3490 174
rect 3550 114 3890 174
rect 3950 114 4300 174
rect 120 -30 290 30
rect 350 -30 690 30
rect 750 -30 1090 30
rect 1150 -30 1490 30
rect 1550 -30 1890 30
rect 1950 -30 2290 30
rect 2350 -30 2690 30
rect 2750 -30 3090 30
rect 3150 -30 3490 30
rect 3550 -30 3890 30
rect 3950 -30 4300 30
<< viali >>
rect 290 1310 350 1370
rect 690 1310 750 1370
rect 1090 1310 1150 1370
rect 1490 1310 1550 1370
rect 1890 1310 1950 1370
rect 2290 1310 2350 1370
rect 2690 1310 2750 1370
rect 3090 1310 3150 1370
rect 3490 1310 3550 1370
rect 3890 1310 3950 1370
rect 132 342 166 1118
rect 590 342 624 1118
rect 1048 342 1082 1118
rect 1506 342 1540 1118
rect 1964 342 1998 1118
rect 2422 342 2456 1118
rect 2880 342 2914 1118
rect 3338 342 3372 1118
rect 3796 342 3830 1118
rect 4254 342 4288 1118
rect 290 -30 350 30
rect 690 -30 750 30
rect 1090 -30 1150 30
rect 1490 -30 1550 30
rect 1890 -30 1950 30
rect 2290 -30 2350 30
rect 2690 -30 2750 30
rect 3090 -30 3150 30
rect 3490 -30 3550 30
rect 3890 -30 3950 30
<< metal1 >>
rect 120 1370 4300 1400
rect 120 1310 290 1370
rect 350 1310 690 1370
rect 750 1310 1090 1370
rect 1150 1310 1490 1370
rect 1550 1310 1890 1370
rect 1950 1310 2290 1370
rect 2350 1310 2690 1370
rect 2750 1310 3090 1370
rect 3150 1310 3490 1370
rect 3550 1310 3890 1370
rect 3950 1310 4300 1370
rect 120 1280 4300 1310
rect 126 1118 172 1130
rect 126 342 132 1118
rect 166 342 172 1118
rect 126 330 172 342
rect 584 1118 630 1130
rect 584 342 590 1118
rect 624 342 630 1118
rect 584 330 630 342
rect 1042 1118 1088 1130
rect 1042 342 1048 1118
rect 1082 342 1088 1118
rect 1042 330 1088 342
rect 1500 1118 1546 1130
rect 1500 342 1506 1118
rect 1540 342 1546 1118
rect 1500 330 1546 342
rect 1958 1118 2004 1130
rect 1958 342 1964 1118
rect 1998 342 2004 1118
rect 1958 330 2004 342
rect 2416 1118 2462 1130
rect 2416 342 2422 1118
rect 2456 342 2462 1118
rect 2416 330 2462 342
rect 2874 1118 2920 1130
rect 2874 342 2880 1118
rect 2914 342 2920 1118
rect 2874 330 2920 342
rect 3332 1118 3378 1130
rect 3332 342 3338 1118
rect 3372 342 3378 1118
rect 3332 330 3378 342
rect 3790 1118 3836 1130
rect 3790 342 3796 1118
rect 3830 342 3836 1118
rect 3790 330 3836 342
rect 4248 1118 4294 1130
rect 4248 342 4254 1118
rect 4288 342 4294 1118
rect 4248 330 4294 342
rect 120 30 4300 60
rect 120 -30 290 30
rect 350 -30 690 30
rect 750 -30 1090 30
rect 1150 -30 1490 30
rect 1550 -30 1890 30
rect 1950 -30 2290 30
rect 2350 -30 2690 30
rect 2750 -30 3090 30
rect 3150 -30 3490 30
rect 3550 -30 3890 30
rect 3950 -30 4300 30
rect 120 -60 4300 -30
<< labels >>
flabel metal1 120 1310 180 1370 1 FreeSans 480 0 0 0 VPWR
port 4 n power bidirectional
flabel metal1 120 -30 180 30 1 FreeSans 480 0 0 0 VGND
port 5 n ground bidirectional
flabel locali 4240 1190 4300 1250 1 FreeSans 480 0 0 0 SOURCE
port 2 n default bidirectional
flabel locali 4240 210 4300 270 1 FreeSans 480 0 0 0 DRAIN
port 3 n default bidirectional
flabel locali 4240 114 4300 174 1 FreeSans 480 0 0 0 GATE
port 1 n default bidirectional
<< properties >>
string FIXED_BBOX 0 0 4518 1880
string LEFclass CORE
string LEFsite unitasc
<< end >>
