* NGSPICE file created from my_analog_mux.ext - technology: sky130A

.subckt sky130_fd_pr__pfet_01v8_UNG2NQ a_n416_n136# a_352_n136# a_n128_n136# a_n224_n136#
+ a_64_n136# a_160_n136# a_n320_n136# w_n646_n356# a_n32_n136# a_n508_n136# a_448_n136#
+ a_n512_n234# a_256_n136#
X0 a_n224_n136# a_n512_n234# a_n320_n136# w_n646_n356# sky130_fd_pr__pfet_01v8 ad=4.488e+11p pd=3.38e+06u as=4.488e+11p ps=3.38e+06u w=1.36e+06u l=150000u
X1 a_352_n136# a_n512_n234# a_256_n136# w_n646_n356# sky130_fd_pr__pfet_01v8 ad=4.488e+11p pd=3.38e+06u as=4.488e+11p ps=3.38e+06u w=1.36e+06u l=150000u
X2 a_n128_n136# a_n512_n234# a_n224_n136# w_n646_n356# sky130_fd_pr__pfet_01v8 ad=4.488e+11p pd=3.38e+06u as=0p ps=0u w=1.36e+06u l=150000u
X3 a_256_n136# a_n512_n234# a_160_n136# w_n646_n356# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=4.488e+11p ps=3.38e+06u w=1.36e+06u l=150000u
X4 a_n416_n136# a_n512_n234# a_n508_n136# w_n646_n356# sky130_fd_pr__pfet_01v8 ad=4.488e+11p pd=3.38e+06u as=4.216e+11p ps=3.34e+06u w=1.36e+06u l=150000u
X5 a_n320_n136# a_n512_n234# a_n416_n136# w_n646_n356# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.36e+06u l=150000u
X6 a_n32_n136# a_n512_n234# a_n128_n136# w_n646_n356# sky130_fd_pr__pfet_01v8 ad=4.488e+11p pd=3.38e+06u as=0p ps=0u w=1.36e+06u l=150000u
X7 a_448_n136# a_n512_n234# a_352_n136# w_n646_n356# sky130_fd_pr__pfet_01v8 ad=4.216e+11p pd=3.34e+06u as=0p ps=0u w=1.36e+06u l=150000u
X8 a_64_n136# a_n512_n234# a_n32_n136# w_n646_n356# sky130_fd_pr__pfet_01v8 ad=4.488e+11p pd=3.38e+06u as=0p ps=0u w=1.36e+06u l=150000u
X9 a_160_n136# a_n512_n234# a_64_n136# w_n646_n356# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.36e+06u l=150000u
.ends

.subckt sky130_fd_pr__nfet_01v8_6J4AMR a_256_n52# a_n32_n52# a_n224_n52# a_448_n52#
+ a_n416_n52# a_160_n52# a_n610_n226# a_n128_n52# a_n512_n140# a_352_n52# a_n320_n52#
+ a_n508_n52# a_64_n52#
X0 a_n32_n52# a_n512_n140# a_n128_n52# a_n610_n226# sky130_fd_pr__nfet_01v8 ad=1.716e+11p pd=1.7e+06u as=1.716e+11p ps=1.7e+06u w=520000u l=150000u
X1 a_n416_n52# a_n512_n140# a_n508_n52# a_n610_n226# sky130_fd_pr__nfet_01v8 ad=1.716e+11p pd=1.7e+06u as=1.612e+11p ps=1.66e+06u w=520000u l=150000u
X2 a_n224_n52# a_n512_n140# a_n320_n52# a_n610_n226# sky130_fd_pr__nfet_01v8 ad=1.716e+11p pd=1.7e+06u as=1.716e+11p ps=1.7e+06u w=520000u l=150000u
X3 a_n128_n52# a_n512_n140# a_n224_n52# a_n610_n226# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X4 a_n320_n52# a_n512_n140# a_n416_n52# a_n610_n226# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X5 a_160_n52# a_n512_n140# a_64_n52# a_n610_n226# sky130_fd_pr__nfet_01v8 ad=1.716e+11p pd=1.7e+06u as=1.716e+11p ps=1.7e+06u w=520000u l=150000u
X6 a_352_n52# a_n512_n140# a_256_n52# a_n610_n226# sky130_fd_pr__nfet_01v8 ad=1.716e+11p pd=1.7e+06u as=1.716e+11p ps=1.7e+06u w=520000u l=150000u
X7 a_256_n52# a_n512_n140# a_160_n52# a_n610_n226# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X8 a_448_n52# a_n512_n140# a_352_n52# a_n610_n226# sky130_fd_pr__nfet_01v8 ad=1.612e+11p pd=1.66e+06u as=0p ps=0u w=520000u l=150000u
X9 a_64_n52# a_n512_n140# a_n32_n52# a_n610_n226# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
.ends

.subckt transmission_gate m1_n216_396# m1_78_883# VSUBS li_1171_545# m1_97_253# m1_78_76#
Xsky130_fd_pr__pfet_01v8_UNG2NQ_0 m1_n216_396# m1_n216_396# m1_97_253# m1_n216_396#
+ m1_97_253# m1_n216_396# m1_97_253# li_1171_545# m1_n216_396# m1_97_253# m1_97_253#
+ m1_78_883# m1_97_253# sky130_fd_pr__pfet_01v8_UNG2NQ
Xsky130_fd_pr__nfet_01v8_6J4AMR_0 m1_97_253# m1_n216_396# m1_n216_396# m1_97_253#
+ m1_n216_396# m1_n216_396# VSUBS m1_97_253# m1_78_76# m1_n216_396# m1_97_253# m1_97_253#
+ m1_97_253# sky130_fd_pr__nfet_01v8_6J4AMR
.ends

.subckt sky130_fd_pr__nfet_01v8_E56BNL a_n72_n90# a_16_n90# a_n32_32# VSUBS
X0 a_16_n90# a_n32_32# a_n72_n90# VSUBS sky130_fd_pr__nfet_01v8 ad=1.45e+11p pd=1.58e+06u as=1.45e+11p ps=1.58e+06u w=500000u l=150000u
.ends

.subckt switch_5t m1_n53_451# m2_1263_131# m1_1517_361# w_1427_468# m1_2985_451# VSUBS
Xtransmission_gate_0 m1_n53_451# m1_1517_361# VSUBS w_1427_468# m1_1580_239# m2_1263_131#
+ transmission_gate
Xtransmission_gate_1 m1_1580_239# m1_1517_361# VSUBS w_1427_468# m1_2985_451# m2_1263_131#
+ transmission_gate
Xsky130_fd_pr__nfet_01v8_E56BNL_0 VSUBS m1_1580_239# m1_1517_361# VSUBS sky130_fd_pr__nfet_01v8_E56BNL
.ends

.subckt sky130_fd_sc_hd__inv_1 Y A VGND VPWR VNB VPB
X0 Y A VGND VNB sky130_fd_pr__nfet_01v8 ad=1.69e+11p pd=1.82e+06u as=1.69e+11p ps=1.82e+06u w=650000u l=150000u
X1 Y A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=2.6e+11p pd=2.52e+06u as=2.6e+11p ps=2.52e+06u w=1e+06u l=150000u
.ends

.subckt my_one_line sky130_fd_sc_hd__inv_1_0/VPB transmission_gate_0/m1_n216_396#
+ m1_934_370# m1_916_n436# sky130_fd_sc_hd__inv_1_0/A m1_4613_n111# VSUBS
Xswitch_5t_0 m1_915_n115# sky130_fd_sc_hd__inv_1_0/Y sky130_fd_sc_hd__inv_1_0/A sky130_fd_sc_hd__inv_1_0/VPB
+ m1_4613_n111# VSUBS switch_5t
Xtransmission_gate_0 transmission_gate_0/m1_n216_396# m1_934_370# VSUBS sky130_fd_sc_hd__inv_1_0/VPB
+ m1_915_n115# m1_916_n436# transmission_gate
Xsky130_fd_sc_hd__inv_1_0 sky130_fd_sc_hd__inv_1_0/Y sky130_fd_sc_hd__inv_1_0/A VSUBS
+ sky130_fd_sc_hd__inv_1_0/VPB VSUBS sky130_fd_sc_hd__inv_1_0/VPB sky130_fd_sc_hd__inv_1
.ends

.subckt my_analog_mux out en31_b in_31 en30_b in_30 en29_b in_29 en28_b in_28 en27_b
+ in_27 en26_b in_26 en25_b in_25 en24_b in_24 en23_b in_23 en22_b in_22 en21_b in_21
+ en20_b in_20 en19_b in_19 en18_b in_18 en17_b in_17 en16_b in_16 en15_b in_15 en14_b
+ in_14 en13_b in_13 en12_b in_12 en11_b in_11 en10_b in_10 en9_b in_9 en8_b in_8
+ en7_b in_7 en6_b in_6 en5_b in_5 en4_b in_4 en3_b in_3 en2_b in_2 en1_b in_1 en0_b
+ in_0 en_b en  VSS  VDD
Xmy_one_line_0  VDD in_31 en_b en en31_b out  VSS my_one_line
Xmy_one_line_1  VDD in_30 en_b en en30_b out  VSS my_one_line
Xmy_one_line_2  VDD in_29 en_b en en29_b out  VSS my_one_line
Xmy_one_line_4  VDD in_27 en_b en en27_b out  VSS my_one_line
Xmy_one_line_3  VDD in_28 en_b en en28_b out  VSS my_one_line
Xmy_one_line_5  VDD in_26 en_b en en26_b out  VSS my_one_line
Xmy_one_line_6  VDD in_25 en_b en en25_b out  VSS my_one_line
Xmy_one_line_7  VDD in_24 en_b en en24_b out  VSS my_one_line
Xmy_one_line_8  VDD in_23 en_b en en23_b out  VSS my_one_line
Xmy_one_line_9  VDD in_22 en_b en en22_b out  VSS my_one_line
Xmy_one_line_30  VDD in_1 en_b en en1_b out  VSS my_one_line
Xmy_one_line_31  VDD in_0 en_b en en0_b out  VSS my_one_line
Xmy_one_line_20  VDD in_11 en_b en en11_b out  VSS my_one_line
Xmy_one_line_22  VDD in_9 en_b en en9_b out  VSS my_one_line
Xmy_one_line_21  VDD in_10 en_b en en10_b out  VSS my_one_line
Xmy_one_line_11  VDD in_20 en_b en en20_b out  VSS my_one_line
Xmy_one_line_10  VDD in_21 en_b en en21_b out  VSS my_one_line
Xmy_one_line_23  VDD in_8 en_b en en8_b out  VSS my_one_line
Xmy_one_line_12  VDD in_19 en_b en en19_b out  VSS my_one_line
Xmy_one_line_24  VDD in_7 en_b en en7_b out  VSS my_one_line
Xmy_one_line_13  VDD in_18 en_b en en18_b out  VSS my_one_line
Xmy_one_line_25  VDD in_6 en_b en en6_b out  VSS my_one_line
Xmy_one_line_14  VDD in_17 en_b en en17_b out  VSS my_one_line
Xmy_one_line_26  VDD in_5 en_b en en5_b out  VSS my_one_line
Xmy_one_line_15  VDD in_16 en_b en en16_b out  VSS my_one_line
Xmy_one_line_27  VDD in_4 en_b en en4_b out  VSS my_one_line
Xmy_one_line_16  VDD in_15 en_b en en15_b out  VSS my_one_line
Xmy_one_line_28  VDD in_3 en_b en en3_b out  VSS my_one_line
Xmy_one_line_17  VDD in_14 en_b en en14_b out  VSS my_one_line
Xmy_one_line_29  VDD in_2 en_b en en2_b out  VSS my_one_line
Xmy_one_line_19  VDD in_12 en_b en en12_b out  VSS my_one_line
Xmy_one_line_18  VDD in_13 en_b en en13_b out  VSS my_one_line
.ends

