VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO sky130_asc_pnp_05v5_W3p40L3p40_8
  CLASS CORE ;
  FOREIGN sky130_asc_pnp_05v5_W3p40L3p40_8 ;
  ORIGIN 0.000 0.000 ;
  SIZE 54.500 BY 9.400 ;
  SITE unitasc ;
  PIN Emitter
    DIRECTION INOUT ;
    ANTENNADIFFAREA 92.479996 ;
    PORT
      LAYER li1 ;
        RECT 2.065 2.965 5.535 6.435 ;
        RECT 8.765 2.965 12.235 6.435 ;
        RECT 15.465 2.965 18.935 6.435 ;
        RECT 22.165 2.965 25.635 6.435 ;
        RECT 28.865 2.965 32.335 6.435 ;
        RECT 35.565 2.965 39.035 6.435 ;
        RECT 42.265 2.965 45.735 6.435 ;
        RECT 48.965 2.965 52.435 6.435 ;
      LAYER mcon ;
        RECT 2.430 5.830 2.600 6.000 ;
        RECT 2.930 5.830 3.100 6.000 ;
        RECT 3.430 5.830 3.600 6.000 ;
        RECT 3.930 5.830 4.100 6.000 ;
        RECT 4.430 5.830 4.600 6.000 ;
        RECT 4.930 5.830 5.100 6.000 ;
        RECT 2.430 5.330 2.600 5.500 ;
        RECT 2.930 5.330 3.100 5.500 ;
        RECT 3.430 5.330 3.600 5.500 ;
        RECT 3.930 5.330 4.100 5.500 ;
        RECT 4.430 5.330 4.600 5.500 ;
        RECT 4.930 5.330 5.100 5.500 ;
        RECT 2.430 4.830 2.600 5.000 ;
        RECT 2.930 4.830 3.100 5.000 ;
        RECT 3.430 4.830 3.600 5.000 ;
        RECT 3.930 4.830 4.100 5.000 ;
        RECT 4.430 4.830 4.600 5.000 ;
        RECT 4.930 4.830 5.100 5.000 ;
        RECT 2.430 4.330 2.600 4.500 ;
        RECT 2.930 4.330 3.100 4.500 ;
        RECT 3.430 4.330 3.600 4.500 ;
        RECT 3.930 4.330 4.100 4.500 ;
        RECT 4.430 4.330 4.600 4.500 ;
        RECT 4.930 4.330 5.100 4.500 ;
        RECT 2.430 3.830 2.600 4.000 ;
        RECT 2.930 3.830 3.100 4.000 ;
        RECT 3.430 3.830 3.600 4.000 ;
        RECT 3.930 3.830 4.100 4.000 ;
        RECT 4.430 3.830 4.600 4.000 ;
        RECT 4.930 3.830 5.100 4.000 ;
        RECT 2.430 3.330 2.600 3.500 ;
        RECT 2.930 3.330 3.100 3.500 ;
        RECT 3.430 3.330 3.600 3.500 ;
        RECT 3.930 3.330 4.100 3.500 ;
        RECT 4.430 3.330 4.600 3.500 ;
        RECT 4.930 3.330 5.100 3.500 ;
        RECT 9.130 5.830 9.300 6.000 ;
        RECT 9.630 5.830 9.800 6.000 ;
        RECT 10.130 5.830 10.300 6.000 ;
        RECT 10.630 5.830 10.800 6.000 ;
        RECT 11.130 5.830 11.300 6.000 ;
        RECT 11.630 5.830 11.800 6.000 ;
        RECT 9.130 5.330 9.300 5.500 ;
        RECT 9.630 5.330 9.800 5.500 ;
        RECT 10.130 5.330 10.300 5.500 ;
        RECT 10.630 5.330 10.800 5.500 ;
        RECT 11.130 5.330 11.300 5.500 ;
        RECT 11.630 5.330 11.800 5.500 ;
        RECT 9.130 4.830 9.300 5.000 ;
        RECT 9.630 4.830 9.800 5.000 ;
        RECT 10.130 4.830 10.300 5.000 ;
        RECT 10.630 4.830 10.800 5.000 ;
        RECT 11.130 4.830 11.300 5.000 ;
        RECT 11.630 4.830 11.800 5.000 ;
        RECT 9.130 4.330 9.300 4.500 ;
        RECT 9.630 4.330 9.800 4.500 ;
        RECT 10.130 4.330 10.300 4.500 ;
        RECT 10.630 4.330 10.800 4.500 ;
        RECT 11.130 4.330 11.300 4.500 ;
        RECT 11.630 4.330 11.800 4.500 ;
        RECT 9.130 3.830 9.300 4.000 ;
        RECT 9.630 3.830 9.800 4.000 ;
        RECT 10.130 3.830 10.300 4.000 ;
        RECT 10.630 3.830 10.800 4.000 ;
        RECT 11.130 3.830 11.300 4.000 ;
        RECT 11.630 3.830 11.800 4.000 ;
        RECT 9.130 3.330 9.300 3.500 ;
        RECT 9.630 3.330 9.800 3.500 ;
        RECT 10.130 3.330 10.300 3.500 ;
        RECT 10.630 3.330 10.800 3.500 ;
        RECT 11.130 3.330 11.300 3.500 ;
        RECT 11.630 3.330 11.800 3.500 ;
        RECT 15.830 5.830 16.000 6.000 ;
        RECT 16.330 5.830 16.500 6.000 ;
        RECT 16.830 5.830 17.000 6.000 ;
        RECT 17.330 5.830 17.500 6.000 ;
        RECT 17.830 5.830 18.000 6.000 ;
        RECT 18.330 5.830 18.500 6.000 ;
        RECT 15.830 5.330 16.000 5.500 ;
        RECT 16.330 5.330 16.500 5.500 ;
        RECT 16.830 5.330 17.000 5.500 ;
        RECT 17.330 5.330 17.500 5.500 ;
        RECT 17.830 5.330 18.000 5.500 ;
        RECT 18.330 5.330 18.500 5.500 ;
        RECT 15.830 4.830 16.000 5.000 ;
        RECT 16.330 4.830 16.500 5.000 ;
        RECT 16.830 4.830 17.000 5.000 ;
        RECT 17.330 4.830 17.500 5.000 ;
        RECT 17.830 4.830 18.000 5.000 ;
        RECT 18.330 4.830 18.500 5.000 ;
        RECT 15.830 4.330 16.000 4.500 ;
        RECT 16.330 4.330 16.500 4.500 ;
        RECT 16.830 4.330 17.000 4.500 ;
        RECT 17.330 4.330 17.500 4.500 ;
        RECT 17.830 4.330 18.000 4.500 ;
        RECT 18.330 4.330 18.500 4.500 ;
        RECT 15.830 3.830 16.000 4.000 ;
        RECT 16.330 3.830 16.500 4.000 ;
        RECT 16.830 3.830 17.000 4.000 ;
        RECT 17.330 3.830 17.500 4.000 ;
        RECT 17.830 3.830 18.000 4.000 ;
        RECT 18.330 3.830 18.500 4.000 ;
        RECT 15.830 3.330 16.000 3.500 ;
        RECT 16.330 3.330 16.500 3.500 ;
        RECT 16.830 3.330 17.000 3.500 ;
        RECT 17.330 3.330 17.500 3.500 ;
        RECT 17.830 3.330 18.000 3.500 ;
        RECT 18.330 3.330 18.500 3.500 ;
        RECT 22.530 5.830 22.700 6.000 ;
        RECT 23.030 5.830 23.200 6.000 ;
        RECT 23.530 5.830 23.700 6.000 ;
        RECT 24.030 5.830 24.200 6.000 ;
        RECT 24.530 5.830 24.700 6.000 ;
        RECT 25.030 5.830 25.200 6.000 ;
        RECT 22.530 5.330 22.700 5.500 ;
        RECT 23.030 5.330 23.200 5.500 ;
        RECT 23.530 5.330 23.700 5.500 ;
        RECT 24.030 5.330 24.200 5.500 ;
        RECT 24.530 5.330 24.700 5.500 ;
        RECT 25.030 5.330 25.200 5.500 ;
        RECT 22.530 4.830 22.700 5.000 ;
        RECT 23.030 4.830 23.200 5.000 ;
        RECT 23.530 4.830 23.700 5.000 ;
        RECT 24.030 4.830 24.200 5.000 ;
        RECT 24.530 4.830 24.700 5.000 ;
        RECT 25.030 4.830 25.200 5.000 ;
        RECT 22.530 4.330 22.700 4.500 ;
        RECT 23.030 4.330 23.200 4.500 ;
        RECT 23.530 4.330 23.700 4.500 ;
        RECT 24.030 4.330 24.200 4.500 ;
        RECT 24.530 4.330 24.700 4.500 ;
        RECT 25.030 4.330 25.200 4.500 ;
        RECT 22.530 3.830 22.700 4.000 ;
        RECT 23.030 3.830 23.200 4.000 ;
        RECT 23.530 3.830 23.700 4.000 ;
        RECT 24.030 3.830 24.200 4.000 ;
        RECT 24.530 3.830 24.700 4.000 ;
        RECT 25.030 3.830 25.200 4.000 ;
        RECT 22.530 3.330 22.700 3.500 ;
        RECT 23.030 3.330 23.200 3.500 ;
        RECT 23.530 3.330 23.700 3.500 ;
        RECT 24.030 3.330 24.200 3.500 ;
        RECT 24.530 3.330 24.700 3.500 ;
        RECT 25.030 3.330 25.200 3.500 ;
        RECT 29.230 5.830 29.400 6.000 ;
        RECT 29.730 5.830 29.900 6.000 ;
        RECT 30.230 5.830 30.400 6.000 ;
        RECT 30.730 5.830 30.900 6.000 ;
        RECT 31.230 5.830 31.400 6.000 ;
        RECT 31.730 5.830 31.900 6.000 ;
        RECT 29.230 5.330 29.400 5.500 ;
        RECT 29.730 5.330 29.900 5.500 ;
        RECT 30.230 5.330 30.400 5.500 ;
        RECT 30.730 5.330 30.900 5.500 ;
        RECT 31.230 5.330 31.400 5.500 ;
        RECT 31.730 5.330 31.900 5.500 ;
        RECT 29.230 4.830 29.400 5.000 ;
        RECT 29.730 4.830 29.900 5.000 ;
        RECT 30.230 4.830 30.400 5.000 ;
        RECT 30.730 4.830 30.900 5.000 ;
        RECT 31.230 4.830 31.400 5.000 ;
        RECT 31.730 4.830 31.900 5.000 ;
        RECT 29.230 4.330 29.400 4.500 ;
        RECT 29.730 4.330 29.900 4.500 ;
        RECT 30.230 4.330 30.400 4.500 ;
        RECT 30.730 4.330 30.900 4.500 ;
        RECT 31.230 4.330 31.400 4.500 ;
        RECT 31.730 4.330 31.900 4.500 ;
        RECT 29.230 3.830 29.400 4.000 ;
        RECT 29.730 3.830 29.900 4.000 ;
        RECT 30.230 3.830 30.400 4.000 ;
        RECT 30.730 3.830 30.900 4.000 ;
        RECT 31.230 3.830 31.400 4.000 ;
        RECT 31.730 3.830 31.900 4.000 ;
        RECT 29.230 3.330 29.400 3.500 ;
        RECT 29.730 3.330 29.900 3.500 ;
        RECT 30.230 3.330 30.400 3.500 ;
        RECT 30.730 3.330 30.900 3.500 ;
        RECT 31.230 3.330 31.400 3.500 ;
        RECT 31.730 3.330 31.900 3.500 ;
        RECT 35.930 5.830 36.100 6.000 ;
        RECT 36.430 5.830 36.600 6.000 ;
        RECT 36.930 5.830 37.100 6.000 ;
        RECT 37.430 5.830 37.600 6.000 ;
        RECT 37.930 5.830 38.100 6.000 ;
        RECT 38.430 5.830 38.600 6.000 ;
        RECT 35.930 5.330 36.100 5.500 ;
        RECT 36.430 5.330 36.600 5.500 ;
        RECT 36.930 5.330 37.100 5.500 ;
        RECT 37.430 5.330 37.600 5.500 ;
        RECT 37.930 5.330 38.100 5.500 ;
        RECT 38.430 5.330 38.600 5.500 ;
        RECT 35.930 4.830 36.100 5.000 ;
        RECT 36.430 4.830 36.600 5.000 ;
        RECT 36.930 4.830 37.100 5.000 ;
        RECT 37.430 4.830 37.600 5.000 ;
        RECT 37.930 4.830 38.100 5.000 ;
        RECT 38.430 4.830 38.600 5.000 ;
        RECT 35.930 4.330 36.100 4.500 ;
        RECT 36.430 4.330 36.600 4.500 ;
        RECT 36.930 4.330 37.100 4.500 ;
        RECT 37.430 4.330 37.600 4.500 ;
        RECT 37.930 4.330 38.100 4.500 ;
        RECT 38.430 4.330 38.600 4.500 ;
        RECT 35.930 3.830 36.100 4.000 ;
        RECT 36.430 3.830 36.600 4.000 ;
        RECT 36.930 3.830 37.100 4.000 ;
        RECT 37.430 3.830 37.600 4.000 ;
        RECT 37.930 3.830 38.100 4.000 ;
        RECT 38.430 3.830 38.600 4.000 ;
        RECT 35.930 3.330 36.100 3.500 ;
        RECT 36.430 3.330 36.600 3.500 ;
        RECT 36.930 3.330 37.100 3.500 ;
        RECT 37.430 3.330 37.600 3.500 ;
        RECT 37.930 3.330 38.100 3.500 ;
        RECT 38.430 3.330 38.600 3.500 ;
        RECT 42.630 5.830 42.800 6.000 ;
        RECT 43.130 5.830 43.300 6.000 ;
        RECT 43.630 5.830 43.800 6.000 ;
        RECT 44.130 5.830 44.300 6.000 ;
        RECT 44.630 5.830 44.800 6.000 ;
        RECT 45.130 5.830 45.300 6.000 ;
        RECT 42.630 5.330 42.800 5.500 ;
        RECT 43.130 5.330 43.300 5.500 ;
        RECT 43.630 5.330 43.800 5.500 ;
        RECT 44.130 5.330 44.300 5.500 ;
        RECT 44.630 5.330 44.800 5.500 ;
        RECT 45.130 5.330 45.300 5.500 ;
        RECT 42.630 4.830 42.800 5.000 ;
        RECT 43.130 4.830 43.300 5.000 ;
        RECT 43.630 4.830 43.800 5.000 ;
        RECT 44.130 4.830 44.300 5.000 ;
        RECT 44.630 4.830 44.800 5.000 ;
        RECT 45.130 4.830 45.300 5.000 ;
        RECT 42.630 4.330 42.800 4.500 ;
        RECT 43.130 4.330 43.300 4.500 ;
        RECT 43.630 4.330 43.800 4.500 ;
        RECT 44.130 4.330 44.300 4.500 ;
        RECT 44.630 4.330 44.800 4.500 ;
        RECT 45.130 4.330 45.300 4.500 ;
        RECT 42.630 3.830 42.800 4.000 ;
        RECT 43.130 3.830 43.300 4.000 ;
        RECT 43.630 3.830 43.800 4.000 ;
        RECT 44.130 3.830 44.300 4.000 ;
        RECT 44.630 3.830 44.800 4.000 ;
        RECT 45.130 3.830 45.300 4.000 ;
        RECT 42.630 3.330 42.800 3.500 ;
        RECT 43.130 3.330 43.300 3.500 ;
        RECT 43.630 3.330 43.800 3.500 ;
        RECT 44.130 3.330 44.300 3.500 ;
        RECT 44.630 3.330 44.800 3.500 ;
        RECT 45.130 3.330 45.300 3.500 ;
        RECT 49.330 5.830 49.500 6.000 ;
        RECT 49.830 5.830 50.000 6.000 ;
        RECT 50.330 5.830 50.500 6.000 ;
        RECT 50.830 5.830 51.000 6.000 ;
        RECT 51.330 5.830 51.500 6.000 ;
        RECT 51.830 5.830 52.000 6.000 ;
        RECT 49.330 5.330 49.500 5.500 ;
        RECT 49.830 5.330 50.000 5.500 ;
        RECT 50.330 5.330 50.500 5.500 ;
        RECT 50.830 5.330 51.000 5.500 ;
        RECT 51.330 5.330 51.500 5.500 ;
        RECT 51.830 5.330 52.000 5.500 ;
        RECT 49.330 4.830 49.500 5.000 ;
        RECT 49.830 4.830 50.000 5.000 ;
        RECT 50.330 4.830 50.500 5.000 ;
        RECT 50.830 4.830 51.000 5.000 ;
        RECT 51.330 4.830 51.500 5.000 ;
        RECT 51.830 4.830 52.000 5.000 ;
        RECT 49.330 4.330 49.500 4.500 ;
        RECT 49.830 4.330 50.000 4.500 ;
        RECT 50.330 4.330 50.500 4.500 ;
        RECT 50.830 4.330 51.000 4.500 ;
        RECT 51.330 4.330 51.500 4.500 ;
        RECT 51.830 4.330 52.000 4.500 ;
        RECT 49.330 3.830 49.500 4.000 ;
        RECT 49.830 3.830 50.000 4.000 ;
        RECT 50.330 3.830 50.500 4.000 ;
        RECT 50.830 3.830 51.000 4.000 ;
        RECT 51.330 3.830 51.500 4.000 ;
        RECT 51.830 3.830 52.000 4.000 ;
        RECT 49.330 3.330 49.500 3.500 ;
        RECT 49.830 3.330 50.000 3.500 ;
        RECT 50.330 3.330 50.500 3.500 ;
        RECT 50.830 3.330 51.000 3.500 ;
        RECT 51.330 3.330 51.500 3.500 ;
        RECT 51.830 3.330 52.000 3.500 ;
      LAYER met1 ;
        RECT 2.270 3.170 52.230 6.230 ;
    END
  END Emitter
  PIN Base
    DIRECTION INOUT ;
    ANTENNAGATEAREA 213.831192 ;
    ANTENNADIFFAREA 51.264000 ;
    PORT
      LAYER li1 ;
        RECT 1.395 6.745 6.205 7.105 ;
        RECT 1.395 2.655 1.755 6.745 ;
        RECT 5.845 2.655 6.205 6.745 ;
        RECT 1.395 2.295 6.205 2.655 ;
        RECT 8.095 6.745 12.905 7.105 ;
        RECT 8.095 2.655 8.455 6.745 ;
        RECT 12.545 2.655 12.905 6.745 ;
        RECT 8.095 2.295 12.905 2.655 ;
        RECT 14.795 6.745 19.605 7.105 ;
        RECT 14.795 2.655 15.155 6.745 ;
        RECT 19.245 2.655 19.605 6.745 ;
        RECT 14.795 2.295 19.605 2.655 ;
        RECT 21.495 6.745 26.305 7.105 ;
        RECT 21.495 2.655 21.855 6.745 ;
        RECT 25.945 2.655 26.305 6.745 ;
        RECT 21.495 2.295 26.305 2.655 ;
        RECT 28.195 6.745 33.005 7.105 ;
        RECT 28.195 2.655 28.555 6.745 ;
        RECT 32.645 2.655 33.005 6.745 ;
        RECT 28.195 2.295 33.005 2.655 ;
        RECT 34.895 6.745 39.705 7.105 ;
        RECT 34.895 2.655 35.255 6.745 ;
        RECT 39.345 2.655 39.705 6.745 ;
        RECT 34.895 2.295 39.705 2.655 ;
        RECT 41.595 6.745 46.405 7.105 ;
        RECT 41.595 2.655 41.955 6.745 ;
        RECT 46.045 2.655 46.405 6.745 ;
        RECT 41.595 2.295 46.405 2.655 ;
        RECT 48.295 6.745 53.105 7.105 ;
        RECT 48.295 2.655 48.655 6.745 ;
        RECT 52.745 2.655 53.105 6.745 ;
        RECT 48.295 2.295 53.105 2.655 ;
      LAYER mcon ;
        RECT 1.500 6.850 1.670 7.020 ;
        RECT 1.950 6.850 2.120 7.020 ;
        RECT 2.400 6.850 2.570 7.020 ;
        RECT 2.850 6.850 3.020 7.020 ;
        RECT 3.300 6.850 3.470 7.020 ;
        RECT 3.750 6.850 3.920 7.020 ;
        RECT 4.200 6.850 4.370 7.020 ;
        RECT 4.650 6.850 4.820 7.020 ;
        RECT 5.100 6.850 5.270 7.020 ;
        RECT 5.550 6.850 5.720 7.020 ;
        RECT 6.000 6.850 6.170 7.020 ;
        RECT 8.200 6.850 8.370 7.020 ;
        RECT 8.650 6.850 8.820 7.020 ;
        RECT 9.100 6.850 9.270 7.020 ;
        RECT 9.550 6.850 9.720 7.020 ;
        RECT 10.000 6.850 10.170 7.020 ;
        RECT 10.450 6.850 10.620 7.020 ;
        RECT 10.900 6.850 11.070 7.020 ;
        RECT 11.350 6.850 11.520 7.020 ;
        RECT 11.800 6.850 11.970 7.020 ;
        RECT 12.250 6.850 12.420 7.020 ;
        RECT 12.700 6.850 12.870 7.020 ;
        RECT 14.900 6.850 15.070 7.020 ;
        RECT 15.350 6.850 15.520 7.020 ;
        RECT 15.800 6.850 15.970 7.020 ;
        RECT 16.250 6.850 16.420 7.020 ;
        RECT 16.700 6.850 16.870 7.020 ;
        RECT 17.150 6.850 17.320 7.020 ;
        RECT 17.600 6.850 17.770 7.020 ;
        RECT 18.050 6.850 18.220 7.020 ;
        RECT 18.500 6.850 18.670 7.020 ;
        RECT 18.950 6.850 19.120 7.020 ;
        RECT 19.400 6.850 19.570 7.020 ;
        RECT 21.600 6.850 21.770 7.020 ;
        RECT 22.050 6.850 22.220 7.020 ;
        RECT 22.500 6.850 22.670 7.020 ;
        RECT 22.950 6.850 23.120 7.020 ;
        RECT 23.400 6.850 23.570 7.020 ;
        RECT 23.850 6.850 24.020 7.020 ;
        RECT 24.300 6.850 24.470 7.020 ;
        RECT 24.750 6.850 24.920 7.020 ;
        RECT 25.200 6.850 25.370 7.020 ;
        RECT 25.650 6.850 25.820 7.020 ;
        RECT 26.100 6.850 26.270 7.020 ;
        RECT 28.300 6.850 28.470 7.020 ;
        RECT 28.750 6.850 28.920 7.020 ;
        RECT 29.200 6.850 29.370 7.020 ;
        RECT 29.650 6.850 29.820 7.020 ;
        RECT 30.100 6.850 30.270 7.020 ;
        RECT 30.550 6.850 30.720 7.020 ;
        RECT 31.000 6.850 31.170 7.020 ;
        RECT 31.450 6.850 31.620 7.020 ;
        RECT 31.900 6.850 32.070 7.020 ;
        RECT 32.350 6.850 32.520 7.020 ;
        RECT 32.800 6.850 32.970 7.020 ;
        RECT 35.000 6.850 35.170 7.020 ;
        RECT 35.450 6.850 35.620 7.020 ;
        RECT 35.900 6.850 36.070 7.020 ;
        RECT 36.350 6.850 36.520 7.020 ;
        RECT 36.800 6.850 36.970 7.020 ;
        RECT 37.250 6.850 37.420 7.020 ;
        RECT 37.700 6.850 37.870 7.020 ;
        RECT 38.150 6.850 38.320 7.020 ;
        RECT 38.600 6.850 38.770 7.020 ;
        RECT 39.050 6.850 39.220 7.020 ;
        RECT 39.500 6.850 39.670 7.020 ;
        RECT 41.700 6.850 41.870 7.020 ;
        RECT 42.150 6.850 42.320 7.020 ;
        RECT 42.600 6.850 42.770 7.020 ;
        RECT 43.050 6.850 43.220 7.020 ;
        RECT 43.500 6.850 43.670 7.020 ;
        RECT 43.950 6.850 44.120 7.020 ;
        RECT 44.400 6.850 44.570 7.020 ;
        RECT 44.850 6.850 45.020 7.020 ;
        RECT 45.300 6.850 45.470 7.020 ;
        RECT 45.750 6.850 45.920 7.020 ;
        RECT 46.200 6.850 46.370 7.020 ;
        RECT 48.400 6.850 48.570 7.020 ;
        RECT 48.850 6.850 49.020 7.020 ;
        RECT 49.300 6.850 49.470 7.020 ;
        RECT 49.750 6.850 49.920 7.020 ;
        RECT 50.200 6.850 50.370 7.020 ;
        RECT 50.650 6.850 50.820 7.020 ;
        RECT 51.100 6.850 51.270 7.020 ;
        RECT 51.550 6.850 51.720 7.020 ;
        RECT 52.000 6.850 52.170 7.020 ;
        RECT 52.450 6.850 52.620 7.020 ;
        RECT 52.900 6.850 53.070 7.020 ;
      LAYER met1 ;
        RECT 1.400 6.750 53.100 7.100 ;
    END
  END Base
  PIN Collector
    DIRECTION INOUT ;
    ANTENNADIFFAREA 107.630394 ;
    PORT
      LAYER pwell ;
        RECT 0.450 7.285 54.050 8.050 ;
        RECT 0.450 2.115 1.215 7.285 ;
        RECT 6.385 2.115 7.915 7.285 ;
        RECT 13.085 2.115 14.615 7.285 ;
        RECT 19.785 2.115 21.315 7.285 ;
        RECT 26.485 2.115 28.015 7.285 ;
        RECT 33.185 2.115 34.715 7.285 ;
        RECT 39.885 2.115 41.415 7.285 ;
        RECT 46.585 2.115 48.115 7.285 ;
        RECT 53.285 2.115 54.050 7.285 ;
        RECT 0.450 1.350 54.050 2.115 ;
      LAYER li1 ;
        RECT 0.580 7.425 53.920 7.920 ;
        RECT 0.580 1.975 1.075 7.425 ;
        RECT 6.525 1.975 7.775 7.425 ;
        RECT 13.225 1.975 14.475 7.425 ;
        RECT 19.925 1.975 21.175 7.425 ;
        RECT 26.625 1.975 27.875 7.425 ;
        RECT 33.325 1.975 34.575 7.425 ;
        RECT 40.025 1.975 41.275 7.425 ;
        RECT 46.725 1.975 47.975 7.425 ;
        RECT 53.425 1.975 53.920 7.425 ;
        RECT 0.580 1.480 53.920 1.975 ;
      LAYER mcon ;
        RECT 0.680 7.650 0.850 7.820 ;
        RECT 1.130 7.650 1.300 7.820 ;
        RECT 1.580 7.650 1.750 7.820 ;
        RECT 2.030 7.650 2.200 7.820 ;
        RECT 2.480 7.650 2.650 7.820 ;
        RECT 2.930 7.650 3.100 7.820 ;
        RECT 3.380 7.650 3.550 7.820 ;
        RECT 3.830 7.650 4.000 7.820 ;
        RECT 4.280 7.650 4.450 7.820 ;
        RECT 4.730 7.650 4.900 7.820 ;
        RECT 5.180 7.650 5.350 7.820 ;
        RECT 5.630 7.650 5.800 7.820 ;
        RECT 6.080 7.650 6.250 7.820 ;
        RECT 6.530 7.650 6.700 7.820 ;
        RECT 7.380 7.650 7.550 7.820 ;
        RECT 7.830 7.650 8.000 7.820 ;
        RECT 8.280 7.650 8.450 7.820 ;
        RECT 8.730 7.650 8.900 7.820 ;
        RECT 9.180 7.650 9.350 7.820 ;
        RECT 9.630 7.650 9.800 7.820 ;
        RECT 10.080 7.650 10.250 7.820 ;
        RECT 10.530 7.650 10.700 7.820 ;
        RECT 10.980 7.650 11.150 7.820 ;
        RECT 11.430 7.650 11.600 7.820 ;
        RECT 11.880 7.650 12.050 7.820 ;
        RECT 12.330 7.650 12.500 7.820 ;
        RECT 12.780 7.650 12.950 7.820 ;
        RECT 13.230 7.650 13.400 7.820 ;
        RECT 14.080 7.650 14.250 7.820 ;
        RECT 14.530 7.650 14.700 7.820 ;
        RECT 14.980 7.650 15.150 7.820 ;
        RECT 15.430 7.650 15.600 7.820 ;
        RECT 15.880 7.650 16.050 7.820 ;
        RECT 16.330 7.650 16.500 7.820 ;
        RECT 16.780 7.650 16.950 7.820 ;
        RECT 17.230 7.650 17.400 7.820 ;
        RECT 17.680 7.650 17.850 7.820 ;
        RECT 18.130 7.650 18.300 7.820 ;
        RECT 18.580 7.650 18.750 7.820 ;
        RECT 19.030 7.650 19.200 7.820 ;
        RECT 19.480 7.650 19.650 7.820 ;
        RECT 19.930 7.650 20.100 7.820 ;
        RECT 20.780 7.650 20.950 7.820 ;
        RECT 21.230 7.650 21.400 7.820 ;
        RECT 21.680 7.650 21.850 7.820 ;
        RECT 22.130 7.650 22.300 7.820 ;
        RECT 22.580 7.650 22.750 7.820 ;
        RECT 23.030 7.650 23.200 7.820 ;
        RECT 23.480 7.650 23.650 7.820 ;
        RECT 23.930 7.650 24.100 7.820 ;
        RECT 24.380 7.650 24.550 7.820 ;
        RECT 24.830 7.650 25.000 7.820 ;
        RECT 25.280 7.650 25.450 7.820 ;
        RECT 25.730 7.650 25.900 7.820 ;
        RECT 26.180 7.650 26.350 7.820 ;
        RECT 26.630 7.650 26.800 7.820 ;
        RECT 27.480 7.650 27.650 7.820 ;
        RECT 27.930 7.650 28.100 7.820 ;
        RECT 28.380 7.650 28.550 7.820 ;
        RECT 28.830 7.650 29.000 7.820 ;
        RECT 29.280 7.650 29.450 7.820 ;
        RECT 29.730 7.650 29.900 7.820 ;
        RECT 30.180 7.650 30.350 7.820 ;
        RECT 30.630 7.650 30.800 7.820 ;
        RECT 31.080 7.650 31.250 7.820 ;
        RECT 31.530 7.650 31.700 7.820 ;
        RECT 31.980 7.650 32.150 7.820 ;
        RECT 32.430 7.650 32.600 7.820 ;
        RECT 32.880 7.650 33.050 7.820 ;
        RECT 33.330 7.650 33.500 7.820 ;
        RECT 34.180 7.650 34.350 7.820 ;
        RECT 34.630 7.650 34.800 7.820 ;
        RECT 35.080 7.650 35.250 7.820 ;
        RECT 35.530 7.650 35.700 7.820 ;
        RECT 35.980 7.650 36.150 7.820 ;
        RECT 36.430 7.650 36.600 7.820 ;
        RECT 36.880 7.650 37.050 7.820 ;
        RECT 37.330 7.650 37.500 7.820 ;
        RECT 37.780 7.650 37.950 7.820 ;
        RECT 38.230 7.650 38.400 7.820 ;
        RECT 38.680 7.650 38.850 7.820 ;
        RECT 39.130 7.650 39.300 7.820 ;
        RECT 39.580 7.650 39.750 7.820 ;
        RECT 40.030 7.650 40.200 7.820 ;
        RECT 40.880 7.650 41.050 7.820 ;
        RECT 41.330 7.650 41.500 7.820 ;
        RECT 41.780 7.650 41.950 7.820 ;
        RECT 42.230 7.650 42.400 7.820 ;
        RECT 42.680 7.650 42.850 7.820 ;
        RECT 43.130 7.650 43.300 7.820 ;
        RECT 43.580 7.650 43.750 7.820 ;
        RECT 44.030 7.650 44.200 7.820 ;
        RECT 44.480 7.650 44.650 7.820 ;
        RECT 44.930 7.650 45.100 7.820 ;
        RECT 45.380 7.650 45.550 7.820 ;
        RECT 45.830 7.650 46.000 7.820 ;
        RECT 46.280 7.650 46.450 7.820 ;
        RECT 46.730 7.650 46.900 7.820 ;
        RECT 47.580 7.650 47.750 7.820 ;
        RECT 48.030 7.650 48.200 7.820 ;
        RECT 48.480 7.650 48.650 7.820 ;
        RECT 48.930 7.650 49.100 7.820 ;
        RECT 49.380 7.650 49.550 7.820 ;
        RECT 49.830 7.650 50.000 7.820 ;
        RECT 50.280 7.650 50.450 7.820 ;
        RECT 50.730 7.650 50.900 7.820 ;
        RECT 51.180 7.650 51.350 7.820 ;
        RECT 51.630 7.650 51.800 7.820 ;
        RECT 52.080 7.650 52.250 7.820 ;
        RECT 52.530 7.650 52.700 7.820 ;
        RECT 52.980 7.650 53.150 7.820 ;
        RECT 53.430 7.650 53.600 7.820 ;
      LAYER met1 ;
        RECT 0.580 7.500 53.920 7.850 ;
    END
  END Collector
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER li1 ;
        RECT 0.450 9.250 54.050 9.550 ;
      LAYER mcon ;
        RECT 1.300 9.250 1.600 9.550 ;
        RECT 2.300 9.250 2.600 9.550 ;
        RECT 3.300 9.250 3.600 9.550 ;
        RECT 4.300 9.250 4.600 9.550 ;
        RECT 5.300 9.250 5.600 9.550 ;
        RECT 6.300 9.250 6.600 9.550 ;
        RECT 7.300 9.250 7.600 9.550 ;
        RECT 8.300 9.250 8.600 9.550 ;
        RECT 9.300 9.250 9.600 9.550 ;
        RECT 10.300 9.250 10.600 9.550 ;
        RECT 11.300 9.250 11.600 9.550 ;
        RECT 12.300 9.250 12.600 9.550 ;
        RECT 13.300 9.250 13.600 9.550 ;
        RECT 14.300 9.250 14.600 9.550 ;
        RECT 15.300 9.250 15.600 9.550 ;
        RECT 16.300 9.250 16.600 9.550 ;
        RECT 17.300 9.250 17.600 9.550 ;
        RECT 18.300 9.250 18.600 9.550 ;
        RECT 19.300 9.250 19.600 9.550 ;
        RECT 20.300 9.250 20.600 9.550 ;
        RECT 21.300 9.250 21.600 9.550 ;
        RECT 22.300 9.250 22.600 9.550 ;
        RECT 23.300 9.250 23.600 9.550 ;
        RECT 24.300 9.250 24.600 9.550 ;
        RECT 25.300 9.250 25.600 9.550 ;
        RECT 26.300 9.250 26.600 9.550 ;
        RECT 27.300 9.250 27.600 9.550 ;
        RECT 28.300 9.250 28.600 9.550 ;
        RECT 29.300 9.250 29.600 9.550 ;
        RECT 30.300 9.250 30.600 9.550 ;
        RECT 31.300 9.250 31.600 9.550 ;
        RECT 32.300 9.250 32.600 9.550 ;
        RECT 33.300 9.250 33.600 9.550 ;
        RECT 34.300 9.250 34.600 9.550 ;
        RECT 35.300 9.250 35.600 9.550 ;
        RECT 36.300 9.250 36.600 9.550 ;
        RECT 37.300 9.250 37.600 9.550 ;
        RECT 38.300 9.250 38.600 9.550 ;
        RECT 39.300 9.250 39.600 9.550 ;
        RECT 40.300 9.250 40.600 9.550 ;
        RECT 41.300 9.250 41.600 9.550 ;
        RECT 42.300 9.250 42.600 9.550 ;
        RECT 43.300 9.250 43.600 9.550 ;
        RECT 44.300 9.250 44.600 9.550 ;
        RECT 45.300 9.250 45.600 9.550 ;
        RECT 46.300 9.250 46.600 9.550 ;
        RECT 47.300 9.250 47.600 9.550 ;
        RECT 48.300 9.250 48.600 9.550 ;
        RECT 49.300 9.250 49.600 9.550 ;
        RECT 50.300 9.250 50.600 9.550 ;
        RECT 51.300 9.250 51.600 9.550 ;
        RECT 52.300 9.250 52.600 9.550 ;
        RECT 53.300 9.250 53.600 9.550 ;
      LAYER met1 ;
        RECT 0.450 9.100 54.050 9.700 ;
    END
  END VPWR
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER li1 ;
        RECT 0.450 -0.150 54.050 0.150 ;
      LAYER mcon ;
        RECT 1.300 -0.150 1.600 0.150 ;
        RECT 2.300 -0.150 2.600 0.150 ;
        RECT 3.300 -0.150 3.600 0.150 ;
        RECT 4.300 -0.150 4.600 0.150 ;
        RECT 5.300 -0.150 5.600 0.150 ;
        RECT 6.300 -0.150 6.600 0.150 ;
        RECT 7.300 -0.150 7.600 0.150 ;
        RECT 8.300 -0.150 8.600 0.150 ;
        RECT 9.300 -0.150 9.600 0.150 ;
        RECT 10.300 -0.150 10.600 0.150 ;
        RECT 11.300 -0.150 11.600 0.150 ;
        RECT 12.300 -0.150 12.600 0.150 ;
        RECT 13.300 -0.150 13.600 0.150 ;
        RECT 14.300 -0.150 14.600 0.150 ;
        RECT 15.300 -0.150 15.600 0.150 ;
        RECT 16.300 -0.150 16.600 0.150 ;
        RECT 17.300 -0.150 17.600 0.150 ;
        RECT 18.300 -0.150 18.600 0.150 ;
        RECT 19.300 -0.150 19.600 0.150 ;
        RECT 20.300 -0.150 20.600 0.150 ;
        RECT 21.300 -0.150 21.600 0.150 ;
        RECT 22.300 -0.150 22.600 0.150 ;
        RECT 23.300 -0.150 23.600 0.150 ;
        RECT 24.300 -0.150 24.600 0.150 ;
        RECT 25.300 -0.150 25.600 0.150 ;
        RECT 26.300 -0.150 26.600 0.150 ;
        RECT 27.300 -0.150 27.600 0.150 ;
        RECT 28.300 -0.150 28.600 0.150 ;
        RECT 29.300 -0.150 29.600 0.150 ;
        RECT 30.300 -0.150 30.600 0.150 ;
        RECT 31.300 -0.150 31.600 0.150 ;
        RECT 32.300 -0.150 32.600 0.150 ;
        RECT 33.300 -0.150 33.600 0.150 ;
        RECT 34.300 -0.150 34.600 0.150 ;
        RECT 35.300 -0.150 35.600 0.150 ;
        RECT 36.300 -0.150 36.600 0.150 ;
        RECT 37.300 -0.150 37.600 0.150 ;
        RECT 38.300 -0.150 38.600 0.150 ;
        RECT 39.300 -0.150 39.600 0.150 ;
        RECT 40.300 -0.150 40.600 0.150 ;
        RECT 41.300 -0.150 41.600 0.150 ;
        RECT 42.300 -0.150 42.600 0.150 ;
        RECT 43.300 -0.150 43.600 0.150 ;
        RECT 44.300 -0.150 44.600 0.150 ;
        RECT 45.300 -0.150 45.600 0.150 ;
        RECT 46.300 -0.150 46.600 0.150 ;
        RECT 47.300 -0.150 47.600 0.150 ;
        RECT 48.300 -0.150 48.600 0.150 ;
        RECT 49.300 -0.150 49.600 0.150 ;
        RECT 50.300 -0.150 50.600 0.150 ;
        RECT 51.300 -0.150 51.600 0.150 ;
        RECT 52.300 -0.150 52.600 0.150 ;
        RECT 53.300 -0.150 53.600 0.150 ;
      LAYER met1 ;
        RECT 0.450 -0.300 54.050 0.300 ;
    END
  END VGND
END sky130_asc_pnp_05v5_W3p40L3p40_8

#--------EOF---------

MACRO sky130_asc_nfet_01v8_lvt_1
  CLASS CORE ;
  FOREIGN sky130_asc_nfet_01v8_lvt_1 ;
  ORIGIN 0.000 0.000 ;
  SIZE 3.970 BY 9.400 ;
  SITE unitasc ;
  PIN GATE
    DIRECTION INOUT ;
    ANTENNAGATEAREA 8.000000 ;
    PORT
      LAYER li1 ;
        RECT 1.340 0.720 3.520 1.020 ;
    END
  END GATE
  PIN SOURCE
    DIRECTION INOUT ;
    ANTENNADIFFAREA 1.160000 ;
    PORT
      LAYER li1 ;
        RECT 0.940 8.450 3.520 8.750 ;
        RECT 3.285 7.020 3.455 8.450 ;
        RECT 3.285 6.930 3.460 7.020 ;
        RECT 3.290 2.980 3.460 6.930 ;
      LAYER mcon ;
        RECT 3.290 3.060 3.460 6.940 ;
      LAYER met1 ;
        RECT 3.260 3.000 3.490 7.000 ;
    END
  END SOURCE
  PIN DRAIN
    DIRECTION INOUT ;
    ANTENNADIFFAREA 1.160000 ;
    PORT
      LAYER li1 ;
        RECT 1.000 3.270 1.170 7.020 ;
        RECT 0.995 2.980 1.170 3.270 ;
        RECT 0.995 2.150 1.165 2.980 ;
        RECT 0.940 1.850 3.520 2.150 ;
      LAYER mcon ;
        RECT 1.000 3.060 1.170 6.940 ;
      LAYER met1 ;
        RECT 0.970 3.000 1.200 7.000 ;
    END
  END DRAIN
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER li1 ;
        RECT 0.450 9.250 3.520 9.550 ;
      LAYER mcon ;
        RECT 1.790 9.250 2.090 9.550 ;
      LAYER met1 ;
        RECT 0.450 9.100 3.520 9.700 ;
    END
  END VPWR
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.450 0.150 3.520 7.130 ;
      LAYER li1 ;
        RECT 0.590 0.150 0.890 1.200 ;
        RECT 0.450 -0.150 3.520 0.150 ;
      LAYER mcon ;
        RECT 1.790 -0.150 2.090 0.150 ;
      LAYER met1 ;
        RECT 0.450 -0.300 3.520 0.300 ;
    END
  END VGND
END sky130_asc_nfet_01v8_lvt_1

#--------EOF---------

MACRO sky130_asc_pfet_01v8_lvt_1
  CLASS CORE ;
  FOREIGN sky130_asc_pfet_01v8_lvt_1 ;
  ORIGIN 0.000 0.000 ;
  SIZE 4.330 BY 9.400 ;
  SITE unitasc ;
  PIN GATE
    DIRECTION INOUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 12.900000 ;
    PORT
      LAYER li1 ;
        RECT 0.940 0.520 3.880 0.820 ;
    END
  END GATE
  PIN SOURCE
    DIRECTION INOUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.870500 ;
    PORT
      LAYER li1 ;
        RECT 1.240 8.450 3.880 8.650 ;
        RECT 3.465 8.245 3.635 8.450 ;
        RECT 3.465 8.130 3.640 8.245 ;
        RECT 3.470 1.755 3.640 8.130 ;
      LAYER mcon ;
        RECT 3.470 1.835 3.640 8.165 ;
      LAYER met1 ;
        RECT 3.440 1.775 3.670 8.225 ;
    END
  END SOURCE
  PIN DRAIN
    DIRECTION INOUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.870500 ;
    PORT
      LAYER li1 ;
        RECT 1.180 1.870 1.350 8.245 ;
        RECT 1.175 1.755 1.350 1.870 ;
        RECT 1.175 1.350 1.345 1.755 ;
        RECT 0.940 1.050 3.880 1.350 ;
      LAYER mcon ;
        RECT 1.180 1.835 1.350 8.165 ;
      LAYER met1 ;
        RECT 1.150 1.775 1.380 8.225 ;
    END
  END DRAIN
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT 0.450 1.470 3.880 9.700 ;
        RECT 0.940 1.465 3.880 1.470 ;
      LAYER li1 ;
        RECT 0.450 9.250 3.880 9.550 ;
        RECT 0.590 8.200 0.890 9.250 ;
      LAYER mcon ;
        RECT 1.790 9.250 2.090 9.550 ;
      LAYER met1 ;
        RECT 0.450 9.100 3.880 9.700 ;
    END
  END VPWR
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER li1 ;
        RECT 0.450 -0.150 3.880 0.150 ;
      LAYER mcon ;
        RECT 1.790 -0.150 2.090 0.150 ;
      LAYER met1 ;
        RECT 0.450 -0.300 3.880 0.300 ;
    END
  END VGND
END sky130_asc_pfet_01v8_lvt_1

#--------EOF---------

MACRO sky130_asc_res_xhigh_po_2p85_1
  CLASS CORE ;
  FOREIGN sky130_asc_res_xhigh_po_2p85_1 ;
  ORIGIN 0.000 0.000 ;
  SIZE 13.600 BY 9.400 ;
  SITE unitasc ;
  PIN Rin
    DIRECTION INOUT ;
    PORT
      LAYER li1 ;
        RECT 0.700 5.375 2.860 8.225 ;
      LAYER mcon ;
        RECT 0.790 5.455 2.775 8.145 ;
      LAYER met1 ;
        RECT 0.755 5.395 2.805 8.205 ;
    END
  END Rin
  PIN Rout
    DIRECTION INOUT ;
    PORT
      LAYER li1 ;
        RECT 0.700 0.575 2.860 3.425 ;
      LAYER mcon ;
        RECT 0.790 0.655 2.775 3.345 ;
      LAYER met1 ;
        RECT 0.755 0.595 2.805 3.405 ;
    END
  END Rout
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER li1 ;
        RECT 0.700 9.250 12.900 9.550 ;
      LAYER mcon ;
        RECT 1.550 9.250 1.850 9.550 ;
        RECT 2.550 9.250 2.850 9.550 ;
        RECT 3.550 9.250 3.850 9.550 ;
        RECT 4.550 9.250 4.850 9.550 ;
        RECT 5.550 9.250 5.850 9.550 ;
        RECT 6.550 9.250 6.850 9.550 ;
        RECT 7.550 9.250 7.850 9.550 ;
        RECT 8.550 9.250 8.850 9.550 ;
        RECT 9.550 9.250 9.850 9.550 ;
        RECT 10.550 9.250 10.850 9.550 ;
        RECT 11.550 9.250 11.850 9.550 ;
      LAYER met1 ;
        RECT 0.700 9.100 12.900 9.700 ;
    END
  END VPWR
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.700 -0.300 12.900 8.250 ;
      LAYER li1 ;
        RECT 5.260 0.150 8.340 4.850 ;
        RECT 0.700 -0.150 12.900 0.150 ;
      LAYER mcon ;
        RECT 1.550 -0.150 1.850 0.150 ;
        RECT 2.550 -0.150 2.850 0.150 ;
        RECT 3.550 -0.150 3.850 0.150 ;
        RECT 4.550 -0.150 4.850 0.150 ;
        RECT 5.550 -0.150 5.850 0.150 ;
        RECT 6.550 -0.150 6.850 0.150 ;
        RECT 7.550 -0.150 7.850 0.150 ;
        RECT 8.550 -0.150 8.850 0.150 ;
        RECT 9.550 -0.150 9.850 0.150 ;
        RECT 10.550 -0.150 10.850 0.150 ;
        RECT 11.550 -0.150 11.850 0.150 ;
      LAYER met1 ;
        RECT 0.700 -0.300 12.900 0.300 ;
    END
  END VGND
  OBS
      LAYER li1 ;
        RECT 10.740 0.575 12.900 8.225 ;
      LAYER mcon ;
        RECT 10.825 5.455 12.810 8.145 ;
        RECT 10.825 0.655 12.810 3.345 ;
      LAYER met1 ;
        RECT 10.795 5.395 12.845 8.205 ;
        RECT 10.740 0.575 12.900 5.395 ;
  END
END sky130_asc_res_xhigh_po_2p85_1

#--------EOF---------

MACRO sky130_asc_pfet_01v8_lvt_60
  CLASS CORE ;
  FOREIGN sky130_asc_pfet_01v8_lvt_60 ;
  ORIGIN 0.000 0.000 ;
  SIZE 139.435 BY 9.400 ;
  SITE unitasc ;
  PIN GATE
    DIRECTION INOUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 774.000000 ;
    PORT
      LAYER li1 ;
        RECT 0.940 0.520 138.980 0.820 ;
    END
  END GATE
  PIN SOURCE
    DIRECTION INOUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 56.114998 ;
    PORT
      LAYER li1 ;
        RECT 1.240 8.450 138.980 8.650 ;
        RECT 3.465 1.755 3.635 8.450 ;
        RECT 8.045 1.755 8.215 8.450 ;
        RECT 12.625 1.755 12.795 8.450 ;
        RECT 17.205 1.755 17.375 8.450 ;
        RECT 21.785 1.755 21.955 8.450 ;
        RECT 26.365 1.755 26.535 8.450 ;
        RECT 30.945 1.755 31.115 8.450 ;
        RECT 35.525 1.755 35.695 8.450 ;
        RECT 40.105 1.755 40.275 8.450 ;
        RECT 44.685 1.755 44.855 8.450 ;
        RECT 49.265 1.755 49.435 8.450 ;
        RECT 53.845 1.755 54.015 8.450 ;
        RECT 58.425 1.755 58.595 8.450 ;
        RECT 63.005 1.755 63.175 8.450 ;
        RECT 67.585 1.755 67.755 8.450 ;
        RECT 72.165 1.755 72.335 8.450 ;
        RECT 76.745 1.755 76.915 8.450 ;
        RECT 81.325 1.755 81.495 8.450 ;
        RECT 85.905 1.755 86.075 8.450 ;
        RECT 90.485 1.755 90.655 8.450 ;
        RECT 95.065 1.755 95.235 8.450 ;
        RECT 99.645 1.755 99.815 8.450 ;
        RECT 104.225 1.755 104.395 8.450 ;
        RECT 108.805 1.755 108.975 8.450 ;
        RECT 113.385 1.755 113.555 8.450 ;
        RECT 117.965 1.755 118.135 8.450 ;
        RECT 122.545 1.755 122.715 8.450 ;
        RECT 127.125 1.755 127.295 8.450 ;
        RECT 131.705 1.755 131.875 8.450 ;
        RECT 136.285 1.755 136.455 8.450 ;
      LAYER mcon ;
        RECT 3.465 1.835 3.635 8.165 ;
        RECT 8.045 1.835 8.215 8.165 ;
        RECT 12.625 1.835 12.795 8.165 ;
        RECT 17.205 1.835 17.375 8.165 ;
        RECT 21.785 1.835 21.955 8.165 ;
        RECT 26.365 1.835 26.535 8.165 ;
        RECT 30.945 1.835 31.115 8.165 ;
        RECT 35.525 1.835 35.695 8.165 ;
        RECT 40.105 1.835 40.275 8.165 ;
        RECT 44.685 1.835 44.855 8.165 ;
        RECT 49.265 1.835 49.435 8.165 ;
        RECT 53.845 1.835 54.015 8.165 ;
        RECT 58.425 1.835 58.595 8.165 ;
        RECT 63.005 1.835 63.175 8.165 ;
        RECT 67.585 1.835 67.755 8.165 ;
        RECT 72.165 1.835 72.335 8.165 ;
        RECT 76.745 1.835 76.915 8.165 ;
        RECT 81.325 1.835 81.495 8.165 ;
        RECT 85.905 1.835 86.075 8.165 ;
        RECT 90.485 1.835 90.655 8.165 ;
        RECT 95.065 1.835 95.235 8.165 ;
        RECT 99.645 1.835 99.815 8.165 ;
        RECT 104.225 1.835 104.395 8.165 ;
        RECT 108.805 1.835 108.975 8.165 ;
        RECT 113.385 1.835 113.555 8.165 ;
        RECT 117.965 1.835 118.135 8.165 ;
        RECT 122.545 1.835 122.715 8.165 ;
        RECT 127.125 1.835 127.295 8.165 ;
        RECT 131.705 1.835 131.875 8.165 ;
        RECT 136.285 1.835 136.455 8.165 ;
      LAYER met1 ;
        RECT 3.435 1.775 3.665 8.225 ;
        RECT 8.015 1.775 8.245 8.225 ;
        RECT 12.595 1.775 12.825 8.225 ;
        RECT 17.175 1.775 17.405 8.225 ;
        RECT 21.755 1.775 21.985 8.225 ;
        RECT 26.335 1.775 26.565 8.225 ;
        RECT 30.915 1.775 31.145 8.225 ;
        RECT 35.495 1.775 35.725 8.225 ;
        RECT 40.075 1.775 40.305 8.225 ;
        RECT 44.655 1.775 44.885 8.225 ;
        RECT 49.235 1.775 49.465 8.225 ;
        RECT 53.815 1.775 54.045 8.225 ;
        RECT 58.395 1.775 58.625 8.225 ;
        RECT 62.975 1.775 63.205 8.225 ;
        RECT 67.555 1.775 67.785 8.225 ;
        RECT 72.135 1.775 72.365 8.225 ;
        RECT 76.715 1.775 76.945 8.225 ;
        RECT 81.295 1.775 81.525 8.225 ;
        RECT 85.875 1.775 86.105 8.225 ;
        RECT 90.455 1.775 90.685 8.225 ;
        RECT 95.035 1.775 95.265 8.225 ;
        RECT 99.615 1.775 99.845 8.225 ;
        RECT 104.195 1.775 104.425 8.225 ;
        RECT 108.775 1.775 109.005 8.225 ;
        RECT 113.355 1.775 113.585 8.225 ;
        RECT 117.935 1.775 118.165 8.225 ;
        RECT 122.515 1.775 122.745 8.225 ;
        RECT 127.095 1.775 127.325 8.225 ;
        RECT 131.675 1.775 131.905 8.225 ;
        RECT 136.255 1.775 136.485 8.225 ;
    END
  END SOURCE
  PIN DRAIN
    DIRECTION INOUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 57.985500 ;
    PORT
      LAYER li1 ;
        RECT 1.175 1.350 1.345 8.245 ;
        RECT 5.755 1.350 5.925 8.245 ;
        RECT 10.335 1.350 10.505 8.245 ;
        RECT 14.915 1.350 15.085 8.245 ;
        RECT 19.495 1.350 19.665 8.245 ;
        RECT 24.075 1.350 24.245 8.245 ;
        RECT 28.655 1.350 28.825 8.245 ;
        RECT 33.235 1.350 33.405 8.245 ;
        RECT 37.815 1.350 37.985 8.245 ;
        RECT 42.395 1.350 42.565 8.245 ;
        RECT 46.975 1.350 47.145 8.245 ;
        RECT 51.555 1.350 51.725 8.245 ;
        RECT 56.135 1.350 56.305 8.245 ;
        RECT 60.715 1.350 60.885 8.245 ;
        RECT 65.295 1.350 65.465 8.245 ;
        RECT 69.875 1.350 70.045 8.245 ;
        RECT 74.455 1.350 74.625 8.245 ;
        RECT 79.035 1.350 79.205 8.245 ;
        RECT 83.615 1.350 83.785 8.245 ;
        RECT 88.195 1.350 88.365 8.245 ;
        RECT 92.775 1.350 92.945 8.245 ;
        RECT 97.355 1.350 97.525 8.245 ;
        RECT 101.935 1.350 102.105 8.245 ;
        RECT 106.515 1.350 106.685 8.245 ;
        RECT 111.095 1.350 111.265 8.245 ;
        RECT 115.675 1.350 115.845 8.245 ;
        RECT 120.255 1.350 120.425 8.245 ;
        RECT 124.835 1.350 125.005 8.245 ;
        RECT 129.415 1.350 129.585 8.245 ;
        RECT 133.995 1.350 134.165 8.245 ;
        RECT 138.575 1.350 138.745 8.245 ;
        RECT 0.940 1.050 138.980 1.350 ;
      LAYER mcon ;
        RECT 1.175 1.835 1.345 8.165 ;
        RECT 5.755 1.835 5.925 8.165 ;
        RECT 10.335 1.835 10.505 8.165 ;
        RECT 14.915 1.835 15.085 8.165 ;
        RECT 19.495 1.835 19.665 8.165 ;
        RECT 24.075 1.835 24.245 8.165 ;
        RECT 28.655 1.835 28.825 8.165 ;
        RECT 33.235 1.835 33.405 8.165 ;
        RECT 37.815 1.835 37.985 8.165 ;
        RECT 42.395 1.835 42.565 8.165 ;
        RECT 46.975 1.835 47.145 8.165 ;
        RECT 51.555 1.835 51.725 8.165 ;
        RECT 56.135 1.835 56.305 8.165 ;
        RECT 60.715 1.835 60.885 8.165 ;
        RECT 65.295 1.835 65.465 8.165 ;
        RECT 69.875 1.835 70.045 8.165 ;
        RECT 74.455 1.835 74.625 8.165 ;
        RECT 79.035 1.835 79.205 8.165 ;
        RECT 83.615 1.835 83.785 8.165 ;
        RECT 88.195 1.835 88.365 8.165 ;
        RECT 92.775 1.835 92.945 8.165 ;
        RECT 97.355 1.835 97.525 8.165 ;
        RECT 101.935 1.835 102.105 8.165 ;
        RECT 106.515 1.835 106.685 8.165 ;
        RECT 111.095 1.835 111.265 8.165 ;
        RECT 115.675 1.835 115.845 8.165 ;
        RECT 120.255 1.835 120.425 8.165 ;
        RECT 124.835 1.835 125.005 8.165 ;
        RECT 129.415 1.835 129.585 8.165 ;
        RECT 133.995 1.835 134.165 8.165 ;
        RECT 138.575 1.835 138.745 8.165 ;
      LAYER met1 ;
        RECT 1.145 1.775 1.375 8.225 ;
        RECT 5.725 1.775 5.955 8.225 ;
        RECT 10.305 1.775 10.535 8.225 ;
        RECT 14.885 1.775 15.115 8.225 ;
        RECT 19.465 1.775 19.695 8.225 ;
        RECT 24.045 1.775 24.275 8.225 ;
        RECT 28.625 1.775 28.855 8.225 ;
        RECT 33.205 1.775 33.435 8.225 ;
        RECT 37.785 1.775 38.015 8.225 ;
        RECT 42.365 1.775 42.595 8.225 ;
        RECT 46.945 1.775 47.175 8.225 ;
        RECT 51.525 1.775 51.755 8.225 ;
        RECT 56.105 1.775 56.335 8.225 ;
        RECT 60.685 1.775 60.915 8.225 ;
        RECT 65.265 1.775 65.495 8.225 ;
        RECT 69.845 1.775 70.075 8.225 ;
        RECT 74.425 1.775 74.655 8.225 ;
        RECT 79.005 1.775 79.235 8.225 ;
        RECT 83.585 1.775 83.815 8.225 ;
        RECT 88.165 1.775 88.395 8.225 ;
        RECT 92.745 1.775 92.975 8.225 ;
        RECT 97.325 1.775 97.555 8.225 ;
        RECT 101.905 1.775 102.135 8.225 ;
        RECT 106.485 1.775 106.715 8.225 ;
        RECT 111.065 1.775 111.295 8.225 ;
        RECT 115.645 1.775 115.875 8.225 ;
        RECT 120.225 1.775 120.455 8.225 ;
        RECT 124.805 1.775 125.035 8.225 ;
        RECT 129.385 1.775 129.615 8.225 ;
        RECT 133.965 1.775 134.195 8.225 ;
        RECT 138.545 1.775 138.775 8.225 ;
    END
  END DRAIN
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT 0.450 8.535 138.980 9.700 ;
        RECT 0.450 1.470 138.985 8.535 ;
        RECT 0.935 1.465 138.985 1.470 ;
      LAYER li1 ;
        RECT 0.450 9.250 138.980 9.550 ;
        RECT 0.590 8.200 0.890 9.250 ;
        RECT 5.830 8.850 6.630 9.250 ;
        RECT 12.330 8.850 13.130 9.250 ;
        RECT 18.830 8.850 19.630 9.250 ;
        RECT 25.330 8.850 26.130 9.250 ;
        RECT 31.830 8.850 32.630 9.250 ;
        RECT 38.330 8.850 39.130 9.250 ;
        RECT 44.830 8.850 45.630 9.250 ;
        RECT 51.330 8.850 52.130 9.250 ;
        RECT 57.830 8.850 58.630 9.250 ;
        RECT 64.330 8.850 65.130 9.250 ;
        RECT 70.830 8.850 71.630 9.250 ;
        RECT 77.330 8.850 78.130 9.250 ;
        RECT 83.830 8.850 84.630 9.250 ;
        RECT 90.330 8.850 91.130 9.250 ;
        RECT 96.830 8.850 97.630 9.250 ;
        RECT 103.330 8.850 104.130 9.250 ;
        RECT 109.830 8.850 110.630 9.250 ;
        RECT 116.330 8.850 117.130 9.250 ;
        RECT 122.830 8.850 123.630 9.250 ;
        RECT 129.330 8.850 130.130 9.250 ;
      LAYER mcon ;
        RECT 1.790 9.250 2.090 9.550 ;
        RECT 3.790 9.250 4.090 9.550 ;
        RECT 5.790 9.250 6.090 9.550 ;
        RECT 7.790 9.250 8.090 9.550 ;
        RECT 9.790 9.250 10.090 9.550 ;
        RECT 11.790 9.250 12.090 9.550 ;
        RECT 13.790 9.250 14.090 9.550 ;
        RECT 15.790 9.250 16.090 9.550 ;
        RECT 17.790 9.250 18.090 9.550 ;
        RECT 19.790 9.250 20.090 9.550 ;
        RECT 21.790 9.250 22.090 9.550 ;
        RECT 23.790 9.250 24.090 9.550 ;
        RECT 25.790 9.250 26.090 9.550 ;
        RECT 27.790 9.250 28.090 9.550 ;
        RECT 29.790 9.250 30.090 9.550 ;
        RECT 31.790 9.250 32.090 9.550 ;
        RECT 33.790 9.250 34.090 9.550 ;
        RECT 35.790 9.250 36.090 9.550 ;
        RECT 37.790 9.250 38.090 9.550 ;
        RECT 39.790 9.250 40.090 9.550 ;
        RECT 41.790 9.250 42.090 9.550 ;
        RECT 43.790 9.250 44.090 9.550 ;
        RECT 45.790 9.250 46.090 9.550 ;
        RECT 47.790 9.250 48.090 9.550 ;
        RECT 49.790 9.250 50.090 9.550 ;
        RECT 51.790 9.250 52.090 9.550 ;
        RECT 53.790 9.250 54.090 9.550 ;
        RECT 55.790 9.250 56.090 9.550 ;
        RECT 57.790 9.250 58.090 9.550 ;
        RECT 59.790 9.250 60.090 9.550 ;
        RECT 61.790 9.250 62.090 9.550 ;
        RECT 63.790 9.250 64.090 9.550 ;
        RECT 65.790 9.250 66.090 9.550 ;
        RECT 67.790 9.250 68.090 9.550 ;
        RECT 69.790 9.250 70.090 9.550 ;
        RECT 71.790 9.250 72.090 9.550 ;
        RECT 73.790 9.250 74.090 9.550 ;
        RECT 75.790 9.250 76.090 9.550 ;
        RECT 77.790 9.250 78.090 9.550 ;
        RECT 79.790 9.250 80.090 9.550 ;
        RECT 81.790 9.250 82.090 9.550 ;
        RECT 83.790 9.250 84.090 9.550 ;
        RECT 85.790 9.250 86.090 9.550 ;
        RECT 87.790 9.250 88.090 9.550 ;
        RECT 89.790 9.250 90.090 9.550 ;
        RECT 91.790 9.250 92.090 9.550 ;
        RECT 93.790 9.250 94.090 9.550 ;
        RECT 95.790 9.250 96.090 9.550 ;
        RECT 97.790 9.250 98.090 9.550 ;
        RECT 99.790 9.250 100.090 9.550 ;
        RECT 101.790 9.250 102.090 9.550 ;
        RECT 103.790 9.250 104.090 9.550 ;
        RECT 105.790 9.250 106.090 9.550 ;
        RECT 107.790 9.250 108.090 9.550 ;
        RECT 109.790 9.250 110.090 9.550 ;
        RECT 111.790 9.250 112.090 9.550 ;
        RECT 113.790 9.250 114.090 9.550 ;
        RECT 115.790 9.250 116.090 9.550 ;
        RECT 117.790 9.250 118.090 9.550 ;
        RECT 119.790 9.250 120.090 9.550 ;
        RECT 121.790 9.250 122.090 9.550 ;
        RECT 123.790 9.250 124.090 9.550 ;
        RECT 125.790 9.250 126.090 9.550 ;
        RECT 127.790 9.250 128.090 9.550 ;
        RECT 129.790 9.250 130.090 9.550 ;
        RECT 131.790 9.250 132.090 9.550 ;
        RECT 133.790 9.250 134.090 9.550 ;
        RECT 135.790 9.250 136.090 9.550 ;
        RECT 137.790 9.250 138.090 9.550 ;
      LAYER met1 ;
        RECT 0.450 9.100 138.980 9.700 ;
    END
  END VPWR
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER li1 ;
        RECT 0.450 -0.150 138.980 0.150 ;
      LAYER mcon ;
        RECT 1.790 -0.150 2.090 0.150 ;
        RECT 3.790 -0.150 4.090 0.150 ;
        RECT 5.790 -0.150 6.090 0.150 ;
        RECT 7.790 -0.150 8.090 0.150 ;
        RECT 9.790 -0.150 10.090 0.150 ;
        RECT 11.790 -0.150 12.090 0.150 ;
        RECT 13.790 -0.150 14.090 0.150 ;
        RECT 15.790 -0.150 16.090 0.150 ;
        RECT 17.790 -0.150 18.090 0.150 ;
        RECT 19.790 -0.150 20.090 0.150 ;
        RECT 21.790 -0.150 22.090 0.150 ;
        RECT 23.790 -0.150 24.090 0.150 ;
        RECT 25.790 -0.150 26.090 0.150 ;
        RECT 27.790 -0.150 28.090 0.150 ;
        RECT 29.790 -0.150 30.090 0.150 ;
        RECT 31.790 -0.150 32.090 0.150 ;
        RECT 33.790 -0.150 34.090 0.150 ;
        RECT 35.790 -0.150 36.090 0.150 ;
        RECT 37.790 -0.150 38.090 0.150 ;
        RECT 39.790 -0.150 40.090 0.150 ;
        RECT 41.790 -0.150 42.090 0.150 ;
        RECT 43.790 -0.150 44.090 0.150 ;
        RECT 45.790 -0.150 46.090 0.150 ;
        RECT 47.790 -0.150 48.090 0.150 ;
        RECT 49.790 -0.150 50.090 0.150 ;
        RECT 51.790 -0.150 52.090 0.150 ;
        RECT 53.790 -0.150 54.090 0.150 ;
        RECT 55.790 -0.150 56.090 0.150 ;
        RECT 57.790 -0.150 58.090 0.150 ;
        RECT 59.790 -0.150 60.090 0.150 ;
        RECT 61.790 -0.150 62.090 0.150 ;
        RECT 63.790 -0.150 64.090 0.150 ;
        RECT 65.790 -0.150 66.090 0.150 ;
        RECT 67.790 -0.150 68.090 0.150 ;
        RECT 69.790 -0.150 70.090 0.150 ;
        RECT 71.790 -0.150 72.090 0.150 ;
        RECT 73.790 -0.150 74.090 0.150 ;
        RECT 75.790 -0.150 76.090 0.150 ;
        RECT 77.790 -0.150 78.090 0.150 ;
        RECT 79.790 -0.150 80.090 0.150 ;
        RECT 81.790 -0.150 82.090 0.150 ;
        RECT 83.790 -0.150 84.090 0.150 ;
        RECT 85.790 -0.150 86.090 0.150 ;
        RECT 87.790 -0.150 88.090 0.150 ;
        RECT 89.790 -0.150 90.090 0.150 ;
        RECT 91.790 -0.150 92.090 0.150 ;
        RECT 93.790 -0.150 94.090 0.150 ;
        RECT 95.790 -0.150 96.090 0.150 ;
        RECT 97.790 -0.150 98.090 0.150 ;
        RECT 99.790 -0.150 100.090 0.150 ;
        RECT 101.790 -0.150 102.090 0.150 ;
        RECT 103.790 -0.150 104.090 0.150 ;
        RECT 105.790 -0.150 106.090 0.150 ;
        RECT 107.790 -0.150 108.090 0.150 ;
        RECT 109.790 -0.150 110.090 0.150 ;
        RECT 111.790 -0.150 112.090 0.150 ;
        RECT 113.790 -0.150 114.090 0.150 ;
        RECT 115.790 -0.150 116.090 0.150 ;
        RECT 117.790 -0.150 118.090 0.150 ;
        RECT 119.790 -0.150 120.090 0.150 ;
        RECT 121.790 -0.150 122.090 0.150 ;
        RECT 123.790 -0.150 124.090 0.150 ;
        RECT 125.790 -0.150 126.090 0.150 ;
        RECT 127.790 -0.150 128.090 0.150 ;
        RECT 129.790 -0.150 130.090 0.150 ;
        RECT 131.790 -0.150 132.090 0.150 ;
        RECT 133.790 -0.150 134.090 0.150 ;
        RECT 135.790 -0.150 136.090 0.150 ;
        RECT 137.790 -0.150 138.090 0.150 ;
      LAYER met1 ;
        RECT 0.450 -0.300 138.980 0.300 ;
    END
  END VGND
END sky130_asc_pfet_01v8_lvt_60

#--------EOF---------

MACRO sky130_asc_res_xhigh_po_2p85_2
  CLASS CORE ;
  FOREIGN sky130_asc_res_xhigh_po_2p85_2 ;
  ORIGIN 0.000 0.000 ;
  SIZE 16.470 BY 9.400 ;
  SITE unitasc ;
  PIN Rin
    DIRECTION INOUT ;
    PORT
      LAYER li1 ;
        RECT 0.705 5.375 2.865 8.225 ;
      LAYER mcon ;
        RECT 0.795 5.455 2.780 8.145 ;
      LAYER met1 ;
        RECT 0.760 5.395 2.810 8.205 ;
    END
  END Rin
  PIN Rout
    DIRECTION INOUT ;
    PORT
      LAYER li1 ;
        RECT 0.705 0.575 2.865 3.425 ;
      LAYER mcon ;
        RECT 0.795 0.655 2.780 3.345 ;
      LAYER met1 ;
        RECT 0.760 0.595 2.810 3.405 ;
    END
  END Rout
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER li1 ;
        RECT 0.710 9.250 15.770 9.550 ;
      LAYER mcon ;
        RECT 1.560 9.250 1.860 9.550 ;
        RECT 2.560 9.250 2.860 9.550 ;
        RECT 3.560 9.250 3.860 9.550 ;
        RECT 4.560 9.250 4.860 9.550 ;
        RECT 5.560 9.250 5.860 9.550 ;
        RECT 6.560 9.250 6.860 9.550 ;
        RECT 7.560 9.250 7.860 9.550 ;
        RECT 8.560 9.250 8.860 9.550 ;
        RECT 9.560 9.250 9.860 9.550 ;
        RECT 10.560 9.250 10.860 9.550 ;
        RECT 11.560 9.250 11.860 9.550 ;
        RECT 12.560 9.250 12.860 9.550 ;
        RECT 13.560 9.250 13.860 9.550 ;
        RECT 14.560 9.250 14.860 9.550 ;
      LAYER met1 ;
        RECT 0.710 9.100 15.770 9.700 ;
    END
  END VPWR
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 2.140 -0.300 14.340 8.250 ;
      LAYER li1 ;
        RECT 6.700 0.150 9.780 4.850 ;
        RECT 0.710 -0.150 15.770 0.150 ;
      LAYER mcon ;
        RECT 1.560 -0.150 1.860 0.150 ;
        RECT 2.560 -0.150 2.860 0.150 ;
        RECT 3.560 -0.150 3.860 0.150 ;
        RECT 4.560 -0.150 4.860 0.150 ;
        RECT 5.560 -0.150 5.860 0.150 ;
        RECT 6.560 -0.150 6.860 0.150 ;
        RECT 7.560 -0.150 7.860 0.150 ;
        RECT 8.560 -0.150 8.860 0.150 ;
        RECT 9.560 -0.150 9.860 0.150 ;
        RECT 10.560 -0.150 10.860 0.150 ;
        RECT 11.560 -0.150 11.860 0.150 ;
        RECT 12.560 -0.150 12.860 0.150 ;
        RECT 13.560 -0.150 13.860 0.150 ;
        RECT 14.560 -0.150 14.860 0.150 ;
      LAYER met1 ;
        RECT 0.710 -0.300 15.770 0.300 ;
    END
  END VGND
  OBS
      LAYER li1 ;
        RECT 13.615 0.575 15.775 8.225 ;
      LAYER mcon ;
        RECT 13.700 5.455 15.685 8.145 ;
        RECT 13.700 0.655 15.685 3.345 ;
      LAYER met1 ;
        RECT 13.670 5.395 15.720 8.205 ;
        RECT 13.615 0.575 15.775 5.395 ;
  END
END sky130_asc_res_xhigh_po_2p85_2

#--------EOF---------

MACRO sky130_asc_pnp_05v5_W3p40L3p40_1
  CLASS CORE ;
  FOREIGN sky130_asc_pnp_05v5_W3p40L3p40_1 ;
  ORIGIN 0.000 0.000 ;
  SIZE 7.600 BY 9.400 ;
  SITE unitasc ;
  PIN Emitter
    DIRECTION INOUT ;
    ANTENNADIFFAREA 11.559999 ;
    PORT
      LAYER li1 ;
        RECT 2.065 2.965 5.535 6.435 ;
      LAYER mcon ;
        RECT 2.430 5.830 2.600 6.000 ;
        RECT 2.930 5.830 3.100 6.000 ;
        RECT 3.430 5.830 3.600 6.000 ;
        RECT 3.930 5.830 4.100 6.000 ;
        RECT 4.430 5.830 4.600 6.000 ;
        RECT 4.930 5.830 5.100 6.000 ;
        RECT 2.430 5.330 2.600 5.500 ;
        RECT 2.930 5.330 3.100 5.500 ;
        RECT 3.430 5.330 3.600 5.500 ;
        RECT 3.930 5.330 4.100 5.500 ;
        RECT 4.430 5.330 4.600 5.500 ;
        RECT 4.930 5.330 5.100 5.500 ;
        RECT 2.430 4.830 2.600 5.000 ;
        RECT 2.930 4.830 3.100 5.000 ;
        RECT 3.430 4.830 3.600 5.000 ;
        RECT 3.930 4.830 4.100 5.000 ;
        RECT 4.430 4.830 4.600 5.000 ;
        RECT 4.930 4.830 5.100 5.000 ;
        RECT 2.430 4.330 2.600 4.500 ;
        RECT 2.930 4.330 3.100 4.500 ;
        RECT 3.430 4.330 3.600 4.500 ;
        RECT 3.930 4.330 4.100 4.500 ;
        RECT 4.430 4.330 4.600 4.500 ;
        RECT 4.930 4.330 5.100 4.500 ;
        RECT 2.430 3.830 2.600 4.000 ;
        RECT 2.930 3.830 3.100 4.000 ;
        RECT 3.430 3.830 3.600 4.000 ;
        RECT 3.930 3.830 4.100 4.000 ;
        RECT 4.430 3.830 4.600 4.000 ;
        RECT 4.930 3.830 5.100 4.000 ;
        RECT 2.430 3.330 2.600 3.500 ;
        RECT 2.930 3.330 3.100 3.500 ;
        RECT 3.430 3.330 3.600 3.500 ;
        RECT 3.930 3.330 4.100 3.500 ;
        RECT 4.430 3.330 4.600 3.500 ;
        RECT 4.930 3.330 5.100 3.500 ;
      LAYER met1 ;
        RECT 2.275 3.175 5.325 6.225 ;
    END
  END Emitter
  PIN Base
    DIRECTION INOUT ;
    ANTENNAGATEAREA 26.728899 ;
    ANTENNADIFFAREA 6.408000 ;
    PORT
      LAYER li1 ;
        RECT 1.395 6.745 6.205 7.105 ;
        RECT 1.395 2.655 1.755 6.745 ;
        RECT 5.845 2.655 6.205 6.745 ;
        RECT 1.395 2.295 6.205 2.655 ;
    END
  END Base
  PIN Collector
    DIRECTION INOUT ;
    ANTENNADIFFAREA 11.988700 ;
    PORT
      LAYER pwell ;
        RECT 0.450 7.285 7.150 8.050 ;
        RECT 0.450 2.115 1.215 7.285 ;
        RECT 6.385 2.115 7.150 7.285 ;
        RECT 0.450 1.350 7.150 2.115 ;
      LAYER li1 ;
        RECT 0.580 7.425 7.020 7.920 ;
        RECT 0.580 1.975 1.075 7.425 ;
        RECT 6.525 1.975 7.020 7.425 ;
        RECT 0.580 1.480 7.020 1.975 ;
    END
  END Collector
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER li1 ;
        RECT 0.450 9.250 7.150 9.550 ;
      LAYER mcon ;
        RECT 1.300 9.250 1.600 9.550 ;
        RECT 2.300 9.250 2.600 9.550 ;
        RECT 3.300 9.250 3.600 9.550 ;
        RECT 4.300 9.250 4.600 9.550 ;
        RECT 5.300 9.250 5.600 9.550 ;
        RECT 6.300 9.250 6.600 9.550 ;
      LAYER met1 ;
        RECT 0.450 9.100 7.150 9.700 ;
    END
  END VPWR
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER li1 ;
        RECT 0.450 -0.150 7.150 0.150 ;
      LAYER mcon ;
        RECT 1.300 -0.150 1.600 0.150 ;
        RECT 2.300 -0.150 2.600 0.150 ;
        RECT 3.300 -0.150 3.600 0.150 ;
        RECT 4.300 -0.150 4.600 0.150 ;
        RECT 5.300 -0.150 5.600 0.150 ;
        RECT 6.300 -0.150 6.600 0.150 ;
      LAYER met1 ;
        RECT 0.450 -0.300 7.150 0.300 ;
    END
  END VGND
END sky130_asc_pnp_05v5_W3p40L3p40_1

#--------EOF---------

MACRO sky130_asc_pfet_01v8_lvt_12
  CLASS CORE ;
  FOREIGN sky130_asc_pfet_01v8_lvt_12 ;
  ORIGIN 0.000 0.000 ;
  SIZE 29.515 BY 9.400 ;
  SITE unitasc ;
  PIN GATE
    DIRECTION INOUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 154.800003 ;
    PORT
      LAYER li1 ;
        RECT 0.940 0.520 29.060 0.820 ;
    END
  END GATE
  PIN SOURCE
    DIRECTION INOUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 11.223000 ;
    PORT
      LAYER li1 ;
        RECT 1.240 8.450 29.060 8.650 ;
        RECT 3.465 1.755 3.635 8.450 ;
        RECT 8.045 1.755 8.215 8.450 ;
        RECT 12.625 1.755 12.795 8.450 ;
        RECT 17.205 1.755 17.375 8.450 ;
        RECT 21.785 1.755 21.955 8.450 ;
        RECT 26.365 1.755 26.535 8.450 ;
      LAYER mcon ;
        RECT 3.465 1.835 3.635 8.165 ;
        RECT 8.045 1.835 8.215 8.165 ;
        RECT 12.625 1.835 12.795 8.165 ;
        RECT 17.205 1.835 17.375 8.165 ;
        RECT 21.785 1.835 21.955 8.165 ;
        RECT 26.365 1.835 26.535 8.165 ;
      LAYER met1 ;
        RECT 3.435 1.775 3.665 8.225 ;
        RECT 8.015 1.775 8.245 8.225 ;
        RECT 12.595 1.775 12.825 8.225 ;
        RECT 17.175 1.775 17.405 8.225 ;
        RECT 21.755 1.775 21.985 8.225 ;
        RECT 26.335 1.775 26.565 8.225 ;
    END
  END SOURCE
  PIN DRAIN
    DIRECTION INOUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 13.093500 ;
    PORT
      LAYER li1 ;
        RECT 1.175 1.350 1.345 8.245 ;
        RECT 5.755 1.350 5.925 8.245 ;
        RECT 10.335 1.350 10.505 8.245 ;
        RECT 14.915 1.350 15.085 8.245 ;
        RECT 19.495 1.350 19.665 8.245 ;
        RECT 24.075 1.350 24.245 8.245 ;
        RECT 28.655 1.350 28.825 8.245 ;
        RECT 0.940 1.050 29.060 1.350 ;
      LAYER mcon ;
        RECT 1.175 1.835 1.345 8.165 ;
        RECT 5.755 1.835 5.925 8.165 ;
        RECT 10.335 1.835 10.505 8.165 ;
        RECT 14.915 1.835 15.085 8.165 ;
        RECT 19.495 1.835 19.665 8.165 ;
        RECT 24.075 1.835 24.245 8.165 ;
        RECT 28.655 1.835 28.825 8.165 ;
      LAYER met1 ;
        RECT 1.145 1.775 1.375 8.225 ;
        RECT 5.725 1.775 5.955 8.225 ;
        RECT 10.305 1.775 10.535 8.225 ;
        RECT 14.885 1.775 15.115 8.225 ;
        RECT 19.465 1.775 19.695 8.225 ;
        RECT 24.045 1.775 24.275 8.225 ;
        RECT 28.625 1.775 28.855 8.225 ;
    END
  END DRAIN
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT 0.450 8.535 29.060 9.700 ;
        RECT 0.450 1.470 29.065 8.535 ;
        RECT 0.935 1.465 29.065 1.470 ;
      LAYER li1 ;
        RECT 0.450 9.250 29.060 9.550 ;
        RECT 0.590 8.200 0.890 9.250 ;
        RECT 5.830 8.850 6.630 9.250 ;
        RECT 12.330 8.850 13.130 9.250 ;
        RECT 18.830 8.850 19.630 9.250 ;
      LAYER mcon ;
        RECT 1.790 9.250 2.090 9.550 ;
        RECT 3.790 9.250 4.090 9.550 ;
        RECT 5.790 9.250 6.090 9.550 ;
        RECT 7.790 9.250 8.090 9.550 ;
        RECT 9.790 9.250 10.090 9.550 ;
        RECT 11.790 9.250 12.090 9.550 ;
        RECT 13.790 9.250 14.090 9.550 ;
        RECT 15.790 9.250 16.090 9.550 ;
        RECT 17.790 9.250 18.090 9.550 ;
        RECT 19.790 9.250 20.090 9.550 ;
        RECT 21.790 9.250 22.090 9.550 ;
        RECT 23.790 9.250 24.090 9.550 ;
        RECT 25.790 9.250 26.090 9.550 ;
        RECT 27.790 9.250 28.090 9.550 ;
      LAYER met1 ;
        RECT 0.450 9.100 29.060 9.700 ;
    END
  END VPWR
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER li1 ;
        RECT 0.450 -0.150 29.060 0.150 ;
      LAYER mcon ;
        RECT 1.790 -0.150 2.090 0.150 ;
        RECT 3.790 -0.150 4.090 0.150 ;
        RECT 5.790 -0.150 6.090 0.150 ;
        RECT 7.790 -0.150 8.090 0.150 ;
        RECT 9.790 -0.150 10.090 0.150 ;
        RECT 11.790 -0.150 12.090 0.150 ;
        RECT 13.790 -0.150 14.090 0.150 ;
        RECT 15.790 -0.150 16.090 0.150 ;
        RECT 17.790 -0.150 18.090 0.150 ;
        RECT 19.790 -0.150 20.090 0.150 ;
        RECT 21.790 -0.150 22.090 0.150 ;
        RECT 23.790 -0.150 24.090 0.150 ;
        RECT 25.790 -0.150 26.090 0.150 ;
        RECT 27.790 -0.150 28.090 0.150 ;
      LAYER met1 ;
        RECT 0.450 -0.300 29.060 0.300 ;
    END
  END VGND
END sky130_asc_pfet_01v8_lvt_12

#--------EOF---------

MACRO sky130_asc_pfet_01v8_lvt_6
  CLASS CORE ;
  FOREIGN sky130_asc_pfet_01v8_lvt_6 ;
  ORIGIN 0.000 0.000 ;
  SIZE 15.775 BY 9.400 ;
  SITE unitasc ;
  PIN GATE
    DIRECTION INOUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 77.400002 ;
    PORT
      LAYER li1 ;
        RECT 0.940 0.520 15.320 0.820 ;
    END
  END GATE
  PIN SOURCE
    DIRECTION INOUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 5.611500 ;
    PORT
      LAYER li1 ;
        RECT 1.240 8.450 15.320 8.650 ;
        RECT 3.465 1.755 3.635 8.450 ;
        RECT 8.045 1.755 8.215 8.450 ;
        RECT 12.625 1.755 12.795 8.450 ;
      LAYER mcon ;
        RECT 3.465 1.835 3.635 8.165 ;
        RECT 8.045 1.835 8.215 8.165 ;
        RECT 12.625 1.835 12.795 8.165 ;
      LAYER met1 ;
        RECT 3.435 1.775 3.665 8.225 ;
        RECT 8.015 1.775 8.245 8.225 ;
        RECT 12.595 1.775 12.825 8.225 ;
    END
  END SOURCE
  PIN DRAIN
    DIRECTION INOUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 7.482000 ;
    PORT
      LAYER li1 ;
        RECT 1.175 1.350 1.345 8.245 ;
        RECT 5.755 1.350 5.925 8.245 ;
        RECT 10.335 1.350 10.505 8.245 ;
        RECT 14.915 1.350 15.085 8.245 ;
        RECT 0.940 1.050 15.320 1.350 ;
      LAYER mcon ;
        RECT 1.175 1.835 1.345 8.165 ;
        RECT 5.755 1.835 5.925 8.165 ;
        RECT 10.335 1.835 10.505 8.165 ;
        RECT 14.915 1.835 15.085 8.165 ;
      LAYER met1 ;
        RECT 1.145 1.775 1.375 8.225 ;
        RECT 5.725 1.775 5.955 8.225 ;
        RECT 10.305 1.775 10.535 8.225 ;
        RECT 14.885 1.775 15.115 8.225 ;
    END
  END DRAIN
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT 0.450 8.535 15.320 9.700 ;
        RECT 0.450 1.470 15.325 8.535 ;
        RECT 0.935 1.465 15.325 1.470 ;
      LAYER li1 ;
        RECT 0.450 9.250 15.320 9.550 ;
        RECT 0.590 8.200 0.890 9.250 ;
        RECT 5.830 8.850 6.630 9.250 ;
      LAYER mcon ;
        RECT 1.790 9.250 2.090 9.550 ;
        RECT 3.790 9.250 4.090 9.550 ;
        RECT 5.790 9.250 6.090 9.550 ;
        RECT 7.790 9.250 8.090 9.550 ;
        RECT 9.790 9.250 10.090 9.550 ;
        RECT 11.790 9.250 12.090 9.550 ;
        RECT 13.790 9.250 14.090 9.550 ;
      LAYER met1 ;
        RECT 0.450 9.100 15.320 9.700 ;
    END
  END VPWR
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER li1 ;
        RECT 0.450 -0.150 15.320 0.150 ;
      LAYER mcon ;
        RECT 1.790 -0.150 2.090 0.150 ;
        RECT 3.790 -0.150 4.090 0.150 ;
        RECT 5.790 -0.150 6.090 0.150 ;
        RECT 7.790 -0.150 8.090 0.150 ;
        RECT 9.790 -0.150 10.090 0.150 ;
        RECT 11.790 -0.150 12.090 0.150 ;
        RECT 13.790 -0.150 14.090 0.150 ;
      LAYER met1 ;
        RECT 0.450 -0.300 15.320 0.300 ;
    END
  END VGND
END sky130_asc_pfet_01v8_lvt_6

#--------EOF---------

MACRO sky130_asc_pnp_05v5_W3p40L3p40_7
  CLASS CORE ;
  FOREIGN sky130_asc_pnp_05v5_W3p40L3p40_7 ;
  ORIGIN 0.000 0.000 ;
  SIZE 47.800 BY 9.400 ;
  SITE unitasc ;
  PIN Emitter
    DIRECTION INOUT ;
    ANTENNADIFFAREA 80.919998 ;
    PORT
      LAYER li1 ;
        RECT 2.065 2.965 5.535 6.435 ;
        RECT 8.765 2.965 12.235 6.435 ;
        RECT 15.465 2.965 18.935 6.435 ;
        RECT 22.165 2.965 25.635 6.435 ;
        RECT 28.865 2.965 32.335 6.435 ;
        RECT 35.565 2.965 39.035 6.435 ;
        RECT 42.265 2.965 45.735 6.435 ;
      LAYER mcon ;
        RECT 2.430 5.830 2.600 6.000 ;
        RECT 2.930 5.830 3.100 6.000 ;
        RECT 3.430 5.830 3.600 6.000 ;
        RECT 3.930 5.830 4.100 6.000 ;
        RECT 4.430 5.830 4.600 6.000 ;
        RECT 4.930 5.830 5.100 6.000 ;
        RECT 2.430 5.330 2.600 5.500 ;
        RECT 2.930 5.330 3.100 5.500 ;
        RECT 3.430 5.330 3.600 5.500 ;
        RECT 3.930 5.330 4.100 5.500 ;
        RECT 4.430 5.330 4.600 5.500 ;
        RECT 4.930 5.330 5.100 5.500 ;
        RECT 2.430 4.830 2.600 5.000 ;
        RECT 2.930 4.830 3.100 5.000 ;
        RECT 3.430 4.830 3.600 5.000 ;
        RECT 3.930 4.830 4.100 5.000 ;
        RECT 4.430 4.830 4.600 5.000 ;
        RECT 4.930 4.830 5.100 5.000 ;
        RECT 2.430 4.330 2.600 4.500 ;
        RECT 2.930 4.330 3.100 4.500 ;
        RECT 3.430 4.330 3.600 4.500 ;
        RECT 3.930 4.330 4.100 4.500 ;
        RECT 4.430 4.330 4.600 4.500 ;
        RECT 4.930 4.330 5.100 4.500 ;
        RECT 2.430 3.830 2.600 4.000 ;
        RECT 2.930 3.830 3.100 4.000 ;
        RECT 3.430 3.830 3.600 4.000 ;
        RECT 3.930 3.830 4.100 4.000 ;
        RECT 4.430 3.830 4.600 4.000 ;
        RECT 4.930 3.830 5.100 4.000 ;
        RECT 2.430 3.330 2.600 3.500 ;
        RECT 2.930 3.330 3.100 3.500 ;
        RECT 3.430 3.330 3.600 3.500 ;
        RECT 3.930 3.330 4.100 3.500 ;
        RECT 4.430 3.330 4.600 3.500 ;
        RECT 4.930 3.330 5.100 3.500 ;
        RECT 9.130 5.830 9.300 6.000 ;
        RECT 9.630 5.830 9.800 6.000 ;
        RECT 10.130 5.830 10.300 6.000 ;
        RECT 10.630 5.830 10.800 6.000 ;
        RECT 11.130 5.830 11.300 6.000 ;
        RECT 11.630 5.830 11.800 6.000 ;
        RECT 9.130 5.330 9.300 5.500 ;
        RECT 9.630 5.330 9.800 5.500 ;
        RECT 10.130 5.330 10.300 5.500 ;
        RECT 10.630 5.330 10.800 5.500 ;
        RECT 11.130 5.330 11.300 5.500 ;
        RECT 11.630 5.330 11.800 5.500 ;
        RECT 9.130 4.830 9.300 5.000 ;
        RECT 9.630 4.830 9.800 5.000 ;
        RECT 10.130 4.830 10.300 5.000 ;
        RECT 10.630 4.830 10.800 5.000 ;
        RECT 11.130 4.830 11.300 5.000 ;
        RECT 11.630 4.830 11.800 5.000 ;
        RECT 9.130 4.330 9.300 4.500 ;
        RECT 9.630 4.330 9.800 4.500 ;
        RECT 10.130 4.330 10.300 4.500 ;
        RECT 10.630 4.330 10.800 4.500 ;
        RECT 11.130 4.330 11.300 4.500 ;
        RECT 11.630 4.330 11.800 4.500 ;
        RECT 9.130 3.830 9.300 4.000 ;
        RECT 9.630 3.830 9.800 4.000 ;
        RECT 10.130 3.830 10.300 4.000 ;
        RECT 10.630 3.830 10.800 4.000 ;
        RECT 11.130 3.830 11.300 4.000 ;
        RECT 11.630 3.830 11.800 4.000 ;
        RECT 9.130 3.330 9.300 3.500 ;
        RECT 9.630 3.330 9.800 3.500 ;
        RECT 10.130 3.330 10.300 3.500 ;
        RECT 10.630 3.330 10.800 3.500 ;
        RECT 11.130 3.330 11.300 3.500 ;
        RECT 11.630 3.330 11.800 3.500 ;
        RECT 15.830 5.830 16.000 6.000 ;
        RECT 16.330 5.830 16.500 6.000 ;
        RECT 16.830 5.830 17.000 6.000 ;
        RECT 17.330 5.830 17.500 6.000 ;
        RECT 17.830 5.830 18.000 6.000 ;
        RECT 18.330 5.830 18.500 6.000 ;
        RECT 15.830 5.330 16.000 5.500 ;
        RECT 16.330 5.330 16.500 5.500 ;
        RECT 16.830 5.330 17.000 5.500 ;
        RECT 17.330 5.330 17.500 5.500 ;
        RECT 17.830 5.330 18.000 5.500 ;
        RECT 18.330 5.330 18.500 5.500 ;
        RECT 15.830 4.830 16.000 5.000 ;
        RECT 16.330 4.830 16.500 5.000 ;
        RECT 16.830 4.830 17.000 5.000 ;
        RECT 17.330 4.830 17.500 5.000 ;
        RECT 17.830 4.830 18.000 5.000 ;
        RECT 18.330 4.830 18.500 5.000 ;
        RECT 15.830 4.330 16.000 4.500 ;
        RECT 16.330 4.330 16.500 4.500 ;
        RECT 16.830 4.330 17.000 4.500 ;
        RECT 17.330 4.330 17.500 4.500 ;
        RECT 17.830 4.330 18.000 4.500 ;
        RECT 18.330 4.330 18.500 4.500 ;
        RECT 15.830 3.830 16.000 4.000 ;
        RECT 16.330 3.830 16.500 4.000 ;
        RECT 16.830 3.830 17.000 4.000 ;
        RECT 17.330 3.830 17.500 4.000 ;
        RECT 17.830 3.830 18.000 4.000 ;
        RECT 18.330 3.830 18.500 4.000 ;
        RECT 15.830 3.330 16.000 3.500 ;
        RECT 16.330 3.330 16.500 3.500 ;
        RECT 16.830 3.330 17.000 3.500 ;
        RECT 17.330 3.330 17.500 3.500 ;
        RECT 17.830 3.330 18.000 3.500 ;
        RECT 18.330 3.330 18.500 3.500 ;
        RECT 22.530 5.830 22.700 6.000 ;
        RECT 23.030 5.830 23.200 6.000 ;
        RECT 23.530 5.830 23.700 6.000 ;
        RECT 24.030 5.830 24.200 6.000 ;
        RECT 24.530 5.830 24.700 6.000 ;
        RECT 25.030 5.830 25.200 6.000 ;
        RECT 22.530 5.330 22.700 5.500 ;
        RECT 23.030 5.330 23.200 5.500 ;
        RECT 23.530 5.330 23.700 5.500 ;
        RECT 24.030 5.330 24.200 5.500 ;
        RECT 24.530 5.330 24.700 5.500 ;
        RECT 25.030 5.330 25.200 5.500 ;
        RECT 22.530 4.830 22.700 5.000 ;
        RECT 23.030 4.830 23.200 5.000 ;
        RECT 23.530 4.830 23.700 5.000 ;
        RECT 24.030 4.830 24.200 5.000 ;
        RECT 24.530 4.830 24.700 5.000 ;
        RECT 25.030 4.830 25.200 5.000 ;
        RECT 22.530 4.330 22.700 4.500 ;
        RECT 23.030 4.330 23.200 4.500 ;
        RECT 23.530 4.330 23.700 4.500 ;
        RECT 24.030 4.330 24.200 4.500 ;
        RECT 24.530 4.330 24.700 4.500 ;
        RECT 25.030 4.330 25.200 4.500 ;
        RECT 22.530 3.830 22.700 4.000 ;
        RECT 23.030 3.830 23.200 4.000 ;
        RECT 23.530 3.830 23.700 4.000 ;
        RECT 24.030 3.830 24.200 4.000 ;
        RECT 24.530 3.830 24.700 4.000 ;
        RECT 25.030 3.830 25.200 4.000 ;
        RECT 22.530 3.330 22.700 3.500 ;
        RECT 23.030 3.330 23.200 3.500 ;
        RECT 23.530 3.330 23.700 3.500 ;
        RECT 24.030 3.330 24.200 3.500 ;
        RECT 24.530 3.330 24.700 3.500 ;
        RECT 25.030 3.330 25.200 3.500 ;
        RECT 29.230 5.830 29.400 6.000 ;
        RECT 29.730 5.830 29.900 6.000 ;
        RECT 30.230 5.830 30.400 6.000 ;
        RECT 30.730 5.830 30.900 6.000 ;
        RECT 31.230 5.830 31.400 6.000 ;
        RECT 31.730 5.830 31.900 6.000 ;
        RECT 29.230 5.330 29.400 5.500 ;
        RECT 29.730 5.330 29.900 5.500 ;
        RECT 30.230 5.330 30.400 5.500 ;
        RECT 30.730 5.330 30.900 5.500 ;
        RECT 31.230 5.330 31.400 5.500 ;
        RECT 31.730 5.330 31.900 5.500 ;
        RECT 29.230 4.830 29.400 5.000 ;
        RECT 29.730 4.830 29.900 5.000 ;
        RECT 30.230 4.830 30.400 5.000 ;
        RECT 30.730 4.830 30.900 5.000 ;
        RECT 31.230 4.830 31.400 5.000 ;
        RECT 31.730 4.830 31.900 5.000 ;
        RECT 29.230 4.330 29.400 4.500 ;
        RECT 29.730 4.330 29.900 4.500 ;
        RECT 30.230 4.330 30.400 4.500 ;
        RECT 30.730 4.330 30.900 4.500 ;
        RECT 31.230 4.330 31.400 4.500 ;
        RECT 31.730 4.330 31.900 4.500 ;
        RECT 29.230 3.830 29.400 4.000 ;
        RECT 29.730 3.830 29.900 4.000 ;
        RECT 30.230 3.830 30.400 4.000 ;
        RECT 30.730 3.830 30.900 4.000 ;
        RECT 31.230 3.830 31.400 4.000 ;
        RECT 31.730 3.830 31.900 4.000 ;
        RECT 29.230 3.330 29.400 3.500 ;
        RECT 29.730 3.330 29.900 3.500 ;
        RECT 30.230 3.330 30.400 3.500 ;
        RECT 30.730 3.330 30.900 3.500 ;
        RECT 31.230 3.330 31.400 3.500 ;
        RECT 31.730 3.330 31.900 3.500 ;
        RECT 35.930 5.830 36.100 6.000 ;
        RECT 36.430 5.830 36.600 6.000 ;
        RECT 36.930 5.830 37.100 6.000 ;
        RECT 37.430 5.830 37.600 6.000 ;
        RECT 37.930 5.830 38.100 6.000 ;
        RECT 38.430 5.830 38.600 6.000 ;
        RECT 35.930 5.330 36.100 5.500 ;
        RECT 36.430 5.330 36.600 5.500 ;
        RECT 36.930 5.330 37.100 5.500 ;
        RECT 37.430 5.330 37.600 5.500 ;
        RECT 37.930 5.330 38.100 5.500 ;
        RECT 38.430 5.330 38.600 5.500 ;
        RECT 35.930 4.830 36.100 5.000 ;
        RECT 36.430 4.830 36.600 5.000 ;
        RECT 36.930 4.830 37.100 5.000 ;
        RECT 37.430 4.830 37.600 5.000 ;
        RECT 37.930 4.830 38.100 5.000 ;
        RECT 38.430 4.830 38.600 5.000 ;
        RECT 35.930 4.330 36.100 4.500 ;
        RECT 36.430 4.330 36.600 4.500 ;
        RECT 36.930 4.330 37.100 4.500 ;
        RECT 37.430 4.330 37.600 4.500 ;
        RECT 37.930 4.330 38.100 4.500 ;
        RECT 38.430 4.330 38.600 4.500 ;
        RECT 35.930 3.830 36.100 4.000 ;
        RECT 36.430 3.830 36.600 4.000 ;
        RECT 36.930 3.830 37.100 4.000 ;
        RECT 37.430 3.830 37.600 4.000 ;
        RECT 37.930 3.830 38.100 4.000 ;
        RECT 38.430 3.830 38.600 4.000 ;
        RECT 35.930 3.330 36.100 3.500 ;
        RECT 36.430 3.330 36.600 3.500 ;
        RECT 36.930 3.330 37.100 3.500 ;
        RECT 37.430 3.330 37.600 3.500 ;
        RECT 37.930 3.330 38.100 3.500 ;
        RECT 38.430 3.330 38.600 3.500 ;
        RECT 42.630 5.830 42.800 6.000 ;
        RECT 43.130 5.830 43.300 6.000 ;
        RECT 43.630 5.830 43.800 6.000 ;
        RECT 44.130 5.830 44.300 6.000 ;
        RECT 44.630 5.830 44.800 6.000 ;
        RECT 45.130 5.830 45.300 6.000 ;
        RECT 42.630 5.330 42.800 5.500 ;
        RECT 43.130 5.330 43.300 5.500 ;
        RECT 43.630 5.330 43.800 5.500 ;
        RECT 44.130 5.330 44.300 5.500 ;
        RECT 44.630 5.330 44.800 5.500 ;
        RECT 45.130 5.330 45.300 5.500 ;
        RECT 42.630 4.830 42.800 5.000 ;
        RECT 43.130 4.830 43.300 5.000 ;
        RECT 43.630 4.830 43.800 5.000 ;
        RECT 44.130 4.830 44.300 5.000 ;
        RECT 44.630 4.830 44.800 5.000 ;
        RECT 45.130 4.830 45.300 5.000 ;
        RECT 42.630 4.330 42.800 4.500 ;
        RECT 43.130 4.330 43.300 4.500 ;
        RECT 43.630 4.330 43.800 4.500 ;
        RECT 44.130 4.330 44.300 4.500 ;
        RECT 44.630 4.330 44.800 4.500 ;
        RECT 45.130 4.330 45.300 4.500 ;
        RECT 42.630 3.830 42.800 4.000 ;
        RECT 43.130 3.830 43.300 4.000 ;
        RECT 43.630 3.830 43.800 4.000 ;
        RECT 44.130 3.830 44.300 4.000 ;
        RECT 44.630 3.830 44.800 4.000 ;
        RECT 45.130 3.830 45.300 4.000 ;
        RECT 42.630 3.330 42.800 3.500 ;
        RECT 43.130 3.330 43.300 3.500 ;
        RECT 43.630 3.330 43.800 3.500 ;
        RECT 44.130 3.330 44.300 3.500 ;
        RECT 44.630 3.330 44.800 3.500 ;
        RECT 45.130 3.330 45.300 3.500 ;
      LAYER met1 ;
        RECT 2.270 3.170 45.530 6.230 ;
    END
  END Emitter
  PIN Base
    DIRECTION INOUT ;
    ANTENNAGATEAREA 187.102295 ;
    ANTENNADIFFAREA 44.855999 ;
    PORT
      LAYER li1 ;
        RECT 1.395 6.745 6.205 7.105 ;
        RECT 1.395 2.655 1.755 6.745 ;
        RECT 5.845 2.655 6.205 6.745 ;
        RECT 1.395 2.295 6.205 2.655 ;
        RECT 8.095 6.745 12.905 7.105 ;
        RECT 8.095 2.655 8.455 6.745 ;
        RECT 12.545 2.655 12.905 6.745 ;
        RECT 8.095 2.295 12.905 2.655 ;
        RECT 14.795 6.745 19.605 7.105 ;
        RECT 14.795 2.655 15.155 6.745 ;
        RECT 19.245 2.655 19.605 6.745 ;
        RECT 14.795 2.295 19.605 2.655 ;
        RECT 21.495 6.745 26.305 7.105 ;
        RECT 21.495 2.655 21.855 6.745 ;
        RECT 25.945 2.655 26.305 6.745 ;
        RECT 21.495 2.295 26.305 2.655 ;
        RECT 28.195 6.745 33.005 7.105 ;
        RECT 28.195 2.655 28.555 6.745 ;
        RECT 32.645 2.655 33.005 6.745 ;
        RECT 28.195 2.295 33.005 2.655 ;
        RECT 34.895 6.745 39.705 7.105 ;
        RECT 34.895 2.655 35.255 6.745 ;
        RECT 39.345 2.655 39.705 6.745 ;
        RECT 34.895 2.295 39.705 2.655 ;
        RECT 41.595 6.745 46.405 7.105 ;
        RECT 41.595 2.655 41.955 6.745 ;
        RECT 46.045 2.655 46.405 6.745 ;
        RECT 41.595 2.295 46.405 2.655 ;
      LAYER mcon ;
        RECT 1.500 6.850 1.670 7.020 ;
        RECT 1.950 6.850 2.120 7.020 ;
        RECT 2.400 6.850 2.570 7.020 ;
        RECT 2.850 6.850 3.020 7.020 ;
        RECT 3.300 6.850 3.470 7.020 ;
        RECT 3.750 6.850 3.920 7.020 ;
        RECT 4.200 6.850 4.370 7.020 ;
        RECT 4.650 6.850 4.820 7.020 ;
        RECT 5.100 6.850 5.270 7.020 ;
        RECT 5.550 6.850 5.720 7.020 ;
        RECT 6.000 6.850 6.170 7.020 ;
        RECT 8.200 6.850 8.370 7.020 ;
        RECT 8.650 6.850 8.820 7.020 ;
        RECT 9.100 6.850 9.270 7.020 ;
        RECT 9.550 6.850 9.720 7.020 ;
        RECT 10.000 6.850 10.170 7.020 ;
        RECT 10.450 6.850 10.620 7.020 ;
        RECT 10.900 6.850 11.070 7.020 ;
        RECT 11.350 6.850 11.520 7.020 ;
        RECT 11.800 6.850 11.970 7.020 ;
        RECT 12.250 6.850 12.420 7.020 ;
        RECT 12.700 6.850 12.870 7.020 ;
        RECT 14.900 6.850 15.070 7.020 ;
        RECT 15.350 6.850 15.520 7.020 ;
        RECT 15.800 6.850 15.970 7.020 ;
        RECT 16.250 6.850 16.420 7.020 ;
        RECT 16.700 6.850 16.870 7.020 ;
        RECT 17.150 6.850 17.320 7.020 ;
        RECT 17.600 6.850 17.770 7.020 ;
        RECT 18.050 6.850 18.220 7.020 ;
        RECT 18.500 6.850 18.670 7.020 ;
        RECT 18.950 6.850 19.120 7.020 ;
        RECT 19.400 6.850 19.570 7.020 ;
        RECT 21.600 6.850 21.770 7.020 ;
        RECT 22.050 6.850 22.220 7.020 ;
        RECT 22.500 6.850 22.670 7.020 ;
        RECT 22.950 6.850 23.120 7.020 ;
        RECT 23.400 6.850 23.570 7.020 ;
        RECT 23.850 6.850 24.020 7.020 ;
        RECT 24.300 6.850 24.470 7.020 ;
        RECT 24.750 6.850 24.920 7.020 ;
        RECT 25.200 6.850 25.370 7.020 ;
        RECT 25.650 6.850 25.820 7.020 ;
        RECT 26.100 6.850 26.270 7.020 ;
        RECT 28.300 6.850 28.470 7.020 ;
        RECT 28.750 6.850 28.920 7.020 ;
        RECT 29.200 6.850 29.370 7.020 ;
        RECT 29.650 6.850 29.820 7.020 ;
        RECT 30.100 6.850 30.270 7.020 ;
        RECT 30.550 6.850 30.720 7.020 ;
        RECT 31.000 6.850 31.170 7.020 ;
        RECT 31.450 6.850 31.620 7.020 ;
        RECT 31.900 6.850 32.070 7.020 ;
        RECT 32.350 6.850 32.520 7.020 ;
        RECT 32.800 6.850 32.970 7.020 ;
        RECT 35.000 6.850 35.170 7.020 ;
        RECT 35.450 6.850 35.620 7.020 ;
        RECT 35.900 6.850 36.070 7.020 ;
        RECT 36.350 6.850 36.520 7.020 ;
        RECT 36.800 6.850 36.970 7.020 ;
        RECT 37.250 6.850 37.420 7.020 ;
        RECT 37.700 6.850 37.870 7.020 ;
        RECT 38.150 6.850 38.320 7.020 ;
        RECT 38.600 6.850 38.770 7.020 ;
        RECT 39.050 6.850 39.220 7.020 ;
        RECT 39.500 6.850 39.670 7.020 ;
        RECT 41.700 6.850 41.870 7.020 ;
        RECT 42.150 6.850 42.320 7.020 ;
        RECT 42.600 6.850 42.770 7.020 ;
        RECT 43.050 6.850 43.220 7.020 ;
        RECT 43.500 6.850 43.670 7.020 ;
        RECT 43.950 6.850 44.120 7.020 ;
        RECT 44.400 6.850 44.570 7.020 ;
        RECT 44.850 6.850 45.020 7.020 ;
        RECT 45.300 6.850 45.470 7.020 ;
        RECT 45.750 6.850 45.920 7.020 ;
        RECT 46.200 6.850 46.370 7.020 ;
      LAYER met1 ;
        RECT 1.400 6.750 46.400 7.100 ;
    END
  END Base
  PIN Collector
    DIRECTION INOUT ;
    ANTENNADIFFAREA 93.967300 ;
    PORT
      LAYER pwell ;
        RECT 0.450 7.285 47.350 8.050 ;
        RECT 0.450 2.115 1.215 7.285 ;
        RECT 6.385 2.115 7.915 7.285 ;
        RECT 13.085 2.115 14.615 7.285 ;
        RECT 19.785 2.115 21.315 7.285 ;
        RECT 26.485 2.115 28.015 7.285 ;
        RECT 33.185 2.115 34.715 7.285 ;
        RECT 39.885 2.115 41.415 7.285 ;
        RECT 46.585 2.115 47.350 7.285 ;
        RECT 0.450 1.350 47.350 2.115 ;
      LAYER li1 ;
        RECT 0.580 7.425 47.220 7.920 ;
        RECT 0.580 1.975 1.075 7.425 ;
        RECT 6.525 1.975 7.775 7.425 ;
        RECT 13.225 1.975 14.475 7.425 ;
        RECT 19.925 1.975 21.175 7.425 ;
        RECT 26.625 1.975 27.875 7.425 ;
        RECT 33.325 1.975 34.575 7.425 ;
        RECT 40.025 1.975 41.275 7.425 ;
        RECT 46.725 1.975 47.220 7.425 ;
        RECT 0.580 1.480 47.220 1.975 ;
      LAYER mcon ;
        RECT 0.680 7.650 0.850 7.820 ;
        RECT 1.130 7.650 1.300 7.820 ;
        RECT 1.580 7.650 1.750 7.820 ;
        RECT 2.030 7.650 2.200 7.820 ;
        RECT 2.480 7.650 2.650 7.820 ;
        RECT 2.930 7.650 3.100 7.820 ;
        RECT 3.380 7.650 3.550 7.820 ;
        RECT 3.830 7.650 4.000 7.820 ;
        RECT 4.280 7.650 4.450 7.820 ;
        RECT 4.730 7.650 4.900 7.820 ;
        RECT 5.180 7.650 5.350 7.820 ;
        RECT 5.630 7.650 5.800 7.820 ;
        RECT 6.080 7.650 6.250 7.820 ;
        RECT 6.530 7.650 6.700 7.820 ;
        RECT 7.380 7.650 7.550 7.820 ;
        RECT 7.830 7.650 8.000 7.820 ;
        RECT 8.280 7.650 8.450 7.820 ;
        RECT 8.730 7.650 8.900 7.820 ;
        RECT 9.180 7.650 9.350 7.820 ;
        RECT 9.630 7.650 9.800 7.820 ;
        RECT 10.080 7.650 10.250 7.820 ;
        RECT 10.530 7.650 10.700 7.820 ;
        RECT 10.980 7.650 11.150 7.820 ;
        RECT 11.430 7.650 11.600 7.820 ;
        RECT 11.880 7.650 12.050 7.820 ;
        RECT 12.330 7.650 12.500 7.820 ;
        RECT 12.780 7.650 12.950 7.820 ;
        RECT 13.230 7.650 13.400 7.820 ;
        RECT 14.080 7.650 14.250 7.820 ;
        RECT 14.530 7.650 14.700 7.820 ;
        RECT 14.980 7.650 15.150 7.820 ;
        RECT 15.430 7.650 15.600 7.820 ;
        RECT 15.880 7.650 16.050 7.820 ;
        RECT 16.330 7.650 16.500 7.820 ;
        RECT 16.780 7.650 16.950 7.820 ;
        RECT 17.230 7.650 17.400 7.820 ;
        RECT 17.680 7.650 17.850 7.820 ;
        RECT 18.130 7.650 18.300 7.820 ;
        RECT 18.580 7.650 18.750 7.820 ;
        RECT 19.030 7.650 19.200 7.820 ;
        RECT 19.480 7.650 19.650 7.820 ;
        RECT 19.930 7.650 20.100 7.820 ;
        RECT 20.780 7.650 20.950 7.820 ;
        RECT 21.230 7.650 21.400 7.820 ;
        RECT 21.680 7.650 21.850 7.820 ;
        RECT 22.130 7.650 22.300 7.820 ;
        RECT 22.580 7.650 22.750 7.820 ;
        RECT 23.030 7.650 23.200 7.820 ;
        RECT 23.480 7.650 23.650 7.820 ;
        RECT 23.930 7.650 24.100 7.820 ;
        RECT 24.380 7.650 24.550 7.820 ;
        RECT 24.830 7.650 25.000 7.820 ;
        RECT 25.280 7.650 25.450 7.820 ;
        RECT 25.730 7.650 25.900 7.820 ;
        RECT 26.180 7.650 26.350 7.820 ;
        RECT 26.630 7.650 26.800 7.820 ;
        RECT 27.480 7.650 27.650 7.820 ;
        RECT 27.930 7.650 28.100 7.820 ;
        RECT 28.380 7.650 28.550 7.820 ;
        RECT 28.830 7.650 29.000 7.820 ;
        RECT 29.280 7.650 29.450 7.820 ;
        RECT 29.730 7.650 29.900 7.820 ;
        RECT 30.180 7.650 30.350 7.820 ;
        RECT 30.630 7.650 30.800 7.820 ;
        RECT 31.080 7.650 31.250 7.820 ;
        RECT 31.530 7.650 31.700 7.820 ;
        RECT 31.980 7.650 32.150 7.820 ;
        RECT 32.430 7.650 32.600 7.820 ;
        RECT 32.880 7.650 33.050 7.820 ;
        RECT 33.330 7.650 33.500 7.820 ;
        RECT 34.180 7.650 34.350 7.820 ;
        RECT 34.630 7.650 34.800 7.820 ;
        RECT 35.080 7.650 35.250 7.820 ;
        RECT 35.530 7.650 35.700 7.820 ;
        RECT 35.980 7.650 36.150 7.820 ;
        RECT 36.430 7.650 36.600 7.820 ;
        RECT 36.880 7.650 37.050 7.820 ;
        RECT 37.330 7.650 37.500 7.820 ;
        RECT 37.780 7.650 37.950 7.820 ;
        RECT 38.230 7.650 38.400 7.820 ;
        RECT 38.680 7.650 38.850 7.820 ;
        RECT 39.130 7.650 39.300 7.820 ;
        RECT 39.580 7.650 39.750 7.820 ;
        RECT 40.030 7.650 40.200 7.820 ;
        RECT 40.880 7.650 41.050 7.820 ;
        RECT 41.330 7.650 41.500 7.820 ;
        RECT 41.780 7.650 41.950 7.820 ;
        RECT 42.230 7.650 42.400 7.820 ;
        RECT 42.680 7.650 42.850 7.820 ;
        RECT 43.130 7.650 43.300 7.820 ;
        RECT 43.580 7.650 43.750 7.820 ;
        RECT 44.030 7.650 44.200 7.820 ;
        RECT 44.480 7.650 44.650 7.820 ;
        RECT 44.930 7.650 45.100 7.820 ;
        RECT 45.380 7.650 45.550 7.820 ;
        RECT 45.830 7.650 46.000 7.820 ;
        RECT 46.280 7.650 46.450 7.820 ;
        RECT 46.730 7.650 46.900 7.820 ;
      LAYER met1 ;
        RECT 0.580 7.500 47.220 7.850 ;
    END
  END Collector
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER li1 ;
        RECT 0.450 9.250 47.350 9.550 ;
      LAYER mcon ;
        RECT 1.300 9.250 1.600 9.550 ;
        RECT 2.300 9.250 2.600 9.550 ;
        RECT 3.300 9.250 3.600 9.550 ;
        RECT 4.300 9.250 4.600 9.550 ;
        RECT 5.300 9.250 5.600 9.550 ;
        RECT 6.300 9.250 6.600 9.550 ;
        RECT 7.300 9.250 7.600 9.550 ;
        RECT 8.300 9.250 8.600 9.550 ;
        RECT 9.300 9.250 9.600 9.550 ;
        RECT 10.300 9.250 10.600 9.550 ;
        RECT 11.300 9.250 11.600 9.550 ;
        RECT 12.300 9.250 12.600 9.550 ;
        RECT 13.300 9.250 13.600 9.550 ;
        RECT 14.300 9.250 14.600 9.550 ;
        RECT 15.300 9.250 15.600 9.550 ;
        RECT 16.300 9.250 16.600 9.550 ;
        RECT 17.300 9.250 17.600 9.550 ;
        RECT 18.300 9.250 18.600 9.550 ;
        RECT 19.300 9.250 19.600 9.550 ;
        RECT 20.300 9.250 20.600 9.550 ;
        RECT 21.300 9.250 21.600 9.550 ;
        RECT 22.300 9.250 22.600 9.550 ;
        RECT 23.300 9.250 23.600 9.550 ;
        RECT 24.300 9.250 24.600 9.550 ;
        RECT 25.300 9.250 25.600 9.550 ;
        RECT 26.300 9.250 26.600 9.550 ;
        RECT 27.300 9.250 27.600 9.550 ;
        RECT 28.300 9.250 28.600 9.550 ;
        RECT 29.300 9.250 29.600 9.550 ;
        RECT 30.300 9.250 30.600 9.550 ;
        RECT 31.300 9.250 31.600 9.550 ;
        RECT 32.300 9.250 32.600 9.550 ;
        RECT 33.300 9.250 33.600 9.550 ;
        RECT 34.300 9.250 34.600 9.550 ;
        RECT 35.300 9.250 35.600 9.550 ;
        RECT 36.300 9.250 36.600 9.550 ;
        RECT 37.300 9.250 37.600 9.550 ;
        RECT 38.300 9.250 38.600 9.550 ;
        RECT 39.300 9.250 39.600 9.550 ;
        RECT 40.300 9.250 40.600 9.550 ;
        RECT 41.300 9.250 41.600 9.550 ;
        RECT 42.300 9.250 42.600 9.550 ;
        RECT 43.300 9.250 43.600 9.550 ;
        RECT 44.300 9.250 44.600 9.550 ;
        RECT 45.300 9.250 45.600 9.550 ;
        RECT 46.300 9.250 46.600 9.550 ;
      LAYER met1 ;
        RECT 0.450 9.100 47.350 9.700 ;
    END
  END VPWR
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER li1 ;
        RECT 0.450 -0.150 47.350 0.150 ;
      LAYER mcon ;
        RECT 1.300 -0.150 1.600 0.150 ;
        RECT 2.300 -0.150 2.600 0.150 ;
        RECT 3.300 -0.150 3.600 0.150 ;
        RECT 4.300 -0.150 4.600 0.150 ;
        RECT 5.300 -0.150 5.600 0.150 ;
        RECT 6.300 -0.150 6.600 0.150 ;
        RECT 7.300 -0.150 7.600 0.150 ;
        RECT 8.300 -0.150 8.600 0.150 ;
        RECT 9.300 -0.150 9.600 0.150 ;
        RECT 10.300 -0.150 10.600 0.150 ;
        RECT 11.300 -0.150 11.600 0.150 ;
        RECT 12.300 -0.150 12.600 0.150 ;
        RECT 13.300 -0.150 13.600 0.150 ;
        RECT 14.300 -0.150 14.600 0.150 ;
        RECT 15.300 -0.150 15.600 0.150 ;
        RECT 16.300 -0.150 16.600 0.150 ;
        RECT 17.300 -0.150 17.600 0.150 ;
        RECT 18.300 -0.150 18.600 0.150 ;
        RECT 19.300 -0.150 19.600 0.150 ;
        RECT 20.300 -0.150 20.600 0.150 ;
        RECT 21.300 -0.150 21.600 0.150 ;
        RECT 22.300 -0.150 22.600 0.150 ;
        RECT 23.300 -0.150 23.600 0.150 ;
        RECT 24.300 -0.150 24.600 0.150 ;
        RECT 25.300 -0.150 25.600 0.150 ;
        RECT 26.300 -0.150 26.600 0.150 ;
        RECT 27.300 -0.150 27.600 0.150 ;
        RECT 28.300 -0.150 28.600 0.150 ;
        RECT 29.300 -0.150 29.600 0.150 ;
        RECT 30.300 -0.150 30.600 0.150 ;
        RECT 31.300 -0.150 31.600 0.150 ;
        RECT 32.300 -0.150 32.600 0.150 ;
        RECT 33.300 -0.150 33.600 0.150 ;
        RECT 34.300 -0.150 34.600 0.150 ;
        RECT 35.300 -0.150 35.600 0.150 ;
        RECT 36.300 -0.150 36.600 0.150 ;
        RECT 37.300 -0.150 37.600 0.150 ;
        RECT 38.300 -0.150 38.600 0.150 ;
        RECT 39.300 -0.150 39.600 0.150 ;
        RECT 40.300 -0.150 40.600 0.150 ;
        RECT 41.300 -0.150 41.600 0.150 ;
        RECT 42.300 -0.150 42.600 0.150 ;
        RECT 43.300 -0.150 43.600 0.150 ;
        RECT 44.300 -0.150 44.600 0.150 ;
        RECT 45.300 -0.150 45.600 0.150 ;
        RECT 46.300 -0.150 46.600 0.150 ;
      LAYER met1 ;
        RECT 0.450 -0.300 47.350 0.300 ;
    END
  END VGND
END sky130_asc_pnp_05v5_W3p40L3p40_7

#--------EOF---------

MACRO sky130_asc_cap_mim_m3_1
  CLASS CORE ;
  FOREIGN sky130_asc_cap_mim_m3_1 ;
  ORIGIN 0.000 0.000 ;
  SIZE 36.855 BY 9.400 ;
  SITE unitasc ;
  PIN Cin
    DIRECTION INOUT ;
    PORT
      LAYER met4 ;
        RECT 3.450 5.310 3.930 8.190 ;
        RECT 7.045 5.310 7.525 8.190 ;
        RECT 10.640 5.310 11.120 8.190 ;
        RECT 14.235 5.310 14.715 8.190 ;
        RECT 17.830 5.310 18.310 8.190 ;
        RECT 21.425 5.310 21.905 8.190 ;
        RECT 25.020 5.310 25.500 8.190 ;
        RECT 28.615 5.310 29.095 8.190 ;
        RECT 32.210 5.310 32.690 8.190 ;
        RECT 35.805 5.310 36.285 8.190 ;
        RECT 3.450 1.810 3.930 4.690 ;
        RECT 7.045 1.810 7.525 4.690 ;
        RECT 10.640 1.810 11.120 4.690 ;
        RECT 14.235 1.810 14.715 4.690 ;
        RECT 17.830 1.810 18.310 4.690 ;
        RECT 21.425 1.810 21.905 4.690 ;
        RECT 25.020 1.810 25.500 4.690 ;
        RECT 28.615 1.810 29.095 4.690 ;
        RECT 32.210 1.810 32.690 4.690 ;
        RECT 35.805 1.810 36.285 4.690 ;
    END
  END Cin
  PIN Cout
    DIRECTION INOUT ;
    PORT
      LAYER met4 ;
        RECT 1.150 7.555 2.750 7.650 ;
        RECT 4.750 7.555 6.350 7.650 ;
        RECT 8.350 7.555 9.950 7.650 ;
        RECT 11.950 7.555 13.550 7.650 ;
        RECT 15.550 7.555 17.150 7.650 ;
        RECT 19.150 7.555 20.750 7.650 ;
        RECT 22.750 7.555 24.350 7.650 ;
        RECT 26.350 7.555 27.950 7.650 ;
        RECT 29.950 7.555 31.550 7.650 ;
        RECT 33.550 7.555 35.150 7.650 ;
        RECT 1.150 5.945 2.760 7.555 ;
        RECT 4.745 5.945 6.355 7.555 ;
        RECT 8.340 5.945 9.950 7.555 ;
        RECT 11.935 5.945 13.550 7.555 ;
        RECT 15.530 5.945 17.150 7.555 ;
        RECT 19.125 5.945 20.750 7.555 ;
        RECT 22.720 5.945 24.350 7.555 ;
        RECT 26.315 5.945 27.950 7.555 ;
        RECT 29.910 5.945 31.550 7.555 ;
        RECT 33.505 5.945 35.150 7.555 ;
        RECT 1.150 4.055 2.750 5.945 ;
        RECT 4.750 4.055 6.350 5.945 ;
        RECT 8.350 4.055 9.950 5.945 ;
        RECT 11.950 4.055 13.550 5.945 ;
        RECT 15.550 4.055 17.150 5.945 ;
        RECT 19.150 4.055 20.750 5.945 ;
        RECT 22.750 4.055 24.350 5.945 ;
        RECT 26.350 4.055 27.950 5.945 ;
        RECT 29.950 4.055 31.550 5.945 ;
        RECT 33.550 4.055 35.150 5.945 ;
        RECT 1.150 2.445 2.760 4.055 ;
        RECT 4.745 2.445 6.355 4.055 ;
        RECT 8.340 2.445 9.950 4.055 ;
        RECT 11.935 2.445 13.550 4.055 ;
        RECT 15.530 2.445 17.150 4.055 ;
        RECT 19.125 2.445 20.750 4.055 ;
        RECT 22.720 2.445 24.350 4.055 ;
        RECT 26.315 2.445 27.950 4.055 ;
        RECT 29.910 2.445 31.550 4.055 ;
        RECT 33.505 2.445 35.150 4.055 ;
        RECT 1.150 1.450 2.750 2.445 ;
        RECT 4.750 1.450 6.350 2.445 ;
        RECT 8.350 1.450 9.950 2.445 ;
        RECT 11.950 1.450 13.550 2.445 ;
        RECT 15.550 1.450 17.150 2.445 ;
        RECT 19.150 1.450 20.750 2.445 ;
        RECT 22.750 1.450 24.350 2.445 ;
        RECT 26.350 1.450 27.950 2.445 ;
        RECT 29.950 1.450 31.550 2.445 ;
        RECT 33.550 1.450 35.150 2.445 ;
        RECT 0.460 0.750 36.300 1.450 ;
    END
  END Cout
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.460 9.100 36.300 9.700 ;
    END
  END VPWR
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.460 -0.300 36.300 0.300 ;
    END
  END VGND
  OBS
      LAYER li1 ;
        RECT 0.460 9.250 36.300 9.550 ;
        RECT 0.460 -0.150 36.300 0.150 ;
      LAYER mcon ;
        RECT 1.310 9.250 1.610 9.550 ;
        RECT 3.310 9.250 3.610 9.550 ;
        RECT 5.310 9.250 5.610 9.550 ;
        RECT 7.310 9.250 7.610 9.550 ;
        RECT 9.310 9.250 9.610 9.550 ;
        RECT 11.310 9.250 11.610 9.550 ;
        RECT 13.310 9.250 13.610 9.550 ;
        RECT 15.310 9.250 15.610 9.550 ;
        RECT 17.310 9.250 17.610 9.550 ;
        RECT 19.310 9.250 19.610 9.550 ;
        RECT 21.310 9.250 21.610 9.550 ;
        RECT 23.310 9.250 23.610 9.550 ;
        RECT 25.310 9.250 25.610 9.550 ;
        RECT 27.310 9.250 27.610 9.550 ;
        RECT 29.310 9.250 29.610 9.550 ;
        RECT 31.310 9.250 31.610 9.550 ;
        RECT 33.310 9.250 33.610 9.550 ;
        RECT 35.310 9.250 35.610 9.550 ;
        RECT 1.310 -0.150 1.610 0.150 ;
        RECT 3.310 -0.150 3.610 0.150 ;
        RECT 5.310 -0.150 5.610 0.150 ;
        RECT 7.310 -0.150 7.610 0.150 ;
        RECT 9.310 -0.150 9.610 0.150 ;
        RECT 11.310 -0.150 11.610 0.150 ;
        RECT 13.310 -0.150 13.610 0.150 ;
        RECT 15.310 -0.150 15.610 0.150 ;
        RECT 17.310 -0.150 17.610 0.150 ;
        RECT 19.310 -0.150 19.610 0.150 ;
        RECT 21.310 -0.150 21.610 0.150 ;
        RECT 23.310 -0.150 23.610 0.150 ;
        RECT 25.310 -0.150 25.610 0.150 ;
        RECT 27.310 -0.150 27.610 0.150 ;
        RECT 29.310 -0.150 29.610 0.150 ;
        RECT 31.310 -0.150 31.610 0.150 ;
        RECT 33.310 -0.150 33.610 0.150 ;
        RECT 35.310 -0.150 35.610 0.150 ;
      LAYER met2 ;
        RECT 0.450 7.850 1.450 8.250 ;
        RECT 0.560 0.800 1.360 1.300 ;
      LAYER via2 ;
        RECT 0.550 7.900 1.350 8.200 ;
        RECT 0.660 0.850 1.260 1.250 ;
      LAYER met3 ;
        RECT 0.450 1.750 36.310 8.250 ;
        RECT 0.460 0.750 1.460 1.350 ;
      LAYER via3 ;
        RECT 3.530 5.390 3.850 8.110 ;
        RECT 7.125 5.390 7.445 8.110 ;
        RECT 10.720 5.390 11.040 8.110 ;
        RECT 14.315 5.390 14.635 8.110 ;
        RECT 17.910 5.390 18.230 8.110 ;
        RECT 21.505 5.390 21.825 8.110 ;
        RECT 25.100 5.390 25.420 8.110 ;
        RECT 28.695 5.390 29.015 8.110 ;
        RECT 32.290 5.390 32.610 8.110 ;
        RECT 35.885 5.390 36.205 8.110 ;
        RECT 3.530 1.890 3.850 4.610 ;
        RECT 7.125 1.890 7.445 4.610 ;
        RECT 10.720 1.890 11.040 4.610 ;
        RECT 14.315 1.890 14.635 4.610 ;
        RECT 17.910 1.890 18.230 4.610 ;
        RECT 21.505 1.890 21.825 4.610 ;
        RECT 25.100 1.890 25.420 4.610 ;
        RECT 28.695 1.890 29.015 4.610 ;
        RECT 32.290 1.890 32.610 4.610 ;
        RECT 35.885 1.890 36.205 4.610 ;
        RECT 0.560 0.800 1.360 1.300 ;
  END
END sky130_asc_cap_mim_m3_1

#--------EOF---------

MACRO sky130_asc_pfet_01v8_lvt_9
  CLASS CORE ;
  FOREIGN sky130_asc_pfet_01v8_lvt_9 ;
  ORIGIN 0.000 0.000 ;
  SIZE 22.650 BY 9.400 ;
  SITE unitasc ;
  PIN GATE
    DIRECTION INOUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 116.099998 ;
    PORT
      LAYER li1 ;
        RECT 0.940 0.520 22.200 0.820 ;
    END
  END GATE
  PIN SOURCE
    DIRECTION INOUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 9.352500 ;
    PORT
      LAYER li1 ;
        RECT 1.240 8.450 22.200 8.650 ;
        RECT 3.465 8.245 3.635 8.450 ;
        RECT 8.045 8.245 8.215 8.450 ;
        RECT 12.625 8.245 12.795 8.450 ;
        RECT 17.205 8.245 17.375 8.450 ;
        RECT 21.785 8.245 21.955 8.450 ;
        RECT 3.465 8.130 3.640 8.245 ;
        RECT 8.045 8.130 8.220 8.245 ;
        RECT 12.625 8.130 12.800 8.245 ;
        RECT 17.205 8.130 17.380 8.245 ;
        RECT 21.785 8.130 21.960 8.245 ;
        RECT 3.470 1.755 3.640 8.130 ;
        RECT 8.050 1.755 8.220 8.130 ;
        RECT 12.630 1.755 12.800 8.130 ;
        RECT 17.210 1.755 17.380 8.130 ;
        RECT 21.790 1.755 21.960 8.130 ;
      LAYER mcon ;
        RECT 3.470 1.835 3.640 8.165 ;
        RECT 8.050 1.835 8.220 8.165 ;
        RECT 12.630 1.835 12.800 8.165 ;
        RECT 17.210 1.835 17.380 8.165 ;
        RECT 21.790 1.835 21.960 8.165 ;
      LAYER met1 ;
        RECT 3.440 1.775 3.670 8.225 ;
        RECT 8.020 1.775 8.250 8.225 ;
        RECT 12.600 1.775 12.830 8.225 ;
        RECT 17.180 1.775 17.410 8.225 ;
        RECT 21.760 1.775 21.990 8.225 ;
    END
  END SOURCE
  PIN DRAIN
    DIRECTION INOUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 9.352500 ;
    PORT
      LAYER li1 ;
        RECT 1.180 1.870 1.350 8.245 ;
        RECT 5.760 1.870 5.930 8.245 ;
        RECT 10.340 1.870 10.510 8.245 ;
        RECT 14.920 1.870 15.090 8.245 ;
        RECT 19.500 1.870 19.670 8.245 ;
        RECT 1.175 1.755 1.350 1.870 ;
        RECT 5.755 1.755 5.930 1.870 ;
        RECT 10.335 1.755 10.510 1.870 ;
        RECT 14.915 1.755 15.090 1.870 ;
        RECT 19.495 1.755 19.670 1.870 ;
        RECT 1.175 1.350 1.345 1.755 ;
        RECT 5.755 1.350 5.925 1.755 ;
        RECT 10.335 1.350 10.505 1.755 ;
        RECT 14.915 1.350 15.085 1.755 ;
        RECT 19.495 1.350 19.665 1.755 ;
        RECT 0.940 1.050 22.200 1.350 ;
      LAYER mcon ;
        RECT 1.180 1.835 1.350 8.165 ;
        RECT 5.760 1.835 5.930 8.165 ;
        RECT 10.340 1.835 10.510 8.165 ;
        RECT 14.920 1.835 15.090 8.165 ;
        RECT 19.500 1.835 19.670 8.165 ;
      LAYER met1 ;
        RECT 1.150 1.775 1.380 8.225 ;
        RECT 5.730 1.775 5.960 8.225 ;
        RECT 10.310 1.775 10.540 8.225 ;
        RECT 14.890 1.775 15.120 8.225 ;
        RECT 19.470 1.775 19.700 8.225 ;
    END
  END DRAIN
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT 0.450 1.470 22.200 9.700 ;
        RECT 0.940 1.465 22.200 1.470 ;
      LAYER li1 ;
        RECT 0.450 9.250 22.200 9.550 ;
        RECT 0.590 8.200 0.890 9.250 ;
        RECT 5.840 8.850 6.640 9.250 ;
        RECT 12.340 8.850 13.140 9.250 ;
      LAYER mcon ;
        RECT 1.790 9.250 2.090 9.550 ;
        RECT 3.790 9.250 4.090 9.550 ;
        RECT 5.790 9.250 6.090 9.550 ;
        RECT 7.790 9.250 8.090 9.550 ;
        RECT 9.790 9.250 10.090 9.550 ;
        RECT 11.790 9.250 12.090 9.550 ;
        RECT 13.790 9.250 14.090 9.550 ;
        RECT 15.790 9.250 16.090 9.550 ;
        RECT 17.790 9.250 18.090 9.550 ;
        RECT 19.790 9.250 20.090 9.550 ;
      LAYER met1 ;
        RECT 0.450 9.100 22.200 9.700 ;
    END
  END VPWR
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER li1 ;
        RECT 0.450 -0.150 22.200 0.150 ;
      LAYER mcon ;
        RECT 1.790 -0.150 2.090 0.150 ;
        RECT 3.790 -0.150 4.090 0.150 ;
        RECT 5.790 -0.150 6.090 0.150 ;
        RECT 7.790 -0.150 8.090 0.150 ;
        RECT 9.790 -0.150 10.090 0.150 ;
        RECT 11.790 -0.150 12.090 0.150 ;
        RECT 13.790 -0.150 14.090 0.150 ;
        RECT 15.790 -0.150 16.090 0.150 ;
        RECT 17.790 -0.150 18.090 0.150 ;
        RECT 19.790 -0.150 20.090 0.150 ;
      LAYER met1 ;
        RECT 0.450 -0.300 22.200 0.300 ;
    END
  END VGND
END sky130_asc_pfet_01v8_lvt_9

#--------EOF---------

END LIBRARY