VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO sky130_asc_pfet_01v8_lvt_6
  CLASS CORE ;
  FOREIGN sky130_asc_pfet_01v8_lvt_6 ;
  ORIGIN 0.000 0.000 ;
  SIZE 15.775 BY 9.400 ;
  SITE unitasc ;
  PIN GATE
    DIRECTION INOUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 77.400002 ;
    PORT
      LAYER li1 ;
        RECT 0.940 0.520 15.320 0.820 ;
    END
  END GATE
  PIN SOURCE
    DIRECTION INOUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 5.611500 ;
    PORT
      LAYER li1 ;
        RECT 1.240 8.450 15.320 8.650 ;
        RECT 3.465 1.755 3.635 8.450 ;
        RECT 8.045 1.755 8.215 8.450 ;
        RECT 12.625 1.755 12.795 8.450 ;
      LAYER mcon ;
        RECT 3.465 1.835 3.635 8.165 ;
        RECT 8.045 1.835 8.215 8.165 ;
        RECT 12.625 1.835 12.795 8.165 ;
      LAYER met1 ;
        RECT 3.435 1.775 3.665 8.225 ;
        RECT 8.015 1.775 8.245 8.225 ;
        RECT 12.595 1.775 12.825 8.225 ;
    END
  END SOURCE
  PIN DRAIN
    DIRECTION INOUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 7.482000 ;
    PORT
      LAYER li1 ;
        RECT 1.175 1.350 1.345 8.245 ;
        RECT 5.755 1.350 5.925 8.245 ;
        RECT 10.335 1.350 10.505 8.245 ;
        RECT 14.915 1.350 15.085 8.245 ;
        RECT 0.940 1.050 15.320 1.350 ;
      LAYER mcon ;
        RECT 1.175 1.835 1.345 8.165 ;
        RECT 5.755 1.835 5.925 8.165 ;
        RECT 10.335 1.835 10.505 8.165 ;
        RECT 14.915 1.835 15.085 8.165 ;
      LAYER met1 ;
        RECT 1.145 1.775 1.375 8.225 ;
        RECT 5.725 1.775 5.955 8.225 ;
        RECT 10.305 1.775 10.535 8.225 ;
        RECT 14.885 1.775 15.115 8.225 ;
    END
  END DRAIN
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT 0.450 8.535 15.320 9.700 ;
        RECT 0.450 1.470 15.325 8.535 ;
        RECT 0.935 1.465 15.325 1.470 ;
      LAYER li1 ;
        RECT 0.450 9.250 15.320 9.550 ;
        RECT 0.590 8.200 0.890 9.250 ;
        RECT 5.830 8.850 6.630 9.250 ;
      LAYER mcon ;
        RECT 1.790 9.250 2.090 9.550 ;
        RECT 3.790 9.250 4.090 9.550 ;
        RECT 5.790 9.250 6.090 9.550 ;
        RECT 7.790 9.250 8.090 9.550 ;
        RECT 9.790 9.250 10.090 9.550 ;
        RECT 11.790 9.250 12.090 9.550 ;
        RECT 13.790 9.250 14.090 9.550 ;
      LAYER met1 ;
        RECT 0.450 9.100 15.320 9.700 ;
    END
  END VPWR
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER li1 ;
        RECT 0.450 -0.150 15.320 0.150 ;
      LAYER mcon ;
        RECT 1.790 -0.150 2.090 0.150 ;
        RECT 3.790 -0.150 4.090 0.150 ;
        RECT 5.790 -0.150 6.090 0.150 ;
        RECT 7.790 -0.150 8.090 0.150 ;
        RECT 9.790 -0.150 10.090 0.150 ;
        RECT 11.790 -0.150 12.090 0.150 ;
        RECT 13.790 -0.150 14.090 0.150 ;
      LAYER met1 ;
        RECT 0.450 -0.300 15.320 0.300 ;
    END
  END VGND
END sky130_asc_pfet_01v8_lvt_6
END LIBRARY

