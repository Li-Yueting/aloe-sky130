magic
tech sky130A
magscale 1 2
timestamp 1654325418
<< nwell >>
rect 1257 863 2551 1513
<< pwell >>
rect 1267 409 2541 851
<< nmos >>
rect 1457 609 1487 713
rect 1553 609 1583 713
rect 1649 609 1679 713
rect 1745 609 1775 713
rect 1841 609 1871 713
rect 1937 609 1967 713
rect 2033 609 2063 713
rect 2129 609 2159 713
rect 2225 609 2255 713
rect 2321 609 2351 713
<< pmos >>
rect 1457 1021 1487 1293
rect 1553 1021 1583 1293
rect 1649 1021 1679 1293
rect 1745 1021 1775 1293
rect 1841 1021 1871 1293
rect 1937 1021 1967 1293
rect 2033 1021 2063 1293
rect 2129 1021 2159 1293
rect 2225 1021 2255 1293
rect 2321 1021 2351 1293
<< ndiff >>
rect 1395 678 1457 713
rect 1395 644 1407 678
rect 1441 644 1457 678
rect 1395 609 1457 644
rect 1487 678 1553 713
rect 1487 644 1503 678
rect 1537 644 1553 678
rect 1487 609 1553 644
rect 1583 678 1649 713
rect 1583 644 1599 678
rect 1633 644 1649 678
rect 1583 609 1649 644
rect 1679 678 1745 713
rect 1679 644 1695 678
rect 1729 644 1745 678
rect 1679 609 1745 644
rect 1775 678 1841 713
rect 1775 644 1791 678
rect 1825 644 1841 678
rect 1775 609 1841 644
rect 1871 678 1937 713
rect 1871 644 1887 678
rect 1921 644 1937 678
rect 1871 609 1937 644
rect 1967 678 2033 713
rect 1967 644 1983 678
rect 2017 644 2033 678
rect 1967 609 2033 644
rect 2063 678 2129 713
rect 2063 644 2079 678
rect 2113 644 2129 678
rect 2063 609 2129 644
rect 2159 678 2225 713
rect 2159 644 2175 678
rect 2209 644 2225 678
rect 2159 609 2225 644
rect 2255 678 2321 713
rect 2255 644 2271 678
rect 2305 644 2321 678
rect 2255 609 2321 644
rect 2351 678 2413 713
rect 2351 644 2367 678
rect 2401 644 2413 678
rect 2351 609 2413 644
<< pdiff >>
rect 1395 1276 1457 1293
rect 1395 1242 1407 1276
rect 1441 1242 1457 1276
rect 1395 1208 1457 1242
rect 1395 1174 1407 1208
rect 1441 1174 1457 1208
rect 1395 1140 1457 1174
rect 1395 1106 1407 1140
rect 1441 1106 1457 1140
rect 1395 1072 1457 1106
rect 1395 1038 1407 1072
rect 1441 1038 1457 1072
rect 1395 1021 1457 1038
rect 1487 1276 1553 1293
rect 1487 1242 1503 1276
rect 1537 1242 1553 1276
rect 1487 1208 1553 1242
rect 1487 1174 1503 1208
rect 1537 1174 1553 1208
rect 1487 1140 1553 1174
rect 1487 1106 1503 1140
rect 1537 1106 1553 1140
rect 1487 1072 1553 1106
rect 1487 1038 1503 1072
rect 1537 1038 1553 1072
rect 1487 1021 1553 1038
rect 1583 1276 1649 1293
rect 1583 1242 1599 1276
rect 1633 1242 1649 1276
rect 1583 1208 1649 1242
rect 1583 1174 1599 1208
rect 1633 1174 1649 1208
rect 1583 1140 1649 1174
rect 1583 1106 1599 1140
rect 1633 1106 1649 1140
rect 1583 1072 1649 1106
rect 1583 1038 1599 1072
rect 1633 1038 1649 1072
rect 1583 1021 1649 1038
rect 1679 1276 1745 1293
rect 1679 1242 1695 1276
rect 1729 1242 1745 1276
rect 1679 1208 1745 1242
rect 1679 1174 1695 1208
rect 1729 1174 1745 1208
rect 1679 1140 1745 1174
rect 1679 1106 1695 1140
rect 1729 1106 1745 1140
rect 1679 1072 1745 1106
rect 1679 1038 1695 1072
rect 1729 1038 1745 1072
rect 1679 1021 1745 1038
rect 1775 1276 1841 1293
rect 1775 1242 1791 1276
rect 1825 1242 1841 1276
rect 1775 1208 1841 1242
rect 1775 1174 1791 1208
rect 1825 1174 1841 1208
rect 1775 1140 1841 1174
rect 1775 1106 1791 1140
rect 1825 1106 1841 1140
rect 1775 1072 1841 1106
rect 1775 1038 1791 1072
rect 1825 1038 1841 1072
rect 1775 1021 1841 1038
rect 1871 1276 1937 1293
rect 1871 1242 1887 1276
rect 1921 1242 1937 1276
rect 1871 1208 1937 1242
rect 1871 1174 1887 1208
rect 1921 1174 1937 1208
rect 1871 1140 1937 1174
rect 1871 1106 1887 1140
rect 1921 1106 1937 1140
rect 1871 1072 1937 1106
rect 1871 1038 1887 1072
rect 1921 1038 1937 1072
rect 1871 1021 1937 1038
rect 1967 1276 2033 1293
rect 1967 1242 1983 1276
rect 2017 1242 2033 1276
rect 1967 1208 2033 1242
rect 1967 1174 1983 1208
rect 2017 1174 2033 1208
rect 1967 1140 2033 1174
rect 1967 1106 1983 1140
rect 2017 1106 2033 1140
rect 1967 1072 2033 1106
rect 1967 1038 1983 1072
rect 2017 1038 2033 1072
rect 1967 1021 2033 1038
rect 2063 1276 2129 1293
rect 2063 1242 2079 1276
rect 2113 1242 2129 1276
rect 2063 1208 2129 1242
rect 2063 1174 2079 1208
rect 2113 1174 2129 1208
rect 2063 1140 2129 1174
rect 2063 1106 2079 1140
rect 2113 1106 2129 1140
rect 2063 1072 2129 1106
rect 2063 1038 2079 1072
rect 2113 1038 2129 1072
rect 2063 1021 2129 1038
rect 2159 1276 2225 1293
rect 2159 1242 2175 1276
rect 2209 1242 2225 1276
rect 2159 1208 2225 1242
rect 2159 1174 2175 1208
rect 2209 1174 2225 1208
rect 2159 1140 2225 1174
rect 2159 1106 2175 1140
rect 2209 1106 2225 1140
rect 2159 1072 2225 1106
rect 2159 1038 2175 1072
rect 2209 1038 2225 1072
rect 2159 1021 2225 1038
rect 2255 1276 2321 1293
rect 2255 1242 2271 1276
rect 2305 1242 2321 1276
rect 2255 1208 2321 1242
rect 2255 1174 2271 1208
rect 2305 1174 2321 1208
rect 2255 1140 2321 1174
rect 2255 1106 2271 1140
rect 2305 1106 2321 1140
rect 2255 1072 2321 1106
rect 2255 1038 2271 1072
rect 2305 1038 2321 1072
rect 2255 1021 2321 1038
rect 2351 1276 2413 1293
rect 2351 1242 2367 1276
rect 2401 1242 2413 1276
rect 2351 1208 2413 1242
rect 2351 1174 2367 1208
rect 2401 1174 2413 1208
rect 2351 1140 2413 1174
rect 2351 1106 2367 1140
rect 2401 1106 2413 1140
rect 2351 1072 2413 1106
rect 2351 1038 2367 1072
rect 2401 1038 2413 1072
rect 2351 1021 2413 1038
<< ndiffc >>
rect 1407 644 1441 678
rect 1503 644 1537 678
rect 1599 644 1633 678
rect 1695 644 1729 678
rect 1791 644 1825 678
rect 1887 644 1921 678
rect 1983 644 2017 678
rect 2079 644 2113 678
rect 2175 644 2209 678
rect 2271 644 2305 678
rect 2367 644 2401 678
<< pdiffc >>
rect 1407 1242 1441 1276
rect 1407 1174 1441 1208
rect 1407 1106 1441 1140
rect 1407 1038 1441 1072
rect 1503 1242 1537 1276
rect 1503 1174 1537 1208
rect 1503 1106 1537 1140
rect 1503 1038 1537 1072
rect 1599 1242 1633 1276
rect 1599 1174 1633 1208
rect 1599 1106 1633 1140
rect 1599 1038 1633 1072
rect 1695 1242 1729 1276
rect 1695 1174 1729 1208
rect 1695 1106 1729 1140
rect 1695 1038 1729 1072
rect 1791 1242 1825 1276
rect 1791 1174 1825 1208
rect 1791 1106 1825 1140
rect 1791 1038 1825 1072
rect 1887 1242 1921 1276
rect 1887 1174 1921 1208
rect 1887 1106 1921 1140
rect 1887 1038 1921 1072
rect 1983 1242 2017 1276
rect 1983 1174 2017 1208
rect 1983 1106 2017 1140
rect 1983 1038 2017 1072
rect 2079 1242 2113 1276
rect 2079 1174 2113 1208
rect 2079 1106 2113 1140
rect 2079 1038 2113 1072
rect 2175 1242 2209 1276
rect 2175 1174 2209 1208
rect 2175 1106 2209 1140
rect 2175 1038 2209 1072
rect 2271 1242 2305 1276
rect 2271 1174 2305 1208
rect 2271 1106 2305 1140
rect 2271 1038 2305 1072
rect 2367 1242 2401 1276
rect 2367 1174 2401 1208
rect 2367 1106 2401 1140
rect 2367 1038 2401 1072
<< psubdiff >>
rect 1293 791 1411 825
rect 1445 791 1479 825
rect 1513 791 1547 825
rect 1581 791 1615 825
rect 1649 791 1683 825
rect 1717 791 1751 825
rect 1785 791 1819 825
rect 1853 791 1887 825
rect 1921 791 1955 825
rect 1989 791 2023 825
rect 2057 791 2091 825
rect 2125 791 2159 825
rect 2193 791 2227 825
rect 2261 791 2295 825
rect 2329 791 2363 825
rect 2397 791 2515 825
rect 1293 715 1327 791
rect 2481 715 2515 791
rect 1293 647 1327 681
rect 1293 579 1327 613
rect 2481 647 2515 681
rect 1293 469 1327 545
rect 2481 579 2515 613
rect 2481 469 2515 545
rect 1293 435 1411 469
rect 1445 435 1479 469
rect 1513 435 1547 469
rect 1581 435 1615 469
rect 1649 435 1683 469
rect 1717 435 1751 469
rect 1785 435 1819 469
rect 1853 435 1887 469
rect 1921 435 1955 469
rect 1989 435 2023 469
rect 2057 435 2091 469
rect 2125 435 2159 469
rect 2193 435 2227 469
rect 2261 435 2295 469
rect 2329 435 2363 469
rect 2397 435 2515 469
<< nsubdiff >>
rect 1293 1443 1411 1477
rect 1445 1443 1479 1477
rect 1513 1443 1547 1477
rect 1581 1443 1615 1477
rect 1649 1443 1683 1477
rect 1717 1443 1751 1477
rect 1785 1443 1819 1477
rect 1853 1443 1887 1477
rect 1921 1443 1955 1477
rect 1989 1443 2023 1477
rect 2057 1443 2091 1477
rect 2125 1443 2159 1477
rect 2193 1443 2227 1477
rect 2261 1443 2295 1477
rect 2329 1443 2363 1477
rect 2397 1443 2515 1477
rect 1293 1375 1327 1443
rect 1293 1307 1327 1341
rect 2481 1375 2515 1443
rect 2481 1307 2515 1341
rect 1293 1239 1327 1273
rect 1293 1171 1327 1205
rect 1293 1103 1327 1137
rect 1293 1035 1327 1069
rect 2481 1239 2515 1273
rect 2481 1171 2515 1205
rect 2481 1103 2515 1137
rect 2481 1035 2515 1069
rect 1293 933 1327 1001
rect 2481 933 2515 1001
rect 1293 899 1411 933
rect 1445 899 1479 933
rect 1513 899 1547 933
rect 1581 899 1615 933
rect 1649 899 1683 933
rect 1717 899 1751 933
rect 1785 899 1819 933
rect 1853 899 1887 933
rect 1921 899 1955 933
rect 1989 899 2023 933
rect 2057 899 2091 933
rect 2125 899 2159 933
rect 2193 899 2227 933
rect 2261 899 2295 933
rect 2329 899 2363 933
rect 2397 899 2515 933
<< psubdiffcont >>
rect 1411 791 1445 825
rect 1479 791 1513 825
rect 1547 791 1581 825
rect 1615 791 1649 825
rect 1683 791 1717 825
rect 1751 791 1785 825
rect 1819 791 1853 825
rect 1887 791 1921 825
rect 1955 791 1989 825
rect 2023 791 2057 825
rect 2091 791 2125 825
rect 2159 791 2193 825
rect 2227 791 2261 825
rect 2295 791 2329 825
rect 2363 791 2397 825
rect 1293 681 1327 715
rect 1293 613 1327 647
rect 2481 681 2515 715
rect 2481 613 2515 647
rect 1293 545 1327 579
rect 2481 545 2515 579
rect 1411 435 1445 469
rect 1479 435 1513 469
rect 1547 435 1581 469
rect 1615 435 1649 469
rect 1683 435 1717 469
rect 1751 435 1785 469
rect 1819 435 1853 469
rect 1887 435 1921 469
rect 1955 435 1989 469
rect 2023 435 2057 469
rect 2091 435 2125 469
rect 2159 435 2193 469
rect 2227 435 2261 469
rect 2295 435 2329 469
rect 2363 435 2397 469
<< nsubdiffcont >>
rect 1411 1443 1445 1477
rect 1479 1443 1513 1477
rect 1547 1443 1581 1477
rect 1615 1443 1649 1477
rect 1683 1443 1717 1477
rect 1751 1443 1785 1477
rect 1819 1443 1853 1477
rect 1887 1443 1921 1477
rect 1955 1443 1989 1477
rect 2023 1443 2057 1477
rect 2091 1443 2125 1477
rect 2159 1443 2193 1477
rect 2227 1443 2261 1477
rect 2295 1443 2329 1477
rect 2363 1443 2397 1477
rect 1293 1341 1327 1375
rect 2481 1341 2515 1375
rect 1293 1273 1327 1307
rect 1293 1205 1327 1239
rect 1293 1137 1327 1171
rect 1293 1069 1327 1103
rect 1293 1001 1327 1035
rect 2481 1273 2515 1307
rect 2481 1205 2515 1239
rect 2481 1137 2515 1171
rect 2481 1069 2515 1103
rect 2481 1001 2515 1035
rect 1411 899 1445 933
rect 1479 899 1513 933
rect 1547 899 1581 933
rect 1615 899 1649 933
rect 1683 899 1717 933
rect 1751 899 1785 933
rect 1819 899 1853 933
rect 1887 899 1921 933
rect 1955 899 1989 933
rect 2023 899 2057 933
rect 2091 899 2125 933
rect 2159 899 2193 933
rect 2227 899 2261 933
rect 2295 899 2329 933
rect 2363 899 2397 933
<< poly >>
rect 1391 1375 2417 1391
rect 1391 1341 1407 1375
rect 1441 1341 1599 1375
rect 1633 1341 1791 1375
rect 1825 1341 1983 1375
rect 2017 1341 2175 1375
rect 2209 1341 2367 1375
rect 2401 1341 2417 1375
rect 1391 1325 2417 1341
rect 1457 1293 1487 1325
rect 1553 1293 1583 1325
rect 1649 1293 1679 1325
rect 1745 1293 1775 1325
rect 1841 1293 1871 1325
rect 1937 1293 1967 1325
rect 2033 1293 2063 1325
rect 2129 1293 2159 1325
rect 2225 1293 2255 1325
rect 2321 1293 2351 1325
rect 1457 995 1487 1021
rect 1553 995 1583 1021
rect 1649 995 1679 1021
rect 1745 995 1775 1021
rect 1841 995 1871 1021
rect 1937 995 1967 1021
rect 2033 995 2063 1021
rect 2129 995 2159 1021
rect 2225 995 2255 1021
rect 2321 995 2351 1021
rect 1457 713 1487 739
rect 1553 713 1583 739
rect 1649 713 1679 739
rect 1745 713 1775 739
rect 1841 713 1871 739
rect 1937 713 1967 739
rect 2033 713 2063 739
rect 2129 713 2159 739
rect 2225 713 2255 739
rect 2321 713 2351 739
rect 1457 587 1487 609
rect 1553 587 1583 609
rect 1649 587 1679 609
rect 1745 587 1775 609
rect 1841 587 1871 609
rect 1937 587 1967 609
rect 2033 587 2063 609
rect 2129 587 2159 609
rect 2225 587 2255 609
rect 2321 587 2351 609
rect 1391 567 2417 587
rect 1391 533 1407 567
rect 1441 533 1599 567
rect 1633 533 1791 567
rect 1825 533 1983 567
rect 2017 533 2175 567
rect 2209 533 2367 567
rect 2401 533 2417 567
rect 1391 521 2417 533
<< polycont >>
rect 1407 1341 1441 1375
rect 1599 1341 1633 1375
rect 1791 1341 1825 1375
rect 1983 1341 2017 1375
rect 2175 1341 2209 1375
rect 2367 1341 2401 1375
rect 1407 533 1441 567
rect 1599 533 1633 567
rect 1791 533 1825 567
rect 1983 533 2017 567
rect 2175 533 2209 567
rect 2367 533 2401 567
<< locali >>
rect 1293 1443 1411 1477
rect 1445 1443 1479 1477
rect 1513 1443 1547 1477
rect 1581 1443 1615 1477
rect 1649 1443 1683 1477
rect 1717 1443 1751 1477
rect 1785 1443 1819 1477
rect 1853 1443 1887 1477
rect 1921 1443 1955 1477
rect 1989 1443 2023 1477
rect 2057 1443 2091 1477
rect 2125 1443 2159 1477
rect 2193 1443 2227 1477
rect 2261 1443 2295 1477
rect 2329 1443 2363 1477
rect 2397 1443 2515 1477
rect 1293 1375 1327 1443
rect 2481 1375 2515 1443
rect 1391 1341 1407 1375
rect 1441 1341 1457 1375
rect 1583 1341 1599 1375
rect 1633 1341 1649 1375
rect 1775 1341 1791 1375
rect 1825 1341 1841 1375
rect 1967 1341 1983 1375
rect 2017 1341 2033 1375
rect 2159 1341 2175 1375
rect 2209 1341 2225 1375
rect 2351 1341 2367 1375
rect 2401 1341 2417 1375
rect 1293 1307 1327 1341
rect 2481 1307 2515 1315
rect 1293 1239 1327 1273
rect 1293 1171 1327 1205
rect 1293 1103 1327 1137
rect 1293 1035 1327 1069
rect 1407 1276 1441 1297
rect 1407 1208 1441 1212
rect 1407 1102 1441 1106
rect 1407 1017 1441 1038
rect 1503 1276 1537 1297
rect 1503 1208 1537 1212
rect 1503 1102 1537 1106
rect 1503 1017 1537 1038
rect 1599 1276 1633 1297
rect 1599 1208 1633 1212
rect 1599 1102 1633 1106
rect 1599 1017 1633 1038
rect 1695 1276 1729 1297
rect 1695 1208 1729 1212
rect 1695 1102 1729 1106
rect 1695 1017 1729 1038
rect 1791 1276 1825 1297
rect 1791 1208 1825 1212
rect 1791 1102 1825 1106
rect 1791 1017 1825 1038
rect 1887 1276 1921 1297
rect 1887 1208 1921 1212
rect 1887 1102 1921 1106
rect 1887 1017 1921 1038
rect 1983 1276 2017 1297
rect 1983 1208 2017 1212
rect 1983 1102 2017 1106
rect 1983 1017 2017 1038
rect 2079 1276 2113 1297
rect 2079 1208 2113 1212
rect 2079 1102 2113 1106
rect 2079 1017 2113 1038
rect 2175 1276 2209 1297
rect 2175 1208 2209 1212
rect 2175 1102 2209 1106
rect 2175 1017 2209 1038
rect 2271 1276 2305 1297
rect 2271 1208 2305 1212
rect 2271 1102 2305 1106
rect 2271 1017 2305 1038
rect 2367 1276 2401 1297
rect 2367 1208 2401 1212
rect 2367 1102 2401 1106
rect 2367 1017 2401 1038
rect 2481 1239 2515 1243
rect 2481 1133 2515 1137
rect 2481 1061 2515 1069
rect 1293 933 1327 1001
rect 2481 933 2515 1001
rect 1293 899 1411 933
rect 1445 899 1479 933
rect 1513 899 1547 933
rect 1581 899 1615 933
rect 1649 899 1683 933
rect 1717 899 1751 933
rect 1785 899 1819 933
rect 1853 899 1887 933
rect 1921 899 1955 933
rect 1989 899 2023 933
rect 2057 899 2091 933
rect 2125 899 2159 933
rect 2193 899 2227 933
rect 2261 899 2295 933
rect 2329 899 2363 933
rect 2397 899 2515 933
rect 1293 791 1411 825
rect 1445 791 1479 825
rect 1513 791 1547 825
rect 1581 791 1615 825
rect 1649 791 1683 825
rect 1717 791 1751 825
rect 1785 791 1819 825
rect 1853 791 1887 825
rect 1921 791 1955 825
rect 1989 791 2023 825
rect 2057 791 2091 825
rect 2125 791 2159 825
rect 2193 791 2227 825
rect 2261 791 2295 825
rect 2329 791 2363 825
rect 2397 791 2515 825
rect 1293 715 1327 791
rect 2481 720 2515 791
rect 1293 647 1327 681
rect 1293 579 1327 613
rect 1407 678 1441 717
rect 1407 605 1441 644
rect 1503 678 1537 717
rect 1503 605 1537 644
rect 1599 678 1633 717
rect 1599 605 1633 644
rect 1695 678 1729 717
rect 1695 605 1729 644
rect 1791 678 1825 717
rect 1791 605 1825 644
rect 1887 678 1921 717
rect 1887 605 1921 644
rect 1983 678 2017 717
rect 1983 605 2017 644
rect 2079 678 2113 717
rect 2079 605 2113 644
rect 2175 678 2209 717
rect 2175 605 2209 644
rect 2271 678 2305 717
rect 2271 605 2305 644
rect 2367 678 2401 717
rect 2367 605 2401 644
rect 2481 648 2515 681
rect 2481 579 2515 613
rect 1293 469 1327 545
rect 1391 533 1407 567
rect 1441 533 1457 567
rect 1583 533 1599 567
rect 1633 533 1649 567
rect 1775 533 1791 567
rect 1825 533 1841 567
rect 1967 533 1983 567
rect 2017 533 2033 567
rect 2159 533 2175 567
rect 2209 533 2225 567
rect 2351 533 2367 567
rect 2401 533 2417 567
rect 2481 469 2515 542
rect 1293 435 1411 469
rect 1445 435 1479 469
rect 1513 435 1547 469
rect 1581 435 1615 469
rect 1649 435 1683 469
rect 1717 435 1751 469
rect 1785 435 1819 469
rect 1853 435 1887 469
rect 1921 435 1955 469
rect 1989 435 2023 469
rect 2057 435 2091 469
rect 2125 435 2159 469
rect 2193 435 2227 469
rect 2261 435 2295 469
rect 2329 435 2363 469
rect 2397 435 2515 469
<< viali >>
rect 1407 1341 1441 1375
rect 1599 1341 1633 1375
rect 1791 1341 1825 1375
rect 1983 1341 2017 1375
rect 2175 1341 2209 1375
rect 2367 1341 2401 1375
rect 2481 1341 2515 1349
rect 2481 1315 2515 1341
rect 1407 1242 1441 1246
rect 1407 1212 1441 1242
rect 1407 1140 1441 1174
rect 1407 1072 1441 1102
rect 1407 1068 1441 1072
rect 1503 1242 1537 1246
rect 1503 1212 1537 1242
rect 1503 1140 1537 1174
rect 1503 1072 1537 1102
rect 1503 1068 1537 1072
rect 1599 1242 1633 1246
rect 1599 1212 1633 1242
rect 1599 1140 1633 1174
rect 1599 1072 1633 1102
rect 1599 1068 1633 1072
rect 1695 1242 1729 1246
rect 1695 1212 1729 1242
rect 1695 1140 1729 1174
rect 1695 1072 1729 1102
rect 1695 1068 1729 1072
rect 1791 1242 1825 1246
rect 1791 1212 1825 1242
rect 1791 1140 1825 1174
rect 1791 1072 1825 1102
rect 1791 1068 1825 1072
rect 1887 1242 1921 1246
rect 1887 1212 1921 1242
rect 1887 1140 1921 1174
rect 1887 1072 1921 1102
rect 1887 1068 1921 1072
rect 1983 1242 2017 1246
rect 1983 1212 2017 1242
rect 1983 1140 2017 1174
rect 1983 1072 2017 1102
rect 1983 1068 2017 1072
rect 2079 1242 2113 1246
rect 2079 1212 2113 1242
rect 2079 1140 2113 1174
rect 2079 1072 2113 1102
rect 2079 1068 2113 1072
rect 2175 1242 2209 1246
rect 2175 1212 2209 1242
rect 2175 1140 2209 1174
rect 2175 1072 2209 1102
rect 2175 1068 2209 1072
rect 2271 1242 2305 1246
rect 2271 1212 2305 1242
rect 2271 1140 2305 1174
rect 2271 1072 2305 1102
rect 2271 1068 2305 1072
rect 2367 1242 2401 1246
rect 2367 1212 2401 1242
rect 2367 1140 2401 1174
rect 2367 1072 2401 1102
rect 2367 1068 2401 1072
rect 2481 1273 2515 1277
rect 2481 1243 2515 1273
rect 2481 1171 2515 1205
rect 2481 1103 2515 1133
rect 2481 1099 2515 1103
rect 2481 1035 2515 1061
rect 2481 1027 2515 1035
rect 1407 644 1441 678
rect 1503 644 1537 678
rect 1599 644 1633 678
rect 1695 644 1729 678
rect 1791 644 1825 678
rect 1887 644 1921 678
rect 1983 644 2017 678
rect 2079 644 2113 678
rect 2175 644 2209 678
rect 2271 644 2305 678
rect 2367 644 2401 678
rect 2481 715 2515 720
rect 2481 686 2515 715
rect 2481 647 2515 648
rect 2481 614 2515 647
rect 1407 533 1441 567
rect 1599 533 1633 567
rect 1791 533 1825 567
rect 1983 533 2017 567
rect 2175 533 2209 567
rect 2367 533 2401 567
rect 2481 545 2515 576
rect 2481 542 2515 545
<< metal1 >>
rect 1223 1443 2305 1477
rect 1223 880 1257 1443
rect 1388 1333 1398 1385
rect 1450 1333 1460 1385
rect 1503 1293 1537 1443
rect 1581 1333 1591 1385
rect 1643 1333 1653 1385
rect 1695 1293 1729 1443
rect 1772 1333 1782 1385
rect 1834 1333 1844 1385
rect 1887 1293 1921 1443
rect 1964 1333 1974 1385
rect 2026 1333 2036 1385
rect 2079 1293 2113 1443
rect 2156 1333 2166 1385
rect 2218 1333 2228 1385
rect 2271 1293 2305 1443
rect 2348 1333 2358 1385
rect 2410 1333 2420 1385
rect 2475 1349 2521 1513
rect 2475 1315 2481 1349
rect 2515 1315 2521 1349
rect 2606 1326 2616 1386
rect 2672 1326 2886 1386
rect 2946 1326 2956 1386
rect 1401 1246 1447 1293
rect 1401 1212 1407 1246
rect 1441 1212 1447 1246
rect 1401 1174 1447 1212
rect 1401 1140 1407 1174
rect 1441 1140 1447 1174
rect 1401 1102 1447 1140
rect 1401 1068 1407 1102
rect 1441 1068 1447 1102
rect 1401 1021 1447 1068
rect 1497 1246 1543 1293
rect 1497 1212 1503 1246
rect 1537 1212 1543 1246
rect 1497 1174 1543 1212
rect 1497 1140 1503 1174
rect 1537 1140 1543 1174
rect 1497 1102 1543 1140
rect 1497 1068 1503 1102
rect 1537 1068 1543 1102
rect 1497 1021 1543 1068
rect 1593 1246 1639 1293
rect 1593 1212 1599 1246
rect 1633 1212 1639 1246
rect 1593 1174 1639 1212
rect 1593 1140 1599 1174
rect 1633 1140 1639 1174
rect 1593 1102 1639 1140
rect 1593 1068 1599 1102
rect 1633 1068 1639 1102
rect 1593 1021 1639 1068
rect 1689 1246 1735 1293
rect 1689 1212 1695 1246
rect 1729 1212 1735 1246
rect 1689 1174 1735 1212
rect 1689 1140 1695 1174
rect 1729 1140 1735 1174
rect 1689 1102 1735 1140
rect 1689 1068 1695 1102
rect 1729 1068 1735 1102
rect 1689 1021 1735 1068
rect 1785 1246 1831 1293
rect 1785 1212 1791 1246
rect 1825 1212 1831 1246
rect 1785 1174 1831 1212
rect 1785 1140 1791 1174
rect 1825 1140 1831 1174
rect 1785 1102 1831 1140
rect 1785 1068 1791 1102
rect 1825 1068 1831 1102
rect 1785 1021 1831 1068
rect 1881 1246 1927 1293
rect 1881 1212 1887 1246
rect 1921 1212 1927 1246
rect 1881 1174 1927 1212
rect 1881 1140 1887 1174
rect 1921 1140 1927 1174
rect 1881 1102 1927 1140
rect 1881 1068 1887 1102
rect 1921 1068 1927 1102
rect 1881 1021 1927 1068
rect 1977 1246 2023 1293
rect 1977 1212 1983 1246
rect 2017 1212 2023 1246
rect 1977 1174 2023 1212
rect 1977 1140 1983 1174
rect 2017 1140 2023 1174
rect 1977 1102 2023 1140
rect 1977 1068 1983 1102
rect 2017 1068 2023 1102
rect 1977 1021 2023 1068
rect 2073 1246 2119 1293
rect 2073 1212 2079 1246
rect 2113 1212 2119 1246
rect 2073 1174 2119 1212
rect 2073 1140 2079 1174
rect 2113 1140 2119 1174
rect 2073 1102 2119 1140
rect 2073 1068 2079 1102
rect 2113 1068 2119 1102
rect 2073 1021 2119 1068
rect 2169 1246 2215 1293
rect 2169 1212 2175 1246
rect 2209 1212 2215 1246
rect 2169 1174 2215 1212
rect 2169 1140 2175 1174
rect 2209 1140 2215 1174
rect 2169 1102 2215 1140
rect 2169 1068 2175 1102
rect 2209 1068 2215 1102
rect 2169 1021 2215 1068
rect 2265 1246 2311 1293
rect 2265 1212 2271 1246
rect 2305 1212 2311 1246
rect 2265 1174 2311 1212
rect 2265 1140 2271 1174
rect 2305 1140 2311 1174
rect 2265 1102 2311 1140
rect 2265 1068 2271 1102
rect 2305 1068 2311 1102
rect 2265 1021 2311 1068
rect 2361 1246 2407 1293
rect 2361 1212 2367 1246
rect 2401 1212 2407 1246
rect 2361 1174 2407 1212
rect 2361 1140 2367 1174
rect 2401 1140 2407 1174
rect 2361 1102 2407 1140
rect 2361 1068 2367 1102
rect 2401 1068 2407 1102
rect 2361 1021 2407 1068
rect 2475 1277 2521 1315
rect 2475 1243 2481 1277
rect 2515 1243 2521 1277
rect 2475 1205 2521 1243
rect 2475 1171 2481 1205
rect 2515 1171 2521 1205
rect 2475 1133 2521 1171
rect 2475 1099 2481 1133
rect 2515 1099 2521 1133
rect 2475 1061 2521 1099
rect 2475 1027 2481 1061
rect 2515 1027 2521 1061
rect 1094 846 1257 880
rect 1223 469 1257 846
rect 1407 880 1441 1021
rect 1599 880 1633 1021
rect 1791 880 1825 1021
rect 1983 880 2017 1021
rect 2175 880 2209 1021
rect 2367 880 2401 1021
rect 2475 983 2521 1027
rect 1407 846 2593 880
rect 1407 713 1441 846
rect 1599 713 1633 846
rect 1791 713 1825 846
rect 1983 713 2017 846
rect 2175 713 2209 846
rect 2367 713 2401 846
rect 2475 720 2521 743
rect 1401 678 1447 713
rect 1401 644 1407 678
rect 1441 644 1447 678
rect 1401 609 1447 644
rect 1497 678 1543 713
rect 1497 644 1503 678
rect 1537 644 1543 678
rect 1497 609 1543 644
rect 1593 678 1639 713
rect 1593 644 1599 678
rect 1633 644 1639 678
rect 1593 609 1639 644
rect 1689 678 1735 713
rect 1689 644 1695 678
rect 1729 644 1735 678
rect 1689 609 1735 644
rect 1785 678 1831 713
rect 1785 644 1791 678
rect 1825 644 1831 678
rect 1785 609 1831 644
rect 1881 678 1927 713
rect 1881 644 1887 678
rect 1921 644 1927 678
rect 1881 609 1927 644
rect 1977 678 2023 713
rect 1977 644 1983 678
rect 2017 644 2023 678
rect 1977 609 2023 644
rect 2073 678 2119 713
rect 2073 644 2079 678
rect 2113 644 2119 678
rect 2073 609 2119 644
rect 2169 678 2215 713
rect 2169 644 2175 678
rect 2209 644 2215 678
rect 2169 609 2215 644
rect 2265 678 2311 713
rect 2265 644 2271 678
rect 2305 644 2311 678
rect 2265 609 2311 644
rect 2361 678 2407 713
rect 2361 644 2367 678
rect 2401 644 2407 678
rect 2361 609 2407 644
rect 2475 686 2481 720
rect 2515 686 2521 720
rect 2475 648 2521 686
rect 2475 614 2481 648
rect 2515 614 2521 648
rect 1391 578 1457 581
rect 1388 526 1398 578
rect 1450 526 1460 578
rect 1391 521 1457 526
rect 1503 469 1537 609
rect 1583 578 1649 581
rect 1579 526 1589 578
rect 1641 526 1651 578
rect 1583 521 1649 526
rect 1695 469 1729 609
rect 1775 578 1841 581
rect 1771 526 1781 578
rect 1833 526 1843 578
rect 1775 521 1841 526
rect 1887 469 1921 609
rect 1967 578 2033 581
rect 1963 526 1973 578
rect 2025 526 2035 578
rect 1967 521 2033 526
rect 2079 469 2113 609
rect 2159 577 2225 581
rect 2156 525 2166 577
rect 2218 525 2228 577
rect 2159 521 2225 525
rect 2271 469 2305 609
rect 2351 577 2417 581
rect 2348 525 2358 577
rect 2410 525 2420 577
rect 2475 576 2521 614
rect 2475 542 2481 576
rect 2515 542 2521 576
rect 2351 521 2417 525
rect 1223 435 2305 469
rect 2475 399 2521 542
<< via1 >>
rect 1398 1375 1450 1385
rect 1398 1341 1407 1375
rect 1407 1341 1441 1375
rect 1441 1341 1450 1375
rect 1398 1333 1450 1341
rect 1591 1375 1643 1385
rect 1591 1341 1599 1375
rect 1599 1341 1633 1375
rect 1633 1341 1643 1375
rect 1591 1333 1643 1341
rect 1782 1375 1834 1385
rect 1782 1341 1791 1375
rect 1791 1341 1825 1375
rect 1825 1341 1834 1375
rect 1782 1333 1834 1341
rect 1974 1375 2026 1385
rect 1974 1341 1983 1375
rect 1983 1341 2017 1375
rect 2017 1341 2026 1375
rect 1974 1333 2026 1341
rect 2166 1375 2218 1385
rect 2166 1341 2175 1375
rect 2175 1341 2209 1375
rect 2209 1341 2218 1375
rect 2166 1333 2218 1341
rect 2358 1375 2410 1385
rect 2358 1341 2367 1375
rect 2367 1341 2401 1375
rect 2401 1341 2410 1375
rect 2358 1333 2410 1341
rect 2616 1326 2672 1386
rect 2886 1326 2946 1386
rect 1398 567 1450 578
rect 1398 533 1407 567
rect 1407 533 1441 567
rect 1441 533 1450 567
rect 1398 526 1450 533
rect 1589 567 1641 578
rect 1589 533 1599 567
rect 1599 533 1633 567
rect 1633 533 1641 567
rect 1589 526 1641 533
rect 1781 567 1833 578
rect 1781 533 1791 567
rect 1791 533 1825 567
rect 1825 533 1833 567
rect 1781 526 1833 533
rect 1973 567 2025 578
rect 1973 533 1983 567
rect 1983 533 2017 567
rect 2017 533 2025 567
rect 1973 526 2025 533
rect 2166 567 2218 577
rect 2166 533 2175 567
rect 2175 533 2209 567
rect 2209 533 2218 567
rect 2166 525 2218 533
rect 2358 567 2410 577
rect 2358 533 2367 567
rect 2367 533 2401 567
rect 2401 533 2410 567
rect 2358 525 2410 533
<< metal2 >>
rect 1398 1385 1450 1395
rect 1591 1385 1643 1395
rect 1782 1385 1834 1395
rect 1974 1385 2026 1395
rect 2166 1385 2218 1395
rect 2358 1385 2410 1395
rect 2616 1386 2672 1396
rect 1120 1333 1398 1385
rect 1450 1333 1591 1385
rect 1643 1333 1782 1385
rect 1834 1333 1974 1385
rect 2026 1333 2166 1385
rect 2218 1333 2358 1385
rect 2410 1333 2616 1385
rect 1398 1323 1450 1333
rect 1591 1323 1643 1333
rect 1782 1323 1834 1333
rect 1974 1323 2026 1333
rect 2166 1323 2218 1333
rect 2358 1323 2410 1333
rect 2616 1316 2672 1326
rect 2886 1386 2946 1396
rect 2886 1190 2946 1326
rect 1398 578 1450 588
rect 1589 578 1641 588
rect 1781 578 1833 588
rect 1973 578 2025 588
rect 2166 578 2218 587
rect 2358 578 2410 587
rect 1121 526 1398 578
rect 1450 526 1589 578
rect 1641 526 1781 578
rect 1833 526 1973 578
rect 2025 577 2596 578
rect 2025 526 2166 577
rect 1398 516 1450 526
rect 1589 516 1641 526
rect 1781 516 1833 526
rect 1973 516 2025 526
rect 2218 526 2358 577
rect 2166 515 2218 525
rect 2410 526 2596 577
rect 2358 515 2410 525
<< labels >>
flabel metal2 1120 1333 1172 1385 1 FreeSans 480 0 0 0 en_b
flabel metal2 1122 526 1182 578 1 FreeSans 480 0 0 0 en
flabel metal1 s 2498 402 2498 402 1 FreeSans 500 0 0 0 VSS
port 6 nsew
flabel metal1 s 2498 1508 2498 1508 5 FreeSans 500 0 0 0 VDD
port 5 nsew
flabel metal1 s 2589 862 2589 862 7 FreeSans 500 0 0 0 out
port 4 nsew
flabel metal1 s 1098 863 1098 863 3 FreeSans 500 0 0 0 in
port 2 nsew
<< end >>
