magic
tech sky130A
magscale 1 2
timestamp 1654744774
<< nwell >>
rect 24732 48779 52438 49012
rect 24732 47366 52439 48779
rect 24829 47365 52439 47366
rect 14932 45019 42638 45252
rect 14932 43606 42639 45019
rect 15029 43605 42639 43606
rect 22576 41259 28298 41492
rect 29240 41259 34962 41492
rect 22576 39846 28299 41259
rect 29240 39846 34963 41259
rect 22673 39845 28299 39846
rect 29337 39845 34963 39846
rect 37374 37499 40348 37732
rect 37374 36086 40349 37499
rect 37471 36085 40349 36086
rect 37374 29979 40348 30212
rect 37374 28566 40349 29979
rect 37471 28565 40349 28566
rect 24732 18699 52438 18932
rect 24732 17286 52439 18699
rect 24829 17285 52439 17286
<< pwell >>
rect 21718 47836 22386 48068
rect 23892 47646 24460 48498
rect 23832 47126 23924 47298
rect 14092 43886 14660 44738
rect 42960 44769 52340 44922
rect 42960 43735 43113 44769
rect 44147 43735 44453 44769
rect 45487 43735 45793 44769
rect 46827 43735 47133 44769
rect 48167 43735 48473 44769
rect 49507 43735 49813 44769
rect 50847 43735 51153 44769
rect 52187 43735 52340 44769
rect 42960 43582 52340 43735
rect 14032 43366 14124 43538
rect 41784 41009 52504 41162
rect 37250 40126 41482 40978
rect 41784 39975 41937 41009
rect 42971 39975 43277 41009
rect 44311 39975 44617 41009
rect 45651 39975 45957 41009
rect 46991 39975 47297 41009
rect 48331 39975 48637 41009
rect 49671 39975 49977 41009
rect 51011 39975 51317 41009
rect 52351 39975 52504 41009
rect 41784 39822 52504 39975
rect 37190 39606 37282 39778
rect 38250 39606 38422 39708
rect 39550 39606 39722 39708
rect 11992 37249 13332 37402
rect 11992 36215 12145 37249
rect 13179 36215 13332 37249
rect 14564 36556 15232 36788
rect 17308 36556 17976 36788
rect 20340 36556 21008 36788
rect 23384 36556 24052 36788
rect 25392 36366 29624 37218
rect 11992 36062 13332 36215
rect 41784 37249 52504 37402
rect 41784 36215 41937 37249
rect 42971 36215 43277 37249
rect 44311 36215 44617 37249
rect 45651 36215 45957 37249
rect 46991 36215 47297 37249
rect 48331 36215 48637 37249
rect 49671 36215 49977 37249
rect 51011 36215 51317 37249
rect 52351 36215 52504 37249
rect 41784 36062 52504 36215
rect 25332 35846 25424 36018
rect 26392 35846 26564 35948
rect 27692 35846 27864 35948
rect 41784 33489 52504 33642
rect 20150 32796 20818 33028
rect 23182 32796 23850 33028
rect 41784 32455 41937 33489
rect 42971 32455 43277 33489
rect 44311 32455 44617 33489
rect 45651 32455 45957 33489
rect 46991 32455 47297 33489
rect 48331 32455 48637 33489
rect 49671 32455 49977 33489
rect 51011 32455 51317 33489
rect 52351 32455 52504 33489
rect 41784 32302 52504 32455
rect 17406 29036 18074 29268
rect 20150 29036 20818 29268
rect 22894 29036 23562 29268
rect 28088 29036 28756 29268
rect 41784 29729 52504 29882
rect 41784 28695 41937 29729
rect 42971 28695 43277 29729
rect 44311 28695 44617 29729
rect 45651 28695 45957 29729
rect 46991 28695 47297 29729
rect 48331 28695 48637 29729
rect 49671 28695 49977 29729
rect 51011 28695 51317 29729
rect 52351 28695 52504 29729
rect 41784 28542 52504 28695
rect 23286 25276 23954 25508
rect 25392 25086 29624 25938
rect 38280 25276 38948 25508
rect 41024 25276 41692 25508
rect 43768 25276 44436 25508
rect 46512 25276 47180 25508
rect 49256 25276 49924 25508
rect 25332 24566 25424 24738
rect 26392 24566 26564 24668
rect 27692 24566 27864 24668
rect 24756 21516 25424 21748
rect 28088 21516 28756 21748
rect 30832 21516 31500 21748
rect 34066 21516 34734 21748
rect 38280 21516 38948 21748
rect 41024 21516 41692 21748
rect 49256 21516 49924 21748
rect 44748 13996 45416 14228
rect 47492 13996 48160 14228
rect 50236 13996 50904 14228
rect 44650 10236 45318 10468
rect 47394 10236 48062 10468
rect 50138 10236 50806 10468
rect 45434 6476 46102 6708
rect 48178 6476 48846 6708
rect 50922 6476 51590 6708
<< nbase >>
rect 43113 43735 44147 44769
rect 44453 43735 45487 44769
rect 45793 43735 46827 44769
rect 47133 43735 48167 44769
rect 48473 43735 49507 44769
rect 49813 43735 50847 44769
rect 51153 43735 52187 44769
rect 41937 39975 42971 41009
rect 43277 39975 44311 41009
rect 44617 39975 45651 41009
rect 45957 39975 46991 41009
rect 47297 39975 48331 41009
rect 48637 39975 49671 41009
rect 49977 39975 51011 41009
rect 51317 39975 52351 41009
rect 12145 36215 13179 37249
rect 41937 36215 42971 37249
rect 43277 36215 44311 37249
rect 44617 36215 45651 37249
rect 45957 36215 46991 37249
rect 47297 36215 48331 37249
rect 48637 36215 49671 37249
rect 49977 36215 51011 37249
rect 51317 36215 52351 37249
rect 41937 32455 42971 33489
rect 43277 32455 44311 33489
rect 44617 32455 45651 33489
rect 45957 32455 46991 33489
rect 47297 32455 48331 33489
rect 48637 32455 49671 33489
rect 49977 32455 51011 33489
rect 51317 32455 52351 33489
rect 41937 28695 42971 29729
rect 43277 28695 44311 29729
rect 44617 28695 45651 29729
rect 45957 28695 46991 29729
rect 47297 28695 48331 29729
rect 48637 28695 49671 29729
rect 49977 28695 51011 29729
rect 51317 28695 52351 29729
<< pmoslvt >>
rect 24923 47427 25323 48717
rect 25381 47427 25781 48717
rect 25839 47427 26239 48717
rect 26297 47427 26697 48717
rect 26755 47427 27155 48717
rect 27213 47427 27613 48717
rect 27671 47427 28071 48717
rect 28129 47427 28529 48717
rect 28587 47427 28987 48717
rect 29045 47427 29445 48717
rect 29503 47427 29903 48717
rect 29961 47427 30361 48717
rect 30419 47427 30819 48717
rect 30877 47427 31277 48717
rect 31335 47427 31735 48717
rect 31793 47427 32193 48717
rect 32251 47427 32651 48717
rect 32709 47427 33109 48717
rect 33167 47427 33567 48717
rect 33625 47427 34025 48717
rect 34083 47427 34483 48717
rect 34541 47427 34941 48717
rect 34999 47427 35399 48717
rect 35457 47427 35857 48717
rect 35915 47427 36315 48717
rect 36373 47427 36773 48717
rect 36831 47427 37231 48717
rect 37289 47427 37689 48717
rect 37747 47427 38147 48717
rect 38205 47427 38605 48717
rect 38663 47427 39063 48717
rect 39121 47427 39521 48717
rect 39579 47427 39979 48717
rect 40037 47427 40437 48717
rect 40495 47427 40895 48717
rect 40953 47427 41353 48717
rect 41411 47427 41811 48717
rect 41869 47427 42269 48717
rect 42327 47427 42727 48717
rect 42785 47427 43185 48717
rect 43243 47427 43643 48717
rect 43701 47427 44101 48717
rect 44159 47427 44559 48717
rect 44617 47427 45017 48717
rect 45075 47427 45475 48717
rect 45533 47427 45933 48717
rect 45991 47427 46391 48717
rect 46449 47427 46849 48717
rect 46907 47427 47307 48717
rect 47365 47427 47765 48717
rect 47823 47427 48223 48717
rect 48281 47427 48681 48717
rect 48739 47427 49139 48717
rect 49197 47427 49597 48717
rect 49655 47427 50055 48717
rect 50113 47427 50513 48717
rect 50571 47427 50971 48717
rect 51029 47427 51429 48717
rect 51487 47427 51887 48717
rect 51945 47427 52345 48717
rect 15123 43667 15523 44957
rect 15581 43667 15981 44957
rect 16039 43667 16439 44957
rect 16497 43667 16897 44957
rect 16955 43667 17355 44957
rect 17413 43667 17813 44957
rect 17871 43667 18271 44957
rect 18329 43667 18729 44957
rect 18787 43667 19187 44957
rect 19245 43667 19645 44957
rect 19703 43667 20103 44957
rect 20161 43667 20561 44957
rect 20619 43667 21019 44957
rect 21077 43667 21477 44957
rect 21535 43667 21935 44957
rect 21993 43667 22393 44957
rect 22451 43667 22851 44957
rect 22909 43667 23309 44957
rect 23367 43667 23767 44957
rect 23825 43667 24225 44957
rect 24283 43667 24683 44957
rect 24741 43667 25141 44957
rect 25199 43667 25599 44957
rect 25657 43667 26057 44957
rect 26115 43667 26515 44957
rect 26573 43667 26973 44957
rect 27031 43667 27431 44957
rect 27489 43667 27889 44957
rect 27947 43667 28347 44957
rect 28405 43667 28805 44957
rect 28863 43667 29263 44957
rect 29321 43667 29721 44957
rect 29779 43667 30179 44957
rect 30237 43667 30637 44957
rect 30695 43667 31095 44957
rect 31153 43667 31553 44957
rect 31611 43667 32011 44957
rect 32069 43667 32469 44957
rect 32527 43667 32927 44957
rect 32985 43667 33385 44957
rect 33443 43667 33843 44957
rect 33901 43667 34301 44957
rect 34359 43667 34759 44957
rect 34817 43667 35217 44957
rect 35275 43667 35675 44957
rect 35733 43667 36133 44957
rect 36191 43667 36591 44957
rect 36649 43667 37049 44957
rect 37107 43667 37507 44957
rect 37565 43667 37965 44957
rect 38023 43667 38423 44957
rect 38481 43667 38881 44957
rect 38939 43667 39339 44957
rect 39397 43667 39797 44957
rect 39855 43667 40255 44957
rect 40313 43667 40713 44957
rect 40771 43667 41171 44957
rect 41229 43667 41629 44957
rect 41687 43667 42087 44957
rect 42145 43667 42545 44957
rect 22767 39907 23167 41197
rect 23225 39907 23625 41197
rect 23683 39907 24083 41197
rect 24141 39907 24541 41197
rect 24599 39907 24999 41197
rect 25057 39907 25457 41197
rect 25515 39907 25915 41197
rect 25973 39907 26373 41197
rect 26431 39907 26831 41197
rect 26889 39907 27289 41197
rect 27347 39907 27747 41197
rect 27805 39907 28205 41197
rect 29431 39907 29831 41197
rect 29889 39907 30289 41197
rect 30347 39907 30747 41197
rect 30805 39907 31205 41197
rect 31263 39907 31663 41197
rect 31721 39907 32121 41197
rect 32179 39907 32579 41197
rect 32637 39907 33037 41197
rect 33095 39907 33495 41197
rect 33553 39907 33953 41197
rect 34011 39907 34411 41197
rect 34469 39907 34869 41197
rect 37565 36147 37965 37437
rect 38023 36147 38423 37437
rect 38481 36147 38881 37437
rect 38939 36147 39339 37437
rect 39397 36147 39797 37437
rect 39855 36147 40255 37437
rect 37565 28627 37965 29917
rect 38023 28627 38423 29917
rect 38481 28627 38881 29917
rect 38939 28627 39339 29917
rect 39397 28627 39797 29917
rect 39855 28627 40255 29917
rect 24923 17347 25323 18637
rect 25381 17347 25781 18637
rect 25839 17347 26239 18637
rect 26297 17347 26697 18637
rect 26755 17347 27155 18637
rect 27213 17347 27613 18637
rect 27671 17347 28071 18637
rect 28129 17347 28529 18637
rect 28587 17347 28987 18637
rect 29045 17347 29445 18637
rect 29503 17347 29903 18637
rect 29961 17347 30361 18637
rect 30419 17347 30819 18637
rect 30877 17347 31277 18637
rect 31335 17347 31735 18637
rect 31793 17347 32193 18637
rect 32251 17347 32651 18637
rect 32709 17347 33109 18637
rect 33167 17347 33567 18637
rect 33625 17347 34025 18637
rect 34083 17347 34483 18637
rect 34541 17347 34941 18637
rect 34999 17347 35399 18637
rect 35457 17347 35857 18637
rect 35915 17347 36315 18637
rect 36373 17347 36773 18637
rect 36831 17347 37231 18637
rect 37289 17347 37689 18637
rect 37747 17347 38147 18637
rect 38205 17347 38605 18637
rect 38663 17347 39063 18637
rect 39121 17347 39521 18637
rect 39579 17347 39979 18637
rect 40037 17347 40437 18637
rect 40495 17347 40895 18637
rect 40953 17347 41353 18637
rect 41411 17347 41811 18637
rect 41869 17347 42269 18637
rect 42327 17347 42727 18637
rect 42785 17347 43185 18637
rect 43243 17347 43643 18637
rect 43701 17347 44101 18637
rect 44159 17347 44559 18637
rect 44617 17347 45017 18637
rect 45075 17347 45475 18637
rect 45533 17347 45933 18637
rect 45991 17347 46391 18637
rect 46449 17347 46849 18637
rect 46907 17347 47307 18637
rect 47365 17347 47765 18637
rect 47823 17347 48223 18637
rect 48281 17347 48681 18637
rect 48739 17347 49139 18637
rect 49197 17347 49597 18637
rect 49655 17347 50055 18637
rect 50113 17347 50513 18637
rect 50571 17347 50971 18637
rect 51029 17347 51429 18637
rect 51487 17347 51887 18637
rect 51945 17347 52345 18637
<< nmoslvt >>
rect 23976 47672 24376 48472
rect 14176 43912 14576 44712
rect 37334 40152 37734 40952
rect 37792 40152 38192 40952
rect 38250 40152 38650 40952
rect 38708 40152 39108 40952
rect 39166 40152 39566 40952
rect 39624 40152 40024 40952
rect 40082 40152 40482 40952
rect 40540 40152 40940 40952
rect 40998 40152 41398 40952
rect 25476 36392 25876 37192
rect 25934 36392 26334 37192
rect 26392 36392 26792 37192
rect 26850 36392 27250 37192
rect 27308 36392 27708 37192
rect 27766 36392 28166 37192
rect 28224 36392 28624 37192
rect 28682 36392 29082 37192
rect 29140 36392 29540 37192
rect 25476 25112 25876 25912
rect 25934 25112 26334 25912
rect 26392 25112 26792 25912
rect 26850 25112 27250 25912
rect 27308 25112 27708 25912
rect 27766 25112 28166 25912
rect 28224 25112 28624 25912
rect 28682 25112 29082 25912
rect 29140 25112 29540 25912
<< ndiff >>
rect 23918 48429 23976 48472
rect 23918 48395 23930 48429
rect 23964 48395 23976 48429
rect 23918 48361 23976 48395
rect 23918 48327 23930 48361
rect 23964 48327 23976 48361
rect 23918 48293 23976 48327
rect 23918 48259 23930 48293
rect 23964 48259 23976 48293
rect 23918 48225 23976 48259
rect 23918 48191 23930 48225
rect 23964 48191 23976 48225
rect 23918 48157 23976 48191
rect 23918 48123 23930 48157
rect 23964 48123 23976 48157
rect 23918 48089 23976 48123
rect 23918 48055 23930 48089
rect 23964 48055 23976 48089
rect 23918 48021 23976 48055
rect 23918 47987 23930 48021
rect 23964 47987 23976 48021
rect 23918 47953 23976 47987
rect 23918 47919 23930 47953
rect 23964 47919 23976 47953
rect 23918 47885 23976 47919
rect 23918 47851 23930 47885
rect 23964 47851 23976 47885
rect 23918 47817 23976 47851
rect 23918 47783 23930 47817
rect 23964 47783 23976 47817
rect 23918 47749 23976 47783
rect 23918 47715 23930 47749
rect 23964 47715 23976 47749
rect 23918 47672 23976 47715
rect 24376 48429 24434 48472
rect 24376 48395 24388 48429
rect 24422 48395 24434 48429
rect 24376 48361 24434 48395
rect 24376 48327 24388 48361
rect 24422 48327 24434 48361
rect 24376 48293 24434 48327
rect 24376 48259 24388 48293
rect 24422 48259 24434 48293
rect 24376 48225 24434 48259
rect 24376 48191 24388 48225
rect 24422 48191 24434 48225
rect 24376 48157 24434 48191
rect 24376 48123 24388 48157
rect 24422 48123 24434 48157
rect 24376 48089 24434 48123
rect 24376 48055 24388 48089
rect 24422 48055 24434 48089
rect 24376 48021 24434 48055
rect 24376 47987 24388 48021
rect 24422 47987 24434 48021
rect 24376 47953 24434 47987
rect 24376 47919 24388 47953
rect 24422 47919 24434 47953
rect 24376 47885 24434 47919
rect 24376 47851 24388 47885
rect 24422 47851 24434 47885
rect 24376 47817 24434 47851
rect 24376 47783 24388 47817
rect 24422 47783 24434 47817
rect 24376 47749 24434 47783
rect 24376 47715 24388 47749
rect 24422 47715 24434 47749
rect 24376 47672 24434 47715
rect 14118 44669 14176 44712
rect 14118 44635 14130 44669
rect 14164 44635 14176 44669
rect 14118 44601 14176 44635
rect 14118 44567 14130 44601
rect 14164 44567 14176 44601
rect 14118 44533 14176 44567
rect 14118 44499 14130 44533
rect 14164 44499 14176 44533
rect 14118 44465 14176 44499
rect 14118 44431 14130 44465
rect 14164 44431 14176 44465
rect 14118 44397 14176 44431
rect 14118 44363 14130 44397
rect 14164 44363 14176 44397
rect 14118 44329 14176 44363
rect 14118 44295 14130 44329
rect 14164 44295 14176 44329
rect 14118 44261 14176 44295
rect 14118 44227 14130 44261
rect 14164 44227 14176 44261
rect 14118 44193 14176 44227
rect 14118 44159 14130 44193
rect 14164 44159 14176 44193
rect 14118 44125 14176 44159
rect 14118 44091 14130 44125
rect 14164 44091 14176 44125
rect 14118 44057 14176 44091
rect 14118 44023 14130 44057
rect 14164 44023 14176 44057
rect 14118 43989 14176 44023
rect 14118 43955 14130 43989
rect 14164 43955 14176 43989
rect 14118 43912 14176 43955
rect 14576 44669 14634 44712
rect 14576 44635 14588 44669
rect 14622 44635 14634 44669
rect 14576 44601 14634 44635
rect 14576 44567 14588 44601
rect 14622 44567 14634 44601
rect 14576 44533 14634 44567
rect 14576 44499 14588 44533
rect 14622 44499 14634 44533
rect 14576 44465 14634 44499
rect 14576 44431 14588 44465
rect 14622 44431 14634 44465
rect 14576 44397 14634 44431
rect 14576 44363 14588 44397
rect 14622 44363 14634 44397
rect 14576 44329 14634 44363
rect 14576 44295 14588 44329
rect 14622 44295 14634 44329
rect 14576 44261 14634 44295
rect 14576 44227 14588 44261
rect 14622 44227 14634 44261
rect 14576 44193 14634 44227
rect 14576 44159 14588 44193
rect 14622 44159 14634 44193
rect 14576 44125 14634 44159
rect 14576 44091 14588 44125
rect 14622 44091 14634 44125
rect 14576 44057 14634 44091
rect 14576 44023 14588 44057
rect 14622 44023 14634 44057
rect 14576 43989 14634 44023
rect 14576 43955 14588 43989
rect 14622 43955 14634 43989
rect 14576 43912 14634 43955
rect 37276 40909 37334 40952
rect 37276 40875 37288 40909
rect 37322 40875 37334 40909
rect 37276 40841 37334 40875
rect 37276 40807 37288 40841
rect 37322 40807 37334 40841
rect 37276 40773 37334 40807
rect 37276 40739 37288 40773
rect 37322 40739 37334 40773
rect 37276 40705 37334 40739
rect 37276 40671 37288 40705
rect 37322 40671 37334 40705
rect 37276 40637 37334 40671
rect 37276 40603 37288 40637
rect 37322 40603 37334 40637
rect 37276 40569 37334 40603
rect 37276 40535 37288 40569
rect 37322 40535 37334 40569
rect 37276 40501 37334 40535
rect 37276 40467 37288 40501
rect 37322 40467 37334 40501
rect 37276 40433 37334 40467
rect 37276 40399 37288 40433
rect 37322 40399 37334 40433
rect 37276 40365 37334 40399
rect 37276 40331 37288 40365
rect 37322 40331 37334 40365
rect 37276 40297 37334 40331
rect 37276 40263 37288 40297
rect 37322 40263 37334 40297
rect 37276 40229 37334 40263
rect 37276 40195 37288 40229
rect 37322 40195 37334 40229
rect 37276 40152 37334 40195
rect 37734 40909 37792 40952
rect 37734 40875 37746 40909
rect 37780 40875 37792 40909
rect 37734 40841 37792 40875
rect 37734 40807 37746 40841
rect 37780 40807 37792 40841
rect 37734 40773 37792 40807
rect 37734 40739 37746 40773
rect 37780 40739 37792 40773
rect 37734 40705 37792 40739
rect 37734 40671 37746 40705
rect 37780 40671 37792 40705
rect 37734 40637 37792 40671
rect 37734 40603 37746 40637
rect 37780 40603 37792 40637
rect 37734 40569 37792 40603
rect 37734 40535 37746 40569
rect 37780 40535 37792 40569
rect 37734 40501 37792 40535
rect 37734 40467 37746 40501
rect 37780 40467 37792 40501
rect 37734 40433 37792 40467
rect 37734 40399 37746 40433
rect 37780 40399 37792 40433
rect 37734 40365 37792 40399
rect 37734 40331 37746 40365
rect 37780 40331 37792 40365
rect 37734 40297 37792 40331
rect 37734 40263 37746 40297
rect 37780 40263 37792 40297
rect 37734 40229 37792 40263
rect 37734 40195 37746 40229
rect 37780 40195 37792 40229
rect 37734 40152 37792 40195
rect 38192 40909 38250 40952
rect 38192 40875 38204 40909
rect 38238 40875 38250 40909
rect 38192 40841 38250 40875
rect 38192 40807 38204 40841
rect 38238 40807 38250 40841
rect 38192 40773 38250 40807
rect 38192 40739 38204 40773
rect 38238 40739 38250 40773
rect 38192 40705 38250 40739
rect 38192 40671 38204 40705
rect 38238 40671 38250 40705
rect 38192 40637 38250 40671
rect 38192 40603 38204 40637
rect 38238 40603 38250 40637
rect 38192 40569 38250 40603
rect 38192 40535 38204 40569
rect 38238 40535 38250 40569
rect 38192 40501 38250 40535
rect 38192 40467 38204 40501
rect 38238 40467 38250 40501
rect 38192 40433 38250 40467
rect 38192 40399 38204 40433
rect 38238 40399 38250 40433
rect 38192 40365 38250 40399
rect 38192 40331 38204 40365
rect 38238 40331 38250 40365
rect 38192 40297 38250 40331
rect 38192 40263 38204 40297
rect 38238 40263 38250 40297
rect 38192 40229 38250 40263
rect 38192 40195 38204 40229
rect 38238 40195 38250 40229
rect 38192 40152 38250 40195
rect 38650 40909 38708 40952
rect 38650 40875 38662 40909
rect 38696 40875 38708 40909
rect 38650 40841 38708 40875
rect 38650 40807 38662 40841
rect 38696 40807 38708 40841
rect 38650 40773 38708 40807
rect 38650 40739 38662 40773
rect 38696 40739 38708 40773
rect 38650 40705 38708 40739
rect 38650 40671 38662 40705
rect 38696 40671 38708 40705
rect 38650 40637 38708 40671
rect 38650 40603 38662 40637
rect 38696 40603 38708 40637
rect 38650 40569 38708 40603
rect 38650 40535 38662 40569
rect 38696 40535 38708 40569
rect 38650 40501 38708 40535
rect 38650 40467 38662 40501
rect 38696 40467 38708 40501
rect 38650 40433 38708 40467
rect 38650 40399 38662 40433
rect 38696 40399 38708 40433
rect 38650 40365 38708 40399
rect 38650 40331 38662 40365
rect 38696 40331 38708 40365
rect 38650 40297 38708 40331
rect 38650 40263 38662 40297
rect 38696 40263 38708 40297
rect 38650 40229 38708 40263
rect 38650 40195 38662 40229
rect 38696 40195 38708 40229
rect 38650 40152 38708 40195
rect 39108 40909 39166 40952
rect 39108 40875 39120 40909
rect 39154 40875 39166 40909
rect 39108 40841 39166 40875
rect 39108 40807 39120 40841
rect 39154 40807 39166 40841
rect 39108 40773 39166 40807
rect 39108 40739 39120 40773
rect 39154 40739 39166 40773
rect 39108 40705 39166 40739
rect 39108 40671 39120 40705
rect 39154 40671 39166 40705
rect 39108 40637 39166 40671
rect 39108 40603 39120 40637
rect 39154 40603 39166 40637
rect 39108 40569 39166 40603
rect 39108 40535 39120 40569
rect 39154 40535 39166 40569
rect 39108 40501 39166 40535
rect 39108 40467 39120 40501
rect 39154 40467 39166 40501
rect 39108 40433 39166 40467
rect 39108 40399 39120 40433
rect 39154 40399 39166 40433
rect 39108 40365 39166 40399
rect 39108 40331 39120 40365
rect 39154 40331 39166 40365
rect 39108 40297 39166 40331
rect 39108 40263 39120 40297
rect 39154 40263 39166 40297
rect 39108 40229 39166 40263
rect 39108 40195 39120 40229
rect 39154 40195 39166 40229
rect 39108 40152 39166 40195
rect 39566 40909 39624 40952
rect 39566 40875 39578 40909
rect 39612 40875 39624 40909
rect 39566 40841 39624 40875
rect 39566 40807 39578 40841
rect 39612 40807 39624 40841
rect 39566 40773 39624 40807
rect 39566 40739 39578 40773
rect 39612 40739 39624 40773
rect 39566 40705 39624 40739
rect 39566 40671 39578 40705
rect 39612 40671 39624 40705
rect 39566 40637 39624 40671
rect 39566 40603 39578 40637
rect 39612 40603 39624 40637
rect 39566 40569 39624 40603
rect 39566 40535 39578 40569
rect 39612 40535 39624 40569
rect 39566 40501 39624 40535
rect 39566 40467 39578 40501
rect 39612 40467 39624 40501
rect 39566 40433 39624 40467
rect 39566 40399 39578 40433
rect 39612 40399 39624 40433
rect 39566 40365 39624 40399
rect 39566 40331 39578 40365
rect 39612 40331 39624 40365
rect 39566 40297 39624 40331
rect 39566 40263 39578 40297
rect 39612 40263 39624 40297
rect 39566 40229 39624 40263
rect 39566 40195 39578 40229
rect 39612 40195 39624 40229
rect 39566 40152 39624 40195
rect 40024 40909 40082 40952
rect 40024 40875 40036 40909
rect 40070 40875 40082 40909
rect 40024 40841 40082 40875
rect 40024 40807 40036 40841
rect 40070 40807 40082 40841
rect 40024 40773 40082 40807
rect 40024 40739 40036 40773
rect 40070 40739 40082 40773
rect 40024 40705 40082 40739
rect 40024 40671 40036 40705
rect 40070 40671 40082 40705
rect 40024 40637 40082 40671
rect 40024 40603 40036 40637
rect 40070 40603 40082 40637
rect 40024 40569 40082 40603
rect 40024 40535 40036 40569
rect 40070 40535 40082 40569
rect 40024 40501 40082 40535
rect 40024 40467 40036 40501
rect 40070 40467 40082 40501
rect 40024 40433 40082 40467
rect 40024 40399 40036 40433
rect 40070 40399 40082 40433
rect 40024 40365 40082 40399
rect 40024 40331 40036 40365
rect 40070 40331 40082 40365
rect 40024 40297 40082 40331
rect 40024 40263 40036 40297
rect 40070 40263 40082 40297
rect 40024 40229 40082 40263
rect 40024 40195 40036 40229
rect 40070 40195 40082 40229
rect 40024 40152 40082 40195
rect 40482 40909 40540 40952
rect 40482 40875 40494 40909
rect 40528 40875 40540 40909
rect 40482 40841 40540 40875
rect 40482 40807 40494 40841
rect 40528 40807 40540 40841
rect 40482 40773 40540 40807
rect 40482 40739 40494 40773
rect 40528 40739 40540 40773
rect 40482 40705 40540 40739
rect 40482 40671 40494 40705
rect 40528 40671 40540 40705
rect 40482 40637 40540 40671
rect 40482 40603 40494 40637
rect 40528 40603 40540 40637
rect 40482 40569 40540 40603
rect 40482 40535 40494 40569
rect 40528 40535 40540 40569
rect 40482 40501 40540 40535
rect 40482 40467 40494 40501
rect 40528 40467 40540 40501
rect 40482 40433 40540 40467
rect 40482 40399 40494 40433
rect 40528 40399 40540 40433
rect 40482 40365 40540 40399
rect 40482 40331 40494 40365
rect 40528 40331 40540 40365
rect 40482 40297 40540 40331
rect 40482 40263 40494 40297
rect 40528 40263 40540 40297
rect 40482 40229 40540 40263
rect 40482 40195 40494 40229
rect 40528 40195 40540 40229
rect 40482 40152 40540 40195
rect 40940 40909 40998 40952
rect 40940 40875 40952 40909
rect 40986 40875 40998 40909
rect 40940 40841 40998 40875
rect 40940 40807 40952 40841
rect 40986 40807 40998 40841
rect 40940 40773 40998 40807
rect 40940 40739 40952 40773
rect 40986 40739 40998 40773
rect 40940 40705 40998 40739
rect 40940 40671 40952 40705
rect 40986 40671 40998 40705
rect 40940 40637 40998 40671
rect 40940 40603 40952 40637
rect 40986 40603 40998 40637
rect 40940 40569 40998 40603
rect 40940 40535 40952 40569
rect 40986 40535 40998 40569
rect 40940 40501 40998 40535
rect 40940 40467 40952 40501
rect 40986 40467 40998 40501
rect 40940 40433 40998 40467
rect 40940 40399 40952 40433
rect 40986 40399 40998 40433
rect 40940 40365 40998 40399
rect 40940 40331 40952 40365
rect 40986 40331 40998 40365
rect 40940 40297 40998 40331
rect 40940 40263 40952 40297
rect 40986 40263 40998 40297
rect 40940 40229 40998 40263
rect 40940 40195 40952 40229
rect 40986 40195 40998 40229
rect 40940 40152 40998 40195
rect 41398 40909 41456 40952
rect 41398 40875 41410 40909
rect 41444 40875 41456 40909
rect 41398 40841 41456 40875
rect 41398 40807 41410 40841
rect 41444 40807 41456 40841
rect 41398 40773 41456 40807
rect 41398 40739 41410 40773
rect 41444 40739 41456 40773
rect 41398 40705 41456 40739
rect 41398 40671 41410 40705
rect 41444 40671 41456 40705
rect 41398 40637 41456 40671
rect 41398 40603 41410 40637
rect 41444 40603 41456 40637
rect 41398 40569 41456 40603
rect 41398 40535 41410 40569
rect 41444 40535 41456 40569
rect 41398 40501 41456 40535
rect 41398 40467 41410 40501
rect 41444 40467 41456 40501
rect 41398 40433 41456 40467
rect 41398 40399 41410 40433
rect 41444 40399 41456 40433
rect 41398 40365 41456 40399
rect 41398 40331 41410 40365
rect 41444 40331 41456 40365
rect 41398 40297 41456 40331
rect 41398 40263 41410 40297
rect 41444 40263 41456 40297
rect 41398 40229 41456 40263
rect 41398 40195 41410 40229
rect 41444 40195 41456 40229
rect 41398 40152 41456 40195
rect 25418 37149 25476 37192
rect 25418 37115 25430 37149
rect 25464 37115 25476 37149
rect 25418 37081 25476 37115
rect 25418 37047 25430 37081
rect 25464 37047 25476 37081
rect 25418 37013 25476 37047
rect 25418 36979 25430 37013
rect 25464 36979 25476 37013
rect 25418 36945 25476 36979
rect 25418 36911 25430 36945
rect 25464 36911 25476 36945
rect 25418 36877 25476 36911
rect 25418 36843 25430 36877
rect 25464 36843 25476 36877
rect 25418 36809 25476 36843
rect 25418 36775 25430 36809
rect 25464 36775 25476 36809
rect 25418 36741 25476 36775
rect 25418 36707 25430 36741
rect 25464 36707 25476 36741
rect 25418 36673 25476 36707
rect 25418 36639 25430 36673
rect 25464 36639 25476 36673
rect 25418 36605 25476 36639
rect 25418 36571 25430 36605
rect 25464 36571 25476 36605
rect 25418 36537 25476 36571
rect 25418 36503 25430 36537
rect 25464 36503 25476 36537
rect 25418 36469 25476 36503
rect 25418 36435 25430 36469
rect 25464 36435 25476 36469
rect 25418 36392 25476 36435
rect 25876 37149 25934 37192
rect 25876 37115 25888 37149
rect 25922 37115 25934 37149
rect 25876 37081 25934 37115
rect 25876 37047 25888 37081
rect 25922 37047 25934 37081
rect 25876 37013 25934 37047
rect 25876 36979 25888 37013
rect 25922 36979 25934 37013
rect 25876 36945 25934 36979
rect 25876 36911 25888 36945
rect 25922 36911 25934 36945
rect 25876 36877 25934 36911
rect 25876 36843 25888 36877
rect 25922 36843 25934 36877
rect 25876 36809 25934 36843
rect 25876 36775 25888 36809
rect 25922 36775 25934 36809
rect 25876 36741 25934 36775
rect 25876 36707 25888 36741
rect 25922 36707 25934 36741
rect 25876 36673 25934 36707
rect 25876 36639 25888 36673
rect 25922 36639 25934 36673
rect 25876 36605 25934 36639
rect 25876 36571 25888 36605
rect 25922 36571 25934 36605
rect 25876 36537 25934 36571
rect 25876 36503 25888 36537
rect 25922 36503 25934 36537
rect 25876 36469 25934 36503
rect 25876 36435 25888 36469
rect 25922 36435 25934 36469
rect 25876 36392 25934 36435
rect 26334 37149 26392 37192
rect 26334 37115 26346 37149
rect 26380 37115 26392 37149
rect 26334 37081 26392 37115
rect 26334 37047 26346 37081
rect 26380 37047 26392 37081
rect 26334 37013 26392 37047
rect 26334 36979 26346 37013
rect 26380 36979 26392 37013
rect 26334 36945 26392 36979
rect 26334 36911 26346 36945
rect 26380 36911 26392 36945
rect 26334 36877 26392 36911
rect 26334 36843 26346 36877
rect 26380 36843 26392 36877
rect 26334 36809 26392 36843
rect 26334 36775 26346 36809
rect 26380 36775 26392 36809
rect 26334 36741 26392 36775
rect 26334 36707 26346 36741
rect 26380 36707 26392 36741
rect 26334 36673 26392 36707
rect 26334 36639 26346 36673
rect 26380 36639 26392 36673
rect 26334 36605 26392 36639
rect 26334 36571 26346 36605
rect 26380 36571 26392 36605
rect 26334 36537 26392 36571
rect 26334 36503 26346 36537
rect 26380 36503 26392 36537
rect 26334 36469 26392 36503
rect 26334 36435 26346 36469
rect 26380 36435 26392 36469
rect 26334 36392 26392 36435
rect 26792 37149 26850 37192
rect 26792 37115 26804 37149
rect 26838 37115 26850 37149
rect 26792 37081 26850 37115
rect 26792 37047 26804 37081
rect 26838 37047 26850 37081
rect 26792 37013 26850 37047
rect 26792 36979 26804 37013
rect 26838 36979 26850 37013
rect 26792 36945 26850 36979
rect 26792 36911 26804 36945
rect 26838 36911 26850 36945
rect 26792 36877 26850 36911
rect 26792 36843 26804 36877
rect 26838 36843 26850 36877
rect 26792 36809 26850 36843
rect 26792 36775 26804 36809
rect 26838 36775 26850 36809
rect 26792 36741 26850 36775
rect 26792 36707 26804 36741
rect 26838 36707 26850 36741
rect 26792 36673 26850 36707
rect 26792 36639 26804 36673
rect 26838 36639 26850 36673
rect 26792 36605 26850 36639
rect 26792 36571 26804 36605
rect 26838 36571 26850 36605
rect 26792 36537 26850 36571
rect 26792 36503 26804 36537
rect 26838 36503 26850 36537
rect 26792 36469 26850 36503
rect 26792 36435 26804 36469
rect 26838 36435 26850 36469
rect 26792 36392 26850 36435
rect 27250 37149 27308 37192
rect 27250 37115 27262 37149
rect 27296 37115 27308 37149
rect 27250 37081 27308 37115
rect 27250 37047 27262 37081
rect 27296 37047 27308 37081
rect 27250 37013 27308 37047
rect 27250 36979 27262 37013
rect 27296 36979 27308 37013
rect 27250 36945 27308 36979
rect 27250 36911 27262 36945
rect 27296 36911 27308 36945
rect 27250 36877 27308 36911
rect 27250 36843 27262 36877
rect 27296 36843 27308 36877
rect 27250 36809 27308 36843
rect 27250 36775 27262 36809
rect 27296 36775 27308 36809
rect 27250 36741 27308 36775
rect 27250 36707 27262 36741
rect 27296 36707 27308 36741
rect 27250 36673 27308 36707
rect 27250 36639 27262 36673
rect 27296 36639 27308 36673
rect 27250 36605 27308 36639
rect 27250 36571 27262 36605
rect 27296 36571 27308 36605
rect 27250 36537 27308 36571
rect 27250 36503 27262 36537
rect 27296 36503 27308 36537
rect 27250 36469 27308 36503
rect 27250 36435 27262 36469
rect 27296 36435 27308 36469
rect 27250 36392 27308 36435
rect 27708 37149 27766 37192
rect 27708 37115 27720 37149
rect 27754 37115 27766 37149
rect 27708 37081 27766 37115
rect 27708 37047 27720 37081
rect 27754 37047 27766 37081
rect 27708 37013 27766 37047
rect 27708 36979 27720 37013
rect 27754 36979 27766 37013
rect 27708 36945 27766 36979
rect 27708 36911 27720 36945
rect 27754 36911 27766 36945
rect 27708 36877 27766 36911
rect 27708 36843 27720 36877
rect 27754 36843 27766 36877
rect 27708 36809 27766 36843
rect 27708 36775 27720 36809
rect 27754 36775 27766 36809
rect 27708 36741 27766 36775
rect 27708 36707 27720 36741
rect 27754 36707 27766 36741
rect 27708 36673 27766 36707
rect 27708 36639 27720 36673
rect 27754 36639 27766 36673
rect 27708 36605 27766 36639
rect 27708 36571 27720 36605
rect 27754 36571 27766 36605
rect 27708 36537 27766 36571
rect 27708 36503 27720 36537
rect 27754 36503 27766 36537
rect 27708 36469 27766 36503
rect 27708 36435 27720 36469
rect 27754 36435 27766 36469
rect 27708 36392 27766 36435
rect 28166 37149 28224 37192
rect 28166 37115 28178 37149
rect 28212 37115 28224 37149
rect 28166 37081 28224 37115
rect 28166 37047 28178 37081
rect 28212 37047 28224 37081
rect 28166 37013 28224 37047
rect 28166 36979 28178 37013
rect 28212 36979 28224 37013
rect 28166 36945 28224 36979
rect 28166 36911 28178 36945
rect 28212 36911 28224 36945
rect 28166 36877 28224 36911
rect 28166 36843 28178 36877
rect 28212 36843 28224 36877
rect 28166 36809 28224 36843
rect 28166 36775 28178 36809
rect 28212 36775 28224 36809
rect 28166 36741 28224 36775
rect 28166 36707 28178 36741
rect 28212 36707 28224 36741
rect 28166 36673 28224 36707
rect 28166 36639 28178 36673
rect 28212 36639 28224 36673
rect 28166 36605 28224 36639
rect 28166 36571 28178 36605
rect 28212 36571 28224 36605
rect 28166 36537 28224 36571
rect 28166 36503 28178 36537
rect 28212 36503 28224 36537
rect 28166 36469 28224 36503
rect 28166 36435 28178 36469
rect 28212 36435 28224 36469
rect 28166 36392 28224 36435
rect 28624 37149 28682 37192
rect 28624 37115 28636 37149
rect 28670 37115 28682 37149
rect 28624 37081 28682 37115
rect 28624 37047 28636 37081
rect 28670 37047 28682 37081
rect 28624 37013 28682 37047
rect 28624 36979 28636 37013
rect 28670 36979 28682 37013
rect 28624 36945 28682 36979
rect 28624 36911 28636 36945
rect 28670 36911 28682 36945
rect 28624 36877 28682 36911
rect 28624 36843 28636 36877
rect 28670 36843 28682 36877
rect 28624 36809 28682 36843
rect 28624 36775 28636 36809
rect 28670 36775 28682 36809
rect 28624 36741 28682 36775
rect 28624 36707 28636 36741
rect 28670 36707 28682 36741
rect 28624 36673 28682 36707
rect 28624 36639 28636 36673
rect 28670 36639 28682 36673
rect 28624 36605 28682 36639
rect 28624 36571 28636 36605
rect 28670 36571 28682 36605
rect 28624 36537 28682 36571
rect 28624 36503 28636 36537
rect 28670 36503 28682 36537
rect 28624 36469 28682 36503
rect 28624 36435 28636 36469
rect 28670 36435 28682 36469
rect 28624 36392 28682 36435
rect 29082 37149 29140 37192
rect 29082 37115 29094 37149
rect 29128 37115 29140 37149
rect 29082 37081 29140 37115
rect 29082 37047 29094 37081
rect 29128 37047 29140 37081
rect 29082 37013 29140 37047
rect 29082 36979 29094 37013
rect 29128 36979 29140 37013
rect 29082 36945 29140 36979
rect 29082 36911 29094 36945
rect 29128 36911 29140 36945
rect 29082 36877 29140 36911
rect 29082 36843 29094 36877
rect 29128 36843 29140 36877
rect 29082 36809 29140 36843
rect 29082 36775 29094 36809
rect 29128 36775 29140 36809
rect 29082 36741 29140 36775
rect 29082 36707 29094 36741
rect 29128 36707 29140 36741
rect 29082 36673 29140 36707
rect 29082 36639 29094 36673
rect 29128 36639 29140 36673
rect 29082 36605 29140 36639
rect 29082 36571 29094 36605
rect 29128 36571 29140 36605
rect 29082 36537 29140 36571
rect 29082 36503 29094 36537
rect 29128 36503 29140 36537
rect 29082 36469 29140 36503
rect 29082 36435 29094 36469
rect 29128 36435 29140 36469
rect 29082 36392 29140 36435
rect 29540 37149 29598 37192
rect 29540 37115 29552 37149
rect 29586 37115 29598 37149
rect 29540 37081 29598 37115
rect 29540 37047 29552 37081
rect 29586 37047 29598 37081
rect 29540 37013 29598 37047
rect 29540 36979 29552 37013
rect 29586 36979 29598 37013
rect 29540 36945 29598 36979
rect 29540 36911 29552 36945
rect 29586 36911 29598 36945
rect 29540 36877 29598 36911
rect 29540 36843 29552 36877
rect 29586 36843 29598 36877
rect 29540 36809 29598 36843
rect 29540 36775 29552 36809
rect 29586 36775 29598 36809
rect 29540 36741 29598 36775
rect 29540 36707 29552 36741
rect 29586 36707 29598 36741
rect 29540 36673 29598 36707
rect 29540 36639 29552 36673
rect 29586 36639 29598 36673
rect 29540 36605 29598 36639
rect 29540 36571 29552 36605
rect 29586 36571 29598 36605
rect 29540 36537 29598 36571
rect 29540 36503 29552 36537
rect 29586 36503 29598 36537
rect 29540 36469 29598 36503
rect 29540 36435 29552 36469
rect 29586 36435 29598 36469
rect 29540 36392 29598 36435
rect 25418 25869 25476 25912
rect 25418 25835 25430 25869
rect 25464 25835 25476 25869
rect 25418 25801 25476 25835
rect 25418 25767 25430 25801
rect 25464 25767 25476 25801
rect 25418 25733 25476 25767
rect 25418 25699 25430 25733
rect 25464 25699 25476 25733
rect 25418 25665 25476 25699
rect 25418 25631 25430 25665
rect 25464 25631 25476 25665
rect 25418 25597 25476 25631
rect 25418 25563 25430 25597
rect 25464 25563 25476 25597
rect 25418 25529 25476 25563
rect 25418 25495 25430 25529
rect 25464 25495 25476 25529
rect 25418 25461 25476 25495
rect 25418 25427 25430 25461
rect 25464 25427 25476 25461
rect 25418 25393 25476 25427
rect 25418 25359 25430 25393
rect 25464 25359 25476 25393
rect 25418 25325 25476 25359
rect 25418 25291 25430 25325
rect 25464 25291 25476 25325
rect 25418 25257 25476 25291
rect 25418 25223 25430 25257
rect 25464 25223 25476 25257
rect 25418 25189 25476 25223
rect 25418 25155 25430 25189
rect 25464 25155 25476 25189
rect 25418 25112 25476 25155
rect 25876 25869 25934 25912
rect 25876 25835 25888 25869
rect 25922 25835 25934 25869
rect 25876 25801 25934 25835
rect 25876 25767 25888 25801
rect 25922 25767 25934 25801
rect 25876 25733 25934 25767
rect 25876 25699 25888 25733
rect 25922 25699 25934 25733
rect 25876 25665 25934 25699
rect 25876 25631 25888 25665
rect 25922 25631 25934 25665
rect 25876 25597 25934 25631
rect 25876 25563 25888 25597
rect 25922 25563 25934 25597
rect 25876 25529 25934 25563
rect 25876 25495 25888 25529
rect 25922 25495 25934 25529
rect 25876 25461 25934 25495
rect 25876 25427 25888 25461
rect 25922 25427 25934 25461
rect 25876 25393 25934 25427
rect 25876 25359 25888 25393
rect 25922 25359 25934 25393
rect 25876 25325 25934 25359
rect 25876 25291 25888 25325
rect 25922 25291 25934 25325
rect 25876 25257 25934 25291
rect 25876 25223 25888 25257
rect 25922 25223 25934 25257
rect 25876 25189 25934 25223
rect 25876 25155 25888 25189
rect 25922 25155 25934 25189
rect 25876 25112 25934 25155
rect 26334 25869 26392 25912
rect 26334 25835 26346 25869
rect 26380 25835 26392 25869
rect 26334 25801 26392 25835
rect 26334 25767 26346 25801
rect 26380 25767 26392 25801
rect 26334 25733 26392 25767
rect 26334 25699 26346 25733
rect 26380 25699 26392 25733
rect 26334 25665 26392 25699
rect 26334 25631 26346 25665
rect 26380 25631 26392 25665
rect 26334 25597 26392 25631
rect 26334 25563 26346 25597
rect 26380 25563 26392 25597
rect 26334 25529 26392 25563
rect 26334 25495 26346 25529
rect 26380 25495 26392 25529
rect 26334 25461 26392 25495
rect 26334 25427 26346 25461
rect 26380 25427 26392 25461
rect 26334 25393 26392 25427
rect 26334 25359 26346 25393
rect 26380 25359 26392 25393
rect 26334 25325 26392 25359
rect 26334 25291 26346 25325
rect 26380 25291 26392 25325
rect 26334 25257 26392 25291
rect 26334 25223 26346 25257
rect 26380 25223 26392 25257
rect 26334 25189 26392 25223
rect 26334 25155 26346 25189
rect 26380 25155 26392 25189
rect 26334 25112 26392 25155
rect 26792 25869 26850 25912
rect 26792 25835 26804 25869
rect 26838 25835 26850 25869
rect 26792 25801 26850 25835
rect 26792 25767 26804 25801
rect 26838 25767 26850 25801
rect 26792 25733 26850 25767
rect 26792 25699 26804 25733
rect 26838 25699 26850 25733
rect 26792 25665 26850 25699
rect 26792 25631 26804 25665
rect 26838 25631 26850 25665
rect 26792 25597 26850 25631
rect 26792 25563 26804 25597
rect 26838 25563 26850 25597
rect 26792 25529 26850 25563
rect 26792 25495 26804 25529
rect 26838 25495 26850 25529
rect 26792 25461 26850 25495
rect 26792 25427 26804 25461
rect 26838 25427 26850 25461
rect 26792 25393 26850 25427
rect 26792 25359 26804 25393
rect 26838 25359 26850 25393
rect 26792 25325 26850 25359
rect 26792 25291 26804 25325
rect 26838 25291 26850 25325
rect 26792 25257 26850 25291
rect 26792 25223 26804 25257
rect 26838 25223 26850 25257
rect 26792 25189 26850 25223
rect 26792 25155 26804 25189
rect 26838 25155 26850 25189
rect 26792 25112 26850 25155
rect 27250 25869 27308 25912
rect 27250 25835 27262 25869
rect 27296 25835 27308 25869
rect 27250 25801 27308 25835
rect 27250 25767 27262 25801
rect 27296 25767 27308 25801
rect 27250 25733 27308 25767
rect 27250 25699 27262 25733
rect 27296 25699 27308 25733
rect 27250 25665 27308 25699
rect 27250 25631 27262 25665
rect 27296 25631 27308 25665
rect 27250 25597 27308 25631
rect 27250 25563 27262 25597
rect 27296 25563 27308 25597
rect 27250 25529 27308 25563
rect 27250 25495 27262 25529
rect 27296 25495 27308 25529
rect 27250 25461 27308 25495
rect 27250 25427 27262 25461
rect 27296 25427 27308 25461
rect 27250 25393 27308 25427
rect 27250 25359 27262 25393
rect 27296 25359 27308 25393
rect 27250 25325 27308 25359
rect 27250 25291 27262 25325
rect 27296 25291 27308 25325
rect 27250 25257 27308 25291
rect 27250 25223 27262 25257
rect 27296 25223 27308 25257
rect 27250 25189 27308 25223
rect 27250 25155 27262 25189
rect 27296 25155 27308 25189
rect 27250 25112 27308 25155
rect 27708 25869 27766 25912
rect 27708 25835 27720 25869
rect 27754 25835 27766 25869
rect 27708 25801 27766 25835
rect 27708 25767 27720 25801
rect 27754 25767 27766 25801
rect 27708 25733 27766 25767
rect 27708 25699 27720 25733
rect 27754 25699 27766 25733
rect 27708 25665 27766 25699
rect 27708 25631 27720 25665
rect 27754 25631 27766 25665
rect 27708 25597 27766 25631
rect 27708 25563 27720 25597
rect 27754 25563 27766 25597
rect 27708 25529 27766 25563
rect 27708 25495 27720 25529
rect 27754 25495 27766 25529
rect 27708 25461 27766 25495
rect 27708 25427 27720 25461
rect 27754 25427 27766 25461
rect 27708 25393 27766 25427
rect 27708 25359 27720 25393
rect 27754 25359 27766 25393
rect 27708 25325 27766 25359
rect 27708 25291 27720 25325
rect 27754 25291 27766 25325
rect 27708 25257 27766 25291
rect 27708 25223 27720 25257
rect 27754 25223 27766 25257
rect 27708 25189 27766 25223
rect 27708 25155 27720 25189
rect 27754 25155 27766 25189
rect 27708 25112 27766 25155
rect 28166 25869 28224 25912
rect 28166 25835 28178 25869
rect 28212 25835 28224 25869
rect 28166 25801 28224 25835
rect 28166 25767 28178 25801
rect 28212 25767 28224 25801
rect 28166 25733 28224 25767
rect 28166 25699 28178 25733
rect 28212 25699 28224 25733
rect 28166 25665 28224 25699
rect 28166 25631 28178 25665
rect 28212 25631 28224 25665
rect 28166 25597 28224 25631
rect 28166 25563 28178 25597
rect 28212 25563 28224 25597
rect 28166 25529 28224 25563
rect 28166 25495 28178 25529
rect 28212 25495 28224 25529
rect 28166 25461 28224 25495
rect 28166 25427 28178 25461
rect 28212 25427 28224 25461
rect 28166 25393 28224 25427
rect 28166 25359 28178 25393
rect 28212 25359 28224 25393
rect 28166 25325 28224 25359
rect 28166 25291 28178 25325
rect 28212 25291 28224 25325
rect 28166 25257 28224 25291
rect 28166 25223 28178 25257
rect 28212 25223 28224 25257
rect 28166 25189 28224 25223
rect 28166 25155 28178 25189
rect 28212 25155 28224 25189
rect 28166 25112 28224 25155
rect 28624 25869 28682 25912
rect 28624 25835 28636 25869
rect 28670 25835 28682 25869
rect 28624 25801 28682 25835
rect 28624 25767 28636 25801
rect 28670 25767 28682 25801
rect 28624 25733 28682 25767
rect 28624 25699 28636 25733
rect 28670 25699 28682 25733
rect 28624 25665 28682 25699
rect 28624 25631 28636 25665
rect 28670 25631 28682 25665
rect 28624 25597 28682 25631
rect 28624 25563 28636 25597
rect 28670 25563 28682 25597
rect 28624 25529 28682 25563
rect 28624 25495 28636 25529
rect 28670 25495 28682 25529
rect 28624 25461 28682 25495
rect 28624 25427 28636 25461
rect 28670 25427 28682 25461
rect 28624 25393 28682 25427
rect 28624 25359 28636 25393
rect 28670 25359 28682 25393
rect 28624 25325 28682 25359
rect 28624 25291 28636 25325
rect 28670 25291 28682 25325
rect 28624 25257 28682 25291
rect 28624 25223 28636 25257
rect 28670 25223 28682 25257
rect 28624 25189 28682 25223
rect 28624 25155 28636 25189
rect 28670 25155 28682 25189
rect 28624 25112 28682 25155
rect 29082 25869 29140 25912
rect 29082 25835 29094 25869
rect 29128 25835 29140 25869
rect 29082 25801 29140 25835
rect 29082 25767 29094 25801
rect 29128 25767 29140 25801
rect 29082 25733 29140 25767
rect 29082 25699 29094 25733
rect 29128 25699 29140 25733
rect 29082 25665 29140 25699
rect 29082 25631 29094 25665
rect 29128 25631 29140 25665
rect 29082 25597 29140 25631
rect 29082 25563 29094 25597
rect 29128 25563 29140 25597
rect 29082 25529 29140 25563
rect 29082 25495 29094 25529
rect 29128 25495 29140 25529
rect 29082 25461 29140 25495
rect 29082 25427 29094 25461
rect 29128 25427 29140 25461
rect 29082 25393 29140 25427
rect 29082 25359 29094 25393
rect 29128 25359 29140 25393
rect 29082 25325 29140 25359
rect 29082 25291 29094 25325
rect 29128 25291 29140 25325
rect 29082 25257 29140 25291
rect 29082 25223 29094 25257
rect 29128 25223 29140 25257
rect 29082 25189 29140 25223
rect 29082 25155 29094 25189
rect 29128 25155 29140 25189
rect 29082 25112 29140 25155
rect 29540 25869 29598 25912
rect 29540 25835 29552 25869
rect 29586 25835 29598 25869
rect 29540 25801 29598 25835
rect 29540 25767 29552 25801
rect 29586 25767 29598 25801
rect 29540 25733 29598 25767
rect 29540 25699 29552 25733
rect 29586 25699 29598 25733
rect 29540 25665 29598 25699
rect 29540 25631 29552 25665
rect 29586 25631 29598 25665
rect 29540 25597 29598 25631
rect 29540 25563 29552 25597
rect 29586 25563 29598 25597
rect 29540 25529 29598 25563
rect 29540 25495 29552 25529
rect 29586 25495 29598 25529
rect 29540 25461 29598 25495
rect 29540 25427 29552 25461
rect 29586 25427 29598 25461
rect 29540 25393 29598 25427
rect 29540 25359 29552 25393
rect 29586 25359 29598 25393
rect 29540 25325 29598 25359
rect 29540 25291 29552 25325
rect 29586 25291 29598 25325
rect 29540 25257 29598 25291
rect 29540 25223 29552 25257
rect 29586 25223 29598 25257
rect 29540 25189 29598 25223
rect 29540 25155 29552 25189
rect 29586 25155 29598 25189
rect 29540 25112 29598 25155
<< pdiff >>
rect 24865 48701 24923 48717
rect 24865 48667 24877 48701
rect 24911 48667 24923 48701
rect 24865 48633 24923 48667
rect 24865 48599 24877 48633
rect 24911 48599 24923 48633
rect 24865 48565 24923 48599
rect 24865 48531 24877 48565
rect 24911 48531 24923 48565
rect 24865 48497 24923 48531
rect 24865 48463 24877 48497
rect 24911 48463 24923 48497
rect 24865 48429 24923 48463
rect 24865 48395 24877 48429
rect 24911 48395 24923 48429
rect 24865 48361 24923 48395
rect 24865 48327 24877 48361
rect 24911 48327 24923 48361
rect 24865 48293 24923 48327
rect 24865 48259 24877 48293
rect 24911 48259 24923 48293
rect 24865 48225 24923 48259
rect 24865 48191 24877 48225
rect 24911 48191 24923 48225
rect 24865 48157 24923 48191
rect 24865 48123 24877 48157
rect 24911 48123 24923 48157
rect 24865 48089 24923 48123
rect 24865 48055 24877 48089
rect 24911 48055 24923 48089
rect 24865 48021 24923 48055
rect 24865 47987 24877 48021
rect 24911 47987 24923 48021
rect 24865 47953 24923 47987
rect 24865 47919 24877 47953
rect 24911 47919 24923 47953
rect 24865 47885 24923 47919
rect 24865 47851 24877 47885
rect 24911 47851 24923 47885
rect 24865 47817 24923 47851
rect 24865 47783 24877 47817
rect 24911 47783 24923 47817
rect 24865 47749 24923 47783
rect 24865 47715 24877 47749
rect 24911 47715 24923 47749
rect 24865 47681 24923 47715
rect 24865 47647 24877 47681
rect 24911 47647 24923 47681
rect 24865 47613 24923 47647
rect 24865 47579 24877 47613
rect 24911 47579 24923 47613
rect 24865 47545 24923 47579
rect 24865 47511 24877 47545
rect 24911 47511 24923 47545
rect 24865 47477 24923 47511
rect 24865 47443 24877 47477
rect 24911 47443 24923 47477
rect 24865 47427 24923 47443
rect 25323 48701 25381 48717
rect 25323 48667 25335 48701
rect 25369 48667 25381 48701
rect 25323 48633 25381 48667
rect 25323 48599 25335 48633
rect 25369 48599 25381 48633
rect 25323 48565 25381 48599
rect 25323 48531 25335 48565
rect 25369 48531 25381 48565
rect 25323 48497 25381 48531
rect 25323 48463 25335 48497
rect 25369 48463 25381 48497
rect 25323 48429 25381 48463
rect 25323 48395 25335 48429
rect 25369 48395 25381 48429
rect 25323 48361 25381 48395
rect 25323 48327 25335 48361
rect 25369 48327 25381 48361
rect 25323 48293 25381 48327
rect 25323 48259 25335 48293
rect 25369 48259 25381 48293
rect 25323 48225 25381 48259
rect 25323 48191 25335 48225
rect 25369 48191 25381 48225
rect 25323 48157 25381 48191
rect 25323 48123 25335 48157
rect 25369 48123 25381 48157
rect 25323 48089 25381 48123
rect 25323 48055 25335 48089
rect 25369 48055 25381 48089
rect 25323 48021 25381 48055
rect 25323 47987 25335 48021
rect 25369 47987 25381 48021
rect 25323 47953 25381 47987
rect 25323 47919 25335 47953
rect 25369 47919 25381 47953
rect 25323 47885 25381 47919
rect 25323 47851 25335 47885
rect 25369 47851 25381 47885
rect 25323 47817 25381 47851
rect 25323 47783 25335 47817
rect 25369 47783 25381 47817
rect 25323 47749 25381 47783
rect 25323 47715 25335 47749
rect 25369 47715 25381 47749
rect 25323 47681 25381 47715
rect 25323 47647 25335 47681
rect 25369 47647 25381 47681
rect 25323 47613 25381 47647
rect 25323 47579 25335 47613
rect 25369 47579 25381 47613
rect 25323 47545 25381 47579
rect 25323 47511 25335 47545
rect 25369 47511 25381 47545
rect 25323 47477 25381 47511
rect 25323 47443 25335 47477
rect 25369 47443 25381 47477
rect 25323 47427 25381 47443
rect 25781 48701 25839 48717
rect 25781 48667 25793 48701
rect 25827 48667 25839 48701
rect 25781 48633 25839 48667
rect 25781 48599 25793 48633
rect 25827 48599 25839 48633
rect 25781 48565 25839 48599
rect 25781 48531 25793 48565
rect 25827 48531 25839 48565
rect 25781 48497 25839 48531
rect 25781 48463 25793 48497
rect 25827 48463 25839 48497
rect 25781 48429 25839 48463
rect 25781 48395 25793 48429
rect 25827 48395 25839 48429
rect 25781 48361 25839 48395
rect 25781 48327 25793 48361
rect 25827 48327 25839 48361
rect 25781 48293 25839 48327
rect 25781 48259 25793 48293
rect 25827 48259 25839 48293
rect 25781 48225 25839 48259
rect 25781 48191 25793 48225
rect 25827 48191 25839 48225
rect 25781 48157 25839 48191
rect 25781 48123 25793 48157
rect 25827 48123 25839 48157
rect 25781 48089 25839 48123
rect 25781 48055 25793 48089
rect 25827 48055 25839 48089
rect 25781 48021 25839 48055
rect 25781 47987 25793 48021
rect 25827 47987 25839 48021
rect 25781 47953 25839 47987
rect 25781 47919 25793 47953
rect 25827 47919 25839 47953
rect 25781 47885 25839 47919
rect 25781 47851 25793 47885
rect 25827 47851 25839 47885
rect 25781 47817 25839 47851
rect 25781 47783 25793 47817
rect 25827 47783 25839 47817
rect 25781 47749 25839 47783
rect 25781 47715 25793 47749
rect 25827 47715 25839 47749
rect 25781 47681 25839 47715
rect 25781 47647 25793 47681
rect 25827 47647 25839 47681
rect 25781 47613 25839 47647
rect 25781 47579 25793 47613
rect 25827 47579 25839 47613
rect 25781 47545 25839 47579
rect 25781 47511 25793 47545
rect 25827 47511 25839 47545
rect 25781 47477 25839 47511
rect 25781 47443 25793 47477
rect 25827 47443 25839 47477
rect 25781 47427 25839 47443
rect 26239 48701 26297 48717
rect 26239 48667 26251 48701
rect 26285 48667 26297 48701
rect 26239 48633 26297 48667
rect 26239 48599 26251 48633
rect 26285 48599 26297 48633
rect 26239 48565 26297 48599
rect 26239 48531 26251 48565
rect 26285 48531 26297 48565
rect 26239 48497 26297 48531
rect 26239 48463 26251 48497
rect 26285 48463 26297 48497
rect 26239 48429 26297 48463
rect 26239 48395 26251 48429
rect 26285 48395 26297 48429
rect 26239 48361 26297 48395
rect 26239 48327 26251 48361
rect 26285 48327 26297 48361
rect 26239 48293 26297 48327
rect 26239 48259 26251 48293
rect 26285 48259 26297 48293
rect 26239 48225 26297 48259
rect 26239 48191 26251 48225
rect 26285 48191 26297 48225
rect 26239 48157 26297 48191
rect 26239 48123 26251 48157
rect 26285 48123 26297 48157
rect 26239 48089 26297 48123
rect 26239 48055 26251 48089
rect 26285 48055 26297 48089
rect 26239 48021 26297 48055
rect 26239 47987 26251 48021
rect 26285 47987 26297 48021
rect 26239 47953 26297 47987
rect 26239 47919 26251 47953
rect 26285 47919 26297 47953
rect 26239 47885 26297 47919
rect 26239 47851 26251 47885
rect 26285 47851 26297 47885
rect 26239 47817 26297 47851
rect 26239 47783 26251 47817
rect 26285 47783 26297 47817
rect 26239 47749 26297 47783
rect 26239 47715 26251 47749
rect 26285 47715 26297 47749
rect 26239 47681 26297 47715
rect 26239 47647 26251 47681
rect 26285 47647 26297 47681
rect 26239 47613 26297 47647
rect 26239 47579 26251 47613
rect 26285 47579 26297 47613
rect 26239 47545 26297 47579
rect 26239 47511 26251 47545
rect 26285 47511 26297 47545
rect 26239 47477 26297 47511
rect 26239 47443 26251 47477
rect 26285 47443 26297 47477
rect 26239 47427 26297 47443
rect 26697 48701 26755 48717
rect 26697 48667 26709 48701
rect 26743 48667 26755 48701
rect 26697 48633 26755 48667
rect 26697 48599 26709 48633
rect 26743 48599 26755 48633
rect 26697 48565 26755 48599
rect 26697 48531 26709 48565
rect 26743 48531 26755 48565
rect 26697 48497 26755 48531
rect 26697 48463 26709 48497
rect 26743 48463 26755 48497
rect 26697 48429 26755 48463
rect 26697 48395 26709 48429
rect 26743 48395 26755 48429
rect 26697 48361 26755 48395
rect 26697 48327 26709 48361
rect 26743 48327 26755 48361
rect 26697 48293 26755 48327
rect 26697 48259 26709 48293
rect 26743 48259 26755 48293
rect 26697 48225 26755 48259
rect 26697 48191 26709 48225
rect 26743 48191 26755 48225
rect 26697 48157 26755 48191
rect 26697 48123 26709 48157
rect 26743 48123 26755 48157
rect 26697 48089 26755 48123
rect 26697 48055 26709 48089
rect 26743 48055 26755 48089
rect 26697 48021 26755 48055
rect 26697 47987 26709 48021
rect 26743 47987 26755 48021
rect 26697 47953 26755 47987
rect 26697 47919 26709 47953
rect 26743 47919 26755 47953
rect 26697 47885 26755 47919
rect 26697 47851 26709 47885
rect 26743 47851 26755 47885
rect 26697 47817 26755 47851
rect 26697 47783 26709 47817
rect 26743 47783 26755 47817
rect 26697 47749 26755 47783
rect 26697 47715 26709 47749
rect 26743 47715 26755 47749
rect 26697 47681 26755 47715
rect 26697 47647 26709 47681
rect 26743 47647 26755 47681
rect 26697 47613 26755 47647
rect 26697 47579 26709 47613
rect 26743 47579 26755 47613
rect 26697 47545 26755 47579
rect 26697 47511 26709 47545
rect 26743 47511 26755 47545
rect 26697 47477 26755 47511
rect 26697 47443 26709 47477
rect 26743 47443 26755 47477
rect 26697 47427 26755 47443
rect 27155 48701 27213 48717
rect 27155 48667 27167 48701
rect 27201 48667 27213 48701
rect 27155 48633 27213 48667
rect 27155 48599 27167 48633
rect 27201 48599 27213 48633
rect 27155 48565 27213 48599
rect 27155 48531 27167 48565
rect 27201 48531 27213 48565
rect 27155 48497 27213 48531
rect 27155 48463 27167 48497
rect 27201 48463 27213 48497
rect 27155 48429 27213 48463
rect 27155 48395 27167 48429
rect 27201 48395 27213 48429
rect 27155 48361 27213 48395
rect 27155 48327 27167 48361
rect 27201 48327 27213 48361
rect 27155 48293 27213 48327
rect 27155 48259 27167 48293
rect 27201 48259 27213 48293
rect 27155 48225 27213 48259
rect 27155 48191 27167 48225
rect 27201 48191 27213 48225
rect 27155 48157 27213 48191
rect 27155 48123 27167 48157
rect 27201 48123 27213 48157
rect 27155 48089 27213 48123
rect 27155 48055 27167 48089
rect 27201 48055 27213 48089
rect 27155 48021 27213 48055
rect 27155 47987 27167 48021
rect 27201 47987 27213 48021
rect 27155 47953 27213 47987
rect 27155 47919 27167 47953
rect 27201 47919 27213 47953
rect 27155 47885 27213 47919
rect 27155 47851 27167 47885
rect 27201 47851 27213 47885
rect 27155 47817 27213 47851
rect 27155 47783 27167 47817
rect 27201 47783 27213 47817
rect 27155 47749 27213 47783
rect 27155 47715 27167 47749
rect 27201 47715 27213 47749
rect 27155 47681 27213 47715
rect 27155 47647 27167 47681
rect 27201 47647 27213 47681
rect 27155 47613 27213 47647
rect 27155 47579 27167 47613
rect 27201 47579 27213 47613
rect 27155 47545 27213 47579
rect 27155 47511 27167 47545
rect 27201 47511 27213 47545
rect 27155 47477 27213 47511
rect 27155 47443 27167 47477
rect 27201 47443 27213 47477
rect 27155 47427 27213 47443
rect 27613 48701 27671 48717
rect 27613 48667 27625 48701
rect 27659 48667 27671 48701
rect 27613 48633 27671 48667
rect 27613 48599 27625 48633
rect 27659 48599 27671 48633
rect 27613 48565 27671 48599
rect 27613 48531 27625 48565
rect 27659 48531 27671 48565
rect 27613 48497 27671 48531
rect 27613 48463 27625 48497
rect 27659 48463 27671 48497
rect 27613 48429 27671 48463
rect 27613 48395 27625 48429
rect 27659 48395 27671 48429
rect 27613 48361 27671 48395
rect 27613 48327 27625 48361
rect 27659 48327 27671 48361
rect 27613 48293 27671 48327
rect 27613 48259 27625 48293
rect 27659 48259 27671 48293
rect 27613 48225 27671 48259
rect 27613 48191 27625 48225
rect 27659 48191 27671 48225
rect 27613 48157 27671 48191
rect 27613 48123 27625 48157
rect 27659 48123 27671 48157
rect 27613 48089 27671 48123
rect 27613 48055 27625 48089
rect 27659 48055 27671 48089
rect 27613 48021 27671 48055
rect 27613 47987 27625 48021
rect 27659 47987 27671 48021
rect 27613 47953 27671 47987
rect 27613 47919 27625 47953
rect 27659 47919 27671 47953
rect 27613 47885 27671 47919
rect 27613 47851 27625 47885
rect 27659 47851 27671 47885
rect 27613 47817 27671 47851
rect 27613 47783 27625 47817
rect 27659 47783 27671 47817
rect 27613 47749 27671 47783
rect 27613 47715 27625 47749
rect 27659 47715 27671 47749
rect 27613 47681 27671 47715
rect 27613 47647 27625 47681
rect 27659 47647 27671 47681
rect 27613 47613 27671 47647
rect 27613 47579 27625 47613
rect 27659 47579 27671 47613
rect 27613 47545 27671 47579
rect 27613 47511 27625 47545
rect 27659 47511 27671 47545
rect 27613 47477 27671 47511
rect 27613 47443 27625 47477
rect 27659 47443 27671 47477
rect 27613 47427 27671 47443
rect 28071 48701 28129 48717
rect 28071 48667 28083 48701
rect 28117 48667 28129 48701
rect 28071 48633 28129 48667
rect 28071 48599 28083 48633
rect 28117 48599 28129 48633
rect 28071 48565 28129 48599
rect 28071 48531 28083 48565
rect 28117 48531 28129 48565
rect 28071 48497 28129 48531
rect 28071 48463 28083 48497
rect 28117 48463 28129 48497
rect 28071 48429 28129 48463
rect 28071 48395 28083 48429
rect 28117 48395 28129 48429
rect 28071 48361 28129 48395
rect 28071 48327 28083 48361
rect 28117 48327 28129 48361
rect 28071 48293 28129 48327
rect 28071 48259 28083 48293
rect 28117 48259 28129 48293
rect 28071 48225 28129 48259
rect 28071 48191 28083 48225
rect 28117 48191 28129 48225
rect 28071 48157 28129 48191
rect 28071 48123 28083 48157
rect 28117 48123 28129 48157
rect 28071 48089 28129 48123
rect 28071 48055 28083 48089
rect 28117 48055 28129 48089
rect 28071 48021 28129 48055
rect 28071 47987 28083 48021
rect 28117 47987 28129 48021
rect 28071 47953 28129 47987
rect 28071 47919 28083 47953
rect 28117 47919 28129 47953
rect 28071 47885 28129 47919
rect 28071 47851 28083 47885
rect 28117 47851 28129 47885
rect 28071 47817 28129 47851
rect 28071 47783 28083 47817
rect 28117 47783 28129 47817
rect 28071 47749 28129 47783
rect 28071 47715 28083 47749
rect 28117 47715 28129 47749
rect 28071 47681 28129 47715
rect 28071 47647 28083 47681
rect 28117 47647 28129 47681
rect 28071 47613 28129 47647
rect 28071 47579 28083 47613
rect 28117 47579 28129 47613
rect 28071 47545 28129 47579
rect 28071 47511 28083 47545
rect 28117 47511 28129 47545
rect 28071 47477 28129 47511
rect 28071 47443 28083 47477
rect 28117 47443 28129 47477
rect 28071 47427 28129 47443
rect 28529 48701 28587 48717
rect 28529 48667 28541 48701
rect 28575 48667 28587 48701
rect 28529 48633 28587 48667
rect 28529 48599 28541 48633
rect 28575 48599 28587 48633
rect 28529 48565 28587 48599
rect 28529 48531 28541 48565
rect 28575 48531 28587 48565
rect 28529 48497 28587 48531
rect 28529 48463 28541 48497
rect 28575 48463 28587 48497
rect 28529 48429 28587 48463
rect 28529 48395 28541 48429
rect 28575 48395 28587 48429
rect 28529 48361 28587 48395
rect 28529 48327 28541 48361
rect 28575 48327 28587 48361
rect 28529 48293 28587 48327
rect 28529 48259 28541 48293
rect 28575 48259 28587 48293
rect 28529 48225 28587 48259
rect 28529 48191 28541 48225
rect 28575 48191 28587 48225
rect 28529 48157 28587 48191
rect 28529 48123 28541 48157
rect 28575 48123 28587 48157
rect 28529 48089 28587 48123
rect 28529 48055 28541 48089
rect 28575 48055 28587 48089
rect 28529 48021 28587 48055
rect 28529 47987 28541 48021
rect 28575 47987 28587 48021
rect 28529 47953 28587 47987
rect 28529 47919 28541 47953
rect 28575 47919 28587 47953
rect 28529 47885 28587 47919
rect 28529 47851 28541 47885
rect 28575 47851 28587 47885
rect 28529 47817 28587 47851
rect 28529 47783 28541 47817
rect 28575 47783 28587 47817
rect 28529 47749 28587 47783
rect 28529 47715 28541 47749
rect 28575 47715 28587 47749
rect 28529 47681 28587 47715
rect 28529 47647 28541 47681
rect 28575 47647 28587 47681
rect 28529 47613 28587 47647
rect 28529 47579 28541 47613
rect 28575 47579 28587 47613
rect 28529 47545 28587 47579
rect 28529 47511 28541 47545
rect 28575 47511 28587 47545
rect 28529 47477 28587 47511
rect 28529 47443 28541 47477
rect 28575 47443 28587 47477
rect 28529 47427 28587 47443
rect 28987 48701 29045 48717
rect 28987 48667 28999 48701
rect 29033 48667 29045 48701
rect 28987 48633 29045 48667
rect 28987 48599 28999 48633
rect 29033 48599 29045 48633
rect 28987 48565 29045 48599
rect 28987 48531 28999 48565
rect 29033 48531 29045 48565
rect 28987 48497 29045 48531
rect 28987 48463 28999 48497
rect 29033 48463 29045 48497
rect 28987 48429 29045 48463
rect 28987 48395 28999 48429
rect 29033 48395 29045 48429
rect 28987 48361 29045 48395
rect 28987 48327 28999 48361
rect 29033 48327 29045 48361
rect 28987 48293 29045 48327
rect 28987 48259 28999 48293
rect 29033 48259 29045 48293
rect 28987 48225 29045 48259
rect 28987 48191 28999 48225
rect 29033 48191 29045 48225
rect 28987 48157 29045 48191
rect 28987 48123 28999 48157
rect 29033 48123 29045 48157
rect 28987 48089 29045 48123
rect 28987 48055 28999 48089
rect 29033 48055 29045 48089
rect 28987 48021 29045 48055
rect 28987 47987 28999 48021
rect 29033 47987 29045 48021
rect 28987 47953 29045 47987
rect 28987 47919 28999 47953
rect 29033 47919 29045 47953
rect 28987 47885 29045 47919
rect 28987 47851 28999 47885
rect 29033 47851 29045 47885
rect 28987 47817 29045 47851
rect 28987 47783 28999 47817
rect 29033 47783 29045 47817
rect 28987 47749 29045 47783
rect 28987 47715 28999 47749
rect 29033 47715 29045 47749
rect 28987 47681 29045 47715
rect 28987 47647 28999 47681
rect 29033 47647 29045 47681
rect 28987 47613 29045 47647
rect 28987 47579 28999 47613
rect 29033 47579 29045 47613
rect 28987 47545 29045 47579
rect 28987 47511 28999 47545
rect 29033 47511 29045 47545
rect 28987 47477 29045 47511
rect 28987 47443 28999 47477
rect 29033 47443 29045 47477
rect 28987 47427 29045 47443
rect 29445 48701 29503 48717
rect 29445 48667 29457 48701
rect 29491 48667 29503 48701
rect 29445 48633 29503 48667
rect 29445 48599 29457 48633
rect 29491 48599 29503 48633
rect 29445 48565 29503 48599
rect 29445 48531 29457 48565
rect 29491 48531 29503 48565
rect 29445 48497 29503 48531
rect 29445 48463 29457 48497
rect 29491 48463 29503 48497
rect 29445 48429 29503 48463
rect 29445 48395 29457 48429
rect 29491 48395 29503 48429
rect 29445 48361 29503 48395
rect 29445 48327 29457 48361
rect 29491 48327 29503 48361
rect 29445 48293 29503 48327
rect 29445 48259 29457 48293
rect 29491 48259 29503 48293
rect 29445 48225 29503 48259
rect 29445 48191 29457 48225
rect 29491 48191 29503 48225
rect 29445 48157 29503 48191
rect 29445 48123 29457 48157
rect 29491 48123 29503 48157
rect 29445 48089 29503 48123
rect 29445 48055 29457 48089
rect 29491 48055 29503 48089
rect 29445 48021 29503 48055
rect 29445 47987 29457 48021
rect 29491 47987 29503 48021
rect 29445 47953 29503 47987
rect 29445 47919 29457 47953
rect 29491 47919 29503 47953
rect 29445 47885 29503 47919
rect 29445 47851 29457 47885
rect 29491 47851 29503 47885
rect 29445 47817 29503 47851
rect 29445 47783 29457 47817
rect 29491 47783 29503 47817
rect 29445 47749 29503 47783
rect 29445 47715 29457 47749
rect 29491 47715 29503 47749
rect 29445 47681 29503 47715
rect 29445 47647 29457 47681
rect 29491 47647 29503 47681
rect 29445 47613 29503 47647
rect 29445 47579 29457 47613
rect 29491 47579 29503 47613
rect 29445 47545 29503 47579
rect 29445 47511 29457 47545
rect 29491 47511 29503 47545
rect 29445 47477 29503 47511
rect 29445 47443 29457 47477
rect 29491 47443 29503 47477
rect 29445 47427 29503 47443
rect 29903 48701 29961 48717
rect 29903 48667 29915 48701
rect 29949 48667 29961 48701
rect 29903 48633 29961 48667
rect 29903 48599 29915 48633
rect 29949 48599 29961 48633
rect 29903 48565 29961 48599
rect 29903 48531 29915 48565
rect 29949 48531 29961 48565
rect 29903 48497 29961 48531
rect 29903 48463 29915 48497
rect 29949 48463 29961 48497
rect 29903 48429 29961 48463
rect 29903 48395 29915 48429
rect 29949 48395 29961 48429
rect 29903 48361 29961 48395
rect 29903 48327 29915 48361
rect 29949 48327 29961 48361
rect 29903 48293 29961 48327
rect 29903 48259 29915 48293
rect 29949 48259 29961 48293
rect 29903 48225 29961 48259
rect 29903 48191 29915 48225
rect 29949 48191 29961 48225
rect 29903 48157 29961 48191
rect 29903 48123 29915 48157
rect 29949 48123 29961 48157
rect 29903 48089 29961 48123
rect 29903 48055 29915 48089
rect 29949 48055 29961 48089
rect 29903 48021 29961 48055
rect 29903 47987 29915 48021
rect 29949 47987 29961 48021
rect 29903 47953 29961 47987
rect 29903 47919 29915 47953
rect 29949 47919 29961 47953
rect 29903 47885 29961 47919
rect 29903 47851 29915 47885
rect 29949 47851 29961 47885
rect 29903 47817 29961 47851
rect 29903 47783 29915 47817
rect 29949 47783 29961 47817
rect 29903 47749 29961 47783
rect 29903 47715 29915 47749
rect 29949 47715 29961 47749
rect 29903 47681 29961 47715
rect 29903 47647 29915 47681
rect 29949 47647 29961 47681
rect 29903 47613 29961 47647
rect 29903 47579 29915 47613
rect 29949 47579 29961 47613
rect 29903 47545 29961 47579
rect 29903 47511 29915 47545
rect 29949 47511 29961 47545
rect 29903 47477 29961 47511
rect 29903 47443 29915 47477
rect 29949 47443 29961 47477
rect 29903 47427 29961 47443
rect 30361 48701 30419 48717
rect 30361 48667 30373 48701
rect 30407 48667 30419 48701
rect 30361 48633 30419 48667
rect 30361 48599 30373 48633
rect 30407 48599 30419 48633
rect 30361 48565 30419 48599
rect 30361 48531 30373 48565
rect 30407 48531 30419 48565
rect 30361 48497 30419 48531
rect 30361 48463 30373 48497
rect 30407 48463 30419 48497
rect 30361 48429 30419 48463
rect 30361 48395 30373 48429
rect 30407 48395 30419 48429
rect 30361 48361 30419 48395
rect 30361 48327 30373 48361
rect 30407 48327 30419 48361
rect 30361 48293 30419 48327
rect 30361 48259 30373 48293
rect 30407 48259 30419 48293
rect 30361 48225 30419 48259
rect 30361 48191 30373 48225
rect 30407 48191 30419 48225
rect 30361 48157 30419 48191
rect 30361 48123 30373 48157
rect 30407 48123 30419 48157
rect 30361 48089 30419 48123
rect 30361 48055 30373 48089
rect 30407 48055 30419 48089
rect 30361 48021 30419 48055
rect 30361 47987 30373 48021
rect 30407 47987 30419 48021
rect 30361 47953 30419 47987
rect 30361 47919 30373 47953
rect 30407 47919 30419 47953
rect 30361 47885 30419 47919
rect 30361 47851 30373 47885
rect 30407 47851 30419 47885
rect 30361 47817 30419 47851
rect 30361 47783 30373 47817
rect 30407 47783 30419 47817
rect 30361 47749 30419 47783
rect 30361 47715 30373 47749
rect 30407 47715 30419 47749
rect 30361 47681 30419 47715
rect 30361 47647 30373 47681
rect 30407 47647 30419 47681
rect 30361 47613 30419 47647
rect 30361 47579 30373 47613
rect 30407 47579 30419 47613
rect 30361 47545 30419 47579
rect 30361 47511 30373 47545
rect 30407 47511 30419 47545
rect 30361 47477 30419 47511
rect 30361 47443 30373 47477
rect 30407 47443 30419 47477
rect 30361 47427 30419 47443
rect 30819 48701 30877 48717
rect 30819 48667 30831 48701
rect 30865 48667 30877 48701
rect 30819 48633 30877 48667
rect 30819 48599 30831 48633
rect 30865 48599 30877 48633
rect 30819 48565 30877 48599
rect 30819 48531 30831 48565
rect 30865 48531 30877 48565
rect 30819 48497 30877 48531
rect 30819 48463 30831 48497
rect 30865 48463 30877 48497
rect 30819 48429 30877 48463
rect 30819 48395 30831 48429
rect 30865 48395 30877 48429
rect 30819 48361 30877 48395
rect 30819 48327 30831 48361
rect 30865 48327 30877 48361
rect 30819 48293 30877 48327
rect 30819 48259 30831 48293
rect 30865 48259 30877 48293
rect 30819 48225 30877 48259
rect 30819 48191 30831 48225
rect 30865 48191 30877 48225
rect 30819 48157 30877 48191
rect 30819 48123 30831 48157
rect 30865 48123 30877 48157
rect 30819 48089 30877 48123
rect 30819 48055 30831 48089
rect 30865 48055 30877 48089
rect 30819 48021 30877 48055
rect 30819 47987 30831 48021
rect 30865 47987 30877 48021
rect 30819 47953 30877 47987
rect 30819 47919 30831 47953
rect 30865 47919 30877 47953
rect 30819 47885 30877 47919
rect 30819 47851 30831 47885
rect 30865 47851 30877 47885
rect 30819 47817 30877 47851
rect 30819 47783 30831 47817
rect 30865 47783 30877 47817
rect 30819 47749 30877 47783
rect 30819 47715 30831 47749
rect 30865 47715 30877 47749
rect 30819 47681 30877 47715
rect 30819 47647 30831 47681
rect 30865 47647 30877 47681
rect 30819 47613 30877 47647
rect 30819 47579 30831 47613
rect 30865 47579 30877 47613
rect 30819 47545 30877 47579
rect 30819 47511 30831 47545
rect 30865 47511 30877 47545
rect 30819 47477 30877 47511
rect 30819 47443 30831 47477
rect 30865 47443 30877 47477
rect 30819 47427 30877 47443
rect 31277 48701 31335 48717
rect 31277 48667 31289 48701
rect 31323 48667 31335 48701
rect 31277 48633 31335 48667
rect 31277 48599 31289 48633
rect 31323 48599 31335 48633
rect 31277 48565 31335 48599
rect 31277 48531 31289 48565
rect 31323 48531 31335 48565
rect 31277 48497 31335 48531
rect 31277 48463 31289 48497
rect 31323 48463 31335 48497
rect 31277 48429 31335 48463
rect 31277 48395 31289 48429
rect 31323 48395 31335 48429
rect 31277 48361 31335 48395
rect 31277 48327 31289 48361
rect 31323 48327 31335 48361
rect 31277 48293 31335 48327
rect 31277 48259 31289 48293
rect 31323 48259 31335 48293
rect 31277 48225 31335 48259
rect 31277 48191 31289 48225
rect 31323 48191 31335 48225
rect 31277 48157 31335 48191
rect 31277 48123 31289 48157
rect 31323 48123 31335 48157
rect 31277 48089 31335 48123
rect 31277 48055 31289 48089
rect 31323 48055 31335 48089
rect 31277 48021 31335 48055
rect 31277 47987 31289 48021
rect 31323 47987 31335 48021
rect 31277 47953 31335 47987
rect 31277 47919 31289 47953
rect 31323 47919 31335 47953
rect 31277 47885 31335 47919
rect 31277 47851 31289 47885
rect 31323 47851 31335 47885
rect 31277 47817 31335 47851
rect 31277 47783 31289 47817
rect 31323 47783 31335 47817
rect 31277 47749 31335 47783
rect 31277 47715 31289 47749
rect 31323 47715 31335 47749
rect 31277 47681 31335 47715
rect 31277 47647 31289 47681
rect 31323 47647 31335 47681
rect 31277 47613 31335 47647
rect 31277 47579 31289 47613
rect 31323 47579 31335 47613
rect 31277 47545 31335 47579
rect 31277 47511 31289 47545
rect 31323 47511 31335 47545
rect 31277 47477 31335 47511
rect 31277 47443 31289 47477
rect 31323 47443 31335 47477
rect 31277 47427 31335 47443
rect 31735 48701 31793 48717
rect 31735 48667 31747 48701
rect 31781 48667 31793 48701
rect 31735 48633 31793 48667
rect 31735 48599 31747 48633
rect 31781 48599 31793 48633
rect 31735 48565 31793 48599
rect 31735 48531 31747 48565
rect 31781 48531 31793 48565
rect 31735 48497 31793 48531
rect 31735 48463 31747 48497
rect 31781 48463 31793 48497
rect 31735 48429 31793 48463
rect 31735 48395 31747 48429
rect 31781 48395 31793 48429
rect 31735 48361 31793 48395
rect 31735 48327 31747 48361
rect 31781 48327 31793 48361
rect 31735 48293 31793 48327
rect 31735 48259 31747 48293
rect 31781 48259 31793 48293
rect 31735 48225 31793 48259
rect 31735 48191 31747 48225
rect 31781 48191 31793 48225
rect 31735 48157 31793 48191
rect 31735 48123 31747 48157
rect 31781 48123 31793 48157
rect 31735 48089 31793 48123
rect 31735 48055 31747 48089
rect 31781 48055 31793 48089
rect 31735 48021 31793 48055
rect 31735 47987 31747 48021
rect 31781 47987 31793 48021
rect 31735 47953 31793 47987
rect 31735 47919 31747 47953
rect 31781 47919 31793 47953
rect 31735 47885 31793 47919
rect 31735 47851 31747 47885
rect 31781 47851 31793 47885
rect 31735 47817 31793 47851
rect 31735 47783 31747 47817
rect 31781 47783 31793 47817
rect 31735 47749 31793 47783
rect 31735 47715 31747 47749
rect 31781 47715 31793 47749
rect 31735 47681 31793 47715
rect 31735 47647 31747 47681
rect 31781 47647 31793 47681
rect 31735 47613 31793 47647
rect 31735 47579 31747 47613
rect 31781 47579 31793 47613
rect 31735 47545 31793 47579
rect 31735 47511 31747 47545
rect 31781 47511 31793 47545
rect 31735 47477 31793 47511
rect 31735 47443 31747 47477
rect 31781 47443 31793 47477
rect 31735 47427 31793 47443
rect 32193 48701 32251 48717
rect 32193 48667 32205 48701
rect 32239 48667 32251 48701
rect 32193 48633 32251 48667
rect 32193 48599 32205 48633
rect 32239 48599 32251 48633
rect 32193 48565 32251 48599
rect 32193 48531 32205 48565
rect 32239 48531 32251 48565
rect 32193 48497 32251 48531
rect 32193 48463 32205 48497
rect 32239 48463 32251 48497
rect 32193 48429 32251 48463
rect 32193 48395 32205 48429
rect 32239 48395 32251 48429
rect 32193 48361 32251 48395
rect 32193 48327 32205 48361
rect 32239 48327 32251 48361
rect 32193 48293 32251 48327
rect 32193 48259 32205 48293
rect 32239 48259 32251 48293
rect 32193 48225 32251 48259
rect 32193 48191 32205 48225
rect 32239 48191 32251 48225
rect 32193 48157 32251 48191
rect 32193 48123 32205 48157
rect 32239 48123 32251 48157
rect 32193 48089 32251 48123
rect 32193 48055 32205 48089
rect 32239 48055 32251 48089
rect 32193 48021 32251 48055
rect 32193 47987 32205 48021
rect 32239 47987 32251 48021
rect 32193 47953 32251 47987
rect 32193 47919 32205 47953
rect 32239 47919 32251 47953
rect 32193 47885 32251 47919
rect 32193 47851 32205 47885
rect 32239 47851 32251 47885
rect 32193 47817 32251 47851
rect 32193 47783 32205 47817
rect 32239 47783 32251 47817
rect 32193 47749 32251 47783
rect 32193 47715 32205 47749
rect 32239 47715 32251 47749
rect 32193 47681 32251 47715
rect 32193 47647 32205 47681
rect 32239 47647 32251 47681
rect 32193 47613 32251 47647
rect 32193 47579 32205 47613
rect 32239 47579 32251 47613
rect 32193 47545 32251 47579
rect 32193 47511 32205 47545
rect 32239 47511 32251 47545
rect 32193 47477 32251 47511
rect 32193 47443 32205 47477
rect 32239 47443 32251 47477
rect 32193 47427 32251 47443
rect 32651 48701 32709 48717
rect 32651 48667 32663 48701
rect 32697 48667 32709 48701
rect 32651 48633 32709 48667
rect 32651 48599 32663 48633
rect 32697 48599 32709 48633
rect 32651 48565 32709 48599
rect 32651 48531 32663 48565
rect 32697 48531 32709 48565
rect 32651 48497 32709 48531
rect 32651 48463 32663 48497
rect 32697 48463 32709 48497
rect 32651 48429 32709 48463
rect 32651 48395 32663 48429
rect 32697 48395 32709 48429
rect 32651 48361 32709 48395
rect 32651 48327 32663 48361
rect 32697 48327 32709 48361
rect 32651 48293 32709 48327
rect 32651 48259 32663 48293
rect 32697 48259 32709 48293
rect 32651 48225 32709 48259
rect 32651 48191 32663 48225
rect 32697 48191 32709 48225
rect 32651 48157 32709 48191
rect 32651 48123 32663 48157
rect 32697 48123 32709 48157
rect 32651 48089 32709 48123
rect 32651 48055 32663 48089
rect 32697 48055 32709 48089
rect 32651 48021 32709 48055
rect 32651 47987 32663 48021
rect 32697 47987 32709 48021
rect 32651 47953 32709 47987
rect 32651 47919 32663 47953
rect 32697 47919 32709 47953
rect 32651 47885 32709 47919
rect 32651 47851 32663 47885
rect 32697 47851 32709 47885
rect 32651 47817 32709 47851
rect 32651 47783 32663 47817
rect 32697 47783 32709 47817
rect 32651 47749 32709 47783
rect 32651 47715 32663 47749
rect 32697 47715 32709 47749
rect 32651 47681 32709 47715
rect 32651 47647 32663 47681
rect 32697 47647 32709 47681
rect 32651 47613 32709 47647
rect 32651 47579 32663 47613
rect 32697 47579 32709 47613
rect 32651 47545 32709 47579
rect 32651 47511 32663 47545
rect 32697 47511 32709 47545
rect 32651 47477 32709 47511
rect 32651 47443 32663 47477
rect 32697 47443 32709 47477
rect 32651 47427 32709 47443
rect 33109 48701 33167 48717
rect 33109 48667 33121 48701
rect 33155 48667 33167 48701
rect 33109 48633 33167 48667
rect 33109 48599 33121 48633
rect 33155 48599 33167 48633
rect 33109 48565 33167 48599
rect 33109 48531 33121 48565
rect 33155 48531 33167 48565
rect 33109 48497 33167 48531
rect 33109 48463 33121 48497
rect 33155 48463 33167 48497
rect 33109 48429 33167 48463
rect 33109 48395 33121 48429
rect 33155 48395 33167 48429
rect 33109 48361 33167 48395
rect 33109 48327 33121 48361
rect 33155 48327 33167 48361
rect 33109 48293 33167 48327
rect 33109 48259 33121 48293
rect 33155 48259 33167 48293
rect 33109 48225 33167 48259
rect 33109 48191 33121 48225
rect 33155 48191 33167 48225
rect 33109 48157 33167 48191
rect 33109 48123 33121 48157
rect 33155 48123 33167 48157
rect 33109 48089 33167 48123
rect 33109 48055 33121 48089
rect 33155 48055 33167 48089
rect 33109 48021 33167 48055
rect 33109 47987 33121 48021
rect 33155 47987 33167 48021
rect 33109 47953 33167 47987
rect 33109 47919 33121 47953
rect 33155 47919 33167 47953
rect 33109 47885 33167 47919
rect 33109 47851 33121 47885
rect 33155 47851 33167 47885
rect 33109 47817 33167 47851
rect 33109 47783 33121 47817
rect 33155 47783 33167 47817
rect 33109 47749 33167 47783
rect 33109 47715 33121 47749
rect 33155 47715 33167 47749
rect 33109 47681 33167 47715
rect 33109 47647 33121 47681
rect 33155 47647 33167 47681
rect 33109 47613 33167 47647
rect 33109 47579 33121 47613
rect 33155 47579 33167 47613
rect 33109 47545 33167 47579
rect 33109 47511 33121 47545
rect 33155 47511 33167 47545
rect 33109 47477 33167 47511
rect 33109 47443 33121 47477
rect 33155 47443 33167 47477
rect 33109 47427 33167 47443
rect 33567 48701 33625 48717
rect 33567 48667 33579 48701
rect 33613 48667 33625 48701
rect 33567 48633 33625 48667
rect 33567 48599 33579 48633
rect 33613 48599 33625 48633
rect 33567 48565 33625 48599
rect 33567 48531 33579 48565
rect 33613 48531 33625 48565
rect 33567 48497 33625 48531
rect 33567 48463 33579 48497
rect 33613 48463 33625 48497
rect 33567 48429 33625 48463
rect 33567 48395 33579 48429
rect 33613 48395 33625 48429
rect 33567 48361 33625 48395
rect 33567 48327 33579 48361
rect 33613 48327 33625 48361
rect 33567 48293 33625 48327
rect 33567 48259 33579 48293
rect 33613 48259 33625 48293
rect 33567 48225 33625 48259
rect 33567 48191 33579 48225
rect 33613 48191 33625 48225
rect 33567 48157 33625 48191
rect 33567 48123 33579 48157
rect 33613 48123 33625 48157
rect 33567 48089 33625 48123
rect 33567 48055 33579 48089
rect 33613 48055 33625 48089
rect 33567 48021 33625 48055
rect 33567 47987 33579 48021
rect 33613 47987 33625 48021
rect 33567 47953 33625 47987
rect 33567 47919 33579 47953
rect 33613 47919 33625 47953
rect 33567 47885 33625 47919
rect 33567 47851 33579 47885
rect 33613 47851 33625 47885
rect 33567 47817 33625 47851
rect 33567 47783 33579 47817
rect 33613 47783 33625 47817
rect 33567 47749 33625 47783
rect 33567 47715 33579 47749
rect 33613 47715 33625 47749
rect 33567 47681 33625 47715
rect 33567 47647 33579 47681
rect 33613 47647 33625 47681
rect 33567 47613 33625 47647
rect 33567 47579 33579 47613
rect 33613 47579 33625 47613
rect 33567 47545 33625 47579
rect 33567 47511 33579 47545
rect 33613 47511 33625 47545
rect 33567 47477 33625 47511
rect 33567 47443 33579 47477
rect 33613 47443 33625 47477
rect 33567 47427 33625 47443
rect 34025 48701 34083 48717
rect 34025 48667 34037 48701
rect 34071 48667 34083 48701
rect 34025 48633 34083 48667
rect 34025 48599 34037 48633
rect 34071 48599 34083 48633
rect 34025 48565 34083 48599
rect 34025 48531 34037 48565
rect 34071 48531 34083 48565
rect 34025 48497 34083 48531
rect 34025 48463 34037 48497
rect 34071 48463 34083 48497
rect 34025 48429 34083 48463
rect 34025 48395 34037 48429
rect 34071 48395 34083 48429
rect 34025 48361 34083 48395
rect 34025 48327 34037 48361
rect 34071 48327 34083 48361
rect 34025 48293 34083 48327
rect 34025 48259 34037 48293
rect 34071 48259 34083 48293
rect 34025 48225 34083 48259
rect 34025 48191 34037 48225
rect 34071 48191 34083 48225
rect 34025 48157 34083 48191
rect 34025 48123 34037 48157
rect 34071 48123 34083 48157
rect 34025 48089 34083 48123
rect 34025 48055 34037 48089
rect 34071 48055 34083 48089
rect 34025 48021 34083 48055
rect 34025 47987 34037 48021
rect 34071 47987 34083 48021
rect 34025 47953 34083 47987
rect 34025 47919 34037 47953
rect 34071 47919 34083 47953
rect 34025 47885 34083 47919
rect 34025 47851 34037 47885
rect 34071 47851 34083 47885
rect 34025 47817 34083 47851
rect 34025 47783 34037 47817
rect 34071 47783 34083 47817
rect 34025 47749 34083 47783
rect 34025 47715 34037 47749
rect 34071 47715 34083 47749
rect 34025 47681 34083 47715
rect 34025 47647 34037 47681
rect 34071 47647 34083 47681
rect 34025 47613 34083 47647
rect 34025 47579 34037 47613
rect 34071 47579 34083 47613
rect 34025 47545 34083 47579
rect 34025 47511 34037 47545
rect 34071 47511 34083 47545
rect 34025 47477 34083 47511
rect 34025 47443 34037 47477
rect 34071 47443 34083 47477
rect 34025 47427 34083 47443
rect 34483 48701 34541 48717
rect 34483 48667 34495 48701
rect 34529 48667 34541 48701
rect 34483 48633 34541 48667
rect 34483 48599 34495 48633
rect 34529 48599 34541 48633
rect 34483 48565 34541 48599
rect 34483 48531 34495 48565
rect 34529 48531 34541 48565
rect 34483 48497 34541 48531
rect 34483 48463 34495 48497
rect 34529 48463 34541 48497
rect 34483 48429 34541 48463
rect 34483 48395 34495 48429
rect 34529 48395 34541 48429
rect 34483 48361 34541 48395
rect 34483 48327 34495 48361
rect 34529 48327 34541 48361
rect 34483 48293 34541 48327
rect 34483 48259 34495 48293
rect 34529 48259 34541 48293
rect 34483 48225 34541 48259
rect 34483 48191 34495 48225
rect 34529 48191 34541 48225
rect 34483 48157 34541 48191
rect 34483 48123 34495 48157
rect 34529 48123 34541 48157
rect 34483 48089 34541 48123
rect 34483 48055 34495 48089
rect 34529 48055 34541 48089
rect 34483 48021 34541 48055
rect 34483 47987 34495 48021
rect 34529 47987 34541 48021
rect 34483 47953 34541 47987
rect 34483 47919 34495 47953
rect 34529 47919 34541 47953
rect 34483 47885 34541 47919
rect 34483 47851 34495 47885
rect 34529 47851 34541 47885
rect 34483 47817 34541 47851
rect 34483 47783 34495 47817
rect 34529 47783 34541 47817
rect 34483 47749 34541 47783
rect 34483 47715 34495 47749
rect 34529 47715 34541 47749
rect 34483 47681 34541 47715
rect 34483 47647 34495 47681
rect 34529 47647 34541 47681
rect 34483 47613 34541 47647
rect 34483 47579 34495 47613
rect 34529 47579 34541 47613
rect 34483 47545 34541 47579
rect 34483 47511 34495 47545
rect 34529 47511 34541 47545
rect 34483 47477 34541 47511
rect 34483 47443 34495 47477
rect 34529 47443 34541 47477
rect 34483 47427 34541 47443
rect 34941 48701 34999 48717
rect 34941 48667 34953 48701
rect 34987 48667 34999 48701
rect 34941 48633 34999 48667
rect 34941 48599 34953 48633
rect 34987 48599 34999 48633
rect 34941 48565 34999 48599
rect 34941 48531 34953 48565
rect 34987 48531 34999 48565
rect 34941 48497 34999 48531
rect 34941 48463 34953 48497
rect 34987 48463 34999 48497
rect 34941 48429 34999 48463
rect 34941 48395 34953 48429
rect 34987 48395 34999 48429
rect 34941 48361 34999 48395
rect 34941 48327 34953 48361
rect 34987 48327 34999 48361
rect 34941 48293 34999 48327
rect 34941 48259 34953 48293
rect 34987 48259 34999 48293
rect 34941 48225 34999 48259
rect 34941 48191 34953 48225
rect 34987 48191 34999 48225
rect 34941 48157 34999 48191
rect 34941 48123 34953 48157
rect 34987 48123 34999 48157
rect 34941 48089 34999 48123
rect 34941 48055 34953 48089
rect 34987 48055 34999 48089
rect 34941 48021 34999 48055
rect 34941 47987 34953 48021
rect 34987 47987 34999 48021
rect 34941 47953 34999 47987
rect 34941 47919 34953 47953
rect 34987 47919 34999 47953
rect 34941 47885 34999 47919
rect 34941 47851 34953 47885
rect 34987 47851 34999 47885
rect 34941 47817 34999 47851
rect 34941 47783 34953 47817
rect 34987 47783 34999 47817
rect 34941 47749 34999 47783
rect 34941 47715 34953 47749
rect 34987 47715 34999 47749
rect 34941 47681 34999 47715
rect 34941 47647 34953 47681
rect 34987 47647 34999 47681
rect 34941 47613 34999 47647
rect 34941 47579 34953 47613
rect 34987 47579 34999 47613
rect 34941 47545 34999 47579
rect 34941 47511 34953 47545
rect 34987 47511 34999 47545
rect 34941 47477 34999 47511
rect 34941 47443 34953 47477
rect 34987 47443 34999 47477
rect 34941 47427 34999 47443
rect 35399 48701 35457 48717
rect 35399 48667 35411 48701
rect 35445 48667 35457 48701
rect 35399 48633 35457 48667
rect 35399 48599 35411 48633
rect 35445 48599 35457 48633
rect 35399 48565 35457 48599
rect 35399 48531 35411 48565
rect 35445 48531 35457 48565
rect 35399 48497 35457 48531
rect 35399 48463 35411 48497
rect 35445 48463 35457 48497
rect 35399 48429 35457 48463
rect 35399 48395 35411 48429
rect 35445 48395 35457 48429
rect 35399 48361 35457 48395
rect 35399 48327 35411 48361
rect 35445 48327 35457 48361
rect 35399 48293 35457 48327
rect 35399 48259 35411 48293
rect 35445 48259 35457 48293
rect 35399 48225 35457 48259
rect 35399 48191 35411 48225
rect 35445 48191 35457 48225
rect 35399 48157 35457 48191
rect 35399 48123 35411 48157
rect 35445 48123 35457 48157
rect 35399 48089 35457 48123
rect 35399 48055 35411 48089
rect 35445 48055 35457 48089
rect 35399 48021 35457 48055
rect 35399 47987 35411 48021
rect 35445 47987 35457 48021
rect 35399 47953 35457 47987
rect 35399 47919 35411 47953
rect 35445 47919 35457 47953
rect 35399 47885 35457 47919
rect 35399 47851 35411 47885
rect 35445 47851 35457 47885
rect 35399 47817 35457 47851
rect 35399 47783 35411 47817
rect 35445 47783 35457 47817
rect 35399 47749 35457 47783
rect 35399 47715 35411 47749
rect 35445 47715 35457 47749
rect 35399 47681 35457 47715
rect 35399 47647 35411 47681
rect 35445 47647 35457 47681
rect 35399 47613 35457 47647
rect 35399 47579 35411 47613
rect 35445 47579 35457 47613
rect 35399 47545 35457 47579
rect 35399 47511 35411 47545
rect 35445 47511 35457 47545
rect 35399 47477 35457 47511
rect 35399 47443 35411 47477
rect 35445 47443 35457 47477
rect 35399 47427 35457 47443
rect 35857 48701 35915 48717
rect 35857 48667 35869 48701
rect 35903 48667 35915 48701
rect 35857 48633 35915 48667
rect 35857 48599 35869 48633
rect 35903 48599 35915 48633
rect 35857 48565 35915 48599
rect 35857 48531 35869 48565
rect 35903 48531 35915 48565
rect 35857 48497 35915 48531
rect 35857 48463 35869 48497
rect 35903 48463 35915 48497
rect 35857 48429 35915 48463
rect 35857 48395 35869 48429
rect 35903 48395 35915 48429
rect 35857 48361 35915 48395
rect 35857 48327 35869 48361
rect 35903 48327 35915 48361
rect 35857 48293 35915 48327
rect 35857 48259 35869 48293
rect 35903 48259 35915 48293
rect 35857 48225 35915 48259
rect 35857 48191 35869 48225
rect 35903 48191 35915 48225
rect 35857 48157 35915 48191
rect 35857 48123 35869 48157
rect 35903 48123 35915 48157
rect 35857 48089 35915 48123
rect 35857 48055 35869 48089
rect 35903 48055 35915 48089
rect 35857 48021 35915 48055
rect 35857 47987 35869 48021
rect 35903 47987 35915 48021
rect 35857 47953 35915 47987
rect 35857 47919 35869 47953
rect 35903 47919 35915 47953
rect 35857 47885 35915 47919
rect 35857 47851 35869 47885
rect 35903 47851 35915 47885
rect 35857 47817 35915 47851
rect 35857 47783 35869 47817
rect 35903 47783 35915 47817
rect 35857 47749 35915 47783
rect 35857 47715 35869 47749
rect 35903 47715 35915 47749
rect 35857 47681 35915 47715
rect 35857 47647 35869 47681
rect 35903 47647 35915 47681
rect 35857 47613 35915 47647
rect 35857 47579 35869 47613
rect 35903 47579 35915 47613
rect 35857 47545 35915 47579
rect 35857 47511 35869 47545
rect 35903 47511 35915 47545
rect 35857 47477 35915 47511
rect 35857 47443 35869 47477
rect 35903 47443 35915 47477
rect 35857 47427 35915 47443
rect 36315 48701 36373 48717
rect 36315 48667 36327 48701
rect 36361 48667 36373 48701
rect 36315 48633 36373 48667
rect 36315 48599 36327 48633
rect 36361 48599 36373 48633
rect 36315 48565 36373 48599
rect 36315 48531 36327 48565
rect 36361 48531 36373 48565
rect 36315 48497 36373 48531
rect 36315 48463 36327 48497
rect 36361 48463 36373 48497
rect 36315 48429 36373 48463
rect 36315 48395 36327 48429
rect 36361 48395 36373 48429
rect 36315 48361 36373 48395
rect 36315 48327 36327 48361
rect 36361 48327 36373 48361
rect 36315 48293 36373 48327
rect 36315 48259 36327 48293
rect 36361 48259 36373 48293
rect 36315 48225 36373 48259
rect 36315 48191 36327 48225
rect 36361 48191 36373 48225
rect 36315 48157 36373 48191
rect 36315 48123 36327 48157
rect 36361 48123 36373 48157
rect 36315 48089 36373 48123
rect 36315 48055 36327 48089
rect 36361 48055 36373 48089
rect 36315 48021 36373 48055
rect 36315 47987 36327 48021
rect 36361 47987 36373 48021
rect 36315 47953 36373 47987
rect 36315 47919 36327 47953
rect 36361 47919 36373 47953
rect 36315 47885 36373 47919
rect 36315 47851 36327 47885
rect 36361 47851 36373 47885
rect 36315 47817 36373 47851
rect 36315 47783 36327 47817
rect 36361 47783 36373 47817
rect 36315 47749 36373 47783
rect 36315 47715 36327 47749
rect 36361 47715 36373 47749
rect 36315 47681 36373 47715
rect 36315 47647 36327 47681
rect 36361 47647 36373 47681
rect 36315 47613 36373 47647
rect 36315 47579 36327 47613
rect 36361 47579 36373 47613
rect 36315 47545 36373 47579
rect 36315 47511 36327 47545
rect 36361 47511 36373 47545
rect 36315 47477 36373 47511
rect 36315 47443 36327 47477
rect 36361 47443 36373 47477
rect 36315 47427 36373 47443
rect 36773 48701 36831 48717
rect 36773 48667 36785 48701
rect 36819 48667 36831 48701
rect 36773 48633 36831 48667
rect 36773 48599 36785 48633
rect 36819 48599 36831 48633
rect 36773 48565 36831 48599
rect 36773 48531 36785 48565
rect 36819 48531 36831 48565
rect 36773 48497 36831 48531
rect 36773 48463 36785 48497
rect 36819 48463 36831 48497
rect 36773 48429 36831 48463
rect 36773 48395 36785 48429
rect 36819 48395 36831 48429
rect 36773 48361 36831 48395
rect 36773 48327 36785 48361
rect 36819 48327 36831 48361
rect 36773 48293 36831 48327
rect 36773 48259 36785 48293
rect 36819 48259 36831 48293
rect 36773 48225 36831 48259
rect 36773 48191 36785 48225
rect 36819 48191 36831 48225
rect 36773 48157 36831 48191
rect 36773 48123 36785 48157
rect 36819 48123 36831 48157
rect 36773 48089 36831 48123
rect 36773 48055 36785 48089
rect 36819 48055 36831 48089
rect 36773 48021 36831 48055
rect 36773 47987 36785 48021
rect 36819 47987 36831 48021
rect 36773 47953 36831 47987
rect 36773 47919 36785 47953
rect 36819 47919 36831 47953
rect 36773 47885 36831 47919
rect 36773 47851 36785 47885
rect 36819 47851 36831 47885
rect 36773 47817 36831 47851
rect 36773 47783 36785 47817
rect 36819 47783 36831 47817
rect 36773 47749 36831 47783
rect 36773 47715 36785 47749
rect 36819 47715 36831 47749
rect 36773 47681 36831 47715
rect 36773 47647 36785 47681
rect 36819 47647 36831 47681
rect 36773 47613 36831 47647
rect 36773 47579 36785 47613
rect 36819 47579 36831 47613
rect 36773 47545 36831 47579
rect 36773 47511 36785 47545
rect 36819 47511 36831 47545
rect 36773 47477 36831 47511
rect 36773 47443 36785 47477
rect 36819 47443 36831 47477
rect 36773 47427 36831 47443
rect 37231 48701 37289 48717
rect 37231 48667 37243 48701
rect 37277 48667 37289 48701
rect 37231 48633 37289 48667
rect 37231 48599 37243 48633
rect 37277 48599 37289 48633
rect 37231 48565 37289 48599
rect 37231 48531 37243 48565
rect 37277 48531 37289 48565
rect 37231 48497 37289 48531
rect 37231 48463 37243 48497
rect 37277 48463 37289 48497
rect 37231 48429 37289 48463
rect 37231 48395 37243 48429
rect 37277 48395 37289 48429
rect 37231 48361 37289 48395
rect 37231 48327 37243 48361
rect 37277 48327 37289 48361
rect 37231 48293 37289 48327
rect 37231 48259 37243 48293
rect 37277 48259 37289 48293
rect 37231 48225 37289 48259
rect 37231 48191 37243 48225
rect 37277 48191 37289 48225
rect 37231 48157 37289 48191
rect 37231 48123 37243 48157
rect 37277 48123 37289 48157
rect 37231 48089 37289 48123
rect 37231 48055 37243 48089
rect 37277 48055 37289 48089
rect 37231 48021 37289 48055
rect 37231 47987 37243 48021
rect 37277 47987 37289 48021
rect 37231 47953 37289 47987
rect 37231 47919 37243 47953
rect 37277 47919 37289 47953
rect 37231 47885 37289 47919
rect 37231 47851 37243 47885
rect 37277 47851 37289 47885
rect 37231 47817 37289 47851
rect 37231 47783 37243 47817
rect 37277 47783 37289 47817
rect 37231 47749 37289 47783
rect 37231 47715 37243 47749
rect 37277 47715 37289 47749
rect 37231 47681 37289 47715
rect 37231 47647 37243 47681
rect 37277 47647 37289 47681
rect 37231 47613 37289 47647
rect 37231 47579 37243 47613
rect 37277 47579 37289 47613
rect 37231 47545 37289 47579
rect 37231 47511 37243 47545
rect 37277 47511 37289 47545
rect 37231 47477 37289 47511
rect 37231 47443 37243 47477
rect 37277 47443 37289 47477
rect 37231 47427 37289 47443
rect 37689 48701 37747 48717
rect 37689 48667 37701 48701
rect 37735 48667 37747 48701
rect 37689 48633 37747 48667
rect 37689 48599 37701 48633
rect 37735 48599 37747 48633
rect 37689 48565 37747 48599
rect 37689 48531 37701 48565
rect 37735 48531 37747 48565
rect 37689 48497 37747 48531
rect 37689 48463 37701 48497
rect 37735 48463 37747 48497
rect 37689 48429 37747 48463
rect 37689 48395 37701 48429
rect 37735 48395 37747 48429
rect 37689 48361 37747 48395
rect 37689 48327 37701 48361
rect 37735 48327 37747 48361
rect 37689 48293 37747 48327
rect 37689 48259 37701 48293
rect 37735 48259 37747 48293
rect 37689 48225 37747 48259
rect 37689 48191 37701 48225
rect 37735 48191 37747 48225
rect 37689 48157 37747 48191
rect 37689 48123 37701 48157
rect 37735 48123 37747 48157
rect 37689 48089 37747 48123
rect 37689 48055 37701 48089
rect 37735 48055 37747 48089
rect 37689 48021 37747 48055
rect 37689 47987 37701 48021
rect 37735 47987 37747 48021
rect 37689 47953 37747 47987
rect 37689 47919 37701 47953
rect 37735 47919 37747 47953
rect 37689 47885 37747 47919
rect 37689 47851 37701 47885
rect 37735 47851 37747 47885
rect 37689 47817 37747 47851
rect 37689 47783 37701 47817
rect 37735 47783 37747 47817
rect 37689 47749 37747 47783
rect 37689 47715 37701 47749
rect 37735 47715 37747 47749
rect 37689 47681 37747 47715
rect 37689 47647 37701 47681
rect 37735 47647 37747 47681
rect 37689 47613 37747 47647
rect 37689 47579 37701 47613
rect 37735 47579 37747 47613
rect 37689 47545 37747 47579
rect 37689 47511 37701 47545
rect 37735 47511 37747 47545
rect 37689 47477 37747 47511
rect 37689 47443 37701 47477
rect 37735 47443 37747 47477
rect 37689 47427 37747 47443
rect 38147 48701 38205 48717
rect 38147 48667 38159 48701
rect 38193 48667 38205 48701
rect 38147 48633 38205 48667
rect 38147 48599 38159 48633
rect 38193 48599 38205 48633
rect 38147 48565 38205 48599
rect 38147 48531 38159 48565
rect 38193 48531 38205 48565
rect 38147 48497 38205 48531
rect 38147 48463 38159 48497
rect 38193 48463 38205 48497
rect 38147 48429 38205 48463
rect 38147 48395 38159 48429
rect 38193 48395 38205 48429
rect 38147 48361 38205 48395
rect 38147 48327 38159 48361
rect 38193 48327 38205 48361
rect 38147 48293 38205 48327
rect 38147 48259 38159 48293
rect 38193 48259 38205 48293
rect 38147 48225 38205 48259
rect 38147 48191 38159 48225
rect 38193 48191 38205 48225
rect 38147 48157 38205 48191
rect 38147 48123 38159 48157
rect 38193 48123 38205 48157
rect 38147 48089 38205 48123
rect 38147 48055 38159 48089
rect 38193 48055 38205 48089
rect 38147 48021 38205 48055
rect 38147 47987 38159 48021
rect 38193 47987 38205 48021
rect 38147 47953 38205 47987
rect 38147 47919 38159 47953
rect 38193 47919 38205 47953
rect 38147 47885 38205 47919
rect 38147 47851 38159 47885
rect 38193 47851 38205 47885
rect 38147 47817 38205 47851
rect 38147 47783 38159 47817
rect 38193 47783 38205 47817
rect 38147 47749 38205 47783
rect 38147 47715 38159 47749
rect 38193 47715 38205 47749
rect 38147 47681 38205 47715
rect 38147 47647 38159 47681
rect 38193 47647 38205 47681
rect 38147 47613 38205 47647
rect 38147 47579 38159 47613
rect 38193 47579 38205 47613
rect 38147 47545 38205 47579
rect 38147 47511 38159 47545
rect 38193 47511 38205 47545
rect 38147 47477 38205 47511
rect 38147 47443 38159 47477
rect 38193 47443 38205 47477
rect 38147 47427 38205 47443
rect 38605 48701 38663 48717
rect 38605 48667 38617 48701
rect 38651 48667 38663 48701
rect 38605 48633 38663 48667
rect 38605 48599 38617 48633
rect 38651 48599 38663 48633
rect 38605 48565 38663 48599
rect 38605 48531 38617 48565
rect 38651 48531 38663 48565
rect 38605 48497 38663 48531
rect 38605 48463 38617 48497
rect 38651 48463 38663 48497
rect 38605 48429 38663 48463
rect 38605 48395 38617 48429
rect 38651 48395 38663 48429
rect 38605 48361 38663 48395
rect 38605 48327 38617 48361
rect 38651 48327 38663 48361
rect 38605 48293 38663 48327
rect 38605 48259 38617 48293
rect 38651 48259 38663 48293
rect 38605 48225 38663 48259
rect 38605 48191 38617 48225
rect 38651 48191 38663 48225
rect 38605 48157 38663 48191
rect 38605 48123 38617 48157
rect 38651 48123 38663 48157
rect 38605 48089 38663 48123
rect 38605 48055 38617 48089
rect 38651 48055 38663 48089
rect 38605 48021 38663 48055
rect 38605 47987 38617 48021
rect 38651 47987 38663 48021
rect 38605 47953 38663 47987
rect 38605 47919 38617 47953
rect 38651 47919 38663 47953
rect 38605 47885 38663 47919
rect 38605 47851 38617 47885
rect 38651 47851 38663 47885
rect 38605 47817 38663 47851
rect 38605 47783 38617 47817
rect 38651 47783 38663 47817
rect 38605 47749 38663 47783
rect 38605 47715 38617 47749
rect 38651 47715 38663 47749
rect 38605 47681 38663 47715
rect 38605 47647 38617 47681
rect 38651 47647 38663 47681
rect 38605 47613 38663 47647
rect 38605 47579 38617 47613
rect 38651 47579 38663 47613
rect 38605 47545 38663 47579
rect 38605 47511 38617 47545
rect 38651 47511 38663 47545
rect 38605 47477 38663 47511
rect 38605 47443 38617 47477
rect 38651 47443 38663 47477
rect 38605 47427 38663 47443
rect 39063 48701 39121 48717
rect 39063 48667 39075 48701
rect 39109 48667 39121 48701
rect 39063 48633 39121 48667
rect 39063 48599 39075 48633
rect 39109 48599 39121 48633
rect 39063 48565 39121 48599
rect 39063 48531 39075 48565
rect 39109 48531 39121 48565
rect 39063 48497 39121 48531
rect 39063 48463 39075 48497
rect 39109 48463 39121 48497
rect 39063 48429 39121 48463
rect 39063 48395 39075 48429
rect 39109 48395 39121 48429
rect 39063 48361 39121 48395
rect 39063 48327 39075 48361
rect 39109 48327 39121 48361
rect 39063 48293 39121 48327
rect 39063 48259 39075 48293
rect 39109 48259 39121 48293
rect 39063 48225 39121 48259
rect 39063 48191 39075 48225
rect 39109 48191 39121 48225
rect 39063 48157 39121 48191
rect 39063 48123 39075 48157
rect 39109 48123 39121 48157
rect 39063 48089 39121 48123
rect 39063 48055 39075 48089
rect 39109 48055 39121 48089
rect 39063 48021 39121 48055
rect 39063 47987 39075 48021
rect 39109 47987 39121 48021
rect 39063 47953 39121 47987
rect 39063 47919 39075 47953
rect 39109 47919 39121 47953
rect 39063 47885 39121 47919
rect 39063 47851 39075 47885
rect 39109 47851 39121 47885
rect 39063 47817 39121 47851
rect 39063 47783 39075 47817
rect 39109 47783 39121 47817
rect 39063 47749 39121 47783
rect 39063 47715 39075 47749
rect 39109 47715 39121 47749
rect 39063 47681 39121 47715
rect 39063 47647 39075 47681
rect 39109 47647 39121 47681
rect 39063 47613 39121 47647
rect 39063 47579 39075 47613
rect 39109 47579 39121 47613
rect 39063 47545 39121 47579
rect 39063 47511 39075 47545
rect 39109 47511 39121 47545
rect 39063 47477 39121 47511
rect 39063 47443 39075 47477
rect 39109 47443 39121 47477
rect 39063 47427 39121 47443
rect 39521 48701 39579 48717
rect 39521 48667 39533 48701
rect 39567 48667 39579 48701
rect 39521 48633 39579 48667
rect 39521 48599 39533 48633
rect 39567 48599 39579 48633
rect 39521 48565 39579 48599
rect 39521 48531 39533 48565
rect 39567 48531 39579 48565
rect 39521 48497 39579 48531
rect 39521 48463 39533 48497
rect 39567 48463 39579 48497
rect 39521 48429 39579 48463
rect 39521 48395 39533 48429
rect 39567 48395 39579 48429
rect 39521 48361 39579 48395
rect 39521 48327 39533 48361
rect 39567 48327 39579 48361
rect 39521 48293 39579 48327
rect 39521 48259 39533 48293
rect 39567 48259 39579 48293
rect 39521 48225 39579 48259
rect 39521 48191 39533 48225
rect 39567 48191 39579 48225
rect 39521 48157 39579 48191
rect 39521 48123 39533 48157
rect 39567 48123 39579 48157
rect 39521 48089 39579 48123
rect 39521 48055 39533 48089
rect 39567 48055 39579 48089
rect 39521 48021 39579 48055
rect 39521 47987 39533 48021
rect 39567 47987 39579 48021
rect 39521 47953 39579 47987
rect 39521 47919 39533 47953
rect 39567 47919 39579 47953
rect 39521 47885 39579 47919
rect 39521 47851 39533 47885
rect 39567 47851 39579 47885
rect 39521 47817 39579 47851
rect 39521 47783 39533 47817
rect 39567 47783 39579 47817
rect 39521 47749 39579 47783
rect 39521 47715 39533 47749
rect 39567 47715 39579 47749
rect 39521 47681 39579 47715
rect 39521 47647 39533 47681
rect 39567 47647 39579 47681
rect 39521 47613 39579 47647
rect 39521 47579 39533 47613
rect 39567 47579 39579 47613
rect 39521 47545 39579 47579
rect 39521 47511 39533 47545
rect 39567 47511 39579 47545
rect 39521 47477 39579 47511
rect 39521 47443 39533 47477
rect 39567 47443 39579 47477
rect 39521 47427 39579 47443
rect 39979 48701 40037 48717
rect 39979 48667 39991 48701
rect 40025 48667 40037 48701
rect 39979 48633 40037 48667
rect 39979 48599 39991 48633
rect 40025 48599 40037 48633
rect 39979 48565 40037 48599
rect 39979 48531 39991 48565
rect 40025 48531 40037 48565
rect 39979 48497 40037 48531
rect 39979 48463 39991 48497
rect 40025 48463 40037 48497
rect 39979 48429 40037 48463
rect 39979 48395 39991 48429
rect 40025 48395 40037 48429
rect 39979 48361 40037 48395
rect 39979 48327 39991 48361
rect 40025 48327 40037 48361
rect 39979 48293 40037 48327
rect 39979 48259 39991 48293
rect 40025 48259 40037 48293
rect 39979 48225 40037 48259
rect 39979 48191 39991 48225
rect 40025 48191 40037 48225
rect 39979 48157 40037 48191
rect 39979 48123 39991 48157
rect 40025 48123 40037 48157
rect 39979 48089 40037 48123
rect 39979 48055 39991 48089
rect 40025 48055 40037 48089
rect 39979 48021 40037 48055
rect 39979 47987 39991 48021
rect 40025 47987 40037 48021
rect 39979 47953 40037 47987
rect 39979 47919 39991 47953
rect 40025 47919 40037 47953
rect 39979 47885 40037 47919
rect 39979 47851 39991 47885
rect 40025 47851 40037 47885
rect 39979 47817 40037 47851
rect 39979 47783 39991 47817
rect 40025 47783 40037 47817
rect 39979 47749 40037 47783
rect 39979 47715 39991 47749
rect 40025 47715 40037 47749
rect 39979 47681 40037 47715
rect 39979 47647 39991 47681
rect 40025 47647 40037 47681
rect 39979 47613 40037 47647
rect 39979 47579 39991 47613
rect 40025 47579 40037 47613
rect 39979 47545 40037 47579
rect 39979 47511 39991 47545
rect 40025 47511 40037 47545
rect 39979 47477 40037 47511
rect 39979 47443 39991 47477
rect 40025 47443 40037 47477
rect 39979 47427 40037 47443
rect 40437 48701 40495 48717
rect 40437 48667 40449 48701
rect 40483 48667 40495 48701
rect 40437 48633 40495 48667
rect 40437 48599 40449 48633
rect 40483 48599 40495 48633
rect 40437 48565 40495 48599
rect 40437 48531 40449 48565
rect 40483 48531 40495 48565
rect 40437 48497 40495 48531
rect 40437 48463 40449 48497
rect 40483 48463 40495 48497
rect 40437 48429 40495 48463
rect 40437 48395 40449 48429
rect 40483 48395 40495 48429
rect 40437 48361 40495 48395
rect 40437 48327 40449 48361
rect 40483 48327 40495 48361
rect 40437 48293 40495 48327
rect 40437 48259 40449 48293
rect 40483 48259 40495 48293
rect 40437 48225 40495 48259
rect 40437 48191 40449 48225
rect 40483 48191 40495 48225
rect 40437 48157 40495 48191
rect 40437 48123 40449 48157
rect 40483 48123 40495 48157
rect 40437 48089 40495 48123
rect 40437 48055 40449 48089
rect 40483 48055 40495 48089
rect 40437 48021 40495 48055
rect 40437 47987 40449 48021
rect 40483 47987 40495 48021
rect 40437 47953 40495 47987
rect 40437 47919 40449 47953
rect 40483 47919 40495 47953
rect 40437 47885 40495 47919
rect 40437 47851 40449 47885
rect 40483 47851 40495 47885
rect 40437 47817 40495 47851
rect 40437 47783 40449 47817
rect 40483 47783 40495 47817
rect 40437 47749 40495 47783
rect 40437 47715 40449 47749
rect 40483 47715 40495 47749
rect 40437 47681 40495 47715
rect 40437 47647 40449 47681
rect 40483 47647 40495 47681
rect 40437 47613 40495 47647
rect 40437 47579 40449 47613
rect 40483 47579 40495 47613
rect 40437 47545 40495 47579
rect 40437 47511 40449 47545
rect 40483 47511 40495 47545
rect 40437 47477 40495 47511
rect 40437 47443 40449 47477
rect 40483 47443 40495 47477
rect 40437 47427 40495 47443
rect 40895 48701 40953 48717
rect 40895 48667 40907 48701
rect 40941 48667 40953 48701
rect 40895 48633 40953 48667
rect 40895 48599 40907 48633
rect 40941 48599 40953 48633
rect 40895 48565 40953 48599
rect 40895 48531 40907 48565
rect 40941 48531 40953 48565
rect 40895 48497 40953 48531
rect 40895 48463 40907 48497
rect 40941 48463 40953 48497
rect 40895 48429 40953 48463
rect 40895 48395 40907 48429
rect 40941 48395 40953 48429
rect 40895 48361 40953 48395
rect 40895 48327 40907 48361
rect 40941 48327 40953 48361
rect 40895 48293 40953 48327
rect 40895 48259 40907 48293
rect 40941 48259 40953 48293
rect 40895 48225 40953 48259
rect 40895 48191 40907 48225
rect 40941 48191 40953 48225
rect 40895 48157 40953 48191
rect 40895 48123 40907 48157
rect 40941 48123 40953 48157
rect 40895 48089 40953 48123
rect 40895 48055 40907 48089
rect 40941 48055 40953 48089
rect 40895 48021 40953 48055
rect 40895 47987 40907 48021
rect 40941 47987 40953 48021
rect 40895 47953 40953 47987
rect 40895 47919 40907 47953
rect 40941 47919 40953 47953
rect 40895 47885 40953 47919
rect 40895 47851 40907 47885
rect 40941 47851 40953 47885
rect 40895 47817 40953 47851
rect 40895 47783 40907 47817
rect 40941 47783 40953 47817
rect 40895 47749 40953 47783
rect 40895 47715 40907 47749
rect 40941 47715 40953 47749
rect 40895 47681 40953 47715
rect 40895 47647 40907 47681
rect 40941 47647 40953 47681
rect 40895 47613 40953 47647
rect 40895 47579 40907 47613
rect 40941 47579 40953 47613
rect 40895 47545 40953 47579
rect 40895 47511 40907 47545
rect 40941 47511 40953 47545
rect 40895 47477 40953 47511
rect 40895 47443 40907 47477
rect 40941 47443 40953 47477
rect 40895 47427 40953 47443
rect 41353 48701 41411 48717
rect 41353 48667 41365 48701
rect 41399 48667 41411 48701
rect 41353 48633 41411 48667
rect 41353 48599 41365 48633
rect 41399 48599 41411 48633
rect 41353 48565 41411 48599
rect 41353 48531 41365 48565
rect 41399 48531 41411 48565
rect 41353 48497 41411 48531
rect 41353 48463 41365 48497
rect 41399 48463 41411 48497
rect 41353 48429 41411 48463
rect 41353 48395 41365 48429
rect 41399 48395 41411 48429
rect 41353 48361 41411 48395
rect 41353 48327 41365 48361
rect 41399 48327 41411 48361
rect 41353 48293 41411 48327
rect 41353 48259 41365 48293
rect 41399 48259 41411 48293
rect 41353 48225 41411 48259
rect 41353 48191 41365 48225
rect 41399 48191 41411 48225
rect 41353 48157 41411 48191
rect 41353 48123 41365 48157
rect 41399 48123 41411 48157
rect 41353 48089 41411 48123
rect 41353 48055 41365 48089
rect 41399 48055 41411 48089
rect 41353 48021 41411 48055
rect 41353 47987 41365 48021
rect 41399 47987 41411 48021
rect 41353 47953 41411 47987
rect 41353 47919 41365 47953
rect 41399 47919 41411 47953
rect 41353 47885 41411 47919
rect 41353 47851 41365 47885
rect 41399 47851 41411 47885
rect 41353 47817 41411 47851
rect 41353 47783 41365 47817
rect 41399 47783 41411 47817
rect 41353 47749 41411 47783
rect 41353 47715 41365 47749
rect 41399 47715 41411 47749
rect 41353 47681 41411 47715
rect 41353 47647 41365 47681
rect 41399 47647 41411 47681
rect 41353 47613 41411 47647
rect 41353 47579 41365 47613
rect 41399 47579 41411 47613
rect 41353 47545 41411 47579
rect 41353 47511 41365 47545
rect 41399 47511 41411 47545
rect 41353 47477 41411 47511
rect 41353 47443 41365 47477
rect 41399 47443 41411 47477
rect 41353 47427 41411 47443
rect 41811 48701 41869 48717
rect 41811 48667 41823 48701
rect 41857 48667 41869 48701
rect 41811 48633 41869 48667
rect 41811 48599 41823 48633
rect 41857 48599 41869 48633
rect 41811 48565 41869 48599
rect 41811 48531 41823 48565
rect 41857 48531 41869 48565
rect 41811 48497 41869 48531
rect 41811 48463 41823 48497
rect 41857 48463 41869 48497
rect 41811 48429 41869 48463
rect 41811 48395 41823 48429
rect 41857 48395 41869 48429
rect 41811 48361 41869 48395
rect 41811 48327 41823 48361
rect 41857 48327 41869 48361
rect 41811 48293 41869 48327
rect 41811 48259 41823 48293
rect 41857 48259 41869 48293
rect 41811 48225 41869 48259
rect 41811 48191 41823 48225
rect 41857 48191 41869 48225
rect 41811 48157 41869 48191
rect 41811 48123 41823 48157
rect 41857 48123 41869 48157
rect 41811 48089 41869 48123
rect 41811 48055 41823 48089
rect 41857 48055 41869 48089
rect 41811 48021 41869 48055
rect 41811 47987 41823 48021
rect 41857 47987 41869 48021
rect 41811 47953 41869 47987
rect 41811 47919 41823 47953
rect 41857 47919 41869 47953
rect 41811 47885 41869 47919
rect 41811 47851 41823 47885
rect 41857 47851 41869 47885
rect 41811 47817 41869 47851
rect 41811 47783 41823 47817
rect 41857 47783 41869 47817
rect 41811 47749 41869 47783
rect 41811 47715 41823 47749
rect 41857 47715 41869 47749
rect 41811 47681 41869 47715
rect 41811 47647 41823 47681
rect 41857 47647 41869 47681
rect 41811 47613 41869 47647
rect 41811 47579 41823 47613
rect 41857 47579 41869 47613
rect 41811 47545 41869 47579
rect 41811 47511 41823 47545
rect 41857 47511 41869 47545
rect 41811 47477 41869 47511
rect 41811 47443 41823 47477
rect 41857 47443 41869 47477
rect 41811 47427 41869 47443
rect 42269 48701 42327 48717
rect 42269 48667 42281 48701
rect 42315 48667 42327 48701
rect 42269 48633 42327 48667
rect 42269 48599 42281 48633
rect 42315 48599 42327 48633
rect 42269 48565 42327 48599
rect 42269 48531 42281 48565
rect 42315 48531 42327 48565
rect 42269 48497 42327 48531
rect 42269 48463 42281 48497
rect 42315 48463 42327 48497
rect 42269 48429 42327 48463
rect 42269 48395 42281 48429
rect 42315 48395 42327 48429
rect 42269 48361 42327 48395
rect 42269 48327 42281 48361
rect 42315 48327 42327 48361
rect 42269 48293 42327 48327
rect 42269 48259 42281 48293
rect 42315 48259 42327 48293
rect 42269 48225 42327 48259
rect 42269 48191 42281 48225
rect 42315 48191 42327 48225
rect 42269 48157 42327 48191
rect 42269 48123 42281 48157
rect 42315 48123 42327 48157
rect 42269 48089 42327 48123
rect 42269 48055 42281 48089
rect 42315 48055 42327 48089
rect 42269 48021 42327 48055
rect 42269 47987 42281 48021
rect 42315 47987 42327 48021
rect 42269 47953 42327 47987
rect 42269 47919 42281 47953
rect 42315 47919 42327 47953
rect 42269 47885 42327 47919
rect 42269 47851 42281 47885
rect 42315 47851 42327 47885
rect 42269 47817 42327 47851
rect 42269 47783 42281 47817
rect 42315 47783 42327 47817
rect 42269 47749 42327 47783
rect 42269 47715 42281 47749
rect 42315 47715 42327 47749
rect 42269 47681 42327 47715
rect 42269 47647 42281 47681
rect 42315 47647 42327 47681
rect 42269 47613 42327 47647
rect 42269 47579 42281 47613
rect 42315 47579 42327 47613
rect 42269 47545 42327 47579
rect 42269 47511 42281 47545
rect 42315 47511 42327 47545
rect 42269 47477 42327 47511
rect 42269 47443 42281 47477
rect 42315 47443 42327 47477
rect 42269 47427 42327 47443
rect 42727 48701 42785 48717
rect 42727 48667 42739 48701
rect 42773 48667 42785 48701
rect 42727 48633 42785 48667
rect 42727 48599 42739 48633
rect 42773 48599 42785 48633
rect 42727 48565 42785 48599
rect 42727 48531 42739 48565
rect 42773 48531 42785 48565
rect 42727 48497 42785 48531
rect 42727 48463 42739 48497
rect 42773 48463 42785 48497
rect 42727 48429 42785 48463
rect 42727 48395 42739 48429
rect 42773 48395 42785 48429
rect 42727 48361 42785 48395
rect 42727 48327 42739 48361
rect 42773 48327 42785 48361
rect 42727 48293 42785 48327
rect 42727 48259 42739 48293
rect 42773 48259 42785 48293
rect 42727 48225 42785 48259
rect 42727 48191 42739 48225
rect 42773 48191 42785 48225
rect 42727 48157 42785 48191
rect 42727 48123 42739 48157
rect 42773 48123 42785 48157
rect 42727 48089 42785 48123
rect 42727 48055 42739 48089
rect 42773 48055 42785 48089
rect 42727 48021 42785 48055
rect 42727 47987 42739 48021
rect 42773 47987 42785 48021
rect 42727 47953 42785 47987
rect 42727 47919 42739 47953
rect 42773 47919 42785 47953
rect 42727 47885 42785 47919
rect 42727 47851 42739 47885
rect 42773 47851 42785 47885
rect 42727 47817 42785 47851
rect 42727 47783 42739 47817
rect 42773 47783 42785 47817
rect 42727 47749 42785 47783
rect 42727 47715 42739 47749
rect 42773 47715 42785 47749
rect 42727 47681 42785 47715
rect 42727 47647 42739 47681
rect 42773 47647 42785 47681
rect 42727 47613 42785 47647
rect 42727 47579 42739 47613
rect 42773 47579 42785 47613
rect 42727 47545 42785 47579
rect 42727 47511 42739 47545
rect 42773 47511 42785 47545
rect 42727 47477 42785 47511
rect 42727 47443 42739 47477
rect 42773 47443 42785 47477
rect 42727 47427 42785 47443
rect 43185 48701 43243 48717
rect 43185 48667 43197 48701
rect 43231 48667 43243 48701
rect 43185 48633 43243 48667
rect 43185 48599 43197 48633
rect 43231 48599 43243 48633
rect 43185 48565 43243 48599
rect 43185 48531 43197 48565
rect 43231 48531 43243 48565
rect 43185 48497 43243 48531
rect 43185 48463 43197 48497
rect 43231 48463 43243 48497
rect 43185 48429 43243 48463
rect 43185 48395 43197 48429
rect 43231 48395 43243 48429
rect 43185 48361 43243 48395
rect 43185 48327 43197 48361
rect 43231 48327 43243 48361
rect 43185 48293 43243 48327
rect 43185 48259 43197 48293
rect 43231 48259 43243 48293
rect 43185 48225 43243 48259
rect 43185 48191 43197 48225
rect 43231 48191 43243 48225
rect 43185 48157 43243 48191
rect 43185 48123 43197 48157
rect 43231 48123 43243 48157
rect 43185 48089 43243 48123
rect 43185 48055 43197 48089
rect 43231 48055 43243 48089
rect 43185 48021 43243 48055
rect 43185 47987 43197 48021
rect 43231 47987 43243 48021
rect 43185 47953 43243 47987
rect 43185 47919 43197 47953
rect 43231 47919 43243 47953
rect 43185 47885 43243 47919
rect 43185 47851 43197 47885
rect 43231 47851 43243 47885
rect 43185 47817 43243 47851
rect 43185 47783 43197 47817
rect 43231 47783 43243 47817
rect 43185 47749 43243 47783
rect 43185 47715 43197 47749
rect 43231 47715 43243 47749
rect 43185 47681 43243 47715
rect 43185 47647 43197 47681
rect 43231 47647 43243 47681
rect 43185 47613 43243 47647
rect 43185 47579 43197 47613
rect 43231 47579 43243 47613
rect 43185 47545 43243 47579
rect 43185 47511 43197 47545
rect 43231 47511 43243 47545
rect 43185 47477 43243 47511
rect 43185 47443 43197 47477
rect 43231 47443 43243 47477
rect 43185 47427 43243 47443
rect 43643 48701 43701 48717
rect 43643 48667 43655 48701
rect 43689 48667 43701 48701
rect 43643 48633 43701 48667
rect 43643 48599 43655 48633
rect 43689 48599 43701 48633
rect 43643 48565 43701 48599
rect 43643 48531 43655 48565
rect 43689 48531 43701 48565
rect 43643 48497 43701 48531
rect 43643 48463 43655 48497
rect 43689 48463 43701 48497
rect 43643 48429 43701 48463
rect 43643 48395 43655 48429
rect 43689 48395 43701 48429
rect 43643 48361 43701 48395
rect 43643 48327 43655 48361
rect 43689 48327 43701 48361
rect 43643 48293 43701 48327
rect 43643 48259 43655 48293
rect 43689 48259 43701 48293
rect 43643 48225 43701 48259
rect 43643 48191 43655 48225
rect 43689 48191 43701 48225
rect 43643 48157 43701 48191
rect 43643 48123 43655 48157
rect 43689 48123 43701 48157
rect 43643 48089 43701 48123
rect 43643 48055 43655 48089
rect 43689 48055 43701 48089
rect 43643 48021 43701 48055
rect 43643 47987 43655 48021
rect 43689 47987 43701 48021
rect 43643 47953 43701 47987
rect 43643 47919 43655 47953
rect 43689 47919 43701 47953
rect 43643 47885 43701 47919
rect 43643 47851 43655 47885
rect 43689 47851 43701 47885
rect 43643 47817 43701 47851
rect 43643 47783 43655 47817
rect 43689 47783 43701 47817
rect 43643 47749 43701 47783
rect 43643 47715 43655 47749
rect 43689 47715 43701 47749
rect 43643 47681 43701 47715
rect 43643 47647 43655 47681
rect 43689 47647 43701 47681
rect 43643 47613 43701 47647
rect 43643 47579 43655 47613
rect 43689 47579 43701 47613
rect 43643 47545 43701 47579
rect 43643 47511 43655 47545
rect 43689 47511 43701 47545
rect 43643 47477 43701 47511
rect 43643 47443 43655 47477
rect 43689 47443 43701 47477
rect 43643 47427 43701 47443
rect 44101 48701 44159 48717
rect 44101 48667 44113 48701
rect 44147 48667 44159 48701
rect 44101 48633 44159 48667
rect 44101 48599 44113 48633
rect 44147 48599 44159 48633
rect 44101 48565 44159 48599
rect 44101 48531 44113 48565
rect 44147 48531 44159 48565
rect 44101 48497 44159 48531
rect 44101 48463 44113 48497
rect 44147 48463 44159 48497
rect 44101 48429 44159 48463
rect 44101 48395 44113 48429
rect 44147 48395 44159 48429
rect 44101 48361 44159 48395
rect 44101 48327 44113 48361
rect 44147 48327 44159 48361
rect 44101 48293 44159 48327
rect 44101 48259 44113 48293
rect 44147 48259 44159 48293
rect 44101 48225 44159 48259
rect 44101 48191 44113 48225
rect 44147 48191 44159 48225
rect 44101 48157 44159 48191
rect 44101 48123 44113 48157
rect 44147 48123 44159 48157
rect 44101 48089 44159 48123
rect 44101 48055 44113 48089
rect 44147 48055 44159 48089
rect 44101 48021 44159 48055
rect 44101 47987 44113 48021
rect 44147 47987 44159 48021
rect 44101 47953 44159 47987
rect 44101 47919 44113 47953
rect 44147 47919 44159 47953
rect 44101 47885 44159 47919
rect 44101 47851 44113 47885
rect 44147 47851 44159 47885
rect 44101 47817 44159 47851
rect 44101 47783 44113 47817
rect 44147 47783 44159 47817
rect 44101 47749 44159 47783
rect 44101 47715 44113 47749
rect 44147 47715 44159 47749
rect 44101 47681 44159 47715
rect 44101 47647 44113 47681
rect 44147 47647 44159 47681
rect 44101 47613 44159 47647
rect 44101 47579 44113 47613
rect 44147 47579 44159 47613
rect 44101 47545 44159 47579
rect 44101 47511 44113 47545
rect 44147 47511 44159 47545
rect 44101 47477 44159 47511
rect 44101 47443 44113 47477
rect 44147 47443 44159 47477
rect 44101 47427 44159 47443
rect 44559 48701 44617 48717
rect 44559 48667 44571 48701
rect 44605 48667 44617 48701
rect 44559 48633 44617 48667
rect 44559 48599 44571 48633
rect 44605 48599 44617 48633
rect 44559 48565 44617 48599
rect 44559 48531 44571 48565
rect 44605 48531 44617 48565
rect 44559 48497 44617 48531
rect 44559 48463 44571 48497
rect 44605 48463 44617 48497
rect 44559 48429 44617 48463
rect 44559 48395 44571 48429
rect 44605 48395 44617 48429
rect 44559 48361 44617 48395
rect 44559 48327 44571 48361
rect 44605 48327 44617 48361
rect 44559 48293 44617 48327
rect 44559 48259 44571 48293
rect 44605 48259 44617 48293
rect 44559 48225 44617 48259
rect 44559 48191 44571 48225
rect 44605 48191 44617 48225
rect 44559 48157 44617 48191
rect 44559 48123 44571 48157
rect 44605 48123 44617 48157
rect 44559 48089 44617 48123
rect 44559 48055 44571 48089
rect 44605 48055 44617 48089
rect 44559 48021 44617 48055
rect 44559 47987 44571 48021
rect 44605 47987 44617 48021
rect 44559 47953 44617 47987
rect 44559 47919 44571 47953
rect 44605 47919 44617 47953
rect 44559 47885 44617 47919
rect 44559 47851 44571 47885
rect 44605 47851 44617 47885
rect 44559 47817 44617 47851
rect 44559 47783 44571 47817
rect 44605 47783 44617 47817
rect 44559 47749 44617 47783
rect 44559 47715 44571 47749
rect 44605 47715 44617 47749
rect 44559 47681 44617 47715
rect 44559 47647 44571 47681
rect 44605 47647 44617 47681
rect 44559 47613 44617 47647
rect 44559 47579 44571 47613
rect 44605 47579 44617 47613
rect 44559 47545 44617 47579
rect 44559 47511 44571 47545
rect 44605 47511 44617 47545
rect 44559 47477 44617 47511
rect 44559 47443 44571 47477
rect 44605 47443 44617 47477
rect 44559 47427 44617 47443
rect 45017 48701 45075 48717
rect 45017 48667 45029 48701
rect 45063 48667 45075 48701
rect 45017 48633 45075 48667
rect 45017 48599 45029 48633
rect 45063 48599 45075 48633
rect 45017 48565 45075 48599
rect 45017 48531 45029 48565
rect 45063 48531 45075 48565
rect 45017 48497 45075 48531
rect 45017 48463 45029 48497
rect 45063 48463 45075 48497
rect 45017 48429 45075 48463
rect 45017 48395 45029 48429
rect 45063 48395 45075 48429
rect 45017 48361 45075 48395
rect 45017 48327 45029 48361
rect 45063 48327 45075 48361
rect 45017 48293 45075 48327
rect 45017 48259 45029 48293
rect 45063 48259 45075 48293
rect 45017 48225 45075 48259
rect 45017 48191 45029 48225
rect 45063 48191 45075 48225
rect 45017 48157 45075 48191
rect 45017 48123 45029 48157
rect 45063 48123 45075 48157
rect 45017 48089 45075 48123
rect 45017 48055 45029 48089
rect 45063 48055 45075 48089
rect 45017 48021 45075 48055
rect 45017 47987 45029 48021
rect 45063 47987 45075 48021
rect 45017 47953 45075 47987
rect 45017 47919 45029 47953
rect 45063 47919 45075 47953
rect 45017 47885 45075 47919
rect 45017 47851 45029 47885
rect 45063 47851 45075 47885
rect 45017 47817 45075 47851
rect 45017 47783 45029 47817
rect 45063 47783 45075 47817
rect 45017 47749 45075 47783
rect 45017 47715 45029 47749
rect 45063 47715 45075 47749
rect 45017 47681 45075 47715
rect 45017 47647 45029 47681
rect 45063 47647 45075 47681
rect 45017 47613 45075 47647
rect 45017 47579 45029 47613
rect 45063 47579 45075 47613
rect 45017 47545 45075 47579
rect 45017 47511 45029 47545
rect 45063 47511 45075 47545
rect 45017 47477 45075 47511
rect 45017 47443 45029 47477
rect 45063 47443 45075 47477
rect 45017 47427 45075 47443
rect 45475 48701 45533 48717
rect 45475 48667 45487 48701
rect 45521 48667 45533 48701
rect 45475 48633 45533 48667
rect 45475 48599 45487 48633
rect 45521 48599 45533 48633
rect 45475 48565 45533 48599
rect 45475 48531 45487 48565
rect 45521 48531 45533 48565
rect 45475 48497 45533 48531
rect 45475 48463 45487 48497
rect 45521 48463 45533 48497
rect 45475 48429 45533 48463
rect 45475 48395 45487 48429
rect 45521 48395 45533 48429
rect 45475 48361 45533 48395
rect 45475 48327 45487 48361
rect 45521 48327 45533 48361
rect 45475 48293 45533 48327
rect 45475 48259 45487 48293
rect 45521 48259 45533 48293
rect 45475 48225 45533 48259
rect 45475 48191 45487 48225
rect 45521 48191 45533 48225
rect 45475 48157 45533 48191
rect 45475 48123 45487 48157
rect 45521 48123 45533 48157
rect 45475 48089 45533 48123
rect 45475 48055 45487 48089
rect 45521 48055 45533 48089
rect 45475 48021 45533 48055
rect 45475 47987 45487 48021
rect 45521 47987 45533 48021
rect 45475 47953 45533 47987
rect 45475 47919 45487 47953
rect 45521 47919 45533 47953
rect 45475 47885 45533 47919
rect 45475 47851 45487 47885
rect 45521 47851 45533 47885
rect 45475 47817 45533 47851
rect 45475 47783 45487 47817
rect 45521 47783 45533 47817
rect 45475 47749 45533 47783
rect 45475 47715 45487 47749
rect 45521 47715 45533 47749
rect 45475 47681 45533 47715
rect 45475 47647 45487 47681
rect 45521 47647 45533 47681
rect 45475 47613 45533 47647
rect 45475 47579 45487 47613
rect 45521 47579 45533 47613
rect 45475 47545 45533 47579
rect 45475 47511 45487 47545
rect 45521 47511 45533 47545
rect 45475 47477 45533 47511
rect 45475 47443 45487 47477
rect 45521 47443 45533 47477
rect 45475 47427 45533 47443
rect 45933 48701 45991 48717
rect 45933 48667 45945 48701
rect 45979 48667 45991 48701
rect 45933 48633 45991 48667
rect 45933 48599 45945 48633
rect 45979 48599 45991 48633
rect 45933 48565 45991 48599
rect 45933 48531 45945 48565
rect 45979 48531 45991 48565
rect 45933 48497 45991 48531
rect 45933 48463 45945 48497
rect 45979 48463 45991 48497
rect 45933 48429 45991 48463
rect 45933 48395 45945 48429
rect 45979 48395 45991 48429
rect 45933 48361 45991 48395
rect 45933 48327 45945 48361
rect 45979 48327 45991 48361
rect 45933 48293 45991 48327
rect 45933 48259 45945 48293
rect 45979 48259 45991 48293
rect 45933 48225 45991 48259
rect 45933 48191 45945 48225
rect 45979 48191 45991 48225
rect 45933 48157 45991 48191
rect 45933 48123 45945 48157
rect 45979 48123 45991 48157
rect 45933 48089 45991 48123
rect 45933 48055 45945 48089
rect 45979 48055 45991 48089
rect 45933 48021 45991 48055
rect 45933 47987 45945 48021
rect 45979 47987 45991 48021
rect 45933 47953 45991 47987
rect 45933 47919 45945 47953
rect 45979 47919 45991 47953
rect 45933 47885 45991 47919
rect 45933 47851 45945 47885
rect 45979 47851 45991 47885
rect 45933 47817 45991 47851
rect 45933 47783 45945 47817
rect 45979 47783 45991 47817
rect 45933 47749 45991 47783
rect 45933 47715 45945 47749
rect 45979 47715 45991 47749
rect 45933 47681 45991 47715
rect 45933 47647 45945 47681
rect 45979 47647 45991 47681
rect 45933 47613 45991 47647
rect 45933 47579 45945 47613
rect 45979 47579 45991 47613
rect 45933 47545 45991 47579
rect 45933 47511 45945 47545
rect 45979 47511 45991 47545
rect 45933 47477 45991 47511
rect 45933 47443 45945 47477
rect 45979 47443 45991 47477
rect 45933 47427 45991 47443
rect 46391 48701 46449 48717
rect 46391 48667 46403 48701
rect 46437 48667 46449 48701
rect 46391 48633 46449 48667
rect 46391 48599 46403 48633
rect 46437 48599 46449 48633
rect 46391 48565 46449 48599
rect 46391 48531 46403 48565
rect 46437 48531 46449 48565
rect 46391 48497 46449 48531
rect 46391 48463 46403 48497
rect 46437 48463 46449 48497
rect 46391 48429 46449 48463
rect 46391 48395 46403 48429
rect 46437 48395 46449 48429
rect 46391 48361 46449 48395
rect 46391 48327 46403 48361
rect 46437 48327 46449 48361
rect 46391 48293 46449 48327
rect 46391 48259 46403 48293
rect 46437 48259 46449 48293
rect 46391 48225 46449 48259
rect 46391 48191 46403 48225
rect 46437 48191 46449 48225
rect 46391 48157 46449 48191
rect 46391 48123 46403 48157
rect 46437 48123 46449 48157
rect 46391 48089 46449 48123
rect 46391 48055 46403 48089
rect 46437 48055 46449 48089
rect 46391 48021 46449 48055
rect 46391 47987 46403 48021
rect 46437 47987 46449 48021
rect 46391 47953 46449 47987
rect 46391 47919 46403 47953
rect 46437 47919 46449 47953
rect 46391 47885 46449 47919
rect 46391 47851 46403 47885
rect 46437 47851 46449 47885
rect 46391 47817 46449 47851
rect 46391 47783 46403 47817
rect 46437 47783 46449 47817
rect 46391 47749 46449 47783
rect 46391 47715 46403 47749
rect 46437 47715 46449 47749
rect 46391 47681 46449 47715
rect 46391 47647 46403 47681
rect 46437 47647 46449 47681
rect 46391 47613 46449 47647
rect 46391 47579 46403 47613
rect 46437 47579 46449 47613
rect 46391 47545 46449 47579
rect 46391 47511 46403 47545
rect 46437 47511 46449 47545
rect 46391 47477 46449 47511
rect 46391 47443 46403 47477
rect 46437 47443 46449 47477
rect 46391 47427 46449 47443
rect 46849 48701 46907 48717
rect 46849 48667 46861 48701
rect 46895 48667 46907 48701
rect 46849 48633 46907 48667
rect 46849 48599 46861 48633
rect 46895 48599 46907 48633
rect 46849 48565 46907 48599
rect 46849 48531 46861 48565
rect 46895 48531 46907 48565
rect 46849 48497 46907 48531
rect 46849 48463 46861 48497
rect 46895 48463 46907 48497
rect 46849 48429 46907 48463
rect 46849 48395 46861 48429
rect 46895 48395 46907 48429
rect 46849 48361 46907 48395
rect 46849 48327 46861 48361
rect 46895 48327 46907 48361
rect 46849 48293 46907 48327
rect 46849 48259 46861 48293
rect 46895 48259 46907 48293
rect 46849 48225 46907 48259
rect 46849 48191 46861 48225
rect 46895 48191 46907 48225
rect 46849 48157 46907 48191
rect 46849 48123 46861 48157
rect 46895 48123 46907 48157
rect 46849 48089 46907 48123
rect 46849 48055 46861 48089
rect 46895 48055 46907 48089
rect 46849 48021 46907 48055
rect 46849 47987 46861 48021
rect 46895 47987 46907 48021
rect 46849 47953 46907 47987
rect 46849 47919 46861 47953
rect 46895 47919 46907 47953
rect 46849 47885 46907 47919
rect 46849 47851 46861 47885
rect 46895 47851 46907 47885
rect 46849 47817 46907 47851
rect 46849 47783 46861 47817
rect 46895 47783 46907 47817
rect 46849 47749 46907 47783
rect 46849 47715 46861 47749
rect 46895 47715 46907 47749
rect 46849 47681 46907 47715
rect 46849 47647 46861 47681
rect 46895 47647 46907 47681
rect 46849 47613 46907 47647
rect 46849 47579 46861 47613
rect 46895 47579 46907 47613
rect 46849 47545 46907 47579
rect 46849 47511 46861 47545
rect 46895 47511 46907 47545
rect 46849 47477 46907 47511
rect 46849 47443 46861 47477
rect 46895 47443 46907 47477
rect 46849 47427 46907 47443
rect 47307 48701 47365 48717
rect 47307 48667 47319 48701
rect 47353 48667 47365 48701
rect 47307 48633 47365 48667
rect 47307 48599 47319 48633
rect 47353 48599 47365 48633
rect 47307 48565 47365 48599
rect 47307 48531 47319 48565
rect 47353 48531 47365 48565
rect 47307 48497 47365 48531
rect 47307 48463 47319 48497
rect 47353 48463 47365 48497
rect 47307 48429 47365 48463
rect 47307 48395 47319 48429
rect 47353 48395 47365 48429
rect 47307 48361 47365 48395
rect 47307 48327 47319 48361
rect 47353 48327 47365 48361
rect 47307 48293 47365 48327
rect 47307 48259 47319 48293
rect 47353 48259 47365 48293
rect 47307 48225 47365 48259
rect 47307 48191 47319 48225
rect 47353 48191 47365 48225
rect 47307 48157 47365 48191
rect 47307 48123 47319 48157
rect 47353 48123 47365 48157
rect 47307 48089 47365 48123
rect 47307 48055 47319 48089
rect 47353 48055 47365 48089
rect 47307 48021 47365 48055
rect 47307 47987 47319 48021
rect 47353 47987 47365 48021
rect 47307 47953 47365 47987
rect 47307 47919 47319 47953
rect 47353 47919 47365 47953
rect 47307 47885 47365 47919
rect 47307 47851 47319 47885
rect 47353 47851 47365 47885
rect 47307 47817 47365 47851
rect 47307 47783 47319 47817
rect 47353 47783 47365 47817
rect 47307 47749 47365 47783
rect 47307 47715 47319 47749
rect 47353 47715 47365 47749
rect 47307 47681 47365 47715
rect 47307 47647 47319 47681
rect 47353 47647 47365 47681
rect 47307 47613 47365 47647
rect 47307 47579 47319 47613
rect 47353 47579 47365 47613
rect 47307 47545 47365 47579
rect 47307 47511 47319 47545
rect 47353 47511 47365 47545
rect 47307 47477 47365 47511
rect 47307 47443 47319 47477
rect 47353 47443 47365 47477
rect 47307 47427 47365 47443
rect 47765 48701 47823 48717
rect 47765 48667 47777 48701
rect 47811 48667 47823 48701
rect 47765 48633 47823 48667
rect 47765 48599 47777 48633
rect 47811 48599 47823 48633
rect 47765 48565 47823 48599
rect 47765 48531 47777 48565
rect 47811 48531 47823 48565
rect 47765 48497 47823 48531
rect 47765 48463 47777 48497
rect 47811 48463 47823 48497
rect 47765 48429 47823 48463
rect 47765 48395 47777 48429
rect 47811 48395 47823 48429
rect 47765 48361 47823 48395
rect 47765 48327 47777 48361
rect 47811 48327 47823 48361
rect 47765 48293 47823 48327
rect 47765 48259 47777 48293
rect 47811 48259 47823 48293
rect 47765 48225 47823 48259
rect 47765 48191 47777 48225
rect 47811 48191 47823 48225
rect 47765 48157 47823 48191
rect 47765 48123 47777 48157
rect 47811 48123 47823 48157
rect 47765 48089 47823 48123
rect 47765 48055 47777 48089
rect 47811 48055 47823 48089
rect 47765 48021 47823 48055
rect 47765 47987 47777 48021
rect 47811 47987 47823 48021
rect 47765 47953 47823 47987
rect 47765 47919 47777 47953
rect 47811 47919 47823 47953
rect 47765 47885 47823 47919
rect 47765 47851 47777 47885
rect 47811 47851 47823 47885
rect 47765 47817 47823 47851
rect 47765 47783 47777 47817
rect 47811 47783 47823 47817
rect 47765 47749 47823 47783
rect 47765 47715 47777 47749
rect 47811 47715 47823 47749
rect 47765 47681 47823 47715
rect 47765 47647 47777 47681
rect 47811 47647 47823 47681
rect 47765 47613 47823 47647
rect 47765 47579 47777 47613
rect 47811 47579 47823 47613
rect 47765 47545 47823 47579
rect 47765 47511 47777 47545
rect 47811 47511 47823 47545
rect 47765 47477 47823 47511
rect 47765 47443 47777 47477
rect 47811 47443 47823 47477
rect 47765 47427 47823 47443
rect 48223 48701 48281 48717
rect 48223 48667 48235 48701
rect 48269 48667 48281 48701
rect 48223 48633 48281 48667
rect 48223 48599 48235 48633
rect 48269 48599 48281 48633
rect 48223 48565 48281 48599
rect 48223 48531 48235 48565
rect 48269 48531 48281 48565
rect 48223 48497 48281 48531
rect 48223 48463 48235 48497
rect 48269 48463 48281 48497
rect 48223 48429 48281 48463
rect 48223 48395 48235 48429
rect 48269 48395 48281 48429
rect 48223 48361 48281 48395
rect 48223 48327 48235 48361
rect 48269 48327 48281 48361
rect 48223 48293 48281 48327
rect 48223 48259 48235 48293
rect 48269 48259 48281 48293
rect 48223 48225 48281 48259
rect 48223 48191 48235 48225
rect 48269 48191 48281 48225
rect 48223 48157 48281 48191
rect 48223 48123 48235 48157
rect 48269 48123 48281 48157
rect 48223 48089 48281 48123
rect 48223 48055 48235 48089
rect 48269 48055 48281 48089
rect 48223 48021 48281 48055
rect 48223 47987 48235 48021
rect 48269 47987 48281 48021
rect 48223 47953 48281 47987
rect 48223 47919 48235 47953
rect 48269 47919 48281 47953
rect 48223 47885 48281 47919
rect 48223 47851 48235 47885
rect 48269 47851 48281 47885
rect 48223 47817 48281 47851
rect 48223 47783 48235 47817
rect 48269 47783 48281 47817
rect 48223 47749 48281 47783
rect 48223 47715 48235 47749
rect 48269 47715 48281 47749
rect 48223 47681 48281 47715
rect 48223 47647 48235 47681
rect 48269 47647 48281 47681
rect 48223 47613 48281 47647
rect 48223 47579 48235 47613
rect 48269 47579 48281 47613
rect 48223 47545 48281 47579
rect 48223 47511 48235 47545
rect 48269 47511 48281 47545
rect 48223 47477 48281 47511
rect 48223 47443 48235 47477
rect 48269 47443 48281 47477
rect 48223 47427 48281 47443
rect 48681 48701 48739 48717
rect 48681 48667 48693 48701
rect 48727 48667 48739 48701
rect 48681 48633 48739 48667
rect 48681 48599 48693 48633
rect 48727 48599 48739 48633
rect 48681 48565 48739 48599
rect 48681 48531 48693 48565
rect 48727 48531 48739 48565
rect 48681 48497 48739 48531
rect 48681 48463 48693 48497
rect 48727 48463 48739 48497
rect 48681 48429 48739 48463
rect 48681 48395 48693 48429
rect 48727 48395 48739 48429
rect 48681 48361 48739 48395
rect 48681 48327 48693 48361
rect 48727 48327 48739 48361
rect 48681 48293 48739 48327
rect 48681 48259 48693 48293
rect 48727 48259 48739 48293
rect 48681 48225 48739 48259
rect 48681 48191 48693 48225
rect 48727 48191 48739 48225
rect 48681 48157 48739 48191
rect 48681 48123 48693 48157
rect 48727 48123 48739 48157
rect 48681 48089 48739 48123
rect 48681 48055 48693 48089
rect 48727 48055 48739 48089
rect 48681 48021 48739 48055
rect 48681 47987 48693 48021
rect 48727 47987 48739 48021
rect 48681 47953 48739 47987
rect 48681 47919 48693 47953
rect 48727 47919 48739 47953
rect 48681 47885 48739 47919
rect 48681 47851 48693 47885
rect 48727 47851 48739 47885
rect 48681 47817 48739 47851
rect 48681 47783 48693 47817
rect 48727 47783 48739 47817
rect 48681 47749 48739 47783
rect 48681 47715 48693 47749
rect 48727 47715 48739 47749
rect 48681 47681 48739 47715
rect 48681 47647 48693 47681
rect 48727 47647 48739 47681
rect 48681 47613 48739 47647
rect 48681 47579 48693 47613
rect 48727 47579 48739 47613
rect 48681 47545 48739 47579
rect 48681 47511 48693 47545
rect 48727 47511 48739 47545
rect 48681 47477 48739 47511
rect 48681 47443 48693 47477
rect 48727 47443 48739 47477
rect 48681 47427 48739 47443
rect 49139 48701 49197 48717
rect 49139 48667 49151 48701
rect 49185 48667 49197 48701
rect 49139 48633 49197 48667
rect 49139 48599 49151 48633
rect 49185 48599 49197 48633
rect 49139 48565 49197 48599
rect 49139 48531 49151 48565
rect 49185 48531 49197 48565
rect 49139 48497 49197 48531
rect 49139 48463 49151 48497
rect 49185 48463 49197 48497
rect 49139 48429 49197 48463
rect 49139 48395 49151 48429
rect 49185 48395 49197 48429
rect 49139 48361 49197 48395
rect 49139 48327 49151 48361
rect 49185 48327 49197 48361
rect 49139 48293 49197 48327
rect 49139 48259 49151 48293
rect 49185 48259 49197 48293
rect 49139 48225 49197 48259
rect 49139 48191 49151 48225
rect 49185 48191 49197 48225
rect 49139 48157 49197 48191
rect 49139 48123 49151 48157
rect 49185 48123 49197 48157
rect 49139 48089 49197 48123
rect 49139 48055 49151 48089
rect 49185 48055 49197 48089
rect 49139 48021 49197 48055
rect 49139 47987 49151 48021
rect 49185 47987 49197 48021
rect 49139 47953 49197 47987
rect 49139 47919 49151 47953
rect 49185 47919 49197 47953
rect 49139 47885 49197 47919
rect 49139 47851 49151 47885
rect 49185 47851 49197 47885
rect 49139 47817 49197 47851
rect 49139 47783 49151 47817
rect 49185 47783 49197 47817
rect 49139 47749 49197 47783
rect 49139 47715 49151 47749
rect 49185 47715 49197 47749
rect 49139 47681 49197 47715
rect 49139 47647 49151 47681
rect 49185 47647 49197 47681
rect 49139 47613 49197 47647
rect 49139 47579 49151 47613
rect 49185 47579 49197 47613
rect 49139 47545 49197 47579
rect 49139 47511 49151 47545
rect 49185 47511 49197 47545
rect 49139 47477 49197 47511
rect 49139 47443 49151 47477
rect 49185 47443 49197 47477
rect 49139 47427 49197 47443
rect 49597 48701 49655 48717
rect 49597 48667 49609 48701
rect 49643 48667 49655 48701
rect 49597 48633 49655 48667
rect 49597 48599 49609 48633
rect 49643 48599 49655 48633
rect 49597 48565 49655 48599
rect 49597 48531 49609 48565
rect 49643 48531 49655 48565
rect 49597 48497 49655 48531
rect 49597 48463 49609 48497
rect 49643 48463 49655 48497
rect 49597 48429 49655 48463
rect 49597 48395 49609 48429
rect 49643 48395 49655 48429
rect 49597 48361 49655 48395
rect 49597 48327 49609 48361
rect 49643 48327 49655 48361
rect 49597 48293 49655 48327
rect 49597 48259 49609 48293
rect 49643 48259 49655 48293
rect 49597 48225 49655 48259
rect 49597 48191 49609 48225
rect 49643 48191 49655 48225
rect 49597 48157 49655 48191
rect 49597 48123 49609 48157
rect 49643 48123 49655 48157
rect 49597 48089 49655 48123
rect 49597 48055 49609 48089
rect 49643 48055 49655 48089
rect 49597 48021 49655 48055
rect 49597 47987 49609 48021
rect 49643 47987 49655 48021
rect 49597 47953 49655 47987
rect 49597 47919 49609 47953
rect 49643 47919 49655 47953
rect 49597 47885 49655 47919
rect 49597 47851 49609 47885
rect 49643 47851 49655 47885
rect 49597 47817 49655 47851
rect 49597 47783 49609 47817
rect 49643 47783 49655 47817
rect 49597 47749 49655 47783
rect 49597 47715 49609 47749
rect 49643 47715 49655 47749
rect 49597 47681 49655 47715
rect 49597 47647 49609 47681
rect 49643 47647 49655 47681
rect 49597 47613 49655 47647
rect 49597 47579 49609 47613
rect 49643 47579 49655 47613
rect 49597 47545 49655 47579
rect 49597 47511 49609 47545
rect 49643 47511 49655 47545
rect 49597 47477 49655 47511
rect 49597 47443 49609 47477
rect 49643 47443 49655 47477
rect 49597 47427 49655 47443
rect 50055 48701 50113 48717
rect 50055 48667 50067 48701
rect 50101 48667 50113 48701
rect 50055 48633 50113 48667
rect 50055 48599 50067 48633
rect 50101 48599 50113 48633
rect 50055 48565 50113 48599
rect 50055 48531 50067 48565
rect 50101 48531 50113 48565
rect 50055 48497 50113 48531
rect 50055 48463 50067 48497
rect 50101 48463 50113 48497
rect 50055 48429 50113 48463
rect 50055 48395 50067 48429
rect 50101 48395 50113 48429
rect 50055 48361 50113 48395
rect 50055 48327 50067 48361
rect 50101 48327 50113 48361
rect 50055 48293 50113 48327
rect 50055 48259 50067 48293
rect 50101 48259 50113 48293
rect 50055 48225 50113 48259
rect 50055 48191 50067 48225
rect 50101 48191 50113 48225
rect 50055 48157 50113 48191
rect 50055 48123 50067 48157
rect 50101 48123 50113 48157
rect 50055 48089 50113 48123
rect 50055 48055 50067 48089
rect 50101 48055 50113 48089
rect 50055 48021 50113 48055
rect 50055 47987 50067 48021
rect 50101 47987 50113 48021
rect 50055 47953 50113 47987
rect 50055 47919 50067 47953
rect 50101 47919 50113 47953
rect 50055 47885 50113 47919
rect 50055 47851 50067 47885
rect 50101 47851 50113 47885
rect 50055 47817 50113 47851
rect 50055 47783 50067 47817
rect 50101 47783 50113 47817
rect 50055 47749 50113 47783
rect 50055 47715 50067 47749
rect 50101 47715 50113 47749
rect 50055 47681 50113 47715
rect 50055 47647 50067 47681
rect 50101 47647 50113 47681
rect 50055 47613 50113 47647
rect 50055 47579 50067 47613
rect 50101 47579 50113 47613
rect 50055 47545 50113 47579
rect 50055 47511 50067 47545
rect 50101 47511 50113 47545
rect 50055 47477 50113 47511
rect 50055 47443 50067 47477
rect 50101 47443 50113 47477
rect 50055 47427 50113 47443
rect 50513 48701 50571 48717
rect 50513 48667 50525 48701
rect 50559 48667 50571 48701
rect 50513 48633 50571 48667
rect 50513 48599 50525 48633
rect 50559 48599 50571 48633
rect 50513 48565 50571 48599
rect 50513 48531 50525 48565
rect 50559 48531 50571 48565
rect 50513 48497 50571 48531
rect 50513 48463 50525 48497
rect 50559 48463 50571 48497
rect 50513 48429 50571 48463
rect 50513 48395 50525 48429
rect 50559 48395 50571 48429
rect 50513 48361 50571 48395
rect 50513 48327 50525 48361
rect 50559 48327 50571 48361
rect 50513 48293 50571 48327
rect 50513 48259 50525 48293
rect 50559 48259 50571 48293
rect 50513 48225 50571 48259
rect 50513 48191 50525 48225
rect 50559 48191 50571 48225
rect 50513 48157 50571 48191
rect 50513 48123 50525 48157
rect 50559 48123 50571 48157
rect 50513 48089 50571 48123
rect 50513 48055 50525 48089
rect 50559 48055 50571 48089
rect 50513 48021 50571 48055
rect 50513 47987 50525 48021
rect 50559 47987 50571 48021
rect 50513 47953 50571 47987
rect 50513 47919 50525 47953
rect 50559 47919 50571 47953
rect 50513 47885 50571 47919
rect 50513 47851 50525 47885
rect 50559 47851 50571 47885
rect 50513 47817 50571 47851
rect 50513 47783 50525 47817
rect 50559 47783 50571 47817
rect 50513 47749 50571 47783
rect 50513 47715 50525 47749
rect 50559 47715 50571 47749
rect 50513 47681 50571 47715
rect 50513 47647 50525 47681
rect 50559 47647 50571 47681
rect 50513 47613 50571 47647
rect 50513 47579 50525 47613
rect 50559 47579 50571 47613
rect 50513 47545 50571 47579
rect 50513 47511 50525 47545
rect 50559 47511 50571 47545
rect 50513 47477 50571 47511
rect 50513 47443 50525 47477
rect 50559 47443 50571 47477
rect 50513 47427 50571 47443
rect 50971 48701 51029 48717
rect 50971 48667 50983 48701
rect 51017 48667 51029 48701
rect 50971 48633 51029 48667
rect 50971 48599 50983 48633
rect 51017 48599 51029 48633
rect 50971 48565 51029 48599
rect 50971 48531 50983 48565
rect 51017 48531 51029 48565
rect 50971 48497 51029 48531
rect 50971 48463 50983 48497
rect 51017 48463 51029 48497
rect 50971 48429 51029 48463
rect 50971 48395 50983 48429
rect 51017 48395 51029 48429
rect 50971 48361 51029 48395
rect 50971 48327 50983 48361
rect 51017 48327 51029 48361
rect 50971 48293 51029 48327
rect 50971 48259 50983 48293
rect 51017 48259 51029 48293
rect 50971 48225 51029 48259
rect 50971 48191 50983 48225
rect 51017 48191 51029 48225
rect 50971 48157 51029 48191
rect 50971 48123 50983 48157
rect 51017 48123 51029 48157
rect 50971 48089 51029 48123
rect 50971 48055 50983 48089
rect 51017 48055 51029 48089
rect 50971 48021 51029 48055
rect 50971 47987 50983 48021
rect 51017 47987 51029 48021
rect 50971 47953 51029 47987
rect 50971 47919 50983 47953
rect 51017 47919 51029 47953
rect 50971 47885 51029 47919
rect 50971 47851 50983 47885
rect 51017 47851 51029 47885
rect 50971 47817 51029 47851
rect 50971 47783 50983 47817
rect 51017 47783 51029 47817
rect 50971 47749 51029 47783
rect 50971 47715 50983 47749
rect 51017 47715 51029 47749
rect 50971 47681 51029 47715
rect 50971 47647 50983 47681
rect 51017 47647 51029 47681
rect 50971 47613 51029 47647
rect 50971 47579 50983 47613
rect 51017 47579 51029 47613
rect 50971 47545 51029 47579
rect 50971 47511 50983 47545
rect 51017 47511 51029 47545
rect 50971 47477 51029 47511
rect 50971 47443 50983 47477
rect 51017 47443 51029 47477
rect 50971 47427 51029 47443
rect 51429 48701 51487 48717
rect 51429 48667 51441 48701
rect 51475 48667 51487 48701
rect 51429 48633 51487 48667
rect 51429 48599 51441 48633
rect 51475 48599 51487 48633
rect 51429 48565 51487 48599
rect 51429 48531 51441 48565
rect 51475 48531 51487 48565
rect 51429 48497 51487 48531
rect 51429 48463 51441 48497
rect 51475 48463 51487 48497
rect 51429 48429 51487 48463
rect 51429 48395 51441 48429
rect 51475 48395 51487 48429
rect 51429 48361 51487 48395
rect 51429 48327 51441 48361
rect 51475 48327 51487 48361
rect 51429 48293 51487 48327
rect 51429 48259 51441 48293
rect 51475 48259 51487 48293
rect 51429 48225 51487 48259
rect 51429 48191 51441 48225
rect 51475 48191 51487 48225
rect 51429 48157 51487 48191
rect 51429 48123 51441 48157
rect 51475 48123 51487 48157
rect 51429 48089 51487 48123
rect 51429 48055 51441 48089
rect 51475 48055 51487 48089
rect 51429 48021 51487 48055
rect 51429 47987 51441 48021
rect 51475 47987 51487 48021
rect 51429 47953 51487 47987
rect 51429 47919 51441 47953
rect 51475 47919 51487 47953
rect 51429 47885 51487 47919
rect 51429 47851 51441 47885
rect 51475 47851 51487 47885
rect 51429 47817 51487 47851
rect 51429 47783 51441 47817
rect 51475 47783 51487 47817
rect 51429 47749 51487 47783
rect 51429 47715 51441 47749
rect 51475 47715 51487 47749
rect 51429 47681 51487 47715
rect 51429 47647 51441 47681
rect 51475 47647 51487 47681
rect 51429 47613 51487 47647
rect 51429 47579 51441 47613
rect 51475 47579 51487 47613
rect 51429 47545 51487 47579
rect 51429 47511 51441 47545
rect 51475 47511 51487 47545
rect 51429 47477 51487 47511
rect 51429 47443 51441 47477
rect 51475 47443 51487 47477
rect 51429 47427 51487 47443
rect 51887 48701 51945 48717
rect 51887 48667 51899 48701
rect 51933 48667 51945 48701
rect 51887 48633 51945 48667
rect 51887 48599 51899 48633
rect 51933 48599 51945 48633
rect 51887 48565 51945 48599
rect 51887 48531 51899 48565
rect 51933 48531 51945 48565
rect 51887 48497 51945 48531
rect 51887 48463 51899 48497
rect 51933 48463 51945 48497
rect 51887 48429 51945 48463
rect 51887 48395 51899 48429
rect 51933 48395 51945 48429
rect 51887 48361 51945 48395
rect 51887 48327 51899 48361
rect 51933 48327 51945 48361
rect 51887 48293 51945 48327
rect 51887 48259 51899 48293
rect 51933 48259 51945 48293
rect 51887 48225 51945 48259
rect 51887 48191 51899 48225
rect 51933 48191 51945 48225
rect 51887 48157 51945 48191
rect 51887 48123 51899 48157
rect 51933 48123 51945 48157
rect 51887 48089 51945 48123
rect 51887 48055 51899 48089
rect 51933 48055 51945 48089
rect 51887 48021 51945 48055
rect 51887 47987 51899 48021
rect 51933 47987 51945 48021
rect 51887 47953 51945 47987
rect 51887 47919 51899 47953
rect 51933 47919 51945 47953
rect 51887 47885 51945 47919
rect 51887 47851 51899 47885
rect 51933 47851 51945 47885
rect 51887 47817 51945 47851
rect 51887 47783 51899 47817
rect 51933 47783 51945 47817
rect 51887 47749 51945 47783
rect 51887 47715 51899 47749
rect 51933 47715 51945 47749
rect 51887 47681 51945 47715
rect 51887 47647 51899 47681
rect 51933 47647 51945 47681
rect 51887 47613 51945 47647
rect 51887 47579 51899 47613
rect 51933 47579 51945 47613
rect 51887 47545 51945 47579
rect 51887 47511 51899 47545
rect 51933 47511 51945 47545
rect 51887 47477 51945 47511
rect 51887 47443 51899 47477
rect 51933 47443 51945 47477
rect 51887 47427 51945 47443
rect 52345 48701 52403 48717
rect 52345 48667 52357 48701
rect 52391 48667 52403 48701
rect 52345 48633 52403 48667
rect 52345 48599 52357 48633
rect 52391 48599 52403 48633
rect 52345 48565 52403 48599
rect 52345 48531 52357 48565
rect 52391 48531 52403 48565
rect 52345 48497 52403 48531
rect 52345 48463 52357 48497
rect 52391 48463 52403 48497
rect 52345 48429 52403 48463
rect 52345 48395 52357 48429
rect 52391 48395 52403 48429
rect 52345 48361 52403 48395
rect 52345 48327 52357 48361
rect 52391 48327 52403 48361
rect 52345 48293 52403 48327
rect 52345 48259 52357 48293
rect 52391 48259 52403 48293
rect 52345 48225 52403 48259
rect 52345 48191 52357 48225
rect 52391 48191 52403 48225
rect 52345 48157 52403 48191
rect 52345 48123 52357 48157
rect 52391 48123 52403 48157
rect 52345 48089 52403 48123
rect 52345 48055 52357 48089
rect 52391 48055 52403 48089
rect 52345 48021 52403 48055
rect 52345 47987 52357 48021
rect 52391 47987 52403 48021
rect 52345 47953 52403 47987
rect 52345 47919 52357 47953
rect 52391 47919 52403 47953
rect 52345 47885 52403 47919
rect 52345 47851 52357 47885
rect 52391 47851 52403 47885
rect 52345 47817 52403 47851
rect 52345 47783 52357 47817
rect 52391 47783 52403 47817
rect 52345 47749 52403 47783
rect 52345 47715 52357 47749
rect 52391 47715 52403 47749
rect 52345 47681 52403 47715
rect 52345 47647 52357 47681
rect 52391 47647 52403 47681
rect 52345 47613 52403 47647
rect 52345 47579 52357 47613
rect 52391 47579 52403 47613
rect 52345 47545 52403 47579
rect 52345 47511 52357 47545
rect 52391 47511 52403 47545
rect 52345 47477 52403 47511
rect 52345 47443 52357 47477
rect 52391 47443 52403 47477
rect 52345 47427 52403 47443
rect 15065 44941 15123 44957
rect 15065 44907 15077 44941
rect 15111 44907 15123 44941
rect 15065 44873 15123 44907
rect 15065 44839 15077 44873
rect 15111 44839 15123 44873
rect 15065 44805 15123 44839
rect 15065 44771 15077 44805
rect 15111 44771 15123 44805
rect 15065 44737 15123 44771
rect 15065 44703 15077 44737
rect 15111 44703 15123 44737
rect 15065 44669 15123 44703
rect 15065 44635 15077 44669
rect 15111 44635 15123 44669
rect 15065 44601 15123 44635
rect 15065 44567 15077 44601
rect 15111 44567 15123 44601
rect 15065 44533 15123 44567
rect 15065 44499 15077 44533
rect 15111 44499 15123 44533
rect 15065 44465 15123 44499
rect 15065 44431 15077 44465
rect 15111 44431 15123 44465
rect 15065 44397 15123 44431
rect 15065 44363 15077 44397
rect 15111 44363 15123 44397
rect 15065 44329 15123 44363
rect 15065 44295 15077 44329
rect 15111 44295 15123 44329
rect 15065 44261 15123 44295
rect 15065 44227 15077 44261
rect 15111 44227 15123 44261
rect 15065 44193 15123 44227
rect 15065 44159 15077 44193
rect 15111 44159 15123 44193
rect 15065 44125 15123 44159
rect 15065 44091 15077 44125
rect 15111 44091 15123 44125
rect 15065 44057 15123 44091
rect 15065 44023 15077 44057
rect 15111 44023 15123 44057
rect 15065 43989 15123 44023
rect 15065 43955 15077 43989
rect 15111 43955 15123 43989
rect 15065 43921 15123 43955
rect 15065 43887 15077 43921
rect 15111 43887 15123 43921
rect 15065 43853 15123 43887
rect 15065 43819 15077 43853
rect 15111 43819 15123 43853
rect 15065 43785 15123 43819
rect 15065 43751 15077 43785
rect 15111 43751 15123 43785
rect 15065 43717 15123 43751
rect 15065 43683 15077 43717
rect 15111 43683 15123 43717
rect 15065 43667 15123 43683
rect 15523 44941 15581 44957
rect 15523 44907 15535 44941
rect 15569 44907 15581 44941
rect 15523 44873 15581 44907
rect 15523 44839 15535 44873
rect 15569 44839 15581 44873
rect 15523 44805 15581 44839
rect 15523 44771 15535 44805
rect 15569 44771 15581 44805
rect 15523 44737 15581 44771
rect 15523 44703 15535 44737
rect 15569 44703 15581 44737
rect 15523 44669 15581 44703
rect 15523 44635 15535 44669
rect 15569 44635 15581 44669
rect 15523 44601 15581 44635
rect 15523 44567 15535 44601
rect 15569 44567 15581 44601
rect 15523 44533 15581 44567
rect 15523 44499 15535 44533
rect 15569 44499 15581 44533
rect 15523 44465 15581 44499
rect 15523 44431 15535 44465
rect 15569 44431 15581 44465
rect 15523 44397 15581 44431
rect 15523 44363 15535 44397
rect 15569 44363 15581 44397
rect 15523 44329 15581 44363
rect 15523 44295 15535 44329
rect 15569 44295 15581 44329
rect 15523 44261 15581 44295
rect 15523 44227 15535 44261
rect 15569 44227 15581 44261
rect 15523 44193 15581 44227
rect 15523 44159 15535 44193
rect 15569 44159 15581 44193
rect 15523 44125 15581 44159
rect 15523 44091 15535 44125
rect 15569 44091 15581 44125
rect 15523 44057 15581 44091
rect 15523 44023 15535 44057
rect 15569 44023 15581 44057
rect 15523 43989 15581 44023
rect 15523 43955 15535 43989
rect 15569 43955 15581 43989
rect 15523 43921 15581 43955
rect 15523 43887 15535 43921
rect 15569 43887 15581 43921
rect 15523 43853 15581 43887
rect 15523 43819 15535 43853
rect 15569 43819 15581 43853
rect 15523 43785 15581 43819
rect 15523 43751 15535 43785
rect 15569 43751 15581 43785
rect 15523 43717 15581 43751
rect 15523 43683 15535 43717
rect 15569 43683 15581 43717
rect 15523 43667 15581 43683
rect 15981 44941 16039 44957
rect 15981 44907 15993 44941
rect 16027 44907 16039 44941
rect 15981 44873 16039 44907
rect 15981 44839 15993 44873
rect 16027 44839 16039 44873
rect 15981 44805 16039 44839
rect 15981 44771 15993 44805
rect 16027 44771 16039 44805
rect 15981 44737 16039 44771
rect 15981 44703 15993 44737
rect 16027 44703 16039 44737
rect 15981 44669 16039 44703
rect 15981 44635 15993 44669
rect 16027 44635 16039 44669
rect 15981 44601 16039 44635
rect 15981 44567 15993 44601
rect 16027 44567 16039 44601
rect 15981 44533 16039 44567
rect 15981 44499 15993 44533
rect 16027 44499 16039 44533
rect 15981 44465 16039 44499
rect 15981 44431 15993 44465
rect 16027 44431 16039 44465
rect 15981 44397 16039 44431
rect 15981 44363 15993 44397
rect 16027 44363 16039 44397
rect 15981 44329 16039 44363
rect 15981 44295 15993 44329
rect 16027 44295 16039 44329
rect 15981 44261 16039 44295
rect 15981 44227 15993 44261
rect 16027 44227 16039 44261
rect 15981 44193 16039 44227
rect 15981 44159 15993 44193
rect 16027 44159 16039 44193
rect 15981 44125 16039 44159
rect 15981 44091 15993 44125
rect 16027 44091 16039 44125
rect 15981 44057 16039 44091
rect 15981 44023 15993 44057
rect 16027 44023 16039 44057
rect 15981 43989 16039 44023
rect 15981 43955 15993 43989
rect 16027 43955 16039 43989
rect 15981 43921 16039 43955
rect 15981 43887 15993 43921
rect 16027 43887 16039 43921
rect 15981 43853 16039 43887
rect 15981 43819 15993 43853
rect 16027 43819 16039 43853
rect 15981 43785 16039 43819
rect 15981 43751 15993 43785
rect 16027 43751 16039 43785
rect 15981 43717 16039 43751
rect 15981 43683 15993 43717
rect 16027 43683 16039 43717
rect 15981 43667 16039 43683
rect 16439 44941 16497 44957
rect 16439 44907 16451 44941
rect 16485 44907 16497 44941
rect 16439 44873 16497 44907
rect 16439 44839 16451 44873
rect 16485 44839 16497 44873
rect 16439 44805 16497 44839
rect 16439 44771 16451 44805
rect 16485 44771 16497 44805
rect 16439 44737 16497 44771
rect 16439 44703 16451 44737
rect 16485 44703 16497 44737
rect 16439 44669 16497 44703
rect 16439 44635 16451 44669
rect 16485 44635 16497 44669
rect 16439 44601 16497 44635
rect 16439 44567 16451 44601
rect 16485 44567 16497 44601
rect 16439 44533 16497 44567
rect 16439 44499 16451 44533
rect 16485 44499 16497 44533
rect 16439 44465 16497 44499
rect 16439 44431 16451 44465
rect 16485 44431 16497 44465
rect 16439 44397 16497 44431
rect 16439 44363 16451 44397
rect 16485 44363 16497 44397
rect 16439 44329 16497 44363
rect 16439 44295 16451 44329
rect 16485 44295 16497 44329
rect 16439 44261 16497 44295
rect 16439 44227 16451 44261
rect 16485 44227 16497 44261
rect 16439 44193 16497 44227
rect 16439 44159 16451 44193
rect 16485 44159 16497 44193
rect 16439 44125 16497 44159
rect 16439 44091 16451 44125
rect 16485 44091 16497 44125
rect 16439 44057 16497 44091
rect 16439 44023 16451 44057
rect 16485 44023 16497 44057
rect 16439 43989 16497 44023
rect 16439 43955 16451 43989
rect 16485 43955 16497 43989
rect 16439 43921 16497 43955
rect 16439 43887 16451 43921
rect 16485 43887 16497 43921
rect 16439 43853 16497 43887
rect 16439 43819 16451 43853
rect 16485 43819 16497 43853
rect 16439 43785 16497 43819
rect 16439 43751 16451 43785
rect 16485 43751 16497 43785
rect 16439 43717 16497 43751
rect 16439 43683 16451 43717
rect 16485 43683 16497 43717
rect 16439 43667 16497 43683
rect 16897 44941 16955 44957
rect 16897 44907 16909 44941
rect 16943 44907 16955 44941
rect 16897 44873 16955 44907
rect 16897 44839 16909 44873
rect 16943 44839 16955 44873
rect 16897 44805 16955 44839
rect 16897 44771 16909 44805
rect 16943 44771 16955 44805
rect 16897 44737 16955 44771
rect 16897 44703 16909 44737
rect 16943 44703 16955 44737
rect 16897 44669 16955 44703
rect 16897 44635 16909 44669
rect 16943 44635 16955 44669
rect 16897 44601 16955 44635
rect 16897 44567 16909 44601
rect 16943 44567 16955 44601
rect 16897 44533 16955 44567
rect 16897 44499 16909 44533
rect 16943 44499 16955 44533
rect 16897 44465 16955 44499
rect 16897 44431 16909 44465
rect 16943 44431 16955 44465
rect 16897 44397 16955 44431
rect 16897 44363 16909 44397
rect 16943 44363 16955 44397
rect 16897 44329 16955 44363
rect 16897 44295 16909 44329
rect 16943 44295 16955 44329
rect 16897 44261 16955 44295
rect 16897 44227 16909 44261
rect 16943 44227 16955 44261
rect 16897 44193 16955 44227
rect 16897 44159 16909 44193
rect 16943 44159 16955 44193
rect 16897 44125 16955 44159
rect 16897 44091 16909 44125
rect 16943 44091 16955 44125
rect 16897 44057 16955 44091
rect 16897 44023 16909 44057
rect 16943 44023 16955 44057
rect 16897 43989 16955 44023
rect 16897 43955 16909 43989
rect 16943 43955 16955 43989
rect 16897 43921 16955 43955
rect 16897 43887 16909 43921
rect 16943 43887 16955 43921
rect 16897 43853 16955 43887
rect 16897 43819 16909 43853
rect 16943 43819 16955 43853
rect 16897 43785 16955 43819
rect 16897 43751 16909 43785
rect 16943 43751 16955 43785
rect 16897 43717 16955 43751
rect 16897 43683 16909 43717
rect 16943 43683 16955 43717
rect 16897 43667 16955 43683
rect 17355 44941 17413 44957
rect 17355 44907 17367 44941
rect 17401 44907 17413 44941
rect 17355 44873 17413 44907
rect 17355 44839 17367 44873
rect 17401 44839 17413 44873
rect 17355 44805 17413 44839
rect 17355 44771 17367 44805
rect 17401 44771 17413 44805
rect 17355 44737 17413 44771
rect 17355 44703 17367 44737
rect 17401 44703 17413 44737
rect 17355 44669 17413 44703
rect 17355 44635 17367 44669
rect 17401 44635 17413 44669
rect 17355 44601 17413 44635
rect 17355 44567 17367 44601
rect 17401 44567 17413 44601
rect 17355 44533 17413 44567
rect 17355 44499 17367 44533
rect 17401 44499 17413 44533
rect 17355 44465 17413 44499
rect 17355 44431 17367 44465
rect 17401 44431 17413 44465
rect 17355 44397 17413 44431
rect 17355 44363 17367 44397
rect 17401 44363 17413 44397
rect 17355 44329 17413 44363
rect 17355 44295 17367 44329
rect 17401 44295 17413 44329
rect 17355 44261 17413 44295
rect 17355 44227 17367 44261
rect 17401 44227 17413 44261
rect 17355 44193 17413 44227
rect 17355 44159 17367 44193
rect 17401 44159 17413 44193
rect 17355 44125 17413 44159
rect 17355 44091 17367 44125
rect 17401 44091 17413 44125
rect 17355 44057 17413 44091
rect 17355 44023 17367 44057
rect 17401 44023 17413 44057
rect 17355 43989 17413 44023
rect 17355 43955 17367 43989
rect 17401 43955 17413 43989
rect 17355 43921 17413 43955
rect 17355 43887 17367 43921
rect 17401 43887 17413 43921
rect 17355 43853 17413 43887
rect 17355 43819 17367 43853
rect 17401 43819 17413 43853
rect 17355 43785 17413 43819
rect 17355 43751 17367 43785
rect 17401 43751 17413 43785
rect 17355 43717 17413 43751
rect 17355 43683 17367 43717
rect 17401 43683 17413 43717
rect 17355 43667 17413 43683
rect 17813 44941 17871 44957
rect 17813 44907 17825 44941
rect 17859 44907 17871 44941
rect 17813 44873 17871 44907
rect 17813 44839 17825 44873
rect 17859 44839 17871 44873
rect 17813 44805 17871 44839
rect 17813 44771 17825 44805
rect 17859 44771 17871 44805
rect 17813 44737 17871 44771
rect 17813 44703 17825 44737
rect 17859 44703 17871 44737
rect 17813 44669 17871 44703
rect 17813 44635 17825 44669
rect 17859 44635 17871 44669
rect 17813 44601 17871 44635
rect 17813 44567 17825 44601
rect 17859 44567 17871 44601
rect 17813 44533 17871 44567
rect 17813 44499 17825 44533
rect 17859 44499 17871 44533
rect 17813 44465 17871 44499
rect 17813 44431 17825 44465
rect 17859 44431 17871 44465
rect 17813 44397 17871 44431
rect 17813 44363 17825 44397
rect 17859 44363 17871 44397
rect 17813 44329 17871 44363
rect 17813 44295 17825 44329
rect 17859 44295 17871 44329
rect 17813 44261 17871 44295
rect 17813 44227 17825 44261
rect 17859 44227 17871 44261
rect 17813 44193 17871 44227
rect 17813 44159 17825 44193
rect 17859 44159 17871 44193
rect 17813 44125 17871 44159
rect 17813 44091 17825 44125
rect 17859 44091 17871 44125
rect 17813 44057 17871 44091
rect 17813 44023 17825 44057
rect 17859 44023 17871 44057
rect 17813 43989 17871 44023
rect 17813 43955 17825 43989
rect 17859 43955 17871 43989
rect 17813 43921 17871 43955
rect 17813 43887 17825 43921
rect 17859 43887 17871 43921
rect 17813 43853 17871 43887
rect 17813 43819 17825 43853
rect 17859 43819 17871 43853
rect 17813 43785 17871 43819
rect 17813 43751 17825 43785
rect 17859 43751 17871 43785
rect 17813 43717 17871 43751
rect 17813 43683 17825 43717
rect 17859 43683 17871 43717
rect 17813 43667 17871 43683
rect 18271 44941 18329 44957
rect 18271 44907 18283 44941
rect 18317 44907 18329 44941
rect 18271 44873 18329 44907
rect 18271 44839 18283 44873
rect 18317 44839 18329 44873
rect 18271 44805 18329 44839
rect 18271 44771 18283 44805
rect 18317 44771 18329 44805
rect 18271 44737 18329 44771
rect 18271 44703 18283 44737
rect 18317 44703 18329 44737
rect 18271 44669 18329 44703
rect 18271 44635 18283 44669
rect 18317 44635 18329 44669
rect 18271 44601 18329 44635
rect 18271 44567 18283 44601
rect 18317 44567 18329 44601
rect 18271 44533 18329 44567
rect 18271 44499 18283 44533
rect 18317 44499 18329 44533
rect 18271 44465 18329 44499
rect 18271 44431 18283 44465
rect 18317 44431 18329 44465
rect 18271 44397 18329 44431
rect 18271 44363 18283 44397
rect 18317 44363 18329 44397
rect 18271 44329 18329 44363
rect 18271 44295 18283 44329
rect 18317 44295 18329 44329
rect 18271 44261 18329 44295
rect 18271 44227 18283 44261
rect 18317 44227 18329 44261
rect 18271 44193 18329 44227
rect 18271 44159 18283 44193
rect 18317 44159 18329 44193
rect 18271 44125 18329 44159
rect 18271 44091 18283 44125
rect 18317 44091 18329 44125
rect 18271 44057 18329 44091
rect 18271 44023 18283 44057
rect 18317 44023 18329 44057
rect 18271 43989 18329 44023
rect 18271 43955 18283 43989
rect 18317 43955 18329 43989
rect 18271 43921 18329 43955
rect 18271 43887 18283 43921
rect 18317 43887 18329 43921
rect 18271 43853 18329 43887
rect 18271 43819 18283 43853
rect 18317 43819 18329 43853
rect 18271 43785 18329 43819
rect 18271 43751 18283 43785
rect 18317 43751 18329 43785
rect 18271 43717 18329 43751
rect 18271 43683 18283 43717
rect 18317 43683 18329 43717
rect 18271 43667 18329 43683
rect 18729 44941 18787 44957
rect 18729 44907 18741 44941
rect 18775 44907 18787 44941
rect 18729 44873 18787 44907
rect 18729 44839 18741 44873
rect 18775 44839 18787 44873
rect 18729 44805 18787 44839
rect 18729 44771 18741 44805
rect 18775 44771 18787 44805
rect 18729 44737 18787 44771
rect 18729 44703 18741 44737
rect 18775 44703 18787 44737
rect 18729 44669 18787 44703
rect 18729 44635 18741 44669
rect 18775 44635 18787 44669
rect 18729 44601 18787 44635
rect 18729 44567 18741 44601
rect 18775 44567 18787 44601
rect 18729 44533 18787 44567
rect 18729 44499 18741 44533
rect 18775 44499 18787 44533
rect 18729 44465 18787 44499
rect 18729 44431 18741 44465
rect 18775 44431 18787 44465
rect 18729 44397 18787 44431
rect 18729 44363 18741 44397
rect 18775 44363 18787 44397
rect 18729 44329 18787 44363
rect 18729 44295 18741 44329
rect 18775 44295 18787 44329
rect 18729 44261 18787 44295
rect 18729 44227 18741 44261
rect 18775 44227 18787 44261
rect 18729 44193 18787 44227
rect 18729 44159 18741 44193
rect 18775 44159 18787 44193
rect 18729 44125 18787 44159
rect 18729 44091 18741 44125
rect 18775 44091 18787 44125
rect 18729 44057 18787 44091
rect 18729 44023 18741 44057
rect 18775 44023 18787 44057
rect 18729 43989 18787 44023
rect 18729 43955 18741 43989
rect 18775 43955 18787 43989
rect 18729 43921 18787 43955
rect 18729 43887 18741 43921
rect 18775 43887 18787 43921
rect 18729 43853 18787 43887
rect 18729 43819 18741 43853
rect 18775 43819 18787 43853
rect 18729 43785 18787 43819
rect 18729 43751 18741 43785
rect 18775 43751 18787 43785
rect 18729 43717 18787 43751
rect 18729 43683 18741 43717
rect 18775 43683 18787 43717
rect 18729 43667 18787 43683
rect 19187 44941 19245 44957
rect 19187 44907 19199 44941
rect 19233 44907 19245 44941
rect 19187 44873 19245 44907
rect 19187 44839 19199 44873
rect 19233 44839 19245 44873
rect 19187 44805 19245 44839
rect 19187 44771 19199 44805
rect 19233 44771 19245 44805
rect 19187 44737 19245 44771
rect 19187 44703 19199 44737
rect 19233 44703 19245 44737
rect 19187 44669 19245 44703
rect 19187 44635 19199 44669
rect 19233 44635 19245 44669
rect 19187 44601 19245 44635
rect 19187 44567 19199 44601
rect 19233 44567 19245 44601
rect 19187 44533 19245 44567
rect 19187 44499 19199 44533
rect 19233 44499 19245 44533
rect 19187 44465 19245 44499
rect 19187 44431 19199 44465
rect 19233 44431 19245 44465
rect 19187 44397 19245 44431
rect 19187 44363 19199 44397
rect 19233 44363 19245 44397
rect 19187 44329 19245 44363
rect 19187 44295 19199 44329
rect 19233 44295 19245 44329
rect 19187 44261 19245 44295
rect 19187 44227 19199 44261
rect 19233 44227 19245 44261
rect 19187 44193 19245 44227
rect 19187 44159 19199 44193
rect 19233 44159 19245 44193
rect 19187 44125 19245 44159
rect 19187 44091 19199 44125
rect 19233 44091 19245 44125
rect 19187 44057 19245 44091
rect 19187 44023 19199 44057
rect 19233 44023 19245 44057
rect 19187 43989 19245 44023
rect 19187 43955 19199 43989
rect 19233 43955 19245 43989
rect 19187 43921 19245 43955
rect 19187 43887 19199 43921
rect 19233 43887 19245 43921
rect 19187 43853 19245 43887
rect 19187 43819 19199 43853
rect 19233 43819 19245 43853
rect 19187 43785 19245 43819
rect 19187 43751 19199 43785
rect 19233 43751 19245 43785
rect 19187 43717 19245 43751
rect 19187 43683 19199 43717
rect 19233 43683 19245 43717
rect 19187 43667 19245 43683
rect 19645 44941 19703 44957
rect 19645 44907 19657 44941
rect 19691 44907 19703 44941
rect 19645 44873 19703 44907
rect 19645 44839 19657 44873
rect 19691 44839 19703 44873
rect 19645 44805 19703 44839
rect 19645 44771 19657 44805
rect 19691 44771 19703 44805
rect 19645 44737 19703 44771
rect 19645 44703 19657 44737
rect 19691 44703 19703 44737
rect 19645 44669 19703 44703
rect 19645 44635 19657 44669
rect 19691 44635 19703 44669
rect 19645 44601 19703 44635
rect 19645 44567 19657 44601
rect 19691 44567 19703 44601
rect 19645 44533 19703 44567
rect 19645 44499 19657 44533
rect 19691 44499 19703 44533
rect 19645 44465 19703 44499
rect 19645 44431 19657 44465
rect 19691 44431 19703 44465
rect 19645 44397 19703 44431
rect 19645 44363 19657 44397
rect 19691 44363 19703 44397
rect 19645 44329 19703 44363
rect 19645 44295 19657 44329
rect 19691 44295 19703 44329
rect 19645 44261 19703 44295
rect 19645 44227 19657 44261
rect 19691 44227 19703 44261
rect 19645 44193 19703 44227
rect 19645 44159 19657 44193
rect 19691 44159 19703 44193
rect 19645 44125 19703 44159
rect 19645 44091 19657 44125
rect 19691 44091 19703 44125
rect 19645 44057 19703 44091
rect 19645 44023 19657 44057
rect 19691 44023 19703 44057
rect 19645 43989 19703 44023
rect 19645 43955 19657 43989
rect 19691 43955 19703 43989
rect 19645 43921 19703 43955
rect 19645 43887 19657 43921
rect 19691 43887 19703 43921
rect 19645 43853 19703 43887
rect 19645 43819 19657 43853
rect 19691 43819 19703 43853
rect 19645 43785 19703 43819
rect 19645 43751 19657 43785
rect 19691 43751 19703 43785
rect 19645 43717 19703 43751
rect 19645 43683 19657 43717
rect 19691 43683 19703 43717
rect 19645 43667 19703 43683
rect 20103 44941 20161 44957
rect 20103 44907 20115 44941
rect 20149 44907 20161 44941
rect 20103 44873 20161 44907
rect 20103 44839 20115 44873
rect 20149 44839 20161 44873
rect 20103 44805 20161 44839
rect 20103 44771 20115 44805
rect 20149 44771 20161 44805
rect 20103 44737 20161 44771
rect 20103 44703 20115 44737
rect 20149 44703 20161 44737
rect 20103 44669 20161 44703
rect 20103 44635 20115 44669
rect 20149 44635 20161 44669
rect 20103 44601 20161 44635
rect 20103 44567 20115 44601
rect 20149 44567 20161 44601
rect 20103 44533 20161 44567
rect 20103 44499 20115 44533
rect 20149 44499 20161 44533
rect 20103 44465 20161 44499
rect 20103 44431 20115 44465
rect 20149 44431 20161 44465
rect 20103 44397 20161 44431
rect 20103 44363 20115 44397
rect 20149 44363 20161 44397
rect 20103 44329 20161 44363
rect 20103 44295 20115 44329
rect 20149 44295 20161 44329
rect 20103 44261 20161 44295
rect 20103 44227 20115 44261
rect 20149 44227 20161 44261
rect 20103 44193 20161 44227
rect 20103 44159 20115 44193
rect 20149 44159 20161 44193
rect 20103 44125 20161 44159
rect 20103 44091 20115 44125
rect 20149 44091 20161 44125
rect 20103 44057 20161 44091
rect 20103 44023 20115 44057
rect 20149 44023 20161 44057
rect 20103 43989 20161 44023
rect 20103 43955 20115 43989
rect 20149 43955 20161 43989
rect 20103 43921 20161 43955
rect 20103 43887 20115 43921
rect 20149 43887 20161 43921
rect 20103 43853 20161 43887
rect 20103 43819 20115 43853
rect 20149 43819 20161 43853
rect 20103 43785 20161 43819
rect 20103 43751 20115 43785
rect 20149 43751 20161 43785
rect 20103 43717 20161 43751
rect 20103 43683 20115 43717
rect 20149 43683 20161 43717
rect 20103 43667 20161 43683
rect 20561 44941 20619 44957
rect 20561 44907 20573 44941
rect 20607 44907 20619 44941
rect 20561 44873 20619 44907
rect 20561 44839 20573 44873
rect 20607 44839 20619 44873
rect 20561 44805 20619 44839
rect 20561 44771 20573 44805
rect 20607 44771 20619 44805
rect 20561 44737 20619 44771
rect 20561 44703 20573 44737
rect 20607 44703 20619 44737
rect 20561 44669 20619 44703
rect 20561 44635 20573 44669
rect 20607 44635 20619 44669
rect 20561 44601 20619 44635
rect 20561 44567 20573 44601
rect 20607 44567 20619 44601
rect 20561 44533 20619 44567
rect 20561 44499 20573 44533
rect 20607 44499 20619 44533
rect 20561 44465 20619 44499
rect 20561 44431 20573 44465
rect 20607 44431 20619 44465
rect 20561 44397 20619 44431
rect 20561 44363 20573 44397
rect 20607 44363 20619 44397
rect 20561 44329 20619 44363
rect 20561 44295 20573 44329
rect 20607 44295 20619 44329
rect 20561 44261 20619 44295
rect 20561 44227 20573 44261
rect 20607 44227 20619 44261
rect 20561 44193 20619 44227
rect 20561 44159 20573 44193
rect 20607 44159 20619 44193
rect 20561 44125 20619 44159
rect 20561 44091 20573 44125
rect 20607 44091 20619 44125
rect 20561 44057 20619 44091
rect 20561 44023 20573 44057
rect 20607 44023 20619 44057
rect 20561 43989 20619 44023
rect 20561 43955 20573 43989
rect 20607 43955 20619 43989
rect 20561 43921 20619 43955
rect 20561 43887 20573 43921
rect 20607 43887 20619 43921
rect 20561 43853 20619 43887
rect 20561 43819 20573 43853
rect 20607 43819 20619 43853
rect 20561 43785 20619 43819
rect 20561 43751 20573 43785
rect 20607 43751 20619 43785
rect 20561 43717 20619 43751
rect 20561 43683 20573 43717
rect 20607 43683 20619 43717
rect 20561 43667 20619 43683
rect 21019 44941 21077 44957
rect 21019 44907 21031 44941
rect 21065 44907 21077 44941
rect 21019 44873 21077 44907
rect 21019 44839 21031 44873
rect 21065 44839 21077 44873
rect 21019 44805 21077 44839
rect 21019 44771 21031 44805
rect 21065 44771 21077 44805
rect 21019 44737 21077 44771
rect 21019 44703 21031 44737
rect 21065 44703 21077 44737
rect 21019 44669 21077 44703
rect 21019 44635 21031 44669
rect 21065 44635 21077 44669
rect 21019 44601 21077 44635
rect 21019 44567 21031 44601
rect 21065 44567 21077 44601
rect 21019 44533 21077 44567
rect 21019 44499 21031 44533
rect 21065 44499 21077 44533
rect 21019 44465 21077 44499
rect 21019 44431 21031 44465
rect 21065 44431 21077 44465
rect 21019 44397 21077 44431
rect 21019 44363 21031 44397
rect 21065 44363 21077 44397
rect 21019 44329 21077 44363
rect 21019 44295 21031 44329
rect 21065 44295 21077 44329
rect 21019 44261 21077 44295
rect 21019 44227 21031 44261
rect 21065 44227 21077 44261
rect 21019 44193 21077 44227
rect 21019 44159 21031 44193
rect 21065 44159 21077 44193
rect 21019 44125 21077 44159
rect 21019 44091 21031 44125
rect 21065 44091 21077 44125
rect 21019 44057 21077 44091
rect 21019 44023 21031 44057
rect 21065 44023 21077 44057
rect 21019 43989 21077 44023
rect 21019 43955 21031 43989
rect 21065 43955 21077 43989
rect 21019 43921 21077 43955
rect 21019 43887 21031 43921
rect 21065 43887 21077 43921
rect 21019 43853 21077 43887
rect 21019 43819 21031 43853
rect 21065 43819 21077 43853
rect 21019 43785 21077 43819
rect 21019 43751 21031 43785
rect 21065 43751 21077 43785
rect 21019 43717 21077 43751
rect 21019 43683 21031 43717
rect 21065 43683 21077 43717
rect 21019 43667 21077 43683
rect 21477 44941 21535 44957
rect 21477 44907 21489 44941
rect 21523 44907 21535 44941
rect 21477 44873 21535 44907
rect 21477 44839 21489 44873
rect 21523 44839 21535 44873
rect 21477 44805 21535 44839
rect 21477 44771 21489 44805
rect 21523 44771 21535 44805
rect 21477 44737 21535 44771
rect 21477 44703 21489 44737
rect 21523 44703 21535 44737
rect 21477 44669 21535 44703
rect 21477 44635 21489 44669
rect 21523 44635 21535 44669
rect 21477 44601 21535 44635
rect 21477 44567 21489 44601
rect 21523 44567 21535 44601
rect 21477 44533 21535 44567
rect 21477 44499 21489 44533
rect 21523 44499 21535 44533
rect 21477 44465 21535 44499
rect 21477 44431 21489 44465
rect 21523 44431 21535 44465
rect 21477 44397 21535 44431
rect 21477 44363 21489 44397
rect 21523 44363 21535 44397
rect 21477 44329 21535 44363
rect 21477 44295 21489 44329
rect 21523 44295 21535 44329
rect 21477 44261 21535 44295
rect 21477 44227 21489 44261
rect 21523 44227 21535 44261
rect 21477 44193 21535 44227
rect 21477 44159 21489 44193
rect 21523 44159 21535 44193
rect 21477 44125 21535 44159
rect 21477 44091 21489 44125
rect 21523 44091 21535 44125
rect 21477 44057 21535 44091
rect 21477 44023 21489 44057
rect 21523 44023 21535 44057
rect 21477 43989 21535 44023
rect 21477 43955 21489 43989
rect 21523 43955 21535 43989
rect 21477 43921 21535 43955
rect 21477 43887 21489 43921
rect 21523 43887 21535 43921
rect 21477 43853 21535 43887
rect 21477 43819 21489 43853
rect 21523 43819 21535 43853
rect 21477 43785 21535 43819
rect 21477 43751 21489 43785
rect 21523 43751 21535 43785
rect 21477 43717 21535 43751
rect 21477 43683 21489 43717
rect 21523 43683 21535 43717
rect 21477 43667 21535 43683
rect 21935 44941 21993 44957
rect 21935 44907 21947 44941
rect 21981 44907 21993 44941
rect 21935 44873 21993 44907
rect 21935 44839 21947 44873
rect 21981 44839 21993 44873
rect 21935 44805 21993 44839
rect 21935 44771 21947 44805
rect 21981 44771 21993 44805
rect 21935 44737 21993 44771
rect 21935 44703 21947 44737
rect 21981 44703 21993 44737
rect 21935 44669 21993 44703
rect 21935 44635 21947 44669
rect 21981 44635 21993 44669
rect 21935 44601 21993 44635
rect 21935 44567 21947 44601
rect 21981 44567 21993 44601
rect 21935 44533 21993 44567
rect 21935 44499 21947 44533
rect 21981 44499 21993 44533
rect 21935 44465 21993 44499
rect 21935 44431 21947 44465
rect 21981 44431 21993 44465
rect 21935 44397 21993 44431
rect 21935 44363 21947 44397
rect 21981 44363 21993 44397
rect 21935 44329 21993 44363
rect 21935 44295 21947 44329
rect 21981 44295 21993 44329
rect 21935 44261 21993 44295
rect 21935 44227 21947 44261
rect 21981 44227 21993 44261
rect 21935 44193 21993 44227
rect 21935 44159 21947 44193
rect 21981 44159 21993 44193
rect 21935 44125 21993 44159
rect 21935 44091 21947 44125
rect 21981 44091 21993 44125
rect 21935 44057 21993 44091
rect 21935 44023 21947 44057
rect 21981 44023 21993 44057
rect 21935 43989 21993 44023
rect 21935 43955 21947 43989
rect 21981 43955 21993 43989
rect 21935 43921 21993 43955
rect 21935 43887 21947 43921
rect 21981 43887 21993 43921
rect 21935 43853 21993 43887
rect 21935 43819 21947 43853
rect 21981 43819 21993 43853
rect 21935 43785 21993 43819
rect 21935 43751 21947 43785
rect 21981 43751 21993 43785
rect 21935 43717 21993 43751
rect 21935 43683 21947 43717
rect 21981 43683 21993 43717
rect 21935 43667 21993 43683
rect 22393 44941 22451 44957
rect 22393 44907 22405 44941
rect 22439 44907 22451 44941
rect 22393 44873 22451 44907
rect 22393 44839 22405 44873
rect 22439 44839 22451 44873
rect 22393 44805 22451 44839
rect 22393 44771 22405 44805
rect 22439 44771 22451 44805
rect 22393 44737 22451 44771
rect 22393 44703 22405 44737
rect 22439 44703 22451 44737
rect 22393 44669 22451 44703
rect 22393 44635 22405 44669
rect 22439 44635 22451 44669
rect 22393 44601 22451 44635
rect 22393 44567 22405 44601
rect 22439 44567 22451 44601
rect 22393 44533 22451 44567
rect 22393 44499 22405 44533
rect 22439 44499 22451 44533
rect 22393 44465 22451 44499
rect 22393 44431 22405 44465
rect 22439 44431 22451 44465
rect 22393 44397 22451 44431
rect 22393 44363 22405 44397
rect 22439 44363 22451 44397
rect 22393 44329 22451 44363
rect 22393 44295 22405 44329
rect 22439 44295 22451 44329
rect 22393 44261 22451 44295
rect 22393 44227 22405 44261
rect 22439 44227 22451 44261
rect 22393 44193 22451 44227
rect 22393 44159 22405 44193
rect 22439 44159 22451 44193
rect 22393 44125 22451 44159
rect 22393 44091 22405 44125
rect 22439 44091 22451 44125
rect 22393 44057 22451 44091
rect 22393 44023 22405 44057
rect 22439 44023 22451 44057
rect 22393 43989 22451 44023
rect 22393 43955 22405 43989
rect 22439 43955 22451 43989
rect 22393 43921 22451 43955
rect 22393 43887 22405 43921
rect 22439 43887 22451 43921
rect 22393 43853 22451 43887
rect 22393 43819 22405 43853
rect 22439 43819 22451 43853
rect 22393 43785 22451 43819
rect 22393 43751 22405 43785
rect 22439 43751 22451 43785
rect 22393 43717 22451 43751
rect 22393 43683 22405 43717
rect 22439 43683 22451 43717
rect 22393 43667 22451 43683
rect 22851 44941 22909 44957
rect 22851 44907 22863 44941
rect 22897 44907 22909 44941
rect 22851 44873 22909 44907
rect 22851 44839 22863 44873
rect 22897 44839 22909 44873
rect 22851 44805 22909 44839
rect 22851 44771 22863 44805
rect 22897 44771 22909 44805
rect 22851 44737 22909 44771
rect 22851 44703 22863 44737
rect 22897 44703 22909 44737
rect 22851 44669 22909 44703
rect 22851 44635 22863 44669
rect 22897 44635 22909 44669
rect 22851 44601 22909 44635
rect 22851 44567 22863 44601
rect 22897 44567 22909 44601
rect 22851 44533 22909 44567
rect 22851 44499 22863 44533
rect 22897 44499 22909 44533
rect 22851 44465 22909 44499
rect 22851 44431 22863 44465
rect 22897 44431 22909 44465
rect 22851 44397 22909 44431
rect 22851 44363 22863 44397
rect 22897 44363 22909 44397
rect 22851 44329 22909 44363
rect 22851 44295 22863 44329
rect 22897 44295 22909 44329
rect 22851 44261 22909 44295
rect 22851 44227 22863 44261
rect 22897 44227 22909 44261
rect 22851 44193 22909 44227
rect 22851 44159 22863 44193
rect 22897 44159 22909 44193
rect 22851 44125 22909 44159
rect 22851 44091 22863 44125
rect 22897 44091 22909 44125
rect 22851 44057 22909 44091
rect 22851 44023 22863 44057
rect 22897 44023 22909 44057
rect 22851 43989 22909 44023
rect 22851 43955 22863 43989
rect 22897 43955 22909 43989
rect 22851 43921 22909 43955
rect 22851 43887 22863 43921
rect 22897 43887 22909 43921
rect 22851 43853 22909 43887
rect 22851 43819 22863 43853
rect 22897 43819 22909 43853
rect 22851 43785 22909 43819
rect 22851 43751 22863 43785
rect 22897 43751 22909 43785
rect 22851 43717 22909 43751
rect 22851 43683 22863 43717
rect 22897 43683 22909 43717
rect 22851 43667 22909 43683
rect 23309 44941 23367 44957
rect 23309 44907 23321 44941
rect 23355 44907 23367 44941
rect 23309 44873 23367 44907
rect 23309 44839 23321 44873
rect 23355 44839 23367 44873
rect 23309 44805 23367 44839
rect 23309 44771 23321 44805
rect 23355 44771 23367 44805
rect 23309 44737 23367 44771
rect 23309 44703 23321 44737
rect 23355 44703 23367 44737
rect 23309 44669 23367 44703
rect 23309 44635 23321 44669
rect 23355 44635 23367 44669
rect 23309 44601 23367 44635
rect 23309 44567 23321 44601
rect 23355 44567 23367 44601
rect 23309 44533 23367 44567
rect 23309 44499 23321 44533
rect 23355 44499 23367 44533
rect 23309 44465 23367 44499
rect 23309 44431 23321 44465
rect 23355 44431 23367 44465
rect 23309 44397 23367 44431
rect 23309 44363 23321 44397
rect 23355 44363 23367 44397
rect 23309 44329 23367 44363
rect 23309 44295 23321 44329
rect 23355 44295 23367 44329
rect 23309 44261 23367 44295
rect 23309 44227 23321 44261
rect 23355 44227 23367 44261
rect 23309 44193 23367 44227
rect 23309 44159 23321 44193
rect 23355 44159 23367 44193
rect 23309 44125 23367 44159
rect 23309 44091 23321 44125
rect 23355 44091 23367 44125
rect 23309 44057 23367 44091
rect 23309 44023 23321 44057
rect 23355 44023 23367 44057
rect 23309 43989 23367 44023
rect 23309 43955 23321 43989
rect 23355 43955 23367 43989
rect 23309 43921 23367 43955
rect 23309 43887 23321 43921
rect 23355 43887 23367 43921
rect 23309 43853 23367 43887
rect 23309 43819 23321 43853
rect 23355 43819 23367 43853
rect 23309 43785 23367 43819
rect 23309 43751 23321 43785
rect 23355 43751 23367 43785
rect 23309 43717 23367 43751
rect 23309 43683 23321 43717
rect 23355 43683 23367 43717
rect 23309 43667 23367 43683
rect 23767 44941 23825 44957
rect 23767 44907 23779 44941
rect 23813 44907 23825 44941
rect 23767 44873 23825 44907
rect 23767 44839 23779 44873
rect 23813 44839 23825 44873
rect 23767 44805 23825 44839
rect 23767 44771 23779 44805
rect 23813 44771 23825 44805
rect 23767 44737 23825 44771
rect 23767 44703 23779 44737
rect 23813 44703 23825 44737
rect 23767 44669 23825 44703
rect 23767 44635 23779 44669
rect 23813 44635 23825 44669
rect 23767 44601 23825 44635
rect 23767 44567 23779 44601
rect 23813 44567 23825 44601
rect 23767 44533 23825 44567
rect 23767 44499 23779 44533
rect 23813 44499 23825 44533
rect 23767 44465 23825 44499
rect 23767 44431 23779 44465
rect 23813 44431 23825 44465
rect 23767 44397 23825 44431
rect 23767 44363 23779 44397
rect 23813 44363 23825 44397
rect 23767 44329 23825 44363
rect 23767 44295 23779 44329
rect 23813 44295 23825 44329
rect 23767 44261 23825 44295
rect 23767 44227 23779 44261
rect 23813 44227 23825 44261
rect 23767 44193 23825 44227
rect 23767 44159 23779 44193
rect 23813 44159 23825 44193
rect 23767 44125 23825 44159
rect 23767 44091 23779 44125
rect 23813 44091 23825 44125
rect 23767 44057 23825 44091
rect 23767 44023 23779 44057
rect 23813 44023 23825 44057
rect 23767 43989 23825 44023
rect 23767 43955 23779 43989
rect 23813 43955 23825 43989
rect 23767 43921 23825 43955
rect 23767 43887 23779 43921
rect 23813 43887 23825 43921
rect 23767 43853 23825 43887
rect 23767 43819 23779 43853
rect 23813 43819 23825 43853
rect 23767 43785 23825 43819
rect 23767 43751 23779 43785
rect 23813 43751 23825 43785
rect 23767 43717 23825 43751
rect 23767 43683 23779 43717
rect 23813 43683 23825 43717
rect 23767 43667 23825 43683
rect 24225 44941 24283 44957
rect 24225 44907 24237 44941
rect 24271 44907 24283 44941
rect 24225 44873 24283 44907
rect 24225 44839 24237 44873
rect 24271 44839 24283 44873
rect 24225 44805 24283 44839
rect 24225 44771 24237 44805
rect 24271 44771 24283 44805
rect 24225 44737 24283 44771
rect 24225 44703 24237 44737
rect 24271 44703 24283 44737
rect 24225 44669 24283 44703
rect 24225 44635 24237 44669
rect 24271 44635 24283 44669
rect 24225 44601 24283 44635
rect 24225 44567 24237 44601
rect 24271 44567 24283 44601
rect 24225 44533 24283 44567
rect 24225 44499 24237 44533
rect 24271 44499 24283 44533
rect 24225 44465 24283 44499
rect 24225 44431 24237 44465
rect 24271 44431 24283 44465
rect 24225 44397 24283 44431
rect 24225 44363 24237 44397
rect 24271 44363 24283 44397
rect 24225 44329 24283 44363
rect 24225 44295 24237 44329
rect 24271 44295 24283 44329
rect 24225 44261 24283 44295
rect 24225 44227 24237 44261
rect 24271 44227 24283 44261
rect 24225 44193 24283 44227
rect 24225 44159 24237 44193
rect 24271 44159 24283 44193
rect 24225 44125 24283 44159
rect 24225 44091 24237 44125
rect 24271 44091 24283 44125
rect 24225 44057 24283 44091
rect 24225 44023 24237 44057
rect 24271 44023 24283 44057
rect 24225 43989 24283 44023
rect 24225 43955 24237 43989
rect 24271 43955 24283 43989
rect 24225 43921 24283 43955
rect 24225 43887 24237 43921
rect 24271 43887 24283 43921
rect 24225 43853 24283 43887
rect 24225 43819 24237 43853
rect 24271 43819 24283 43853
rect 24225 43785 24283 43819
rect 24225 43751 24237 43785
rect 24271 43751 24283 43785
rect 24225 43717 24283 43751
rect 24225 43683 24237 43717
rect 24271 43683 24283 43717
rect 24225 43667 24283 43683
rect 24683 44941 24741 44957
rect 24683 44907 24695 44941
rect 24729 44907 24741 44941
rect 24683 44873 24741 44907
rect 24683 44839 24695 44873
rect 24729 44839 24741 44873
rect 24683 44805 24741 44839
rect 24683 44771 24695 44805
rect 24729 44771 24741 44805
rect 24683 44737 24741 44771
rect 24683 44703 24695 44737
rect 24729 44703 24741 44737
rect 24683 44669 24741 44703
rect 24683 44635 24695 44669
rect 24729 44635 24741 44669
rect 24683 44601 24741 44635
rect 24683 44567 24695 44601
rect 24729 44567 24741 44601
rect 24683 44533 24741 44567
rect 24683 44499 24695 44533
rect 24729 44499 24741 44533
rect 24683 44465 24741 44499
rect 24683 44431 24695 44465
rect 24729 44431 24741 44465
rect 24683 44397 24741 44431
rect 24683 44363 24695 44397
rect 24729 44363 24741 44397
rect 24683 44329 24741 44363
rect 24683 44295 24695 44329
rect 24729 44295 24741 44329
rect 24683 44261 24741 44295
rect 24683 44227 24695 44261
rect 24729 44227 24741 44261
rect 24683 44193 24741 44227
rect 24683 44159 24695 44193
rect 24729 44159 24741 44193
rect 24683 44125 24741 44159
rect 24683 44091 24695 44125
rect 24729 44091 24741 44125
rect 24683 44057 24741 44091
rect 24683 44023 24695 44057
rect 24729 44023 24741 44057
rect 24683 43989 24741 44023
rect 24683 43955 24695 43989
rect 24729 43955 24741 43989
rect 24683 43921 24741 43955
rect 24683 43887 24695 43921
rect 24729 43887 24741 43921
rect 24683 43853 24741 43887
rect 24683 43819 24695 43853
rect 24729 43819 24741 43853
rect 24683 43785 24741 43819
rect 24683 43751 24695 43785
rect 24729 43751 24741 43785
rect 24683 43717 24741 43751
rect 24683 43683 24695 43717
rect 24729 43683 24741 43717
rect 24683 43667 24741 43683
rect 25141 44941 25199 44957
rect 25141 44907 25153 44941
rect 25187 44907 25199 44941
rect 25141 44873 25199 44907
rect 25141 44839 25153 44873
rect 25187 44839 25199 44873
rect 25141 44805 25199 44839
rect 25141 44771 25153 44805
rect 25187 44771 25199 44805
rect 25141 44737 25199 44771
rect 25141 44703 25153 44737
rect 25187 44703 25199 44737
rect 25141 44669 25199 44703
rect 25141 44635 25153 44669
rect 25187 44635 25199 44669
rect 25141 44601 25199 44635
rect 25141 44567 25153 44601
rect 25187 44567 25199 44601
rect 25141 44533 25199 44567
rect 25141 44499 25153 44533
rect 25187 44499 25199 44533
rect 25141 44465 25199 44499
rect 25141 44431 25153 44465
rect 25187 44431 25199 44465
rect 25141 44397 25199 44431
rect 25141 44363 25153 44397
rect 25187 44363 25199 44397
rect 25141 44329 25199 44363
rect 25141 44295 25153 44329
rect 25187 44295 25199 44329
rect 25141 44261 25199 44295
rect 25141 44227 25153 44261
rect 25187 44227 25199 44261
rect 25141 44193 25199 44227
rect 25141 44159 25153 44193
rect 25187 44159 25199 44193
rect 25141 44125 25199 44159
rect 25141 44091 25153 44125
rect 25187 44091 25199 44125
rect 25141 44057 25199 44091
rect 25141 44023 25153 44057
rect 25187 44023 25199 44057
rect 25141 43989 25199 44023
rect 25141 43955 25153 43989
rect 25187 43955 25199 43989
rect 25141 43921 25199 43955
rect 25141 43887 25153 43921
rect 25187 43887 25199 43921
rect 25141 43853 25199 43887
rect 25141 43819 25153 43853
rect 25187 43819 25199 43853
rect 25141 43785 25199 43819
rect 25141 43751 25153 43785
rect 25187 43751 25199 43785
rect 25141 43717 25199 43751
rect 25141 43683 25153 43717
rect 25187 43683 25199 43717
rect 25141 43667 25199 43683
rect 25599 44941 25657 44957
rect 25599 44907 25611 44941
rect 25645 44907 25657 44941
rect 25599 44873 25657 44907
rect 25599 44839 25611 44873
rect 25645 44839 25657 44873
rect 25599 44805 25657 44839
rect 25599 44771 25611 44805
rect 25645 44771 25657 44805
rect 25599 44737 25657 44771
rect 25599 44703 25611 44737
rect 25645 44703 25657 44737
rect 25599 44669 25657 44703
rect 25599 44635 25611 44669
rect 25645 44635 25657 44669
rect 25599 44601 25657 44635
rect 25599 44567 25611 44601
rect 25645 44567 25657 44601
rect 25599 44533 25657 44567
rect 25599 44499 25611 44533
rect 25645 44499 25657 44533
rect 25599 44465 25657 44499
rect 25599 44431 25611 44465
rect 25645 44431 25657 44465
rect 25599 44397 25657 44431
rect 25599 44363 25611 44397
rect 25645 44363 25657 44397
rect 25599 44329 25657 44363
rect 25599 44295 25611 44329
rect 25645 44295 25657 44329
rect 25599 44261 25657 44295
rect 25599 44227 25611 44261
rect 25645 44227 25657 44261
rect 25599 44193 25657 44227
rect 25599 44159 25611 44193
rect 25645 44159 25657 44193
rect 25599 44125 25657 44159
rect 25599 44091 25611 44125
rect 25645 44091 25657 44125
rect 25599 44057 25657 44091
rect 25599 44023 25611 44057
rect 25645 44023 25657 44057
rect 25599 43989 25657 44023
rect 25599 43955 25611 43989
rect 25645 43955 25657 43989
rect 25599 43921 25657 43955
rect 25599 43887 25611 43921
rect 25645 43887 25657 43921
rect 25599 43853 25657 43887
rect 25599 43819 25611 43853
rect 25645 43819 25657 43853
rect 25599 43785 25657 43819
rect 25599 43751 25611 43785
rect 25645 43751 25657 43785
rect 25599 43717 25657 43751
rect 25599 43683 25611 43717
rect 25645 43683 25657 43717
rect 25599 43667 25657 43683
rect 26057 44941 26115 44957
rect 26057 44907 26069 44941
rect 26103 44907 26115 44941
rect 26057 44873 26115 44907
rect 26057 44839 26069 44873
rect 26103 44839 26115 44873
rect 26057 44805 26115 44839
rect 26057 44771 26069 44805
rect 26103 44771 26115 44805
rect 26057 44737 26115 44771
rect 26057 44703 26069 44737
rect 26103 44703 26115 44737
rect 26057 44669 26115 44703
rect 26057 44635 26069 44669
rect 26103 44635 26115 44669
rect 26057 44601 26115 44635
rect 26057 44567 26069 44601
rect 26103 44567 26115 44601
rect 26057 44533 26115 44567
rect 26057 44499 26069 44533
rect 26103 44499 26115 44533
rect 26057 44465 26115 44499
rect 26057 44431 26069 44465
rect 26103 44431 26115 44465
rect 26057 44397 26115 44431
rect 26057 44363 26069 44397
rect 26103 44363 26115 44397
rect 26057 44329 26115 44363
rect 26057 44295 26069 44329
rect 26103 44295 26115 44329
rect 26057 44261 26115 44295
rect 26057 44227 26069 44261
rect 26103 44227 26115 44261
rect 26057 44193 26115 44227
rect 26057 44159 26069 44193
rect 26103 44159 26115 44193
rect 26057 44125 26115 44159
rect 26057 44091 26069 44125
rect 26103 44091 26115 44125
rect 26057 44057 26115 44091
rect 26057 44023 26069 44057
rect 26103 44023 26115 44057
rect 26057 43989 26115 44023
rect 26057 43955 26069 43989
rect 26103 43955 26115 43989
rect 26057 43921 26115 43955
rect 26057 43887 26069 43921
rect 26103 43887 26115 43921
rect 26057 43853 26115 43887
rect 26057 43819 26069 43853
rect 26103 43819 26115 43853
rect 26057 43785 26115 43819
rect 26057 43751 26069 43785
rect 26103 43751 26115 43785
rect 26057 43717 26115 43751
rect 26057 43683 26069 43717
rect 26103 43683 26115 43717
rect 26057 43667 26115 43683
rect 26515 44941 26573 44957
rect 26515 44907 26527 44941
rect 26561 44907 26573 44941
rect 26515 44873 26573 44907
rect 26515 44839 26527 44873
rect 26561 44839 26573 44873
rect 26515 44805 26573 44839
rect 26515 44771 26527 44805
rect 26561 44771 26573 44805
rect 26515 44737 26573 44771
rect 26515 44703 26527 44737
rect 26561 44703 26573 44737
rect 26515 44669 26573 44703
rect 26515 44635 26527 44669
rect 26561 44635 26573 44669
rect 26515 44601 26573 44635
rect 26515 44567 26527 44601
rect 26561 44567 26573 44601
rect 26515 44533 26573 44567
rect 26515 44499 26527 44533
rect 26561 44499 26573 44533
rect 26515 44465 26573 44499
rect 26515 44431 26527 44465
rect 26561 44431 26573 44465
rect 26515 44397 26573 44431
rect 26515 44363 26527 44397
rect 26561 44363 26573 44397
rect 26515 44329 26573 44363
rect 26515 44295 26527 44329
rect 26561 44295 26573 44329
rect 26515 44261 26573 44295
rect 26515 44227 26527 44261
rect 26561 44227 26573 44261
rect 26515 44193 26573 44227
rect 26515 44159 26527 44193
rect 26561 44159 26573 44193
rect 26515 44125 26573 44159
rect 26515 44091 26527 44125
rect 26561 44091 26573 44125
rect 26515 44057 26573 44091
rect 26515 44023 26527 44057
rect 26561 44023 26573 44057
rect 26515 43989 26573 44023
rect 26515 43955 26527 43989
rect 26561 43955 26573 43989
rect 26515 43921 26573 43955
rect 26515 43887 26527 43921
rect 26561 43887 26573 43921
rect 26515 43853 26573 43887
rect 26515 43819 26527 43853
rect 26561 43819 26573 43853
rect 26515 43785 26573 43819
rect 26515 43751 26527 43785
rect 26561 43751 26573 43785
rect 26515 43717 26573 43751
rect 26515 43683 26527 43717
rect 26561 43683 26573 43717
rect 26515 43667 26573 43683
rect 26973 44941 27031 44957
rect 26973 44907 26985 44941
rect 27019 44907 27031 44941
rect 26973 44873 27031 44907
rect 26973 44839 26985 44873
rect 27019 44839 27031 44873
rect 26973 44805 27031 44839
rect 26973 44771 26985 44805
rect 27019 44771 27031 44805
rect 26973 44737 27031 44771
rect 26973 44703 26985 44737
rect 27019 44703 27031 44737
rect 26973 44669 27031 44703
rect 26973 44635 26985 44669
rect 27019 44635 27031 44669
rect 26973 44601 27031 44635
rect 26973 44567 26985 44601
rect 27019 44567 27031 44601
rect 26973 44533 27031 44567
rect 26973 44499 26985 44533
rect 27019 44499 27031 44533
rect 26973 44465 27031 44499
rect 26973 44431 26985 44465
rect 27019 44431 27031 44465
rect 26973 44397 27031 44431
rect 26973 44363 26985 44397
rect 27019 44363 27031 44397
rect 26973 44329 27031 44363
rect 26973 44295 26985 44329
rect 27019 44295 27031 44329
rect 26973 44261 27031 44295
rect 26973 44227 26985 44261
rect 27019 44227 27031 44261
rect 26973 44193 27031 44227
rect 26973 44159 26985 44193
rect 27019 44159 27031 44193
rect 26973 44125 27031 44159
rect 26973 44091 26985 44125
rect 27019 44091 27031 44125
rect 26973 44057 27031 44091
rect 26973 44023 26985 44057
rect 27019 44023 27031 44057
rect 26973 43989 27031 44023
rect 26973 43955 26985 43989
rect 27019 43955 27031 43989
rect 26973 43921 27031 43955
rect 26973 43887 26985 43921
rect 27019 43887 27031 43921
rect 26973 43853 27031 43887
rect 26973 43819 26985 43853
rect 27019 43819 27031 43853
rect 26973 43785 27031 43819
rect 26973 43751 26985 43785
rect 27019 43751 27031 43785
rect 26973 43717 27031 43751
rect 26973 43683 26985 43717
rect 27019 43683 27031 43717
rect 26973 43667 27031 43683
rect 27431 44941 27489 44957
rect 27431 44907 27443 44941
rect 27477 44907 27489 44941
rect 27431 44873 27489 44907
rect 27431 44839 27443 44873
rect 27477 44839 27489 44873
rect 27431 44805 27489 44839
rect 27431 44771 27443 44805
rect 27477 44771 27489 44805
rect 27431 44737 27489 44771
rect 27431 44703 27443 44737
rect 27477 44703 27489 44737
rect 27431 44669 27489 44703
rect 27431 44635 27443 44669
rect 27477 44635 27489 44669
rect 27431 44601 27489 44635
rect 27431 44567 27443 44601
rect 27477 44567 27489 44601
rect 27431 44533 27489 44567
rect 27431 44499 27443 44533
rect 27477 44499 27489 44533
rect 27431 44465 27489 44499
rect 27431 44431 27443 44465
rect 27477 44431 27489 44465
rect 27431 44397 27489 44431
rect 27431 44363 27443 44397
rect 27477 44363 27489 44397
rect 27431 44329 27489 44363
rect 27431 44295 27443 44329
rect 27477 44295 27489 44329
rect 27431 44261 27489 44295
rect 27431 44227 27443 44261
rect 27477 44227 27489 44261
rect 27431 44193 27489 44227
rect 27431 44159 27443 44193
rect 27477 44159 27489 44193
rect 27431 44125 27489 44159
rect 27431 44091 27443 44125
rect 27477 44091 27489 44125
rect 27431 44057 27489 44091
rect 27431 44023 27443 44057
rect 27477 44023 27489 44057
rect 27431 43989 27489 44023
rect 27431 43955 27443 43989
rect 27477 43955 27489 43989
rect 27431 43921 27489 43955
rect 27431 43887 27443 43921
rect 27477 43887 27489 43921
rect 27431 43853 27489 43887
rect 27431 43819 27443 43853
rect 27477 43819 27489 43853
rect 27431 43785 27489 43819
rect 27431 43751 27443 43785
rect 27477 43751 27489 43785
rect 27431 43717 27489 43751
rect 27431 43683 27443 43717
rect 27477 43683 27489 43717
rect 27431 43667 27489 43683
rect 27889 44941 27947 44957
rect 27889 44907 27901 44941
rect 27935 44907 27947 44941
rect 27889 44873 27947 44907
rect 27889 44839 27901 44873
rect 27935 44839 27947 44873
rect 27889 44805 27947 44839
rect 27889 44771 27901 44805
rect 27935 44771 27947 44805
rect 27889 44737 27947 44771
rect 27889 44703 27901 44737
rect 27935 44703 27947 44737
rect 27889 44669 27947 44703
rect 27889 44635 27901 44669
rect 27935 44635 27947 44669
rect 27889 44601 27947 44635
rect 27889 44567 27901 44601
rect 27935 44567 27947 44601
rect 27889 44533 27947 44567
rect 27889 44499 27901 44533
rect 27935 44499 27947 44533
rect 27889 44465 27947 44499
rect 27889 44431 27901 44465
rect 27935 44431 27947 44465
rect 27889 44397 27947 44431
rect 27889 44363 27901 44397
rect 27935 44363 27947 44397
rect 27889 44329 27947 44363
rect 27889 44295 27901 44329
rect 27935 44295 27947 44329
rect 27889 44261 27947 44295
rect 27889 44227 27901 44261
rect 27935 44227 27947 44261
rect 27889 44193 27947 44227
rect 27889 44159 27901 44193
rect 27935 44159 27947 44193
rect 27889 44125 27947 44159
rect 27889 44091 27901 44125
rect 27935 44091 27947 44125
rect 27889 44057 27947 44091
rect 27889 44023 27901 44057
rect 27935 44023 27947 44057
rect 27889 43989 27947 44023
rect 27889 43955 27901 43989
rect 27935 43955 27947 43989
rect 27889 43921 27947 43955
rect 27889 43887 27901 43921
rect 27935 43887 27947 43921
rect 27889 43853 27947 43887
rect 27889 43819 27901 43853
rect 27935 43819 27947 43853
rect 27889 43785 27947 43819
rect 27889 43751 27901 43785
rect 27935 43751 27947 43785
rect 27889 43717 27947 43751
rect 27889 43683 27901 43717
rect 27935 43683 27947 43717
rect 27889 43667 27947 43683
rect 28347 44941 28405 44957
rect 28347 44907 28359 44941
rect 28393 44907 28405 44941
rect 28347 44873 28405 44907
rect 28347 44839 28359 44873
rect 28393 44839 28405 44873
rect 28347 44805 28405 44839
rect 28347 44771 28359 44805
rect 28393 44771 28405 44805
rect 28347 44737 28405 44771
rect 28347 44703 28359 44737
rect 28393 44703 28405 44737
rect 28347 44669 28405 44703
rect 28347 44635 28359 44669
rect 28393 44635 28405 44669
rect 28347 44601 28405 44635
rect 28347 44567 28359 44601
rect 28393 44567 28405 44601
rect 28347 44533 28405 44567
rect 28347 44499 28359 44533
rect 28393 44499 28405 44533
rect 28347 44465 28405 44499
rect 28347 44431 28359 44465
rect 28393 44431 28405 44465
rect 28347 44397 28405 44431
rect 28347 44363 28359 44397
rect 28393 44363 28405 44397
rect 28347 44329 28405 44363
rect 28347 44295 28359 44329
rect 28393 44295 28405 44329
rect 28347 44261 28405 44295
rect 28347 44227 28359 44261
rect 28393 44227 28405 44261
rect 28347 44193 28405 44227
rect 28347 44159 28359 44193
rect 28393 44159 28405 44193
rect 28347 44125 28405 44159
rect 28347 44091 28359 44125
rect 28393 44091 28405 44125
rect 28347 44057 28405 44091
rect 28347 44023 28359 44057
rect 28393 44023 28405 44057
rect 28347 43989 28405 44023
rect 28347 43955 28359 43989
rect 28393 43955 28405 43989
rect 28347 43921 28405 43955
rect 28347 43887 28359 43921
rect 28393 43887 28405 43921
rect 28347 43853 28405 43887
rect 28347 43819 28359 43853
rect 28393 43819 28405 43853
rect 28347 43785 28405 43819
rect 28347 43751 28359 43785
rect 28393 43751 28405 43785
rect 28347 43717 28405 43751
rect 28347 43683 28359 43717
rect 28393 43683 28405 43717
rect 28347 43667 28405 43683
rect 28805 44941 28863 44957
rect 28805 44907 28817 44941
rect 28851 44907 28863 44941
rect 28805 44873 28863 44907
rect 28805 44839 28817 44873
rect 28851 44839 28863 44873
rect 28805 44805 28863 44839
rect 28805 44771 28817 44805
rect 28851 44771 28863 44805
rect 28805 44737 28863 44771
rect 28805 44703 28817 44737
rect 28851 44703 28863 44737
rect 28805 44669 28863 44703
rect 28805 44635 28817 44669
rect 28851 44635 28863 44669
rect 28805 44601 28863 44635
rect 28805 44567 28817 44601
rect 28851 44567 28863 44601
rect 28805 44533 28863 44567
rect 28805 44499 28817 44533
rect 28851 44499 28863 44533
rect 28805 44465 28863 44499
rect 28805 44431 28817 44465
rect 28851 44431 28863 44465
rect 28805 44397 28863 44431
rect 28805 44363 28817 44397
rect 28851 44363 28863 44397
rect 28805 44329 28863 44363
rect 28805 44295 28817 44329
rect 28851 44295 28863 44329
rect 28805 44261 28863 44295
rect 28805 44227 28817 44261
rect 28851 44227 28863 44261
rect 28805 44193 28863 44227
rect 28805 44159 28817 44193
rect 28851 44159 28863 44193
rect 28805 44125 28863 44159
rect 28805 44091 28817 44125
rect 28851 44091 28863 44125
rect 28805 44057 28863 44091
rect 28805 44023 28817 44057
rect 28851 44023 28863 44057
rect 28805 43989 28863 44023
rect 28805 43955 28817 43989
rect 28851 43955 28863 43989
rect 28805 43921 28863 43955
rect 28805 43887 28817 43921
rect 28851 43887 28863 43921
rect 28805 43853 28863 43887
rect 28805 43819 28817 43853
rect 28851 43819 28863 43853
rect 28805 43785 28863 43819
rect 28805 43751 28817 43785
rect 28851 43751 28863 43785
rect 28805 43717 28863 43751
rect 28805 43683 28817 43717
rect 28851 43683 28863 43717
rect 28805 43667 28863 43683
rect 29263 44941 29321 44957
rect 29263 44907 29275 44941
rect 29309 44907 29321 44941
rect 29263 44873 29321 44907
rect 29263 44839 29275 44873
rect 29309 44839 29321 44873
rect 29263 44805 29321 44839
rect 29263 44771 29275 44805
rect 29309 44771 29321 44805
rect 29263 44737 29321 44771
rect 29263 44703 29275 44737
rect 29309 44703 29321 44737
rect 29263 44669 29321 44703
rect 29263 44635 29275 44669
rect 29309 44635 29321 44669
rect 29263 44601 29321 44635
rect 29263 44567 29275 44601
rect 29309 44567 29321 44601
rect 29263 44533 29321 44567
rect 29263 44499 29275 44533
rect 29309 44499 29321 44533
rect 29263 44465 29321 44499
rect 29263 44431 29275 44465
rect 29309 44431 29321 44465
rect 29263 44397 29321 44431
rect 29263 44363 29275 44397
rect 29309 44363 29321 44397
rect 29263 44329 29321 44363
rect 29263 44295 29275 44329
rect 29309 44295 29321 44329
rect 29263 44261 29321 44295
rect 29263 44227 29275 44261
rect 29309 44227 29321 44261
rect 29263 44193 29321 44227
rect 29263 44159 29275 44193
rect 29309 44159 29321 44193
rect 29263 44125 29321 44159
rect 29263 44091 29275 44125
rect 29309 44091 29321 44125
rect 29263 44057 29321 44091
rect 29263 44023 29275 44057
rect 29309 44023 29321 44057
rect 29263 43989 29321 44023
rect 29263 43955 29275 43989
rect 29309 43955 29321 43989
rect 29263 43921 29321 43955
rect 29263 43887 29275 43921
rect 29309 43887 29321 43921
rect 29263 43853 29321 43887
rect 29263 43819 29275 43853
rect 29309 43819 29321 43853
rect 29263 43785 29321 43819
rect 29263 43751 29275 43785
rect 29309 43751 29321 43785
rect 29263 43717 29321 43751
rect 29263 43683 29275 43717
rect 29309 43683 29321 43717
rect 29263 43667 29321 43683
rect 29721 44941 29779 44957
rect 29721 44907 29733 44941
rect 29767 44907 29779 44941
rect 29721 44873 29779 44907
rect 29721 44839 29733 44873
rect 29767 44839 29779 44873
rect 29721 44805 29779 44839
rect 29721 44771 29733 44805
rect 29767 44771 29779 44805
rect 29721 44737 29779 44771
rect 29721 44703 29733 44737
rect 29767 44703 29779 44737
rect 29721 44669 29779 44703
rect 29721 44635 29733 44669
rect 29767 44635 29779 44669
rect 29721 44601 29779 44635
rect 29721 44567 29733 44601
rect 29767 44567 29779 44601
rect 29721 44533 29779 44567
rect 29721 44499 29733 44533
rect 29767 44499 29779 44533
rect 29721 44465 29779 44499
rect 29721 44431 29733 44465
rect 29767 44431 29779 44465
rect 29721 44397 29779 44431
rect 29721 44363 29733 44397
rect 29767 44363 29779 44397
rect 29721 44329 29779 44363
rect 29721 44295 29733 44329
rect 29767 44295 29779 44329
rect 29721 44261 29779 44295
rect 29721 44227 29733 44261
rect 29767 44227 29779 44261
rect 29721 44193 29779 44227
rect 29721 44159 29733 44193
rect 29767 44159 29779 44193
rect 29721 44125 29779 44159
rect 29721 44091 29733 44125
rect 29767 44091 29779 44125
rect 29721 44057 29779 44091
rect 29721 44023 29733 44057
rect 29767 44023 29779 44057
rect 29721 43989 29779 44023
rect 29721 43955 29733 43989
rect 29767 43955 29779 43989
rect 29721 43921 29779 43955
rect 29721 43887 29733 43921
rect 29767 43887 29779 43921
rect 29721 43853 29779 43887
rect 29721 43819 29733 43853
rect 29767 43819 29779 43853
rect 29721 43785 29779 43819
rect 29721 43751 29733 43785
rect 29767 43751 29779 43785
rect 29721 43717 29779 43751
rect 29721 43683 29733 43717
rect 29767 43683 29779 43717
rect 29721 43667 29779 43683
rect 30179 44941 30237 44957
rect 30179 44907 30191 44941
rect 30225 44907 30237 44941
rect 30179 44873 30237 44907
rect 30179 44839 30191 44873
rect 30225 44839 30237 44873
rect 30179 44805 30237 44839
rect 30179 44771 30191 44805
rect 30225 44771 30237 44805
rect 30179 44737 30237 44771
rect 30179 44703 30191 44737
rect 30225 44703 30237 44737
rect 30179 44669 30237 44703
rect 30179 44635 30191 44669
rect 30225 44635 30237 44669
rect 30179 44601 30237 44635
rect 30179 44567 30191 44601
rect 30225 44567 30237 44601
rect 30179 44533 30237 44567
rect 30179 44499 30191 44533
rect 30225 44499 30237 44533
rect 30179 44465 30237 44499
rect 30179 44431 30191 44465
rect 30225 44431 30237 44465
rect 30179 44397 30237 44431
rect 30179 44363 30191 44397
rect 30225 44363 30237 44397
rect 30179 44329 30237 44363
rect 30179 44295 30191 44329
rect 30225 44295 30237 44329
rect 30179 44261 30237 44295
rect 30179 44227 30191 44261
rect 30225 44227 30237 44261
rect 30179 44193 30237 44227
rect 30179 44159 30191 44193
rect 30225 44159 30237 44193
rect 30179 44125 30237 44159
rect 30179 44091 30191 44125
rect 30225 44091 30237 44125
rect 30179 44057 30237 44091
rect 30179 44023 30191 44057
rect 30225 44023 30237 44057
rect 30179 43989 30237 44023
rect 30179 43955 30191 43989
rect 30225 43955 30237 43989
rect 30179 43921 30237 43955
rect 30179 43887 30191 43921
rect 30225 43887 30237 43921
rect 30179 43853 30237 43887
rect 30179 43819 30191 43853
rect 30225 43819 30237 43853
rect 30179 43785 30237 43819
rect 30179 43751 30191 43785
rect 30225 43751 30237 43785
rect 30179 43717 30237 43751
rect 30179 43683 30191 43717
rect 30225 43683 30237 43717
rect 30179 43667 30237 43683
rect 30637 44941 30695 44957
rect 30637 44907 30649 44941
rect 30683 44907 30695 44941
rect 30637 44873 30695 44907
rect 30637 44839 30649 44873
rect 30683 44839 30695 44873
rect 30637 44805 30695 44839
rect 30637 44771 30649 44805
rect 30683 44771 30695 44805
rect 30637 44737 30695 44771
rect 30637 44703 30649 44737
rect 30683 44703 30695 44737
rect 30637 44669 30695 44703
rect 30637 44635 30649 44669
rect 30683 44635 30695 44669
rect 30637 44601 30695 44635
rect 30637 44567 30649 44601
rect 30683 44567 30695 44601
rect 30637 44533 30695 44567
rect 30637 44499 30649 44533
rect 30683 44499 30695 44533
rect 30637 44465 30695 44499
rect 30637 44431 30649 44465
rect 30683 44431 30695 44465
rect 30637 44397 30695 44431
rect 30637 44363 30649 44397
rect 30683 44363 30695 44397
rect 30637 44329 30695 44363
rect 30637 44295 30649 44329
rect 30683 44295 30695 44329
rect 30637 44261 30695 44295
rect 30637 44227 30649 44261
rect 30683 44227 30695 44261
rect 30637 44193 30695 44227
rect 30637 44159 30649 44193
rect 30683 44159 30695 44193
rect 30637 44125 30695 44159
rect 30637 44091 30649 44125
rect 30683 44091 30695 44125
rect 30637 44057 30695 44091
rect 30637 44023 30649 44057
rect 30683 44023 30695 44057
rect 30637 43989 30695 44023
rect 30637 43955 30649 43989
rect 30683 43955 30695 43989
rect 30637 43921 30695 43955
rect 30637 43887 30649 43921
rect 30683 43887 30695 43921
rect 30637 43853 30695 43887
rect 30637 43819 30649 43853
rect 30683 43819 30695 43853
rect 30637 43785 30695 43819
rect 30637 43751 30649 43785
rect 30683 43751 30695 43785
rect 30637 43717 30695 43751
rect 30637 43683 30649 43717
rect 30683 43683 30695 43717
rect 30637 43667 30695 43683
rect 31095 44941 31153 44957
rect 31095 44907 31107 44941
rect 31141 44907 31153 44941
rect 31095 44873 31153 44907
rect 31095 44839 31107 44873
rect 31141 44839 31153 44873
rect 31095 44805 31153 44839
rect 31095 44771 31107 44805
rect 31141 44771 31153 44805
rect 31095 44737 31153 44771
rect 31095 44703 31107 44737
rect 31141 44703 31153 44737
rect 31095 44669 31153 44703
rect 31095 44635 31107 44669
rect 31141 44635 31153 44669
rect 31095 44601 31153 44635
rect 31095 44567 31107 44601
rect 31141 44567 31153 44601
rect 31095 44533 31153 44567
rect 31095 44499 31107 44533
rect 31141 44499 31153 44533
rect 31095 44465 31153 44499
rect 31095 44431 31107 44465
rect 31141 44431 31153 44465
rect 31095 44397 31153 44431
rect 31095 44363 31107 44397
rect 31141 44363 31153 44397
rect 31095 44329 31153 44363
rect 31095 44295 31107 44329
rect 31141 44295 31153 44329
rect 31095 44261 31153 44295
rect 31095 44227 31107 44261
rect 31141 44227 31153 44261
rect 31095 44193 31153 44227
rect 31095 44159 31107 44193
rect 31141 44159 31153 44193
rect 31095 44125 31153 44159
rect 31095 44091 31107 44125
rect 31141 44091 31153 44125
rect 31095 44057 31153 44091
rect 31095 44023 31107 44057
rect 31141 44023 31153 44057
rect 31095 43989 31153 44023
rect 31095 43955 31107 43989
rect 31141 43955 31153 43989
rect 31095 43921 31153 43955
rect 31095 43887 31107 43921
rect 31141 43887 31153 43921
rect 31095 43853 31153 43887
rect 31095 43819 31107 43853
rect 31141 43819 31153 43853
rect 31095 43785 31153 43819
rect 31095 43751 31107 43785
rect 31141 43751 31153 43785
rect 31095 43717 31153 43751
rect 31095 43683 31107 43717
rect 31141 43683 31153 43717
rect 31095 43667 31153 43683
rect 31553 44941 31611 44957
rect 31553 44907 31565 44941
rect 31599 44907 31611 44941
rect 31553 44873 31611 44907
rect 31553 44839 31565 44873
rect 31599 44839 31611 44873
rect 31553 44805 31611 44839
rect 31553 44771 31565 44805
rect 31599 44771 31611 44805
rect 31553 44737 31611 44771
rect 31553 44703 31565 44737
rect 31599 44703 31611 44737
rect 31553 44669 31611 44703
rect 31553 44635 31565 44669
rect 31599 44635 31611 44669
rect 31553 44601 31611 44635
rect 31553 44567 31565 44601
rect 31599 44567 31611 44601
rect 31553 44533 31611 44567
rect 31553 44499 31565 44533
rect 31599 44499 31611 44533
rect 31553 44465 31611 44499
rect 31553 44431 31565 44465
rect 31599 44431 31611 44465
rect 31553 44397 31611 44431
rect 31553 44363 31565 44397
rect 31599 44363 31611 44397
rect 31553 44329 31611 44363
rect 31553 44295 31565 44329
rect 31599 44295 31611 44329
rect 31553 44261 31611 44295
rect 31553 44227 31565 44261
rect 31599 44227 31611 44261
rect 31553 44193 31611 44227
rect 31553 44159 31565 44193
rect 31599 44159 31611 44193
rect 31553 44125 31611 44159
rect 31553 44091 31565 44125
rect 31599 44091 31611 44125
rect 31553 44057 31611 44091
rect 31553 44023 31565 44057
rect 31599 44023 31611 44057
rect 31553 43989 31611 44023
rect 31553 43955 31565 43989
rect 31599 43955 31611 43989
rect 31553 43921 31611 43955
rect 31553 43887 31565 43921
rect 31599 43887 31611 43921
rect 31553 43853 31611 43887
rect 31553 43819 31565 43853
rect 31599 43819 31611 43853
rect 31553 43785 31611 43819
rect 31553 43751 31565 43785
rect 31599 43751 31611 43785
rect 31553 43717 31611 43751
rect 31553 43683 31565 43717
rect 31599 43683 31611 43717
rect 31553 43667 31611 43683
rect 32011 44941 32069 44957
rect 32011 44907 32023 44941
rect 32057 44907 32069 44941
rect 32011 44873 32069 44907
rect 32011 44839 32023 44873
rect 32057 44839 32069 44873
rect 32011 44805 32069 44839
rect 32011 44771 32023 44805
rect 32057 44771 32069 44805
rect 32011 44737 32069 44771
rect 32011 44703 32023 44737
rect 32057 44703 32069 44737
rect 32011 44669 32069 44703
rect 32011 44635 32023 44669
rect 32057 44635 32069 44669
rect 32011 44601 32069 44635
rect 32011 44567 32023 44601
rect 32057 44567 32069 44601
rect 32011 44533 32069 44567
rect 32011 44499 32023 44533
rect 32057 44499 32069 44533
rect 32011 44465 32069 44499
rect 32011 44431 32023 44465
rect 32057 44431 32069 44465
rect 32011 44397 32069 44431
rect 32011 44363 32023 44397
rect 32057 44363 32069 44397
rect 32011 44329 32069 44363
rect 32011 44295 32023 44329
rect 32057 44295 32069 44329
rect 32011 44261 32069 44295
rect 32011 44227 32023 44261
rect 32057 44227 32069 44261
rect 32011 44193 32069 44227
rect 32011 44159 32023 44193
rect 32057 44159 32069 44193
rect 32011 44125 32069 44159
rect 32011 44091 32023 44125
rect 32057 44091 32069 44125
rect 32011 44057 32069 44091
rect 32011 44023 32023 44057
rect 32057 44023 32069 44057
rect 32011 43989 32069 44023
rect 32011 43955 32023 43989
rect 32057 43955 32069 43989
rect 32011 43921 32069 43955
rect 32011 43887 32023 43921
rect 32057 43887 32069 43921
rect 32011 43853 32069 43887
rect 32011 43819 32023 43853
rect 32057 43819 32069 43853
rect 32011 43785 32069 43819
rect 32011 43751 32023 43785
rect 32057 43751 32069 43785
rect 32011 43717 32069 43751
rect 32011 43683 32023 43717
rect 32057 43683 32069 43717
rect 32011 43667 32069 43683
rect 32469 44941 32527 44957
rect 32469 44907 32481 44941
rect 32515 44907 32527 44941
rect 32469 44873 32527 44907
rect 32469 44839 32481 44873
rect 32515 44839 32527 44873
rect 32469 44805 32527 44839
rect 32469 44771 32481 44805
rect 32515 44771 32527 44805
rect 32469 44737 32527 44771
rect 32469 44703 32481 44737
rect 32515 44703 32527 44737
rect 32469 44669 32527 44703
rect 32469 44635 32481 44669
rect 32515 44635 32527 44669
rect 32469 44601 32527 44635
rect 32469 44567 32481 44601
rect 32515 44567 32527 44601
rect 32469 44533 32527 44567
rect 32469 44499 32481 44533
rect 32515 44499 32527 44533
rect 32469 44465 32527 44499
rect 32469 44431 32481 44465
rect 32515 44431 32527 44465
rect 32469 44397 32527 44431
rect 32469 44363 32481 44397
rect 32515 44363 32527 44397
rect 32469 44329 32527 44363
rect 32469 44295 32481 44329
rect 32515 44295 32527 44329
rect 32469 44261 32527 44295
rect 32469 44227 32481 44261
rect 32515 44227 32527 44261
rect 32469 44193 32527 44227
rect 32469 44159 32481 44193
rect 32515 44159 32527 44193
rect 32469 44125 32527 44159
rect 32469 44091 32481 44125
rect 32515 44091 32527 44125
rect 32469 44057 32527 44091
rect 32469 44023 32481 44057
rect 32515 44023 32527 44057
rect 32469 43989 32527 44023
rect 32469 43955 32481 43989
rect 32515 43955 32527 43989
rect 32469 43921 32527 43955
rect 32469 43887 32481 43921
rect 32515 43887 32527 43921
rect 32469 43853 32527 43887
rect 32469 43819 32481 43853
rect 32515 43819 32527 43853
rect 32469 43785 32527 43819
rect 32469 43751 32481 43785
rect 32515 43751 32527 43785
rect 32469 43717 32527 43751
rect 32469 43683 32481 43717
rect 32515 43683 32527 43717
rect 32469 43667 32527 43683
rect 32927 44941 32985 44957
rect 32927 44907 32939 44941
rect 32973 44907 32985 44941
rect 32927 44873 32985 44907
rect 32927 44839 32939 44873
rect 32973 44839 32985 44873
rect 32927 44805 32985 44839
rect 32927 44771 32939 44805
rect 32973 44771 32985 44805
rect 32927 44737 32985 44771
rect 32927 44703 32939 44737
rect 32973 44703 32985 44737
rect 32927 44669 32985 44703
rect 32927 44635 32939 44669
rect 32973 44635 32985 44669
rect 32927 44601 32985 44635
rect 32927 44567 32939 44601
rect 32973 44567 32985 44601
rect 32927 44533 32985 44567
rect 32927 44499 32939 44533
rect 32973 44499 32985 44533
rect 32927 44465 32985 44499
rect 32927 44431 32939 44465
rect 32973 44431 32985 44465
rect 32927 44397 32985 44431
rect 32927 44363 32939 44397
rect 32973 44363 32985 44397
rect 32927 44329 32985 44363
rect 32927 44295 32939 44329
rect 32973 44295 32985 44329
rect 32927 44261 32985 44295
rect 32927 44227 32939 44261
rect 32973 44227 32985 44261
rect 32927 44193 32985 44227
rect 32927 44159 32939 44193
rect 32973 44159 32985 44193
rect 32927 44125 32985 44159
rect 32927 44091 32939 44125
rect 32973 44091 32985 44125
rect 32927 44057 32985 44091
rect 32927 44023 32939 44057
rect 32973 44023 32985 44057
rect 32927 43989 32985 44023
rect 32927 43955 32939 43989
rect 32973 43955 32985 43989
rect 32927 43921 32985 43955
rect 32927 43887 32939 43921
rect 32973 43887 32985 43921
rect 32927 43853 32985 43887
rect 32927 43819 32939 43853
rect 32973 43819 32985 43853
rect 32927 43785 32985 43819
rect 32927 43751 32939 43785
rect 32973 43751 32985 43785
rect 32927 43717 32985 43751
rect 32927 43683 32939 43717
rect 32973 43683 32985 43717
rect 32927 43667 32985 43683
rect 33385 44941 33443 44957
rect 33385 44907 33397 44941
rect 33431 44907 33443 44941
rect 33385 44873 33443 44907
rect 33385 44839 33397 44873
rect 33431 44839 33443 44873
rect 33385 44805 33443 44839
rect 33385 44771 33397 44805
rect 33431 44771 33443 44805
rect 33385 44737 33443 44771
rect 33385 44703 33397 44737
rect 33431 44703 33443 44737
rect 33385 44669 33443 44703
rect 33385 44635 33397 44669
rect 33431 44635 33443 44669
rect 33385 44601 33443 44635
rect 33385 44567 33397 44601
rect 33431 44567 33443 44601
rect 33385 44533 33443 44567
rect 33385 44499 33397 44533
rect 33431 44499 33443 44533
rect 33385 44465 33443 44499
rect 33385 44431 33397 44465
rect 33431 44431 33443 44465
rect 33385 44397 33443 44431
rect 33385 44363 33397 44397
rect 33431 44363 33443 44397
rect 33385 44329 33443 44363
rect 33385 44295 33397 44329
rect 33431 44295 33443 44329
rect 33385 44261 33443 44295
rect 33385 44227 33397 44261
rect 33431 44227 33443 44261
rect 33385 44193 33443 44227
rect 33385 44159 33397 44193
rect 33431 44159 33443 44193
rect 33385 44125 33443 44159
rect 33385 44091 33397 44125
rect 33431 44091 33443 44125
rect 33385 44057 33443 44091
rect 33385 44023 33397 44057
rect 33431 44023 33443 44057
rect 33385 43989 33443 44023
rect 33385 43955 33397 43989
rect 33431 43955 33443 43989
rect 33385 43921 33443 43955
rect 33385 43887 33397 43921
rect 33431 43887 33443 43921
rect 33385 43853 33443 43887
rect 33385 43819 33397 43853
rect 33431 43819 33443 43853
rect 33385 43785 33443 43819
rect 33385 43751 33397 43785
rect 33431 43751 33443 43785
rect 33385 43717 33443 43751
rect 33385 43683 33397 43717
rect 33431 43683 33443 43717
rect 33385 43667 33443 43683
rect 33843 44941 33901 44957
rect 33843 44907 33855 44941
rect 33889 44907 33901 44941
rect 33843 44873 33901 44907
rect 33843 44839 33855 44873
rect 33889 44839 33901 44873
rect 33843 44805 33901 44839
rect 33843 44771 33855 44805
rect 33889 44771 33901 44805
rect 33843 44737 33901 44771
rect 33843 44703 33855 44737
rect 33889 44703 33901 44737
rect 33843 44669 33901 44703
rect 33843 44635 33855 44669
rect 33889 44635 33901 44669
rect 33843 44601 33901 44635
rect 33843 44567 33855 44601
rect 33889 44567 33901 44601
rect 33843 44533 33901 44567
rect 33843 44499 33855 44533
rect 33889 44499 33901 44533
rect 33843 44465 33901 44499
rect 33843 44431 33855 44465
rect 33889 44431 33901 44465
rect 33843 44397 33901 44431
rect 33843 44363 33855 44397
rect 33889 44363 33901 44397
rect 33843 44329 33901 44363
rect 33843 44295 33855 44329
rect 33889 44295 33901 44329
rect 33843 44261 33901 44295
rect 33843 44227 33855 44261
rect 33889 44227 33901 44261
rect 33843 44193 33901 44227
rect 33843 44159 33855 44193
rect 33889 44159 33901 44193
rect 33843 44125 33901 44159
rect 33843 44091 33855 44125
rect 33889 44091 33901 44125
rect 33843 44057 33901 44091
rect 33843 44023 33855 44057
rect 33889 44023 33901 44057
rect 33843 43989 33901 44023
rect 33843 43955 33855 43989
rect 33889 43955 33901 43989
rect 33843 43921 33901 43955
rect 33843 43887 33855 43921
rect 33889 43887 33901 43921
rect 33843 43853 33901 43887
rect 33843 43819 33855 43853
rect 33889 43819 33901 43853
rect 33843 43785 33901 43819
rect 33843 43751 33855 43785
rect 33889 43751 33901 43785
rect 33843 43717 33901 43751
rect 33843 43683 33855 43717
rect 33889 43683 33901 43717
rect 33843 43667 33901 43683
rect 34301 44941 34359 44957
rect 34301 44907 34313 44941
rect 34347 44907 34359 44941
rect 34301 44873 34359 44907
rect 34301 44839 34313 44873
rect 34347 44839 34359 44873
rect 34301 44805 34359 44839
rect 34301 44771 34313 44805
rect 34347 44771 34359 44805
rect 34301 44737 34359 44771
rect 34301 44703 34313 44737
rect 34347 44703 34359 44737
rect 34301 44669 34359 44703
rect 34301 44635 34313 44669
rect 34347 44635 34359 44669
rect 34301 44601 34359 44635
rect 34301 44567 34313 44601
rect 34347 44567 34359 44601
rect 34301 44533 34359 44567
rect 34301 44499 34313 44533
rect 34347 44499 34359 44533
rect 34301 44465 34359 44499
rect 34301 44431 34313 44465
rect 34347 44431 34359 44465
rect 34301 44397 34359 44431
rect 34301 44363 34313 44397
rect 34347 44363 34359 44397
rect 34301 44329 34359 44363
rect 34301 44295 34313 44329
rect 34347 44295 34359 44329
rect 34301 44261 34359 44295
rect 34301 44227 34313 44261
rect 34347 44227 34359 44261
rect 34301 44193 34359 44227
rect 34301 44159 34313 44193
rect 34347 44159 34359 44193
rect 34301 44125 34359 44159
rect 34301 44091 34313 44125
rect 34347 44091 34359 44125
rect 34301 44057 34359 44091
rect 34301 44023 34313 44057
rect 34347 44023 34359 44057
rect 34301 43989 34359 44023
rect 34301 43955 34313 43989
rect 34347 43955 34359 43989
rect 34301 43921 34359 43955
rect 34301 43887 34313 43921
rect 34347 43887 34359 43921
rect 34301 43853 34359 43887
rect 34301 43819 34313 43853
rect 34347 43819 34359 43853
rect 34301 43785 34359 43819
rect 34301 43751 34313 43785
rect 34347 43751 34359 43785
rect 34301 43717 34359 43751
rect 34301 43683 34313 43717
rect 34347 43683 34359 43717
rect 34301 43667 34359 43683
rect 34759 44941 34817 44957
rect 34759 44907 34771 44941
rect 34805 44907 34817 44941
rect 34759 44873 34817 44907
rect 34759 44839 34771 44873
rect 34805 44839 34817 44873
rect 34759 44805 34817 44839
rect 34759 44771 34771 44805
rect 34805 44771 34817 44805
rect 34759 44737 34817 44771
rect 34759 44703 34771 44737
rect 34805 44703 34817 44737
rect 34759 44669 34817 44703
rect 34759 44635 34771 44669
rect 34805 44635 34817 44669
rect 34759 44601 34817 44635
rect 34759 44567 34771 44601
rect 34805 44567 34817 44601
rect 34759 44533 34817 44567
rect 34759 44499 34771 44533
rect 34805 44499 34817 44533
rect 34759 44465 34817 44499
rect 34759 44431 34771 44465
rect 34805 44431 34817 44465
rect 34759 44397 34817 44431
rect 34759 44363 34771 44397
rect 34805 44363 34817 44397
rect 34759 44329 34817 44363
rect 34759 44295 34771 44329
rect 34805 44295 34817 44329
rect 34759 44261 34817 44295
rect 34759 44227 34771 44261
rect 34805 44227 34817 44261
rect 34759 44193 34817 44227
rect 34759 44159 34771 44193
rect 34805 44159 34817 44193
rect 34759 44125 34817 44159
rect 34759 44091 34771 44125
rect 34805 44091 34817 44125
rect 34759 44057 34817 44091
rect 34759 44023 34771 44057
rect 34805 44023 34817 44057
rect 34759 43989 34817 44023
rect 34759 43955 34771 43989
rect 34805 43955 34817 43989
rect 34759 43921 34817 43955
rect 34759 43887 34771 43921
rect 34805 43887 34817 43921
rect 34759 43853 34817 43887
rect 34759 43819 34771 43853
rect 34805 43819 34817 43853
rect 34759 43785 34817 43819
rect 34759 43751 34771 43785
rect 34805 43751 34817 43785
rect 34759 43717 34817 43751
rect 34759 43683 34771 43717
rect 34805 43683 34817 43717
rect 34759 43667 34817 43683
rect 35217 44941 35275 44957
rect 35217 44907 35229 44941
rect 35263 44907 35275 44941
rect 35217 44873 35275 44907
rect 35217 44839 35229 44873
rect 35263 44839 35275 44873
rect 35217 44805 35275 44839
rect 35217 44771 35229 44805
rect 35263 44771 35275 44805
rect 35217 44737 35275 44771
rect 35217 44703 35229 44737
rect 35263 44703 35275 44737
rect 35217 44669 35275 44703
rect 35217 44635 35229 44669
rect 35263 44635 35275 44669
rect 35217 44601 35275 44635
rect 35217 44567 35229 44601
rect 35263 44567 35275 44601
rect 35217 44533 35275 44567
rect 35217 44499 35229 44533
rect 35263 44499 35275 44533
rect 35217 44465 35275 44499
rect 35217 44431 35229 44465
rect 35263 44431 35275 44465
rect 35217 44397 35275 44431
rect 35217 44363 35229 44397
rect 35263 44363 35275 44397
rect 35217 44329 35275 44363
rect 35217 44295 35229 44329
rect 35263 44295 35275 44329
rect 35217 44261 35275 44295
rect 35217 44227 35229 44261
rect 35263 44227 35275 44261
rect 35217 44193 35275 44227
rect 35217 44159 35229 44193
rect 35263 44159 35275 44193
rect 35217 44125 35275 44159
rect 35217 44091 35229 44125
rect 35263 44091 35275 44125
rect 35217 44057 35275 44091
rect 35217 44023 35229 44057
rect 35263 44023 35275 44057
rect 35217 43989 35275 44023
rect 35217 43955 35229 43989
rect 35263 43955 35275 43989
rect 35217 43921 35275 43955
rect 35217 43887 35229 43921
rect 35263 43887 35275 43921
rect 35217 43853 35275 43887
rect 35217 43819 35229 43853
rect 35263 43819 35275 43853
rect 35217 43785 35275 43819
rect 35217 43751 35229 43785
rect 35263 43751 35275 43785
rect 35217 43717 35275 43751
rect 35217 43683 35229 43717
rect 35263 43683 35275 43717
rect 35217 43667 35275 43683
rect 35675 44941 35733 44957
rect 35675 44907 35687 44941
rect 35721 44907 35733 44941
rect 35675 44873 35733 44907
rect 35675 44839 35687 44873
rect 35721 44839 35733 44873
rect 35675 44805 35733 44839
rect 35675 44771 35687 44805
rect 35721 44771 35733 44805
rect 35675 44737 35733 44771
rect 35675 44703 35687 44737
rect 35721 44703 35733 44737
rect 35675 44669 35733 44703
rect 35675 44635 35687 44669
rect 35721 44635 35733 44669
rect 35675 44601 35733 44635
rect 35675 44567 35687 44601
rect 35721 44567 35733 44601
rect 35675 44533 35733 44567
rect 35675 44499 35687 44533
rect 35721 44499 35733 44533
rect 35675 44465 35733 44499
rect 35675 44431 35687 44465
rect 35721 44431 35733 44465
rect 35675 44397 35733 44431
rect 35675 44363 35687 44397
rect 35721 44363 35733 44397
rect 35675 44329 35733 44363
rect 35675 44295 35687 44329
rect 35721 44295 35733 44329
rect 35675 44261 35733 44295
rect 35675 44227 35687 44261
rect 35721 44227 35733 44261
rect 35675 44193 35733 44227
rect 35675 44159 35687 44193
rect 35721 44159 35733 44193
rect 35675 44125 35733 44159
rect 35675 44091 35687 44125
rect 35721 44091 35733 44125
rect 35675 44057 35733 44091
rect 35675 44023 35687 44057
rect 35721 44023 35733 44057
rect 35675 43989 35733 44023
rect 35675 43955 35687 43989
rect 35721 43955 35733 43989
rect 35675 43921 35733 43955
rect 35675 43887 35687 43921
rect 35721 43887 35733 43921
rect 35675 43853 35733 43887
rect 35675 43819 35687 43853
rect 35721 43819 35733 43853
rect 35675 43785 35733 43819
rect 35675 43751 35687 43785
rect 35721 43751 35733 43785
rect 35675 43717 35733 43751
rect 35675 43683 35687 43717
rect 35721 43683 35733 43717
rect 35675 43667 35733 43683
rect 36133 44941 36191 44957
rect 36133 44907 36145 44941
rect 36179 44907 36191 44941
rect 36133 44873 36191 44907
rect 36133 44839 36145 44873
rect 36179 44839 36191 44873
rect 36133 44805 36191 44839
rect 36133 44771 36145 44805
rect 36179 44771 36191 44805
rect 36133 44737 36191 44771
rect 36133 44703 36145 44737
rect 36179 44703 36191 44737
rect 36133 44669 36191 44703
rect 36133 44635 36145 44669
rect 36179 44635 36191 44669
rect 36133 44601 36191 44635
rect 36133 44567 36145 44601
rect 36179 44567 36191 44601
rect 36133 44533 36191 44567
rect 36133 44499 36145 44533
rect 36179 44499 36191 44533
rect 36133 44465 36191 44499
rect 36133 44431 36145 44465
rect 36179 44431 36191 44465
rect 36133 44397 36191 44431
rect 36133 44363 36145 44397
rect 36179 44363 36191 44397
rect 36133 44329 36191 44363
rect 36133 44295 36145 44329
rect 36179 44295 36191 44329
rect 36133 44261 36191 44295
rect 36133 44227 36145 44261
rect 36179 44227 36191 44261
rect 36133 44193 36191 44227
rect 36133 44159 36145 44193
rect 36179 44159 36191 44193
rect 36133 44125 36191 44159
rect 36133 44091 36145 44125
rect 36179 44091 36191 44125
rect 36133 44057 36191 44091
rect 36133 44023 36145 44057
rect 36179 44023 36191 44057
rect 36133 43989 36191 44023
rect 36133 43955 36145 43989
rect 36179 43955 36191 43989
rect 36133 43921 36191 43955
rect 36133 43887 36145 43921
rect 36179 43887 36191 43921
rect 36133 43853 36191 43887
rect 36133 43819 36145 43853
rect 36179 43819 36191 43853
rect 36133 43785 36191 43819
rect 36133 43751 36145 43785
rect 36179 43751 36191 43785
rect 36133 43717 36191 43751
rect 36133 43683 36145 43717
rect 36179 43683 36191 43717
rect 36133 43667 36191 43683
rect 36591 44941 36649 44957
rect 36591 44907 36603 44941
rect 36637 44907 36649 44941
rect 36591 44873 36649 44907
rect 36591 44839 36603 44873
rect 36637 44839 36649 44873
rect 36591 44805 36649 44839
rect 36591 44771 36603 44805
rect 36637 44771 36649 44805
rect 36591 44737 36649 44771
rect 36591 44703 36603 44737
rect 36637 44703 36649 44737
rect 36591 44669 36649 44703
rect 36591 44635 36603 44669
rect 36637 44635 36649 44669
rect 36591 44601 36649 44635
rect 36591 44567 36603 44601
rect 36637 44567 36649 44601
rect 36591 44533 36649 44567
rect 36591 44499 36603 44533
rect 36637 44499 36649 44533
rect 36591 44465 36649 44499
rect 36591 44431 36603 44465
rect 36637 44431 36649 44465
rect 36591 44397 36649 44431
rect 36591 44363 36603 44397
rect 36637 44363 36649 44397
rect 36591 44329 36649 44363
rect 36591 44295 36603 44329
rect 36637 44295 36649 44329
rect 36591 44261 36649 44295
rect 36591 44227 36603 44261
rect 36637 44227 36649 44261
rect 36591 44193 36649 44227
rect 36591 44159 36603 44193
rect 36637 44159 36649 44193
rect 36591 44125 36649 44159
rect 36591 44091 36603 44125
rect 36637 44091 36649 44125
rect 36591 44057 36649 44091
rect 36591 44023 36603 44057
rect 36637 44023 36649 44057
rect 36591 43989 36649 44023
rect 36591 43955 36603 43989
rect 36637 43955 36649 43989
rect 36591 43921 36649 43955
rect 36591 43887 36603 43921
rect 36637 43887 36649 43921
rect 36591 43853 36649 43887
rect 36591 43819 36603 43853
rect 36637 43819 36649 43853
rect 36591 43785 36649 43819
rect 36591 43751 36603 43785
rect 36637 43751 36649 43785
rect 36591 43717 36649 43751
rect 36591 43683 36603 43717
rect 36637 43683 36649 43717
rect 36591 43667 36649 43683
rect 37049 44941 37107 44957
rect 37049 44907 37061 44941
rect 37095 44907 37107 44941
rect 37049 44873 37107 44907
rect 37049 44839 37061 44873
rect 37095 44839 37107 44873
rect 37049 44805 37107 44839
rect 37049 44771 37061 44805
rect 37095 44771 37107 44805
rect 37049 44737 37107 44771
rect 37049 44703 37061 44737
rect 37095 44703 37107 44737
rect 37049 44669 37107 44703
rect 37049 44635 37061 44669
rect 37095 44635 37107 44669
rect 37049 44601 37107 44635
rect 37049 44567 37061 44601
rect 37095 44567 37107 44601
rect 37049 44533 37107 44567
rect 37049 44499 37061 44533
rect 37095 44499 37107 44533
rect 37049 44465 37107 44499
rect 37049 44431 37061 44465
rect 37095 44431 37107 44465
rect 37049 44397 37107 44431
rect 37049 44363 37061 44397
rect 37095 44363 37107 44397
rect 37049 44329 37107 44363
rect 37049 44295 37061 44329
rect 37095 44295 37107 44329
rect 37049 44261 37107 44295
rect 37049 44227 37061 44261
rect 37095 44227 37107 44261
rect 37049 44193 37107 44227
rect 37049 44159 37061 44193
rect 37095 44159 37107 44193
rect 37049 44125 37107 44159
rect 37049 44091 37061 44125
rect 37095 44091 37107 44125
rect 37049 44057 37107 44091
rect 37049 44023 37061 44057
rect 37095 44023 37107 44057
rect 37049 43989 37107 44023
rect 37049 43955 37061 43989
rect 37095 43955 37107 43989
rect 37049 43921 37107 43955
rect 37049 43887 37061 43921
rect 37095 43887 37107 43921
rect 37049 43853 37107 43887
rect 37049 43819 37061 43853
rect 37095 43819 37107 43853
rect 37049 43785 37107 43819
rect 37049 43751 37061 43785
rect 37095 43751 37107 43785
rect 37049 43717 37107 43751
rect 37049 43683 37061 43717
rect 37095 43683 37107 43717
rect 37049 43667 37107 43683
rect 37507 44941 37565 44957
rect 37507 44907 37519 44941
rect 37553 44907 37565 44941
rect 37507 44873 37565 44907
rect 37507 44839 37519 44873
rect 37553 44839 37565 44873
rect 37507 44805 37565 44839
rect 37507 44771 37519 44805
rect 37553 44771 37565 44805
rect 37507 44737 37565 44771
rect 37507 44703 37519 44737
rect 37553 44703 37565 44737
rect 37507 44669 37565 44703
rect 37507 44635 37519 44669
rect 37553 44635 37565 44669
rect 37507 44601 37565 44635
rect 37507 44567 37519 44601
rect 37553 44567 37565 44601
rect 37507 44533 37565 44567
rect 37507 44499 37519 44533
rect 37553 44499 37565 44533
rect 37507 44465 37565 44499
rect 37507 44431 37519 44465
rect 37553 44431 37565 44465
rect 37507 44397 37565 44431
rect 37507 44363 37519 44397
rect 37553 44363 37565 44397
rect 37507 44329 37565 44363
rect 37507 44295 37519 44329
rect 37553 44295 37565 44329
rect 37507 44261 37565 44295
rect 37507 44227 37519 44261
rect 37553 44227 37565 44261
rect 37507 44193 37565 44227
rect 37507 44159 37519 44193
rect 37553 44159 37565 44193
rect 37507 44125 37565 44159
rect 37507 44091 37519 44125
rect 37553 44091 37565 44125
rect 37507 44057 37565 44091
rect 37507 44023 37519 44057
rect 37553 44023 37565 44057
rect 37507 43989 37565 44023
rect 37507 43955 37519 43989
rect 37553 43955 37565 43989
rect 37507 43921 37565 43955
rect 37507 43887 37519 43921
rect 37553 43887 37565 43921
rect 37507 43853 37565 43887
rect 37507 43819 37519 43853
rect 37553 43819 37565 43853
rect 37507 43785 37565 43819
rect 37507 43751 37519 43785
rect 37553 43751 37565 43785
rect 37507 43717 37565 43751
rect 37507 43683 37519 43717
rect 37553 43683 37565 43717
rect 37507 43667 37565 43683
rect 37965 44941 38023 44957
rect 37965 44907 37977 44941
rect 38011 44907 38023 44941
rect 37965 44873 38023 44907
rect 37965 44839 37977 44873
rect 38011 44839 38023 44873
rect 37965 44805 38023 44839
rect 37965 44771 37977 44805
rect 38011 44771 38023 44805
rect 37965 44737 38023 44771
rect 37965 44703 37977 44737
rect 38011 44703 38023 44737
rect 37965 44669 38023 44703
rect 37965 44635 37977 44669
rect 38011 44635 38023 44669
rect 37965 44601 38023 44635
rect 37965 44567 37977 44601
rect 38011 44567 38023 44601
rect 37965 44533 38023 44567
rect 37965 44499 37977 44533
rect 38011 44499 38023 44533
rect 37965 44465 38023 44499
rect 37965 44431 37977 44465
rect 38011 44431 38023 44465
rect 37965 44397 38023 44431
rect 37965 44363 37977 44397
rect 38011 44363 38023 44397
rect 37965 44329 38023 44363
rect 37965 44295 37977 44329
rect 38011 44295 38023 44329
rect 37965 44261 38023 44295
rect 37965 44227 37977 44261
rect 38011 44227 38023 44261
rect 37965 44193 38023 44227
rect 37965 44159 37977 44193
rect 38011 44159 38023 44193
rect 37965 44125 38023 44159
rect 37965 44091 37977 44125
rect 38011 44091 38023 44125
rect 37965 44057 38023 44091
rect 37965 44023 37977 44057
rect 38011 44023 38023 44057
rect 37965 43989 38023 44023
rect 37965 43955 37977 43989
rect 38011 43955 38023 43989
rect 37965 43921 38023 43955
rect 37965 43887 37977 43921
rect 38011 43887 38023 43921
rect 37965 43853 38023 43887
rect 37965 43819 37977 43853
rect 38011 43819 38023 43853
rect 37965 43785 38023 43819
rect 37965 43751 37977 43785
rect 38011 43751 38023 43785
rect 37965 43717 38023 43751
rect 37965 43683 37977 43717
rect 38011 43683 38023 43717
rect 37965 43667 38023 43683
rect 38423 44941 38481 44957
rect 38423 44907 38435 44941
rect 38469 44907 38481 44941
rect 38423 44873 38481 44907
rect 38423 44839 38435 44873
rect 38469 44839 38481 44873
rect 38423 44805 38481 44839
rect 38423 44771 38435 44805
rect 38469 44771 38481 44805
rect 38423 44737 38481 44771
rect 38423 44703 38435 44737
rect 38469 44703 38481 44737
rect 38423 44669 38481 44703
rect 38423 44635 38435 44669
rect 38469 44635 38481 44669
rect 38423 44601 38481 44635
rect 38423 44567 38435 44601
rect 38469 44567 38481 44601
rect 38423 44533 38481 44567
rect 38423 44499 38435 44533
rect 38469 44499 38481 44533
rect 38423 44465 38481 44499
rect 38423 44431 38435 44465
rect 38469 44431 38481 44465
rect 38423 44397 38481 44431
rect 38423 44363 38435 44397
rect 38469 44363 38481 44397
rect 38423 44329 38481 44363
rect 38423 44295 38435 44329
rect 38469 44295 38481 44329
rect 38423 44261 38481 44295
rect 38423 44227 38435 44261
rect 38469 44227 38481 44261
rect 38423 44193 38481 44227
rect 38423 44159 38435 44193
rect 38469 44159 38481 44193
rect 38423 44125 38481 44159
rect 38423 44091 38435 44125
rect 38469 44091 38481 44125
rect 38423 44057 38481 44091
rect 38423 44023 38435 44057
rect 38469 44023 38481 44057
rect 38423 43989 38481 44023
rect 38423 43955 38435 43989
rect 38469 43955 38481 43989
rect 38423 43921 38481 43955
rect 38423 43887 38435 43921
rect 38469 43887 38481 43921
rect 38423 43853 38481 43887
rect 38423 43819 38435 43853
rect 38469 43819 38481 43853
rect 38423 43785 38481 43819
rect 38423 43751 38435 43785
rect 38469 43751 38481 43785
rect 38423 43717 38481 43751
rect 38423 43683 38435 43717
rect 38469 43683 38481 43717
rect 38423 43667 38481 43683
rect 38881 44941 38939 44957
rect 38881 44907 38893 44941
rect 38927 44907 38939 44941
rect 38881 44873 38939 44907
rect 38881 44839 38893 44873
rect 38927 44839 38939 44873
rect 38881 44805 38939 44839
rect 38881 44771 38893 44805
rect 38927 44771 38939 44805
rect 38881 44737 38939 44771
rect 38881 44703 38893 44737
rect 38927 44703 38939 44737
rect 38881 44669 38939 44703
rect 38881 44635 38893 44669
rect 38927 44635 38939 44669
rect 38881 44601 38939 44635
rect 38881 44567 38893 44601
rect 38927 44567 38939 44601
rect 38881 44533 38939 44567
rect 38881 44499 38893 44533
rect 38927 44499 38939 44533
rect 38881 44465 38939 44499
rect 38881 44431 38893 44465
rect 38927 44431 38939 44465
rect 38881 44397 38939 44431
rect 38881 44363 38893 44397
rect 38927 44363 38939 44397
rect 38881 44329 38939 44363
rect 38881 44295 38893 44329
rect 38927 44295 38939 44329
rect 38881 44261 38939 44295
rect 38881 44227 38893 44261
rect 38927 44227 38939 44261
rect 38881 44193 38939 44227
rect 38881 44159 38893 44193
rect 38927 44159 38939 44193
rect 38881 44125 38939 44159
rect 38881 44091 38893 44125
rect 38927 44091 38939 44125
rect 38881 44057 38939 44091
rect 38881 44023 38893 44057
rect 38927 44023 38939 44057
rect 38881 43989 38939 44023
rect 38881 43955 38893 43989
rect 38927 43955 38939 43989
rect 38881 43921 38939 43955
rect 38881 43887 38893 43921
rect 38927 43887 38939 43921
rect 38881 43853 38939 43887
rect 38881 43819 38893 43853
rect 38927 43819 38939 43853
rect 38881 43785 38939 43819
rect 38881 43751 38893 43785
rect 38927 43751 38939 43785
rect 38881 43717 38939 43751
rect 38881 43683 38893 43717
rect 38927 43683 38939 43717
rect 38881 43667 38939 43683
rect 39339 44941 39397 44957
rect 39339 44907 39351 44941
rect 39385 44907 39397 44941
rect 39339 44873 39397 44907
rect 39339 44839 39351 44873
rect 39385 44839 39397 44873
rect 39339 44805 39397 44839
rect 39339 44771 39351 44805
rect 39385 44771 39397 44805
rect 39339 44737 39397 44771
rect 39339 44703 39351 44737
rect 39385 44703 39397 44737
rect 39339 44669 39397 44703
rect 39339 44635 39351 44669
rect 39385 44635 39397 44669
rect 39339 44601 39397 44635
rect 39339 44567 39351 44601
rect 39385 44567 39397 44601
rect 39339 44533 39397 44567
rect 39339 44499 39351 44533
rect 39385 44499 39397 44533
rect 39339 44465 39397 44499
rect 39339 44431 39351 44465
rect 39385 44431 39397 44465
rect 39339 44397 39397 44431
rect 39339 44363 39351 44397
rect 39385 44363 39397 44397
rect 39339 44329 39397 44363
rect 39339 44295 39351 44329
rect 39385 44295 39397 44329
rect 39339 44261 39397 44295
rect 39339 44227 39351 44261
rect 39385 44227 39397 44261
rect 39339 44193 39397 44227
rect 39339 44159 39351 44193
rect 39385 44159 39397 44193
rect 39339 44125 39397 44159
rect 39339 44091 39351 44125
rect 39385 44091 39397 44125
rect 39339 44057 39397 44091
rect 39339 44023 39351 44057
rect 39385 44023 39397 44057
rect 39339 43989 39397 44023
rect 39339 43955 39351 43989
rect 39385 43955 39397 43989
rect 39339 43921 39397 43955
rect 39339 43887 39351 43921
rect 39385 43887 39397 43921
rect 39339 43853 39397 43887
rect 39339 43819 39351 43853
rect 39385 43819 39397 43853
rect 39339 43785 39397 43819
rect 39339 43751 39351 43785
rect 39385 43751 39397 43785
rect 39339 43717 39397 43751
rect 39339 43683 39351 43717
rect 39385 43683 39397 43717
rect 39339 43667 39397 43683
rect 39797 44941 39855 44957
rect 39797 44907 39809 44941
rect 39843 44907 39855 44941
rect 39797 44873 39855 44907
rect 39797 44839 39809 44873
rect 39843 44839 39855 44873
rect 39797 44805 39855 44839
rect 39797 44771 39809 44805
rect 39843 44771 39855 44805
rect 39797 44737 39855 44771
rect 39797 44703 39809 44737
rect 39843 44703 39855 44737
rect 39797 44669 39855 44703
rect 39797 44635 39809 44669
rect 39843 44635 39855 44669
rect 39797 44601 39855 44635
rect 39797 44567 39809 44601
rect 39843 44567 39855 44601
rect 39797 44533 39855 44567
rect 39797 44499 39809 44533
rect 39843 44499 39855 44533
rect 39797 44465 39855 44499
rect 39797 44431 39809 44465
rect 39843 44431 39855 44465
rect 39797 44397 39855 44431
rect 39797 44363 39809 44397
rect 39843 44363 39855 44397
rect 39797 44329 39855 44363
rect 39797 44295 39809 44329
rect 39843 44295 39855 44329
rect 39797 44261 39855 44295
rect 39797 44227 39809 44261
rect 39843 44227 39855 44261
rect 39797 44193 39855 44227
rect 39797 44159 39809 44193
rect 39843 44159 39855 44193
rect 39797 44125 39855 44159
rect 39797 44091 39809 44125
rect 39843 44091 39855 44125
rect 39797 44057 39855 44091
rect 39797 44023 39809 44057
rect 39843 44023 39855 44057
rect 39797 43989 39855 44023
rect 39797 43955 39809 43989
rect 39843 43955 39855 43989
rect 39797 43921 39855 43955
rect 39797 43887 39809 43921
rect 39843 43887 39855 43921
rect 39797 43853 39855 43887
rect 39797 43819 39809 43853
rect 39843 43819 39855 43853
rect 39797 43785 39855 43819
rect 39797 43751 39809 43785
rect 39843 43751 39855 43785
rect 39797 43717 39855 43751
rect 39797 43683 39809 43717
rect 39843 43683 39855 43717
rect 39797 43667 39855 43683
rect 40255 44941 40313 44957
rect 40255 44907 40267 44941
rect 40301 44907 40313 44941
rect 40255 44873 40313 44907
rect 40255 44839 40267 44873
rect 40301 44839 40313 44873
rect 40255 44805 40313 44839
rect 40255 44771 40267 44805
rect 40301 44771 40313 44805
rect 40255 44737 40313 44771
rect 40255 44703 40267 44737
rect 40301 44703 40313 44737
rect 40255 44669 40313 44703
rect 40255 44635 40267 44669
rect 40301 44635 40313 44669
rect 40255 44601 40313 44635
rect 40255 44567 40267 44601
rect 40301 44567 40313 44601
rect 40255 44533 40313 44567
rect 40255 44499 40267 44533
rect 40301 44499 40313 44533
rect 40255 44465 40313 44499
rect 40255 44431 40267 44465
rect 40301 44431 40313 44465
rect 40255 44397 40313 44431
rect 40255 44363 40267 44397
rect 40301 44363 40313 44397
rect 40255 44329 40313 44363
rect 40255 44295 40267 44329
rect 40301 44295 40313 44329
rect 40255 44261 40313 44295
rect 40255 44227 40267 44261
rect 40301 44227 40313 44261
rect 40255 44193 40313 44227
rect 40255 44159 40267 44193
rect 40301 44159 40313 44193
rect 40255 44125 40313 44159
rect 40255 44091 40267 44125
rect 40301 44091 40313 44125
rect 40255 44057 40313 44091
rect 40255 44023 40267 44057
rect 40301 44023 40313 44057
rect 40255 43989 40313 44023
rect 40255 43955 40267 43989
rect 40301 43955 40313 43989
rect 40255 43921 40313 43955
rect 40255 43887 40267 43921
rect 40301 43887 40313 43921
rect 40255 43853 40313 43887
rect 40255 43819 40267 43853
rect 40301 43819 40313 43853
rect 40255 43785 40313 43819
rect 40255 43751 40267 43785
rect 40301 43751 40313 43785
rect 40255 43717 40313 43751
rect 40255 43683 40267 43717
rect 40301 43683 40313 43717
rect 40255 43667 40313 43683
rect 40713 44941 40771 44957
rect 40713 44907 40725 44941
rect 40759 44907 40771 44941
rect 40713 44873 40771 44907
rect 40713 44839 40725 44873
rect 40759 44839 40771 44873
rect 40713 44805 40771 44839
rect 40713 44771 40725 44805
rect 40759 44771 40771 44805
rect 40713 44737 40771 44771
rect 40713 44703 40725 44737
rect 40759 44703 40771 44737
rect 40713 44669 40771 44703
rect 40713 44635 40725 44669
rect 40759 44635 40771 44669
rect 40713 44601 40771 44635
rect 40713 44567 40725 44601
rect 40759 44567 40771 44601
rect 40713 44533 40771 44567
rect 40713 44499 40725 44533
rect 40759 44499 40771 44533
rect 40713 44465 40771 44499
rect 40713 44431 40725 44465
rect 40759 44431 40771 44465
rect 40713 44397 40771 44431
rect 40713 44363 40725 44397
rect 40759 44363 40771 44397
rect 40713 44329 40771 44363
rect 40713 44295 40725 44329
rect 40759 44295 40771 44329
rect 40713 44261 40771 44295
rect 40713 44227 40725 44261
rect 40759 44227 40771 44261
rect 40713 44193 40771 44227
rect 40713 44159 40725 44193
rect 40759 44159 40771 44193
rect 40713 44125 40771 44159
rect 40713 44091 40725 44125
rect 40759 44091 40771 44125
rect 40713 44057 40771 44091
rect 40713 44023 40725 44057
rect 40759 44023 40771 44057
rect 40713 43989 40771 44023
rect 40713 43955 40725 43989
rect 40759 43955 40771 43989
rect 40713 43921 40771 43955
rect 40713 43887 40725 43921
rect 40759 43887 40771 43921
rect 40713 43853 40771 43887
rect 40713 43819 40725 43853
rect 40759 43819 40771 43853
rect 40713 43785 40771 43819
rect 40713 43751 40725 43785
rect 40759 43751 40771 43785
rect 40713 43717 40771 43751
rect 40713 43683 40725 43717
rect 40759 43683 40771 43717
rect 40713 43667 40771 43683
rect 41171 44941 41229 44957
rect 41171 44907 41183 44941
rect 41217 44907 41229 44941
rect 41171 44873 41229 44907
rect 41171 44839 41183 44873
rect 41217 44839 41229 44873
rect 41171 44805 41229 44839
rect 41171 44771 41183 44805
rect 41217 44771 41229 44805
rect 41171 44737 41229 44771
rect 41171 44703 41183 44737
rect 41217 44703 41229 44737
rect 41171 44669 41229 44703
rect 41171 44635 41183 44669
rect 41217 44635 41229 44669
rect 41171 44601 41229 44635
rect 41171 44567 41183 44601
rect 41217 44567 41229 44601
rect 41171 44533 41229 44567
rect 41171 44499 41183 44533
rect 41217 44499 41229 44533
rect 41171 44465 41229 44499
rect 41171 44431 41183 44465
rect 41217 44431 41229 44465
rect 41171 44397 41229 44431
rect 41171 44363 41183 44397
rect 41217 44363 41229 44397
rect 41171 44329 41229 44363
rect 41171 44295 41183 44329
rect 41217 44295 41229 44329
rect 41171 44261 41229 44295
rect 41171 44227 41183 44261
rect 41217 44227 41229 44261
rect 41171 44193 41229 44227
rect 41171 44159 41183 44193
rect 41217 44159 41229 44193
rect 41171 44125 41229 44159
rect 41171 44091 41183 44125
rect 41217 44091 41229 44125
rect 41171 44057 41229 44091
rect 41171 44023 41183 44057
rect 41217 44023 41229 44057
rect 41171 43989 41229 44023
rect 41171 43955 41183 43989
rect 41217 43955 41229 43989
rect 41171 43921 41229 43955
rect 41171 43887 41183 43921
rect 41217 43887 41229 43921
rect 41171 43853 41229 43887
rect 41171 43819 41183 43853
rect 41217 43819 41229 43853
rect 41171 43785 41229 43819
rect 41171 43751 41183 43785
rect 41217 43751 41229 43785
rect 41171 43717 41229 43751
rect 41171 43683 41183 43717
rect 41217 43683 41229 43717
rect 41171 43667 41229 43683
rect 41629 44941 41687 44957
rect 41629 44907 41641 44941
rect 41675 44907 41687 44941
rect 41629 44873 41687 44907
rect 41629 44839 41641 44873
rect 41675 44839 41687 44873
rect 41629 44805 41687 44839
rect 41629 44771 41641 44805
rect 41675 44771 41687 44805
rect 41629 44737 41687 44771
rect 41629 44703 41641 44737
rect 41675 44703 41687 44737
rect 41629 44669 41687 44703
rect 41629 44635 41641 44669
rect 41675 44635 41687 44669
rect 41629 44601 41687 44635
rect 41629 44567 41641 44601
rect 41675 44567 41687 44601
rect 41629 44533 41687 44567
rect 41629 44499 41641 44533
rect 41675 44499 41687 44533
rect 41629 44465 41687 44499
rect 41629 44431 41641 44465
rect 41675 44431 41687 44465
rect 41629 44397 41687 44431
rect 41629 44363 41641 44397
rect 41675 44363 41687 44397
rect 41629 44329 41687 44363
rect 41629 44295 41641 44329
rect 41675 44295 41687 44329
rect 41629 44261 41687 44295
rect 41629 44227 41641 44261
rect 41675 44227 41687 44261
rect 41629 44193 41687 44227
rect 41629 44159 41641 44193
rect 41675 44159 41687 44193
rect 41629 44125 41687 44159
rect 41629 44091 41641 44125
rect 41675 44091 41687 44125
rect 41629 44057 41687 44091
rect 41629 44023 41641 44057
rect 41675 44023 41687 44057
rect 41629 43989 41687 44023
rect 41629 43955 41641 43989
rect 41675 43955 41687 43989
rect 41629 43921 41687 43955
rect 41629 43887 41641 43921
rect 41675 43887 41687 43921
rect 41629 43853 41687 43887
rect 41629 43819 41641 43853
rect 41675 43819 41687 43853
rect 41629 43785 41687 43819
rect 41629 43751 41641 43785
rect 41675 43751 41687 43785
rect 41629 43717 41687 43751
rect 41629 43683 41641 43717
rect 41675 43683 41687 43717
rect 41629 43667 41687 43683
rect 42087 44941 42145 44957
rect 42087 44907 42099 44941
rect 42133 44907 42145 44941
rect 42087 44873 42145 44907
rect 42087 44839 42099 44873
rect 42133 44839 42145 44873
rect 42087 44805 42145 44839
rect 42087 44771 42099 44805
rect 42133 44771 42145 44805
rect 42087 44737 42145 44771
rect 42087 44703 42099 44737
rect 42133 44703 42145 44737
rect 42087 44669 42145 44703
rect 42087 44635 42099 44669
rect 42133 44635 42145 44669
rect 42087 44601 42145 44635
rect 42087 44567 42099 44601
rect 42133 44567 42145 44601
rect 42087 44533 42145 44567
rect 42087 44499 42099 44533
rect 42133 44499 42145 44533
rect 42087 44465 42145 44499
rect 42087 44431 42099 44465
rect 42133 44431 42145 44465
rect 42087 44397 42145 44431
rect 42087 44363 42099 44397
rect 42133 44363 42145 44397
rect 42087 44329 42145 44363
rect 42087 44295 42099 44329
rect 42133 44295 42145 44329
rect 42087 44261 42145 44295
rect 42087 44227 42099 44261
rect 42133 44227 42145 44261
rect 42087 44193 42145 44227
rect 42087 44159 42099 44193
rect 42133 44159 42145 44193
rect 42087 44125 42145 44159
rect 42087 44091 42099 44125
rect 42133 44091 42145 44125
rect 42087 44057 42145 44091
rect 42087 44023 42099 44057
rect 42133 44023 42145 44057
rect 42087 43989 42145 44023
rect 42087 43955 42099 43989
rect 42133 43955 42145 43989
rect 42087 43921 42145 43955
rect 42087 43887 42099 43921
rect 42133 43887 42145 43921
rect 42087 43853 42145 43887
rect 42087 43819 42099 43853
rect 42133 43819 42145 43853
rect 42087 43785 42145 43819
rect 42087 43751 42099 43785
rect 42133 43751 42145 43785
rect 42087 43717 42145 43751
rect 42087 43683 42099 43717
rect 42133 43683 42145 43717
rect 42087 43667 42145 43683
rect 42545 44941 42603 44957
rect 42545 44907 42557 44941
rect 42591 44907 42603 44941
rect 42545 44873 42603 44907
rect 42545 44839 42557 44873
rect 42591 44839 42603 44873
rect 42545 44805 42603 44839
rect 42545 44771 42557 44805
rect 42591 44771 42603 44805
rect 42545 44737 42603 44771
rect 42545 44703 42557 44737
rect 42591 44703 42603 44737
rect 42545 44669 42603 44703
rect 42545 44635 42557 44669
rect 42591 44635 42603 44669
rect 42545 44601 42603 44635
rect 42545 44567 42557 44601
rect 42591 44567 42603 44601
rect 42545 44533 42603 44567
rect 42545 44499 42557 44533
rect 42591 44499 42603 44533
rect 42545 44465 42603 44499
rect 42545 44431 42557 44465
rect 42591 44431 42603 44465
rect 42545 44397 42603 44431
rect 42545 44363 42557 44397
rect 42591 44363 42603 44397
rect 42545 44329 42603 44363
rect 42545 44295 42557 44329
rect 42591 44295 42603 44329
rect 42545 44261 42603 44295
rect 42545 44227 42557 44261
rect 42591 44227 42603 44261
rect 42545 44193 42603 44227
rect 42545 44159 42557 44193
rect 42591 44159 42603 44193
rect 42545 44125 42603 44159
rect 42545 44091 42557 44125
rect 42591 44091 42603 44125
rect 42545 44057 42603 44091
rect 42545 44023 42557 44057
rect 42591 44023 42603 44057
rect 42545 43989 42603 44023
rect 42545 43955 42557 43989
rect 42591 43955 42603 43989
rect 42545 43921 42603 43955
rect 42545 43887 42557 43921
rect 42591 43887 42603 43921
rect 42545 43853 42603 43887
rect 42545 43819 42557 43853
rect 42591 43819 42603 43853
rect 42545 43785 42603 43819
rect 42545 43751 42557 43785
rect 42591 43751 42603 43785
rect 42545 43717 42603 43751
rect 42545 43683 42557 43717
rect 42591 43683 42603 43717
rect 42545 43667 42603 43683
rect 43290 44540 43970 44592
rect 43290 44506 43344 44540
rect 43378 44506 43434 44540
rect 43468 44506 43524 44540
rect 43558 44506 43614 44540
rect 43648 44506 43704 44540
rect 43738 44506 43794 44540
rect 43828 44506 43884 44540
rect 43918 44506 43970 44540
rect 43290 44450 43970 44506
rect 43290 44416 43344 44450
rect 43378 44416 43434 44450
rect 43468 44416 43524 44450
rect 43558 44416 43614 44450
rect 43648 44416 43704 44450
rect 43738 44416 43794 44450
rect 43828 44416 43884 44450
rect 43918 44416 43970 44450
rect 43290 44360 43970 44416
rect 43290 44326 43344 44360
rect 43378 44326 43434 44360
rect 43468 44326 43524 44360
rect 43558 44326 43614 44360
rect 43648 44326 43704 44360
rect 43738 44326 43794 44360
rect 43828 44326 43884 44360
rect 43918 44326 43970 44360
rect 43290 44270 43970 44326
rect 43290 44236 43344 44270
rect 43378 44236 43434 44270
rect 43468 44236 43524 44270
rect 43558 44236 43614 44270
rect 43648 44236 43704 44270
rect 43738 44236 43794 44270
rect 43828 44236 43884 44270
rect 43918 44236 43970 44270
rect 43290 44180 43970 44236
rect 43290 44146 43344 44180
rect 43378 44146 43434 44180
rect 43468 44146 43524 44180
rect 43558 44146 43614 44180
rect 43648 44146 43704 44180
rect 43738 44146 43794 44180
rect 43828 44146 43884 44180
rect 43918 44146 43970 44180
rect 43290 44090 43970 44146
rect 43290 44056 43344 44090
rect 43378 44056 43434 44090
rect 43468 44056 43524 44090
rect 43558 44056 43614 44090
rect 43648 44056 43704 44090
rect 43738 44056 43794 44090
rect 43828 44056 43884 44090
rect 43918 44056 43970 44090
rect 43290 44000 43970 44056
rect 43290 43966 43344 44000
rect 43378 43966 43434 44000
rect 43468 43966 43524 44000
rect 43558 43966 43614 44000
rect 43648 43966 43704 44000
rect 43738 43966 43794 44000
rect 43828 43966 43884 44000
rect 43918 43966 43970 44000
rect 43290 43912 43970 43966
rect 44630 44540 45310 44592
rect 44630 44506 44684 44540
rect 44718 44506 44774 44540
rect 44808 44506 44864 44540
rect 44898 44506 44954 44540
rect 44988 44506 45044 44540
rect 45078 44506 45134 44540
rect 45168 44506 45224 44540
rect 45258 44506 45310 44540
rect 44630 44450 45310 44506
rect 44630 44416 44684 44450
rect 44718 44416 44774 44450
rect 44808 44416 44864 44450
rect 44898 44416 44954 44450
rect 44988 44416 45044 44450
rect 45078 44416 45134 44450
rect 45168 44416 45224 44450
rect 45258 44416 45310 44450
rect 44630 44360 45310 44416
rect 44630 44326 44684 44360
rect 44718 44326 44774 44360
rect 44808 44326 44864 44360
rect 44898 44326 44954 44360
rect 44988 44326 45044 44360
rect 45078 44326 45134 44360
rect 45168 44326 45224 44360
rect 45258 44326 45310 44360
rect 44630 44270 45310 44326
rect 44630 44236 44684 44270
rect 44718 44236 44774 44270
rect 44808 44236 44864 44270
rect 44898 44236 44954 44270
rect 44988 44236 45044 44270
rect 45078 44236 45134 44270
rect 45168 44236 45224 44270
rect 45258 44236 45310 44270
rect 44630 44180 45310 44236
rect 44630 44146 44684 44180
rect 44718 44146 44774 44180
rect 44808 44146 44864 44180
rect 44898 44146 44954 44180
rect 44988 44146 45044 44180
rect 45078 44146 45134 44180
rect 45168 44146 45224 44180
rect 45258 44146 45310 44180
rect 44630 44090 45310 44146
rect 44630 44056 44684 44090
rect 44718 44056 44774 44090
rect 44808 44056 44864 44090
rect 44898 44056 44954 44090
rect 44988 44056 45044 44090
rect 45078 44056 45134 44090
rect 45168 44056 45224 44090
rect 45258 44056 45310 44090
rect 44630 44000 45310 44056
rect 44630 43966 44684 44000
rect 44718 43966 44774 44000
rect 44808 43966 44864 44000
rect 44898 43966 44954 44000
rect 44988 43966 45044 44000
rect 45078 43966 45134 44000
rect 45168 43966 45224 44000
rect 45258 43966 45310 44000
rect 44630 43912 45310 43966
rect 45970 44540 46650 44592
rect 45970 44506 46024 44540
rect 46058 44506 46114 44540
rect 46148 44506 46204 44540
rect 46238 44506 46294 44540
rect 46328 44506 46384 44540
rect 46418 44506 46474 44540
rect 46508 44506 46564 44540
rect 46598 44506 46650 44540
rect 45970 44450 46650 44506
rect 45970 44416 46024 44450
rect 46058 44416 46114 44450
rect 46148 44416 46204 44450
rect 46238 44416 46294 44450
rect 46328 44416 46384 44450
rect 46418 44416 46474 44450
rect 46508 44416 46564 44450
rect 46598 44416 46650 44450
rect 45970 44360 46650 44416
rect 45970 44326 46024 44360
rect 46058 44326 46114 44360
rect 46148 44326 46204 44360
rect 46238 44326 46294 44360
rect 46328 44326 46384 44360
rect 46418 44326 46474 44360
rect 46508 44326 46564 44360
rect 46598 44326 46650 44360
rect 45970 44270 46650 44326
rect 45970 44236 46024 44270
rect 46058 44236 46114 44270
rect 46148 44236 46204 44270
rect 46238 44236 46294 44270
rect 46328 44236 46384 44270
rect 46418 44236 46474 44270
rect 46508 44236 46564 44270
rect 46598 44236 46650 44270
rect 45970 44180 46650 44236
rect 45970 44146 46024 44180
rect 46058 44146 46114 44180
rect 46148 44146 46204 44180
rect 46238 44146 46294 44180
rect 46328 44146 46384 44180
rect 46418 44146 46474 44180
rect 46508 44146 46564 44180
rect 46598 44146 46650 44180
rect 45970 44090 46650 44146
rect 45970 44056 46024 44090
rect 46058 44056 46114 44090
rect 46148 44056 46204 44090
rect 46238 44056 46294 44090
rect 46328 44056 46384 44090
rect 46418 44056 46474 44090
rect 46508 44056 46564 44090
rect 46598 44056 46650 44090
rect 45970 44000 46650 44056
rect 45970 43966 46024 44000
rect 46058 43966 46114 44000
rect 46148 43966 46204 44000
rect 46238 43966 46294 44000
rect 46328 43966 46384 44000
rect 46418 43966 46474 44000
rect 46508 43966 46564 44000
rect 46598 43966 46650 44000
rect 45970 43912 46650 43966
rect 47310 44540 47990 44592
rect 47310 44506 47364 44540
rect 47398 44506 47454 44540
rect 47488 44506 47544 44540
rect 47578 44506 47634 44540
rect 47668 44506 47724 44540
rect 47758 44506 47814 44540
rect 47848 44506 47904 44540
rect 47938 44506 47990 44540
rect 47310 44450 47990 44506
rect 47310 44416 47364 44450
rect 47398 44416 47454 44450
rect 47488 44416 47544 44450
rect 47578 44416 47634 44450
rect 47668 44416 47724 44450
rect 47758 44416 47814 44450
rect 47848 44416 47904 44450
rect 47938 44416 47990 44450
rect 47310 44360 47990 44416
rect 47310 44326 47364 44360
rect 47398 44326 47454 44360
rect 47488 44326 47544 44360
rect 47578 44326 47634 44360
rect 47668 44326 47724 44360
rect 47758 44326 47814 44360
rect 47848 44326 47904 44360
rect 47938 44326 47990 44360
rect 47310 44270 47990 44326
rect 47310 44236 47364 44270
rect 47398 44236 47454 44270
rect 47488 44236 47544 44270
rect 47578 44236 47634 44270
rect 47668 44236 47724 44270
rect 47758 44236 47814 44270
rect 47848 44236 47904 44270
rect 47938 44236 47990 44270
rect 47310 44180 47990 44236
rect 47310 44146 47364 44180
rect 47398 44146 47454 44180
rect 47488 44146 47544 44180
rect 47578 44146 47634 44180
rect 47668 44146 47724 44180
rect 47758 44146 47814 44180
rect 47848 44146 47904 44180
rect 47938 44146 47990 44180
rect 47310 44090 47990 44146
rect 47310 44056 47364 44090
rect 47398 44056 47454 44090
rect 47488 44056 47544 44090
rect 47578 44056 47634 44090
rect 47668 44056 47724 44090
rect 47758 44056 47814 44090
rect 47848 44056 47904 44090
rect 47938 44056 47990 44090
rect 47310 44000 47990 44056
rect 47310 43966 47364 44000
rect 47398 43966 47454 44000
rect 47488 43966 47544 44000
rect 47578 43966 47634 44000
rect 47668 43966 47724 44000
rect 47758 43966 47814 44000
rect 47848 43966 47904 44000
rect 47938 43966 47990 44000
rect 47310 43912 47990 43966
rect 48650 44540 49330 44592
rect 48650 44506 48704 44540
rect 48738 44506 48794 44540
rect 48828 44506 48884 44540
rect 48918 44506 48974 44540
rect 49008 44506 49064 44540
rect 49098 44506 49154 44540
rect 49188 44506 49244 44540
rect 49278 44506 49330 44540
rect 48650 44450 49330 44506
rect 48650 44416 48704 44450
rect 48738 44416 48794 44450
rect 48828 44416 48884 44450
rect 48918 44416 48974 44450
rect 49008 44416 49064 44450
rect 49098 44416 49154 44450
rect 49188 44416 49244 44450
rect 49278 44416 49330 44450
rect 48650 44360 49330 44416
rect 48650 44326 48704 44360
rect 48738 44326 48794 44360
rect 48828 44326 48884 44360
rect 48918 44326 48974 44360
rect 49008 44326 49064 44360
rect 49098 44326 49154 44360
rect 49188 44326 49244 44360
rect 49278 44326 49330 44360
rect 48650 44270 49330 44326
rect 48650 44236 48704 44270
rect 48738 44236 48794 44270
rect 48828 44236 48884 44270
rect 48918 44236 48974 44270
rect 49008 44236 49064 44270
rect 49098 44236 49154 44270
rect 49188 44236 49244 44270
rect 49278 44236 49330 44270
rect 48650 44180 49330 44236
rect 48650 44146 48704 44180
rect 48738 44146 48794 44180
rect 48828 44146 48884 44180
rect 48918 44146 48974 44180
rect 49008 44146 49064 44180
rect 49098 44146 49154 44180
rect 49188 44146 49244 44180
rect 49278 44146 49330 44180
rect 48650 44090 49330 44146
rect 48650 44056 48704 44090
rect 48738 44056 48794 44090
rect 48828 44056 48884 44090
rect 48918 44056 48974 44090
rect 49008 44056 49064 44090
rect 49098 44056 49154 44090
rect 49188 44056 49244 44090
rect 49278 44056 49330 44090
rect 48650 44000 49330 44056
rect 48650 43966 48704 44000
rect 48738 43966 48794 44000
rect 48828 43966 48884 44000
rect 48918 43966 48974 44000
rect 49008 43966 49064 44000
rect 49098 43966 49154 44000
rect 49188 43966 49244 44000
rect 49278 43966 49330 44000
rect 48650 43912 49330 43966
rect 49990 44540 50670 44592
rect 49990 44506 50044 44540
rect 50078 44506 50134 44540
rect 50168 44506 50224 44540
rect 50258 44506 50314 44540
rect 50348 44506 50404 44540
rect 50438 44506 50494 44540
rect 50528 44506 50584 44540
rect 50618 44506 50670 44540
rect 49990 44450 50670 44506
rect 49990 44416 50044 44450
rect 50078 44416 50134 44450
rect 50168 44416 50224 44450
rect 50258 44416 50314 44450
rect 50348 44416 50404 44450
rect 50438 44416 50494 44450
rect 50528 44416 50584 44450
rect 50618 44416 50670 44450
rect 49990 44360 50670 44416
rect 49990 44326 50044 44360
rect 50078 44326 50134 44360
rect 50168 44326 50224 44360
rect 50258 44326 50314 44360
rect 50348 44326 50404 44360
rect 50438 44326 50494 44360
rect 50528 44326 50584 44360
rect 50618 44326 50670 44360
rect 49990 44270 50670 44326
rect 49990 44236 50044 44270
rect 50078 44236 50134 44270
rect 50168 44236 50224 44270
rect 50258 44236 50314 44270
rect 50348 44236 50404 44270
rect 50438 44236 50494 44270
rect 50528 44236 50584 44270
rect 50618 44236 50670 44270
rect 49990 44180 50670 44236
rect 49990 44146 50044 44180
rect 50078 44146 50134 44180
rect 50168 44146 50224 44180
rect 50258 44146 50314 44180
rect 50348 44146 50404 44180
rect 50438 44146 50494 44180
rect 50528 44146 50584 44180
rect 50618 44146 50670 44180
rect 49990 44090 50670 44146
rect 49990 44056 50044 44090
rect 50078 44056 50134 44090
rect 50168 44056 50224 44090
rect 50258 44056 50314 44090
rect 50348 44056 50404 44090
rect 50438 44056 50494 44090
rect 50528 44056 50584 44090
rect 50618 44056 50670 44090
rect 49990 44000 50670 44056
rect 49990 43966 50044 44000
rect 50078 43966 50134 44000
rect 50168 43966 50224 44000
rect 50258 43966 50314 44000
rect 50348 43966 50404 44000
rect 50438 43966 50494 44000
rect 50528 43966 50584 44000
rect 50618 43966 50670 44000
rect 49990 43912 50670 43966
rect 51330 44540 52010 44592
rect 51330 44506 51384 44540
rect 51418 44506 51474 44540
rect 51508 44506 51564 44540
rect 51598 44506 51654 44540
rect 51688 44506 51744 44540
rect 51778 44506 51834 44540
rect 51868 44506 51924 44540
rect 51958 44506 52010 44540
rect 51330 44450 52010 44506
rect 51330 44416 51384 44450
rect 51418 44416 51474 44450
rect 51508 44416 51564 44450
rect 51598 44416 51654 44450
rect 51688 44416 51744 44450
rect 51778 44416 51834 44450
rect 51868 44416 51924 44450
rect 51958 44416 52010 44450
rect 51330 44360 52010 44416
rect 51330 44326 51384 44360
rect 51418 44326 51474 44360
rect 51508 44326 51564 44360
rect 51598 44326 51654 44360
rect 51688 44326 51744 44360
rect 51778 44326 51834 44360
rect 51868 44326 51924 44360
rect 51958 44326 52010 44360
rect 51330 44270 52010 44326
rect 51330 44236 51384 44270
rect 51418 44236 51474 44270
rect 51508 44236 51564 44270
rect 51598 44236 51654 44270
rect 51688 44236 51744 44270
rect 51778 44236 51834 44270
rect 51868 44236 51924 44270
rect 51958 44236 52010 44270
rect 51330 44180 52010 44236
rect 51330 44146 51384 44180
rect 51418 44146 51474 44180
rect 51508 44146 51564 44180
rect 51598 44146 51654 44180
rect 51688 44146 51744 44180
rect 51778 44146 51834 44180
rect 51868 44146 51924 44180
rect 51958 44146 52010 44180
rect 51330 44090 52010 44146
rect 51330 44056 51384 44090
rect 51418 44056 51474 44090
rect 51508 44056 51564 44090
rect 51598 44056 51654 44090
rect 51688 44056 51744 44090
rect 51778 44056 51834 44090
rect 51868 44056 51924 44090
rect 51958 44056 52010 44090
rect 51330 44000 52010 44056
rect 51330 43966 51384 44000
rect 51418 43966 51474 44000
rect 51508 43966 51564 44000
rect 51598 43966 51654 44000
rect 51688 43966 51744 44000
rect 51778 43966 51834 44000
rect 51868 43966 51924 44000
rect 51958 43966 52010 44000
rect 51330 43912 52010 43966
rect 22709 41181 22767 41197
rect 22709 41147 22721 41181
rect 22755 41147 22767 41181
rect 22709 41113 22767 41147
rect 22709 41079 22721 41113
rect 22755 41079 22767 41113
rect 22709 41045 22767 41079
rect 22709 41011 22721 41045
rect 22755 41011 22767 41045
rect 22709 40977 22767 41011
rect 22709 40943 22721 40977
rect 22755 40943 22767 40977
rect 22709 40909 22767 40943
rect 22709 40875 22721 40909
rect 22755 40875 22767 40909
rect 22709 40841 22767 40875
rect 22709 40807 22721 40841
rect 22755 40807 22767 40841
rect 22709 40773 22767 40807
rect 22709 40739 22721 40773
rect 22755 40739 22767 40773
rect 22709 40705 22767 40739
rect 22709 40671 22721 40705
rect 22755 40671 22767 40705
rect 22709 40637 22767 40671
rect 22709 40603 22721 40637
rect 22755 40603 22767 40637
rect 22709 40569 22767 40603
rect 22709 40535 22721 40569
rect 22755 40535 22767 40569
rect 22709 40501 22767 40535
rect 22709 40467 22721 40501
rect 22755 40467 22767 40501
rect 22709 40433 22767 40467
rect 22709 40399 22721 40433
rect 22755 40399 22767 40433
rect 22709 40365 22767 40399
rect 22709 40331 22721 40365
rect 22755 40331 22767 40365
rect 22709 40297 22767 40331
rect 22709 40263 22721 40297
rect 22755 40263 22767 40297
rect 22709 40229 22767 40263
rect 22709 40195 22721 40229
rect 22755 40195 22767 40229
rect 22709 40161 22767 40195
rect 22709 40127 22721 40161
rect 22755 40127 22767 40161
rect 22709 40093 22767 40127
rect 22709 40059 22721 40093
rect 22755 40059 22767 40093
rect 22709 40025 22767 40059
rect 22709 39991 22721 40025
rect 22755 39991 22767 40025
rect 22709 39957 22767 39991
rect 22709 39923 22721 39957
rect 22755 39923 22767 39957
rect 22709 39907 22767 39923
rect 23167 41181 23225 41197
rect 23167 41147 23179 41181
rect 23213 41147 23225 41181
rect 23167 41113 23225 41147
rect 23167 41079 23179 41113
rect 23213 41079 23225 41113
rect 23167 41045 23225 41079
rect 23167 41011 23179 41045
rect 23213 41011 23225 41045
rect 23167 40977 23225 41011
rect 23167 40943 23179 40977
rect 23213 40943 23225 40977
rect 23167 40909 23225 40943
rect 23167 40875 23179 40909
rect 23213 40875 23225 40909
rect 23167 40841 23225 40875
rect 23167 40807 23179 40841
rect 23213 40807 23225 40841
rect 23167 40773 23225 40807
rect 23167 40739 23179 40773
rect 23213 40739 23225 40773
rect 23167 40705 23225 40739
rect 23167 40671 23179 40705
rect 23213 40671 23225 40705
rect 23167 40637 23225 40671
rect 23167 40603 23179 40637
rect 23213 40603 23225 40637
rect 23167 40569 23225 40603
rect 23167 40535 23179 40569
rect 23213 40535 23225 40569
rect 23167 40501 23225 40535
rect 23167 40467 23179 40501
rect 23213 40467 23225 40501
rect 23167 40433 23225 40467
rect 23167 40399 23179 40433
rect 23213 40399 23225 40433
rect 23167 40365 23225 40399
rect 23167 40331 23179 40365
rect 23213 40331 23225 40365
rect 23167 40297 23225 40331
rect 23167 40263 23179 40297
rect 23213 40263 23225 40297
rect 23167 40229 23225 40263
rect 23167 40195 23179 40229
rect 23213 40195 23225 40229
rect 23167 40161 23225 40195
rect 23167 40127 23179 40161
rect 23213 40127 23225 40161
rect 23167 40093 23225 40127
rect 23167 40059 23179 40093
rect 23213 40059 23225 40093
rect 23167 40025 23225 40059
rect 23167 39991 23179 40025
rect 23213 39991 23225 40025
rect 23167 39957 23225 39991
rect 23167 39923 23179 39957
rect 23213 39923 23225 39957
rect 23167 39907 23225 39923
rect 23625 41181 23683 41197
rect 23625 41147 23637 41181
rect 23671 41147 23683 41181
rect 23625 41113 23683 41147
rect 23625 41079 23637 41113
rect 23671 41079 23683 41113
rect 23625 41045 23683 41079
rect 23625 41011 23637 41045
rect 23671 41011 23683 41045
rect 23625 40977 23683 41011
rect 23625 40943 23637 40977
rect 23671 40943 23683 40977
rect 23625 40909 23683 40943
rect 23625 40875 23637 40909
rect 23671 40875 23683 40909
rect 23625 40841 23683 40875
rect 23625 40807 23637 40841
rect 23671 40807 23683 40841
rect 23625 40773 23683 40807
rect 23625 40739 23637 40773
rect 23671 40739 23683 40773
rect 23625 40705 23683 40739
rect 23625 40671 23637 40705
rect 23671 40671 23683 40705
rect 23625 40637 23683 40671
rect 23625 40603 23637 40637
rect 23671 40603 23683 40637
rect 23625 40569 23683 40603
rect 23625 40535 23637 40569
rect 23671 40535 23683 40569
rect 23625 40501 23683 40535
rect 23625 40467 23637 40501
rect 23671 40467 23683 40501
rect 23625 40433 23683 40467
rect 23625 40399 23637 40433
rect 23671 40399 23683 40433
rect 23625 40365 23683 40399
rect 23625 40331 23637 40365
rect 23671 40331 23683 40365
rect 23625 40297 23683 40331
rect 23625 40263 23637 40297
rect 23671 40263 23683 40297
rect 23625 40229 23683 40263
rect 23625 40195 23637 40229
rect 23671 40195 23683 40229
rect 23625 40161 23683 40195
rect 23625 40127 23637 40161
rect 23671 40127 23683 40161
rect 23625 40093 23683 40127
rect 23625 40059 23637 40093
rect 23671 40059 23683 40093
rect 23625 40025 23683 40059
rect 23625 39991 23637 40025
rect 23671 39991 23683 40025
rect 23625 39957 23683 39991
rect 23625 39923 23637 39957
rect 23671 39923 23683 39957
rect 23625 39907 23683 39923
rect 24083 41181 24141 41197
rect 24083 41147 24095 41181
rect 24129 41147 24141 41181
rect 24083 41113 24141 41147
rect 24083 41079 24095 41113
rect 24129 41079 24141 41113
rect 24083 41045 24141 41079
rect 24083 41011 24095 41045
rect 24129 41011 24141 41045
rect 24083 40977 24141 41011
rect 24083 40943 24095 40977
rect 24129 40943 24141 40977
rect 24083 40909 24141 40943
rect 24083 40875 24095 40909
rect 24129 40875 24141 40909
rect 24083 40841 24141 40875
rect 24083 40807 24095 40841
rect 24129 40807 24141 40841
rect 24083 40773 24141 40807
rect 24083 40739 24095 40773
rect 24129 40739 24141 40773
rect 24083 40705 24141 40739
rect 24083 40671 24095 40705
rect 24129 40671 24141 40705
rect 24083 40637 24141 40671
rect 24083 40603 24095 40637
rect 24129 40603 24141 40637
rect 24083 40569 24141 40603
rect 24083 40535 24095 40569
rect 24129 40535 24141 40569
rect 24083 40501 24141 40535
rect 24083 40467 24095 40501
rect 24129 40467 24141 40501
rect 24083 40433 24141 40467
rect 24083 40399 24095 40433
rect 24129 40399 24141 40433
rect 24083 40365 24141 40399
rect 24083 40331 24095 40365
rect 24129 40331 24141 40365
rect 24083 40297 24141 40331
rect 24083 40263 24095 40297
rect 24129 40263 24141 40297
rect 24083 40229 24141 40263
rect 24083 40195 24095 40229
rect 24129 40195 24141 40229
rect 24083 40161 24141 40195
rect 24083 40127 24095 40161
rect 24129 40127 24141 40161
rect 24083 40093 24141 40127
rect 24083 40059 24095 40093
rect 24129 40059 24141 40093
rect 24083 40025 24141 40059
rect 24083 39991 24095 40025
rect 24129 39991 24141 40025
rect 24083 39957 24141 39991
rect 24083 39923 24095 39957
rect 24129 39923 24141 39957
rect 24083 39907 24141 39923
rect 24541 41181 24599 41197
rect 24541 41147 24553 41181
rect 24587 41147 24599 41181
rect 24541 41113 24599 41147
rect 24541 41079 24553 41113
rect 24587 41079 24599 41113
rect 24541 41045 24599 41079
rect 24541 41011 24553 41045
rect 24587 41011 24599 41045
rect 24541 40977 24599 41011
rect 24541 40943 24553 40977
rect 24587 40943 24599 40977
rect 24541 40909 24599 40943
rect 24541 40875 24553 40909
rect 24587 40875 24599 40909
rect 24541 40841 24599 40875
rect 24541 40807 24553 40841
rect 24587 40807 24599 40841
rect 24541 40773 24599 40807
rect 24541 40739 24553 40773
rect 24587 40739 24599 40773
rect 24541 40705 24599 40739
rect 24541 40671 24553 40705
rect 24587 40671 24599 40705
rect 24541 40637 24599 40671
rect 24541 40603 24553 40637
rect 24587 40603 24599 40637
rect 24541 40569 24599 40603
rect 24541 40535 24553 40569
rect 24587 40535 24599 40569
rect 24541 40501 24599 40535
rect 24541 40467 24553 40501
rect 24587 40467 24599 40501
rect 24541 40433 24599 40467
rect 24541 40399 24553 40433
rect 24587 40399 24599 40433
rect 24541 40365 24599 40399
rect 24541 40331 24553 40365
rect 24587 40331 24599 40365
rect 24541 40297 24599 40331
rect 24541 40263 24553 40297
rect 24587 40263 24599 40297
rect 24541 40229 24599 40263
rect 24541 40195 24553 40229
rect 24587 40195 24599 40229
rect 24541 40161 24599 40195
rect 24541 40127 24553 40161
rect 24587 40127 24599 40161
rect 24541 40093 24599 40127
rect 24541 40059 24553 40093
rect 24587 40059 24599 40093
rect 24541 40025 24599 40059
rect 24541 39991 24553 40025
rect 24587 39991 24599 40025
rect 24541 39957 24599 39991
rect 24541 39923 24553 39957
rect 24587 39923 24599 39957
rect 24541 39907 24599 39923
rect 24999 41181 25057 41197
rect 24999 41147 25011 41181
rect 25045 41147 25057 41181
rect 24999 41113 25057 41147
rect 24999 41079 25011 41113
rect 25045 41079 25057 41113
rect 24999 41045 25057 41079
rect 24999 41011 25011 41045
rect 25045 41011 25057 41045
rect 24999 40977 25057 41011
rect 24999 40943 25011 40977
rect 25045 40943 25057 40977
rect 24999 40909 25057 40943
rect 24999 40875 25011 40909
rect 25045 40875 25057 40909
rect 24999 40841 25057 40875
rect 24999 40807 25011 40841
rect 25045 40807 25057 40841
rect 24999 40773 25057 40807
rect 24999 40739 25011 40773
rect 25045 40739 25057 40773
rect 24999 40705 25057 40739
rect 24999 40671 25011 40705
rect 25045 40671 25057 40705
rect 24999 40637 25057 40671
rect 24999 40603 25011 40637
rect 25045 40603 25057 40637
rect 24999 40569 25057 40603
rect 24999 40535 25011 40569
rect 25045 40535 25057 40569
rect 24999 40501 25057 40535
rect 24999 40467 25011 40501
rect 25045 40467 25057 40501
rect 24999 40433 25057 40467
rect 24999 40399 25011 40433
rect 25045 40399 25057 40433
rect 24999 40365 25057 40399
rect 24999 40331 25011 40365
rect 25045 40331 25057 40365
rect 24999 40297 25057 40331
rect 24999 40263 25011 40297
rect 25045 40263 25057 40297
rect 24999 40229 25057 40263
rect 24999 40195 25011 40229
rect 25045 40195 25057 40229
rect 24999 40161 25057 40195
rect 24999 40127 25011 40161
rect 25045 40127 25057 40161
rect 24999 40093 25057 40127
rect 24999 40059 25011 40093
rect 25045 40059 25057 40093
rect 24999 40025 25057 40059
rect 24999 39991 25011 40025
rect 25045 39991 25057 40025
rect 24999 39957 25057 39991
rect 24999 39923 25011 39957
rect 25045 39923 25057 39957
rect 24999 39907 25057 39923
rect 25457 41181 25515 41197
rect 25457 41147 25469 41181
rect 25503 41147 25515 41181
rect 25457 41113 25515 41147
rect 25457 41079 25469 41113
rect 25503 41079 25515 41113
rect 25457 41045 25515 41079
rect 25457 41011 25469 41045
rect 25503 41011 25515 41045
rect 25457 40977 25515 41011
rect 25457 40943 25469 40977
rect 25503 40943 25515 40977
rect 25457 40909 25515 40943
rect 25457 40875 25469 40909
rect 25503 40875 25515 40909
rect 25457 40841 25515 40875
rect 25457 40807 25469 40841
rect 25503 40807 25515 40841
rect 25457 40773 25515 40807
rect 25457 40739 25469 40773
rect 25503 40739 25515 40773
rect 25457 40705 25515 40739
rect 25457 40671 25469 40705
rect 25503 40671 25515 40705
rect 25457 40637 25515 40671
rect 25457 40603 25469 40637
rect 25503 40603 25515 40637
rect 25457 40569 25515 40603
rect 25457 40535 25469 40569
rect 25503 40535 25515 40569
rect 25457 40501 25515 40535
rect 25457 40467 25469 40501
rect 25503 40467 25515 40501
rect 25457 40433 25515 40467
rect 25457 40399 25469 40433
rect 25503 40399 25515 40433
rect 25457 40365 25515 40399
rect 25457 40331 25469 40365
rect 25503 40331 25515 40365
rect 25457 40297 25515 40331
rect 25457 40263 25469 40297
rect 25503 40263 25515 40297
rect 25457 40229 25515 40263
rect 25457 40195 25469 40229
rect 25503 40195 25515 40229
rect 25457 40161 25515 40195
rect 25457 40127 25469 40161
rect 25503 40127 25515 40161
rect 25457 40093 25515 40127
rect 25457 40059 25469 40093
rect 25503 40059 25515 40093
rect 25457 40025 25515 40059
rect 25457 39991 25469 40025
rect 25503 39991 25515 40025
rect 25457 39957 25515 39991
rect 25457 39923 25469 39957
rect 25503 39923 25515 39957
rect 25457 39907 25515 39923
rect 25915 41181 25973 41197
rect 25915 41147 25927 41181
rect 25961 41147 25973 41181
rect 25915 41113 25973 41147
rect 25915 41079 25927 41113
rect 25961 41079 25973 41113
rect 25915 41045 25973 41079
rect 25915 41011 25927 41045
rect 25961 41011 25973 41045
rect 25915 40977 25973 41011
rect 25915 40943 25927 40977
rect 25961 40943 25973 40977
rect 25915 40909 25973 40943
rect 25915 40875 25927 40909
rect 25961 40875 25973 40909
rect 25915 40841 25973 40875
rect 25915 40807 25927 40841
rect 25961 40807 25973 40841
rect 25915 40773 25973 40807
rect 25915 40739 25927 40773
rect 25961 40739 25973 40773
rect 25915 40705 25973 40739
rect 25915 40671 25927 40705
rect 25961 40671 25973 40705
rect 25915 40637 25973 40671
rect 25915 40603 25927 40637
rect 25961 40603 25973 40637
rect 25915 40569 25973 40603
rect 25915 40535 25927 40569
rect 25961 40535 25973 40569
rect 25915 40501 25973 40535
rect 25915 40467 25927 40501
rect 25961 40467 25973 40501
rect 25915 40433 25973 40467
rect 25915 40399 25927 40433
rect 25961 40399 25973 40433
rect 25915 40365 25973 40399
rect 25915 40331 25927 40365
rect 25961 40331 25973 40365
rect 25915 40297 25973 40331
rect 25915 40263 25927 40297
rect 25961 40263 25973 40297
rect 25915 40229 25973 40263
rect 25915 40195 25927 40229
rect 25961 40195 25973 40229
rect 25915 40161 25973 40195
rect 25915 40127 25927 40161
rect 25961 40127 25973 40161
rect 25915 40093 25973 40127
rect 25915 40059 25927 40093
rect 25961 40059 25973 40093
rect 25915 40025 25973 40059
rect 25915 39991 25927 40025
rect 25961 39991 25973 40025
rect 25915 39957 25973 39991
rect 25915 39923 25927 39957
rect 25961 39923 25973 39957
rect 25915 39907 25973 39923
rect 26373 41181 26431 41197
rect 26373 41147 26385 41181
rect 26419 41147 26431 41181
rect 26373 41113 26431 41147
rect 26373 41079 26385 41113
rect 26419 41079 26431 41113
rect 26373 41045 26431 41079
rect 26373 41011 26385 41045
rect 26419 41011 26431 41045
rect 26373 40977 26431 41011
rect 26373 40943 26385 40977
rect 26419 40943 26431 40977
rect 26373 40909 26431 40943
rect 26373 40875 26385 40909
rect 26419 40875 26431 40909
rect 26373 40841 26431 40875
rect 26373 40807 26385 40841
rect 26419 40807 26431 40841
rect 26373 40773 26431 40807
rect 26373 40739 26385 40773
rect 26419 40739 26431 40773
rect 26373 40705 26431 40739
rect 26373 40671 26385 40705
rect 26419 40671 26431 40705
rect 26373 40637 26431 40671
rect 26373 40603 26385 40637
rect 26419 40603 26431 40637
rect 26373 40569 26431 40603
rect 26373 40535 26385 40569
rect 26419 40535 26431 40569
rect 26373 40501 26431 40535
rect 26373 40467 26385 40501
rect 26419 40467 26431 40501
rect 26373 40433 26431 40467
rect 26373 40399 26385 40433
rect 26419 40399 26431 40433
rect 26373 40365 26431 40399
rect 26373 40331 26385 40365
rect 26419 40331 26431 40365
rect 26373 40297 26431 40331
rect 26373 40263 26385 40297
rect 26419 40263 26431 40297
rect 26373 40229 26431 40263
rect 26373 40195 26385 40229
rect 26419 40195 26431 40229
rect 26373 40161 26431 40195
rect 26373 40127 26385 40161
rect 26419 40127 26431 40161
rect 26373 40093 26431 40127
rect 26373 40059 26385 40093
rect 26419 40059 26431 40093
rect 26373 40025 26431 40059
rect 26373 39991 26385 40025
rect 26419 39991 26431 40025
rect 26373 39957 26431 39991
rect 26373 39923 26385 39957
rect 26419 39923 26431 39957
rect 26373 39907 26431 39923
rect 26831 41181 26889 41197
rect 26831 41147 26843 41181
rect 26877 41147 26889 41181
rect 26831 41113 26889 41147
rect 26831 41079 26843 41113
rect 26877 41079 26889 41113
rect 26831 41045 26889 41079
rect 26831 41011 26843 41045
rect 26877 41011 26889 41045
rect 26831 40977 26889 41011
rect 26831 40943 26843 40977
rect 26877 40943 26889 40977
rect 26831 40909 26889 40943
rect 26831 40875 26843 40909
rect 26877 40875 26889 40909
rect 26831 40841 26889 40875
rect 26831 40807 26843 40841
rect 26877 40807 26889 40841
rect 26831 40773 26889 40807
rect 26831 40739 26843 40773
rect 26877 40739 26889 40773
rect 26831 40705 26889 40739
rect 26831 40671 26843 40705
rect 26877 40671 26889 40705
rect 26831 40637 26889 40671
rect 26831 40603 26843 40637
rect 26877 40603 26889 40637
rect 26831 40569 26889 40603
rect 26831 40535 26843 40569
rect 26877 40535 26889 40569
rect 26831 40501 26889 40535
rect 26831 40467 26843 40501
rect 26877 40467 26889 40501
rect 26831 40433 26889 40467
rect 26831 40399 26843 40433
rect 26877 40399 26889 40433
rect 26831 40365 26889 40399
rect 26831 40331 26843 40365
rect 26877 40331 26889 40365
rect 26831 40297 26889 40331
rect 26831 40263 26843 40297
rect 26877 40263 26889 40297
rect 26831 40229 26889 40263
rect 26831 40195 26843 40229
rect 26877 40195 26889 40229
rect 26831 40161 26889 40195
rect 26831 40127 26843 40161
rect 26877 40127 26889 40161
rect 26831 40093 26889 40127
rect 26831 40059 26843 40093
rect 26877 40059 26889 40093
rect 26831 40025 26889 40059
rect 26831 39991 26843 40025
rect 26877 39991 26889 40025
rect 26831 39957 26889 39991
rect 26831 39923 26843 39957
rect 26877 39923 26889 39957
rect 26831 39907 26889 39923
rect 27289 41181 27347 41197
rect 27289 41147 27301 41181
rect 27335 41147 27347 41181
rect 27289 41113 27347 41147
rect 27289 41079 27301 41113
rect 27335 41079 27347 41113
rect 27289 41045 27347 41079
rect 27289 41011 27301 41045
rect 27335 41011 27347 41045
rect 27289 40977 27347 41011
rect 27289 40943 27301 40977
rect 27335 40943 27347 40977
rect 27289 40909 27347 40943
rect 27289 40875 27301 40909
rect 27335 40875 27347 40909
rect 27289 40841 27347 40875
rect 27289 40807 27301 40841
rect 27335 40807 27347 40841
rect 27289 40773 27347 40807
rect 27289 40739 27301 40773
rect 27335 40739 27347 40773
rect 27289 40705 27347 40739
rect 27289 40671 27301 40705
rect 27335 40671 27347 40705
rect 27289 40637 27347 40671
rect 27289 40603 27301 40637
rect 27335 40603 27347 40637
rect 27289 40569 27347 40603
rect 27289 40535 27301 40569
rect 27335 40535 27347 40569
rect 27289 40501 27347 40535
rect 27289 40467 27301 40501
rect 27335 40467 27347 40501
rect 27289 40433 27347 40467
rect 27289 40399 27301 40433
rect 27335 40399 27347 40433
rect 27289 40365 27347 40399
rect 27289 40331 27301 40365
rect 27335 40331 27347 40365
rect 27289 40297 27347 40331
rect 27289 40263 27301 40297
rect 27335 40263 27347 40297
rect 27289 40229 27347 40263
rect 27289 40195 27301 40229
rect 27335 40195 27347 40229
rect 27289 40161 27347 40195
rect 27289 40127 27301 40161
rect 27335 40127 27347 40161
rect 27289 40093 27347 40127
rect 27289 40059 27301 40093
rect 27335 40059 27347 40093
rect 27289 40025 27347 40059
rect 27289 39991 27301 40025
rect 27335 39991 27347 40025
rect 27289 39957 27347 39991
rect 27289 39923 27301 39957
rect 27335 39923 27347 39957
rect 27289 39907 27347 39923
rect 27747 41181 27805 41197
rect 27747 41147 27759 41181
rect 27793 41147 27805 41181
rect 27747 41113 27805 41147
rect 27747 41079 27759 41113
rect 27793 41079 27805 41113
rect 27747 41045 27805 41079
rect 27747 41011 27759 41045
rect 27793 41011 27805 41045
rect 27747 40977 27805 41011
rect 27747 40943 27759 40977
rect 27793 40943 27805 40977
rect 27747 40909 27805 40943
rect 27747 40875 27759 40909
rect 27793 40875 27805 40909
rect 27747 40841 27805 40875
rect 27747 40807 27759 40841
rect 27793 40807 27805 40841
rect 27747 40773 27805 40807
rect 27747 40739 27759 40773
rect 27793 40739 27805 40773
rect 27747 40705 27805 40739
rect 27747 40671 27759 40705
rect 27793 40671 27805 40705
rect 27747 40637 27805 40671
rect 27747 40603 27759 40637
rect 27793 40603 27805 40637
rect 27747 40569 27805 40603
rect 27747 40535 27759 40569
rect 27793 40535 27805 40569
rect 27747 40501 27805 40535
rect 27747 40467 27759 40501
rect 27793 40467 27805 40501
rect 27747 40433 27805 40467
rect 27747 40399 27759 40433
rect 27793 40399 27805 40433
rect 27747 40365 27805 40399
rect 27747 40331 27759 40365
rect 27793 40331 27805 40365
rect 27747 40297 27805 40331
rect 27747 40263 27759 40297
rect 27793 40263 27805 40297
rect 27747 40229 27805 40263
rect 27747 40195 27759 40229
rect 27793 40195 27805 40229
rect 27747 40161 27805 40195
rect 27747 40127 27759 40161
rect 27793 40127 27805 40161
rect 27747 40093 27805 40127
rect 27747 40059 27759 40093
rect 27793 40059 27805 40093
rect 27747 40025 27805 40059
rect 27747 39991 27759 40025
rect 27793 39991 27805 40025
rect 27747 39957 27805 39991
rect 27747 39923 27759 39957
rect 27793 39923 27805 39957
rect 27747 39907 27805 39923
rect 28205 41181 28263 41197
rect 28205 41147 28217 41181
rect 28251 41147 28263 41181
rect 28205 41113 28263 41147
rect 28205 41079 28217 41113
rect 28251 41079 28263 41113
rect 28205 41045 28263 41079
rect 28205 41011 28217 41045
rect 28251 41011 28263 41045
rect 28205 40977 28263 41011
rect 28205 40943 28217 40977
rect 28251 40943 28263 40977
rect 28205 40909 28263 40943
rect 28205 40875 28217 40909
rect 28251 40875 28263 40909
rect 28205 40841 28263 40875
rect 28205 40807 28217 40841
rect 28251 40807 28263 40841
rect 28205 40773 28263 40807
rect 28205 40739 28217 40773
rect 28251 40739 28263 40773
rect 28205 40705 28263 40739
rect 28205 40671 28217 40705
rect 28251 40671 28263 40705
rect 28205 40637 28263 40671
rect 28205 40603 28217 40637
rect 28251 40603 28263 40637
rect 28205 40569 28263 40603
rect 28205 40535 28217 40569
rect 28251 40535 28263 40569
rect 28205 40501 28263 40535
rect 28205 40467 28217 40501
rect 28251 40467 28263 40501
rect 28205 40433 28263 40467
rect 28205 40399 28217 40433
rect 28251 40399 28263 40433
rect 28205 40365 28263 40399
rect 28205 40331 28217 40365
rect 28251 40331 28263 40365
rect 28205 40297 28263 40331
rect 28205 40263 28217 40297
rect 28251 40263 28263 40297
rect 28205 40229 28263 40263
rect 28205 40195 28217 40229
rect 28251 40195 28263 40229
rect 28205 40161 28263 40195
rect 28205 40127 28217 40161
rect 28251 40127 28263 40161
rect 28205 40093 28263 40127
rect 28205 40059 28217 40093
rect 28251 40059 28263 40093
rect 28205 40025 28263 40059
rect 28205 39991 28217 40025
rect 28251 39991 28263 40025
rect 28205 39957 28263 39991
rect 28205 39923 28217 39957
rect 28251 39923 28263 39957
rect 28205 39907 28263 39923
rect 29373 41181 29431 41197
rect 29373 41147 29385 41181
rect 29419 41147 29431 41181
rect 29373 41113 29431 41147
rect 29373 41079 29385 41113
rect 29419 41079 29431 41113
rect 29373 41045 29431 41079
rect 29373 41011 29385 41045
rect 29419 41011 29431 41045
rect 29373 40977 29431 41011
rect 29373 40943 29385 40977
rect 29419 40943 29431 40977
rect 29373 40909 29431 40943
rect 29373 40875 29385 40909
rect 29419 40875 29431 40909
rect 29373 40841 29431 40875
rect 29373 40807 29385 40841
rect 29419 40807 29431 40841
rect 29373 40773 29431 40807
rect 29373 40739 29385 40773
rect 29419 40739 29431 40773
rect 29373 40705 29431 40739
rect 29373 40671 29385 40705
rect 29419 40671 29431 40705
rect 29373 40637 29431 40671
rect 29373 40603 29385 40637
rect 29419 40603 29431 40637
rect 29373 40569 29431 40603
rect 29373 40535 29385 40569
rect 29419 40535 29431 40569
rect 29373 40501 29431 40535
rect 29373 40467 29385 40501
rect 29419 40467 29431 40501
rect 29373 40433 29431 40467
rect 29373 40399 29385 40433
rect 29419 40399 29431 40433
rect 29373 40365 29431 40399
rect 29373 40331 29385 40365
rect 29419 40331 29431 40365
rect 29373 40297 29431 40331
rect 29373 40263 29385 40297
rect 29419 40263 29431 40297
rect 29373 40229 29431 40263
rect 29373 40195 29385 40229
rect 29419 40195 29431 40229
rect 29373 40161 29431 40195
rect 29373 40127 29385 40161
rect 29419 40127 29431 40161
rect 29373 40093 29431 40127
rect 29373 40059 29385 40093
rect 29419 40059 29431 40093
rect 29373 40025 29431 40059
rect 29373 39991 29385 40025
rect 29419 39991 29431 40025
rect 29373 39957 29431 39991
rect 29373 39923 29385 39957
rect 29419 39923 29431 39957
rect 29373 39907 29431 39923
rect 29831 41181 29889 41197
rect 29831 41147 29843 41181
rect 29877 41147 29889 41181
rect 29831 41113 29889 41147
rect 29831 41079 29843 41113
rect 29877 41079 29889 41113
rect 29831 41045 29889 41079
rect 29831 41011 29843 41045
rect 29877 41011 29889 41045
rect 29831 40977 29889 41011
rect 29831 40943 29843 40977
rect 29877 40943 29889 40977
rect 29831 40909 29889 40943
rect 29831 40875 29843 40909
rect 29877 40875 29889 40909
rect 29831 40841 29889 40875
rect 29831 40807 29843 40841
rect 29877 40807 29889 40841
rect 29831 40773 29889 40807
rect 29831 40739 29843 40773
rect 29877 40739 29889 40773
rect 29831 40705 29889 40739
rect 29831 40671 29843 40705
rect 29877 40671 29889 40705
rect 29831 40637 29889 40671
rect 29831 40603 29843 40637
rect 29877 40603 29889 40637
rect 29831 40569 29889 40603
rect 29831 40535 29843 40569
rect 29877 40535 29889 40569
rect 29831 40501 29889 40535
rect 29831 40467 29843 40501
rect 29877 40467 29889 40501
rect 29831 40433 29889 40467
rect 29831 40399 29843 40433
rect 29877 40399 29889 40433
rect 29831 40365 29889 40399
rect 29831 40331 29843 40365
rect 29877 40331 29889 40365
rect 29831 40297 29889 40331
rect 29831 40263 29843 40297
rect 29877 40263 29889 40297
rect 29831 40229 29889 40263
rect 29831 40195 29843 40229
rect 29877 40195 29889 40229
rect 29831 40161 29889 40195
rect 29831 40127 29843 40161
rect 29877 40127 29889 40161
rect 29831 40093 29889 40127
rect 29831 40059 29843 40093
rect 29877 40059 29889 40093
rect 29831 40025 29889 40059
rect 29831 39991 29843 40025
rect 29877 39991 29889 40025
rect 29831 39957 29889 39991
rect 29831 39923 29843 39957
rect 29877 39923 29889 39957
rect 29831 39907 29889 39923
rect 30289 41181 30347 41197
rect 30289 41147 30301 41181
rect 30335 41147 30347 41181
rect 30289 41113 30347 41147
rect 30289 41079 30301 41113
rect 30335 41079 30347 41113
rect 30289 41045 30347 41079
rect 30289 41011 30301 41045
rect 30335 41011 30347 41045
rect 30289 40977 30347 41011
rect 30289 40943 30301 40977
rect 30335 40943 30347 40977
rect 30289 40909 30347 40943
rect 30289 40875 30301 40909
rect 30335 40875 30347 40909
rect 30289 40841 30347 40875
rect 30289 40807 30301 40841
rect 30335 40807 30347 40841
rect 30289 40773 30347 40807
rect 30289 40739 30301 40773
rect 30335 40739 30347 40773
rect 30289 40705 30347 40739
rect 30289 40671 30301 40705
rect 30335 40671 30347 40705
rect 30289 40637 30347 40671
rect 30289 40603 30301 40637
rect 30335 40603 30347 40637
rect 30289 40569 30347 40603
rect 30289 40535 30301 40569
rect 30335 40535 30347 40569
rect 30289 40501 30347 40535
rect 30289 40467 30301 40501
rect 30335 40467 30347 40501
rect 30289 40433 30347 40467
rect 30289 40399 30301 40433
rect 30335 40399 30347 40433
rect 30289 40365 30347 40399
rect 30289 40331 30301 40365
rect 30335 40331 30347 40365
rect 30289 40297 30347 40331
rect 30289 40263 30301 40297
rect 30335 40263 30347 40297
rect 30289 40229 30347 40263
rect 30289 40195 30301 40229
rect 30335 40195 30347 40229
rect 30289 40161 30347 40195
rect 30289 40127 30301 40161
rect 30335 40127 30347 40161
rect 30289 40093 30347 40127
rect 30289 40059 30301 40093
rect 30335 40059 30347 40093
rect 30289 40025 30347 40059
rect 30289 39991 30301 40025
rect 30335 39991 30347 40025
rect 30289 39957 30347 39991
rect 30289 39923 30301 39957
rect 30335 39923 30347 39957
rect 30289 39907 30347 39923
rect 30747 41181 30805 41197
rect 30747 41147 30759 41181
rect 30793 41147 30805 41181
rect 30747 41113 30805 41147
rect 30747 41079 30759 41113
rect 30793 41079 30805 41113
rect 30747 41045 30805 41079
rect 30747 41011 30759 41045
rect 30793 41011 30805 41045
rect 30747 40977 30805 41011
rect 30747 40943 30759 40977
rect 30793 40943 30805 40977
rect 30747 40909 30805 40943
rect 30747 40875 30759 40909
rect 30793 40875 30805 40909
rect 30747 40841 30805 40875
rect 30747 40807 30759 40841
rect 30793 40807 30805 40841
rect 30747 40773 30805 40807
rect 30747 40739 30759 40773
rect 30793 40739 30805 40773
rect 30747 40705 30805 40739
rect 30747 40671 30759 40705
rect 30793 40671 30805 40705
rect 30747 40637 30805 40671
rect 30747 40603 30759 40637
rect 30793 40603 30805 40637
rect 30747 40569 30805 40603
rect 30747 40535 30759 40569
rect 30793 40535 30805 40569
rect 30747 40501 30805 40535
rect 30747 40467 30759 40501
rect 30793 40467 30805 40501
rect 30747 40433 30805 40467
rect 30747 40399 30759 40433
rect 30793 40399 30805 40433
rect 30747 40365 30805 40399
rect 30747 40331 30759 40365
rect 30793 40331 30805 40365
rect 30747 40297 30805 40331
rect 30747 40263 30759 40297
rect 30793 40263 30805 40297
rect 30747 40229 30805 40263
rect 30747 40195 30759 40229
rect 30793 40195 30805 40229
rect 30747 40161 30805 40195
rect 30747 40127 30759 40161
rect 30793 40127 30805 40161
rect 30747 40093 30805 40127
rect 30747 40059 30759 40093
rect 30793 40059 30805 40093
rect 30747 40025 30805 40059
rect 30747 39991 30759 40025
rect 30793 39991 30805 40025
rect 30747 39957 30805 39991
rect 30747 39923 30759 39957
rect 30793 39923 30805 39957
rect 30747 39907 30805 39923
rect 31205 41181 31263 41197
rect 31205 41147 31217 41181
rect 31251 41147 31263 41181
rect 31205 41113 31263 41147
rect 31205 41079 31217 41113
rect 31251 41079 31263 41113
rect 31205 41045 31263 41079
rect 31205 41011 31217 41045
rect 31251 41011 31263 41045
rect 31205 40977 31263 41011
rect 31205 40943 31217 40977
rect 31251 40943 31263 40977
rect 31205 40909 31263 40943
rect 31205 40875 31217 40909
rect 31251 40875 31263 40909
rect 31205 40841 31263 40875
rect 31205 40807 31217 40841
rect 31251 40807 31263 40841
rect 31205 40773 31263 40807
rect 31205 40739 31217 40773
rect 31251 40739 31263 40773
rect 31205 40705 31263 40739
rect 31205 40671 31217 40705
rect 31251 40671 31263 40705
rect 31205 40637 31263 40671
rect 31205 40603 31217 40637
rect 31251 40603 31263 40637
rect 31205 40569 31263 40603
rect 31205 40535 31217 40569
rect 31251 40535 31263 40569
rect 31205 40501 31263 40535
rect 31205 40467 31217 40501
rect 31251 40467 31263 40501
rect 31205 40433 31263 40467
rect 31205 40399 31217 40433
rect 31251 40399 31263 40433
rect 31205 40365 31263 40399
rect 31205 40331 31217 40365
rect 31251 40331 31263 40365
rect 31205 40297 31263 40331
rect 31205 40263 31217 40297
rect 31251 40263 31263 40297
rect 31205 40229 31263 40263
rect 31205 40195 31217 40229
rect 31251 40195 31263 40229
rect 31205 40161 31263 40195
rect 31205 40127 31217 40161
rect 31251 40127 31263 40161
rect 31205 40093 31263 40127
rect 31205 40059 31217 40093
rect 31251 40059 31263 40093
rect 31205 40025 31263 40059
rect 31205 39991 31217 40025
rect 31251 39991 31263 40025
rect 31205 39957 31263 39991
rect 31205 39923 31217 39957
rect 31251 39923 31263 39957
rect 31205 39907 31263 39923
rect 31663 41181 31721 41197
rect 31663 41147 31675 41181
rect 31709 41147 31721 41181
rect 31663 41113 31721 41147
rect 31663 41079 31675 41113
rect 31709 41079 31721 41113
rect 31663 41045 31721 41079
rect 31663 41011 31675 41045
rect 31709 41011 31721 41045
rect 31663 40977 31721 41011
rect 31663 40943 31675 40977
rect 31709 40943 31721 40977
rect 31663 40909 31721 40943
rect 31663 40875 31675 40909
rect 31709 40875 31721 40909
rect 31663 40841 31721 40875
rect 31663 40807 31675 40841
rect 31709 40807 31721 40841
rect 31663 40773 31721 40807
rect 31663 40739 31675 40773
rect 31709 40739 31721 40773
rect 31663 40705 31721 40739
rect 31663 40671 31675 40705
rect 31709 40671 31721 40705
rect 31663 40637 31721 40671
rect 31663 40603 31675 40637
rect 31709 40603 31721 40637
rect 31663 40569 31721 40603
rect 31663 40535 31675 40569
rect 31709 40535 31721 40569
rect 31663 40501 31721 40535
rect 31663 40467 31675 40501
rect 31709 40467 31721 40501
rect 31663 40433 31721 40467
rect 31663 40399 31675 40433
rect 31709 40399 31721 40433
rect 31663 40365 31721 40399
rect 31663 40331 31675 40365
rect 31709 40331 31721 40365
rect 31663 40297 31721 40331
rect 31663 40263 31675 40297
rect 31709 40263 31721 40297
rect 31663 40229 31721 40263
rect 31663 40195 31675 40229
rect 31709 40195 31721 40229
rect 31663 40161 31721 40195
rect 31663 40127 31675 40161
rect 31709 40127 31721 40161
rect 31663 40093 31721 40127
rect 31663 40059 31675 40093
rect 31709 40059 31721 40093
rect 31663 40025 31721 40059
rect 31663 39991 31675 40025
rect 31709 39991 31721 40025
rect 31663 39957 31721 39991
rect 31663 39923 31675 39957
rect 31709 39923 31721 39957
rect 31663 39907 31721 39923
rect 32121 41181 32179 41197
rect 32121 41147 32133 41181
rect 32167 41147 32179 41181
rect 32121 41113 32179 41147
rect 32121 41079 32133 41113
rect 32167 41079 32179 41113
rect 32121 41045 32179 41079
rect 32121 41011 32133 41045
rect 32167 41011 32179 41045
rect 32121 40977 32179 41011
rect 32121 40943 32133 40977
rect 32167 40943 32179 40977
rect 32121 40909 32179 40943
rect 32121 40875 32133 40909
rect 32167 40875 32179 40909
rect 32121 40841 32179 40875
rect 32121 40807 32133 40841
rect 32167 40807 32179 40841
rect 32121 40773 32179 40807
rect 32121 40739 32133 40773
rect 32167 40739 32179 40773
rect 32121 40705 32179 40739
rect 32121 40671 32133 40705
rect 32167 40671 32179 40705
rect 32121 40637 32179 40671
rect 32121 40603 32133 40637
rect 32167 40603 32179 40637
rect 32121 40569 32179 40603
rect 32121 40535 32133 40569
rect 32167 40535 32179 40569
rect 32121 40501 32179 40535
rect 32121 40467 32133 40501
rect 32167 40467 32179 40501
rect 32121 40433 32179 40467
rect 32121 40399 32133 40433
rect 32167 40399 32179 40433
rect 32121 40365 32179 40399
rect 32121 40331 32133 40365
rect 32167 40331 32179 40365
rect 32121 40297 32179 40331
rect 32121 40263 32133 40297
rect 32167 40263 32179 40297
rect 32121 40229 32179 40263
rect 32121 40195 32133 40229
rect 32167 40195 32179 40229
rect 32121 40161 32179 40195
rect 32121 40127 32133 40161
rect 32167 40127 32179 40161
rect 32121 40093 32179 40127
rect 32121 40059 32133 40093
rect 32167 40059 32179 40093
rect 32121 40025 32179 40059
rect 32121 39991 32133 40025
rect 32167 39991 32179 40025
rect 32121 39957 32179 39991
rect 32121 39923 32133 39957
rect 32167 39923 32179 39957
rect 32121 39907 32179 39923
rect 32579 41181 32637 41197
rect 32579 41147 32591 41181
rect 32625 41147 32637 41181
rect 32579 41113 32637 41147
rect 32579 41079 32591 41113
rect 32625 41079 32637 41113
rect 32579 41045 32637 41079
rect 32579 41011 32591 41045
rect 32625 41011 32637 41045
rect 32579 40977 32637 41011
rect 32579 40943 32591 40977
rect 32625 40943 32637 40977
rect 32579 40909 32637 40943
rect 32579 40875 32591 40909
rect 32625 40875 32637 40909
rect 32579 40841 32637 40875
rect 32579 40807 32591 40841
rect 32625 40807 32637 40841
rect 32579 40773 32637 40807
rect 32579 40739 32591 40773
rect 32625 40739 32637 40773
rect 32579 40705 32637 40739
rect 32579 40671 32591 40705
rect 32625 40671 32637 40705
rect 32579 40637 32637 40671
rect 32579 40603 32591 40637
rect 32625 40603 32637 40637
rect 32579 40569 32637 40603
rect 32579 40535 32591 40569
rect 32625 40535 32637 40569
rect 32579 40501 32637 40535
rect 32579 40467 32591 40501
rect 32625 40467 32637 40501
rect 32579 40433 32637 40467
rect 32579 40399 32591 40433
rect 32625 40399 32637 40433
rect 32579 40365 32637 40399
rect 32579 40331 32591 40365
rect 32625 40331 32637 40365
rect 32579 40297 32637 40331
rect 32579 40263 32591 40297
rect 32625 40263 32637 40297
rect 32579 40229 32637 40263
rect 32579 40195 32591 40229
rect 32625 40195 32637 40229
rect 32579 40161 32637 40195
rect 32579 40127 32591 40161
rect 32625 40127 32637 40161
rect 32579 40093 32637 40127
rect 32579 40059 32591 40093
rect 32625 40059 32637 40093
rect 32579 40025 32637 40059
rect 32579 39991 32591 40025
rect 32625 39991 32637 40025
rect 32579 39957 32637 39991
rect 32579 39923 32591 39957
rect 32625 39923 32637 39957
rect 32579 39907 32637 39923
rect 33037 41181 33095 41197
rect 33037 41147 33049 41181
rect 33083 41147 33095 41181
rect 33037 41113 33095 41147
rect 33037 41079 33049 41113
rect 33083 41079 33095 41113
rect 33037 41045 33095 41079
rect 33037 41011 33049 41045
rect 33083 41011 33095 41045
rect 33037 40977 33095 41011
rect 33037 40943 33049 40977
rect 33083 40943 33095 40977
rect 33037 40909 33095 40943
rect 33037 40875 33049 40909
rect 33083 40875 33095 40909
rect 33037 40841 33095 40875
rect 33037 40807 33049 40841
rect 33083 40807 33095 40841
rect 33037 40773 33095 40807
rect 33037 40739 33049 40773
rect 33083 40739 33095 40773
rect 33037 40705 33095 40739
rect 33037 40671 33049 40705
rect 33083 40671 33095 40705
rect 33037 40637 33095 40671
rect 33037 40603 33049 40637
rect 33083 40603 33095 40637
rect 33037 40569 33095 40603
rect 33037 40535 33049 40569
rect 33083 40535 33095 40569
rect 33037 40501 33095 40535
rect 33037 40467 33049 40501
rect 33083 40467 33095 40501
rect 33037 40433 33095 40467
rect 33037 40399 33049 40433
rect 33083 40399 33095 40433
rect 33037 40365 33095 40399
rect 33037 40331 33049 40365
rect 33083 40331 33095 40365
rect 33037 40297 33095 40331
rect 33037 40263 33049 40297
rect 33083 40263 33095 40297
rect 33037 40229 33095 40263
rect 33037 40195 33049 40229
rect 33083 40195 33095 40229
rect 33037 40161 33095 40195
rect 33037 40127 33049 40161
rect 33083 40127 33095 40161
rect 33037 40093 33095 40127
rect 33037 40059 33049 40093
rect 33083 40059 33095 40093
rect 33037 40025 33095 40059
rect 33037 39991 33049 40025
rect 33083 39991 33095 40025
rect 33037 39957 33095 39991
rect 33037 39923 33049 39957
rect 33083 39923 33095 39957
rect 33037 39907 33095 39923
rect 33495 41181 33553 41197
rect 33495 41147 33507 41181
rect 33541 41147 33553 41181
rect 33495 41113 33553 41147
rect 33495 41079 33507 41113
rect 33541 41079 33553 41113
rect 33495 41045 33553 41079
rect 33495 41011 33507 41045
rect 33541 41011 33553 41045
rect 33495 40977 33553 41011
rect 33495 40943 33507 40977
rect 33541 40943 33553 40977
rect 33495 40909 33553 40943
rect 33495 40875 33507 40909
rect 33541 40875 33553 40909
rect 33495 40841 33553 40875
rect 33495 40807 33507 40841
rect 33541 40807 33553 40841
rect 33495 40773 33553 40807
rect 33495 40739 33507 40773
rect 33541 40739 33553 40773
rect 33495 40705 33553 40739
rect 33495 40671 33507 40705
rect 33541 40671 33553 40705
rect 33495 40637 33553 40671
rect 33495 40603 33507 40637
rect 33541 40603 33553 40637
rect 33495 40569 33553 40603
rect 33495 40535 33507 40569
rect 33541 40535 33553 40569
rect 33495 40501 33553 40535
rect 33495 40467 33507 40501
rect 33541 40467 33553 40501
rect 33495 40433 33553 40467
rect 33495 40399 33507 40433
rect 33541 40399 33553 40433
rect 33495 40365 33553 40399
rect 33495 40331 33507 40365
rect 33541 40331 33553 40365
rect 33495 40297 33553 40331
rect 33495 40263 33507 40297
rect 33541 40263 33553 40297
rect 33495 40229 33553 40263
rect 33495 40195 33507 40229
rect 33541 40195 33553 40229
rect 33495 40161 33553 40195
rect 33495 40127 33507 40161
rect 33541 40127 33553 40161
rect 33495 40093 33553 40127
rect 33495 40059 33507 40093
rect 33541 40059 33553 40093
rect 33495 40025 33553 40059
rect 33495 39991 33507 40025
rect 33541 39991 33553 40025
rect 33495 39957 33553 39991
rect 33495 39923 33507 39957
rect 33541 39923 33553 39957
rect 33495 39907 33553 39923
rect 33953 41181 34011 41197
rect 33953 41147 33965 41181
rect 33999 41147 34011 41181
rect 33953 41113 34011 41147
rect 33953 41079 33965 41113
rect 33999 41079 34011 41113
rect 33953 41045 34011 41079
rect 33953 41011 33965 41045
rect 33999 41011 34011 41045
rect 33953 40977 34011 41011
rect 33953 40943 33965 40977
rect 33999 40943 34011 40977
rect 33953 40909 34011 40943
rect 33953 40875 33965 40909
rect 33999 40875 34011 40909
rect 33953 40841 34011 40875
rect 33953 40807 33965 40841
rect 33999 40807 34011 40841
rect 33953 40773 34011 40807
rect 33953 40739 33965 40773
rect 33999 40739 34011 40773
rect 33953 40705 34011 40739
rect 33953 40671 33965 40705
rect 33999 40671 34011 40705
rect 33953 40637 34011 40671
rect 33953 40603 33965 40637
rect 33999 40603 34011 40637
rect 33953 40569 34011 40603
rect 33953 40535 33965 40569
rect 33999 40535 34011 40569
rect 33953 40501 34011 40535
rect 33953 40467 33965 40501
rect 33999 40467 34011 40501
rect 33953 40433 34011 40467
rect 33953 40399 33965 40433
rect 33999 40399 34011 40433
rect 33953 40365 34011 40399
rect 33953 40331 33965 40365
rect 33999 40331 34011 40365
rect 33953 40297 34011 40331
rect 33953 40263 33965 40297
rect 33999 40263 34011 40297
rect 33953 40229 34011 40263
rect 33953 40195 33965 40229
rect 33999 40195 34011 40229
rect 33953 40161 34011 40195
rect 33953 40127 33965 40161
rect 33999 40127 34011 40161
rect 33953 40093 34011 40127
rect 33953 40059 33965 40093
rect 33999 40059 34011 40093
rect 33953 40025 34011 40059
rect 33953 39991 33965 40025
rect 33999 39991 34011 40025
rect 33953 39957 34011 39991
rect 33953 39923 33965 39957
rect 33999 39923 34011 39957
rect 33953 39907 34011 39923
rect 34411 41181 34469 41197
rect 34411 41147 34423 41181
rect 34457 41147 34469 41181
rect 34411 41113 34469 41147
rect 34411 41079 34423 41113
rect 34457 41079 34469 41113
rect 34411 41045 34469 41079
rect 34411 41011 34423 41045
rect 34457 41011 34469 41045
rect 34411 40977 34469 41011
rect 34411 40943 34423 40977
rect 34457 40943 34469 40977
rect 34411 40909 34469 40943
rect 34411 40875 34423 40909
rect 34457 40875 34469 40909
rect 34411 40841 34469 40875
rect 34411 40807 34423 40841
rect 34457 40807 34469 40841
rect 34411 40773 34469 40807
rect 34411 40739 34423 40773
rect 34457 40739 34469 40773
rect 34411 40705 34469 40739
rect 34411 40671 34423 40705
rect 34457 40671 34469 40705
rect 34411 40637 34469 40671
rect 34411 40603 34423 40637
rect 34457 40603 34469 40637
rect 34411 40569 34469 40603
rect 34411 40535 34423 40569
rect 34457 40535 34469 40569
rect 34411 40501 34469 40535
rect 34411 40467 34423 40501
rect 34457 40467 34469 40501
rect 34411 40433 34469 40467
rect 34411 40399 34423 40433
rect 34457 40399 34469 40433
rect 34411 40365 34469 40399
rect 34411 40331 34423 40365
rect 34457 40331 34469 40365
rect 34411 40297 34469 40331
rect 34411 40263 34423 40297
rect 34457 40263 34469 40297
rect 34411 40229 34469 40263
rect 34411 40195 34423 40229
rect 34457 40195 34469 40229
rect 34411 40161 34469 40195
rect 34411 40127 34423 40161
rect 34457 40127 34469 40161
rect 34411 40093 34469 40127
rect 34411 40059 34423 40093
rect 34457 40059 34469 40093
rect 34411 40025 34469 40059
rect 34411 39991 34423 40025
rect 34457 39991 34469 40025
rect 34411 39957 34469 39991
rect 34411 39923 34423 39957
rect 34457 39923 34469 39957
rect 34411 39907 34469 39923
rect 34869 41181 34927 41197
rect 34869 41147 34881 41181
rect 34915 41147 34927 41181
rect 34869 41113 34927 41147
rect 34869 41079 34881 41113
rect 34915 41079 34927 41113
rect 34869 41045 34927 41079
rect 34869 41011 34881 41045
rect 34915 41011 34927 41045
rect 34869 40977 34927 41011
rect 34869 40943 34881 40977
rect 34915 40943 34927 40977
rect 34869 40909 34927 40943
rect 34869 40875 34881 40909
rect 34915 40875 34927 40909
rect 34869 40841 34927 40875
rect 34869 40807 34881 40841
rect 34915 40807 34927 40841
rect 34869 40773 34927 40807
rect 34869 40739 34881 40773
rect 34915 40739 34927 40773
rect 34869 40705 34927 40739
rect 34869 40671 34881 40705
rect 34915 40671 34927 40705
rect 34869 40637 34927 40671
rect 34869 40603 34881 40637
rect 34915 40603 34927 40637
rect 34869 40569 34927 40603
rect 34869 40535 34881 40569
rect 34915 40535 34927 40569
rect 34869 40501 34927 40535
rect 34869 40467 34881 40501
rect 34915 40467 34927 40501
rect 34869 40433 34927 40467
rect 34869 40399 34881 40433
rect 34915 40399 34927 40433
rect 34869 40365 34927 40399
rect 34869 40331 34881 40365
rect 34915 40331 34927 40365
rect 34869 40297 34927 40331
rect 34869 40263 34881 40297
rect 34915 40263 34927 40297
rect 34869 40229 34927 40263
rect 34869 40195 34881 40229
rect 34915 40195 34927 40229
rect 34869 40161 34927 40195
rect 34869 40127 34881 40161
rect 34915 40127 34927 40161
rect 34869 40093 34927 40127
rect 34869 40059 34881 40093
rect 34915 40059 34927 40093
rect 34869 40025 34927 40059
rect 34869 39991 34881 40025
rect 34915 39991 34927 40025
rect 34869 39957 34927 39991
rect 34869 39923 34881 39957
rect 34915 39923 34927 39957
rect 42114 40780 42794 40832
rect 42114 40746 42168 40780
rect 42202 40746 42258 40780
rect 42292 40746 42348 40780
rect 42382 40746 42438 40780
rect 42472 40746 42528 40780
rect 42562 40746 42618 40780
rect 42652 40746 42708 40780
rect 42742 40746 42794 40780
rect 42114 40690 42794 40746
rect 42114 40656 42168 40690
rect 42202 40656 42258 40690
rect 42292 40656 42348 40690
rect 42382 40656 42438 40690
rect 42472 40656 42528 40690
rect 42562 40656 42618 40690
rect 42652 40656 42708 40690
rect 42742 40656 42794 40690
rect 42114 40600 42794 40656
rect 42114 40566 42168 40600
rect 42202 40566 42258 40600
rect 42292 40566 42348 40600
rect 42382 40566 42438 40600
rect 42472 40566 42528 40600
rect 42562 40566 42618 40600
rect 42652 40566 42708 40600
rect 42742 40566 42794 40600
rect 42114 40510 42794 40566
rect 42114 40476 42168 40510
rect 42202 40476 42258 40510
rect 42292 40476 42348 40510
rect 42382 40476 42438 40510
rect 42472 40476 42528 40510
rect 42562 40476 42618 40510
rect 42652 40476 42708 40510
rect 42742 40476 42794 40510
rect 42114 40420 42794 40476
rect 42114 40386 42168 40420
rect 42202 40386 42258 40420
rect 42292 40386 42348 40420
rect 42382 40386 42438 40420
rect 42472 40386 42528 40420
rect 42562 40386 42618 40420
rect 42652 40386 42708 40420
rect 42742 40386 42794 40420
rect 42114 40330 42794 40386
rect 42114 40296 42168 40330
rect 42202 40296 42258 40330
rect 42292 40296 42348 40330
rect 42382 40296 42438 40330
rect 42472 40296 42528 40330
rect 42562 40296 42618 40330
rect 42652 40296 42708 40330
rect 42742 40296 42794 40330
rect 42114 40240 42794 40296
rect 42114 40206 42168 40240
rect 42202 40206 42258 40240
rect 42292 40206 42348 40240
rect 42382 40206 42438 40240
rect 42472 40206 42528 40240
rect 42562 40206 42618 40240
rect 42652 40206 42708 40240
rect 42742 40206 42794 40240
rect 42114 40152 42794 40206
rect 43454 40780 44134 40832
rect 43454 40746 43508 40780
rect 43542 40746 43598 40780
rect 43632 40746 43688 40780
rect 43722 40746 43778 40780
rect 43812 40746 43868 40780
rect 43902 40746 43958 40780
rect 43992 40746 44048 40780
rect 44082 40746 44134 40780
rect 43454 40690 44134 40746
rect 43454 40656 43508 40690
rect 43542 40656 43598 40690
rect 43632 40656 43688 40690
rect 43722 40656 43778 40690
rect 43812 40656 43868 40690
rect 43902 40656 43958 40690
rect 43992 40656 44048 40690
rect 44082 40656 44134 40690
rect 43454 40600 44134 40656
rect 43454 40566 43508 40600
rect 43542 40566 43598 40600
rect 43632 40566 43688 40600
rect 43722 40566 43778 40600
rect 43812 40566 43868 40600
rect 43902 40566 43958 40600
rect 43992 40566 44048 40600
rect 44082 40566 44134 40600
rect 43454 40510 44134 40566
rect 43454 40476 43508 40510
rect 43542 40476 43598 40510
rect 43632 40476 43688 40510
rect 43722 40476 43778 40510
rect 43812 40476 43868 40510
rect 43902 40476 43958 40510
rect 43992 40476 44048 40510
rect 44082 40476 44134 40510
rect 43454 40420 44134 40476
rect 43454 40386 43508 40420
rect 43542 40386 43598 40420
rect 43632 40386 43688 40420
rect 43722 40386 43778 40420
rect 43812 40386 43868 40420
rect 43902 40386 43958 40420
rect 43992 40386 44048 40420
rect 44082 40386 44134 40420
rect 43454 40330 44134 40386
rect 43454 40296 43508 40330
rect 43542 40296 43598 40330
rect 43632 40296 43688 40330
rect 43722 40296 43778 40330
rect 43812 40296 43868 40330
rect 43902 40296 43958 40330
rect 43992 40296 44048 40330
rect 44082 40296 44134 40330
rect 43454 40240 44134 40296
rect 43454 40206 43508 40240
rect 43542 40206 43598 40240
rect 43632 40206 43688 40240
rect 43722 40206 43778 40240
rect 43812 40206 43868 40240
rect 43902 40206 43958 40240
rect 43992 40206 44048 40240
rect 44082 40206 44134 40240
rect 43454 40152 44134 40206
rect 44794 40780 45474 40832
rect 44794 40746 44848 40780
rect 44882 40746 44938 40780
rect 44972 40746 45028 40780
rect 45062 40746 45118 40780
rect 45152 40746 45208 40780
rect 45242 40746 45298 40780
rect 45332 40746 45388 40780
rect 45422 40746 45474 40780
rect 44794 40690 45474 40746
rect 44794 40656 44848 40690
rect 44882 40656 44938 40690
rect 44972 40656 45028 40690
rect 45062 40656 45118 40690
rect 45152 40656 45208 40690
rect 45242 40656 45298 40690
rect 45332 40656 45388 40690
rect 45422 40656 45474 40690
rect 44794 40600 45474 40656
rect 44794 40566 44848 40600
rect 44882 40566 44938 40600
rect 44972 40566 45028 40600
rect 45062 40566 45118 40600
rect 45152 40566 45208 40600
rect 45242 40566 45298 40600
rect 45332 40566 45388 40600
rect 45422 40566 45474 40600
rect 44794 40510 45474 40566
rect 44794 40476 44848 40510
rect 44882 40476 44938 40510
rect 44972 40476 45028 40510
rect 45062 40476 45118 40510
rect 45152 40476 45208 40510
rect 45242 40476 45298 40510
rect 45332 40476 45388 40510
rect 45422 40476 45474 40510
rect 44794 40420 45474 40476
rect 44794 40386 44848 40420
rect 44882 40386 44938 40420
rect 44972 40386 45028 40420
rect 45062 40386 45118 40420
rect 45152 40386 45208 40420
rect 45242 40386 45298 40420
rect 45332 40386 45388 40420
rect 45422 40386 45474 40420
rect 44794 40330 45474 40386
rect 44794 40296 44848 40330
rect 44882 40296 44938 40330
rect 44972 40296 45028 40330
rect 45062 40296 45118 40330
rect 45152 40296 45208 40330
rect 45242 40296 45298 40330
rect 45332 40296 45388 40330
rect 45422 40296 45474 40330
rect 44794 40240 45474 40296
rect 44794 40206 44848 40240
rect 44882 40206 44938 40240
rect 44972 40206 45028 40240
rect 45062 40206 45118 40240
rect 45152 40206 45208 40240
rect 45242 40206 45298 40240
rect 45332 40206 45388 40240
rect 45422 40206 45474 40240
rect 44794 40152 45474 40206
rect 46134 40780 46814 40832
rect 46134 40746 46188 40780
rect 46222 40746 46278 40780
rect 46312 40746 46368 40780
rect 46402 40746 46458 40780
rect 46492 40746 46548 40780
rect 46582 40746 46638 40780
rect 46672 40746 46728 40780
rect 46762 40746 46814 40780
rect 46134 40690 46814 40746
rect 46134 40656 46188 40690
rect 46222 40656 46278 40690
rect 46312 40656 46368 40690
rect 46402 40656 46458 40690
rect 46492 40656 46548 40690
rect 46582 40656 46638 40690
rect 46672 40656 46728 40690
rect 46762 40656 46814 40690
rect 46134 40600 46814 40656
rect 46134 40566 46188 40600
rect 46222 40566 46278 40600
rect 46312 40566 46368 40600
rect 46402 40566 46458 40600
rect 46492 40566 46548 40600
rect 46582 40566 46638 40600
rect 46672 40566 46728 40600
rect 46762 40566 46814 40600
rect 46134 40510 46814 40566
rect 46134 40476 46188 40510
rect 46222 40476 46278 40510
rect 46312 40476 46368 40510
rect 46402 40476 46458 40510
rect 46492 40476 46548 40510
rect 46582 40476 46638 40510
rect 46672 40476 46728 40510
rect 46762 40476 46814 40510
rect 46134 40420 46814 40476
rect 46134 40386 46188 40420
rect 46222 40386 46278 40420
rect 46312 40386 46368 40420
rect 46402 40386 46458 40420
rect 46492 40386 46548 40420
rect 46582 40386 46638 40420
rect 46672 40386 46728 40420
rect 46762 40386 46814 40420
rect 46134 40330 46814 40386
rect 46134 40296 46188 40330
rect 46222 40296 46278 40330
rect 46312 40296 46368 40330
rect 46402 40296 46458 40330
rect 46492 40296 46548 40330
rect 46582 40296 46638 40330
rect 46672 40296 46728 40330
rect 46762 40296 46814 40330
rect 46134 40240 46814 40296
rect 46134 40206 46188 40240
rect 46222 40206 46278 40240
rect 46312 40206 46368 40240
rect 46402 40206 46458 40240
rect 46492 40206 46548 40240
rect 46582 40206 46638 40240
rect 46672 40206 46728 40240
rect 46762 40206 46814 40240
rect 46134 40152 46814 40206
rect 47474 40780 48154 40832
rect 47474 40746 47528 40780
rect 47562 40746 47618 40780
rect 47652 40746 47708 40780
rect 47742 40746 47798 40780
rect 47832 40746 47888 40780
rect 47922 40746 47978 40780
rect 48012 40746 48068 40780
rect 48102 40746 48154 40780
rect 47474 40690 48154 40746
rect 47474 40656 47528 40690
rect 47562 40656 47618 40690
rect 47652 40656 47708 40690
rect 47742 40656 47798 40690
rect 47832 40656 47888 40690
rect 47922 40656 47978 40690
rect 48012 40656 48068 40690
rect 48102 40656 48154 40690
rect 47474 40600 48154 40656
rect 47474 40566 47528 40600
rect 47562 40566 47618 40600
rect 47652 40566 47708 40600
rect 47742 40566 47798 40600
rect 47832 40566 47888 40600
rect 47922 40566 47978 40600
rect 48012 40566 48068 40600
rect 48102 40566 48154 40600
rect 47474 40510 48154 40566
rect 47474 40476 47528 40510
rect 47562 40476 47618 40510
rect 47652 40476 47708 40510
rect 47742 40476 47798 40510
rect 47832 40476 47888 40510
rect 47922 40476 47978 40510
rect 48012 40476 48068 40510
rect 48102 40476 48154 40510
rect 47474 40420 48154 40476
rect 47474 40386 47528 40420
rect 47562 40386 47618 40420
rect 47652 40386 47708 40420
rect 47742 40386 47798 40420
rect 47832 40386 47888 40420
rect 47922 40386 47978 40420
rect 48012 40386 48068 40420
rect 48102 40386 48154 40420
rect 47474 40330 48154 40386
rect 47474 40296 47528 40330
rect 47562 40296 47618 40330
rect 47652 40296 47708 40330
rect 47742 40296 47798 40330
rect 47832 40296 47888 40330
rect 47922 40296 47978 40330
rect 48012 40296 48068 40330
rect 48102 40296 48154 40330
rect 47474 40240 48154 40296
rect 47474 40206 47528 40240
rect 47562 40206 47618 40240
rect 47652 40206 47708 40240
rect 47742 40206 47798 40240
rect 47832 40206 47888 40240
rect 47922 40206 47978 40240
rect 48012 40206 48068 40240
rect 48102 40206 48154 40240
rect 47474 40152 48154 40206
rect 48814 40780 49494 40832
rect 48814 40746 48868 40780
rect 48902 40746 48958 40780
rect 48992 40746 49048 40780
rect 49082 40746 49138 40780
rect 49172 40746 49228 40780
rect 49262 40746 49318 40780
rect 49352 40746 49408 40780
rect 49442 40746 49494 40780
rect 48814 40690 49494 40746
rect 48814 40656 48868 40690
rect 48902 40656 48958 40690
rect 48992 40656 49048 40690
rect 49082 40656 49138 40690
rect 49172 40656 49228 40690
rect 49262 40656 49318 40690
rect 49352 40656 49408 40690
rect 49442 40656 49494 40690
rect 48814 40600 49494 40656
rect 48814 40566 48868 40600
rect 48902 40566 48958 40600
rect 48992 40566 49048 40600
rect 49082 40566 49138 40600
rect 49172 40566 49228 40600
rect 49262 40566 49318 40600
rect 49352 40566 49408 40600
rect 49442 40566 49494 40600
rect 48814 40510 49494 40566
rect 48814 40476 48868 40510
rect 48902 40476 48958 40510
rect 48992 40476 49048 40510
rect 49082 40476 49138 40510
rect 49172 40476 49228 40510
rect 49262 40476 49318 40510
rect 49352 40476 49408 40510
rect 49442 40476 49494 40510
rect 48814 40420 49494 40476
rect 48814 40386 48868 40420
rect 48902 40386 48958 40420
rect 48992 40386 49048 40420
rect 49082 40386 49138 40420
rect 49172 40386 49228 40420
rect 49262 40386 49318 40420
rect 49352 40386 49408 40420
rect 49442 40386 49494 40420
rect 48814 40330 49494 40386
rect 48814 40296 48868 40330
rect 48902 40296 48958 40330
rect 48992 40296 49048 40330
rect 49082 40296 49138 40330
rect 49172 40296 49228 40330
rect 49262 40296 49318 40330
rect 49352 40296 49408 40330
rect 49442 40296 49494 40330
rect 48814 40240 49494 40296
rect 48814 40206 48868 40240
rect 48902 40206 48958 40240
rect 48992 40206 49048 40240
rect 49082 40206 49138 40240
rect 49172 40206 49228 40240
rect 49262 40206 49318 40240
rect 49352 40206 49408 40240
rect 49442 40206 49494 40240
rect 48814 40152 49494 40206
rect 50154 40780 50834 40832
rect 50154 40746 50208 40780
rect 50242 40746 50298 40780
rect 50332 40746 50388 40780
rect 50422 40746 50478 40780
rect 50512 40746 50568 40780
rect 50602 40746 50658 40780
rect 50692 40746 50748 40780
rect 50782 40746 50834 40780
rect 50154 40690 50834 40746
rect 50154 40656 50208 40690
rect 50242 40656 50298 40690
rect 50332 40656 50388 40690
rect 50422 40656 50478 40690
rect 50512 40656 50568 40690
rect 50602 40656 50658 40690
rect 50692 40656 50748 40690
rect 50782 40656 50834 40690
rect 50154 40600 50834 40656
rect 50154 40566 50208 40600
rect 50242 40566 50298 40600
rect 50332 40566 50388 40600
rect 50422 40566 50478 40600
rect 50512 40566 50568 40600
rect 50602 40566 50658 40600
rect 50692 40566 50748 40600
rect 50782 40566 50834 40600
rect 50154 40510 50834 40566
rect 50154 40476 50208 40510
rect 50242 40476 50298 40510
rect 50332 40476 50388 40510
rect 50422 40476 50478 40510
rect 50512 40476 50568 40510
rect 50602 40476 50658 40510
rect 50692 40476 50748 40510
rect 50782 40476 50834 40510
rect 50154 40420 50834 40476
rect 50154 40386 50208 40420
rect 50242 40386 50298 40420
rect 50332 40386 50388 40420
rect 50422 40386 50478 40420
rect 50512 40386 50568 40420
rect 50602 40386 50658 40420
rect 50692 40386 50748 40420
rect 50782 40386 50834 40420
rect 50154 40330 50834 40386
rect 50154 40296 50208 40330
rect 50242 40296 50298 40330
rect 50332 40296 50388 40330
rect 50422 40296 50478 40330
rect 50512 40296 50568 40330
rect 50602 40296 50658 40330
rect 50692 40296 50748 40330
rect 50782 40296 50834 40330
rect 50154 40240 50834 40296
rect 50154 40206 50208 40240
rect 50242 40206 50298 40240
rect 50332 40206 50388 40240
rect 50422 40206 50478 40240
rect 50512 40206 50568 40240
rect 50602 40206 50658 40240
rect 50692 40206 50748 40240
rect 50782 40206 50834 40240
rect 50154 40152 50834 40206
rect 51494 40780 52174 40832
rect 51494 40746 51548 40780
rect 51582 40746 51638 40780
rect 51672 40746 51728 40780
rect 51762 40746 51818 40780
rect 51852 40746 51908 40780
rect 51942 40746 51998 40780
rect 52032 40746 52088 40780
rect 52122 40746 52174 40780
rect 51494 40690 52174 40746
rect 51494 40656 51548 40690
rect 51582 40656 51638 40690
rect 51672 40656 51728 40690
rect 51762 40656 51818 40690
rect 51852 40656 51908 40690
rect 51942 40656 51998 40690
rect 52032 40656 52088 40690
rect 52122 40656 52174 40690
rect 51494 40600 52174 40656
rect 51494 40566 51548 40600
rect 51582 40566 51638 40600
rect 51672 40566 51728 40600
rect 51762 40566 51818 40600
rect 51852 40566 51908 40600
rect 51942 40566 51998 40600
rect 52032 40566 52088 40600
rect 52122 40566 52174 40600
rect 51494 40510 52174 40566
rect 51494 40476 51548 40510
rect 51582 40476 51638 40510
rect 51672 40476 51728 40510
rect 51762 40476 51818 40510
rect 51852 40476 51908 40510
rect 51942 40476 51998 40510
rect 52032 40476 52088 40510
rect 52122 40476 52174 40510
rect 51494 40420 52174 40476
rect 51494 40386 51548 40420
rect 51582 40386 51638 40420
rect 51672 40386 51728 40420
rect 51762 40386 51818 40420
rect 51852 40386 51908 40420
rect 51942 40386 51998 40420
rect 52032 40386 52088 40420
rect 52122 40386 52174 40420
rect 51494 40330 52174 40386
rect 51494 40296 51548 40330
rect 51582 40296 51638 40330
rect 51672 40296 51728 40330
rect 51762 40296 51818 40330
rect 51852 40296 51908 40330
rect 51942 40296 51998 40330
rect 52032 40296 52088 40330
rect 52122 40296 52174 40330
rect 51494 40240 52174 40296
rect 51494 40206 51548 40240
rect 51582 40206 51638 40240
rect 51672 40206 51728 40240
rect 51762 40206 51818 40240
rect 51852 40206 51908 40240
rect 51942 40206 51998 40240
rect 52032 40206 52088 40240
rect 52122 40206 52174 40240
rect 51494 40152 52174 40206
rect 34869 39907 34927 39923
rect 12322 37020 13002 37072
rect 12322 36986 12376 37020
rect 12410 36986 12466 37020
rect 12500 36986 12556 37020
rect 12590 36986 12646 37020
rect 12680 36986 12736 37020
rect 12770 36986 12826 37020
rect 12860 36986 12916 37020
rect 12950 36986 13002 37020
rect 12322 36930 13002 36986
rect 12322 36896 12376 36930
rect 12410 36896 12466 36930
rect 12500 36896 12556 36930
rect 12590 36896 12646 36930
rect 12680 36896 12736 36930
rect 12770 36896 12826 36930
rect 12860 36896 12916 36930
rect 12950 36896 13002 36930
rect 12322 36840 13002 36896
rect 12322 36806 12376 36840
rect 12410 36806 12466 36840
rect 12500 36806 12556 36840
rect 12590 36806 12646 36840
rect 12680 36806 12736 36840
rect 12770 36806 12826 36840
rect 12860 36806 12916 36840
rect 12950 36806 13002 36840
rect 12322 36750 13002 36806
rect 12322 36716 12376 36750
rect 12410 36716 12466 36750
rect 12500 36716 12556 36750
rect 12590 36716 12646 36750
rect 12680 36716 12736 36750
rect 12770 36716 12826 36750
rect 12860 36716 12916 36750
rect 12950 36716 13002 36750
rect 12322 36660 13002 36716
rect 12322 36626 12376 36660
rect 12410 36626 12466 36660
rect 12500 36626 12556 36660
rect 12590 36626 12646 36660
rect 12680 36626 12736 36660
rect 12770 36626 12826 36660
rect 12860 36626 12916 36660
rect 12950 36626 13002 36660
rect 12322 36570 13002 36626
rect 12322 36536 12376 36570
rect 12410 36536 12466 36570
rect 12500 36536 12556 36570
rect 12590 36536 12646 36570
rect 12680 36536 12736 36570
rect 12770 36536 12826 36570
rect 12860 36536 12916 36570
rect 12950 36536 13002 36570
rect 12322 36480 13002 36536
rect 12322 36446 12376 36480
rect 12410 36446 12466 36480
rect 12500 36446 12556 36480
rect 12590 36446 12646 36480
rect 12680 36446 12736 36480
rect 12770 36446 12826 36480
rect 12860 36446 12916 36480
rect 12950 36446 13002 36480
rect 12322 36392 13002 36446
rect 37507 37421 37565 37437
rect 37507 37387 37519 37421
rect 37553 37387 37565 37421
rect 37507 37353 37565 37387
rect 37507 37319 37519 37353
rect 37553 37319 37565 37353
rect 37507 37285 37565 37319
rect 37507 37251 37519 37285
rect 37553 37251 37565 37285
rect 37507 37217 37565 37251
rect 37507 37183 37519 37217
rect 37553 37183 37565 37217
rect 37507 37149 37565 37183
rect 37507 37115 37519 37149
rect 37553 37115 37565 37149
rect 37507 37081 37565 37115
rect 37507 37047 37519 37081
rect 37553 37047 37565 37081
rect 37507 37013 37565 37047
rect 37507 36979 37519 37013
rect 37553 36979 37565 37013
rect 37507 36945 37565 36979
rect 37507 36911 37519 36945
rect 37553 36911 37565 36945
rect 37507 36877 37565 36911
rect 37507 36843 37519 36877
rect 37553 36843 37565 36877
rect 37507 36809 37565 36843
rect 37507 36775 37519 36809
rect 37553 36775 37565 36809
rect 37507 36741 37565 36775
rect 37507 36707 37519 36741
rect 37553 36707 37565 36741
rect 37507 36673 37565 36707
rect 37507 36639 37519 36673
rect 37553 36639 37565 36673
rect 37507 36605 37565 36639
rect 37507 36571 37519 36605
rect 37553 36571 37565 36605
rect 37507 36537 37565 36571
rect 37507 36503 37519 36537
rect 37553 36503 37565 36537
rect 37507 36469 37565 36503
rect 37507 36435 37519 36469
rect 37553 36435 37565 36469
rect 37507 36401 37565 36435
rect 37507 36367 37519 36401
rect 37553 36367 37565 36401
rect 37507 36333 37565 36367
rect 37507 36299 37519 36333
rect 37553 36299 37565 36333
rect 37507 36265 37565 36299
rect 37507 36231 37519 36265
rect 37553 36231 37565 36265
rect 37507 36197 37565 36231
rect 37507 36163 37519 36197
rect 37553 36163 37565 36197
rect 37507 36147 37565 36163
rect 37965 37421 38023 37437
rect 37965 37387 37977 37421
rect 38011 37387 38023 37421
rect 37965 37353 38023 37387
rect 37965 37319 37977 37353
rect 38011 37319 38023 37353
rect 37965 37285 38023 37319
rect 37965 37251 37977 37285
rect 38011 37251 38023 37285
rect 37965 37217 38023 37251
rect 37965 37183 37977 37217
rect 38011 37183 38023 37217
rect 37965 37149 38023 37183
rect 37965 37115 37977 37149
rect 38011 37115 38023 37149
rect 37965 37081 38023 37115
rect 37965 37047 37977 37081
rect 38011 37047 38023 37081
rect 37965 37013 38023 37047
rect 37965 36979 37977 37013
rect 38011 36979 38023 37013
rect 37965 36945 38023 36979
rect 37965 36911 37977 36945
rect 38011 36911 38023 36945
rect 37965 36877 38023 36911
rect 37965 36843 37977 36877
rect 38011 36843 38023 36877
rect 37965 36809 38023 36843
rect 37965 36775 37977 36809
rect 38011 36775 38023 36809
rect 37965 36741 38023 36775
rect 37965 36707 37977 36741
rect 38011 36707 38023 36741
rect 37965 36673 38023 36707
rect 37965 36639 37977 36673
rect 38011 36639 38023 36673
rect 37965 36605 38023 36639
rect 37965 36571 37977 36605
rect 38011 36571 38023 36605
rect 37965 36537 38023 36571
rect 37965 36503 37977 36537
rect 38011 36503 38023 36537
rect 37965 36469 38023 36503
rect 37965 36435 37977 36469
rect 38011 36435 38023 36469
rect 37965 36401 38023 36435
rect 37965 36367 37977 36401
rect 38011 36367 38023 36401
rect 37965 36333 38023 36367
rect 37965 36299 37977 36333
rect 38011 36299 38023 36333
rect 37965 36265 38023 36299
rect 37965 36231 37977 36265
rect 38011 36231 38023 36265
rect 37965 36197 38023 36231
rect 37965 36163 37977 36197
rect 38011 36163 38023 36197
rect 37965 36147 38023 36163
rect 38423 37421 38481 37437
rect 38423 37387 38435 37421
rect 38469 37387 38481 37421
rect 38423 37353 38481 37387
rect 38423 37319 38435 37353
rect 38469 37319 38481 37353
rect 38423 37285 38481 37319
rect 38423 37251 38435 37285
rect 38469 37251 38481 37285
rect 38423 37217 38481 37251
rect 38423 37183 38435 37217
rect 38469 37183 38481 37217
rect 38423 37149 38481 37183
rect 38423 37115 38435 37149
rect 38469 37115 38481 37149
rect 38423 37081 38481 37115
rect 38423 37047 38435 37081
rect 38469 37047 38481 37081
rect 38423 37013 38481 37047
rect 38423 36979 38435 37013
rect 38469 36979 38481 37013
rect 38423 36945 38481 36979
rect 38423 36911 38435 36945
rect 38469 36911 38481 36945
rect 38423 36877 38481 36911
rect 38423 36843 38435 36877
rect 38469 36843 38481 36877
rect 38423 36809 38481 36843
rect 38423 36775 38435 36809
rect 38469 36775 38481 36809
rect 38423 36741 38481 36775
rect 38423 36707 38435 36741
rect 38469 36707 38481 36741
rect 38423 36673 38481 36707
rect 38423 36639 38435 36673
rect 38469 36639 38481 36673
rect 38423 36605 38481 36639
rect 38423 36571 38435 36605
rect 38469 36571 38481 36605
rect 38423 36537 38481 36571
rect 38423 36503 38435 36537
rect 38469 36503 38481 36537
rect 38423 36469 38481 36503
rect 38423 36435 38435 36469
rect 38469 36435 38481 36469
rect 38423 36401 38481 36435
rect 38423 36367 38435 36401
rect 38469 36367 38481 36401
rect 38423 36333 38481 36367
rect 38423 36299 38435 36333
rect 38469 36299 38481 36333
rect 38423 36265 38481 36299
rect 38423 36231 38435 36265
rect 38469 36231 38481 36265
rect 38423 36197 38481 36231
rect 38423 36163 38435 36197
rect 38469 36163 38481 36197
rect 38423 36147 38481 36163
rect 38881 37421 38939 37437
rect 38881 37387 38893 37421
rect 38927 37387 38939 37421
rect 38881 37353 38939 37387
rect 38881 37319 38893 37353
rect 38927 37319 38939 37353
rect 38881 37285 38939 37319
rect 38881 37251 38893 37285
rect 38927 37251 38939 37285
rect 38881 37217 38939 37251
rect 38881 37183 38893 37217
rect 38927 37183 38939 37217
rect 38881 37149 38939 37183
rect 38881 37115 38893 37149
rect 38927 37115 38939 37149
rect 38881 37081 38939 37115
rect 38881 37047 38893 37081
rect 38927 37047 38939 37081
rect 38881 37013 38939 37047
rect 38881 36979 38893 37013
rect 38927 36979 38939 37013
rect 38881 36945 38939 36979
rect 38881 36911 38893 36945
rect 38927 36911 38939 36945
rect 38881 36877 38939 36911
rect 38881 36843 38893 36877
rect 38927 36843 38939 36877
rect 38881 36809 38939 36843
rect 38881 36775 38893 36809
rect 38927 36775 38939 36809
rect 38881 36741 38939 36775
rect 38881 36707 38893 36741
rect 38927 36707 38939 36741
rect 38881 36673 38939 36707
rect 38881 36639 38893 36673
rect 38927 36639 38939 36673
rect 38881 36605 38939 36639
rect 38881 36571 38893 36605
rect 38927 36571 38939 36605
rect 38881 36537 38939 36571
rect 38881 36503 38893 36537
rect 38927 36503 38939 36537
rect 38881 36469 38939 36503
rect 38881 36435 38893 36469
rect 38927 36435 38939 36469
rect 38881 36401 38939 36435
rect 38881 36367 38893 36401
rect 38927 36367 38939 36401
rect 38881 36333 38939 36367
rect 38881 36299 38893 36333
rect 38927 36299 38939 36333
rect 38881 36265 38939 36299
rect 38881 36231 38893 36265
rect 38927 36231 38939 36265
rect 38881 36197 38939 36231
rect 38881 36163 38893 36197
rect 38927 36163 38939 36197
rect 38881 36147 38939 36163
rect 39339 37421 39397 37437
rect 39339 37387 39351 37421
rect 39385 37387 39397 37421
rect 39339 37353 39397 37387
rect 39339 37319 39351 37353
rect 39385 37319 39397 37353
rect 39339 37285 39397 37319
rect 39339 37251 39351 37285
rect 39385 37251 39397 37285
rect 39339 37217 39397 37251
rect 39339 37183 39351 37217
rect 39385 37183 39397 37217
rect 39339 37149 39397 37183
rect 39339 37115 39351 37149
rect 39385 37115 39397 37149
rect 39339 37081 39397 37115
rect 39339 37047 39351 37081
rect 39385 37047 39397 37081
rect 39339 37013 39397 37047
rect 39339 36979 39351 37013
rect 39385 36979 39397 37013
rect 39339 36945 39397 36979
rect 39339 36911 39351 36945
rect 39385 36911 39397 36945
rect 39339 36877 39397 36911
rect 39339 36843 39351 36877
rect 39385 36843 39397 36877
rect 39339 36809 39397 36843
rect 39339 36775 39351 36809
rect 39385 36775 39397 36809
rect 39339 36741 39397 36775
rect 39339 36707 39351 36741
rect 39385 36707 39397 36741
rect 39339 36673 39397 36707
rect 39339 36639 39351 36673
rect 39385 36639 39397 36673
rect 39339 36605 39397 36639
rect 39339 36571 39351 36605
rect 39385 36571 39397 36605
rect 39339 36537 39397 36571
rect 39339 36503 39351 36537
rect 39385 36503 39397 36537
rect 39339 36469 39397 36503
rect 39339 36435 39351 36469
rect 39385 36435 39397 36469
rect 39339 36401 39397 36435
rect 39339 36367 39351 36401
rect 39385 36367 39397 36401
rect 39339 36333 39397 36367
rect 39339 36299 39351 36333
rect 39385 36299 39397 36333
rect 39339 36265 39397 36299
rect 39339 36231 39351 36265
rect 39385 36231 39397 36265
rect 39339 36197 39397 36231
rect 39339 36163 39351 36197
rect 39385 36163 39397 36197
rect 39339 36147 39397 36163
rect 39797 37421 39855 37437
rect 39797 37387 39809 37421
rect 39843 37387 39855 37421
rect 39797 37353 39855 37387
rect 39797 37319 39809 37353
rect 39843 37319 39855 37353
rect 39797 37285 39855 37319
rect 39797 37251 39809 37285
rect 39843 37251 39855 37285
rect 39797 37217 39855 37251
rect 39797 37183 39809 37217
rect 39843 37183 39855 37217
rect 39797 37149 39855 37183
rect 39797 37115 39809 37149
rect 39843 37115 39855 37149
rect 39797 37081 39855 37115
rect 39797 37047 39809 37081
rect 39843 37047 39855 37081
rect 39797 37013 39855 37047
rect 39797 36979 39809 37013
rect 39843 36979 39855 37013
rect 39797 36945 39855 36979
rect 39797 36911 39809 36945
rect 39843 36911 39855 36945
rect 39797 36877 39855 36911
rect 39797 36843 39809 36877
rect 39843 36843 39855 36877
rect 39797 36809 39855 36843
rect 39797 36775 39809 36809
rect 39843 36775 39855 36809
rect 39797 36741 39855 36775
rect 39797 36707 39809 36741
rect 39843 36707 39855 36741
rect 39797 36673 39855 36707
rect 39797 36639 39809 36673
rect 39843 36639 39855 36673
rect 39797 36605 39855 36639
rect 39797 36571 39809 36605
rect 39843 36571 39855 36605
rect 39797 36537 39855 36571
rect 39797 36503 39809 36537
rect 39843 36503 39855 36537
rect 39797 36469 39855 36503
rect 39797 36435 39809 36469
rect 39843 36435 39855 36469
rect 39797 36401 39855 36435
rect 39797 36367 39809 36401
rect 39843 36367 39855 36401
rect 39797 36333 39855 36367
rect 39797 36299 39809 36333
rect 39843 36299 39855 36333
rect 39797 36265 39855 36299
rect 39797 36231 39809 36265
rect 39843 36231 39855 36265
rect 39797 36197 39855 36231
rect 39797 36163 39809 36197
rect 39843 36163 39855 36197
rect 39797 36147 39855 36163
rect 40255 37421 40313 37437
rect 40255 37387 40267 37421
rect 40301 37387 40313 37421
rect 40255 37353 40313 37387
rect 40255 37319 40267 37353
rect 40301 37319 40313 37353
rect 40255 37285 40313 37319
rect 40255 37251 40267 37285
rect 40301 37251 40313 37285
rect 40255 37217 40313 37251
rect 40255 37183 40267 37217
rect 40301 37183 40313 37217
rect 40255 37149 40313 37183
rect 40255 37115 40267 37149
rect 40301 37115 40313 37149
rect 40255 37081 40313 37115
rect 40255 37047 40267 37081
rect 40301 37047 40313 37081
rect 40255 37013 40313 37047
rect 40255 36979 40267 37013
rect 40301 36979 40313 37013
rect 40255 36945 40313 36979
rect 40255 36911 40267 36945
rect 40301 36911 40313 36945
rect 40255 36877 40313 36911
rect 40255 36843 40267 36877
rect 40301 36843 40313 36877
rect 40255 36809 40313 36843
rect 40255 36775 40267 36809
rect 40301 36775 40313 36809
rect 40255 36741 40313 36775
rect 40255 36707 40267 36741
rect 40301 36707 40313 36741
rect 40255 36673 40313 36707
rect 40255 36639 40267 36673
rect 40301 36639 40313 36673
rect 40255 36605 40313 36639
rect 40255 36571 40267 36605
rect 40301 36571 40313 36605
rect 40255 36537 40313 36571
rect 40255 36503 40267 36537
rect 40301 36503 40313 36537
rect 40255 36469 40313 36503
rect 40255 36435 40267 36469
rect 40301 36435 40313 36469
rect 40255 36401 40313 36435
rect 40255 36367 40267 36401
rect 40301 36367 40313 36401
rect 40255 36333 40313 36367
rect 40255 36299 40267 36333
rect 40301 36299 40313 36333
rect 40255 36265 40313 36299
rect 40255 36231 40267 36265
rect 40301 36231 40313 36265
rect 40255 36197 40313 36231
rect 40255 36163 40267 36197
rect 40301 36163 40313 36197
rect 40255 36147 40313 36163
rect 42114 37020 42794 37072
rect 42114 36986 42168 37020
rect 42202 36986 42258 37020
rect 42292 36986 42348 37020
rect 42382 36986 42438 37020
rect 42472 36986 42528 37020
rect 42562 36986 42618 37020
rect 42652 36986 42708 37020
rect 42742 36986 42794 37020
rect 42114 36930 42794 36986
rect 42114 36896 42168 36930
rect 42202 36896 42258 36930
rect 42292 36896 42348 36930
rect 42382 36896 42438 36930
rect 42472 36896 42528 36930
rect 42562 36896 42618 36930
rect 42652 36896 42708 36930
rect 42742 36896 42794 36930
rect 42114 36840 42794 36896
rect 42114 36806 42168 36840
rect 42202 36806 42258 36840
rect 42292 36806 42348 36840
rect 42382 36806 42438 36840
rect 42472 36806 42528 36840
rect 42562 36806 42618 36840
rect 42652 36806 42708 36840
rect 42742 36806 42794 36840
rect 42114 36750 42794 36806
rect 42114 36716 42168 36750
rect 42202 36716 42258 36750
rect 42292 36716 42348 36750
rect 42382 36716 42438 36750
rect 42472 36716 42528 36750
rect 42562 36716 42618 36750
rect 42652 36716 42708 36750
rect 42742 36716 42794 36750
rect 42114 36660 42794 36716
rect 42114 36626 42168 36660
rect 42202 36626 42258 36660
rect 42292 36626 42348 36660
rect 42382 36626 42438 36660
rect 42472 36626 42528 36660
rect 42562 36626 42618 36660
rect 42652 36626 42708 36660
rect 42742 36626 42794 36660
rect 42114 36570 42794 36626
rect 42114 36536 42168 36570
rect 42202 36536 42258 36570
rect 42292 36536 42348 36570
rect 42382 36536 42438 36570
rect 42472 36536 42528 36570
rect 42562 36536 42618 36570
rect 42652 36536 42708 36570
rect 42742 36536 42794 36570
rect 42114 36480 42794 36536
rect 42114 36446 42168 36480
rect 42202 36446 42258 36480
rect 42292 36446 42348 36480
rect 42382 36446 42438 36480
rect 42472 36446 42528 36480
rect 42562 36446 42618 36480
rect 42652 36446 42708 36480
rect 42742 36446 42794 36480
rect 42114 36392 42794 36446
rect 43454 37020 44134 37072
rect 43454 36986 43508 37020
rect 43542 36986 43598 37020
rect 43632 36986 43688 37020
rect 43722 36986 43778 37020
rect 43812 36986 43868 37020
rect 43902 36986 43958 37020
rect 43992 36986 44048 37020
rect 44082 36986 44134 37020
rect 43454 36930 44134 36986
rect 43454 36896 43508 36930
rect 43542 36896 43598 36930
rect 43632 36896 43688 36930
rect 43722 36896 43778 36930
rect 43812 36896 43868 36930
rect 43902 36896 43958 36930
rect 43992 36896 44048 36930
rect 44082 36896 44134 36930
rect 43454 36840 44134 36896
rect 43454 36806 43508 36840
rect 43542 36806 43598 36840
rect 43632 36806 43688 36840
rect 43722 36806 43778 36840
rect 43812 36806 43868 36840
rect 43902 36806 43958 36840
rect 43992 36806 44048 36840
rect 44082 36806 44134 36840
rect 43454 36750 44134 36806
rect 43454 36716 43508 36750
rect 43542 36716 43598 36750
rect 43632 36716 43688 36750
rect 43722 36716 43778 36750
rect 43812 36716 43868 36750
rect 43902 36716 43958 36750
rect 43992 36716 44048 36750
rect 44082 36716 44134 36750
rect 43454 36660 44134 36716
rect 43454 36626 43508 36660
rect 43542 36626 43598 36660
rect 43632 36626 43688 36660
rect 43722 36626 43778 36660
rect 43812 36626 43868 36660
rect 43902 36626 43958 36660
rect 43992 36626 44048 36660
rect 44082 36626 44134 36660
rect 43454 36570 44134 36626
rect 43454 36536 43508 36570
rect 43542 36536 43598 36570
rect 43632 36536 43688 36570
rect 43722 36536 43778 36570
rect 43812 36536 43868 36570
rect 43902 36536 43958 36570
rect 43992 36536 44048 36570
rect 44082 36536 44134 36570
rect 43454 36480 44134 36536
rect 43454 36446 43508 36480
rect 43542 36446 43598 36480
rect 43632 36446 43688 36480
rect 43722 36446 43778 36480
rect 43812 36446 43868 36480
rect 43902 36446 43958 36480
rect 43992 36446 44048 36480
rect 44082 36446 44134 36480
rect 43454 36392 44134 36446
rect 44794 37020 45474 37072
rect 44794 36986 44848 37020
rect 44882 36986 44938 37020
rect 44972 36986 45028 37020
rect 45062 36986 45118 37020
rect 45152 36986 45208 37020
rect 45242 36986 45298 37020
rect 45332 36986 45388 37020
rect 45422 36986 45474 37020
rect 44794 36930 45474 36986
rect 44794 36896 44848 36930
rect 44882 36896 44938 36930
rect 44972 36896 45028 36930
rect 45062 36896 45118 36930
rect 45152 36896 45208 36930
rect 45242 36896 45298 36930
rect 45332 36896 45388 36930
rect 45422 36896 45474 36930
rect 44794 36840 45474 36896
rect 44794 36806 44848 36840
rect 44882 36806 44938 36840
rect 44972 36806 45028 36840
rect 45062 36806 45118 36840
rect 45152 36806 45208 36840
rect 45242 36806 45298 36840
rect 45332 36806 45388 36840
rect 45422 36806 45474 36840
rect 44794 36750 45474 36806
rect 44794 36716 44848 36750
rect 44882 36716 44938 36750
rect 44972 36716 45028 36750
rect 45062 36716 45118 36750
rect 45152 36716 45208 36750
rect 45242 36716 45298 36750
rect 45332 36716 45388 36750
rect 45422 36716 45474 36750
rect 44794 36660 45474 36716
rect 44794 36626 44848 36660
rect 44882 36626 44938 36660
rect 44972 36626 45028 36660
rect 45062 36626 45118 36660
rect 45152 36626 45208 36660
rect 45242 36626 45298 36660
rect 45332 36626 45388 36660
rect 45422 36626 45474 36660
rect 44794 36570 45474 36626
rect 44794 36536 44848 36570
rect 44882 36536 44938 36570
rect 44972 36536 45028 36570
rect 45062 36536 45118 36570
rect 45152 36536 45208 36570
rect 45242 36536 45298 36570
rect 45332 36536 45388 36570
rect 45422 36536 45474 36570
rect 44794 36480 45474 36536
rect 44794 36446 44848 36480
rect 44882 36446 44938 36480
rect 44972 36446 45028 36480
rect 45062 36446 45118 36480
rect 45152 36446 45208 36480
rect 45242 36446 45298 36480
rect 45332 36446 45388 36480
rect 45422 36446 45474 36480
rect 44794 36392 45474 36446
rect 46134 37020 46814 37072
rect 46134 36986 46188 37020
rect 46222 36986 46278 37020
rect 46312 36986 46368 37020
rect 46402 36986 46458 37020
rect 46492 36986 46548 37020
rect 46582 36986 46638 37020
rect 46672 36986 46728 37020
rect 46762 36986 46814 37020
rect 46134 36930 46814 36986
rect 46134 36896 46188 36930
rect 46222 36896 46278 36930
rect 46312 36896 46368 36930
rect 46402 36896 46458 36930
rect 46492 36896 46548 36930
rect 46582 36896 46638 36930
rect 46672 36896 46728 36930
rect 46762 36896 46814 36930
rect 46134 36840 46814 36896
rect 46134 36806 46188 36840
rect 46222 36806 46278 36840
rect 46312 36806 46368 36840
rect 46402 36806 46458 36840
rect 46492 36806 46548 36840
rect 46582 36806 46638 36840
rect 46672 36806 46728 36840
rect 46762 36806 46814 36840
rect 46134 36750 46814 36806
rect 46134 36716 46188 36750
rect 46222 36716 46278 36750
rect 46312 36716 46368 36750
rect 46402 36716 46458 36750
rect 46492 36716 46548 36750
rect 46582 36716 46638 36750
rect 46672 36716 46728 36750
rect 46762 36716 46814 36750
rect 46134 36660 46814 36716
rect 46134 36626 46188 36660
rect 46222 36626 46278 36660
rect 46312 36626 46368 36660
rect 46402 36626 46458 36660
rect 46492 36626 46548 36660
rect 46582 36626 46638 36660
rect 46672 36626 46728 36660
rect 46762 36626 46814 36660
rect 46134 36570 46814 36626
rect 46134 36536 46188 36570
rect 46222 36536 46278 36570
rect 46312 36536 46368 36570
rect 46402 36536 46458 36570
rect 46492 36536 46548 36570
rect 46582 36536 46638 36570
rect 46672 36536 46728 36570
rect 46762 36536 46814 36570
rect 46134 36480 46814 36536
rect 46134 36446 46188 36480
rect 46222 36446 46278 36480
rect 46312 36446 46368 36480
rect 46402 36446 46458 36480
rect 46492 36446 46548 36480
rect 46582 36446 46638 36480
rect 46672 36446 46728 36480
rect 46762 36446 46814 36480
rect 46134 36392 46814 36446
rect 47474 37020 48154 37072
rect 47474 36986 47528 37020
rect 47562 36986 47618 37020
rect 47652 36986 47708 37020
rect 47742 36986 47798 37020
rect 47832 36986 47888 37020
rect 47922 36986 47978 37020
rect 48012 36986 48068 37020
rect 48102 36986 48154 37020
rect 47474 36930 48154 36986
rect 47474 36896 47528 36930
rect 47562 36896 47618 36930
rect 47652 36896 47708 36930
rect 47742 36896 47798 36930
rect 47832 36896 47888 36930
rect 47922 36896 47978 36930
rect 48012 36896 48068 36930
rect 48102 36896 48154 36930
rect 47474 36840 48154 36896
rect 47474 36806 47528 36840
rect 47562 36806 47618 36840
rect 47652 36806 47708 36840
rect 47742 36806 47798 36840
rect 47832 36806 47888 36840
rect 47922 36806 47978 36840
rect 48012 36806 48068 36840
rect 48102 36806 48154 36840
rect 47474 36750 48154 36806
rect 47474 36716 47528 36750
rect 47562 36716 47618 36750
rect 47652 36716 47708 36750
rect 47742 36716 47798 36750
rect 47832 36716 47888 36750
rect 47922 36716 47978 36750
rect 48012 36716 48068 36750
rect 48102 36716 48154 36750
rect 47474 36660 48154 36716
rect 47474 36626 47528 36660
rect 47562 36626 47618 36660
rect 47652 36626 47708 36660
rect 47742 36626 47798 36660
rect 47832 36626 47888 36660
rect 47922 36626 47978 36660
rect 48012 36626 48068 36660
rect 48102 36626 48154 36660
rect 47474 36570 48154 36626
rect 47474 36536 47528 36570
rect 47562 36536 47618 36570
rect 47652 36536 47708 36570
rect 47742 36536 47798 36570
rect 47832 36536 47888 36570
rect 47922 36536 47978 36570
rect 48012 36536 48068 36570
rect 48102 36536 48154 36570
rect 47474 36480 48154 36536
rect 47474 36446 47528 36480
rect 47562 36446 47618 36480
rect 47652 36446 47708 36480
rect 47742 36446 47798 36480
rect 47832 36446 47888 36480
rect 47922 36446 47978 36480
rect 48012 36446 48068 36480
rect 48102 36446 48154 36480
rect 47474 36392 48154 36446
rect 48814 37020 49494 37072
rect 48814 36986 48868 37020
rect 48902 36986 48958 37020
rect 48992 36986 49048 37020
rect 49082 36986 49138 37020
rect 49172 36986 49228 37020
rect 49262 36986 49318 37020
rect 49352 36986 49408 37020
rect 49442 36986 49494 37020
rect 48814 36930 49494 36986
rect 48814 36896 48868 36930
rect 48902 36896 48958 36930
rect 48992 36896 49048 36930
rect 49082 36896 49138 36930
rect 49172 36896 49228 36930
rect 49262 36896 49318 36930
rect 49352 36896 49408 36930
rect 49442 36896 49494 36930
rect 48814 36840 49494 36896
rect 48814 36806 48868 36840
rect 48902 36806 48958 36840
rect 48992 36806 49048 36840
rect 49082 36806 49138 36840
rect 49172 36806 49228 36840
rect 49262 36806 49318 36840
rect 49352 36806 49408 36840
rect 49442 36806 49494 36840
rect 48814 36750 49494 36806
rect 48814 36716 48868 36750
rect 48902 36716 48958 36750
rect 48992 36716 49048 36750
rect 49082 36716 49138 36750
rect 49172 36716 49228 36750
rect 49262 36716 49318 36750
rect 49352 36716 49408 36750
rect 49442 36716 49494 36750
rect 48814 36660 49494 36716
rect 48814 36626 48868 36660
rect 48902 36626 48958 36660
rect 48992 36626 49048 36660
rect 49082 36626 49138 36660
rect 49172 36626 49228 36660
rect 49262 36626 49318 36660
rect 49352 36626 49408 36660
rect 49442 36626 49494 36660
rect 48814 36570 49494 36626
rect 48814 36536 48868 36570
rect 48902 36536 48958 36570
rect 48992 36536 49048 36570
rect 49082 36536 49138 36570
rect 49172 36536 49228 36570
rect 49262 36536 49318 36570
rect 49352 36536 49408 36570
rect 49442 36536 49494 36570
rect 48814 36480 49494 36536
rect 48814 36446 48868 36480
rect 48902 36446 48958 36480
rect 48992 36446 49048 36480
rect 49082 36446 49138 36480
rect 49172 36446 49228 36480
rect 49262 36446 49318 36480
rect 49352 36446 49408 36480
rect 49442 36446 49494 36480
rect 48814 36392 49494 36446
rect 50154 37020 50834 37072
rect 50154 36986 50208 37020
rect 50242 36986 50298 37020
rect 50332 36986 50388 37020
rect 50422 36986 50478 37020
rect 50512 36986 50568 37020
rect 50602 36986 50658 37020
rect 50692 36986 50748 37020
rect 50782 36986 50834 37020
rect 50154 36930 50834 36986
rect 50154 36896 50208 36930
rect 50242 36896 50298 36930
rect 50332 36896 50388 36930
rect 50422 36896 50478 36930
rect 50512 36896 50568 36930
rect 50602 36896 50658 36930
rect 50692 36896 50748 36930
rect 50782 36896 50834 36930
rect 50154 36840 50834 36896
rect 50154 36806 50208 36840
rect 50242 36806 50298 36840
rect 50332 36806 50388 36840
rect 50422 36806 50478 36840
rect 50512 36806 50568 36840
rect 50602 36806 50658 36840
rect 50692 36806 50748 36840
rect 50782 36806 50834 36840
rect 50154 36750 50834 36806
rect 50154 36716 50208 36750
rect 50242 36716 50298 36750
rect 50332 36716 50388 36750
rect 50422 36716 50478 36750
rect 50512 36716 50568 36750
rect 50602 36716 50658 36750
rect 50692 36716 50748 36750
rect 50782 36716 50834 36750
rect 50154 36660 50834 36716
rect 50154 36626 50208 36660
rect 50242 36626 50298 36660
rect 50332 36626 50388 36660
rect 50422 36626 50478 36660
rect 50512 36626 50568 36660
rect 50602 36626 50658 36660
rect 50692 36626 50748 36660
rect 50782 36626 50834 36660
rect 50154 36570 50834 36626
rect 50154 36536 50208 36570
rect 50242 36536 50298 36570
rect 50332 36536 50388 36570
rect 50422 36536 50478 36570
rect 50512 36536 50568 36570
rect 50602 36536 50658 36570
rect 50692 36536 50748 36570
rect 50782 36536 50834 36570
rect 50154 36480 50834 36536
rect 50154 36446 50208 36480
rect 50242 36446 50298 36480
rect 50332 36446 50388 36480
rect 50422 36446 50478 36480
rect 50512 36446 50568 36480
rect 50602 36446 50658 36480
rect 50692 36446 50748 36480
rect 50782 36446 50834 36480
rect 50154 36392 50834 36446
rect 51494 37020 52174 37072
rect 51494 36986 51548 37020
rect 51582 36986 51638 37020
rect 51672 36986 51728 37020
rect 51762 36986 51818 37020
rect 51852 36986 51908 37020
rect 51942 36986 51998 37020
rect 52032 36986 52088 37020
rect 52122 36986 52174 37020
rect 51494 36930 52174 36986
rect 51494 36896 51548 36930
rect 51582 36896 51638 36930
rect 51672 36896 51728 36930
rect 51762 36896 51818 36930
rect 51852 36896 51908 36930
rect 51942 36896 51998 36930
rect 52032 36896 52088 36930
rect 52122 36896 52174 36930
rect 51494 36840 52174 36896
rect 51494 36806 51548 36840
rect 51582 36806 51638 36840
rect 51672 36806 51728 36840
rect 51762 36806 51818 36840
rect 51852 36806 51908 36840
rect 51942 36806 51998 36840
rect 52032 36806 52088 36840
rect 52122 36806 52174 36840
rect 51494 36750 52174 36806
rect 51494 36716 51548 36750
rect 51582 36716 51638 36750
rect 51672 36716 51728 36750
rect 51762 36716 51818 36750
rect 51852 36716 51908 36750
rect 51942 36716 51998 36750
rect 52032 36716 52088 36750
rect 52122 36716 52174 36750
rect 51494 36660 52174 36716
rect 51494 36626 51548 36660
rect 51582 36626 51638 36660
rect 51672 36626 51728 36660
rect 51762 36626 51818 36660
rect 51852 36626 51908 36660
rect 51942 36626 51998 36660
rect 52032 36626 52088 36660
rect 52122 36626 52174 36660
rect 51494 36570 52174 36626
rect 51494 36536 51548 36570
rect 51582 36536 51638 36570
rect 51672 36536 51728 36570
rect 51762 36536 51818 36570
rect 51852 36536 51908 36570
rect 51942 36536 51998 36570
rect 52032 36536 52088 36570
rect 52122 36536 52174 36570
rect 51494 36480 52174 36536
rect 51494 36446 51548 36480
rect 51582 36446 51638 36480
rect 51672 36446 51728 36480
rect 51762 36446 51818 36480
rect 51852 36446 51908 36480
rect 51942 36446 51998 36480
rect 52032 36446 52088 36480
rect 52122 36446 52174 36480
rect 51494 36392 52174 36446
rect 42114 33260 42794 33312
rect 42114 33226 42168 33260
rect 42202 33226 42258 33260
rect 42292 33226 42348 33260
rect 42382 33226 42438 33260
rect 42472 33226 42528 33260
rect 42562 33226 42618 33260
rect 42652 33226 42708 33260
rect 42742 33226 42794 33260
rect 42114 33170 42794 33226
rect 42114 33136 42168 33170
rect 42202 33136 42258 33170
rect 42292 33136 42348 33170
rect 42382 33136 42438 33170
rect 42472 33136 42528 33170
rect 42562 33136 42618 33170
rect 42652 33136 42708 33170
rect 42742 33136 42794 33170
rect 42114 33080 42794 33136
rect 42114 33046 42168 33080
rect 42202 33046 42258 33080
rect 42292 33046 42348 33080
rect 42382 33046 42438 33080
rect 42472 33046 42528 33080
rect 42562 33046 42618 33080
rect 42652 33046 42708 33080
rect 42742 33046 42794 33080
rect 42114 32990 42794 33046
rect 42114 32956 42168 32990
rect 42202 32956 42258 32990
rect 42292 32956 42348 32990
rect 42382 32956 42438 32990
rect 42472 32956 42528 32990
rect 42562 32956 42618 32990
rect 42652 32956 42708 32990
rect 42742 32956 42794 32990
rect 42114 32900 42794 32956
rect 42114 32866 42168 32900
rect 42202 32866 42258 32900
rect 42292 32866 42348 32900
rect 42382 32866 42438 32900
rect 42472 32866 42528 32900
rect 42562 32866 42618 32900
rect 42652 32866 42708 32900
rect 42742 32866 42794 32900
rect 42114 32810 42794 32866
rect 42114 32776 42168 32810
rect 42202 32776 42258 32810
rect 42292 32776 42348 32810
rect 42382 32776 42438 32810
rect 42472 32776 42528 32810
rect 42562 32776 42618 32810
rect 42652 32776 42708 32810
rect 42742 32776 42794 32810
rect 42114 32720 42794 32776
rect 42114 32686 42168 32720
rect 42202 32686 42258 32720
rect 42292 32686 42348 32720
rect 42382 32686 42438 32720
rect 42472 32686 42528 32720
rect 42562 32686 42618 32720
rect 42652 32686 42708 32720
rect 42742 32686 42794 32720
rect 42114 32632 42794 32686
rect 43454 33260 44134 33312
rect 43454 33226 43508 33260
rect 43542 33226 43598 33260
rect 43632 33226 43688 33260
rect 43722 33226 43778 33260
rect 43812 33226 43868 33260
rect 43902 33226 43958 33260
rect 43992 33226 44048 33260
rect 44082 33226 44134 33260
rect 43454 33170 44134 33226
rect 43454 33136 43508 33170
rect 43542 33136 43598 33170
rect 43632 33136 43688 33170
rect 43722 33136 43778 33170
rect 43812 33136 43868 33170
rect 43902 33136 43958 33170
rect 43992 33136 44048 33170
rect 44082 33136 44134 33170
rect 43454 33080 44134 33136
rect 43454 33046 43508 33080
rect 43542 33046 43598 33080
rect 43632 33046 43688 33080
rect 43722 33046 43778 33080
rect 43812 33046 43868 33080
rect 43902 33046 43958 33080
rect 43992 33046 44048 33080
rect 44082 33046 44134 33080
rect 43454 32990 44134 33046
rect 43454 32956 43508 32990
rect 43542 32956 43598 32990
rect 43632 32956 43688 32990
rect 43722 32956 43778 32990
rect 43812 32956 43868 32990
rect 43902 32956 43958 32990
rect 43992 32956 44048 32990
rect 44082 32956 44134 32990
rect 43454 32900 44134 32956
rect 43454 32866 43508 32900
rect 43542 32866 43598 32900
rect 43632 32866 43688 32900
rect 43722 32866 43778 32900
rect 43812 32866 43868 32900
rect 43902 32866 43958 32900
rect 43992 32866 44048 32900
rect 44082 32866 44134 32900
rect 43454 32810 44134 32866
rect 43454 32776 43508 32810
rect 43542 32776 43598 32810
rect 43632 32776 43688 32810
rect 43722 32776 43778 32810
rect 43812 32776 43868 32810
rect 43902 32776 43958 32810
rect 43992 32776 44048 32810
rect 44082 32776 44134 32810
rect 43454 32720 44134 32776
rect 43454 32686 43508 32720
rect 43542 32686 43598 32720
rect 43632 32686 43688 32720
rect 43722 32686 43778 32720
rect 43812 32686 43868 32720
rect 43902 32686 43958 32720
rect 43992 32686 44048 32720
rect 44082 32686 44134 32720
rect 43454 32632 44134 32686
rect 44794 33260 45474 33312
rect 44794 33226 44848 33260
rect 44882 33226 44938 33260
rect 44972 33226 45028 33260
rect 45062 33226 45118 33260
rect 45152 33226 45208 33260
rect 45242 33226 45298 33260
rect 45332 33226 45388 33260
rect 45422 33226 45474 33260
rect 44794 33170 45474 33226
rect 44794 33136 44848 33170
rect 44882 33136 44938 33170
rect 44972 33136 45028 33170
rect 45062 33136 45118 33170
rect 45152 33136 45208 33170
rect 45242 33136 45298 33170
rect 45332 33136 45388 33170
rect 45422 33136 45474 33170
rect 44794 33080 45474 33136
rect 44794 33046 44848 33080
rect 44882 33046 44938 33080
rect 44972 33046 45028 33080
rect 45062 33046 45118 33080
rect 45152 33046 45208 33080
rect 45242 33046 45298 33080
rect 45332 33046 45388 33080
rect 45422 33046 45474 33080
rect 44794 32990 45474 33046
rect 44794 32956 44848 32990
rect 44882 32956 44938 32990
rect 44972 32956 45028 32990
rect 45062 32956 45118 32990
rect 45152 32956 45208 32990
rect 45242 32956 45298 32990
rect 45332 32956 45388 32990
rect 45422 32956 45474 32990
rect 44794 32900 45474 32956
rect 44794 32866 44848 32900
rect 44882 32866 44938 32900
rect 44972 32866 45028 32900
rect 45062 32866 45118 32900
rect 45152 32866 45208 32900
rect 45242 32866 45298 32900
rect 45332 32866 45388 32900
rect 45422 32866 45474 32900
rect 44794 32810 45474 32866
rect 44794 32776 44848 32810
rect 44882 32776 44938 32810
rect 44972 32776 45028 32810
rect 45062 32776 45118 32810
rect 45152 32776 45208 32810
rect 45242 32776 45298 32810
rect 45332 32776 45388 32810
rect 45422 32776 45474 32810
rect 44794 32720 45474 32776
rect 44794 32686 44848 32720
rect 44882 32686 44938 32720
rect 44972 32686 45028 32720
rect 45062 32686 45118 32720
rect 45152 32686 45208 32720
rect 45242 32686 45298 32720
rect 45332 32686 45388 32720
rect 45422 32686 45474 32720
rect 44794 32632 45474 32686
rect 46134 33260 46814 33312
rect 46134 33226 46188 33260
rect 46222 33226 46278 33260
rect 46312 33226 46368 33260
rect 46402 33226 46458 33260
rect 46492 33226 46548 33260
rect 46582 33226 46638 33260
rect 46672 33226 46728 33260
rect 46762 33226 46814 33260
rect 46134 33170 46814 33226
rect 46134 33136 46188 33170
rect 46222 33136 46278 33170
rect 46312 33136 46368 33170
rect 46402 33136 46458 33170
rect 46492 33136 46548 33170
rect 46582 33136 46638 33170
rect 46672 33136 46728 33170
rect 46762 33136 46814 33170
rect 46134 33080 46814 33136
rect 46134 33046 46188 33080
rect 46222 33046 46278 33080
rect 46312 33046 46368 33080
rect 46402 33046 46458 33080
rect 46492 33046 46548 33080
rect 46582 33046 46638 33080
rect 46672 33046 46728 33080
rect 46762 33046 46814 33080
rect 46134 32990 46814 33046
rect 46134 32956 46188 32990
rect 46222 32956 46278 32990
rect 46312 32956 46368 32990
rect 46402 32956 46458 32990
rect 46492 32956 46548 32990
rect 46582 32956 46638 32990
rect 46672 32956 46728 32990
rect 46762 32956 46814 32990
rect 46134 32900 46814 32956
rect 46134 32866 46188 32900
rect 46222 32866 46278 32900
rect 46312 32866 46368 32900
rect 46402 32866 46458 32900
rect 46492 32866 46548 32900
rect 46582 32866 46638 32900
rect 46672 32866 46728 32900
rect 46762 32866 46814 32900
rect 46134 32810 46814 32866
rect 46134 32776 46188 32810
rect 46222 32776 46278 32810
rect 46312 32776 46368 32810
rect 46402 32776 46458 32810
rect 46492 32776 46548 32810
rect 46582 32776 46638 32810
rect 46672 32776 46728 32810
rect 46762 32776 46814 32810
rect 46134 32720 46814 32776
rect 46134 32686 46188 32720
rect 46222 32686 46278 32720
rect 46312 32686 46368 32720
rect 46402 32686 46458 32720
rect 46492 32686 46548 32720
rect 46582 32686 46638 32720
rect 46672 32686 46728 32720
rect 46762 32686 46814 32720
rect 46134 32632 46814 32686
rect 47474 33260 48154 33312
rect 47474 33226 47528 33260
rect 47562 33226 47618 33260
rect 47652 33226 47708 33260
rect 47742 33226 47798 33260
rect 47832 33226 47888 33260
rect 47922 33226 47978 33260
rect 48012 33226 48068 33260
rect 48102 33226 48154 33260
rect 47474 33170 48154 33226
rect 47474 33136 47528 33170
rect 47562 33136 47618 33170
rect 47652 33136 47708 33170
rect 47742 33136 47798 33170
rect 47832 33136 47888 33170
rect 47922 33136 47978 33170
rect 48012 33136 48068 33170
rect 48102 33136 48154 33170
rect 47474 33080 48154 33136
rect 47474 33046 47528 33080
rect 47562 33046 47618 33080
rect 47652 33046 47708 33080
rect 47742 33046 47798 33080
rect 47832 33046 47888 33080
rect 47922 33046 47978 33080
rect 48012 33046 48068 33080
rect 48102 33046 48154 33080
rect 47474 32990 48154 33046
rect 47474 32956 47528 32990
rect 47562 32956 47618 32990
rect 47652 32956 47708 32990
rect 47742 32956 47798 32990
rect 47832 32956 47888 32990
rect 47922 32956 47978 32990
rect 48012 32956 48068 32990
rect 48102 32956 48154 32990
rect 47474 32900 48154 32956
rect 47474 32866 47528 32900
rect 47562 32866 47618 32900
rect 47652 32866 47708 32900
rect 47742 32866 47798 32900
rect 47832 32866 47888 32900
rect 47922 32866 47978 32900
rect 48012 32866 48068 32900
rect 48102 32866 48154 32900
rect 47474 32810 48154 32866
rect 47474 32776 47528 32810
rect 47562 32776 47618 32810
rect 47652 32776 47708 32810
rect 47742 32776 47798 32810
rect 47832 32776 47888 32810
rect 47922 32776 47978 32810
rect 48012 32776 48068 32810
rect 48102 32776 48154 32810
rect 47474 32720 48154 32776
rect 47474 32686 47528 32720
rect 47562 32686 47618 32720
rect 47652 32686 47708 32720
rect 47742 32686 47798 32720
rect 47832 32686 47888 32720
rect 47922 32686 47978 32720
rect 48012 32686 48068 32720
rect 48102 32686 48154 32720
rect 47474 32632 48154 32686
rect 48814 33260 49494 33312
rect 48814 33226 48868 33260
rect 48902 33226 48958 33260
rect 48992 33226 49048 33260
rect 49082 33226 49138 33260
rect 49172 33226 49228 33260
rect 49262 33226 49318 33260
rect 49352 33226 49408 33260
rect 49442 33226 49494 33260
rect 48814 33170 49494 33226
rect 48814 33136 48868 33170
rect 48902 33136 48958 33170
rect 48992 33136 49048 33170
rect 49082 33136 49138 33170
rect 49172 33136 49228 33170
rect 49262 33136 49318 33170
rect 49352 33136 49408 33170
rect 49442 33136 49494 33170
rect 48814 33080 49494 33136
rect 48814 33046 48868 33080
rect 48902 33046 48958 33080
rect 48992 33046 49048 33080
rect 49082 33046 49138 33080
rect 49172 33046 49228 33080
rect 49262 33046 49318 33080
rect 49352 33046 49408 33080
rect 49442 33046 49494 33080
rect 48814 32990 49494 33046
rect 48814 32956 48868 32990
rect 48902 32956 48958 32990
rect 48992 32956 49048 32990
rect 49082 32956 49138 32990
rect 49172 32956 49228 32990
rect 49262 32956 49318 32990
rect 49352 32956 49408 32990
rect 49442 32956 49494 32990
rect 48814 32900 49494 32956
rect 48814 32866 48868 32900
rect 48902 32866 48958 32900
rect 48992 32866 49048 32900
rect 49082 32866 49138 32900
rect 49172 32866 49228 32900
rect 49262 32866 49318 32900
rect 49352 32866 49408 32900
rect 49442 32866 49494 32900
rect 48814 32810 49494 32866
rect 48814 32776 48868 32810
rect 48902 32776 48958 32810
rect 48992 32776 49048 32810
rect 49082 32776 49138 32810
rect 49172 32776 49228 32810
rect 49262 32776 49318 32810
rect 49352 32776 49408 32810
rect 49442 32776 49494 32810
rect 48814 32720 49494 32776
rect 48814 32686 48868 32720
rect 48902 32686 48958 32720
rect 48992 32686 49048 32720
rect 49082 32686 49138 32720
rect 49172 32686 49228 32720
rect 49262 32686 49318 32720
rect 49352 32686 49408 32720
rect 49442 32686 49494 32720
rect 48814 32632 49494 32686
rect 50154 33260 50834 33312
rect 50154 33226 50208 33260
rect 50242 33226 50298 33260
rect 50332 33226 50388 33260
rect 50422 33226 50478 33260
rect 50512 33226 50568 33260
rect 50602 33226 50658 33260
rect 50692 33226 50748 33260
rect 50782 33226 50834 33260
rect 50154 33170 50834 33226
rect 50154 33136 50208 33170
rect 50242 33136 50298 33170
rect 50332 33136 50388 33170
rect 50422 33136 50478 33170
rect 50512 33136 50568 33170
rect 50602 33136 50658 33170
rect 50692 33136 50748 33170
rect 50782 33136 50834 33170
rect 50154 33080 50834 33136
rect 50154 33046 50208 33080
rect 50242 33046 50298 33080
rect 50332 33046 50388 33080
rect 50422 33046 50478 33080
rect 50512 33046 50568 33080
rect 50602 33046 50658 33080
rect 50692 33046 50748 33080
rect 50782 33046 50834 33080
rect 50154 32990 50834 33046
rect 50154 32956 50208 32990
rect 50242 32956 50298 32990
rect 50332 32956 50388 32990
rect 50422 32956 50478 32990
rect 50512 32956 50568 32990
rect 50602 32956 50658 32990
rect 50692 32956 50748 32990
rect 50782 32956 50834 32990
rect 50154 32900 50834 32956
rect 50154 32866 50208 32900
rect 50242 32866 50298 32900
rect 50332 32866 50388 32900
rect 50422 32866 50478 32900
rect 50512 32866 50568 32900
rect 50602 32866 50658 32900
rect 50692 32866 50748 32900
rect 50782 32866 50834 32900
rect 50154 32810 50834 32866
rect 50154 32776 50208 32810
rect 50242 32776 50298 32810
rect 50332 32776 50388 32810
rect 50422 32776 50478 32810
rect 50512 32776 50568 32810
rect 50602 32776 50658 32810
rect 50692 32776 50748 32810
rect 50782 32776 50834 32810
rect 50154 32720 50834 32776
rect 50154 32686 50208 32720
rect 50242 32686 50298 32720
rect 50332 32686 50388 32720
rect 50422 32686 50478 32720
rect 50512 32686 50568 32720
rect 50602 32686 50658 32720
rect 50692 32686 50748 32720
rect 50782 32686 50834 32720
rect 50154 32632 50834 32686
rect 51494 33260 52174 33312
rect 51494 33226 51548 33260
rect 51582 33226 51638 33260
rect 51672 33226 51728 33260
rect 51762 33226 51818 33260
rect 51852 33226 51908 33260
rect 51942 33226 51998 33260
rect 52032 33226 52088 33260
rect 52122 33226 52174 33260
rect 51494 33170 52174 33226
rect 51494 33136 51548 33170
rect 51582 33136 51638 33170
rect 51672 33136 51728 33170
rect 51762 33136 51818 33170
rect 51852 33136 51908 33170
rect 51942 33136 51998 33170
rect 52032 33136 52088 33170
rect 52122 33136 52174 33170
rect 51494 33080 52174 33136
rect 51494 33046 51548 33080
rect 51582 33046 51638 33080
rect 51672 33046 51728 33080
rect 51762 33046 51818 33080
rect 51852 33046 51908 33080
rect 51942 33046 51998 33080
rect 52032 33046 52088 33080
rect 52122 33046 52174 33080
rect 51494 32990 52174 33046
rect 51494 32956 51548 32990
rect 51582 32956 51638 32990
rect 51672 32956 51728 32990
rect 51762 32956 51818 32990
rect 51852 32956 51908 32990
rect 51942 32956 51998 32990
rect 52032 32956 52088 32990
rect 52122 32956 52174 32990
rect 51494 32900 52174 32956
rect 51494 32866 51548 32900
rect 51582 32866 51638 32900
rect 51672 32866 51728 32900
rect 51762 32866 51818 32900
rect 51852 32866 51908 32900
rect 51942 32866 51998 32900
rect 52032 32866 52088 32900
rect 52122 32866 52174 32900
rect 51494 32810 52174 32866
rect 51494 32776 51548 32810
rect 51582 32776 51638 32810
rect 51672 32776 51728 32810
rect 51762 32776 51818 32810
rect 51852 32776 51908 32810
rect 51942 32776 51998 32810
rect 52032 32776 52088 32810
rect 52122 32776 52174 32810
rect 51494 32720 52174 32776
rect 51494 32686 51548 32720
rect 51582 32686 51638 32720
rect 51672 32686 51728 32720
rect 51762 32686 51818 32720
rect 51852 32686 51908 32720
rect 51942 32686 51998 32720
rect 52032 32686 52088 32720
rect 52122 32686 52174 32720
rect 51494 32632 52174 32686
rect 37507 29901 37565 29917
rect 37507 29867 37519 29901
rect 37553 29867 37565 29901
rect 37507 29833 37565 29867
rect 37507 29799 37519 29833
rect 37553 29799 37565 29833
rect 37507 29765 37565 29799
rect 37507 29731 37519 29765
rect 37553 29731 37565 29765
rect 37507 29697 37565 29731
rect 37507 29663 37519 29697
rect 37553 29663 37565 29697
rect 37507 29629 37565 29663
rect 37507 29595 37519 29629
rect 37553 29595 37565 29629
rect 37507 29561 37565 29595
rect 37507 29527 37519 29561
rect 37553 29527 37565 29561
rect 37507 29493 37565 29527
rect 37507 29459 37519 29493
rect 37553 29459 37565 29493
rect 37507 29425 37565 29459
rect 37507 29391 37519 29425
rect 37553 29391 37565 29425
rect 37507 29357 37565 29391
rect 37507 29323 37519 29357
rect 37553 29323 37565 29357
rect 37507 29289 37565 29323
rect 37507 29255 37519 29289
rect 37553 29255 37565 29289
rect 37507 29221 37565 29255
rect 37507 29187 37519 29221
rect 37553 29187 37565 29221
rect 37507 29153 37565 29187
rect 37507 29119 37519 29153
rect 37553 29119 37565 29153
rect 37507 29085 37565 29119
rect 37507 29051 37519 29085
rect 37553 29051 37565 29085
rect 37507 29017 37565 29051
rect 37507 28983 37519 29017
rect 37553 28983 37565 29017
rect 37507 28949 37565 28983
rect 37507 28915 37519 28949
rect 37553 28915 37565 28949
rect 37507 28881 37565 28915
rect 37507 28847 37519 28881
rect 37553 28847 37565 28881
rect 37507 28813 37565 28847
rect 37507 28779 37519 28813
rect 37553 28779 37565 28813
rect 37507 28745 37565 28779
rect 37507 28711 37519 28745
rect 37553 28711 37565 28745
rect 37507 28677 37565 28711
rect 37507 28643 37519 28677
rect 37553 28643 37565 28677
rect 37507 28627 37565 28643
rect 37965 29901 38023 29917
rect 37965 29867 37977 29901
rect 38011 29867 38023 29901
rect 37965 29833 38023 29867
rect 37965 29799 37977 29833
rect 38011 29799 38023 29833
rect 37965 29765 38023 29799
rect 37965 29731 37977 29765
rect 38011 29731 38023 29765
rect 37965 29697 38023 29731
rect 37965 29663 37977 29697
rect 38011 29663 38023 29697
rect 37965 29629 38023 29663
rect 37965 29595 37977 29629
rect 38011 29595 38023 29629
rect 37965 29561 38023 29595
rect 37965 29527 37977 29561
rect 38011 29527 38023 29561
rect 37965 29493 38023 29527
rect 37965 29459 37977 29493
rect 38011 29459 38023 29493
rect 37965 29425 38023 29459
rect 37965 29391 37977 29425
rect 38011 29391 38023 29425
rect 37965 29357 38023 29391
rect 37965 29323 37977 29357
rect 38011 29323 38023 29357
rect 37965 29289 38023 29323
rect 37965 29255 37977 29289
rect 38011 29255 38023 29289
rect 37965 29221 38023 29255
rect 37965 29187 37977 29221
rect 38011 29187 38023 29221
rect 37965 29153 38023 29187
rect 37965 29119 37977 29153
rect 38011 29119 38023 29153
rect 37965 29085 38023 29119
rect 37965 29051 37977 29085
rect 38011 29051 38023 29085
rect 37965 29017 38023 29051
rect 37965 28983 37977 29017
rect 38011 28983 38023 29017
rect 37965 28949 38023 28983
rect 37965 28915 37977 28949
rect 38011 28915 38023 28949
rect 37965 28881 38023 28915
rect 37965 28847 37977 28881
rect 38011 28847 38023 28881
rect 37965 28813 38023 28847
rect 37965 28779 37977 28813
rect 38011 28779 38023 28813
rect 37965 28745 38023 28779
rect 37965 28711 37977 28745
rect 38011 28711 38023 28745
rect 37965 28677 38023 28711
rect 37965 28643 37977 28677
rect 38011 28643 38023 28677
rect 37965 28627 38023 28643
rect 38423 29901 38481 29917
rect 38423 29867 38435 29901
rect 38469 29867 38481 29901
rect 38423 29833 38481 29867
rect 38423 29799 38435 29833
rect 38469 29799 38481 29833
rect 38423 29765 38481 29799
rect 38423 29731 38435 29765
rect 38469 29731 38481 29765
rect 38423 29697 38481 29731
rect 38423 29663 38435 29697
rect 38469 29663 38481 29697
rect 38423 29629 38481 29663
rect 38423 29595 38435 29629
rect 38469 29595 38481 29629
rect 38423 29561 38481 29595
rect 38423 29527 38435 29561
rect 38469 29527 38481 29561
rect 38423 29493 38481 29527
rect 38423 29459 38435 29493
rect 38469 29459 38481 29493
rect 38423 29425 38481 29459
rect 38423 29391 38435 29425
rect 38469 29391 38481 29425
rect 38423 29357 38481 29391
rect 38423 29323 38435 29357
rect 38469 29323 38481 29357
rect 38423 29289 38481 29323
rect 38423 29255 38435 29289
rect 38469 29255 38481 29289
rect 38423 29221 38481 29255
rect 38423 29187 38435 29221
rect 38469 29187 38481 29221
rect 38423 29153 38481 29187
rect 38423 29119 38435 29153
rect 38469 29119 38481 29153
rect 38423 29085 38481 29119
rect 38423 29051 38435 29085
rect 38469 29051 38481 29085
rect 38423 29017 38481 29051
rect 38423 28983 38435 29017
rect 38469 28983 38481 29017
rect 38423 28949 38481 28983
rect 38423 28915 38435 28949
rect 38469 28915 38481 28949
rect 38423 28881 38481 28915
rect 38423 28847 38435 28881
rect 38469 28847 38481 28881
rect 38423 28813 38481 28847
rect 38423 28779 38435 28813
rect 38469 28779 38481 28813
rect 38423 28745 38481 28779
rect 38423 28711 38435 28745
rect 38469 28711 38481 28745
rect 38423 28677 38481 28711
rect 38423 28643 38435 28677
rect 38469 28643 38481 28677
rect 38423 28627 38481 28643
rect 38881 29901 38939 29917
rect 38881 29867 38893 29901
rect 38927 29867 38939 29901
rect 38881 29833 38939 29867
rect 38881 29799 38893 29833
rect 38927 29799 38939 29833
rect 38881 29765 38939 29799
rect 38881 29731 38893 29765
rect 38927 29731 38939 29765
rect 38881 29697 38939 29731
rect 38881 29663 38893 29697
rect 38927 29663 38939 29697
rect 38881 29629 38939 29663
rect 38881 29595 38893 29629
rect 38927 29595 38939 29629
rect 38881 29561 38939 29595
rect 38881 29527 38893 29561
rect 38927 29527 38939 29561
rect 38881 29493 38939 29527
rect 38881 29459 38893 29493
rect 38927 29459 38939 29493
rect 38881 29425 38939 29459
rect 38881 29391 38893 29425
rect 38927 29391 38939 29425
rect 38881 29357 38939 29391
rect 38881 29323 38893 29357
rect 38927 29323 38939 29357
rect 38881 29289 38939 29323
rect 38881 29255 38893 29289
rect 38927 29255 38939 29289
rect 38881 29221 38939 29255
rect 38881 29187 38893 29221
rect 38927 29187 38939 29221
rect 38881 29153 38939 29187
rect 38881 29119 38893 29153
rect 38927 29119 38939 29153
rect 38881 29085 38939 29119
rect 38881 29051 38893 29085
rect 38927 29051 38939 29085
rect 38881 29017 38939 29051
rect 38881 28983 38893 29017
rect 38927 28983 38939 29017
rect 38881 28949 38939 28983
rect 38881 28915 38893 28949
rect 38927 28915 38939 28949
rect 38881 28881 38939 28915
rect 38881 28847 38893 28881
rect 38927 28847 38939 28881
rect 38881 28813 38939 28847
rect 38881 28779 38893 28813
rect 38927 28779 38939 28813
rect 38881 28745 38939 28779
rect 38881 28711 38893 28745
rect 38927 28711 38939 28745
rect 38881 28677 38939 28711
rect 38881 28643 38893 28677
rect 38927 28643 38939 28677
rect 38881 28627 38939 28643
rect 39339 29901 39397 29917
rect 39339 29867 39351 29901
rect 39385 29867 39397 29901
rect 39339 29833 39397 29867
rect 39339 29799 39351 29833
rect 39385 29799 39397 29833
rect 39339 29765 39397 29799
rect 39339 29731 39351 29765
rect 39385 29731 39397 29765
rect 39339 29697 39397 29731
rect 39339 29663 39351 29697
rect 39385 29663 39397 29697
rect 39339 29629 39397 29663
rect 39339 29595 39351 29629
rect 39385 29595 39397 29629
rect 39339 29561 39397 29595
rect 39339 29527 39351 29561
rect 39385 29527 39397 29561
rect 39339 29493 39397 29527
rect 39339 29459 39351 29493
rect 39385 29459 39397 29493
rect 39339 29425 39397 29459
rect 39339 29391 39351 29425
rect 39385 29391 39397 29425
rect 39339 29357 39397 29391
rect 39339 29323 39351 29357
rect 39385 29323 39397 29357
rect 39339 29289 39397 29323
rect 39339 29255 39351 29289
rect 39385 29255 39397 29289
rect 39339 29221 39397 29255
rect 39339 29187 39351 29221
rect 39385 29187 39397 29221
rect 39339 29153 39397 29187
rect 39339 29119 39351 29153
rect 39385 29119 39397 29153
rect 39339 29085 39397 29119
rect 39339 29051 39351 29085
rect 39385 29051 39397 29085
rect 39339 29017 39397 29051
rect 39339 28983 39351 29017
rect 39385 28983 39397 29017
rect 39339 28949 39397 28983
rect 39339 28915 39351 28949
rect 39385 28915 39397 28949
rect 39339 28881 39397 28915
rect 39339 28847 39351 28881
rect 39385 28847 39397 28881
rect 39339 28813 39397 28847
rect 39339 28779 39351 28813
rect 39385 28779 39397 28813
rect 39339 28745 39397 28779
rect 39339 28711 39351 28745
rect 39385 28711 39397 28745
rect 39339 28677 39397 28711
rect 39339 28643 39351 28677
rect 39385 28643 39397 28677
rect 39339 28627 39397 28643
rect 39797 29901 39855 29917
rect 39797 29867 39809 29901
rect 39843 29867 39855 29901
rect 39797 29833 39855 29867
rect 39797 29799 39809 29833
rect 39843 29799 39855 29833
rect 39797 29765 39855 29799
rect 39797 29731 39809 29765
rect 39843 29731 39855 29765
rect 39797 29697 39855 29731
rect 39797 29663 39809 29697
rect 39843 29663 39855 29697
rect 39797 29629 39855 29663
rect 39797 29595 39809 29629
rect 39843 29595 39855 29629
rect 39797 29561 39855 29595
rect 39797 29527 39809 29561
rect 39843 29527 39855 29561
rect 39797 29493 39855 29527
rect 39797 29459 39809 29493
rect 39843 29459 39855 29493
rect 39797 29425 39855 29459
rect 39797 29391 39809 29425
rect 39843 29391 39855 29425
rect 39797 29357 39855 29391
rect 39797 29323 39809 29357
rect 39843 29323 39855 29357
rect 39797 29289 39855 29323
rect 39797 29255 39809 29289
rect 39843 29255 39855 29289
rect 39797 29221 39855 29255
rect 39797 29187 39809 29221
rect 39843 29187 39855 29221
rect 39797 29153 39855 29187
rect 39797 29119 39809 29153
rect 39843 29119 39855 29153
rect 39797 29085 39855 29119
rect 39797 29051 39809 29085
rect 39843 29051 39855 29085
rect 39797 29017 39855 29051
rect 39797 28983 39809 29017
rect 39843 28983 39855 29017
rect 39797 28949 39855 28983
rect 39797 28915 39809 28949
rect 39843 28915 39855 28949
rect 39797 28881 39855 28915
rect 39797 28847 39809 28881
rect 39843 28847 39855 28881
rect 39797 28813 39855 28847
rect 39797 28779 39809 28813
rect 39843 28779 39855 28813
rect 39797 28745 39855 28779
rect 39797 28711 39809 28745
rect 39843 28711 39855 28745
rect 39797 28677 39855 28711
rect 39797 28643 39809 28677
rect 39843 28643 39855 28677
rect 39797 28627 39855 28643
rect 40255 29901 40313 29917
rect 40255 29867 40267 29901
rect 40301 29867 40313 29901
rect 40255 29833 40313 29867
rect 40255 29799 40267 29833
rect 40301 29799 40313 29833
rect 40255 29765 40313 29799
rect 40255 29731 40267 29765
rect 40301 29731 40313 29765
rect 40255 29697 40313 29731
rect 40255 29663 40267 29697
rect 40301 29663 40313 29697
rect 40255 29629 40313 29663
rect 40255 29595 40267 29629
rect 40301 29595 40313 29629
rect 40255 29561 40313 29595
rect 40255 29527 40267 29561
rect 40301 29527 40313 29561
rect 40255 29493 40313 29527
rect 40255 29459 40267 29493
rect 40301 29459 40313 29493
rect 40255 29425 40313 29459
rect 40255 29391 40267 29425
rect 40301 29391 40313 29425
rect 40255 29357 40313 29391
rect 40255 29323 40267 29357
rect 40301 29323 40313 29357
rect 40255 29289 40313 29323
rect 40255 29255 40267 29289
rect 40301 29255 40313 29289
rect 40255 29221 40313 29255
rect 40255 29187 40267 29221
rect 40301 29187 40313 29221
rect 40255 29153 40313 29187
rect 40255 29119 40267 29153
rect 40301 29119 40313 29153
rect 40255 29085 40313 29119
rect 40255 29051 40267 29085
rect 40301 29051 40313 29085
rect 40255 29017 40313 29051
rect 40255 28983 40267 29017
rect 40301 28983 40313 29017
rect 40255 28949 40313 28983
rect 40255 28915 40267 28949
rect 40301 28915 40313 28949
rect 40255 28881 40313 28915
rect 40255 28847 40267 28881
rect 40301 28847 40313 28881
rect 40255 28813 40313 28847
rect 40255 28779 40267 28813
rect 40301 28779 40313 28813
rect 40255 28745 40313 28779
rect 40255 28711 40267 28745
rect 40301 28711 40313 28745
rect 40255 28677 40313 28711
rect 40255 28643 40267 28677
rect 40301 28643 40313 28677
rect 40255 28627 40313 28643
rect 42114 29500 42794 29552
rect 42114 29466 42168 29500
rect 42202 29466 42258 29500
rect 42292 29466 42348 29500
rect 42382 29466 42438 29500
rect 42472 29466 42528 29500
rect 42562 29466 42618 29500
rect 42652 29466 42708 29500
rect 42742 29466 42794 29500
rect 42114 29410 42794 29466
rect 42114 29376 42168 29410
rect 42202 29376 42258 29410
rect 42292 29376 42348 29410
rect 42382 29376 42438 29410
rect 42472 29376 42528 29410
rect 42562 29376 42618 29410
rect 42652 29376 42708 29410
rect 42742 29376 42794 29410
rect 42114 29320 42794 29376
rect 42114 29286 42168 29320
rect 42202 29286 42258 29320
rect 42292 29286 42348 29320
rect 42382 29286 42438 29320
rect 42472 29286 42528 29320
rect 42562 29286 42618 29320
rect 42652 29286 42708 29320
rect 42742 29286 42794 29320
rect 42114 29230 42794 29286
rect 42114 29196 42168 29230
rect 42202 29196 42258 29230
rect 42292 29196 42348 29230
rect 42382 29196 42438 29230
rect 42472 29196 42528 29230
rect 42562 29196 42618 29230
rect 42652 29196 42708 29230
rect 42742 29196 42794 29230
rect 42114 29140 42794 29196
rect 42114 29106 42168 29140
rect 42202 29106 42258 29140
rect 42292 29106 42348 29140
rect 42382 29106 42438 29140
rect 42472 29106 42528 29140
rect 42562 29106 42618 29140
rect 42652 29106 42708 29140
rect 42742 29106 42794 29140
rect 42114 29050 42794 29106
rect 42114 29016 42168 29050
rect 42202 29016 42258 29050
rect 42292 29016 42348 29050
rect 42382 29016 42438 29050
rect 42472 29016 42528 29050
rect 42562 29016 42618 29050
rect 42652 29016 42708 29050
rect 42742 29016 42794 29050
rect 42114 28960 42794 29016
rect 42114 28926 42168 28960
rect 42202 28926 42258 28960
rect 42292 28926 42348 28960
rect 42382 28926 42438 28960
rect 42472 28926 42528 28960
rect 42562 28926 42618 28960
rect 42652 28926 42708 28960
rect 42742 28926 42794 28960
rect 42114 28872 42794 28926
rect 43454 29500 44134 29552
rect 43454 29466 43508 29500
rect 43542 29466 43598 29500
rect 43632 29466 43688 29500
rect 43722 29466 43778 29500
rect 43812 29466 43868 29500
rect 43902 29466 43958 29500
rect 43992 29466 44048 29500
rect 44082 29466 44134 29500
rect 43454 29410 44134 29466
rect 43454 29376 43508 29410
rect 43542 29376 43598 29410
rect 43632 29376 43688 29410
rect 43722 29376 43778 29410
rect 43812 29376 43868 29410
rect 43902 29376 43958 29410
rect 43992 29376 44048 29410
rect 44082 29376 44134 29410
rect 43454 29320 44134 29376
rect 43454 29286 43508 29320
rect 43542 29286 43598 29320
rect 43632 29286 43688 29320
rect 43722 29286 43778 29320
rect 43812 29286 43868 29320
rect 43902 29286 43958 29320
rect 43992 29286 44048 29320
rect 44082 29286 44134 29320
rect 43454 29230 44134 29286
rect 43454 29196 43508 29230
rect 43542 29196 43598 29230
rect 43632 29196 43688 29230
rect 43722 29196 43778 29230
rect 43812 29196 43868 29230
rect 43902 29196 43958 29230
rect 43992 29196 44048 29230
rect 44082 29196 44134 29230
rect 43454 29140 44134 29196
rect 43454 29106 43508 29140
rect 43542 29106 43598 29140
rect 43632 29106 43688 29140
rect 43722 29106 43778 29140
rect 43812 29106 43868 29140
rect 43902 29106 43958 29140
rect 43992 29106 44048 29140
rect 44082 29106 44134 29140
rect 43454 29050 44134 29106
rect 43454 29016 43508 29050
rect 43542 29016 43598 29050
rect 43632 29016 43688 29050
rect 43722 29016 43778 29050
rect 43812 29016 43868 29050
rect 43902 29016 43958 29050
rect 43992 29016 44048 29050
rect 44082 29016 44134 29050
rect 43454 28960 44134 29016
rect 43454 28926 43508 28960
rect 43542 28926 43598 28960
rect 43632 28926 43688 28960
rect 43722 28926 43778 28960
rect 43812 28926 43868 28960
rect 43902 28926 43958 28960
rect 43992 28926 44048 28960
rect 44082 28926 44134 28960
rect 43454 28872 44134 28926
rect 44794 29500 45474 29552
rect 44794 29466 44848 29500
rect 44882 29466 44938 29500
rect 44972 29466 45028 29500
rect 45062 29466 45118 29500
rect 45152 29466 45208 29500
rect 45242 29466 45298 29500
rect 45332 29466 45388 29500
rect 45422 29466 45474 29500
rect 44794 29410 45474 29466
rect 44794 29376 44848 29410
rect 44882 29376 44938 29410
rect 44972 29376 45028 29410
rect 45062 29376 45118 29410
rect 45152 29376 45208 29410
rect 45242 29376 45298 29410
rect 45332 29376 45388 29410
rect 45422 29376 45474 29410
rect 44794 29320 45474 29376
rect 44794 29286 44848 29320
rect 44882 29286 44938 29320
rect 44972 29286 45028 29320
rect 45062 29286 45118 29320
rect 45152 29286 45208 29320
rect 45242 29286 45298 29320
rect 45332 29286 45388 29320
rect 45422 29286 45474 29320
rect 44794 29230 45474 29286
rect 44794 29196 44848 29230
rect 44882 29196 44938 29230
rect 44972 29196 45028 29230
rect 45062 29196 45118 29230
rect 45152 29196 45208 29230
rect 45242 29196 45298 29230
rect 45332 29196 45388 29230
rect 45422 29196 45474 29230
rect 44794 29140 45474 29196
rect 44794 29106 44848 29140
rect 44882 29106 44938 29140
rect 44972 29106 45028 29140
rect 45062 29106 45118 29140
rect 45152 29106 45208 29140
rect 45242 29106 45298 29140
rect 45332 29106 45388 29140
rect 45422 29106 45474 29140
rect 44794 29050 45474 29106
rect 44794 29016 44848 29050
rect 44882 29016 44938 29050
rect 44972 29016 45028 29050
rect 45062 29016 45118 29050
rect 45152 29016 45208 29050
rect 45242 29016 45298 29050
rect 45332 29016 45388 29050
rect 45422 29016 45474 29050
rect 44794 28960 45474 29016
rect 44794 28926 44848 28960
rect 44882 28926 44938 28960
rect 44972 28926 45028 28960
rect 45062 28926 45118 28960
rect 45152 28926 45208 28960
rect 45242 28926 45298 28960
rect 45332 28926 45388 28960
rect 45422 28926 45474 28960
rect 44794 28872 45474 28926
rect 46134 29500 46814 29552
rect 46134 29466 46188 29500
rect 46222 29466 46278 29500
rect 46312 29466 46368 29500
rect 46402 29466 46458 29500
rect 46492 29466 46548 29500
rect 46582 29466 46638 29500
rect 46672 29466 46728 29500
rect 46762 29466 46814 29500
rect 46134 29410 46814 29466
rect 46134 29376 46188 29410
rect 46222 29376 46278 29410
rect 46312 29376 46368 29410
rect 46402 29376 46458 29410
rect 46492 29376 46548 29410
rect 46582 29376 46638 29410
rect 46672 29376 46728 29410
rect 46762 29376 46814 29410
rect 46134 29320 46814 29376
rect 46134 29286 46188 29320
rect 46222 29286 46278 29320
rect 46312 29286 46368 29320
rect 46402 29286 46458 29320
rect 46492 29286 46548 29320
rect 46582 29286 46638 29320
rect 46672 29286 46728 29320
rect 46762 29286 46814 29320
rect 46134 29230 46814 29286
rect 46134 29196 46188 29230
rect 46222 29196 46278 29230
rect 46312 29196 46368 29230
rect 46402 29196 46458 29230
rect 46492 29196 46548 29230
rect 46582 29196 46638 29230
rect 46672 29196 46728 29230
rect 46762 29196 46814 29230
rect 46134 29140 46814 29196
rect 46134 29106 46188 29140
rect 46222 29106 46278 29140
rect 46312 29106 46368 29140
rect 46402 29106 46458 29140
rect 46492 29106 46548 29140
rect 46582 29106 46638 29140
rect 46672 29106 46728 29140
rect 46762 29106 46814 29140
rect 46134 29050 46814 29106
rect 46134 29016 46188 29050
rect 46222 29016 46278 29050
rect 46312 29016 46368 29050
rect 46402 29016 46458 29050
rect 46492 29016 46548 29050
rect 46582 29016 46638 29050
rect 46672 29016 46728 29050
rect 46762 29016 46814 29050
rect 46134 28960 46814 29016
rect 46134 28926 46188 28960
rect 46222 28926 46278 28960
rect 46312 28926 46368 28960
rect 46402 28926 46458 28960
rect 46492 28926 46548 28960
rect 46582 28926 46638 28960
rect 46672 28926 46728 28960
rect 46762 28926 46814 28960
rect 46134 28872 46814 28926
rect 47474 29500 48154 29552
rect 47474 29466 47528 29500
rect 47562 29466 47618 29500
rect 47652 29466 47708 29500
rect 47742 29466 47798 29500
rect 47832 29466 47888 29500
rect 47922 29466 47978 29500
rect 48012 29466 48068 29500
rect 48102 29466 48154 29500
rect 47474 29410 48154 29466
rect 47474 29376 47528 29410
rect 47562 29376 47618 29410
rect 47652 29376 47708 29410
rect 47742 29376 47798 29410
rect 47832 29376 47888 29410
rect 47922 29376 47978 29410
rect 48012 29376 48068 29410
rect 48102 29376 48154 29410
rect 47474 29320 48154 29376
rect 47474 29286 47528 29320
rect 47562 29286 47618 29320
rect 47652 29286 47708 29320
rect 47742 29286 47798 29320
rect 47832 29286 47888 29320
rect 47922 29286 47978 29320
rect 48012 29286 48068 29320
rect 48102 29286 48154 29320
rect 47474 29230 48154 29286
rect 47474 29196 47528 29230
rect 47562 29196 47618 29230
rect 47652 29196 47708 29230
rect 47742 29196 47798 29230
rect 47832 29196 47888 29230
rect 47922 29196 47978 29230
rect 48012 29196 48068 29230
rect 48102 29196 48154 29230
rect 47474 29140 48154 29196
rect 47474 29106 47528 29140
rect 47562 29106 47618 29140
rect 47652 29106 47708 29140
rect 47742 29106 47798 29140
rect 47832 29106 47888 29140
rect 47922 29106 47978 29140
rect 48012 29106 48068 29140
rect 48102 29106 48154 29140
rect 47474 29050 48154 29106
rect 47474 29016 47528 29050
rect 47562 29016 47618 29050
rect 47652 29016 47708 29050
rect 47742 29016 47798 29050
rect 47832 29016 47888 29050
rect 47922 29016 47978 29050
rect 48012 29016 48068 29050
rect 48102 29016 48154 29050
rect 47474 28960 48154 29016
rect 47474 28926 47528 28960
rect 47562 28926 47618 28960
rect 47652 28926 47708 28960
rect 47742 28926 47798 28960
rect 47832 28926 47888 28960
rect 47922 28926 47978 28960
rect 48012 28926 48068 28960
rect 48102 28926 48154 28960
rect 47474 28872 48154 28926
rect 48814 29500 49494 29552
rect 48814 29466 48868 29500
rect 48902 29466 48958 29500
rect 48992 29466 49048 29500
rect 49082 29466 49138 29500
rect 49172 29466 49228 29500
rect 49262 29466 49318 29500
rect 49352 29466 49408 29500
rect 49442 29466 49494 29500
rect 48814 29410 49494 29466
rect 48814 29376 48868 29410
rect 48902 29376 48958 29410
rect 48992 29376 49048 29410
rect 49082 29376 49138 29410
rect 49172 29376 49228 29410
rect 49262 29376 49318 29410
rect 49352 29376 49408 29410
rect 49442 29376 49494 29410
rect 48814 29320 49494 29376
rect 48814 29286 48868 29320
rect 48902 29286 48958 29320
rect 48992 29286 49048 29320
rect 49082 29286 49138 29320
rect 49172 29286 49228 29320
rect 49262 29286 49318 29320
rect 49352 29286 49408 29320
rect 49442 29286 49494 29320
rect 48814 29230 49494 29286
rect 48814 29196 48868 29230
rect 48902 29196 48958 29230
rect 48992 29196 49048 29230
rect 49082 29196 49138 29230
rect 49172 29196 49228 29230
rect 49262 29196 49318 29230
rect 49352 29196 49408 29230
rect 49442 29196 49494 29230
rect 48814 29140 49494 29196
rect 48814 29106 48868 29140
rect 48902 29106 48958 29140
rect 48992 29106 49048 29140
rect 49082 29106 49138 29140
rect 49172 29106 49228 29140
rect 49262 29106 49318 29140
rect 49352 29106 49408 29140
rect 49442 29106 49494 29140
rect 48814 29050 49494 29106
rect 48814 29016 48868 29050
rect 48902 29016 48958 29050
rect 48992 29016 49048 29050
rect 49082 29016 49138 29050
rect 49172 29016 49228 29050
rect 49262 29016 49318 29050
rect 49352 29016 49408 29050
rect 49442 29016 49494 29050
rect 48814 28960 49494 29016
rect 48814 28926 48868 28960
rect 48902 28926 48958 28960
rect 48992 28926 49048 28960
rect 49082 28926 49138 28960
rect 49172 28926 49228 28960
rect 49262 28926 49318 28960
rect 49352 28926 49408 28960
rect 49442 28926 49494 28960
rect 48814 28872 49494 28926
rect 50154 29500 50834 29552
rect 50154 29466 50208 29500
rect 50242 29466 50298 29500
rect 50332 29466 50388 29500
rect 50422 29466 50478 29500
rect 50512 29466 50568 29500
rect 50602 29466 50658 29500
rect 50692 29466 50748 29500
rect 50782 29466 50834 29500
rect 50154 29410 50834 29466
rect 50154 29376 50208 29410
rect 50242 29376 50298 29410
rect 50332 29376 50388 29410
rect 50422 29376 50478 29410
rect 50512 29376 50568 29410
rect 50602 29376 50658 29410
rect 50692 29376 50748 29410
rect 50782 29376 50834 29410
rect 50154 29320 50834 29376
rect 50154 29286 50208 29320
rect 50242 29286 50298 29320
rect 50332 29286 50388 29320
rect 50422 29286 50478 29320
rect 50512 29286 50568 29320
rect 50602 29286 50658 29320
rect 50692 29286 50748 29320
rect 50782 29286 50834 29320
rect 50154 29230 50834 29286
rect 50154 29196 50208 29230
rect 50242 29196 50298 29230
rect 50332 29196 50388 29230
rect 50422 29196 50478 29230
rect 50512 29196 50568 29230
rect 50602 29196 50658 29230
rect 50692 29196 50748 29230
rect 50782 29196 50834 29230
rect 50154 29140 50834 29196
rect 50154 29106 50208 29140
rect 50242 29106 50298 29140
rect 50332 29106 50388 29140
rect 50422 29106 50478 29140
rect 50512 29106 50568 29140
rect 50602 29106 50658 29140
rect 50692 29106 50748 29140
rect 50782 29106 50834 29140
rect 50154 29050 50834 29106
rect 50154 29016 50208 29050
rect 50242 29016 50298 29050
rect 50332 29016 50388 29050
rect 50422 29016 50478 29050
rect 50512 29016 50568 29050
rect 50602 29016 50658 29050
rect 50692 29016 50748 29050
rect 50782 29016 50834 29050
rect 50154 28960 50834 29016
rect 50154 28926 50208 28960
rect 50242 28926 50298 28960
rect 50332 28926 50388 28960
rect 50422 28926 50478 28960
rect 50512 28926 50568 28960
rect 50602 28926 50658 28960
rect 50692 28926 50748 28960
rect 50782 28926 50834 28960
rect 50154 28872 50834 28926
rect 51494 29500 52174 29552
rect 51494 29466 51548 29500
rect 51582 29466 51638 29500
rect 51672 29466 51728 29500
rect 51762 29466 51818 29500
rect 51852 29466 51908 29500
rect 51942 29466 51998 29500
rect 52032 29466 52088 29500
rect 52122 29466 52174 29500
rect 51494 29410 52174 29466
rect 51494 29376 51548 29410
rect 51582 29376 51638 29410
rect 51672 29376 51728 29410
rect 51762 29376 51818 29410
rect 51852 29376 51908 29410
rect 51942 29376 51998 29410
rect 52032 29376 52088 29410
rect 52122 29376 52174 29410
rect 51494 29320 52174 29376
rect 51494 29286 51548 29320
rect 51582 29286 51638 29320
rect 51672 29286 51728 29320
rect 51762 29286 51818 29320
rect 51852 29286 51908 29320
rect 51942 29286 51998 29320
rect 52032 29286 52088 29320
rect 52122 29286 52174 29320
rect 51494 29230 52174 29286
rect 51494 29196 51548 29230
rect 51582 29196 51638 29230
rect 51672 29196 51728 29230
rect 51762 29196 51818 29230
rect 51852 29196 51908 29230
rect 51942 29196 51998 29230
rect 52032 29196 52088 29230
rect 52122 29196 52174 29230
rect 51494 29140 52174 29196
rect 51494 29106 51548 29140
rect 51582 29106 51638 29140
rect 51672 29106 51728 29140
rect 51762 29106 51818 29140
rect 51852 29106 51908 29140
rect 51942 29106 51998 29140
rect 52032 29106 52088 29140
rect 52122 29106 52174 29140
rect 51494 29050 52174 29106
rect 51494 29016 51548 29050
rect 51582 29016 51638 29050
rect 51672 29016 51728 29050
rect 51762 29016 51818 29050
rect 51852 29016 51908 29050
rect 51942 29016 51998 29050
rect 52032 29016 52088 29050
rect 52122 29016 52174 29050
rect 51494 28960 52174 29016
rect 51494 28926 51548 28960
rect 51582 28926 51638 28960
rect 51672 28926 51728 28960
rect 51762 28926 51818 28960
rect 51852 28926 51908 28960
rect 51942 28926 51998 28960
rect 52032 28926 52088 28960
rect 52122 28926 52174 28960
rect 51494 28872 52174 28926
rect 24865 18621 24923 18637
rect 24865 18587 24877 18621
rect 24911 18587 24923 18621
rect 24865 18553 24923 18587
rect 24865 18519 24877 18553
rect 24911 18519 24923 18553
rect 24865 18485 24923 18519
rect 24865 18451 24877 18485
rect 24911 18451 24923 18485
rect 24865 18417 24923 18451
rect 24865 18383 24877 18417
rect 24911 18383 24923 18417
rect 24865 18349 24923 18383
rect 24865 18315 24877 18349
rect 24911 18315 24923 18349
rect 24865 18281 24923 18315
rect 24865 18247 24877 18281
rect 24911 18247 24923 18281
rect 24865 18213 24923 18247
rect 24865 18179 24877 18213
rect 24911 18179 24923 18213
rect 24865 18145 24923 18179
rect 24865 18111 24877 18145
rect 24911 18111 24923 18145
rect 24865 18077 24923 18111
rect 24865 18043 24877 18077
rect 24911 18043 24923 18077
rect 24865 18009 24923 18043
rect 24865 17975 24877 18009
rect 24911 17975 24923 18009
rect 24865 17941 24923 17975
rect 24865 17907 24877 17941
rect 24911 17907 24923 17941
rect 24865 17873 24923 17907
rect 24865 17839 24877 17873
rect 24911 17839 24923 17873
rect 24865 17805 24923 17839
rect 24865 17771 24877 17805
rect 24911 17771 24923 17805
rect 24865 17737 24923 17771
rect 24865 17703 24877 17737
rect 24911 17703 24923 17737
rect 24865 17669 24923 17703
rect 24865 17635 24877 17669
rect 24911 17635 24923 17669
rect 24865 17601 24923 17635
rect 24865 17567 24877 17601
rect 24911 17567 24923 17601
rect 24865 17533 24923 17567
rect 24865 17499 24877 17533
rect 24911 17499 24923 17533
rect 24865 17465 24923 17499
rect 24865 17431 24877 17465
rect 24911 17431 24923 17465
rect 24865 17397 24923 17431
rect 24865 17363 24877 17397
rect 24911 17363 24923 17397
rect 24865 17347 24923 17363
rect 25323 18621 25381 18637
rect 25323 18587 25335 18621
rect 25369 18587 25381 18621
rect 25323 18553 25381 18587
rect 25323 18519 25335 18553
rect 25369 18519 25381 18553
rect 25323 18485 25381 18519
rect 25323 18451 25335 18485
rect 25369 18451 25381 18485
rect 25323 18417 25381 18451
rect 25323 18383 25335 18417
rect 25369 18383 25381 18417
rect 25323 18349 25381 18383
rect 25323 18315 25335 18349
rect 25369 18315 25381 18349
rect 25323 18281 25381 18315
rect 25323 18247 25335 18281
rect 25369 18247 25381 18281
rect 25323 18213 25381 18247
rect 25323 18179 25335 18213
rect 25369 18179 25381 18213
rect 25323 18145 25381 18179
rect 25323 18111 25335 18145
rect 25369 18111 25381 18145
rect 25323 18077 25381 18111
rect 25323 18043 25335 18077
rect 25369 18043 25381 18077
rect 25323 18009 25381 18043
rect 25323 17975 25335 18009
rect 25369 17975 25381 18009
rect 25323 17941 25381 17975
rect 25323 17907 25335 17941
rect 25369 17907 25381 17941
rect 25323 17873 25381 17907
rect 25323 17839 25335 17873
rect 25369 17839 25381 17873
rect 25323 17805 25381 17839
rect 25323 17771 25335 17805
rect 25369 17771 25381 17805
rect 25323 17737 25381 17771
rect 25323 17703 25335 17737
rect 25369 17703 25381 17737
rect 25323 17669 25381 17703
rect 25323 17635 25335 17669
rect 25369 17635 25381 17669
rect 25323 17601 25381 17635
rect 25323 17567 25335 17601
rect 25369 17567 25381 17601
rect 25323 17533 25381 17567
rect 25323 17499 25335 17533
rect 25369 17499 25381 17533
rect 25323 17465 25381 17499
rect 25323 17431 25335 17465
rect 25369 17431 25381 17465
rect 25323 17397 25381 17431
rect 25323 17363 25335 17397
rect 25369 17363 25381 17397
rect 25323 17347 25381 17363
rect 25781 18621 25839 18637
rect 25781 18587 25793 18621
rect 25827 18587 25839 18621
rect 25781 18553 25839 18587
rect 25781 18519 25793 18553
rect 25827 18519 25839 18553
rect 25781 18485 25839 18519
rect 25781 18451 25793 18485
rect 25827 18451 25839 18485
rect 25781 18417 25839 18451
rect 25781 18383 25793 18417
rect 25827 18383 25839 18417
rect 25781 18349 25839 18383
rect 25781 18315 25793 18349
rect 25827 18315 25839 18349
rect 25781 18281 25839 18315
rect 25781 18247 25793 18281
rect 25827 18247 25839 18281
rect 25781 18213 25839 18247
rect 25781 18179 25793 18213
rect 25827 18179 25839 18213
rect 25781 18145 25839 18179
rect 25781 18111 25793 18145
rect 25827 18111 25839 18145
rect 25781 18077 25839 18111
rect 25781 18043 25793 18077
rect 25827 18043 25839 18077
rect 25781 18009 25839 18043
rect 25781 17975 25793 18009
rect 25827 17975 25839 18009
rect 25781 17941 25839 17975
rect 25781 17907 25793 17941
rect 25827 17907 25839 17941
rect 25781 17873 25839 17907
rect 25781 17839 25793 17873
rect 25827 17839 25839 17873
rect 25781 17805 25839 17839
rect 25781 17771 25793 17805
rect 25827 17771 25839 17805
rect 25781 17737 25839 17771
rect 25781 17703 25793 17737
rect 25827 17703 25839 17737
rect 25781 17669 25839 17703
rect 25781 17635 25793 17669
rect 25827 17635 25839 17669
rect 25781 17601 25839 17635
rect 25781 17567 25793 17601
rect 25827 17567 25839 17601
rect 25781 17533 25839 17567
rect 25781 17499 25793 17533
rect 25827 17499 25839 17533
rect 25781 17465 25839 17499
rect 25781 17431 25793 17465
rect 25827 17431 25839 17465
rect 25781 17397 25839 17431
rect 25781 17363 25793 17397
rect 25827 17363 25839 17397
rect 25781 17347 25839 17363
rect 26239 18621 26297 18637
rect 26239 18587 26251 18621
rect 26285 18587 26297 18621
rect 26239 18553 26297 18587
rect 26239 18519 26251 18553
rect 26285 18519 26297 18553
rect 26239 18485 26297 18519
rect 26239 18451 26251 18485
rect 26285 18451 26297 18485
rect 26239 18417 26297 18451
rect 26239 18383 26251 18417
rect 26285 18383 26297 18417
rect 26239 18349 26297 18383
rect 26239 18315 26251 18349
rect 26285 18315 26297 18349
rect 26239 18281 26297 18315
rect 26239 18247 26251 18281
rect 26285 18247 26297 18281
rect 26239 18213 26297 18247
rect 26239 18179 26251 18213
rect 26285 18179 26297 18213
rect 26239 18145 26297 18179
rect 26239 18111 26251 18145
rect 26285 18111 26297 18145
rect 26239 18077 26297 18111
rect 26239 18043 26251 18077
rect 26285 18043 26297 18077
rect 26239 18009 26297 18043
rect 26239 17975 26251 18009
rect 26285 17975 26297 18009
rect 26239 17941 26297 17975
rect 26239 17907 26251 17941
rect 26285 17907 26297 17941
rect 26239 17873 26297 17907
rect 26239 17839 26251 17873
rect 26285 17839 26297 17873
rect 26239 17805 26297 17839
rect 26239 17771 26251 17805
rect 26285 17771 26297 17805
rect 26239 17737 26297 17771
rect 26239 17703 26251 17737
rect 26285 17703 26297 17737
rect 26239 17669 26297 17703
rect 26239 17635 26251 17669
rect 26285 17635 26297 17669
rect 26239 17601 26297 17635
rect 26239 17567 26251 17601
rect 26285 17567 26297 17601
rect 26239 17533 26297 17567
rect 26239 17499 26251 17533
rect 26285 17499 26297 17533
rect 26239 17465 26297 17499
rect 26239 17431 26251 17465
rect 26285 17431 26297 17465
rect 26239 17397 26297 17431
rect 26239 17363 26251 17397
rect 26285 17363 26297 17397
rect 26239 17347 26297 17363
rect 26697 18621 26755 18637
rect 26697 18587 26709 18621
rect 26743 18587 26755 18621
rect 26697 18553 26755 18587
rect 26697 18519 26709 18553
rect 26743 18519 26755 18553
rect 26697 18485 26755 18519
rect 26697 18451 26709 18485
rect 26743 18451 26755 18485
rect 26697 18417 26755 18451
rect 26697 18383 26709 18417
rect 26743 18383 26755 18417
rect 26697 18349 26755 18383
rect 26697 18315 26709 18349
rect 26743 18315 26755 18349
rect 26697 18281 26755 18315
rect 26697 18247 26709 18281
rect 26743 18247 26755 18281
rect 26697 18213 26755 18247
rect 26697 18179 26709 18213
rect 26743 18179 26755 18213
rect 26697 18145 26755 18179
rect 26697 18111 26709 18145
rect 26743 18111 26755 18145
rect 26697 18077 26755 18111
rect 26697 18043 26709 18077
rect 26743 18043 26755 18077
rect 26697 18009 26755 18043
rect 26697 17975 26709 18009
rect 26743 17975 26755 18009
rect 26697 17941 26755 17975
rect 26697 17907 26709 17941
rect 26743 17907 26755 17941
rect 26697 17873 26755 17907
rect 26697 17839 26709 17873
rect 26743 17839 26755 17873
rect 26697 17805 26755 17839
rect 26697 17771 26709 17805
rect 26743 17771 26755 17805
rect 26697 17737 26755 17771
rect 26697 17703 26709 17737
rect 26743 17703 26755 17737
rect 26697 17669 26755 17703
rect 26697 17635 26709 17669
rect 26743 17635 26755 17669
rect 26697 17601 26755 17635
rect 26697 17567 26709 17601
rect 26743 17567 26755 17601
rect 26697 17533 26755 17567
rect 26697 17499 26709 17533
rect 26743 17499 26755 17533
rect 26697 17465 26755 17499
rect 26697 17431 26709 17465
rect 26743 17431 26755 17465
rect 26697 17397 26755 17431
rect 26697 17363 26709 17397
rect 26743 17363 26755 17397
rect 26697 17347 26755 17363
rect 27155 18621 27213 18637
rect 27155 18587 27167 18621
rect 27201 18587 27213 18621
rect 27155 18553 27213 18587
rect 27155 18519 27167 18553
rect 27201 18519 27213 18553
rect 27155 18485 27213 18519
rect 27155 18451 27167 18485
rect 27201 18451 27213 18485
rect 27155 18417 27213 18451
rect 27155 18383 27167 18417
rect 27201 18383 27213 18417
rect 27155 18349 27213 18383
rect 27155 18315 27167 18349
rect 27201 18315 27213 18349
rect 27155 18281 27213 18315
rect 27155 18247 27167 18281
rect 27201 18247 27213 18281
rect 27155 18213 27213 18247
rect 27155 18179 27167 18213
rect 27201 18179 27213 18213
rect 27155 18145 27213 18179
rect 27155 18111 27167 18145
rect 27201 18111 27213 18145
rect 27155 18077 27213 18111
rect 27155 18043 27167 18077
rect 27201 18043 27213 18077
rect 27155 18009 27213 18043
rect 27155 17975 27167 18009
rect 27201 17975 27213 18009
rect 27155 17941 27213 17975
rect 27155 17907 27167 17941
rect 27201 17907 27213 17941
rect 27155 17873 27213 17907
rect 27155 17839 27167 17873
rect 27201 17839 27213 17873
rect 27155 17805 27213 17839
rect 27155 17771 27167 17805
rect 27201 17771 27213 17805
rect 27155 17737 27213 17771
rect 27155 17703 27167 17737
rect 27201 17703 27213 17737
rect 27155 17669 27213 17703
rect 27155 17635 27167 17669
rect 27201 17635 27213 17669
rect 27155 17601 27213 17635
rect 27155 17567 27167 17601
rect 27201 17567 27213 17601
rect 27155 17533 27213 17567
rect 27155 17499 27167 17533
rect 27201 17499 27213 17533
rect 27155 17465 27213 17499
rect 27155 17431 27167 17465
rect 27201 17431 27213 17465
rect 27155 17397 27213 17431
rect 27155 17363 27167 17397
rect 27201 17363 27213 17397
rect 27155 17347 27213 17363
rect 27613 18621 27671 18637
rect 27613 18587 27625 18621
rect 27659 18587 27671 18621
rect 27613 18553 27671 18587
rect 27613 18519 27625 18553
rect 27659 18519 27671 18553
rect 27613 18485 27671 18519
rect 27613 18451 27625 18485
rect 27659 18451 27671 18485
rect 27613 18417 27671 18451
rect 27613 18383 27625 18417
rect 27659 18383 27671 18417
rect 27613 18349 27671 18383
rect 27613 18315 27625 18349
rect 27659 18315 27671 18349
rect 27613 18281 27671 18315
rect 27613 18247 27625 18281
rect 27659 18247 27671 18281
rect 27613 18213 27671 18247
rect 27613 18179 27625 18213
rect 27659 18179 27671 18213
rect 27613 18145 27671 18179
rect 27613 18111 27625 18145
rect 27659 18111 27671 18145
rect 27613 18077 27671 18111
rect 27613 18043 27625 18077
rect 27659 18043 27671 18077
rect 27613 18009 27671 18043
rect 27613 17975 27625 18009
rect 27659 17975 27671 18009
rect 27613 17941 27671 17975
rect 27613 17907 27625 17941
rect 27659 17907 27671 17941
rect 27613 17873 27671 17907
rect 27613 17839 27625 17873
rect 27659 17839 27671 17873
rect 27613 17805 27671 17839
rect 27613 17771 27625 17805
rect 27659 17771 27671 17805
rect 27613 17737 27671 17771
rect 27613 17703 27625 17737
rect 27659 17703 27671 17737
rect 27613 17669 27671 17703
rect 27613 17635 27625 17669
rect 27659 17635 27671 17669
rect 27613 17601 27671 17635
rect 27613 17567 27625 17601
rect 27659 17567 27671 17601
rect 27613 17533 27671 17567
rect 27613 17499 27625 17533
rect 27659 17499 27671 17533
rect 27613 17465 27671 17499
rect 27613 17431 27625 17465
rect 27659 17431 27671 17465
rect 27613 17397 27671 17431
rect 27613 17363 27625 17397
rect 27659 17363 27671 17397
rect 27613 17347 27671 17363
rect 28071 18621 28129 18637
rect 28071 18587 28083 18621
rect 28117 18587 28129 18621
rect 28071 18553 28129 18587
rect 28071 18519 28083 18553
rect 28117 18519 28129 18553
rect 28071 18485 28129 18519
rect 28071 18451 28083 18485
rect 28117 18451 28129 18485
rect 28071 18417 28129 18451
rect 28071 18383 28083 18417
rect 28117 18383 28129 18417
rect 28071 18349 28129 18383
rect 28071 18315 28083 18349
rect 28117 18315 28129 18349
rect 28071 18281 28129 18315
rect 28071 18247 28083 18281
rect 28117 18247 28129 18281
rect 28071 18213 28129 18247
rect 28071 18179 28083 18213
rect 28117 18179 28129 18213
rect 28071 18145 28129 18179
rect 28071 18111 28083 18145
rect 28117 18111 28129 18145
rect 28071 18077 28129 18111
rect 28071 18043 28083 18077
rect 28117 18043 28129 18077
rect 28071 18009 28129 18043
rect 28071 17975 28083 18009
rect 28117 17975 28129 18009
rect 28071 17941 28129 17975
rect 28071 17907 28083 17941
rect 28117 17907 28129 17941
rect 28071 17873 28129 17907
rect 28071 17839 28083 17873
rect 28117 17839 28129 17873
rect 28071 17805 28129 17839
rect 28071 17771 28083 17805
rect 28117 17771 28129 17805
rect 28071 17737 28129 17771
rect 28071 17703 28083 17737
rect 28117 17703 28129 17737
rect 28071 17669 28129 17703
rect 28071 17635 28083 17669
rect 28117 17635 28129 17669
rect 28071 17601 28129 17635
rect 28071 17567 28083 17601
rect 28117 17567 28129 17601
rect 28071 17533 28129 17567
rect 28071 17499 28083 17533
rect 28117 17499 28129 17533
rect 28071 17465 28129 17499
rect 28071 17431 28083 17465
rect 28117 17431 28129 17465
rect 28071 17397 28129 17431
rect 28071 17363 28083 17397
rect 28117 17363 28129 17397
rect 28071 17347 28129 17363
rect 28529 18621 28587 18637
rect 28529 18587 28541 18621
rect 28575 18587 28587 18621
rect 28529 18553 28587 18587
rect 28529 18519 28541 18553
rect 28575 18519 28587 18553
rect 28529 18485 28587 18519
rect 28529 18451 28541 18485
rect 28575 18451 28587 18485
rect 28529 18417 28587 18451
rect 28529 18383 28541 18417
rect 28575 18383 28587 18417
rect 28529 18349 28587 18383
rect 28529 18315 28541 18349
rect 28575 18315 28587 18349
rect 28529 18281 28587 18315
rect 28529 18247 28541 18281
rect 28575 18247 28587 18281
rect 28529 18213 28587 18247
rect 28529 18179 28541 18213
rect 28575 18179 28587 18213
rect 28529 18145 28587 18179
rect 28529 18111 28541 18145
rect 28575 18111 28587 18145
rect 28529 18077 28587 18111
rect 28529 18043 28541 18077
rect 28575 18043 28587 18077
rect 28529 18009 28587 18043
rect 28529 17975 28541 18009
rect 28575 17975 28587 18009
rect 28529 17941 28587 17975
rect 28529 17907 28541 17941
rect 28575 17907 28587 17941
rect 28529 17873 28587 17907
rect 28529 17839 28541 17873
rect 28575 17839 28587 17873
rect 28529 17805 28587 17839
rect 28529 17771 28541 17805
rect 28575 17771 28587 17805
rect 28529 17737 28587 17771
rect 28529 17703 28541 17737
rect 28575 17703 28587 17737
rect 28529 17669 28587 17703
rect 28529 17635 28541 17669
rect 28575 17635 28587 17669
rect 28529 17601 28587 17635
rect 28529 17567 28541 17601
rect 28575 17567 28587 17601
rect 28529 17533 28587 17567
rect 28529 17499 28541 17533
rect 28575 17499 28587 17533
rect 28529 17465 28587 17499
rect 28529 17431 28541 17465
rect 28575 17431 28587 17465
rect 28529 17397 28587 17431
rect 28529 17363 28541 17397
rect 28575 17363 28587 17397
rect 28529 17347 28587 17363
rect 28987 18621 29045 18637
rect 28987 18587 28999 18621
rect 29033 18587 29045 18621
rect 28987 18553 29045 18587
rect 28987 18519 28999 18553
rect 29033 18519 29045 18553
rect 28987 18485 29045 18519
rect 28987 18451 28999 18485
rect 29033 18451 29045 18485
rect 28987 18417 29045 18451
rect 28987 18383 28999 18417
rect 29033 18383 29045 18417
rect 28987 18349 29045 18383
rect 28987 18315 28999 18349
rect 29033 18315 29045 18349
rect 28987 18281 29045 18315
rect 28987 18247 28999 18281
rect 29033 18247 29045 18281
rect 28987 18213 29045 18247
rect 28987 18179 28999 18213
rect 29033 18179 29045 18213
rect 28987 18145 29045 18179
rect 28987 18111 28999 18145
rect 29033 18111 29045 18145
rect 28987 18077 29045 18111
rect 28987 18043 28999 18077
rect 29033 18043 29045 18077
rect 28987 18009 29045 18043
rect 28987 17975 28999 18009
rect 29033 17975 29045 18009
rect 28987 17941 29045 17975
rect 28987 17907 28999 17941
rect 29033 17907 29045 17941
rect 28987 17873 29045 17907
rect 28987 17839 28999 17873
rect 29033 17839 29045 17873
rect 28987 17805 29045 17839
rect 28987 17771 28999 17805
rect 29033 17771 29045 17805
rect 28987 17737 29045 17771
rect 28987 17703 28999 17737
rect 29033 17703 29045 17737
rect 28987 17669 29045 17703
rect 28987 17635 28999 17669
rect 29033 17635 29045 17669
rect 28987 17601 29045 17635
rect 28987 17567 28999 17601
rect 29033 17567 29045 17601
rect 28987 17533 29045 17567
rect 28987 17499 28999 17533
rect 29033 17499 29045 17533
rect 28987 17465 29045 17499
rect 28987 17431 28999 17465
rect 29033 17431 29045 17465
rect 28987 17397 29045 17431
rect 28987 17363 28999 17397
rect 29033 17363 29045 17397
rect 28987 17347 29045 17363
rect 29445 18621 29503 18637
rect 29445 18587 29457 18621
rect 29491 18587 29503 18621
rect 29445 18553 29503 18587
rect 29445 18519 29457 18553
rect 29491 18519 29503 18553
rect 29445 18485 29503 18519
rect 29445 18451 29457 18485
rect 29491 18451 29503 18485
rect 29445 18417 29503 18451
rect 29445 18383 29457 18417
rect 29491 18383 29503 18417
rect 29445 18349 29503 18383
rect 29445 18315 29457 18349
rect 29491 18315 29503 18349
rect 29445 18281 29503 18315
rect 29445 18247 29457 18281
rect 29491 18247 29503 18281
rect 29445 18213 29503 18247
rect 29445 18179 29457 18213
rect 29491 18179 29503 18213
rect 29445 18145 29503 18179
rect 29445 18111 29457 18145
rect 29491 18111 29503 18145
rect 29445 18077 29503 18111
rect 29445 18043 29457 18077
rect 29491 18043 29503 18077
rect 29445 18009 29503 18043
rect 29445 17975 29457 18009
rect 29491 17975 29503 18009
rect 29445 17941 29503 17975
rect 29445 17907 29457 17941
rect 29491 17907 29503 17941
rect 29445 17873 29503 17907
rect 29445 17839 29457 17873
rect 29491 17839 29503 17873
rect 29445 17805 29503 17839
rect 29445 17771 29457 17805
rect 29491 17771 29503 17805
rect 29445 17737 29503 17771
rect 29445 17703 29457 17737
rect 29491 17703 29503 17737
rect 29445 17669 29503 17703
rect 29445 17635 29457 17669
rect 29491 17635 29503 17669
rect 29445 17601 29503 17635
rect 29445 17567 29457 17601
rect 29491 17567 29503 17601
rect 29445 17533 29503 17567
rect 29445 17499 29457 17533
rect 29491 17499 29503 17533
rect 29445 17465 29503 17499
rect 29445 17431 29457 17465
rect 29491 17431 29503 17465
rect 29445 17397 29503 17431
rect 29445 17363 29457 17397
rect 29491 17363 29503 17397
rect 29445 17347 29503 17363
rect 29903 18621 29961 18637
rect 29903 18587 29915 18621
rect 29949 18587 29961 18621
rect 29903 18553 29961 18587
rect 29903 18519 29915 18553
rect 29949 18519 29961 18553
rect 29903 18485 29961 18519
rect 29903 18451 29915 18485
rect 29949 18451 29961 18485
rect 29903 18417 29961 18451
rect 29903 18383 29915 18417
rect 29949 18383 29961 18417
rect 29903 18349 29961 18383
rect 29903 18315 29915 18349
rect 29949 18315 29961 18349
rect 29903 18281 29961 18315
rect 29903 18247 29915 18281
rect 29949 18247 29961 18281
rect 29903 18213 29961 18247
rect 29903 18179 29915 18213
rect 29949 18179 29961 18213
rect 29903 18145 29961 18179
rect 29903 18111 29915 18145
rect 29949 18111 29961 18145
rect 29903 18077 29961 18111
rect 29903 18043 29915 18077
rect 29949 18043 29961 18077
rect 29903 18009 29961 18043
rect 29903 17975 29915 18009
rect 29949 17975 29961 18009
rect 29903 17941 29961 17975
rect 29903 17907 29915 17941
rect 29949 17907 29961 17941
rect 29903 17873 29961 17907
rect 29903 17839 29915 17873
rect 29949 17839 29961 17873
rect 29903 17805 29961 17839
rect 29903 17771 29915 17805
rect 29949 17771 29961 17805
rect 29903 17737 29961 17771
rect 29903 17703 29915 17737
rect 29949 17703 29961 17737
rect 29903 17669 29961 17703
rect 29903 17635 29915 17669
rect 29949 17635 29961 17669
rect 29903 17601 29961 17635
rect 29903 17567 29915 17601
rect 29949 17567 29961 17601
rect 29903 17533 29961 17567
rect 29903 17499 29915 17533
rect 29949 17499 29961 17533
rect 29903 17465 29961 17499
rect 29903 17431 29915 17465
rect 29949 17431 29961 17465
rect 29903 17397 29961 17431
rect 29903 17363 29915 17397
rect 29949 17363 29961 17397
rect 29903 17347 29961 17363
rect 30361 18621 30419 18637
rect 30361 18587 30373 18621
rect 30407 18587 30419 18621
rect 30361 18553 30419 18587
rect 30361 18519 30373 18553
rect 30407 18519 30419 18553
rect 30361 18485 30419 18519
rect 30361 18451 30373 18485
rect 30407 18451 30419 18485
rect 30361 18417 30419 18451
rect 30361 18383 30373 18417
rect 30407 18383 30419 18417
rect 30361 18349 30419 18383
rect 30361 18315 30373 18349
rect 30407 18315 30419 18349
rect 30361 18281 30419 18315
rect 30361 18247 30373 18281
rect 30407 18247 30419 18281
rect 30361 18213 30419 18247
rect 30361 18179 30373 18213
rect 30407 18179 30419 18213
rect 30361 18145 30419 18179
rect 30361 18111 30373 18145
rect 30407 18111 30419 18145
rect 30361 18077 30419 18111
rect 30361 18043 30373 18077
rect 30407 18043 30419 18077
rect 30361 18009 30419 18043
rect 30361 17975 30373 18009
rect 30407 17975 30419 18009
rect 30361 17941 30419 17975
rect 30361 17907 30373 17941
rect 30407 17907 30419 17941
rect 30361 17873 30419 17907
rect 30361 17839 30373 17873
rect 30407 17839 30419 17873
rect 30361 17805 30419 17839
rect 30361 17771 30373 17805
rect 30407 17771 30419 17805
rect 30361 17737 30419 17771
rect 30361 17703 30373 17737
rect 30407 17703 30419 17737
rect 30361 17669 30419 17703
rect 30361 17635 30373 17669
rect 30407 17635 30419 17669
rect 30361 17601 30419 17635
rect 30361 17567 30373 17601
rect 30407 17567 30419 17601
rect 30361 17533 30419 17567
rect 30361 17499 30373 17533
rect 30407 17499 30419 17533
rect 30361 17465 30419 17499
rect 30361 17431 30373 17465
rect 30407 17431 30419 17465
rect 30361 17397 30419 17431
rect 30361 17363 30373 17397
rect 30407 17363 30419 17397
rect 30361 17347 30419 17363
rect 30819 18621 30877 18637
rect 30819 18587 30831 18621
rect 30865 18587 30877 18621
rect 30819 18553 30877 18587
rect 30819 18519 30831 18553
rect 30865 18519 30877 18553
rect 30819 18485 30877 18519
rect 30819 18451 30831 18485
rect 30865 18451 30877 18485
rect 30819 18417 30877 18451
rect 30819 18383 30831 18417
rect 30865 18383 30877 18417
rect 30819 18349 30877 18383
rect 30819 18315 30831 18349
rect 30865 18315 30877 18349
rect 30819 18281 30877 18315
rect 30819 18247 30831 18281
rect 30865 18247 30877 18281
rect 30819 18213 30877 18247
rect 30819 18179 30831 18213
rect 30865 18179 30877 18213
rect 30819 18145 30877 18179
rect 30819 18111 30831 18145
rect 30865 18111 30877 18145
rect 30819 18077 30877 18111
rect 30819 18043 30831 18077
rect 30865 18043 30877 18077
rect 30819 18009 30877 18043
rect 30819 17975 30831 18009
rect 30865 17975 30877 18009
rect 30819 17941 30877 17975
rect 30819 17907 30831 17941
rect 30865 17907 30877 17941
rect 30819 17873 30877 17907
rect 30819 17839 30831 17873
rect 30865 17839 30877 17873
rect 30819 17805 30877 17839
rect 30819 17771 30831 17805
rect 30865 17771 30877 17805
rect 30819 17737 30877 17771
rect 30819 17703 30831 17737
rect 30865 17703 30877 17737
rect 30819 17669 30877 17703
rect 30819 17635 30831 17669
rect 30865 17635 30877 17669
rect 30819 17601 30877 17635
rect 30819 17567 30831 17601
rect 30865 17567 30877 17601
rect 30819 17533 30877 17567
rect 30819 17499 30831 17533
rect 30865 17499 30877 17533
rect 30819 17465 30877 17499
rect 30819 17431 30831 17465
rect 30865 17431 30877 17465
rect 30819 17397 30877 17431
rect 30819 17363 30831 17397
rect 30865 17363 30877 17397
rect 30819 17347 30877 17363
rect 31277 18621 31335 18637
rect 31277 18587 31289 18621
rect 31323 18587 31335 18621
rect 31277 18553 31335 18587
rect 31277 18519 31289 18553
rect 31323 18519 31335 18553
rect 31277 18485 31335 18519
rect 31277 18451 31289 18485
rect 31323 18451 31335 18485
rect 31277 18417 31335 18451
rect 31277 18383 31289 18417
rect 31323 18383 31335 18417
rect 31277 18349 31335 18383
rect 31277 18315 31289 18349
rect 31323 18315 31335 18349
rect 31277 18281 31335 18315
rect 31277 18247 31289 18281
rect 31323 18247 31335 18281
rect 31277 18213 31335 18247
rect 31277 18179 31289 18213
rect 31323 18179 31335 18213
rect 31277 18145 31335 18179
rect 31277 18111 31289 18145
rect 31323 18111 31335 18145
rect 31277 18077 31335 18111
rect 31277 18043 31289 18077
rect 31323 18043 31335 18077
rect 31277 18009 31335 18043
rect 31277 17975 31289 18009
rect 31323 17975 31335 18009
rect 31277 17941 31335 17975
rect 31277 17907 31289 17941
rect 31323 17907 31335 17941
rect 31277 17873 31335 17907
rect 31277 17839 31289 17873
rect 31323 17839 31335 17873
rect 31277 17805 31335 17839
rect 31277 17771 31289 17805
rect 31323 17771 31335 17805
rect 31277 17737 31335 17771
rect 31277 17703 31289 17737
rect 31323 17703 31335 17737
rect 31277 17669 31335 17703
rect 31277 17635 31289 17669
rect 31323 17635 31335 17669
rect 31277 17601 31335 17635
rect 31277 17567 31289 17601
rect 31323 17567 31335 17601
rect 31277 17533 31335 17567
rect 31277 17499 31289 17533
rect 31323 17499 31335 17533
rect 31277 17465 31335 17499
rect 31277 17431 31289 17465
rect 31323 17431 31335 17465
rect 31277 17397 31335 17431
rect 31277 17363 31289 17397
rect 31323 17363 31335 17397
rect 31277 17347 31335 17363
rect 31735 18621 31793 18637
rect 31735 18587 31747 18621
rect 31781 18587 31793 18621
rect 31735 18553 31793 18587
rect 31735 18519 31747 18553
rect 31781 18519 31793 18553
rect 31735 18485 31793 18519
rect 31735 18451 31747 18485
rect 31781 18451 31793 18485
rect 31735 18417 31793 18451
rect 31735 18383 31747 18417
rect 31781 18383 31793 18417
rect 31735 18349 31793 18383
rect 31735 18315 31747 18349
rect 31781 18315 31793 18349
rect 31735 18281 31793 18315
rect 31735 18247 31747 18281
rect 31781 18247 31793 18281
rect 31735 18213 31793 18247
rect 31735 18179 31747 18213
rect 31781 18179 31793 18213
rect 31735 18145 31793 18179
rect 31735 18111 31747 18145
rect 31781 18111 31793 18145
rect 31735 18077 31793 18111
rect 31735 18043 31747 18077
rect 31781 18043 31793 18077
rect 31735 18009 31793 18043
rect 31735 17975 31747 18009
rect 31781 17975 31793 18009
rect 31735 17941 31793 17975
rect 31735 17907 31747 17941
rect 31781 17907 31793 17941
rect 31735 17873 31793 17907
rect 31735 17839 31747 17873
rect 31781 17839 31793 17873
rect 31735 17805 31793 17839
rect 31735 17771 31747 17805
rect 31781 17771 31793 17805
rect 31735 17737 31793 17771
rect 31735 17703 31747 17737
rect 31781 17703 31793 17737
rect 31735 17669 31793 17703
rect 31735 17635 31747 17669
rect 31781 17635 31793 17669
rect 31735 17601 31793 17635
rect 31735 17567 31747 17601
rect 31781 17567 31793 17601
rect 31735 17533 31793 17567
rect 31735 17499 31747 17533
rect 31781 17499 31793 17533
rect 31735 17465 31793 17499
rect 31735 17431 31747 17465
rect 31781 17431 31793 17465
rect 31735 17397 31793 17431
rect 31735 17363 31747 17397
rect 31781 17363 31793 17397
rect 31735 17347 31793 17363
rect 32193 18621 32251 18637
rect 32193 18587 32205 18621
rect 32239 18587 32251 18621
rect 32193 18553 32251 18587
rect 32193 18519 32205 18553
rect 32239 18519 32251 18553
rect 32193 18485 32251 18519
rect 32193 18451 32205 18485
rect 32239 18451 32251 18485
rect 32193 18417 32251 18451
rect 32193 18383 32205 18417
rect 32239 18383 32251 18417
rect 32193 18349 32251 18383
rect 32193 18315 32205 18349
rect 32239 18315 32251 18349
rect 32193 18281 32251 18315
rect 32193 18247 32205 18281
rect 32239 18247 32251 18281
rect 32193 18213 32251 18247
rect 32193 18179 32205 18213
rect 32239 18179 32251 18213
rect 32193 18145 32251 18179
rect 32193 18111 32205 18145
rect 32239 18111 32251 18145
rect 32193 18077 32251 18111
rect 32193 18043 32205 18077
rect 32239 18043 32251 18077
rect 32193 18009 32251 18043
rect 32193 17975 32205 18009
rect 32239 17975 32251 18009
rect 32193 17941 32251 17975
rect 32193 17907 32205 17941
rect 32239 17907 32251 17941
rect 32193 17873 32251 17907
rect 32193 17839 32205 17873
rect 32239 17839 32251 17873
rect 32193 17805 32251 17839
rect 32193 17771 32205 17805
rect 32239 17771 32251 17805
rect 32193 17737 32251 17771
rect 32193 17703 32205 17737
rect 32239 17703 32251 17737
rect 32193 17669 32251 17703
rect 32193 17635 32205 17669
rect 32239 17635 32251 17669
rect 32193 17601 32251 17635
rect 32193 17567 32205 17601
rect 32239 17567 32251 17601
rect 32193 17533 32251 17567
rect 32193 17499 32205 17533
rect 32239 17499 32251 17533
rect 32193 17465 32251 17499
rect 32193 17431 32205 17465
rect 32239 17431 32251 17465
rect 32193 17397 32251 17431
rect 32193 17363 32205 17397
rect 32239 17363 32251 17397
rect 32193 17347 32251 17363
rect 32651 18621 32709 18637
rect 32651 18587 32663 18621
rect 32697 18587 32709 18621
rect 32651 18553 32709 18587
rect 32651 18519 32663 18553
rect 32697 18519 32709 18553
rect 32651 18485 32709 18519
rect 32651 18451 32663 18485
rect 32697 18451 32709 18485
rect 32651 18417 32709 18451
rect 32651 18383 32663 18417
rect 32697 18383 32709 18417
rect 32651 18349 32709 18383
rect 32651 18315 32663 18349
rect 32697 18315 32709 18349
rect 32651 18281 32709 18315
rect 32651 18247 32663 18281
rect 32697 18247 32709 18281
rect 32651 18213 32709 18247
rect 32651 18179 32663 18213
rect 32697 18179 32709 18213
rect 32651 18145 32709 18179
rect 32651 18111 32663 18145
rect 32697 18111 32709 18145
rect 32651 18077 32709 18111
rect 32651 18043 32663 18077
rect 32697 18043 32709 18077
rect 32651 18009 32709 18043
rect 32651 17975 32663 18009
rect 32697 17975 32709 18009
rect 32651 17941 32709 17975
rect 32651 17907 32663 17941
rect 32697 17907 32709 17941
rect 32651 17873 32709 17907
rect 32651 17839 32663 17873
rect 32697 17839 32709 17873
rect 32651 17805 32709 17839
rect 32651 17771 32663 17805
rect 32697 17771 32709 17805
rect 32651 17737 32709 17771
rect 32651 17703 32663 17737
rect 32697 17703 32709 17737
rect 32651 17669 32709 17703
rect 32651 17635 32663 17669
rect 32697 17635 32709 17669
rect 32651 17601 32709 17635
rect 32651 17567 32663 17601
rect 32697 17567 32709 17601
rect 32651 17533 32709 17567
rect 32651 17499 32663 17533
rect 32697 17499 32709 17533
rect 32651 17465 32709 17499
rect 32651 17431 32663 17465
rect 32697 17431 32709 17465
rect 32651 17397 32709 17431
rect 32651 17363 32663 17397
rect 32697 17363 32709 17397
rect 32651 17347 32709 17363
rect 33109 18621 33167 18637
rect 33109 18587 33121 18621
rect 33155 18587 33167 18621
rect 33109 18553 33167 18587
rect 33109 18519 33121 18553
rect 33155 18519 33167 18553
rect 33109 18485 33167 18519
rect 33109 18451 33121 18485
rect 33155 18451 33167 18485
rect 33109 18417 33167 18451
rect 33109 18383 33121 18417
rect 33155 18383 33167 18417
rect 33109 18349 33167 18383
rect 33109 18315 33121 18349
rect 33155 18315 33167 18349
rect 33109 18281 33167 18315
rect 33109 18247 33121 18281
rect 33155 18247 33167 18281
rect 33109 18213 33167 18247
rect 33109 18179 33121 18213
rect 33155 18179 33167 18213
rect 33109 18145 33167 18179
rect 33109 18111 33121 18145
rect 33155 18111 33167 18145
rect 33109 18077 33167 18111
rect 33109 18043 33121 18077
rect 33155 18043 33167 18077
rect 33109 18009 33167 18043
rect 33109 17975 33121 18009
rect 33155 17975 33167 18009
rect 33109 17941 33167 17975
rect 33109 17907 33121 17941
rect 33155 17907 33167 17941
rect 33109 17873 33167 17907
rect 33109 17839 33121 17873
rect 33155 17839 33167 17873
rect 33109 17805 33167 17839
rect 33109 17771 33121 17805
rect 33155 17771 33167 17805
rect 33109 17737 33167 17771
rect 33109 17703 33121 17737
rect 33155 17703 33167 17737
rect 33109 17669 33167 17703
rect 33109 17635 33121 17669
rect 33155 17635 33167 17669
rect 33109 17601 33167 17635
rect 33109 17567 33121 17601
rect 33155 17567 33167 17601
rect 33109 17533 33167 17567
rect 33109 17499 33121 17533
rect 33155 17499 33167 17533
rect 33109 17465 33167 17499
rect 33109 17431 33121 17465
rect 33155 17431 33167 17465
rect 33109 17397 33167 17431
rect 33109 17363 33121 17397
rect 33155 17363 33167 17397
rect 33109 17347 33167 17363
rect 33567 18621 33625 18637
rect 33567 18587 33579 18621
rect 33613 18587 33625 18621
rect 33567 18553 33625 18587
rect 33567 18519 33579 18553
rect 33613 18519 33625 18553
rect 33567 18485 33625 18519
rect 33567 18451 33579 18485
rect 33613 18451 33625 18485
rect 33567 18417 33625 18451
rect 33567 18383 33579 18417
rect 33613 18383 33625 18417
rect 33567 18349 33625 18383
rect 33567 18315 33579 18349
rect 33613 18315 33625 18349
rect 33567 18281 33625 18315
rect 33567 18247 33579 18281
rect 33613 18247 33625 18281
rect 33567 18213 33625 18247
rect 33567 18179 33579 18213
rect 33613 18179 33625 18213
rect 33567 18145 33625 18179
rect 33567 18111 33579 18145
rect 33613 18111 33625 18145
rect 33567 18077 33625 18111
rect 33567 18043 33579 18077
rect 33613 18043 33625 18077
rect 33567 18009 33625 18043
rect 33567 17975 33579 18009
rect 33613 17975 33625 18009
rect 33567 17941 33625 17975
rect 33567 17907 33579 17941
rect 33613 17907 33625 17941
rect 33567 17873 33625 17907
rect 33567 17839 33579 17873
rect 33613 17839 33625 17873
rect 33567 17805 33625 17839
rect 33567 17771 33579 17805
rect 33613 17771 33625 17805
rect 33567 17737 33625 17771
rect 33567 17703 33579 17737
rect 33613 17703 33625 17737
rect 33567 17669 33625 17703
rect 33567 17635 33579 17669
rect 33613 17635 33625 17669
rect 33567 17601 33625 17635
rect 33567 17567 33579 17601
rect 33613 17567 33625 17601
rect 33567 17533 33625 17567
rect 33567 17499 33579 17533
rect 33613 17499 33625 17533
rect 33567 17465 33625 17499
rect 33567 17431 33579 17465
rect 33613 17431 33625 17465
rect 33567 17397 33625 17431
rect 33567 17363 33579 17397
rect 33613 17363 33625 17397
rect 33567 17347 33625 17363
rect 34025 18621 34083 18637
rect 34025 18587 34037 18621
rect 34071 18587 34083 18621
rect 34025 18553 34083 18587
rect 34025 18519 34037 18553
rect 34071 18519 34083 18553
rect 34025 18485 34083 18519
rect 34025 18451 34037 18485
rect 34071 18451 34083 18485
rect 34025 18417 34083 18451
rect 34025 18383 34037 18417
rect 34071 18383 34083 18417
rect 34025 18349 34083 18383
rect 34025 18315 34037 18349
rect 34071 18315 34083 18349
rect 34025 18281 34083 18315
rect 34025 18247 34037 18281
rect 34071 18247 34083 18281
rect 34025 18213 34083 18247
rect 34025 18179 34037 18213
rect 34071 18179 34083 18213
rect 34025 18145 34083 18179
rect 34025 18111 34037 18145
rect 34071 18111 34083 18145
rect 34025 18077 34083 18111
rect 34025 18043 34037 18077
rect 34071 18043 34083 18077
rect 34025 18009 34083 18043
rect 34025 17975 34037 18009
rect 34071 17975 34083 18009
rect 34025 17941 34083 17975
rect 34025 17907 34037 17941
rect 34071 17907 34083 17941
rect 34025 17873 34083 17907
rect 34025 17839 34037 17873
rect 34071 17839 34083 17873
rect 34025 17805 34083 17839
rect 34025 17771 34037 17805
rect 34071 17771 34083 17805
rect 34025 17737 34083 17771
rect 34025 17703 34037 17737
rect 34071 17703 34083 17737
rect 34025 17669 34083 17703
rect 34025 17635 34037 17669
rect 34071 17635 34083 17669
rect 34025 17601 34083 17635
rect 34025 17567 34037 17601
rect 34071 17567 34083 17601
rect 34025 17533 34083 17567
rect 34025 17499 34037 17533
rect 34071 17499 34083 17533
rect 34025 17465 34083 17499
rect 34025 17431 34037 17465
rect 34071 17431 34083 17465
rect 34025 17397 34083 17431
rect 34025 17363 34037 17397
rect 34071 17363 34083 17397
rect 34025 17347 34083 17363
rect 34483 18621 34541 18637
rect 34483 18587 34495 18621
rect 34529 18587 34541 18621
rect 34483 18553 34541 18587
rect 34483 18519 34495 18553
rect 34529 18519 34541 18553
rect 34483 18485 34541 18519
rect 34483 18451 34495 18485
rect 34529 18451 34541 18485
rect 34483 18417 34541 18451
rect 34483 18383 34495 18417
rect 34529 18383 34541 18417
rect 34483 18349 34541 18383
rect 34483 18315 34495 18349
rect 34529 18315 34541 18349
rect 34483 18281 34541 18315
rect 34483 18247 34495 18281
rect 34529 18247 34541 18281
rect 34483 18213 34541 18247
rect 34483 18179 34495 18213
rect 34529 18179 34541 18213
rect 34483 18145 34541 18179
rect 34483 18111 34495 18145
rect 34529 18111 34541 18145
rect 34483 18077 34541 18111
rect 34483 18043 34495 18077
rect 34529 18043 34541 18077
rect 34483 18009 34541 18043
rect 34483 17975 34495 18009
rect 34529 17975 34541 18009
rect 34483 17941 34541 17975
rect 34483 17907 34495 17941
rect 34529 17907 34541 17941
rect 34483 17873 34541 17907
rect 34483 17839 34495 17873
rect 34529 17839 34541 17873
rect 34483 17805 34541 17839
rect 34483 17771 34495 17805
rect 34529 17771 34541 17805
rect 34483 17737 34541 17771
rect 34483 17703 34495 17737
rect 34529 17703 34541 17737
rect 34483 17669 34541 17703
rect 34483 17635 34495 17669
rect 34529 17635 34541 17669
rect 34483 17601 34541 17635
rect 34483 17567 34495 17601
rect 34529 17567 34541 17601
rect 34483 17533 34541 17567
rect 34483 17499 34495 17533
rect 34529 17499 34541 17533
rect 34483 17465 34541 17499
rect 34483 17431 34495 17465
rect 34529 17431 34541 17465
rect 34483 17397 34541 17431
rect 34483 17363 34495 17397
rect 34529 17363 34541 17397
rect 34483 17347 34541 17363
rect 34941 18621 34999 18637
rect 34941 18587 34953 18621
rect 34987 18587 34999 18621
rect 34941 18553 34999 18587
rect 34941 18519 34953 18553
rect 34987 18519 34999 18553
rect 34941 18485 34999 18519
rect 34941 18451 34953 18485
rect 34987 18451 34999 18485
rect 34941 18417 34999 18451
rect 34941 18383 34953 18417
rect 34987 18383 34999 18417
rect 34941 18349 34999 18383
rect 34941 18315 34953 18349
rect 34987 18315 34999 18349
rect 34941 18281 34999 18315
rect 34941 18247 34953 18281
rect 34987 18247 34999 18281
rect 34941 18213 34999 18247
rect 34941 18179 34953 18213
rect 34987 18179 34999 18213
rect 34941 18145 34999 18179
rect 34941 18111 34953 18145
rect 34987 18111 34999 18145
rect 34941 18077 34999 18111
rect 34941 18043 34953 18077
rect 34987 18043 34999 18077
rect 34941 18009 34999 18043
rect 34941 17975 34953 18009
rect 34987 17975 34999 18009
rect 34941 17941 34999 17975
rect 34941 17907 34953 17941
rect 34987 17907 34999 17941
rect 34941 17873 34999 17907
rect 34941 17839 34953 17873
rect 34987 17839 34999 17873
rect 34941 17805 34999 17839
rect 34941 17771 34953 17805
rect 34987 17771 34999 17805
rect 34941 17737 34999 17771
rect 34941 17703 34953 17737
rect 34987 17703 34999 17737
rect 34941 17669 34999 17703
rect 34941 17635 34953 17669
rect 34987 17635 34999 17669
rect 34941 17601 34999 17635
rect 34941 17567 34953 17601
rect 34987 17567 34999 17601
rect 34941 17533 34999 17567
rect 34941 17499 34953 17533
rect 34987 17499 34999 17533
rect 34941 17465 34999 17499
rect 34941 17431 34953 17465
rect 34987 17431 34999 17465
rect 34941 17397 34999 17431
rect 34941 17363 34953 17397
rect 34987 17363 34999 17397
rect 34941 17347 34999 17363
rect 35399 18621 35457 18637
rect 35399 18587 35411 18621
rect 35445 18587 35457 18621
rect 35399 18553 35457 18587
rect 35399 18519 35411 18553
rect 35445 18519 35457 18553
rect 35399 18485 35457 18519
rect 35399 18451 35411 18485
rect 35445 18451 35457 18485
rect 35399 18417 35457 18451
rect 35399 18383 35411 18417
rect 35445 18383 35457 18417
rect 35399 18349 35457 18383
rect 35399 18315 35411 18349
rect 35445 18315 35457 18349
rect 35399 18281 35457 18315
rect 35399 18247 35411 18281
rect 35445 18247 35457 18281
rect 35399 18213 35457 18247
rect 35399 18179 35411 18213
rect 35445 18179 35457 18213
rect 35399 18145 35457 18179
rect 35399 18111 35411 18145
rect 35445 18111 35457 18145
rect 35399 18077 35457 18111
rect 35399 18043 35411 18077
rect 35445 18043 35457 18077
rect 35399 18009 35457 18043
rect 35399 17975 35411 18009
rect 35445 17975 35457 18009
rect 35399 17941 35457 17975
rect 35399 17907 35411 17941
rect 35445 17907 35457 17941
rect 35399 17873 35457 17907
rect 35399 17839 35411 17873
rect 35445 17839 35457 17873
rect 35399 17805 35457 17839
rect 35399 17771 35411 17805
rect 35445 17771 35457 17805
rect 35399 17737 35457 17771
rect 35399 17703 35411 17737
rect 35445 17703 35457 17737
rect 35399 17669 35457 17703
rect 35399 17635 35411 17669
rect 35445 17635 35457 17669
rect 35399 17601 35457 17635
rect 35399 17567 35411 17601
rect 35445 17567 35457 17601
rect 35399 17533 35457 17567
rect 35399 17499 35411 17533
rect 35445 17499 35457 17533
rect 35399 17465 35457 17499
rect 35399 17431 35411 17465
rect 35445 17431 35457 17465
rect 35399 17397 35457 17431
rect 35399 17363 35411 17397
rect 35445 17363 35457 17397
rect 35399 17347 35457 17363
rect 35857 18621 35915 18637
rect 35857 18587 35869 18621
rect 35903 18587 35915 18621
rect 35857 18553 35915 18587
rect 35857 18519 35869 18553
rect 35903 18519 35915 18553
rect 35857 18485 35915 18519
rect 35857 18451 35869 18485
rect 35903 18451 35915 18485
rect 35857 18417 35915 18451
rect 35857 18383 35869 18417
rect 35903 18383 35915 18417
rect 35857 18349 35915 18383
rect 35857 18315 35869 18349
rect 35903 18315 35915 18349
rect 35857 18281 35915 18315
rect 35857 18247 35869 18281
rect 35903 18247 35915 18281
rect 35857 18213 35915 18247
rect 35857 18179 35869 18213
rect 35903 18179 35915 18213
rect 35857 18145 35915 18179
rect 35857 18111 35869 18145
rect 35903 18111 35915 18145
rect 35857 18077 35915 18111
rect 35857 18043 35869 18077
rect 35903 18043 35915 18077
rect 35857 18009 35915 18043
rect 35857 17975 35869 18009
rect 35903 17975 35915 18009
rect 35857 17941 35915 17975
rect 35857 17907 35869 17941
rect 35903 17907 35915 17941
rect 35857 17873 35915 17907
rect 35857 17839 35869 17873
rect 35903 17839 35915 17873
rect 35857 17805 35915 17839
rect 35857 17771 35869 17805
rect 35903 17771 35915 17805
rect 35857 17737 35915 17771
rect 35857 17703 35869 17737
rect 35903 17703 35915 17737
rect 35857 17669 35915 17703
rect 35857 17635 35869 17669
rect 35903 17635 35915 17669
rect 35857 17601 35915 17635
rect 35857 17567 35869 17601
rect 35903 17567 35915 17601
rect 35857 17533 35915 17567
rect 35857 17499 35869 17533
rect 35903 17499 35915 17533
rect 35857 17465 35915 17499
rect 35857 17431 35869 17465
rect 35903 17431 35915 17465
rect 35857 17397 35915 17431
rect 35857 17363 35869 17397
rect 35903 17363 35915 17397
rect 35857 17347 35915 17363
rect 36315 18621 36373 18637
rect 36315 18587 36327 18621
rect 36361 18587 36373 18621
rect 36315 18553 36373 18587
rect 36315 18519 36327 18553
rect 36361 18519 36373 18553
rect 36315 18485 36373 18519
rect 36315 18451 36327 18485
rect 36361 18451 36373 18485
rect 36315 18417 36373 18451
rect 36315 18383 36327 18417
rect 36361 18383 36373 18417
rect 36315 18349 36373 18383
rect 36315 18315 36327 18349
rect 36361 18315 36373 18349
rect 36315 18281 36373 18315
rect 36315 18247 36327 18281
rect 36361 18247 36373 18281
rect 36315 18213 36373 18247
rect 36315 18179 36327 18213
rect 36361 18179 36373 18213
rect 36315 18145 36373 18179
rect 36315 18111 36327 18145
rect 36361 18111 36373 18145
rect 36315 18077 36373 18111
rect 36315 18043 36327 18077
rect 36361 18043 36373 18077
rect 36315 18009 36373 18043
rect 36315 17975 36327 18009
rect 36361 17975 36373 18009
rect 36315 17941 36373 17975
rect 36315 17907 36327 17941
rect 36361 17907 36373 17941
rect 36315 17873 36373 17907
rect 36315 17839 36327 17873
rect 36361 17839 36373 17873
rect 36315 17805 36373 17839
rect 36315 17771 36327 17805
rect 36361 17771 36373 17805
rect 36315 17737 36373 17771
rect 36315 17703 36327 17737
rect 36361 17703 36373 17737
rect 36315 17669 36373 17703
rect 36315 17635 36327 17669
rect 36361 17635 36373 17669
rect 36315 17601 36373 17635
rect 36315 17567 36327 17601
rect 36361 17567 36373 17601
rect 36315 17533 36373 17567
rect 36315 17499 36327 17533
rect 36361 17499 36373 17533
rect 36315 17465 36373 17499
rect 36315 17431 36327 17465
rect 36361 17431 36373 17465
rect 36315 17397 36373 17431
rect 36315 17363 36327 17397
rect 36361 17363 36373 17397
rect 36315 17347 36373 17363
rect 36773 18621 36831 18637
rect 36773 18587 36785 18621
rect 36819 18587 36831 18621
rect 36773 18553 36831 18587
rect 36773 18519 36785 18553
rect 36819 18519 36831 18553
rect 36773 18485 36831 18519
rect 36773 18451 36785 18485
rect 36819 18451 36831 18485
rect 36773 18417 36831 18451
rect 36773 18383 36785 18417
rect 36819 18383 36831 18417
rect 36773 18349 36831 18383
rect 36773 18315 36785 18349
rect 36819 18315 36831 18349
rect 36773 18281 36831 18315
rect 36773 18247 36785 18281
rect 36819 18247 36831 18281
rect 36773 18213 36831 18247
rect 36773 18179 36785 18213
rect 36819 18179 36831 18213
rect 36773 18145 36831 18179
rect 36773 18111 36785 18145
rect 36819 18111 36831 18145
rect 36773 18077 36831 18111
rect 36773 18043 36785 18077
rect 36819 18043 36831 18077
rect 36773 18009 36831 18043
rect 36773 17975 36785 18009
rect 36819 17975 36831 18009
rect 36773 17941 36831 17975
rect 36773 17907 36785 17941
rect 36819 17907 36831 17941
rect 36773 17873 36831 17907
rect 36773 17839 36785 17873
rect 36819 17839 36831 17873
rect 36773 17805 36831 17839
rect 36773 17771 36785 17805
rect 36819 17771 36831 17805
rect 36773 17737 36831 17771
rect 36773 17703 36785 17737
rect 36819 17703 36831 17737
rect 36773 17669 36831 17703
rect 36773 17635 36785 17669
rect 36819 17635 36831 17669
rect 36773 17601 36831 17635
rect 36773 17567 36785 17601
rect 36819 17567 36831 17601
rect 36773 17533 36831 17567
rect 36773 17499 36785 17533
rect 36819 17499 36831 17533
rect 36773 17465 36831 17499
rect 36773 17431 36785 17465
rect 36819 17431 36831 17465
rect 36773 17397 36831 17431
rect 36773 17363 36785 17397
rect 36819 17363 36831 17397
rect 36773 17347 36831 17363
rect 37231 18621 37289 18637
rect 37231 18587 37243 18621
rect 37277 18587 37289 18621
rect 37231 18553 37289 18587
rect 37231 18519 37243 18553
rect 37277 18519 37289 18553
rect 37231 18485 37289 18519
rect 37231 18451 37243 18485
rect 37277 18451 37289 18485
rect 37231 18417 37289 18451
rect 37231 18383 37243 18417
rect 37277 18383 37289 18417
rect 37231 18349 37289 18383
rect 37231 18315 37243 18349
rect 37277 18315 37289 18349
rect 37231 18281 37289 18315
rect 37231 18247 37243 18281
rect 37277 18247 37289 18281
rect 37231 18213 37289 18247
rect 37231 18179 37243 18213
rect 37277 18179 37289 18213
rect 37231 18145 37289 18179
rect 37231 18111 37243 18145
rect 37277 18111 37289 18145
rect 37231 18077 37289 18111
rect 37231 18043 37243 18077
rect 37277 18043 37289 18077
rect 37231 18009 37289 18043
rect 37231 17975 37243 18009
rect 37277 17975 37289 18009
rect 37231 17941 37289 17975
rect 37231 17907 37243 17941
rect 37277 17907 37289 17941
rect 37231 17873 37289 17907
rect 37231 17839 37243 17873
rect 37277 17839 37289 17873
rect 37231 17805 37289 17839
rect 37231 17771 37243 17805
rect 37277 17771 37289 17805
rect 37231 17737 37289 17771
rect 37231 17703 37243 17737
rect 37277 17703 37289 17737
rect 37231 17669 37289 17703
rect 37231 17635 37243 17669
rect 37277 17635 37289 17669
rect 37231 17601 37289 17635
rect 37231 17567 37243 17601
rect 37277 17567 37289 17601
rect 37231 17533 37289 17567
rect 37231 17499 37243 17533
rect 37277 17499 37289 17533
rect 37231 17465 37289 17499
rect 37231 17431 37243 17465
rect 37277 17431 37289 17465
rect 37231 17397 37289 17431
rect 37231 17363 37243 17397
rect 37277 17363 37289 17397
rect 37231 17347 37289 17363
rect 37689 18621 37747 18637
rect 37689 18587 37701 18621
rect 37735 18587 37747 18621
rect 37689 18553 37747 18587
rect 37689 18519 37701 18553
rect 37735 18519 37747 18553
rect 37689 18485 37747 18519
rect 37689 18451 37701 18485
rect 37735 18451 37747 18485
rect 37689 18417 37747 18451
rect 37689 18383 37701 18417
rect 37735 18383 37747 18417
rect 37689 18349 37747 18383
rect 37689 18315 37701 18349
rect 37735 18315 37747 18349
rect 37689 18281 37747 18315
rect 37689 18247 37701 18281
rect 37735 18247 37747 18281
rect 37689 18213 37747 18247
rect 37689 18179 37701 18213
rect 37735 18179 37747 18213
rect 37689 18145 37747 18179
rect 37689 18111 37701 18145
rect 37735 18111 37747 18145
rect 37689 18077 37747 18111
rect 37689 18043 37701 18077
rect 37735 18043 37747 18077
rect 37689 18009 37747 18043
rect 37689 17975 37701 18009
rect 37735 17975 37747 18009
rect 37689 17941 37747 17975
rect 37689 17907 37701 17941
rect 37735 17907 37747 17941
rect 37689 17873 37747 17907
rect 37689 17839 37701 17873
rect 37735 17839 37747 17873
rect 37689 17805 37747 17839
rect 37689 17771 37701 17805
rect 37735 17771 37747 17805
rect 37689 17737 37747 17771
rect 37689 17703 37701 17737
rect 37735 17703 37747 17737
rect 37689 17669 37747 17703
rect 37689 17635 37701 17669
rect 37735 17635 37747 17669
rect 37689 17601 37747 17635
rect 37689 17567 37701 17601
rect 37735 17567 37747 17601
rect 37689 17533 37747 17567
rect 37689 17499 37701 17533
rect 37735 17499 37747 17533
rect 37689 17465 37747 17499
rect 37689 17431 37701 17465
rect 37735 17431 37747 17465
rect 37689 17397 37747 17431
rect 37689 17363 37701 17397
rect 37735 17363 37747 17397
rect 37689 17347 37747 17363
rect 38147 18621 38205 18637
rect 38147 18587 38159 18621
rect 38193 18587 38205 18621
rect 38147 18553 38205 18587
rect 38147 18519 38159 18553
rect 38193 18519 38205 18553
rect 38147 18485 38205 18519
rect 38147 18451 38159 18485
rect 38193 18451 38205 18485
rect 38147 18417 38205 18451
rect 38147 18383 38159 18417
rect 38193 18383 38205 18417
rect 38147 18349 38205 18383
rect 38147 18315 38159 18349
rect 38193 18315 38205 18349
rect 38147 18281 38205 18315
rect 38147 18247 38159 18281
rect 38193 18247 38205 18281
rect 38147 18213 38205 18247
rect 38147 18179 38159 18213
rect 38193 18179 38205 18213
rect 38147 18145 38205 18179
rect 38147 18111 38159 18145
rect 38193 18111 38205 18145
rect 38147 18077 38205 18111
rect 38147 18043 38159 18077
rect 38193 18043 38205 18077
rect 38147 18009 38205 18043
rect 38147 17975 38159 18009
rect 38193 17975 38205 18009
rect 38147 17941 38205 17975
rect 38147 17907 38159 17941
rect 38193 17907 38205 17941
rect 38147 17873 38205 17907
rect 38147 17839 38159 17873
rect 38193 17839 38205 17873
rect 38147 17805 38205 17839
rect 38147 17771 38159 17805
rect 38193 17771 38205 17805
rect 38147 17737 38205 17771
rect 38147 17703 38159 17737
rect 38193 17703 38205 17737
rect 38147 17669 38205 17703
rect 38147 17635 38159 17669
rect 38193 17635 38205 17669
rect 38147 17601 38205 17635
rect 38147 17567 38159 17601
rect 38193 17567 38205 17601
rect 38147 17533 38205 17567
rect 38147 17499 38159 17533
rect 38193 17499 38205 17533
rect 38147 17465 38205 17499
rect 38147 17431 38159 17465
rect 38193 17431 38205 17465
rect 38147 17397 38205 17431
rect 38147 17363 38159 17397
rect 38193 17363 38205 17397
rect 38147 17347 38205 17363
rect 38605 18621 38663 18637
rect 38605 18587 38617 18621
rect 38651 18587 38663 18621
rect 38605 18553 38663 18587
rect 38605 18519 38617 18553
rect 38651 18519 38663 18553
rect 38605 18485 38663 18519
rect 38605 18451 38617 18485
rect 38651 18451 38663 18485
rect 38605 18417 38663 18451
rect 38605 18383 38617 18417
rect 38651 18383 38663 18417
rect 38605 18349 38663 18383
rect 38605 18315 38617 18349
rect 38651 18315 38663 18349
rect 38605 18281 38663 18315
rect 38605 18247 38617 18281
rect 38651 18247 38663 18281
rect 38605 18213 38663 18247
rect 38605 18179 38617 18213
rect 38651 18179 38663 18213
rect 38605 18145 38663 18179
rect 38605 18111 38617 18145
rect 38651 18111 38663 18145
rect 38605 18077 38663 18111
rect 38605 18043 38617 18077
rect 38651 18043 38663 18077
rect 38605 18009 38663 18043
rect 38605 17975 38617 18009
rect 38651 17975 38663 18009
rect 38605 17941 38663 17975
rect 38605 17907 38617 17941
rect 38651 17907 38663 17941
rect 38605 17873 38663 17907
rect 38605 17839 38617 17873
rect 38651 17839 38663 17873
rect 38605 17805 38663 17839
rect 38605 17771 38617 17805
rect 38651 17771 38663 17805
rect 38605 17737 38663 17771
rect 38605 17703 38617 17737
rect 38651 17703 38663 17737
rect 38605 17669 38663 17703
rect 38605 17635 38617 17669
rect 38651 17635 38663 17669
rect 38605 17601 38663 17635
rect 38605 17567 38617 17601
rect 38651 17567 38663 17601
rect 38605 17533 38663 17567
rect 38605 17499 38617 17533
rect 38651 17499 38663 17533
rect 38605 17465 38663 17499
rect 38605 17431 38617 17465
rect 38651 17431 38663 17465
rect 38605 17397 38663 17431
rect 38605 17363 38617 17397
rect 38651 17363 38663 17397
rect 38605 17347 38663 17363
rect 39063 18621 39121 18637
rect 39063 18587 39075 18621
rect 39109 18587 39121 18621
rect 39063 18553 39121 18587
rect 39063 18519 39075 18553
rect 39109 18519 39121 18553
rect 39063 18485 39121 18519
rect 39063 18451 39075 18485
rect 39109 18451 39121 18485
rect 39063 18417 39121 18451
rect 39063 18383 39075 18417
rect 39109 18383 39121 18417
rect 39063 18349 39121 18383
rect 39063 18315 39075 18349
rect 39109 18315 39121 18349
rect 39063 18281 39121 18315
rect 39063 18247 39075 18281
rect 39109 18247 39121 18281
rect 39063 18213 39121 18247
rect 39063 18179 39075 18213
rect 39109 18179 39121 18213
rect 39063 18145 39121 18179
rect 39063 18111 39075 18145
rect 39109 18111 39121 18145
rect 39063 18077 39121 18111
rect 39063 18043 39075 18077
rect 39109 18043 39121 18077
rect 39063 18009 39121 18043
rect 39063 17975 39075 18009
rect 39109 17975 39121 18009
rect 39063 17941 39121 17975
rect 39063 17907 39075 17941
rect 39109 17907 39121 17941
rect 39063 17873 39121 17907
rect 39063 17839 39075 17873
rect 39109 17839 39121 17873
rect 39063 17805 39121 17839
rect 39063 17771 39075 17805
rect 39109 17771 39121 17805
rect 39063 17737 39121 17771
rect 39063 17703 39075 17737
rect 39109 17703 39121 17737
rect 39063 17669 39121 17703
rect 39063 17635 39075 17669
rect 39109 17635 39121 17669
rect 39063 17601 39121 17635
rect 39063 17567 39075 17601
rect 39109 17567 39121 17601
rect 39063 17533 39121 17567
rect 39063 17499 39075 17533
rect 39109 17499 39121 17533
rect 39063 17465 39121 17499
rect 39063 17431 39075 17465
rect 39109 17431 39121 17465
rect 39063 17397 39121 17431
rect 39063 17363 39075 17397
rect 39109 17363 39121 17397
rect 39063 17347 39121 17363
rect 39521 18621 39579 18637
rect 39521 18587 39533 18621
rect 39567 18587 39579 18621
rect 39521 18553 39579 18587
rect 39521 18519 39533 18553
rect 39567 18519 39579 18553
rect 39521 18485 39579 18519
rect 39521 18451 39533 18485
rect 39567 18451 39579 18485
rect 39521 18417 39579 18451
rect 39521 18383 39533 18417
rect 39567 18383 39579 18417
rect 39521 18349 39579 18383
rect 39521 18315 39533 18349
rect 39567 18315 39579 18349
rect 39521 18281 39579 18315
rect 39521 18247 39533 18281
rect 39567 18247 39579 18281
rect 39521 18213 39579 18247
rect 39521 18179 39533 18213
rect 39567 18179 39579 18213
rect 39521 18145 39579 18179
rect 39521 18111 39533 18145
rect 39567 18111 39579 18145
rect 39521 18077 39579 18111
rect 39521 18043 39533 18077
rect 39567 18043 39579 18077
rect 39521 18009 39579 18043
rect 39521 17975 39533 18009
rect 39567 17975 39579 18009
rect 39521 17941 39579 17975
rect 39521 17907 39533 17941
rect 39567 17907 39579 17941
rect 39521 17873 39579 17907
rect 39521 17839 39533 17873
rect 39567 17839 39579 17873
rect 39521 17805 39579 17839
rect 39521 17771 39533 17805
rect 39567 17771 39579 17805
rect 39521 17737 39579 17771
rect 39521 17703 39533 17737
rect 39567 17703 39579 17737
rect 39521 17669 39579 17703
rect 39521 17635 39533 17669
rect 39567 17635 39579 17669
rect 39521 17601 39579 17635
rect 39521 17567 39533 17601
rect 39567 17567 39579 17601
rect 39521 17533 39579 17567
rect 39521 17499 39533 17533
rect 39567 17499 39579 17533
rect 39521 17465 39579 17499
rect 39521 17431 39533 17465
rect 39567 17431 39579 17465
rect 39521 17397 39579 17431
rect 39521 17363 39533 17397
rect 39567 17363 39579 17397
rect 39521 17347 39579 17363
rect 39979 18621 40037 18637
rect 39979 18587 39991 18621
rect 40025 18587 40037 18621
rect 39979 18553 40037 18587
rect 39979 18519 39991 18553
rect 40025 18519 40037 18553
rect 39979 18485 40037 18519
rect 39979 18451 39991 18485
rect 40025 18451 40037 18485
rect 39979 18417 40037 18451
rect 39979 18383 39991 18417
rect 40025 18383 40037 18417
rect 39979 18349 40037 18383
rect 39979 18315 39991 18349
rect 40025 18315 40037 18349
rect 39979 18281 40037 18315
rect 39979 18247 39991 18281
rect 40025 18247 40037 18281
rect 39979 18213 40037 18247
rect 39979 18179 39991 18213
rect 40025 18179 40037 18213
rect 39979 18145 40037 18179
rect 39979 18111 39991 18145
rect 40025 18111 40037 18145
rect 39979 18077 40037 18111
rect 39979 18043 39991 18077
rect 40025 18043 40037 18077
rect 39979 18009 40037 18043
rect 39979 17975 39991 18009
rect 40025 17975 40037 18009
rect 39979 17941 40037 17975
rect 39979 17907 39991 17941
rect 40025 17907 40037 17941
rect 39979 17873 40037 17907
rect 39979 17839 39991 17873
rect 40025 17839 40037 17873
rect 39979 17805 40037 17839
rect 39979 17771 39991 17805
rect 40025 17771 40037 17805
rect 39979 17737 40037 17771
rect 39979 17703 39991 17737
rect 40025 17703 40037 17737
rect 39979 17669 40037 17703
rect 39979 17635 39991 17669
rect 40025 17635 40037 17669
rect 39979 17601 40037 17635
rect 39979 17567 39991 17601
rect 40025 17567 40037 17601
rect 39979 17533 40037 17567
rect 39979 17499 39991 17533
rect 40025 17499 40037 17533
rect 39979 17465 40037 17499
rect 39979 17431 39991 17465
rect 40025 17431 40037 17465
rect 39979 17397 40037 17431
rect 39979 17363 39991 17397
rect 40025 17363 40037 17397
rect 39979 17347 40037 17363
rect 40437 18621 40495 18637
rect 40437 18587 40449 18621
rect 40483 18587 40495 18621
rect 40437 18553 40495 18587
rect 40437 18519 40449 18553
rect 40483 18519 40495 18553
rect 40437 18485 40495 18519
rect 40437 18451 40449 18485
rect 40483 18451 40495 18485
rect 40437 18417 40495 18451
rect 40437 18383 40449 18417
rect 40483 18383 40495 18417
rect 40437 18349 40495 18383
rect 40437 18315 40449 18349
rect 40483 18315 40495 18349
rect 40437 18281 40495 18315
rect 40437 18247 40449 18281
rect 40483 18247 40495 18281
rect 40437 18213 40495 18247
rect 40437 18179 40449 18213
rect 40483 18179 40495 18213
rect 40437 18145 40495 18179
rect 40437 18111 40449 18145
rect 40483 18111 40495 18145
rect 40437 18077 40495 18111
rect 40437 18043 40449 18077
rect 40483 18043 40495 18077
rect 40437 18009 40495 18043
rect 40437 17975 40449 18009
rect 40483 17975 40495 18009
rect 40437 17941 40495 17975
rect 40437 17907 40449 17941
rect 40483 17907 40495 17941
rect 40437 17873 40495 17907
rect 40437 17839 40449 17873
rect 40483 17839 40495 17873
rect 40437 17805 40495 17839
rect 40437 17771 40449 17805
rect 40483 17771 40495 17805
rect 40437 17737 40495 17771
rect 40437 17703 40449 17737
rect 40483 17703 40495 17737
rect 40437 17669 40495 17703
rect 40437 17635 40449 17669
rect 40483 17635 40495 17669
rect 40437 17601 40495 17635
rect 40437 17567 40449 17601
rect 40483 17567 40495 17601
rect 40437 17533 40495 17567
rect 40437 17499 40449 17533
rect 40483 17499 40495 17533
rect 40437 17465 40495 17499
rect 40437 17431 40449 17465
rect 40483 17431 40495 17465
rect 40437 17397 40495 17431
rect 40437 17363 40449 17397
rect 40483 17363 40495 17397
rect 40437 17347 40495 17363
rect 40895 18621 40953 18637
rect 40895 18587 40907 18621
rect 40941 18587 40953 18621
rect 40895 18553 40953 18587
rect 40895 18519 40907 18553
rect 40941 18519 40953 18553
rect 40895 18485 40953 18519
rect 40895 18451 40907 18485
rect 40941 18451 40953 18485
rect 40895 18417 40953 18451
rect 40895 18383 40907 18417
rect 40941 18383 40953 18417
rect 40895 18349 40953 18383
rect 40895 18315 40907 18349
rect 40941 18315 40953 18349
rect 40895 18281 40953 18315
rect 40895 18247 40907 18281
rect 40941 18247 40953 18281
rect 40895 18213 40953 18247
rect 40895 18179 40907 18213
rect 40941 18179 40953 18213
rect 40895 18145 40953 18179
rect 40895 18111 40907 18145
rect 40941 18111 40953 18145
rect 40895 18077 40953 18111
rect 40895 18043 40907 18077
rect 40941 18043 40953 18077
rect 40895 18009 40953 18043
rect 40895 17975 40907 18009
rect 40941 17975 40953 18009
rect 40895 17941 40953 17975
rect 40895 17907 40907 17941
rect 40941 17907 40953 17941
rect 40895 17873 40953 17907
rect 40895 17839 40907 17873
rect 40941 17839 40953 17873
rect 40895 17805 40953 17839
rect 40895 17771 40907 17805
rect 40941 17771 40953 17805
rect 40895 17737 40953 17771
rect 40895 17703 40907 17737
rect 40941 17703 40953 17737
rect 40895 17669 40953 17703
rect 40895 17635 40907 17669
rect 40941 17635 40953 17669
rect 40895 17601 40953 17635
rect 40895 17567 40907 17601
rect 40941 17567 40953 17601
rect 40895 17533 40953 17567
rect 40895 17499 40907 17533
rect 40941 17499 40953 17533
rect 40895 17465 40953 17499
rect 40895 17431 40907 17465
rect 40941 17431 40953 17465
rect 40895 17397 40953 17431
rect 40895 17363 40907 17397
rect 40941 17363 40953 17397
rect 40895 17347 40953 17363
rect 41353 18621 41411 18637
rect 41353 18587 41365 18621
rect 41399 18587 41411 18621
rect 41353 18553 41411 18587
rect 41353 18519 41365 18553
rect 41399 18519 41411 18553
rect 41353 18485 41411 18519
rect 41353 18451 41365 18485
rect 41399 18451 41411 18485
rect 41353 18417 41411 18451
rect 41353 18383 41365 18417
rect 41399 18383 41411 18417
rect 41353 18349 41411 18383
rect 41353 18315 41365 18349
rect 41399 18315 41411 18349
rect 41353 18281 41411 18315
rect 41353 18247 41365 18281
rect 41399 18247 41411 18281
rect 41353 18213 41411 18247
rect 41353 18179 41365 18213
rect 41399 18179 41411 18213
rect 41353 18145 41411 18179
rect 41353 18111 41365 18145
rect 41399 18111 41411 18145
rect 41353 18077 41411 18111
rect 41353 18043 41365 18077
rect 41399 18043 41411 18077
rect 41353 18009 41411 18043
rect 41353 17975 41365 18009
rect 41399 17975 41411 18009
rect 41353 17941 41411 17975
rect 41353 17907 41365 17941
rect 41399 17907 41411 17941
rect 41353 17873 41411 17907
rect 41353 17839 41365 17873
rect 41399 17839 41411 17873
rect 41353 17805 41411 17839
rect 41353 17771 41365 17805
rect 41399 17771 41411 17805
rect 41353 17737 41411 17771
rect 41353 17703 41365 17737
rect 41399 17703 41411 17737
rect 41353 17669 41411 17703
rect 41353 17635 41365 17669
rect 41399 17635 41411 17669
rect 41353 17601 41411 17635
rect 41353 17567 41365 17601
rect 41399 17567 41411 17601
rect 41353 17533 41411 17567
rect 41353 17499 41365 17533
rect 41399 17499 41411 17533
rect 41353 17465 41411 17499
rect 41353 17431 41365 17465
rect 41399 17431 41411 17465
rect 41353 17397 41411 17431
rect 41353 17363 41365 17397
rect 41399 17363 41411 17397
rect 41353 17347 41411 17363
rect 41811 18621 41869 18637
rect 41811 18587 41823 18621
rect 41857 18587 41869 18621
rect 41811 18553 41869 18587
rect 41811 18519 41823 18553
rect 41857 18519 41869 18553
rect 41811 18485 41869 18519
rect 41811 18451 41823 18485
rect 41857 18451 41869 18485
rect 41811 18417 41869 18451
rect 41811 18383 41823 18417
rect 41857 18383 41869 18417
rect 41811 18349 41869 18383
rect 41811 18315 41823 18349
rect 41857 18315 41869 18349
rect 41811 18281 41869 18315
rect 41811 18247 41823 18281
rect 41857 18247 41869 18281
rect 41811 18213 41869 18247
rect 41811 18179 41823 18213
rect 41857 18179 41869 18213
rect 41811 18145 41869 18179
rect 41811 18111 41823 18145
rect 41857 18111 41869 18145
rect 41811 18077 41869 18111
rect 41811 18043 41823 18077
rect 41857 18043 41869 18077
rect 41811 18009 41869 18043
rect 41811 17975 41823 18009
rect 41857 17975 41869 18009
rect 41811 17941 41869 17975
rect 41811 17907 41823 17941
rect 41857 17907 41869 17941
rect 41811 17873 41869 17907
rect 41811 17839 41823 17873
rect 41857 17839 41869 17873
rect 41811 17805 41869 17839
rect 41811 17771 41823 17805
rect 41857 17771 41869 17805
rect 41811 17737 41869 17771
rect 41811 17703 41823 17737
rect 41857 17703 41869 17737
rect 41811 17669 41869 17703
rect 41811 17635 41823 17669
rect 41857 17635 41869 17669
rect 41811 17601 41869 17635
rect 41811 17567 41823 17601
rect 41857 17567 41869 17601
rect 41811 17533 41869 17567
rect 41811 17499 41823 17533
rect 41857 17499 41869 17533
rect 41811 17465 41869 17499
rect 41811 17431 41823 17465
rect 41857 17431 41869 17465
rect 41811 17397 41869 17431
rect 41811 17363 41823 17397
rect 41857 17363 41869 17397
rect 41811 17347 41869 17363
rect 42269 18621 42327 18637
rect 42269 18587 42281 18621
rect 42315 18587 42327 18621
rect 42269 18553 42327 18587
rect 42269 18519 42281 18553
rect 42315 18519 42327 18553
rect 42269 18485 42327 18519
rect 42269 18451 42281 18485
rect 42315 18451 42327 18485
rect 42269 18417 42327 18451
rect 42269 18383 42281 18417
rect 42315 18383 42327 18417
rect 42269 18349 42327 18383
rect 42269 18315 42281 18349
rect 42315 18315 42327 18349
rect 42269 18281 42327 18315
rect 42269 18247 42281 18281
rect 42315 18247 42327 18281
rect 42269 18213 42327 18247
rect 42269 18179 42281 18213
rect 42315 18179 42327 18213
rect 42269 18145 42327 18179
rect 42269 18111 42281 18145
rect 42315 18111 42327 18145
rect 42269 18077 42327 18111
rect 42269 18043 42281 18077
rect 42315 18043 42327 18077
rect 42269 18009 42327 18043
rect 42269 17975 42281 18009
rect 42315 17975 42327 18009
rect 42269 17941 42327 17975
rect 42269 17907 42281 17941
rect 42315 17907 42327 17941
rect 42269 17873 42327 17907
rect 42269 17839 42281 17873
rect 42315 17839 42327 17873
rect 42269 17805 42327 17839
rect 42269 17771 42281 17805
rect 42315 17771 42327 17805
rect 42269 17737 42327 17771
rect 42269 17703 42281 17737
rect 42315 17703 42327 17737
rect 42269 17669 42327 17703
rect 42269 17635 42281 17669
rect 42315 17635 42327 17669
rect 42269 17601 42327 17635
rect 42269 17567 42281 17601
rect 42315 17567 42327 17601
rect 42269 17533 42327 17567
rect 42269 17499 42281 17533
rect 42315 17499 42327 17533
rect 42269 17465 42327 17499
rect 42269 17431 42281 17465
rect 42315 17431 42327 17465
rect 42269 17397 42327 17431
rect 42269 17363 42281 17397
rect 42315 17363 42327 17397
rect 42269 17347 42327 17363
rect 42727 18621 42785 18637
rect 42727 18587 42739 18621
rect 42773 18587 42785 18621
rect 42727 18553 42785 18587
rect 42727 18519 42739 18553
rect 42773 18519 42785 18553
rect 42727 18485 42785 18519
rect 42727 18451 42739 18485
rect 42773 18451 42785 18485
rect 42727 18417 42785 18451
rect 42727 18383 42739 18417
rect 42773 18383 42785 18417
rect 42727 18349 42785 18383
rect 42727 18315 42739 18349
rect 42773 18315 42785 18349
rect 42727 18281 42785 18315
rect 42727 18247 42739 18281
rect 42773 18247 42785 18281
rect 42727 18213 42785 18247
rect 42727 18179 42739 18213
rect 42773 18179 42785 18213
rect 42727 18145 42785 18179
rect 42727 18111 42739 18145
rect 42773 18111 42785 18145
rect 42727 18077 42785 18111
rect 42727 18043 42739 18077
rect 42773 18043 42785 18077
rect 42727 18009 42785 18043
rect 42727 17975 42739 18009
rect 42773 17975 42785 18009
rect 42727 17941 42785 17975
rect 42727 17907 42739 17941
rect 42773 17907 42785 17941
rect 42727 17873 42785 17907
rect 42727 17839 42739 17873
rect 42773 17839 42785 17873
rect 42727 17805 42785 17839
rect 42727 17771 42739 17805
rect 42773 17771 42785 17805
rect 42727 17737 42785 17771
rect 42727 17703 42739 17737
rect 42773 17703 42785 17737
rect 42727 17669 42785 17703
rect 42727 17635 42739 17669
rect 42773 17635 42785 17669
rect 42727 17601 42785 17635
rect 42727 17567 42739 17601
rect 42773 17567 42785 17601
rect 42727 17533 42785 17567
rect 42727 17499 42739 17533
rect 42773 17499 42785 17533
rect 42727 17465 42785 17499
rect 42727 17431 42739 17465
rect 42773 17431 42785 17465
rect 42727 17397 42785 17431
rect 42727 17363 42739 17397
rect 42773 17363 42785 17397
rect 42727 17347 42785 17363
rect 43185 18621 43243 18637
rect 43185 18587 43197 18621
rect 43231 18587 43243 18621
rect 43185 18553 43243 18587
rect 43185 18519 43197 18553
rect 43231 18519 43243 18553
rect 43185 18485 43243 18519
rect 43185 18451 43197 18485
rect 43231 18451 43243 18485
rect 43185 18417 43243 18451
rect 43185 18383 43197 18417
rect 43231 18383 43243 18417
rect 43185 18349 43243 18383
rect 43185 18315 43197 18349
rect 43231 18315 43243 18349
rect 43185 18281 43243 18315
rect 43185 18247 43197 18281
rect 43231 18247 43243 18281
rect 43185 18213 43243 18247
rect 43185 18179 43197 18213
rect 43231 18179 43243 18213
rect 43185 18145 43243 18179
rect 43185 18111 43197 18145
rect 43231 18111 43243 18145
rect 43185 18077 43243 18111
rect 43185 18043 43197 18077
rect 43231 18043 43243 18077
rect 43185 18009 43243 18043
rect 43185 17975 43197 18009
rect 43231 17975 43243 18009
rect 43185 17941 43243 17975
rect 43185 17907 43197 17941
rect 43231 17907 43243 17941
rect 43185 17873 43243 17907
rect 43185 17839 43197 17873
rect 43231 17839 43243 17873
rect 43185 17805 43243 17839
rect 43185 17771 43197 17805
rect 43231 17771 43243 17805
rect 43185 17737 43243 17771
rect 43185 17703 43197 17737
rect 43231 17703 43243 17737
rect 43185 17669 43243 17703
rect 43185 17635 43197 17669
rect 43231 17635 43243 17669
rect 43185 17601 43243 17635
rect 43185 17567 43197 17601
rect 43231 17567 43243 17601
rect 43185 17533 43243 17567
rect 43185 17499 43197 17533
rect 43231 17499 43243 17533
rect 43185 17465 43243 17499
rect 43185 17431 43197 17465
rect 43231 17431 43243 17465
rect 43185 17397 43243 17431
rect 43185 17363 43197 17397
rect 43231 17363 43243 17397
rect 43185 17347 43243 17363
rect 43643 18621 43701 18637
rect 43643 18587 43655 18621
rect 43689 18587 43701 18621
rect 43643 18553 43701 18587
rect 43643 18519 43655 18553
rect 43689 18519 43701 18553
rect 43643 18485 43701 18519
rect 43643 18451 43655 18485
rect 43689 18451 43701 18485
rect 43643 18417 43701 18451
rect 43643 18383 43655 18417
rect 43689 18383 43701 18417
rect 43643 18349 43701 18383
rect 43643 18315 43655 18349
rect 43689 18315 43701 18349
rect 43643 18281 43701 18315
rect 43643 18247 43655 18281
rect 43689 18247 43701 18281
rect 43643 18213 43701 18247
rect 43643 18179 43655 18213
rect 43689 18179 43701 18213
rect 43643 18145 43701 18179
rect 43643 18111 43655 18145
rect 43689 18111 43701 18145
rect 43643 18077 43701 18111
rect 43643 18043 43655 18077
rect 43689 18043 43701 18077
rect 43643 18009 43701 18043
rect 43643 17975 43655 18009
rect 43689 17975 43701 18009
rect 43643 17941 43701 17975
rect 43643 17907 43655 17941
rect 43689 17907 43701 17941
rect 43643 17873 43701 17907
rect 43643 17839 43655 17873
rect 43689 17839 43701 17873
rect 43643 17805 43701 17839
rect 43643 17771 43655 17805
rect 43689 17771 43701 17805
rect 43643 17737 43701 17771
rect 43643 17703 43655 17737
rect 43689 17703 43701 17737
rect 43643 17669 43701 17703
rect 43643 17635 43655 17669
rect 43689 17635 43701 17669
rect 43643 17601 43701 17635
rect 43643 17567 43655 17601
rect 43689 17567 43701 17601
rect 43643 17533 43701 17567
rect 43643 17499 43655 17533
rect 43689 17499 43701 17533
rect 43643 17465 43701 17499
rect 43643 17431 43655 17465
rect 43689 17431 43701 17465
rect 43643 17397 43701 17431
rect 43643 17363 43655 17397
rect 43689 17363 43701 17397
rect 43643 17347 43701 17363
rect 44101 18621 44159 18637
rect 44101 18587 44113 18621
rect 44147 18587 44159 18621
rect 44101 18553 44159 18587
rect 44101 18519 44113 18553
rect 44147 18519 44159 18553
rect 44101 18485 44159 18519
rect 44101 18451 44113 18485
rect 44147 18451 44159 18485
rect 44101 18417 44159 18451
rect 44101 18383 44113 18417
rect 44147 18383 44159 18417
rect 44101 18349 44159 18383
rect 44101 18315 44113 18349
rect 44147 18315 44159 18349
rect 44101 18281 44159 18315
rect 44101 18247 44113 18281
rect 44147 18247 44159 18281
rect 44101 18213 44159 18247
rect 44101 18179 44113 18213
rect 44147 18179 44159 18213
rect 44101 18145 44159 18179
rect 44101 18111 44113 18145
rect 44147 18111 44159 18145
rect 44101 18077 44159 18111
rect 44101 18043 44113 18077
rect 44147 18043 44159 18077
rect 44101 18009 44159 18043
rect 44101 17975 44113 18009
rect 44147 17975 44159 18009
rect 44101 17941 44159 17975
rect 44101 17907 44113 17941
rect 44147 17907 44159 17941
rect 44101 17873 44159 17907
rect 44101 17839 44113 17873
rect 44147 17839 44159 17873
rect 44101 17805 44159 17839
rect 44101 17771 44113 17805
rect 44147 17771 44159 17805
rect 44101 17737 44159 17771
rect 44101 17703 44113 17737
rect 44147 17703 44159 17737
rect 44101 17669 44159 17703
rect 44101 17635 44113 17669
rect 44147 17635 44159 17669
rect 44101 17601 44159 17635
rect 44101 17567 44113 17601
rect 44147 17567 44159 17601
rect 44101 17533 44159 17567
rect 44101 17499 44113 17533
rect 44147 17499 44159 17533
rect 44101 17465 44159 17499
rect 44101 17431 44113 17465
rect 44147 17431 44159 17465
rect 44101 17397 44159 17431
rect 44101 17363 44113 17397
rect 44147 17363 44159 17397
rect 44101 17347 44159 17363
rect 44559 18621 44617 18637
rect 44559 18587 44571 18621
rect 44605 18587 44617 18621
rect 44559 18553 44617 18587
rect 44559 18519 44571 18553
rect 44605 18519 44617 18553
rect 44559 18485 44617 18519
rect 44559 18451 44571 18485
rect 44605 18451 44617 18485
rect 44559 18417 44617 18451
rect 44559 18383 44571 18417
rect 44605 18383 44617 18417
rect 44559 18349 44617 18383
rect 44559 18315 44571 18349
rect 44605 18315 44617 18349
rect 44559 18281 44617 18315
rect 44559 18247 44571 18281
rect 44605 18247 44617 18281
rect 44559 18213 44617 18247
rect 44559 18179 44571 18213
rect 44605 18179 44617 18213
rect 44559 18145 44617 18179
rect 44559 18111 44571 18145
rect 44605 18111 44617 18145
rect 44559 18077 44617 18111
rect 44559 18043 44571 18077
rect 44605 18043 44617 18077
rect 44559 18009 44617 18043
rect 44559 17975 44571 18009
rect 44605 17975 44617 18009
rect 44559 17941 44617 17975
rect 44559 17907 44571 17941
rect 44605 17907 44617 17941
rect 44559 17873 44617 17907
rect 44559 17839 44571 17873
rect 44605 17839 44617 17873
rect 44559 17805 44617 17839
rect 44559 17771 44571 17805
rect 44605 17771 44617 17805
rect 44559 17737 44617 17771
rect 44559 17703 44571 17737
rect 44605 17703 44617 17737
rect 44559 17669 44617 17703
rect 44559 17635 44571 17669
rect 44605 17635 44617 17669
rect 44559 17601 44617 17635
rect 44559 17567 44571 17601
rect 44605 17567 44617 17601
rect 44559 17533 44617 17567
rect 44559 17499 44571 17533
rect 44605 17499 44617 17533
rect 44559 17465 44617 17499
rect 44559 17431 44571 17465
rect 44605 17431 44617 17465
rect 44559 17397 44617 17431
rect 44559 17363 44571 17397
rect 44605 17363 44617 17397
rect 44559 17347 44617 17363
rect 45017 18621 45075 18637
rect 45017 18587 45029 18621
rect 45063 18587 45075 18621
rect 45017 18553 45075 18587
rect 45017 18519 45029 18553
rect 45063 18519 45075 18553
rect 45017 18485 45075 18519
rect 45017 18451 45029 18485
rect 45063 18451 45075 18485
rect 45017 18417 45075 18451
rect 45017 18383 45029 18417
rect 45063 18383 45075 18417
rect 45017 18349 45075 18383
rect 45017 18315 45029 18349
rect 45063 18315 45075 18349
rect 45017 18281 45075 18315
rect 45017 18247 45029 18281
rect 45063 18247 45075 18281
rect 45017 18213 45075 18247
rect 45017 18179 45029 18213
rect 45063 18179 45075 18213
rect 45017 18145 45075 18179
rect 45017 18111 45029 18145
rect 45063 18111 45075 18145
rect 45017 18077 45075 18111
rect 45017 18043 45029 18077
rect 45063 18043 45075 18077
rect 45017 18009 45075 18043
rect 45017 17975 45029 18009
rect 45063 17975 45075 18009
rect 45017 17941 45075 17975
rect 45017 17907 45029 17941
rect 45063 17907 45075 17941
rect 45017 17873 45075 17907
rect 45017 17839 45029 17873
rect 45063 17839 45075 17873
rect 45017 17805 45075 17839
rect 45017 17771 45029 17805
rect 45063 17771 45075 17805
rect 45017 17737 45075 17771
rect 45017 17703 45029 17737
rect 45063 17703 45075 17737
rect 45017 17669 45075 17703
rect 45017 17635 45029 17669
rect 45063 17635 45075 17669
rect 45017 17601 45075 17635
rect 45017 17567 45029 17601
rect 45063 17567 45075 17601
rect 45017 17533 45075 17567
rect 45017 17499 45029 17533
rect 45063 17499 45075 17533
rect 45017 17465 45075 17499
rect 45017 17431 45029 17465
rect 45063 17431 45075 17465
rect 45017 17397 45075 17431
rect 45017 17363 45029 17397
rect 45063 17363 45075 17397
rect 45017 17347 45075 17363
rect 45475 18621 45533 18637
rect 45475 18587 45487 18621
rect 45521 18587 45533 18621
rect 45475 18553 45533 18587
rect 45475 18519 45487 18553
rect 45521 18519 45533 18553
rect 45475 18485 45533 18519
rect 45475 18451 45487 18485
rect 45521 18451 45533 18485
rect 45475 18417 45533 18451
rect 45475 18383 45487 18417
rect 45521 18383 45533 18417
rect 45475 18349 45533 18383
rect 45475 18315 45487 18349
rect 45521 18315 45533 18349
rect 45475 18281 45533 18315
rect 45475 18247 45487 18281
rect 45521 18247 45533 18281
rect 45475 18213 45533 18247
rect 45475 18179 45487 18213
rect 45521 18179 45533 18213
rect 45475 18145 45533 18179
rect 45475 18111 45487 18145
rect 45521 18111 45533 18145
rect 45475 18077 45533 18111
rect 45475 18043 45487 18077
rect 45521 18043 45533 18077
rect 45475 18009 45533 18043
rect 45475 17975 45487 18009
rect 45521 17975 45533 18009
rect 45475 17941 45533 17975
rect 45475 17907 45487 17941
rect 45521 17907 45533 17941
rect 45475 17873 45533 17907
rect 45475 17839 45487 17873
rect 45521 17839 45533 17873
rect 45475 17805 45533 17839
rect 45475 17771 45487 17805
rect 45521 17771 45533 17805
rect 45475 17737 45533 17771
rect 45475 17703 45487 17737
rect 45521 17703 45533 17737
rect 45475 17669 45533 17703
rect 45475 17635 45487 17669
rect 45521 17635 45533 17669
rect 45475 17601 45533 17635
rect 45475 17567 45487 17601
rect 45521 17567 45533 17601
rect 45475 17533 45533 17567
rect 45475 17499 45487 17533
rect 45521 17499 45533 17533
rect 45475 17465 45533 17499
rect 45475 17431 45487 17465
rect 45521 17431 45533 17465
rect 45475 17397 45533 17431
rect 45475 17363 45487 17397
rect 45521 17363 45533 17397
rect 45475 17347 45533 17363
rect 45933 18621 45991 18637
rect 45933 18587 45945 18621
rect 45979 18587 45991 18621
rect 45933 18553 45991 18587
rect 45933 18519 45945 18553
rect 45979 18519 45991 18553
rect 45933 18485 45991 18519
rect 45933 18451 45945 18485
rect 45979 18451 45991 18485
rect 45933 18417 45991 18451
rect 45933 18383 45945 18417
rect 45979 18383 45991 18417
rect 45933 18349 45991 18383
rect 45933 18315 45945 18349
rect 45979 18315 45991 18349
rect 45933 18281 45991 18315
rect 45933 18247 45945 18281
rect 45979 18247 45991 18281
rect 45933 18213 45991 18247
rect 45933 18179 45945 18213
rect 45979 18179 45991 18213
rect 45933 18145 45991 18179
rect 45933 18111 45945 18145
rect 45979 18111 45991 18145
rect 45933 18077 45991 18111
rect 45933 18043 45945 18077
rect 45979 18043 45991 18077
rect 45933 18009 45991 18043
rect 45933 17975 45945 18009
rect 45979 17975 45991 18009
rect 45933 17941 45991 17975
rect 45933 17907 45945 17941
rect 45979 17907 45991 17941
rect 45933 17873 45991 17907
rect 45933 17839 45945 17873
rect 45979 17839 45991 17873
rect 45933 17805 45991 17839
rect 45933 17771 45945 17805
rect 45979 17771 45991 17805
rect 45933 17737 45991 17771
rect 45933 17703 45945 17737
rect 45979 17703 45991 17737
rect 45933 17669 45991 17703
rect 45933 17635 45945 17669
rect 45979 17635 45991 17669
rect 45933 17601 45991 17635
rect 45933 17567 45945 17601
rect 45979 17567 45991 17601
rect 45933 17533 45991 17567
rect 45933 17499 45945 17533
rect 45979 17499 45991 17533
rect 45933 17465 45991 17499
rect 45933 17431 45945 17465
rect 45979 17431 45991 17465
rect 45933 17397 45991 17431
rect 45933 17363 45945 17397
rect 45979 17363 45991 17397
rect 45933 17347 45991 17363
rect 46391 18621 46449 18637
rect 46391 18587 46403 18621
rect 46437 18587 46449 18621
rect 46391 18553 46449 18587
rect 46391 18519 46403 18553
rect 46437 18519 46449 18553
rect 46391 18485 46449 18519
rect 46391 18451 46403 18485
rect 46437 18451 46449 18485
rect 46391 18417 46449 18451
rect 46391 18383 46403 18417
rect 46437 18383 46449 18417
rect 46391 18349 46449 18383
rect 46391 18315 46403 18349
rect 46437 18315 46449 18349
rect 46391 18281 46449 18315
rect 46391 18247 46403 18281
rect 46437 18247 46449 18281
rect 46391 18213 46449 18247
rect 46391 18179 46403 18213
rect 46437 18179 46449 18213
rect 46391 18145 46449 18179
rect 46391 18111 46403 18145
rect 46437 18111 46449 18145
rect 46391 18077 46449 18111
rect 46391 18043 46403 18077
rect 46437 18043 46449 18077
rect 46391 18009 46449 18043
rect 46391 17975 46403 18009
rect 46437 17975 46449 18009
rect 46391 17941 46449 17975
rect 46391 17907 46403 17941
rect 46437 17907 46449 17941
rect 46391 17873 46449 17907
rect 46391 17839 46403 17873
rect 46437 17839 46449 17873
rect 46391 17805 46449 17839
rect 46391 17771 46403 17805
rect 46437 17771 46449 17805
rect 46391 17737 46449 17771
rect 46391 17703 46403 17737
rect 46437 17703 46449 17737
rect 46391 17669 46449 17703
rect 46391 17635 46403 17669
rect 46437 17635 46449 17669
rect 46391 17601 46449 17635
rect 46391 17567 46403 17601
rect 46437 17567 46449 17601
rect 46391 17533 46449 17567
rect 46391 17499 46403 17533
rect 46437 17499 46449 17533
rect 46391 17465 46449 17499
rect 46391 17431 46403 17465
rect 46437 17431 46449 17465
rect 46391 17397 46449 17431
rect 46391 17363 46403 17397
rect 46437 17363 46449 17397
rect 46391 17347 46449 17363
rect 46849 18621 46907 18637
rect 46849 18587 46861 18621
rect 46895 18587 46907 18621
rect 46849 18553 46907 18587
rect 46849 18519 46861 18553
rect 46895 18519 46907 18553
rect 46849 18485 46907 18519
rect 46849 18451 46861 18485
rect 46895 18451 46907 18485
rect 46849 18417 46907 18451
rect 46849 18383 46861 18417
rect 46895 18383 46907 18417
rect 46849 18349 46907 18383
rect 46849 18315 46861 18349
rect 46895 18315 46907 18349
rect 46849 18281 46907 18315
rect 46849 18247 46861 18281
rect 46895 18247 46907 18281
rect 46849 18213 46907 18247
rect 46849 18179 46861 18213
rect 46895 18179 46907 18213
rect 46849 18145 46907 18179
rect 46849 18111 46861 18145
rect 46895 18111 46907 18145
rect 46849 18077 46907 18111
rect 46849 18043 46861 18077
rect 46895 18043 46907 18077
rect 46849 18009 46907 18043
rect 46849 17975 46861 18009
rect 46895 17975 46907 18009
rect 46849 17941 46907 17975
rect 46849 17907 46861 17941
rect 46895 17907 46907 17941
rect 46849 17873 46907 17907
rect 46849 17839 46861 17873
rect 46895 17839 46907 17873
rect 46849 17805 46907 17839
rect 46849 17771 46861 17805
rect 46895 17771 46907 17805
rect 46849 17737 46907 17771
rect 46849 17703 46861 17737
rect 46895 17703 46907 17737
rect 46849 17669 46907 17703
rect 46849 17635 46861 17669
rect 46895 17635 46907 17669
rect 46849 17601 46907 17635
rect 46849 17567 46861 17601
rect 46895 17567 46907 17601
rect 46849 17533 46907 17567
rect 46849 17499 46861 17533
rect 46895 17499 46907 17533
rect 46849 17465 46907 17499
rect 46849 17431 46861 17465
rect 46895 17431 46907 17465
rect 46849 17397 46907 17431
rect 46849 17363 46861 17397
rect 46895 17363 46907 17397
rect 46849 17347 46907 17363
rect 47307 18621 47365 18637
rect 47307 18587 47319 18621
rect 47353 18587 47365 18621
rect 47307 18553 47365 18587
rect 47307 18519 47319 18553
rect 47353 18519 47365 18553
rect 47307 18485 47365 18519
rect 47307 18451 47319 18485
rect 47353 18451 47365 18485
rect 47307 18417 47365 18451
rect 47307 18383 47319 18417
rect 47353 18383 47365 18417
rect 47307 18349 47365 18383
rect 47307 18315 47319 18349
rect 47353 18315 47365 18349
rect 47307 18281 47365 18315
rect 47307 18247 47319 18281
rect 47353 18247 47365 18281
rect 47307 18213 47365 18247
rect 47307 18179 47319 18213
rect 47353 18179 47365 18213
rect 47307 18145 47365 18179
rect 47307 18111 47319 18145
rect 47353 18111 47365 18145
rect 47307 18077 47365 18111
rect 47307 18043 47319 18077
rect 47353 18043 47365 18077
rect 47307 18009 47365 18043
rect 47307 17975 47319 18009
rect 47353 17975 47365 18009
rect 47307 17941 47365 17975
rect 47307 17907 47319 17941
rect 47353 17907 47365 17941
rect 47307 17873 47365 17907
rect 47307 17839 47319 17873
rect 47353 17839 47365 17873
rect 47307 17805 47365 17839
rect 47307 17771 47319 17805
rect 47353 17771 47365 17805
rect 47307 17737 47365 17771
rect 47307 17703 47319 17737
rect 47353 17703 47365 17737
rect 47307 17669 47365 17703
rect 47307 17635 47319 17669
rect 47353 17635 47365 17669
rect 47307 17601 47365 17635
rect 47307 17567 47319 17601
rect 47353 17567 47365 17601
rect 47307 17533 47365 17567
rect 47307 17499 47319 17533
rect 47353 17499 47365 17533
rect 47307 17465 47365 17499
rect 47307 17431 47319 17465
rect 47353 17431 47365 17465
rect 47307 17397 47365 17431
rect 47307 17363 47319 17397
rect 47353 17363 47365 17397
rect 47307 17347 47365 17363
rect 47765 18621 47823 18637
rect 47765 18587 47777 18621
rect 47811 18587 47823 18621
rect 47765 18553 47823 18587
rect 47765 18519 47777 18553
rect 47811 18519 47823 18553
rect 47765 18485 47823 18519
rect 47765 18451 47777 18485
rect 47811 18451 47823 18485
rect 47765 18417 47823 18451
rect 47765 18383 47777 18417
rect 47811 18383 47823 18417
rect 47765 18349 47823 18383
rect 47765 18315 47777 18349
rect 47811 18315 47823 18349
rect 47765 18281 47823 18315
rect 47765 18247 47777 18281
rect 47811 18247 47823 18281
rect 47765 18213 47823 18247
rect 47765 18179 47777 18213
rect 47811 18179 47823 18213
rect 47765 18145 47823 18179
rect 47765 18111 47777 18145
rect 47811 18111 47823 18145
rect 47765 18077 47823 18111
rect 47765 18043 47777 18077
rect 47811 18043 47823 18077
rect 47765 18009 47823 18043
rect 47765 17975 47777 18009
rect 47811 17975 47823 18009
rect 47765 17941 47823 17975
rect 47765 17907 47777 17941
rect 47811 17907 47823 17941
rect 47765 17873 47823 17907
rect 47765 17839 47777 17873
rect 47811 17839 47823 17873
rect 47765 17805 47823 17839
rect 47765 17771 47777 17805
rect 47811 17771 47823 17805
rect 47765 17737 47823 17771
rect 47765 17703 47777 17737
rect 47811 17703 47823 17737
rect 47765 17669 47823 17703
rect 47765 17635 47777 17669
rect 47811 17635 47823 17669
rect 47765 17601 47823 17635
rect 47765 17567 47777 17601
rect 47811 17567 47823 17601
rect 47765 17533 47823 17567
rect 47765 17499 47777 17533
rect 47811 17499 47823 17533
rect 47765 17465 47823 17499
rect 47765 17431 47777 17465
rect 47811 17431 47823 17465
rect 47765 17397 47823 17431
rect 47765 17363 47777 17397
rect 47811 17363 47823 17397
rect 47765 17347 47823 17363
rect 48223 18621 48281 18637
rect 48223 18587 48235 18621
rect 48269 18587 48281 18621
rect 48223 18553 48281 18587
rect 48223 18519 48235 18553
rect 48269 18519 48281 18553
rect 48223 18485 48281 18519
rect 48223 18451 48235 18485
rect 48269 18451 48281 18485
rect 48223 18417 48281 18451
rect 48223 18383 48235 18417
rect 48269 18383 48281 18417
rect 48223 18349 48281 18383
rect 48223 18315 48235 18349
rect 48269 18315 48281 18349
rect 48223 18281 48281 18315
rect 48223 18247 48235 18281
rect 48269 18247 48281 18281
rect 48223 18213 48281 18247
rect 48223 18179 48235 18213
rect 48269 18179 48281 18213
rect 48223 18145 48281 18179
rect 48223 18111 48235 18145
rect 48269 18111 48281 18145
rect 48223 18077 48281 18111
rect 48223 18043 48235 18077
rect 48269 18043 48281 18077
rect 48223 18009 48281 18043
rect 48223 17975 48235 18009
rect 48269 17975 48281 18009
rect 48223 17941 48281 17975
rect 48223 17907 48235 17941
rect 48269 17907 48281 17941
rect 48223 17873 48281 17907
rect 48223 17839 48235 17873
rect 48269 17839 48281 17873
rect 48223 17805 48281 17839
rect 48223 17771 48235 17805
rect 48269 17771 48281 17805
rect 48223 17737 48281 17771
rect 48223 17703 48235 17737
rect 48269 17703 48281 17737
rect 48223 17669 48281 17703
rect 48223 17635 48235 17669
rect 48269 17635 48281 17669
rect 48223 17601 48281 17635
rect 48223 17567 48235 17601
rect 48269 17567 48281 17601
rect 48223 17533 48281 17567
rect 48223 17499 48235 17533
rect 48269 17499 48281 17533
rect 48223 17465 48281 17499
rect 48223 17431 48235 17465
rect 48269 17431 48281 17465
rect 48223 17397 48281 17431
rect 48223 17363 48235 17397
rect 48269 17363 48281 17397
rect 48223 17347 48281 17363
rect 48681 18621 48739 18637
rect 48681 18587 48693 18621
rect 48727 18587 48739 18621
rect 48681 18553 48739 18587
rect 48681 18519 48693 18553
rect 48727 18519 48739 18553
rect 48681 18485 48739 18519
rect 48681 18451 48693 18485
rect 48727 18451 48739 18485
rect 48681 18417 48739 18451
rect 48681 18383 48693 18417
rect 48727 18383 48739 18417
rect 48681 18349 48739 18383
rect 48681 18315 48693 18349
rect 48727 18315 48739 18349
rect 48681 18281 48739 18315
rect 48681 18247 48693 18281
rect 48727 18247 48739 18281
rect 48681 18213 48739 18247
rect 48681 18179 48693 18213
rect 48727 18179 48739 18213
rect 48681 18145 48739 18179
rect 48681 18111 48693 18145
rect 48727 18111 48739 18145
rect 48681 18077 48739 18111
rect 48681 18043 48693 18077
rect 48727 18043 48739 18077
rect 48681 18009 48739 18043
rect 48681 17975 48693 18009
rect 48727 17975 48739 18009
rect 48681 17941 48739 17975
rect 48681 17907 48693 17941
rect 48727 17907 48739 17941
rect 48681 17873 48739 17907
rect 48681 17839 48693 17873
rect 48727 17839 48739 17873
rect 48681 17805 48739 17839
rect 48681 17771 48693 17805
rect 48727 17771 48739 17805
rect 48681 17737 48739 17771
rect 48681 17703 48693 17737
rect 48727 17703 48739 17737
rect 48681 17669 48739 17703
rect 48681 17635 48693 17669
rect 48727 17635 48739 17669
rect 48681 17601 48739 17635
rect 48681 17567 48693 17601
rect 48727 17567 48739 17601
rect 48681 17533 48739 17567
rect 48681 17499 48693 17533
rect 48727 17499 48739 17533
rect 48681 17465 48739 17499
rect 48681 17431 48693 17465
rect 48727 17431 48739 17465
rect 48681 17397 48739 17431
rect 48681 17363 48693 17397
rect 48727 17363 48739 17397
rect 48681 17347 48739 17363
rect 49139 18621 49197 18637
rect 49139 18587 49151 18621
rect 49185 18587 49197 18621
rect 49139 18553 49197 18587
rect 49139 18519 49151 18553
rect 49185 18519 49197 18553
rect 49139 18485 49197 18519
rect 49139 18451 49151 18485
rect 49185 18451 49197 18485
rect 49139 18417 49197 18451
rect 49139 18383 49151 18417
rect 49185 18383 49197 18417
rect 49139 18349 49197 18383
rect 49139 18315 49151 18349
rect 49185 18315 49197 18349
rect 49139 18281 49197 18315
rect 49139 18247 49151 18281
rect 49185 18247 49197 18281
rect 49139 18213 49197 18247
rect 49139 18179 49151 18213
rect 49185 18179 49197 18213
rect 49139 18145 49197 18179
rect 49139 18111 49151 18145
rect 49185 18111 49197 18145
rect 49139 18077 49197 18111
rect 49139 18043 49151 18077
rect 49185 18043 49197 18077
rect 49139 18009 49197 18043
rect 49139 17975 49151 18009
rect 49185 17975 49197 18009
rect 49139 17941 49197 17975
rect 49139 17907 49151 17941
rect 49185 17907 49197 17941
rect 49139 17873 49197 17907
rect 49139 17839 49151 17873
rect 49185 17839 49197 17873
rect 49139 17805 49197 17839
rect 49139 17771 49151 17805
rect 49185 17771 49197 17805
rect 49139 17737 49197 17771
rect 49139 17703 49151 17737
rect 49185 17703 49197 17737
rect 49139 17669 49197 17703
rect 49139 17635 49151 17669
rect 49185 17635 49197 17669
rect 49139 17601 49197 17635
rect 49139 17567 49151 17601
rect 49185 17567 49197 17601
rect 49139 17533 49197 17567
rect 49139 17499 49151 17533
rect 49185 17499 49197 17533
rect 49139 17465 49197 17499
rect 49139 17431 49151 17465
rect 49185 17431 49197 17465
rect 49139 17397 49197 17431
rect 49139 17363 49151 17397
rect 49185 17363 49197 17397
rect 49139 17347 49197 17363
rect 49597 18621 49655 18637
rect 49597 18587 49609 18621
rect 49643 18587 49655 18621
rect 49597 18553 49655 18587
rect 49597 18519 49609 18553
rect 49643 18519 49655 18553
rect 49597 18485 49655 18519
rect 49597 18451 49609 18485
rect 49643 18451 49655 18485
rect 49597 18417 49655 18451
rect 49597 18383 49609 18417
rect 49643 18383 49655 18417
rect 49597 18349 49655 18383
rect 49597 18315 49609 18349
rect 49643 18315 49655 18349
rect 49597 18281 49655 18315
rect 49597 18247 49609 18281
rect 49643 18247 49655 18281
rect 49597 18213 49655 18247
rect 49597 18179 49609 18213
rect 49643 18179 49655 18213
rect 49597 18145 49655 18179
rect 49597 18111 49609 18145
rect 49643 18111 49655 18145
rect 49597 18077 49655 18111
rect 49597 18043 49609 18077
rect 49643 18043 49655 18077
rect 49597 18009 49655 18043
rect 49597 17975 49609 18009
rect 49643 17975 49655 18009
rect 49597 17941 49655 17975
rect 49597 17907 49609 17941
rect 49643 17907 49655 17941
rect 49597 17873 49655 17907
rect 49597 17839 49609 17873
rect 49643 17839 49655 17873
rect 49597 17805 49655 17839
rect 49597 17771 49609 17805
rect 49643 17771 49655 17805
rect 49597 17737 49655 17771
rect 49597 17703 49609 17737
rect 49643 17703 49655 17737
rect 49597 17669 49655 17703
rect 49597 17635 49609 17669
rect 49643 17635 49655 17669
rect 49597 17601 49655 17635
rect 49597 17567 49609 17601
rect 49643 17567 49655 17601
rect 49597 17533 49655 17567
rect 49597 17499 49609 17533
rect 49643 17499 49655 17533
rect 49597 17465 49655 17499
rect 49597 17431 49609 17465
rect 49643 17431 49655 17465
rect 49597 17397 49655 17431
rect 49597 17363 49609 17397
rect 49643 17363 49655 17397
rect 49597 17347 49655 17363
rect 50055 18621 50113 18637
rect 50055 18587 50067 18621
rect 50101 18587 50113 18621
rect 50055 18553 50113 18587
rect 50055 18519 50067 18553
rect 50101 18519 50113 18553
rect 50055 18485 50113 18519
rect 50055 18451 50067 18485
rect 50101 18451 50113 18485
rect 50055 18417 50113 18451
rect 50055 18383 50067 18417
rect 50101 18383 50113 18417
rect 50055 18349 50113 18383
rect 50055 18315 50067 18349
rect 50101 18315 50113 18349
rect 50055 18281 50113 18315
rect 50055 18247 50067 18281
rect 50101 18247 50113 18281
rect 50055 18213 50113 18247
rect 50055 18179 50067 18213
rect 50101 18179 50113 18213
rect 50055 18145 50113 18179
rect 50055 18111 50067 18145
rect 50101 18111 50113 18145
rect 50055 18077 50113 18111
rect 50055 18043 50067 18077
rect 50101 18043 50113 18077
rect 50055 18009 50113 18043
rect 50055 17975 50067 18009
rect 50101 17975 50113 18009
rect 50055 17941 50113 17975
rect 50055 17907 50067 17941
rect 50101 17907 50113 17941
rect 50055 17873 50113 17907
rect 50055 17839 50067 17873
rect 50101 17839 50113 17873
rect 50055 17805 50113 17839
rect 50055 17771 50067 17805
rect 50101 17771 50113 17805
rect 50055 17737 50113 17771
rect 50055 17703 50067 17737
rect 50101 17703 50113 17737
rect 50055 17669 50113 17703
rect 50055 17635 50067 17669
rect 50101 17635 50113 17669
rect 50055 17601 50113 17635
rect 50055 17567 50067 17601
rect 50101 17567 50113 17601
rect 50055 17533 50113 17567
rect 50055 17499 50067 17533
rect 50101 17499 50113 17533
rect 50055 17465 50113 17499
rect 50055 17431 50067 17465
rect 50101 17431 50113 17465
rect 50055 17397 50113 17431
rect 50055 17363 50067 17397
rect 50101 17363 50113 17397
rect 50055 17347 50113 17363
rect 50513 18621 50571 18637
rect 50513 18587 50525 18621
rect 50559 18587 50571 18621
rect 50513 18553 50571 18587
rect 50513 18519 50525 18553
rect 50559 18519 50571 18553
rect 50513 18485 50571 18519
rect 50513 18451 50525 18485
rect 50559 18451 50571 18485
rect 50513 18417 50571 18451
rect 50513 18383 50525 18417
rect 50559 18383 50571 18417
rect 50513 18349 50571 18383
rect 50513 18315 50525 18349
rect 50559 18315 50571 18349
rect 50513 18281 50571 18315
rect 50513 18247 50525 18281
rect 50559 18247 50571 18281
rect 50513 18213 50571 18247
rect 50513 18179 50525 18213
rect 50559 18179 50571 18213
rect 50513 18145 50571 18179
rect 50513 18111 50525 18145
rect 50559 18111 50571 18145
rect 50513 18077 50571 18111
rect 50513 18043 50525 18077
rect 50559 18043 50571 18077
rect 50513 18009 50571 18043
rect 50513 17975 50525 18009
rect 50559 17975 50571 18009
rect 50513 17941 50571 17975
rect 50513 17907 50525 17941
rect 50559 17907 50571 17941
rect 50513 17873 50571 17907
rect 50513 17839 50525 17873
rect 50559 17839 50571 17873
rect 50513 17805 50571 17839
rect 50513 17771 50525 17805
rect 50559 17771 50571 17805
rect 50513 17737 50571 17771
rect 50513 17703 50525 17737
rect 50559 17703 50571 17737
rect 50513 17669 50571 17703
rect 50513 17635 50525 17669
rect 50559 17635 50571 17669
rect 50513 17601 50571 17635
rect 50513 17567 50525 17601
rect 50559 17567 50571 17601
rect 50513 17533 50571 17567
rect 50513 17499 50525 17533
rect 50559 17499 50571 17533
rect 50513 17465 50571 17499
rect 50513 17431 50525 17465
rect 50559 17431 50571 17465
rect 50513 17397 50571 17431
rect 50513 17363 50525 17397
rect 50559 17363 50571 17397
rect 50513 17347 50571 17363
rect 50971 18621 51029 18637
rect 50971 18587 50983 18621
rect 51017 18587 51029 18621
rect 50971 18553 51029 18587
rect 50971 18519 50983 18553
rect 51017 18519 51029 18553
rect 50971 18485 51029 18519
rect 50971 18451 50983 18485
rect 51017 18451 51029 18485
rect 50971 18417 51029 18451
rect 50971 18383 50983 18417
rect 51017 18383 51029 18417
rect 50971 18349 51029 18383
rect 50971 18315 50983 18349
rect 51017 18315 51029 18349
rect 50971 18281 51029 18315
rect 50971 18247 50983 18281
rect 51017 18247 51029 18281
rect 50971 18213 51029 18247
rect 50971 18179 50983 18213
rect 51017 18179 51029 18213
rect 50971 18145 51029 18179
rect 50971 18111 50983 18145
rect 51017 18111 51029 18145
rect 50971 18077 51029 18111
rect 50971 18043 50983 18077
rect 51017 18043 51029 18077
rect 50971 18009 51029 18043
rect 50971 17975 50983 18009
rect 51017 17975 51029 18009
rect 50971 17941 51029 17975
rect 50971 17907 50983 17941
rect 51017 17907 51029 17941
rect 50971 17873 51029 17907
rect 50971 17839 50983 17873
rect 51017 17839 51029 17873
rect 50971 17805 51029 17839
rect 50971 17771 50983 17805
rect 51017 17771 51029 17805
rect 50971 17737 51029 17771
rect 50971 17703 50983 17737
rect 51017 17703 51029 17737
rect 50971 17669 51029 17703
rect 50971 17635 50983 17669
rect 51017 17635 51029 17669
rect 50971 17601 51029 17635
rect 50971 17567 50983 17601
rect 51017 17567 51029 17601
rect 50971 17533 51029 17567
rect 50971 17499 50983 17533
rect 51017 17499 51029 17533
rect 50971 17465 51029 17499
rect 50971 17431 50983 17465
rect 51017 17431 51029 17465
rect 50971 17397 51029 17431
rect 50971 17363 50983 17397
rect 51017 17363 51029 17397
rect 50971 17347 51029 17363
rect 51429 18621 51487 18637
rect 51429 18587 51441 18621
rect 51475 18587 51487 18621
rect 51429 18553 51487 18587
rect 51429 18519 51441 18553
rect 51475 18519 51487 18553
rect 51429 18485 51487 18519
rect 51429 18451 51441 18485
rect 51475 18451 51487 18485
rect 51429 18417 51487 18451
rect 51429 18383 51441 18417
rect 51475 18383 51487 18417
rect 51429 18349 51487 18383
rect 51429 18315 51441 18349
rect 51475 18315 51487 18349
rect 51429 18281 51487 18315
rect 51429 18247 51441 18281
rect 51475 18247 51487 18281
rect 51429 18213 51487 18247
rect 51429 18179 51441 18213
rect 51475 18179 51487 18213
rect 51429 18145 51487 18179
rect 51429 18111 51441 18145
rect 51475 18111 51487 18145
rect 51429 18077 51487 18111
rect 51429 18043 51441 18077
rect 51475 18043 51487 18077
rect 51429 18009 51487 18043
rect 51429 17975 51441 18009
rect 51475 17975 51487 18009
rect 51429 17941 51487 17975
rect 51429 17907 51441 17941
rect 51475 17907 51487 17941
rect 51429 17873 51487 17907
rect 51429 17839 51441 17873
rect 51475 17839 51487 17873
rect 51429 17805 51487 17839
rect 51429 17771 51441 17805
rect 51475 17771 51487 17805
rect 51429 17737 51487 17771
rect 51429 17703 51441 17737
rect 51475 17703 51487 17737
rect 51429 17669 51487 17703
rect 51429 17635 51441 17669
rect 51475 17635 51487 17669
rect 51429 17601 51487 17635
rect 51429 17567 51441 17601
rect 51475 17567 51487 17601
rect 51429 17533 51487 17567
rect 51429 17499 51441 17533
rect 51475 17499 51487 17533
rect 51429 17465 51487 17499
rect 51429 17431 51441 17465
rect 51475 17431 51487 17465
rect 51429 17397 51487 17431
rect 51429 17363 51441 17397
rect 51475 17363 51487 17397
rect 51429 17347 51487 17363
rect 51887 18621 51945 18637
rect 51887 18587 51899 18621
rect 51933 18587 51945 18621
rect 51887 18553 51945 18587
rect 51887 18519 51899 18553
rect 51933 18519 51945 18553
rect 51887 18485 51945 18519
rect 51887 18451 51899 18485
rect 51933 18451 51945 18485
rect 51887 18417 51945 18451
rect 51887 18383 51899 18417
rect 51933 18383 51945 18417
rect 51887 18349 51945 18383
rect 51887 18315 51899 18349
rect 51933 18315 51945 18349
rect 51887 18281 51945 18315
rect 51887 18247 51899 18281
rect 51933 18247 51945 18281
rect 51887 18213 51945 18247
rect 51887 18179 51899 18213
rect 51933 18179 51945 18213
rect 51887 18145 51945 18179
rect 51887 18111 51899 18145
rect 51933 18111 51945 18145
rect 51887 18077 51945 18111
rect 51887 18043 51899 18077
rect 51933 18043 51945 18077
rect 51887 18009 51945 18043
rect 51887 17975 51899 18009
rect 51933 17975 51945 18009
rect 51887 17941 51945 17975
rect 51887 17907 51899 17941
rect 51933 17907 51945 17941
rect 51887 17873 51945 17907
rect 51887 17839 51899 17873
rect 51933 17839 51945 17873
rect 51887 17805 51945 17839
rect 51887 17771 51899 17805
rect 51933 17771 51945 17805
rect 51887 17737 51945 17771
rect 51887 17703 51899 17737
rect 51933 17703 51945 17737
rect 51887 17669 51945 17703
rect 51887 17635 51899 17669
rect 51933 17635 51945 17669
rect 51887 17601 51945 17635
rect 51887 17567 51899 17601
rect 51933 17567 51945 17601
rect 51887 17533 51945 17567
rect 51887 17499 51899 17533
rect 51933 17499 51945 17533
rect 51887 17465 51945 17499
rect 51887 17431 51899 17465
rect 51933 17431 51945 17465
rect 51887 17397 51945 17431
rect 51887 17363 51899 17397
rect 51933 17363 51945 17397
rect 51887 17347 51945 17363
rect 52345 18621 52403 18637
rect 52345 18587 52357 18621
rect 52391 18587 52403 18621
rect 52345 18553 52403 18587
rect 52345 18519 52357 18553
rect 52391 18519 52403 18553
rect 52345 18485 52403 18519
rect 52345 18451 52357 18485
rect 52391 18451 52403 18485
rect 52345 18417 52403 18451
rect 52345 18383 52357 18417
rect 52391 18383 52403 18417
rect 52345 18349 52403 18383
rect 52345 18315 52357 18349
rect 52391 18315 52403 18349
rect 52345 18281 52403 18315
rect 52345 18247 52357 18281
rect 52391 18247 52403 18281
rect 52345 18213 52403 18247
rect 52345 18179 52357 18213
rect 52391 18179 52403 18213
rect 52345 18145 52403 18179
rect 52345 18111 52357 18145
rect 52391 18111 52403 18145
rect 52345 18077 52403 18111
rect 52345 18043 52357 18077
rect 52391 18043 52403 18077
rect 52345 18009 52403 18043
rect 52345 17975 52357 18009
rect 52391 17975 52403 18009
rect 52345 17941 52403 17975
rect 52345 17907 52357 17941
rect 52391 17907 52403 17941
rect 52345 17873 52403 17907
rect 52345 17839 52357 17873
rect 52391 17839 52403 17873
rect 52345 17805 52403 17839
rect 52345 17771 52357 17805
rect 52391 17771 52403 17805
rect 52345 17737 52403 17771
rect 52345 17703 52357 17737
rect 52391 17703 52403 17737
rect 52345 17669 52403 17703
rect 52345 17635 52357 17669
rect 52391 17635 52403 17669
rect 52345 17601 52403 17635
rect 52345 17567 52357 17601
rect 52391 17567 52403 17601
rect 52345 17533 52403 17567
rect 52345 17499 52357 17533
rect 52391 17499 52403 17533
rect 52345 17465 52403 17499
rect 52345 17431 52357 17465
rect 52391 17431 52403 17465
rect 52345 17397 52403 17431
rect 52345 17363 52357 17397
rect 52391 17363 52403 17397
rect 52345 17347 52403 17363
<< ndiffc >>
rect 23930 48395 23964 48429
rect 23930 48327 23964 48361
rect 23930 48259 23964 48293
rect 23930 48191 23964 48225
rect 23930 48123 23964 48157
rect 23930 48055 23964 48089
rect 23930 47987 23964 48021
rect 23930 47919 23964 47953
rect 23930 47851 23964 47885
rect 23930 47783 23964 47817
rect 23930 47715 23964 47749
rect 24388 48395 24422 48429
rect 24388 48327 24422 48361
rect 24388 48259 24422 48293
rect 24388 48191 24422 48225
rect 24388 48123 24422 48157
rect 24388 48055 24422 48089
rect 24388 47987 24422 48021
rect 24388 47919 24422 47953
rect 24388 47851 24422 47885
rect 24388 47783 24422 47817
rect 24388 47715 24422 47749
rect 14130 44635 14164 44669
rect 14130 44567 14164 44601
rect 14130 44499 14164 44533
rect 14130 44431 14164 44465
rect 14130 44363 14164 44397
rect 14130 44295 14164 44329
rect 14130 44227 14164 44261
rect 14130 44159 14164 44193
rect 14130 44091 14164 44125
rect 14130 44023 14164 44057
rect 14130 43955 14164 43989
rect 14588 44635 14622 44669
rect 14588 44567 14622 44601
rect 14588 44499 14622 44533
rect 14588 44431 14622 44465
rect 14588 44363 14622 44397
rect 14588 44295 14622 44329
rect 14588 44227 14622 44261
rect 14588 44159 14622 44193
rect 14588 44091 14622 44125
rect 14588 44023 14622 44057
rect 14588 43955 14622 43989
rect 37288 40875 37322 40909
rect 37288 40807 37322 40841
rect 37288 40739 37322 40773
rect 37288 40671 37322 40705
rect 37288 40603 37322 40637
rect 37288 40535 37322 40569
rect 37288 40467 37322 40501
rect 37288 40399 37322 40433
rect 37288 40331 37322 40365
rect 37288 40263 37322 40297
rect 37288 40195 37322 40229
rect 37746 40875 37780 40909
rect 37746 40807 37780 40841
rect 37746 40739 37780 40773
rect 37746 40671 37780 40705
rect 37746 40603 37780 40637
rect 37746 40535 37780 40569
rect 37746 40467 37780 40501
rect 37746 40399 37780 40433
rect 37746 40331 37780 40365
rect 37746 40263 37780 40297
rect 37746 40195 37780 40229
rect 38204 40875 38238 40909
rect 38204 40807 38238 40841
rect 38204 40739 38238 40773
rect 38204 40671 38238 40705
rect 38204 40603 38238 40637
rect 38204 40535 38238 40569
rect 38204 40467 38238 40501
rect 38204 40399 38238 40433
rect 38204 40331 38238 40365
rect 38204 40263 38238 40297
rect 38204 40195 38238 40229
rect 38662 40875 38696 40909
rect 38662 40807 38696 40841
rect 38662 40739 38696 40773
rect 38662 40671 38696 40705
rect 38662 40603 38696 40637
rect 38662 40535 38696 40569
rect 38662 40467 38696 40501
rect 38662 40399 38696 40433
rect 38662 40331 38696 40365
rect 38662 40263 38696 40297
rect 38662 40195 38696 40229
rect 39120 40875 39154 40909
rect 39120 40807 39154 40841
rect 39120 40739 39154 40773
rect 39120 40671 39154 40705
rect 39120 40603 39154 40637
rect 39120 40535 39154 40569
rect 39120 40467 39154 40501
rect 39120 40399 39154 40433
rect 39120 40331 39154 40365
rect 39120 40263 39154 40297
rect 39120 40195 39154 40229
rect 39578 40875 39612 40909
rect 39578 40807 39612 40841
rect 39578 40739 39612 40773
rect 39578 40671 39612 40705
rect 39578 40603 39612 40637
rect 39578 40535 39612 40569
rect 39578 40467 39612 40501
rect 39578 40399 39612 40433
rect 39578 40331 39612 40365
rect 39578 40263 39612 40297
rect 39578 40195 39612 40229
rect 40036 40875 40070 40909
rect 40036 40807 40070 40841
rect 40036 40739 40070 40773
rect 40036 40671 40070 40705
rect 40036 40603 40070 40637
rect 40036 40535 40070 40569
rect 40036 40467 40070 40501
rect 40036 40399 40070 40433
rect 40036 40331 40070 40365
rect 40036 40263 40070 40297
rect 40036 40195 40070 40229
rect 40494 40875 40528 40909
rect 40494 40807 40528 40841
rect 40494 40739 40528 40773
rect 40494 40671 40528 40705
rect 40494 40603 40528 40637
rect 40494 40535 40528 40569
rect 40494 40467 40528 40501
rect 40494 40399 40528 40433
rect 40494 40331 40528 40365
rect 40494 40263 40528 40297
rect 40494 40195 40528 40229
rect 40952 40875 40986 40909
rect 40952 40807 40986 40841
rect 40952 40739 40986 40773
rect 40952 40671 40986 40705
rect 40952 40603 40986 40637
rect 40952 40535 40986 40569
rect 40952 40467 40986 40501
rect 40952 40399 40986 40433
rect 40952 40331 40986 40365
rect 40952 40263 40986 40297
rect 40952 40195 40986 40229
rect 41410 40875 41444 40909
rect 41410 40807 41444 40841
rect 41410 40739 41444 40773
rect 41410 40671 41444 40705
rect 41410 40603 41444 40637
rect 41410 40535 41444 40569
rect 41410 40467 41444 40501
rect 41410 40399 41444 40433
rect 41410 40331 41444 40365
rect 41410 40263 41444 40297
rect 41410 40195 41444 40229
rect 25430 37115 25464 37149
rect 25430 37047 25464 37081
rect 25430 36979 25464 37013
rect 25430 36911 25464 36945
rect 25430 36843 25464 36877
rect 25430 36775 25464 36809
rect 25430 36707 25464 36741
rect 25430 36639 25464 36673
rect 25430 36571 25464 36605
rect 25430 36503 25464 36537
rect 25430 36435 25464 36469
rect 25888 37115 25922 37149
rect 25888 37047 25922 37081
rect 25888 36979 25922 37013
rect 25888 36911 25922 36945
rect 25888 36843 25922 36877
rect 25888 36775 25922 36809
rect 25888 36707 25922 36741
rect 25888 36639 25922 36673
rect 25888 36571 25922 36605
rect 25888 36503 25922 36537
rect 25888 36435 25922 36469
rect 26346 37115 26380 37149
rect 26346 37047 26380 37081
rect 26346 36979 26380 37013
rect 26346 36911 26380 36945
rect 26346 36843 26380 36877
rect 26346 36775 26380 36809
rect 26346 36707 26380 36741
rect 26346 36639 26380 36673
rect 26346 36571 26380 36605
rect 26346 36503 26380 36537
rect 26346 36435 26380 36469
rect 26804 37115 26838 37149
rect 26804 37047 26838 37081
rect 26804 36979 26838 37013
rect 26804 36911 26838 36945
rect 26804 36843 26838 36877
rect 26804 36775 26838 36809
rect 26804 36707 26838 36741
rect 26804 36639 26838 36673
rect 26804 36571 26838 36605
rect 26804 36503 26838 36537
rect 26804 36435 26838 36469
rect 27262 37115 27296 37149
rect 27262 37047 27296 37081
rect 27262 36979 27296 37013
rect 27262 36911 27296 36945
rect 27262 36843 27296 36877
rect 27262 36775 27296 36809
rect 27262 36707 27296 36741
rect 27262 36639 27296 36673
rect 27262 36571 27296 36605
rect 27262 36503 27296 36537
rect 27262 36435 27296 36469
rect 27720 37115 27754 37149
rect 27720 37047 27754 37081
rect 27720 36979 27754 37013
rect 27720 36911 27754 36945
rect 27720 36843 27754 36877
rect 27720 36775 27754 36809
rect 27720 36707 27754 36741
rect 27720 36639 27754 36673
rect 27720 36571 27754 36605
rect 27720 36503 27754 36537
rect 27720 36435 27754 36469
rect 28178 37115 28212 37149
rect 28178 37047 28212 37081
rect 28178 36979 28212 37013
rect 28178 36911 28212 36945
rect 28178 36843 28212 36877
rect 28178 36775 28212 36809
rect 28178 36707 28212 36741
rect 28178 36639 28212 36673
rect 28178 36571 28212 36605
rect 28178 36503 28212 36537
rect 28178 36435 28212 36469
rect 28636 37115 28670 37149
rect 28636 37047 28670 37081
rect 28636 36979 28670 37013
rect 28636 36911 28670 36945
rect 28636 36843 28670 36877
rect 28636 36775 28670 36809
rect 28636 36707 28670 36741
rect 28636 36639 28670 36673
rect 28636 36571 28670 36605
rect 28636 36503 28670 36537
rect 28636 36435 28670 36469
rect 29094 37115 29128 37149
rect 29094 37047 29128 37081
rect 29094 36979 29128 37013
rect 29094 36911 29128 36945
rect 29094 36843 29128 36877
rect 29094 36775 29128 36809
rect 29094 36707 29128 36741
rect 29094 36639 29128 36673
rect 29094 36571 29128 36605
rect 29094 36503 29128 36537
rect 29094 36435 29128 36469
rect 29552 37115 29586 37149
rect 29552 37047 29586 37081
rect 29552 36979 29586 37013
rect 29552 36911 29586 36945
rect 29552 36843 29586 36877
rect 29552 36775 29586 36809
rect 29552 36707 29586 36741
rect 29552 36639 29586 36673
rect 29552 36571 29586 36605
rect 29552 36503 29586 36537
rect 29552 36435 29586 36469
rect 25430 25835 25464 25869
rect 25430 25767 25464 25801
rect 25430 25699 25464 25733
rect 25430 25631 25464 25665
rect 25430 25563 25464 25597
rect 25430 25495 25464 25529
rect 25430 25427 25464 25461
rect 25430 25359 25464 25393
rect 25430 25291 25464 25325
rect 25430 25223 25464 25257
rect 25430 25155 25464 25189
rect 25888 25835 25922 25869
rect 25888 25767 25922 25801
rect 25888 25699 25922 25733
rect 25888 25631 25922 25665
rect 25888 25563 25922 25597
rect 25888 25495 25922 25529
rect 25888 25427 25922 25461
rect 25888 25359 25922 25393
rect 25888 25291 25922 25325
rect 25888 25223 25922 25257
rect 25888 25155 25922 25189
rect 26346 25835 26380 25869
rect 26346 25767 26380 25801
rect 26346 25699 26380 25733
rect 26346 25631 26380 25665
rect 26346 25563 26380 25597
rect 26346 25495 26380 25529
rect 26346 25427 26380 25461
rect 26346 25359 26380 25393
rect 26346 25291 26380 25325
rect 26346 25223 26380 25257
rect 26346 25155 26380 25189
rect 26804 25835 26838 25869
rect 26804 25767 26838 25801
rect 26804 25699 26838 25733
rect 26804 25631 26838 25665
rect 26804 25563 26838 25597
rect 26804 25495 26838 25529
rect 26804 25427 26838 25461
rect 26804 25359 26838 25393
rect 26804 25291 26838 25325
rect 26804 25223 26838 25257
rect 26804 25155 26838 25189
rect 27262 25835 27296 25869
rect 27262 25767 27296 25801
rect 27262 25699 27296 25733
rect 27262 25631 27296 25665
rect 27262 25563 27296 25597
rect 27262 25495 27296 25529
rect 27262 25427 27296 25461
rect 27262 25359 27296 25393
rect 27262 25291 27296 25325
rect 27262 25223 27296 25257
rect 27262 25155 27296 25189
rect 27720 25835 27754 25869
rect 27720 25767 27754 25801
rect 27720 25699 27754 25733
rect 27720 25631 27754 25665
rect 27720 25563 27754 25597
rect 27720 25495 27754 25529
rect 27720 25427 27754 25461
rect 27720 25359 27754 25393
rect 27720 25291 27754 25325
rect 27720 25223 27754 25257
rect 27720 25155 27754 25189
rect 28178 25835 28212 25869
rect 28178 25767 28212 25801
rect 28178 25699 28212 25733
rect 28178 25631 28212 25665
rect 28178 25563 28212 25597
rect 28178 25495 28212 25529
rect 28178 25427 28212 25461
rect 28178 25359 28212 25393
rect 28178 25291 28212 25325
rect 28178 25223 28212 25257
rect 28178 25155 28212 25189
rect 28636 25835 28670 25869
rect 28636 25767 28670 25801
rect 28636 25699 28670 25733
rect 28636 25631 28670 25665
rect 28636 25563 28670 25597
rect 28636 25495 28670 25529
rect 28636 25427 28670 25461
rect 28636 25359 28670 25393
rect 28636 25291 28670 25325
rect 28636 25223 28670 25257
rect 28636 25155 28670 25189
rect 29094 25835 29128 25869
rect 29094 25767 29128 25801
rect 29094 25699 29128 25733
rect 29094 25631 29128 25665
rect 29094 25563 29128 25597
rect 29094 25495 29128 25529
rect 29094 25427 29128 25461
rect 29094 25359 29128 25393
rect 29094 25291 29128 25325
rect 29094 25223 29128 25257
rect 29094 25155 29128 25189
rect 29552 25835 29586 25869
rect 29552 25767 29586 25801
rect 29552 25699 29586 25733
rect 29552 25631 29586 25665
rect 29552 25563 29586 25597
rect 29552 25495 29586 25529
rect 29552 25427 29586 25461
rect 29552 25359 29586 25393
rect 29552 25291 29586 25325
rect 29552 25223 29586 25257
rect 29552 25155 29586 25189
<< pdiffc >>
rect 24877 48667 24911 48701
rect 24877 48599 24911 48633
rect 24877 48531 24911 48565
rect 24877 48463 24911 48497
rect 24877 48395 24911 48429
rect 24877 48327 24911 48361
rect 24877 48259 24911 48293
rect 24877 48191 24911 48225
rect 24877 48123 24911 48157
rect 24877 48055 24911 48089
rect 24877 47987 24911 48021
rect 24877 47919 24911 47953
rect 24877 47851 24911 47885
rect 24877 47783 24911 47817
rect 24877 47715 24911 47749
rect 24877 47647 24911 47681
rect 24877 47579 24911 47613
rect 24877 47511 24911 47545
rect 24877 47443 24911 47477
rect 25335 48667 25369 48701
rect 25335 48599 25369 48633
rect 25335 48531 25369 48565
rect 25335 48463 25369 48497
rect 25335 48395 25369 48429
rect 25335 48327 25369 48361
rect 25335 48259 25369 48293
rect 25335 48191 25369 48225
rect 25335 48123 25369 48157
rect 25335 48055 25369 48089
rect 25335 47987 25369 48021
rect 25335 47919 25369 47953
rect 25335 47851 25369 47885
rect 25335 47783 25369 47817
rect 25335 47715 25369 47749
rect 25335 47647 25369 47681
rect 25335 47579 25369 47613
rect 25335 47511 25369 47545
rect 25335 47443 25369 47477
rect 25793 48667 25827 48701
rect 25793 48599 25827 48633
rect 25793 48531 25827 48565
rect 25793 48463 25827 48497
rect 25793 48395 25827 48429
rect 25793 48327 25827 48361
rect 25793 48259 25827 48293
rect 25793 48191 25827 48225
rect 25793 48123 25827 48157
rect 25793 48055 25827 48089
rect 25793 47987 25827 48021
rect 25793 47919 25827 47953
rect 25793 47851 25827 47885
rect 25793 47783 25827 47817
rect 25793 47715 25827 47749
rect 25793 47647 25827 47681
rect 25793 47579 25827 47613
rect 25793 47511 25827 47545
rect 25793 47443 25827 47477
rect 26251 48667 26285 48701
rect 26251 48599 26285 48633
rect 26251 48531 26285 48565
rect 26251 48463 26285 48497
rect 26251 48395 26285 48429
rect 26251 48327 26285 48361
rect 26251 48259 26285 48293
rect 26251 48191 26285 48225
rect 26251 48123 26285 48157
rect 26251 48055 26285 48089
rect 26251 47987 26285 48021
rect 26251 47919 26285 47953
rect 26251 47851 26285 47885
rect 26251 47783 26285 47817
rect 26251 47715 26285 47749
rect 26251 47647 26285 47681
rect 26251 47579 26285 47613
rect 26251 47511 26285 47545
rect 26251 47443 26285 47477
rect 26709 48667 26743 48701
rect 26709 48599 26743 48633
rect 26709 48531 26743 48565
rect 26709 48463 26743 48497
rect 26709 48395 26743 48429
rect 26709 48327 26743 48361
rect 26709 48259 26743 48293
rect 26709 48191 26743 48225
rect 26709 48123 26743 48157
rect 26709 48055 26743 48089
rect 26709 47987 26743 48021
rect 26709 47919 26743 47953
rect 26709 47851 26743 47885
rect 26709 47783 26743 47817
rect 26709 47715 26743 47749
rect 26709 47647 26743 47681
rect 26709 47579 26743 47613
rect 26709 47511 26743 47545
rect 26709 47443 26743 47477
rect 27167 48667 27201 48701
rect 27167 48599 27201 48633
rect 27167 48531 27201 48565
rect 27167 48463 27201 48497
rect 27167 48395 27201 48429
rect 27167 48327 27201 48361
rect 27167 48259 27201 48293
rect 27167 48191 27201 48225
rect 27167 48123 27201 48157
rect 27167 48055 27201 48089
rect 27167 47987 27201 48021
rect 27167 47919 27201 47953
rect 27167 47851 27201 47885
rect 27167 47783 27201 47817
rect 27167 47715 27201 47749
rect 27167 47647 27201 47681
rect 27167 47579 27201 47613
rect 27167 47511 27201 47545
rect 27167 47443 27201 47477
rect 27625 48667 27659 48701
rect 27625 48599 27659 48633
rect 27625 48531 27659 48565
rect 27625 48463 27659 48497
rect 27625 48395 27659 48429
rect 27625 48327 27659 48361
rect 27625 48259 27659 48293
rect 27625 48191 27659 48225
rect 27625 48123 27659 48157
rect 27625 48055 27659 48089
rect 27625 47987 27659 48021
rect 27625 47919 27659 47953
rect 27625 47851 27659 47885
rect 27625 47783 27659 47817
rect 27625 47715 27659 47749
rect 27625 47647 27659 47681
rect 27625 47579 27659 47613
rect 27625 47511 27659 47545
rect 27625 47443 27659 47477
rect 28083 48667 28117 48701
rect 28083 48599 28117 48633
rect 28083 48531 28117 48565
rect 28083 48463 28117 48497
rect 28083 48395 28117 48429
rect 28083 48327 28117 48361
rect 28083 48259 28117 48293
rect 28083 48191 28117 48225
rect 28083 48123 28117 48157
rect 28083 48055 28117 48089
rect 28083 47987 28117 48021
rect 28083 47919 28117 47953
rect 28083 47851 28117 47885
rect 28083 47783 28117 47817
rect 28083 47715 28117 47749
rect 28083 47647 28117 47681
rect 28083 47579 28117 47613
rect 28083 47511 28117 47545
rect 28083 47443 28117 47477
rect 28541 48667 28575 48701
rect 28541 48599 28575 48633
rect 28541 48531 28575 48565
rect 28541 48463 28575 48497
rect 28541 48395 28575 48429
rect 28541 48327 28575 48361
rect 28541 48259 28575 48293
rect 28541 48191 28575 48225
rect 28541 48123 28575 48157
rect 28541 48055 28575 48089
rect 28541 47987 28575 48021
rect 28541 47919 28575 47953
rect 28541 47851 28575 47885
rect 28541 47783 28575 47817
rect 28541 47715 28575 47749
rect 28541 47647 28575 47681
rect 28541 47579 28575 47613
rect 28541 47511 28575 47545
rect 28541 47443 28575 47477
rect 28999 48667 29033 48701
rect 28999 48599 29033 48633
rect 28999 48531 29033 48565
rect 28999 48463 29033 48497
rect 28999 48395 29033 48429
rect 28999 48327 29033 48361
rect 28999 48259 29033 48293
rect 28999 48191 29033 48225
rect 28999 48123 29033 48157
rect 28999 48055 29033 48089
rect 28999 47987 29033 48021
rect 28999 47919 29033 47953
rect 28999 47851 29033 47885
rect 28999 47783 29033 47817
rect 28999 47715 29033 47749
rect 28999 47647 29033 47681
rect 28999 47579 29033 47613
rect 28999 47511 29033 47545
rect 28999 47443 29033 47477
rect 29457 48667 29491 48701
rect 29457 48599 29491 48633
rect 29457 48531 29491 48565
rect 29457 48463 29491 48497
rect 29457 48395 29491 48429
rect 29457 48327 29491 48361
rect 29457 48259 29491 48293
rect 29457 48191 29491 48225
rect 29457 48123 29491 48157
rect 29457 48055 29491 48089
rect 29457 47987 29491 48021
rect 29457 47919 29491 47953
rect 29457 47851 29491 47885
rect 29457 47783 29491 47817
rect 29457 47715 29491 47749
rect 29457 47647 29491 47681
rect 29457 47579 29491 47613
rect 29457 47511 29491 47545
rect 29457 47443 29491 47477
rect 29915 48667 29949 48701
rect 29915 48599 29949 48633
rect 29915 48531 29949 48565
rect 29915 48463 29949 48497
rect 29915 48395 29949 48429
rect 29915 48327 29949 48361
rect 29915 48259 29949 48293
rect 29915 48191 29949 48225
rect 29915 48123 29949 48157
rect 29915 48055 29949 48089
rect 29915 47987 29949 48021
rect 29915 47919 29949 47953
rect 29915 47851 29949 47885
rect 29915 47783 29949 47817
rect 29915 47715 29949 47749
rect 29915 47647 29949 47681
rect 29915 47579 29949 47613
rect 29915 47511 29949 47545
rect 29915 47443 29949 47477
rect 30373 48667 30407 48701
rect 30373 48599 30407 48633
rect 30373 48531 30407 48565
rect 30373 48463 30407 48497
rect 30373 48395 30407 48429
rect 30373 48327 30407 48361
rect 30373 48259 30407 48293
rect 30373 48191 30407 48225
rect 30373 48123 30407 48157
rect 30373 48055 30407 48089
rect 30373 47987 30407 48021
rect 30373 47919 30407 47953
rect 30373 47851 30407 47885
rect 30373 47783 30407 47817
rect 30373 47715 30407 47749
rect 30373 47647 30407 47681
rect 30373 47579 30407 47613
rect 30373 47511 30407 47545
rect 30373 47443 30407 47477
rect 30831 48667 30865 48701
rect 30831 48599 30865 48633
rect 30831 48531 30865 48565
rect 30831 48463 30865 48497
rect 30831 48395 30865 48429
rect 30831 48327 30865 48361
rect 30831 48259 30865 48293
rect 30831 48191 30865 48225
rect 30831 48123 30865 48157
rect 30831 48055 30865 48089
rect 30831 47987 30865 48021
rect 30831 47919 30865 47953
rect 30831 47851 30865 47885
rect 30831 47783 30865 47817
rect 30831 47715 30865 47749
rect 30831 47647 30865 47681
rect 30831 47579 30865 47613
rect 30831 47511 30865 47545
rect 30831 47443 30865 47477
rect 31289 48667 31323 48701
rect 31289 48599 31323 48633
rect 31289 48531 31323 48565
rect 31289 48463 31323 48497
rect 31289 48395 31323 48429
rect 31289 48327 31323 48361
rect 31289 48259 31323 48293
rect 31289 48191 31323 48225
rect 31289 48123 31323 48157
rect 31289 48055 31323 48089
rect 31289 47987 31323 48021
rect 31289 47919 31323 47953
rect 31289 47851 31323 47885
rect 31289 47783 31323 47817
rect 31289 47715 31323 47749
rect 31289 47647 31323 47681
rect 31289 47579 31323 47613
rect 31289 47511 31323 47545
rect 31289 47443 31323 47477
rect 31747 48667 31781 48701
rect 31747 48599 31781 48633
rect 31747 48531 31781 48565
rect 31747 48463 31781 48497
rect 31747 48395 31781 48429
rect 31747 48327 31781 48361
rect 31747 48259 31781 48293
rect 31747 48191 31781 48225
rect 31747 48123 31781 48157
rect 31747 48055 31781 48089
rect 31747 47987 31781 48021
rect 31747 47919 31781 47953
rect 31747 47851 31781 47885
rect 31747 47783 31781 47817
rect 31747 47715 31781 47749
rect 31747 47647 31781 47681
rect 31747 47579 31781 47613
rect 31747 47511 31781 47545
rect 31747 47443 31781 47477
rect 32205 48667 32239 48701
rect 32205 48599 32239 48633
rect 32205 48531 32239 48565
rect 32205 48463 32239 48497
rect 32205 48395 32239 48429
rect 32205 48327 32239 48361
rect 32205 48259 32239 48293
rect 32205 48191 32239 48225
rect 32205 48123 32239 48157
rect 32205 48055 32239 48089
rect 32205 47987 32239 48021
rect 32205 47919 32239 47953
rect 32205 47851 32239 47885
rect 32205 47783 32239 47817
rect 32205 47715 32239 47749
rect 32205 47647 32239 47681
rect 32205 47579 32239 47613
rect 32205 47511 32239 47545
rect 32205 47443 32239 47477
rect 32663 48667 32697 48701
rect 32663 48599 32697 48633
rect 32663 48531 32697 48565
rect 32663 48463 32697 48497
rect 32663 48395 32697 48429
rect 32663 48327 32697 48361
rect 32663 48259 32697 48293
rect 32663 48191 32697 48225
rect 32663 48123 32697 48157
rect 32663 48055 32697 48089
rect 32663 47987 32697 48021
rect 32663 47919 32697 47953
rect 32663 47851 32697 47885
rect 32663 47783 32697 47817
rect 32663 47715 32697 47749
rect 32663 47647 32697 47681
rect 32663 47579 32697 47613
rect 32663 47511 32697 47545
rect 32663 47443 32697 47477
rect 33121 48667 33155 48701
rect 33121 48599 33155 48633
rect 33121 48531 33155 48565
rect 33121 48463 33155 48497
rect 33121 48395 33155 48429
rect 33121 48327 33155 48361
rect 33121 48259 33155 48293
rect 33121 48191 33155 48225
rect 33121 48123 33155 48157
rect 33121 48055 33155 48089
rect 33121 47987 33155 48021
rect 33121 47919 33155 47953
rect 33121 47851 33155 47885
rect 33121 47783 33155 47817
rect 33121 47715 33155 47749
rect 33121 47647 33155 47681
rect 33121 47579 33155 47613
rect 33121 47511 33155 47545
rect 33121 47443 33155 47477
rect 33579 48667 33613 48701
rect 33579 48599 33613 48633
rect 33579 48531 33613 48565
rect 33579 48463 33613 48497
rect 33579 48395 33613 48429
rect 33579 48327 33613 48361
rect 33579 48259 33613 48293
rect 33579 48191 33613 48225
rect 33579 48123 33613 48157
rect 33579 48055 33613 48089
rect 33579 47987 33613 48021
rect 33579 47919 33613 47953
rect 33579 47851 33613 47885
rect 33579 47783 33613 47817
rect 33579 47715 33613 47749
rect 33579 47647 33613 47681
rect 33579 47579 33613 47613
rect 33579 47511 33613 47545
rect 33579 47443 33613 47477
rect 34037 48667 34071 48701
rect 34037 48599 34071 48633
rect 34037 48531 34071 48565
rect 34037 48463 34071 48497
rect 34037 48395 34071 48429
rect 34037 48327 34071 48361
rect 34037 48259 34071 48293
rect 34037 48191 34071 48225
rect 34037 48123 34071 48157
rect 34037 48055 34071 48089
rect 34037 47987 34071 48021
rect 34037 47919 34071 47953
rect 34037 47851 34071 47885
rect 34037 47783 34071 47817
rect 34037 47715 34071 47749
rect 34037 47647 34071 47681
rect 34037 47579 34071 47613
rect 34037 47511 34071 47545
rect 34037 47443 34071 47477
rect 34495 48667 34529 48701
rect 34495 48599 34529 48633
rect 34495 48531 34529 48565
rect 34495 48463 34529 48497
rect 34495 48395 34529 48429
rect 34495 48327 34529 48361
rect 34495 48259 34529 48293
rect 34495 48191 34529 48225
rect 34495 48123 34529 48157
rect 34495 48055 34529 48089
rect 34495 47987 34529 48021
rect 34495 47919 34529 47953
rect 34495 47851 34529 47885
rect 34495 47783 34529 47817
rect 34495 47715 34529 47749
rect 34495 47647 34529 47681
rect 34495 47579 34529 47613
rect 34495 47511 34529 47545
rect 34495 47443 34529 47477
rect 34953 48667 34987 48701
rect 34953 48599 34987 48633
rect 34953 48531 34987 48565
rect 34953 48463 34987 48497
rect 34953 48395 34987 48429
rect 34953 48327 34987 48361
rect 34953 48259 34987 48293
rect 34953 48191 34987 48225
rect 34953 48123 34987 48157
rect 34953 48055 34987 48089
rect 34953 47987 34987 48021
rect 34953 47919 34987 47953
rect 34953 47851 34987 47885
rect 34953 47783 34987 47817
rect 34953 47715 34987 47749
rect 34953 47647 34987 47681
rect 34953 47579 34987 47613
rect 34953 47511 34987 47545
rect 34953 47443 34987 47477
rect 35411 48667 35445 48701
rect 35411 48599 35445 48633
rect 35411 48531 35445 48565
rect 35411 48463 35445 48497
rect 35411 48395 35445 48429
rect 35411 48327 35445 48361
rect 35411 48259 35445 48293
rect 35411 48191 35445 48225
rect 35411 48123 35445 48157
rect 35411 48055 35445 48089
rect 35411 47987 35445 48021
rect 35411 47919 35445 47953
rect 35411 47851 35445 47885
rect 35411 47783 35445 47817
rect 35411 47715 35445 47749
rect 35411 47647 35445 47681
rect 35411 47579 35445 47613
rect 35411 47511 35445 47545
rect 35411 47443 35445 47477
rect 35869 48667 35903 48701
rect 35869 48599 35903 48633
rect 35869 48531 35903 48565
rect 35869 48463 35903 48497
rect 35869 48395 35903 48429
rect 35869 48327 35903 48361
rect 35869 48259 35903 48293
rect 35869 48191 35903 48225
rect 35869 48123 35903 48157
rect 35869 48055 35903 48089
rect 35869 47987 35903 48021
rect 35869 47919 35903 47953
rect 35869 47851 35903 47885
rect 35869 47783 35903 47817
rect 35869 47715 35903 47749
rect 35869 47647 35903 47681
rect 35869 47579 35903 47613
rect 35869 47511 35903 47545
rect 35869 47443 35903 47477
rect 36327 48667 36361 48701
rect 36327 48599 36361 48633
rect 36327 48531 36361 48565
rect 36327 48463 36361 48497
rect 36327 48395 36361 48429
rect 36327 48327 36361 48361
rect 36327 48259 36361 48293
rect 36327 48191 36361 48225
rect 36327 48123 36361 48157
rect 36327 48055 36361 48089
rect 36327 47987 36361 48021
rect 36327 47919 36361 47953
rect 36327 47851 36361 47885
rect 36327 47783 36361 47817
rect 36327 47715 36361 47749
rect 36327 47647 36361 47681
rect 36327 47579 36361 47613
rect 36327 47511 36361 47545
rect 36327 47443 36361 47477
rect 36785 48667 36819 48701
rect 36785 48599 36819 48633
rect 36785 48531 36819 48565
rect 36785 48463 36819 48497
rect 36785 48395 36819 48429
rect 36785 48327 36819 48361
rect 36785 48259 36819 48293
rect 36785 48191 36819 48225
rect 36785 48123 36819 48157
rect 36785 48055 36819 48089
rect 36785 47987 36819 48021
rect 36785 47919 36819 47953
rect 36785 47851 36819 47885
rect 36785 47783 36819 47817
rect 36785 47715 36819 47749
rect 36785 47647 36819 47681
rect 36785 47579 36819 47613
rect 36785 47511 36819 47545
rect 36785 47443 36819 47477
rect 37243 48667 37277 48701
rect 37243 48599 37277 48633
rect 37243 48531 37277 48565
rect 37243 48463 37277 48497
rect 37243 48395 37277 48429
rect 37243 48327 37277 48361
rect 37243 48259 37277 48293
rect 37243 48191 37277 48225
rect 37243 48123 37277 48157
rect 37243 48055 37277 48089
rect 37243 47987 37277 48021
rect 37243 47919 37277 47953
rect 37243 47851 37277 47885
rect 37243 47783 37277 47817
rect 37243 47715 37277 47749
rect 37243 47647 37277 47681
rect 37243 47579 37277 47613
rect 37243 47511 37277 47545
rect 37243 47443 37277 47477
rect 37701 48667 37735 48701
rect 37701 48599 37735 48633
rect 37701 48531 37735 48565
rect 37701 48463 37735 48497
rect 37701 48395 37735 48429
rect 37701 48327 37735 48361
rect 37701 48259 37735 48293
rect 37701 48191 37735 48225
rect 37701 48123 37735 48157
rect 37701 48055 37735 48089
rect 37701 47987 37735 48021
rect 37701 47919 37735 47953
rect 37701 47851 37735 47885
rect 37701 47783 37735 47817
rect 37701 47715 37735 47749
rect 37701 47647 37735 47681
rect 37701 47579 37735 47613
rect 37701 47511 37735 47545
rect 37701 47443 37735 47477
rect 38159 48667 38193 48701
rect 38159 48599 38193 48633
rect 38159 48531 38193 48565
rect 38159 48463 38193 48497
rect 38159 48395 38193 48429
rect 38159 48327 38193 48361
rect 38159 48259 38193 48293
rect 38159 48191 38193 48225
rect 38159 48123 38193 48157
rect 38159 48055 38193 48089
rect 38159 47987 38193 48021
rect 38159 47919 38193 47953
rect 38159 47851 38193 47885
rect 38159 47783 38193 47817
rect 38159 47715 38193 47749
rect 38159 47647 38193 47681
rect 38159 47579 38193 47613
rect 38159 47511 38193 47545
rect 38159 47443 38193 47477
rect 38617 48667 38651 48701
rect 38617 48599 38651 48633
rect 38617 48531 38651 48565
rect 38617 48463 38651 48497
rect 38617 48395 38651 48429
rect 38617 48327 38651 48361
rect 38617 48259 38651 48293
rect 38617 48191 38651 48225
rect 38617 48123 38651 48157
rect 38617 48055 38651 48089
rect 38617 47987 38651 48021
rect 38617 47919 38651 47953
rect 38617 47851 38651 47885
rect 38617 47783 38651 47817
rect 38617 47715 38651 47749
rect 38617 47647 38651 47681
rect 38617 47579 38651 47613
rect 38617 47511 38651 47545
rect 38617 47443 38651 47477
rect 39075 48667 39109 48701
rect 39075 48599 39109 48633
rect 39075 48531 39109 48565
rect 39075 48463 39109 48497
rect 39075 48395 39109 48429
rect 39075 48327 39109 48361
rect 39075 48259 39109 48293
rect 39075 48191 39109 48225
rect 39075 48123 39109 48157
rect 39075 48055 39109 48089
rect 39075 47987 39109 48021
rect 39075 47919 39109 47953
rect 39075 47851 39109 47885
rect 39075 47783 39109 47817
rect 39075 47715 39109 47749
rect 39075 47647 39109 47681
rect 39075 47579 39109 47613
rect 39075 47511 39109 47545
rect 39075 47443 39109 47477
rect 39533 48667 39567 48701
rect 39533 48599 39567 48633
rect 39533 48531 39567 48565
rect 39533 48463 39567 48497
rect 39533 48395 39567 48429
rect 39533 48327 39567 48361
rect 39533 48259 39567 48293
rect 39533 48191 39567 48225
rect 39533 48123 39567 48157
rect 39533 48055 39567 48089
rect 39533 47987 39567 48021
rect 39533 47919 39567 47953
rect 39533 47851 39567 47885
rect 39533 47783 39567 47817
rect 39533 47715 39567 47749
rect 39533 47647 39567 47681
rect 39533 47579 39567 47613
rect 39533 47511 39567 47545
rect 39533 47443 39567 47477
rect 39991 48667 40025 48701
rect 39991 48599 40025 48633
rect 39991 48531 40025 48565
rect 39991 48463 40025 48497
rect 39991 48395 40025 48429
rect 39991 48327 40025 48361
rect 39991 48259 40025 48293
rect 39991 48191 40025 48225
rect 39991 48123 40025 48157
rect 39991 48055 40025 48089
rect 39991 47987 40025 48021
rect 39991 47919 40025 47953
rect 39991 47851 40025 47885
rect 39991 47783 40025 47817
rect 39991 47715 40025 47749
rect 39991 47647 40025 47681
rect 39991 47579 40025 47613
rect 39991 47511 40025 47545
rect 39991 47443 40025 47477
rect 40449 48667 40483 48701
rect 40449 48599 40483 48633
rect 40449 48531 40483 48565
rect 40449 48463 40483 48497
rect 40449 48395 40483 48429
rect 40449 48327 40483 48361
rect 40449 48259 40483 48293
rect 40449 48191 40483 48225
rect 40449 48123 40483 48157
rect 40449 48055 40483 48089
rect 40449 47987 40483 48021
rect 40449 47919 40483 47953
rect 40449 47851 40483 47885
rect 40449 47783 40483 47817
rect 40449 47715 40483 47749
rect 40449 47647 40483 47681
rect 40449 47579 40483 47613
rect 40449 47511 40483 47545
rect 40449 47443 40483 47477
rect 40907 48667 40941 48701
rect 40907 48599 40941 48633
rect 40907 48531 40941 48565
rect 40907 48463 40941 48497
rect 40907 48395 40941 48429
rect 40907 48327 40941 48361
rect 40907 48259 40941 48293
rect 40907 48191 40941 48225
rect 40907 48123 40941 48157
rect 40907 48055 40941 48089
rect 40907 47987 40941 48021
rect 40907 47919 40941 47953
rect 40907 47851 40941 47885
rect 40907 47783 40941 47817
rect 40907 47715 40941 47749
rect 40907 47647 40941 47681
rect 40907 47579 40941 47613
rect 40907 47511 40941 47545
rect 40907 47443 40941 47477
rect 41365 48667 41399 48701
rect 41365 48599 41399 48633
rect 41365 48531 41399 48565
rect 41365 48463 41399 48497
rect 41365 48395 41399 48429
rect 41365 48327 41399 48361
rect 41365 48259 41399 48293
rect 41365 48191 41399 48225
rect 41365 48123 41399 48157
rect 41365 48055 41399 48089
rect 41365 47987 41399 48021
rect 41365 47919 41399 47953
rect 41365 47851 41399 47885
rect 41365 47783 41399 47817
rect 41365 47715 41399 47749
rect 41365 47647 41399 47681
rect 41365 47579 41399 47613
rect 41365 47511 41399 47545
rect 41365 47443 41399 47477
rect 41823 48667 41857 48701
rect 41823 48599 41857 48633
rect 41823 48531 41857 48565
rect 41823 48463 41857 48497
rect 41823 48395 41857 48429
rect 41823 48327 41857 48361
rect 41823 48259 41857 48293
rect 41823 48191 41857 48225
rect 41823 48123 41857 48157
rect 41823 48055 41857 48089
rect 41823 47987 41857 48021
rect 41823 47919 41857 47953
rect 41823 47851 41857 47885
rect 41823 47783 41857 47817
rect 41823 47715 41857 47749
rect 41823 47647 41857 47681
rect 41823 47579 41857 47613
rect 41823 47511 41857 47545
rect 41823 47443 41857 47477
rect 42281 48667 42315 48701
rect 42281 48599 42315 48633
rect 42281 48531 42315 48565
rect 42281 48463 42315 48497
rect 42281 48395 42315 48429
rect 42281 48327 42315 48361
rect 42281 48259 42315 48293
rect 42281 48191 42315 48225
rect 42281 48123 42315 48157
rect 42281 48055 42315 48089
rect 42281 47987 42315 48021
rect 42281 47919 42315 47953
rect 42281 47851 42315 47885
rect 42281 47783 42315 47817
rect 42281 47715 42315 47749
rect 42281 47647 42315 47681
rect 42281 47579 42315 47613
rect 42281 47511 42315 47545
rect 42281 47443 42315 47477
rect 42739 48667 42773 48701
rect 42739 48599 42773 48633
rect 42739 48531 42773 48565
rect 42739 48463 42773 48497
rect 42739 48395 42773 48429
rect 42739 48327 42773 48361
rect 42739 48259 42773 48293
rect 42739 48191 42773 48225
rect 42739 48123 42773 48157
rect 42739 48055 42773 48089
rect 42739 47987 42773 48021
rect 42739 47919 42773 47953
rect 42739 47851 42773 47885
rect 42739 47783 42773 47817
rect 42739 47715 42773 47749
rect 42739 47647 42773 47681
rect 42739 47579 42773 47613
rect 42739 47511 42773 47545
rect 42739 47443 42773 47477
rect 43197 48667 43231 48701
rect 43197 48599 43231 48633
rect 43197 48531 43231 48565
rect 43197 48463 43231 48497
rect 43197 48395 43231 48429
rect 43197 48327 43231 48361
rect 43197 48259 43231 48293
rect 43197 48191 43231 48225
rect 43197 48123 43231 48157
rect 43197 48055 43231 48089
rect 43197 47987 43231 48021
rect 43197 47919 43231 47953
rect 43197 47851 43231 47885
rect 43197 47783 43231 47817
rect 43197 47715 43231 47749
rect 43197 47647 43231 47681
rect 43197 47579 43231 47613
rect 43197 47511 43231 47545
rect 43197 47443 43231 47477
rect 43655 48667 43689 48701
rect 43655 48599 43689 48633
rect 43655 48531 43689 48565
rect 43655 48463 43689 48497
rect 43655 48395 43689 48429
rect 43655 48327 43689 48361
rect 43655 48259 43689 48293
rect 43655 48191 43689 48225
rect 43655 48123 43689 48157
rect 43655 48055 43689 48089
rect 43655 47987 43689 48021
rect 43655 47919 43689 47953
rect 43655 47851 43689 47885
rect 43655 47783 43689 47817
rect 43655 47715 43689 47749
rect 43655 47647 43689 47681
rect 43655 47579 43689 47613
rect 43655 47511 43689 47545
rect 43655 47443 43689 47477
rect 44113 48667 44147 48701
rect 44113 48599 44147 48633
rect 44113 48531 44147 48565
rect 44113 48463 44147 48497
rect 44113 48395 44147 48429
rect 44113 48327 44147 48361
rect 44113 48259 44147 48293
rect 44113 48191 44147 48225
rect 44113 48123 44147 48157
rect 44113 48055 44147 48089
rect 44113 47987 44147 48021
rect 44113 47919 44147 47953
rect 44113 47851 44147 47885
rect 44113 47783 44147 47817
rect 44113 47715 44147 47749
rect 44113 47647 44147 47681
rect 44113 47579 44147 47613
rect 44113 47511 44147 47545
rect 44113 47443 44147 47477
rect 44571 48667 44605 48701
rect 44571 48599 44605 48633
rect 44571 48531 44605 48565
rect 44571 48463 44605 48497
rect 44571 48395 44605 48429
rect 44571 48327 44605 48361
rect 44571 48259 44605 48293
rect 44571 48191 44605 48225
rect 44571 48123 44605 48157
rect 44571 48055 44605 48089
rect 44571 47987 44605 48021
rect 44571 47919 44605 47953
rect 44571 47851 44605 47885
rect 44571 47783 44605 47817
rect 44571 47715 44605 47749
rect 44571 47647 44605 47681
rect 44571 47579 44605 47613
rect 44571 47511 44605 47545
rect 44571 47443 44605 47477
rect 45029 48667 45063 48701
rect 45029 48599 45063 48633
rect 45029 48531 45063 48565
rect 45029 48463 45063 48497
rect 45029 48395 45063 48429
rect 45029 48327 45063 48361
rect 45029 48259 45063 48293
rect 45029 48191 45063 48225
rect 45029 48123 45063 48157
rect 45029 48055 45063 48089
rect 45029 47987 45063 48021
rect 45029 47919 45063 47953
rect 45029 47851 45063 47885
rect 45029 47783 45063 47817
rect 45029 47715 45063 47749
rect 45029 47647 45063 47681
rect 45029 47579 45063 47613
rect 45029 47511 45063 47545
rect 45029 47443 45063 47477
rect 45487 48667 45521 48701
rect 45487 48599 45521 48633
rect 45487 48531 45521 48565
rect 45487 48463 45521 48497
rect 45487 48395 45521 48429
rect 45487 48327 45521 48361
rect 45487 48259 45521 48293
rect 45487 48191 45521 48225
rect 45487 48123 45521 48157
rect 45487 48055 45521 48089
rect 45487 47987 45521 48021
rect 45487 47919 45521 47953
rect 45487 47851 45521 47885
rect 45487 47783 45521 47817
rect 45487 47715 45521 47749
rect 45487 47647 45521 47681
rect 45487 47579 45521 47613
rect 45487 47511 45521 47545
rect 45487 47443 45521 47477
rect 45945 48667 45979 48701
rect 45945 48599 45979 48633
rect 45945 48531 45979 48565
rect 45945 48463 45979 48497
rect 45945 48395 45979 48429
rect 45945 48327 45979 48361
rect 45945 48259 45979 48293
rect 45945 48191 45979 48225
rect 45945 48123 45979 48157
rect 45945 48055 45979 48089
rect 45945 47987 45979 48021
rect 45945 47919 45979 47953
rect 45945 47851 45979 47885
rect 45945 47783 45979 47817
rect 45945 47715 45979 47749
rect 45945 47647 45979 47681
rect 45945 47579 45979 47613
rect 45945 47511 45979 47545
rect 45945 47443 45979 47477
rect 46403 48667 46437 48701
rect 46403 48599 46437 48633
rect 46403 48531 46437 48565
rect 46403 48463 46437 48497
rect 46403 48395 46437 48429
rect 46403 48327 46437 48361
rect 46403 48259 46437 48293
rect 46403 48191 46437 48225
rect 46403 48123 46437 48157
rect 46403 48055 46437 48089
rect 46403 47987 46437 48021
rect 46403 47919 46437 47953
rect 46403 47851 46437 47885
rect 46403 47783 46437 47817
rect 46403 47715 46437 47749
rect 46403 47647 46437 47681
rect 46403 47579 46437 47613
rect 46403 47511 46437 47545
rect 46403 47443 46437 47477
rect 46861 48667 46895 48701
rect 46861 48599 46895 48633
rect 46861 48531 46895 48565
rect 46861 48463 46895 48497
rect 46861 48395 46895 48429
rect 46861 48327 46895 48361
rect 46861 48259 46895 48293
rect 46861 48191 46895 48225
rect 46861 48123 46895 48157
rect 46861 48055 46895 48089
rect 46861 47987 46895 48021
rect 46861 47919 46895 47953
rect 46861 47851 46895 47885
rect 46861 47783 46895 47817
rect 46861 47715 46895 47749
rect 46861 47647 46895 47681
rect 46861 47579 46895 47613
rect 46861 47511 46895 47545
rect 46861 47443 46895 47477
rect 47319 48667 47353 48701
rect 47319 48599 47353 48633
rect 47319 48531 47353 48565
rect 47319 48463 47353 48497
rect 47319 48395 47353 48429
rect 47319 48327 47353 48361
rect 47319 48259 47353 48293
rect 47319 48191 47353 48225
rect 47319 48123 47353 48157
rect 47319 48055 47353 48089
rect 47319 47987 47353 48021
rect 47319 47919 47353 47953
rect 47319 47851 47353 47885
rect 47319 47783 47353 47817
rect 47319 47715 47353 47749
rect 47319 47647 47353 47681
rect 47319 47579 47353 47613
rect 47319 47511 47353 47545
rect 47319 47443 47353 47477
rect 47777 48667 47811 48701
rect 47777 48599 47811 48633
rect 47777 48531 47811 48565
rect 47777 48463 47811 48497
rect 47777 48395 47811 48429
rect 47777 48327 47811 48361
rect 47777 48259 47811 48293
rect 47777 48191 47811 48225
rect 47777 48123 47811 48157
rect 47777 48055 47811 48089
rect 47777 47987 47811 48021
rect 47777 47919 47811 47953
rect 47777 47851 47811 47885
rect 47777 47783 47811 47817
rect 47777 47715 47811 47749
rect 47777 47647 47811 47681
rect 47777 47579 47811 47613
rect 47777 47511 47811 47545
rect 47777 47443 47811 47477
rect 48235 48667 48269 48701
rect 48235 48599 48269 48633
rect 48235 48531 48269 48565
rect 48235 48463 48269 48497
rect 48235 48395 48269 48429
rect 48235 48327 48269 48361
rect 48235 48259 48269 48293
rect 48235 48191 48269 48225
rect 48235 48123 48269 48157
rect 48235 48055 48269 48089
rect 48235 47987 48269 48021
rect 48235 47919 48269 47953
rect 48235 47851 48269 47885
rect 48235 47783 48269 47817
rect 48235 47715 48269 47749
rect 48235 47647 48269 47681
rect 48235 47579 48269 47613
rect 48235 47511 48269 47545
rect 48235 47443 48269 47477
rect 48693 48667 48727 48701
rect 48693 48599 48727 48633
rect 48693 48531 48727 48565
rect 48693 48463 48727 48497
rect 48693 48395 48727 48429
rect 48693 48327 48727 48361
rect 48693 48259 48727 48293
rect 48693 48191 48727 48225
rect 48693 48123 48727 48157
rect 48693 48055 48727 48089
rect 48693 47987 48727 48021
rect 48693 47919 48727 47953
rect 48693 47851 48727 47885
rect 48693 47783 48727 47817
rect 48693 47715 48727 47749
rect 48693 47647 48727 47681
rect 48693 47579 48727 47613
rect 48693 47511 48727 47545
rect 48693 47443 48727 47477
rect 49151 48667 49185 48701
rect 49151 48599 49185 48633
rect 49151 48531 49185 48565
rect 49151 48463 49185 48497
rect 49151 48395 49185 48429
rect 49151 48327 49185 48361
rect 49151 48259 49185 48293
rect 49151 48191 49185 48225
rect 49151 48123 49185 48157
rect 49151 48055 49185 48089
rect 49151 47987 49185 48021
rect 49151 47919 49185 47953
rect 49151 47851 49185 47885
rect 49151 47783 49185 47817
rect 49151 47715 49185 47749
rect 49151 47647 49185 47681
rect 49151 47579 49185 47613
rect 49151 47511 49185 47545
rect 49151 47443 49185 47477
rect 49609 48667 49643 48701
rect 49609 48599 49643 48633
rect 49609 48531 49643 48565
rect 49609 48463 49643 48497
rect 49609 48395 49643 48429
rect 49609 48327 49643 48361
rect 49609 48259 49643 48293
rect 49609 48191 49643 48225
rect 49609 48123 49643 48157
rect 49609 48055 49643 48089
rect 49609 47987 49643 48021
rect 49609 47919 49643 47953
rect 49609 47851 49643 47885
rect 49609 47783 49643 47817
rect 49609 47715 49643 47749
rect 49609 47647 49643 47681
rect 49609 47579 49643 47613
rect 49609 47511 49643 47545
rect 49609 47443 49643 47477
rect 50067 48667 50101 48701
rect 50067 48599 50101 48633
rect 50067 48531 50101 48565
rect 50067 48463 50101 48497
rect 50067 48395 50101 48429
rect 50067 48327 50101 48361
rect 50067 48259 50101 48293
rect 50067 48191 50101 48225
rect 50067 48123 50101 48157
rect 50067 48055 50101 48089
rect 50067 47987 50101 48021
rect 50067 47919 50101 47953
rect 50067 47851 50101 47885
rect 50067 47783 50101 47817
rect 50067 47715 50101 47749
rect 50067 47647 50101 47681
rect 50067 47579 50101 47613
rect 50067 47511 50101 47545
rect 50067 47443 50101 47477
rect 50525 48667 50559 48701
rect 50525 48599 50559 48633
rect 50525 48531 50559 48565
rect 50525 48463 50559 48497
rect 50525 48395 50559 48429
rect 50525 48327 50559 48361
rect 50525 48259 50559 48293
rect 50525 48191 50559 48225
rect 50525 48123 50559 48157
rect 50525 48055 50559 48089
rect 50525 47987 50559 48021
rect 50525 47919 50559 47953
rect 50525 47851 50559 47885
rect 50525 47783 50559 47817
rect 50525 47715 50559 47749
rect 50525 47647 50559 47681
rect 50525 47579 50559 47613
rect 50525 47511 50559 47545
rect 50525 47443 50559 47477
rect 50983 48667 51017 48701
rect 50983 48599 51017 48633
rect 50983 48531 51017 48565
rect 50983 48463 51017 48497
rect 50983 48395 51017 48429
rect 50983 48327 51017 48361
rect 50983 48259 51017 48293
rect 50983 48191 51017 48225
rect 50983 48123 51017 48157
rect 50983 48055 51017 48089
rect 50983 47987 51017 48021
rect 50983 47919 51017 47953
rect 50983 47851 51017 47885
rect 50983 47783 51017 47817
rect 50983 47715 51017 47749
rect 50983 47647 51017 47681
rect 50983 47579 51017 47613
rect 50983 47511 51017 47545
rect 50983 47443 51017 47477
rect 51441 48667 51475 48701
rect 51441 48599 51475 48633
rect 51441 48531 51475 48565
rect 51441 48463 51475 48497
rect 51441 48395 51475 48429
rect 51441 48327 51475 48361
rect 51441 48259 51475 48293
rect 51441 48191 51475 48225
rect 51441 48123 51475 48157
rect 51441 48055 51475 48089
rect 51441 47987 51475 48021
rect 51441 47919 51475 47953
rect 51441 47851 51475 47885
rect 51441 47783 51475 47817
rect 51441 47715 51475 47749
rect 51441 47647 51475 47681
rect 51441 47579 51475 47613
rect 51441 47511 51475 47545
rect 51441 47443 51475 47477
rect 51899 48667 51933 48701
rect 51899 48599 51933 48633
rect 51899 48531 51933 48565
rect 51899 48463 51933 48497
rect 51899 48395 51933 48429
rect 51899 48327 51933 48361
rect 51899 48259 51933 48293
rect 51899 48191 51933 48225
rect 51899 48123 51933 48157
rect 51899 48055 51933 48089
rect 51899 47987 51933 48021
rect 51899 47919 51933 47953
rect 51899 47851 51933 47885
rect 51899 47783 51933 47817
rect 51899 47715 51933 47749
rect 51899 47647 51933 47681
rect 51899 47579 51933 47613
rect 51899 47511 51933 47545
rect 51899 47443 51933 47477
rect 52357 48667 52391 48701
rect 52357 48599 52391 48633
rect 52357 48531 52391 48565
rect 52357 48463 52391 48497
rect 52357 48395 52391 48429
rect 52357 48327 52391 48361
rect 52357 48259 52391 48293
rect 52357 48191 52391 48225
rect 52357 48123 52391 48157
rect 52357 48055 52391 48089
rect 52357 47987 52391 48021
rect 52357 47919 52391 47953
rect 52357 47851 52391 47885
rect 52357 47783 52391 47817
rect 52357 47715 52391 47749
rect 52357 47647 52391 47681
rect 52357 47579 52391 47613
rect 52357 47511 52391 47545
rect 52357 47443 52391 47477
rect 15077 44907 15111 44941
rect 15077 44839 15111 44873
rect 15077 44771 15111 44805
rect 15077 44703 15111 44737
rect 15077 44635 15111 44669
rect 15077 44567 15111 44601
rect 15077 44499 15111 44533
rect 15077 44431 15111 44465
rect 15077 44363 15111 44397
rect 15077 44295 15111 44329
rect 15077 44227 15111 44261
rect 15077 44159 15111 44193
rect 15077 44091 15111 44125
rect 15077 44023 15111 44057
rect 15077 43955 15111 43989
rect 15077 43887 15111 43921
rect 15077 43819 15111 43853
rect 15077 43751 15111 43785
rect 15077 43683 15111 43717
rect 15535 44907 15569 44941
rect 15535 44839 15569 44873
rect 15535 44771 15569 44805
rect 15535 44703 15569 44737
rect 15535 44635 15569 44669
rect 15535 44567 15569 44601
rect 15535 44499 15569 44533
rect 15535 44431 15569 44465
rect 15535 44363 15569 44397
rect 15535 44295 15569 44329
rect 15535 44227 15569 44261
rect 15535 44159 15569 44193
rect 15535 44091 15569 44125
rect 15535 44023 15569 44057
rect 15535 43955 15569 43989
rect 15535 43887 15569 43921
rect 15535 43819 15569 43853
rect 15535 43751 15569 43785
rect 15535 43683 15569 43717
rect 15993 44907 16027 44941
rect 15993 44839 16027 44873
rect 15993 44771 16027 44805
rect 15993 44703 16027 44737
rect 15993 44635 16027 44669
rect 15993 44567 16027 44601
rect 15993 44499 16027 44533
rect 15993 44431 16027 44465
rect 15993 44363 16027 44397
rect 15993 44295 16027 44329
rect 15993 44227 16027 44261
rect 15993 44159 16027 44193
rect 15993 44091 16027 44125
rect 15993 44023 16027 44057
rect 15993 43955 16027 43989
rect 15993 43887 16027 43921
rect 15993 43819 16027 43853
rect 15993 43751 16027 43785
rect 15993 43683 16027 43717
rect 16451 44907 16485 44941
rect 16451 44839 16485 44873
rect 16451 44771 16485 44805
rect 16451 44703 16485 44737
rect 16451 44635 16485 44669
rect 16451 44567 16485 44601
rect 16451 44499 16485 44533
rect 16451 44431 16485 44465
rect 16451 44363 16485 44397
rect 16451 44295 16485 44329
rect 16451 44227 16485 44261
rect 16451 44159 16485 44193
rect 16451 44091 16485 44125
rect 16451 44023 16485 44057
rect 16451 43955 16485 43989
rect 16451 43887 16485 43921
rect 16451 43819 16485 43853
rect 16451 43751 16485 43785
rect 16451 43683 16485 43717
rect 16909 44907 16943 44941
rect 16909 44839 16943 44873
rect 16909 44771 16943 44805
rect 16909 44703 16943 44737
rect 16909 44635 16943 44669
rect 16909 44567 16943 44601
rect 16909 44499 16943 44533
rect 16909 44431 16943 44465
rect 16909 44363 16943 44397
rect 16909 44295 16943 44329
rect 16909 44227 16943 44261
rect 16909 44159 16943 44193
rect 16909 44091 16943 44125
rect 16909 44023 16943 44057
rect 16909 43955 16943 43989
rect 16909 43887 16943 43921
rect 16909 43819 16943 43853
rect 16909 43751 16943 43785
rect 16909 43683 16943 43717
rect 17367 44907 17401 44941
rect 17367 44839 17401 44873
rect 17367 44771 17401 44805
rect 17367 44703 17401 44737
rect 17367 44635 17401 44669
rect 17367 44567 17401 44601
rect 17367 44499 17401 44533
rect 17367 44431 17401 44465
rect 17367 44363 17401 44397
rect 17367 44295 17401 44329
rect 17367 44227 17401 44261
rect 17367 44159 17401 44193
rect 17367 44091 17401 44125
rect 17367 44023 17401 44057
rect 17367 43955 17401 43989
rect 17367 43887 17401 43921
rect 17367 43819 17401 43853
rect 17367 43751 17401 43785
rect 17367 43683 17401 43717
rect 17825 44907 17859 44941
rect 17825 44839 17859 44873
rect 17825 44771 17859 44805
rect 17825 44703 17859 44737
rect 17825 44635 17859 44669
rect 17825 44567 17859 44601
rect 17825 44499 17859 44533
rect 17825 44431 17859 44465
rect 17825 44363 17859 44397
rect 17825 44295 17859 44329
rect 17825 44227 17859 44261
rect 17825 44159 17859 44193
rect 17825 44091 17859 44125
rect 17825 44023 17859 44057
rect 17825 43955 17859 43989
rect 17825 43887 17859 43921
rect 17825 43819 17859 43853
rect 17825 43751 17859 43785
rect 17825 43683 17859 43717
rect 18283 44907 18317 44941
rect 18283 44839 18317 44873
rect 18283 44771 18317 44805
rect 18283 44703 18317 44737
rect 18283 44635 18317 44669
rect 18283 44567 18317 44601
rect 18283 44499 18317 44533
rect 18283 44431 18317 44465
rect 18283 44363 18317 44397
rect 18283 44295 18317 44329
rect 18283 44227 18317 44261
rect 18283 44159 18317 44193
rect 18283 44091 18317 44125
rect 18283 44023 18317 44057
rect 18283 43955 18317 43989
rect 18283 43887 18317 43921
rect 18283 43819 18317 43853
rect 18283 43751 18317 43785
rect 18283 43683 18317 43717
rect 18741 44907 18775 44941
rect 18741 44839 18775 44873
rect 18741 44771 18775 44805
rect 18741 44703 18775 44737
rect 18741 44635 18775 44669
rect 18741 44567 18775 44601
rect 18741 44499 18775 44533
rect 18741 44431 18775 44465
rect 18741 44363 18775 44397
rect 18741 44295 18775 44329
rect 18741 44227 18775 44261
rect 18741 44159 18775 44193
rect 18741 44091 18775 44125
rect 18741 44023 18775 44057
rect 18741 43955 18775 43989
rect 18741 43887 18775 43921
rect 18741 43819 18775 43853
rect 18741 43751 18775 43785
rect 18741 43683 18775 43717
rect 19199 44907 19233 44941
rect 19199 44839 19233 44873
rect 19199 44771 19233 44805
rect 19199 44703 19233 44737
rect 19199 44635 19233 44669
rect 19199 44567 19233 44601
rect 19199 44499 19233 44533
rect 19199 44431 19233 44465
rect 19199 44363 19233 44397
rect 19199 44295 19233 44329
rect 19199 44227 19233 44261
rect 19199 44159 19233 44193
rect 19199 44091 19233 44125
rect 19199 44023 19233 44057
rect 19199 43955 19233 43989
rect 19199 43887 19233 43921
rect 19199 43819 19233 43853
rect 19199 43751 19233 43785
rect 19199 43683 19233 43717
rect 19657 44907 19691 44941
rect 19657 44839 19691 44873
rect 19657 44771 19691 44805
rect 19657 44703 19691 44737
rect 19657 44635 19691 44669
rect 19657 44567 19691 44601
rect 19657 44499 19691 44533
rect 19657 44431 19691 44465
rect 19657 44363 19691 44397
rect 19657 44295 19691 44329
rect 19657 44227 19691 44261
rect 19657 44159 19691 44193
rect 19657 44091 19691 44125
rect 19657 44023 19691 44057
rect 19657 43955 19691 43989
rect 19657 43887 19691 43921
rect 19657 43819 19691 43853
rect 19657 43751 19691 43785
rect 19657 43683 19691 43717
rect 20115 44907 20149 44941
rect 20115 44839 20149 44873
rect 20115 44771 20149 44805
rect 20115 44703 20149 44737
rect 20115 44635 20149 44669
rect 20115 44567 20149 44601
rect 20115 44499 20149 44533
rect 20115 44431 20149 44465
rect 20115 44363 20149 44397
rect 20115 44295 20149 44329
rect 20115 44227 20149 44261
rect 20115 44159 20149 44193
rect 20115 44091 20149 44125
rect 20115 44023 20149 44057
rect 20115 43955 20149 43989
rect 20115 43887 20149 43921
rect 20115 43819 20149 43853
rect 20115 43751 20149 43785
rect 20115 43683 20149 43717
rect 20573 44907 20607 44941
rect 20573 44839 20607 44873
rect 20573 44771 20607 44805
rect 20573 44703 20607 44737
rect 20573 44635 20607 44669
rect 20573 44567 20607 44601
rect 20573 44499 20607 44533
rect 20573 44431 20607 44465
rect 20573 44363 20607 44397
rect 20573 44295 20607 44329
rect 20573 44227 20607 44261
rect 20573 44159 20607 44193
rect 20573 44091 20607 44125
rect 20573 44023 20607 44057
rect 20573 43955 20607 43989
rect 20573 43887 20607 43921
rect 20573 43819 20607 43853
rect 20573 43751 20607 43785
rect 20573 43683 20607 43717
rect 21031 44907 21065 44941
rect 21031 44839 21065 44873
rect 21031 44771 21065 44805
rect 21031 44703 21065 44737
rect 21031 44635 21065 44669
rect 21031 44567 21065 44601
rect 21031 44499 21065 44533
rect 21031 44431 21065 44465
rect 21031 44363 21065 44397
rect 21031 44295 21065 44329
rect 21031 44227 21065 44261
rect 21031 44159 21065 44193
rect 21031 44091 21065 44125
rect 21031 44023 21065 44057
rect 21031 43955 21065 43989
rect 21031 43887 21065 43921
rect 21031 43819 21065 43853
rect 21031 43751 21065 43785
rect 21031 43683 21065 43717
rect 21489 44907 21523 44941
rect 21489 44839 21523 44873
rect 21489 44771 21523 44805
rect 21489 44703 21523 44737
rect 21489 44635 21523 44669
rect 21489 44567 21523 44601
rect 21489 44499 21523 44533
rect 21489 44431 21523 44465
rect 21489 44363 21523 44397
rect 21489 44295 21523 44329
rect 21489 44227 21523 44261
rect 21489 44159 21523 44193
rect 21489 44091 21523 44125
rect 21489 44023 21523 44057
rect 21489 43955 21523 43989
rect 21489 43887 21523 43921
rect 21489 43819 21523 43853
rect 21489 43751 21523 43785
rect 21489 43683 21523 43717
rect 21947 44907 21981 44941
rect 21947 44839 21981 44873
rect 21947 44771 21981 44805
rect 21947 44703 21981 44737
rect 21947 44635 21981 44669
rect 21947 44567 21981 44601
rect 21947 44499 21981 44533
rect 21947 44431 21981 44465
rect 21947 44363 21981 44397
rect 21947 44295 21981 44329
rect 21947 44227 21981 44261
rect 21947 44159 21981 44193
rect 21947 44091 21981 44125
rect 21947 44023 21981 44057
rect 21947 43955 21981 43989
rect 21947 43887 21981 43921
rect 21947 43819 21981 43853
rect 21947 43751 21981 43785
rect 21947 43683 21981 43717
rect 22405 44907 22439 44941
rect 22405 44839 22439 44873
rect 22405 44771 22439 44805
rect 22405 44703 22439 44737
rect 22405 44635 22439 44669
rect 22405 44567 22439 44601
rect 22405 44499 22439 44533
rect 22405 44431 22439 44465
rect 22405 44363 22439 44397
rect 22405 44295 22439 44329
rect 22405 44227 22439 44261
rect 22405 44159 22439 44193
rect 22405 44091 22439 44125
rect 22405 44023 22439 44057
rect 22405 43955 22439 43989
rect 22405 43887 22439 43921
rect 22405 43819 22439 43853
rect 22405 43751 22439 43785
rect 22405 43683 22439 43717
rect 22863 44907 22897 44941
rect 22863 44839 22897 44873
rect 22863 44771 22897 44805
rect 22863 44703 22897 44737
rect 22863 44635 22897 44669
rect 22863 44567 22897 44601
rect 22863 44499 22897 44533
rect 22863 44431 22897 44465
rect 22863 44363 22897 44397
rect 22863 44295 22897 44329
rect 22863 44227 22897 44261
rect 22863 44159 22897 44193
rect 22863 44091 22897 44125
rect 22863 44023 22897 44057
rect 22863 43955 22897 43989
rect 22863 43887 22897 43921
rect 22863 43819 22897 43853
rect 22863 43751 22897 43785
rect 22863 43683 22897 43717
rect 23321 44907 23355 44941
rect 23321 44839 23355 44873
rect 23321 44771 23355 44805
rect 23321 44703 23355 44737
rect 23321 44635 23355 44669
rect 23321 44567 23355 44601
rect 23321 44499 23355 44533
rect 23321 44431 23355 44465
rect 23321 44363 23355 44397
rect 23321 44295 23355 44329
rect 23321 44227 23355 44261
rect 23321 44159 23355 44193
rect 23321 44091 23355 44125
rect 23321 44023 23355 44057
rect 23321 43955 23355 43989
rect 23321 43887 23355 43921
rect 23321 43819 23355 43853
rect 23321 43751 23355 43785
rect 23321 43683 23355 43717
rect 23779 44907 23813 44941
rect 23779 44839 23813 44873
rect 23779 44771 23813 44805
rect 23779 44703 23813 44737
rect 23779 44635 23813 44669
rect 23779 44567 23813 44601
rect 23779 44499 23813 44533
rect 23779 44431 23813 44465
rect 23779 44363 23813 44397
rect 23779 44295 23813 44329
rect 23779 44227 23813 44261
rect 23779 44159 23813 44193
rect 23779 44091 23813 44125
rect 23779 44023 23813 44057
rect 23779 43955 23813 43989
rect 23779 43887 23813 43921
rect 23779 43819 23813 43853
rect 23779 43751 23813 43785
rect 23779 43683 23813 43717
rect 24237 44907 24271 44941
rect 24237 44839 24271 44873
rect 24237 44771 24271 44805
rect 24237 44703 24271 44737
rect 24237 44635 24271 44669
rect 24237 44567 24271 44601
rect 24237 44499 24271 44533
rect 24237 44431 24271 44465
rect 24237 44363 24271 44397
rect 24237 44295 24271 44329
rect 24237 44227 24271 44261
rect 24237 44159 24271 44193
rect 24237 44091 24271 44125
rect 24237 44023 24271 44057
rect 24237 43955 24271 43989
rect 24237 43887 24271 43921
rect 24237 43819 24271 43853
rect 24237 43751 24271 43785
rect 24237 43683 24271 43717
rect 24695 44907 24729 44941
rect 24695 44839 24729 44873
rect 24695 44771 24729 44805
rect 24695 44703 24729 44737
rect 24695 44635 24729 44669
rect 24695 44567 24729 44601
rect 24695 44499 24729 44533
rect 24695 44431 24729 44465
rect 24695 44363 24729 44397
rect 24695 44295 24729 44329
rect 24695 44227 24729 44261
rect 24695 44159 24729 44193
rect 24695 44091 24729 44125
rect 24695 44023 24729 44057
rect 24695 43955 24729 43989
rect 24695 43887 24729 43921
rect 24695 43819 24729 43853
rect 24695 43751 24729 43785
rect 24695 43683 24729 43717
rect 25153 44907 25187 44941
rect 25153 44839 25187 44873
rect 25153 44771 25187 44805
rect 25153 44703 25187 44737
rect 25153 44635 25187 44669
rect 25153 44567 25187 44601
rect 25153 44499 25187 44533
rect 25153 44431 25187 44465
rect 25153 44363 25187 44397
rect 25153 44295 25187 44329
rect 25153 44227 25187 44261
rect 25153 44159 25187 44193
rect 25153 44091 25187 44125
rect 25153 44023 25187 44057
rect 25153 43955 25187 43989
rect 25153 43887 25187 43921
rect 25153 43819 25187 43853
rect 25153 43751 25187 43785
rect 25153 43683 25187 43717
rect 25611 44907 25645 44941
rect 25611 44839 25645 44873
rect 25611 44771 25645 44805
rect 25611 44703 25645 44737
rect 25611 44635 25645 44669
rect 25611 44567 25645 44601
rect 25611 44499 25645 44533
rect 25611 44431 25645 44465
rect 25611 44363 25645 44397
rect 25611 44295 25645 44329
rect 25611 44227 25645 44261
rect 25611 44159 25645 44193
rect 25611 44091 25645 44125
rect 25611 44023 25645 44057
rect 25611 43955 25645 43989
rect 25611 43887 25645 43921
rect 25611 43819 25645 43853
rect 25611 43751 25645 43785
rect 25611 43683 25645 43717
rect 26069 44907 26103 44941
rect 26069 44839 26103 44873
rect 26069 44771 26103 44805
rect 26069 44703 26103 44737
rect 26069 44635 26103 44669
rect 26069 44567 26103 44601
rect 26069 44499 26103 44533
rect 26069 44431 26103 44465
rect 26069 44363 26103 44397
rect 26069 44295 26103 44329
rect 26069 44227 26103 44261
rect 26069 44159 26103 44193
rect 26069 44091 26103 44125
rect 26069 44023 26103 44057
rect 26069 43955 26103 43989
rect 26069 43887 26103 43921
rect 26069 43819 26103 43853
rect 26069 43751 26103 43785
rect 26069 43683 26103 43717
rect 26527 44907 26561 44941
rect 26527 44839 26561 44873
rect 26527 44771 26561 44805
rect 26527 44703 26561 44737
rect 26527 44635 26561 44669
rect 26527 44567 26561 44601
rect 26527 44499 26561 44533
rect 26527 44431 26561 44465
rect 26527 44363 26561 44397
rect 26527 44295 26561 44329
rect 26527 44227 26561 44261
rect 26527 44159 26561 44193
rect 26527 44091 26561 44125
rect 26527 44023 26561 44057
rect 26527 43955 26561 43989
rect 26527 43887 26561 43921
rect 26527 43819 26561 43853
rect 26527 43751 26561 43785
rect 26527 43683 26561 43717
rect 26985 44907 27019 44941
rect 26985 44839 27019 44873
rect 26985 44771 27019 44805
rect 26985 44703 27019 44737
rect 26985 44635 27019 44669
rect 26985 44567 27019 44601
rect 26985 44499 27019 44533
rect 26985 44431 27019 44465
rect 26985 44363 27019 44397
rect 26985 44295 27019 44329
rect 26985 44227 27019 44261
rect 26985 44159 27019 44193
rect 26985 44091 27019 44125
rect 26985 44023 27019 44057
rect 26985 43955 27019 43989
rect 26985 43887 27019 43921
rect 26985 43819 27019 43853
rect 26985 43751 27019 43785
rect 26985 43683 27019 43717
rect 27443 44907 27477 44941
rect 27443 44839 27477 44873
rect 27443 44771 27477 44805
rect 27443 44703 27477 44737
rect 27443 44635 27477 44669
rect 27443 44567 27477 44601
rect 27443 44499 27477 44533
rect 27443 44431 27477 44465
rect 27443 44363 27477 44397
rect 27443 44295 27477 44329
rect 27443 44227 27477 44261
rect 27443 44159 27477 44193
rect 27443 44091 27477 44125
rect 27443 44023 27477 44057
rect 27443 43955 27477 43989
rect 27443 43887 27477 43921
rect 27443 43819 27477 43853
rect 27443 43751 27477 43785
rect 27443 43683 27477 43717
rect 27901 44907 27935 44941
rect 27901 44839 27935 44873
rect 27901 44771 27935 44805
rect 27901 44703 27935 44737
rect 27901 44635 27935 44669
rect 27901 44567 27935 44601
rect 27901 44499 27935 44533
rect 27901 44431 27935 44465
rect 27901 44363 27935 44397
rect 27901 44295 27935 44329
rect 27901 44227 27935 44261
rect 27901 44159 27935 44193
rect 27901 44091 27935 44125
rect 27901 44023 27935 44057
rect 27901 43955 27935 43989
rect 27901 43887 27935 43921
rect 27901 43819 27935 43853
rect 27901 43751 27935 43785
rect 27901 43683 27935 43717
rect 28359 44907 28393 44941
rect 28359 44839 28393 44873
rect 28359 44771 28393 44805
rect 28359 44703 28393 44737
rect 28359 44635 28393 44669
rect 28359 44567 28393 44601
rect 28359 44499 28393 44533
rect 28359 44431 28393 44465
rect 28359 44363 28393 44397
rect 28359 44295 28393 44329
rect 28359 44227 28393 44261
rect 28359 44159 28393 44193
rect 28359 44091 28393 44125
rect 28359 44023 28393 44057
rect 28359 43955 28393 43989
rect 28359 43887 28393 43921
rect 28359 43819 28393 43853
rect 28359 43751 28393 43785
rect 28359 43683 28393 43717
rect 28817 44907 28851 44941
rect 28817 44839 28851 44873
rect 28817 44771 28851 44805
rect 28817 44703 28851 44737
rect 28817 44635 28851 44669
rect 28817 44567 28851 44601
rect 28817 44499 28851 44533
rect 28817 44431 28851 44465
rect 28817 44363 28851 44397
rect 28817 44295 28851 44329
rect 28817 44227 28851 44261
rect 28817 44159 28851 44193
rect 28817 44091 28851 44125
rect 28817 44023 28851 44057
rect 28817 43955 28851 43989
rect 28817 43887 28851 43921
rect 28817 43819 28851 43853
rect 28817 43751 28851 43785
rect 28817 43683 28851 43717
rect 29275 44907 29309 44941
rect 29275 44839 29309 44873
rect 29275 44771 29309 44805
rect 29275 44703 29309 44737
rect 29275 44635 29309 44669
rect 29275 44567 29309 44601
rect 29275 44499 29309 44533
rect 29275 44431 29309 44465
rect 29275 44363 29309 44397
rect 29275 44295 29309 44329
rect 29275 44227 29309 44261
rect 29275 44159 29309 44193
rect 29275 44091 29309 44125
rect 29275 44023 29309 44057
rect 29275 43955 29309 43989
rect 29275 43887 29309 43921
rect 29275 43819 29309 43853
rect 29275 43751 29309 43785
rect 29275 43683 29309 43717
rect 29733 44907 29767 44941
rect 29733 44839 29767 44873
rect 29733 44771 29767 44805
rect 29733 44703 29767 44737
rect 29733 44635 29767 44669
rect 29733 44567 29767 44601
rect 29733 44499 29767 44533
rect 29733 44431 29767 44465
rect 29733 44363 29767 44397
rect 29733 44295 29767 44329
rect 29733 44227 29767 44261
rect 29733 44159 29767 44193
rect 29733 44091 29767 44125
rect 29733 44023 29767 44057
rect 29733 43955 29767 43989
rect 29733 43887 29767 43921
rect 29733 43819 29767 43853
rect 29733 43751 29767 43785
rect 29733 43683 29767 43717
rect 30191 44907 30225 44941
rect 30191 44839 30225 44873
rect 30191 44771 30225 44805
rect 30191 44703 30225 44737
rect 30191 44635 30225 44669
rect 30191 44567 30225 44601
rect 30191 44499 30225 44533
rect 30191 44431 30225 44465
rect 30191 44363 30225 44397
rect 30191 44295 30225 44329
rect 30191 44227 30225 44261
rect 30191 44159 30225 44193
rect 30191 44091 30225 44125
rect 30191 44023 30225 44057
rect 30191 43955 30225 43989
rect 30191 43887 30225 43921
rect 30191 43819 30225 43853
rect 30191 43751 30225 43785
rect 30191 43683 30225 43717
rect 30649 44907 30683 44941
rect 30649 44839 30683 44873
rect 30649 44771 30683 44805
rect 30649 44703 30683 44737
rect 30649 44635 30683 44669
rect 30649 44567 30683 44601
rect 30649 44499 30683 44533
rect 30649 44431 30683 44465
rect 30649 44363 30683 44397
rect 30649 44295 30683 44329
rect 30649 44227 30683 44261
rect 30649 44159 30683 44193
rect 30649 44091 30683 44125
rect 30649 44023 30683 44057
rect 30649 43955 30683 43989
rect 30649 43887 30683 43921
rect 30649 43819 30683 43853
rect 30649 43751 30683 43785
rect 30649 43683 30683 43717
rect 31107 44907 31141 44941
rect 31107 44839 31141 44873
rect 31107 44771 31141 44805
rect 31107 44703 31141 44737
rect 31107 44635 31141 44669
rect 31107 44567 31141 44601
rect 31107 44499 31141 44533
rect 31107 44431 31141 44465
rect 31107 44363 31141 44397
rect 31107 44295 31141 44329
rect 31107 44227 31141 44261
rect 31107 44159 31141 44193
rect 31107 44091 31141 44125
rect 31107 44023 31141 44057
rect 31107 43955 31141 43989
rect 31107 43887 31141 43921
rect 31107 43819 31141 43853
rect 31107 43751 31141 43785
rect 31107 43683 31141 43717
rect 31565 44907 31599 44941
rect 31565 44839 31599 44873
rect 31565 44771 31599 44805
rect 31565 44703 31599 44737
rect 31565 44635 31599 44669
rect 31565 44567 31599 44601
rect 31565 44499 31599 44533
rect 31565 44431 31599 44465
rect 31565 44363 31599 44397
rect 31565 44295 31599 44329
rect 31565 44227 31599 44261
rect 31565 44159 31599 44193
rect 31565 44091 31599 44125
rect 31565 44023 31599 44057
rect 31565 43955 31599 43989
rect 31565 43887 31599 43921
rect 31565 43819 31599 43853
rect 31565 43751 31599 43785
rect 31565 43683 31599 43717
rect 32023 44907 32057 44941
rect 32023 44839 32057 44873
rect 32023 44771 32057 44805
rect 32023 44703 32057 44737
rect 32023 44635 32057 44669
rect 32023 44567 32057 44601
rect 32023 44499 32057 44533
rect 32023 44431 32057 44465
rect 32023 44363 32057 44397
rect 32023 44295 32057 44329
rect 32023 44227 32057 44261
rect 32023 44159 32057 44193
rect 32023 44091 32057 44125
rect 32023 44023 32057 44057
rect 32023 43955 32057 43989
rect 32023 43887 32057 43921
rect 32023 43819 32057 43853
rect 32023 43751 32057 43785
rect 32023 43683 32057 43717
rect 32481 44907 32515 44941
rect 32481 44839 32515 44873
rect 32481 44771 32515 44805
rect 32481 44703 32515 44737
rect 32481 44635 32515 44669
rect 32481 44567 32515 44601
rect 32481 44499 32515 44533
rect 32481 44431 32515 44465
rect 32481 44363 32515 44397
rect 32481 44295 32515 44329
rect 32481 44227 32515 44261
rect 32481 44159 32515 44193
rect 32481 44091 32515 44125
rect 32481 44023 32515 44057
rect 32481 43955 32515 43989
rect 32481 43887 32515 43921
rect 32481 43819 32515 43853
rect 32481 43751 32515 43785
rect 32481 43683 32515 43717
rect 32939 44907 32973 44941
rect 32939 44839 32973 44873
rect 32939 44771 32973 44805
rect 32939 44703 32973 44737
rect 32939 44635 32973 44669
rect 32939 44567 32973 44601
rect 32939 44499 32973 44533
rect 32939 44431 32973 44465
rect 32939 44363 32973 44397
rect 32939 44295 32973 44329
rect 32939 44227 32973 44261
rect 32939 44159 32973 44193
rect 32939 44091 32973 44125
rect 32939 44023 32973 44057
rect 32939 43955 32973 43989
rect 32939 43887 32973 43921
rect 32939 43819 32973 43853
rect 32939 43751 32973 43785
rect 32939 43683 32973 43717
rect 33397 44907 33431 44941
rect 33397 44839 33431 44873
rect 33397 44771 33431 44805
rect 33397 44703 33431 44737
rect 33397 44635 33431 44669
rect 33397 44567 33431 44601
rect 33397 44499 33431 44533
rect 33397 44431 33431 44465
rect 33397 44363 33431 44397
rect 33397 44295 33431 44329
rect 33397 44227 33431 44261
rect 33397 44159 33431 44193
rect 33397 44091 33431 44125
rect 33397 44023 33431 44057
rect 33397 43955 33431 43989
rect 33397 43887 33431 43921
rect 33397 43819 33431 43853
rect 33397 43751 33431 43785
rect 33397 43683 33431 43717
rect 33855 44907 33889 44941
rect 33855 44839 33889 44873
rect 33855 44771 33889 44805
rect 33855 44703 33889 44737
rect 33855 44635 33889 44669
rect 33855 44567 33889 44601
rect 33855 44499 33889 44533
rect 33855 44431 33889 44465
rect 33855 44363 33889 44397
rect 33855 44295 33889 44329
rect 33855 44227 33889 44261
rect 33855 44159 33889 44193
rect 33855 44091 33889 44125
rect 33855 44023 33889 44057
rect 33855 43955 33889 43989
rect 33855 43887 33889 43921
rect 33855 43819 33889 43853
rect 33855 43751 33889 43785
rect 33855 43683 33889 43717
rect 34313 44907 34347 44941
rect 34313 44839 34347 44873
rect 34313 44771 34347 44805
rect 34313 44703 34347 44737
rect 34313 44635 34347 44669
rect 34313 44567 34347 44601
rect 34313 44499 34347 44533
rect 34313 44431 34347 44465
rect 34313 44363 34347 44397
rect 34313 44295 34347 44329
rect 34313 44227 34347 44261
rect 34313 44159 34347 44193
rect 34313 44091 34347 44125
rect 34313 44023 34347 44057
rect 34313 43955 34347 43989
rect 34313 43887 34347 43921
rect 34313 43819 34347 43853
rect 34313 43751 34347 43785
rect 34313 43683 34347 43717
rect 34771 44907 34805 44941
rect 34771 44839 34805 44873
rect 34771 44771 34805 44805
rect 34771 44703 34805 44737
rect 34771 44635 34805 44669
rect 34771 44567 34805 44601
rect 34771 44499 34805 44533
rect 34771 44431 34805 44465
rect 34771 44363 34805 44397
rect 34771 44295 34805 44329
rect 34771 44227 34805 44261
rect 34771 44159 34805 44193
rect 34771 44091 34805 44125
rect 34771 44023 34805 44057
rect 34771 43955 34805 43989
rect 34771 43887 34805 43921
rect 34771 43819 34805 43853
rect 34771 43751 34805 43785
rect 34771 43683 34805 43717
rect 35229 44907 35263 44941
rect 35229 44839 35263 44873
rect 35229 44771 35263 44805
rect 35229 44703 35263 44737
rect 35229 44635 35263 44669
rect 35229 44567 35263 44601
rect 35229 44499 35263 44533
rect 35229 44431 35263 44465
rect 35229 44363 35263 44397
rect 35229 44295 35263 44329
rect 35229 44227 35263 44261
rect 35229 44159 35263 44193
rect 35229 44091 35263 44125
rect 35229 44023 35263 44057
rect 35229 43955 35263 43989
rect 35229 43887 35263 43921
rect 35229 43819 35263 43853
rect 35229 43751 35263 43785
rect 35229 43683 35263 43717
rect 35687 44907 35721 44941
rect 35687 44839 35721 44873
rect 35687 44771 35721 44805
rect 35687 44703 35721 44737
rect 35687 44635 35721 44669
rect 35687 44567 35721 44601
rect 35687 44499 35721 44533
rect 35687 44431 35721 44465
rect 35687 44363 35721 44397
rect 35687 44295 35721 44329
rect 35687 44227 35721 44261
rect 35687 44159 35721 44193
rect 35687 44091 35721 44125
rect 35687 44023 35721 44057
rect 35687 43955 35721 43989
rect 35687 43887 35721 43921
rect 35687 43819 35721 43853
rect 35687 43751 35721 43785
rect 35687 43683 35721 43717
rect 36145 44907 36179 44941
rect 36145 44839 36179 44873
rect 36145 44771 36179 44805
rect 36145 44703 36179 44737
rect 36145 44635 36179 44669
rect 36145 44567 36179 44601
rect 36145 44499 36179 44533
rect 36145 44431 36179 44465
rect 36145 44363 36179 44397
rect 36145 44295 36179 44329
rect 36145 44227 36179 44261
rect 36145 44159 36179 44193
rect 36145 44091 36179 44125
rect 36145 44023 36179 44057
rect 36145 43955 36179 43989
rect 36145 43887 36179 43921
rect 36145 43819 36179 43853
rect 36145 43751 36179 43785
rect 36145 43683 36179 43717
rect 36603 44907 36637 44941
rect 36603 44839 36637 44873
rect 36603 44771 36637 44805
rect 36603 44703 36637 44737
rect 36603 44635 36637 44669
rect 36603 44567 36637 44601
rect 36603 44499 36637 44533
rect 36603 44431 36637 44465
rect 36603 44363 36637 44397
rect 36603 44295 36637 44329
rect 36603 44227 36637 44261
rect 36603 44159 36637 44193
rect 36603 44091 36637 44125
rect 36603 44023 36637 44057
rect 36603 43955 36637 43989
rect 36603 43887 36637 43921
rect 36603 43819 36637 43853
rect 36603 43751 36637 43785
rect 36603 43683 36637 43717
rect 37061 44907 37095 44941
rect 37061 44839 37095 44873
rect 37061 44771 37095 44805
rect 37061 44703 37095 44737
rect 37061 44635 37095 44669
rect 37061 44567 37095 44601
rect 37061 44499 37095 44533
rect 37061 44431 37095 44465
rect 37061 44363 37095 44397
rect 37061 44295 37095 44329
rect 37061 44227 37095 44261
rect 37061 44159 37095 44193
rect 37061 44091 37095 44125
rect 37061 44023 37095 44057
rect 37061 43955 37095 43989
rect 37061 43887 37095 43921
rect 37061 43819 37095 43853
rect 37061 43751 37095 43785
rect 37061 43683 37095 43717
rect 37519 44907 37553 44941
rect 37519 44839 37553 44873
rect 37519 44771 37553 44805
rect 37519 44703 37553 44737
rect 37519 44635 37553 44669
rect 37519 44567 37553 44601
rect 37519 44499 37553 44533
rect 37519 44431 37553 44465
rect 37519 44363 37553 44397
rect 37519 44295 37553 44329
rect 37519 44227 37553 44261
rect 37519 44159 37553 44193
rect 37519 44091 37553 44125
rect 37519 44023 37553 44057
rect 37519 43955 37553 43989
rect 37519 43887 37553 43921
rect 37519 43819 37553 43853
rect 37519 43751 37553 43785
rect 37519 43683 37553 43717
rect 37977 44907 38011 44941
rect 37977 44839 38011 44873
rect 37977 44771 38011 44805
rect 37977 44703 38011 44737
rect 37977 44635 38011 44669
rect 37977 44567 38011 44601
rect 37977 44499 38011 44533
rect 37977 44431 38011 44465
rect 37977 44363 38011 44397
rect 37977 44295 38011 44329
rect 37977 44227 38011 44261
rect 37977 44159 38011 44193
rect 37977 44091 38011 44125
rect 37977 44023 38011 44057
rect 37977 43955 38011 43989
rect 37977 43887 38011 43921
rect 37977 43819 38011 43853
rect 37977 43751 38011 43785
rect 37977 43683 38011 43717
rect 38435 44907 38469 44941
rect 38435 44839 38469 44873
rect 38435 44771 38469 44805
rect 38435 44703 38469 44737
rect 38435 44635 38469 44669
rect 38435 44567 38469 44601
rect 38435 44499 38469 44533
rect 38435 44431 38469 44465
rect 38435 44363 38469 44397
rect 38435 44295 38469 44329
rect 38435 44227 38469 44261
rect 38435 44159 38469 44193
rect 38435 44091 38469 44125
rect 38435 44023 38469 44057
rect 38435 43955 38469 43989
rect 38435 43887 38469 43921
rect 38435 43819 38469 43853
rect 38435 43751 38469 43785
rect 38435 43683 38469 43717
rect 38893 44907 38927 44941
rect 38893 44839 38927 44873
rect 38893 44771 38927 44805
rect 38893 44703 38927 44737
rect 38893 44635 38927 44669
rect 38893 44567 38927 44601
rect 38893 44499 38927 44533
rect 38893 44431 38927 44465
rect 38893 44363 38927 44397
rect 38893 44295 38927 44329
rect 38893 44227 38927 44261
rect 38893 44159 38927 44193
rect 38893 44091 38927 44125
rect 38893 44023 38927 44057
rect 38893 43955 38927 43989
rect 38893 43887 38927 43921
rect 38893 43819 38927 43853
rect 38893 43751 38927 43785
rect 38893 43683 38927 43717
rect 39351 44907 39385 44941
rect 39351 44839 39385 44873
rect 39351 44771 39385 44805
rect 39351 44703 39385 44737
rect 39351 44635 39385 44669
rect 39351 44567 39385 44601
rect 39351 44499 39385 44533
rect 39351 44431 39385 44465
rect 39351 44363 39385 44397
rect 39351 44295 39385 44329
rect 39351 44227 39385 44261
rect 39351 44159 39385 44193
rect 39351 44091 39385 44125
rect 39351 44023 39385 44057
rect 39351 43955 39385 43989
rect 39351 43887 39385 43921
rect 39351 43819 39385 43853
rect 39351 43751 39385 43785
rect 39351 43683 39385 43717
rect 39809 44907 39843 44941
rect 39809 44839 39843 44873
rect 39809 44771 39843 44805
rect 39809 44703 39843 44737
rect 39809 44635 39843 44669
rect 39809 44567 39843 44601
rect 39809 44499 39843 44533
rect 39809 44431 39843 44465
rect 39809 44363 39843 44397
rect 39809 44295 39843 44329
rect 39809 44227 39843 44261
rect 39809 44159 39843 44193
rect 39809 44091 39843 44125
rect 39809 44023 39843 44057
rect 39809 43955 39843 43989
rect 39809 43887 39843 43921
rect 39809 43819 39843 43853
rect 39809 43751 39843 43785
rect 39809 43683 39843 43717
rect 40267 44907 40301 44941
rect 40267 44839 40301 44873
rect 40267 44771 40301 44805
rect 40267 44703 40301 44737
rect 40267 44635 40301 44669
rect 40267 44567 40301 44601
rect 40267 44499 40301 44533
rect 40267 44431 40301 44465
rect 40267 44363 40301 44397
rect 40267 44295 40301 44329
rect 40267 44227 40301 44261
rect 40267 44159 40301 44193
rect 40267 44091 40301 44125
rect 40267 44023 40301 44057
rect 40267 43955 40301 43989
rect 40267 43887 40301 43921
rect 40267 43819 40301 43853
rect 40267 43751 40301 43785
rect 40267 43683 40301 43717
rect 40725 44907 40759 44941
rect 40725 44839 40759 44873
rect 40725 44771 40759 44805
rect 40725 44703 40759 44737
rect 40725 44635 40759 44669
rect 40725 44567 40759 44601
rect 40725 44499 40759 44533
rect 40725 44431 40759 44465
rect 40725 44363 40759 44397
rect 40725 44295 40759 44329
rect 40725 44227 40759 44261
rect 40725 44159 40759 44193
rect 40725 44091 40759 44125
rect 40725 44023 40759 44057
rect 40725 43955 40759 43989
rect 40725 43887 40759 43921
rect 40725 43819 40759 43853
rect 40725 43751 40759 43785
rect 40725 43683 40759 43717
rect 41183 44907 41217 44941
rect 41183 44839 41217 44873
rect 41183 44771 41217 44805
rect 41183 44703 41217 44737
rect 41183 44635 41217 44669
rect 41183 44567 41217 44601
rect 41183 44499 41217 44533
rect 41183 44431 41217 44465
rect 41183 44363 41217 44397
rect 41183 44295 41217 44329
rect 41183 44227 41217 44261
rect 41183 44159 41217 44193
rect 41183 44091 41217 44125
rect 41183 44023 41217 44057
rect 41183 43955 41217 43989
rect 41183 43887 41217 43921
rect 41183 43819 41217 43853
rect 41183 43751 41217 43785
rect 41183 43683 41217 43717
rect 41641 44907 41675 44941
rect 41641 44839 41675 44873
rect 41641 44771 41675 44805
rect 41641 44703 41675 44737
rect 41641 44635 41675 44669
rect 41641 44567 41675 44601
rect 41641 44499 41675 44533
rect 41641 44431 41675 44465
rect 41641 44363 41675 44397
rect 41641 44295 41675 44329
rect 41641 44227 41675 44261
rect 41641 44159 41675 44193
rect 41641 44091 41675 44125
rect 41641 44023 41675 44057
rect 41641 43955 41675 43989
rect 41641 43887 41675 43921
rect 41641 43819 41675 43853
rect 41641 43751 41675 43785
rect 41641 43683 41675 43717
rect 42099 44907 42133 44941
rect 42099 44839 42133 44873
rect 42099 44771 42133 44805
rect 42099 44703 42133 44737
rect 42099 44635 42133 44669
rect 42099 44567 42133 44601
rect 42099 44499 42133 44533
rect 42099 44431 42133 44465
rect 42099 44363 42133 44397
rect 42099 44295 42133 44329
rect 42099 44227 42133 44261
rect 42099 44159 42133 44193
rect 42099 44091 42133 44125
rect 42099 44023 42133 44057
rect 42099 43955 42133 43989
rect 42099 43887 42133 43921
rect 42099 43819 42133 43853
rect 42099 43751 42133 43785
rect 42099 43683 42133 43717
rect 42557 44907 42591 44941
rect 42557 44839 42591 44873
rect 42557 44771 42591 44805
rect 42557 44703 42591 44737
rect 42557 44635 42591 44669
rect 42557 44567 42591 44601
rect 42557 44499 42591 44533
rect 42557 44431 42591 44465
rect 42557 44363 42591 44397
rect 42557 44295 42591 44329
rect 42557 44227 42591 44261
rect 42557 44159 42591 44193
rect 42557 44091 42591 44125
rect 42557 44023 42591 44057
rect 42557 43955 42591 43989
rect 42557 43887 42591 43921
rect 42557 43819 42591 43853
rect 42557 43751 42591 43785
rect 42557 43683 42591 43717
rect 43344 44506 43378 44540
rect 43434 44506 43468 44540
rect 43524 44506 43558 44540
rect 43614 44506 43648 44540
rect 43704 44506 43738 44540
rect 43794 44506 43828 44540
rect 43884 44506 43918 44540
rect 43344 44416 43378 44450
rect 43434 44416 43468 44450
rect 43524 44416 43558 44450
rect 43614 44416 43648 44450
rect 43704 44416 43738 44450
rect 43794 44416 43828 44450
rect 43884 44416 43918 44450
rect 43344 44326 43378 44360
rect 43434 44326 43468 44360
rect 43524 44326 43558 44360
rect 43614 44326 43648 44360
rect 43704 44326 43738 44360
rect 43794 44326 43828 44360
rect 43884 44326 43918 44360
rect 43344 44236 43378 44270
rect 43434 44236 43468 44270
rect 43524 44236 43558 44270
rect 43614 44236 43648 44270
rect 43704 44236 43738 44270
rect 43794 44236 43828 44270
rect 43884 44236 43918 44270
rect 43344 44146 43378 44180
rect 43434 44146 43468 44180
rect 43524 44146 43558 44180
rect 43614 44146 43648 44180
rect 43704 44146 43738 44180
rect 43794 44146 43828 44180
rect 43884 44146 43918 44180
rect 43344 44056 43378 44090
rect 43434 44056 43468 44090
rect 43524 44056 43558 44090
rect 43614 44056 43648 44090
rect 43704 44056 43738 44090
rect 43794 44056 43828 44090
rect 43884 44056 43918 44090
rect 43344 43966 43378 44000
rect 43434 43966 43468 44000
rect 43524 43966 43558 44000
rect 43614 43966 43648 44000
rect 43704 43966 43738 44000
rect 43794 43966 43828 44000
rect 43884 43966 43918 44000
rect 44684 44506 44718 44540
rect 44774 44506 44808 44540
rect 44864 44506 44898 44540
rect 44954 44506 44988 44540
rect 45044 44506 45078 44540
rect 45134 44506 45168 44540
rect 45224 44506 45258 44540
rect 44684 44416 44718 44450
rect 44774 44416 44808 44450
rect 44864 44416 44898 44450
rect 44954 44416 44988 44450
rect 45044 44416 45078 44450
rect 45134 44416 45168 44450
rect 45224 44416 45258 44450
rect 44684 44326 44718 44360
rect 44774 44326 44808 44360
rect 44864 44326 44898 44360
rect 44954 44326 44988 44360
rect 45044 44326 45078 44360
rect 45134 44326 45168 44360
rect 45224 44326 45258 44360
rect 44684 44236 44718 44270
rect 44774 44236 44808 44270
rect 44864 44236 44898 44270
rect 44954 44236 44988 44270
rect 45044 44236 45078 44270
rect 45134 44236 45168 44270
rect 45224 44236 45258 44270
rect 44684 44146 44718 44180
rect 44774 44146 44808 44180
rect 44864 44146 44898 44180
rect 44954 44146 44988 44180
rect 45044 44146 45078 44180
rect 45134 44146 45168 44180
rect 45224 44146 45258 44180
rect 44684 44056 44718 44090
rect 44774 44056 44808 44090
rect 44864 44056 44898 44090
rect 44954 44056 44988 44090
rect 45044 44056 45078 44090
rect 45134 44056 45168 44090
rect 45224 44056 45258 44090
rect 44684 43966 44718 44000
rect 44774 43966 44808 44000
rect 44864 43966 44898 44000
rect 44954 43966 44988 44000
rect 45044 43966 45078 44000
rect 45134 43966 45168 44000
rect 45224 43966 45258 44000
rect 46024 44506 46058 44540
rect 46114 44506 46148 44540
rect 46204 44506 46238 44540
rect 46294 44506 46328 44540
rect 46384 44506 46418 44540
rect 46474 44506 46508 44540
rect 46564 44506 46598 44540
rect 46024 44416 46058 44450
rect 46114 44416 46148 44450
rect 46204 44416 46238 44450
rect 46294 44416 46328 44450
rect 46384 44416 46418 44450
rect 46474 44416 46508 44450
rect 46564 44416 46598 44450
rect 46024 44326 46058 44360
rect 46114 44326 46148 44360
rect 46204 44326 46238 44360
rect 46294 44326 46328 44360
rect 46384 44326 46418 44360
rect 46474 44326 46508 44360
rect 46564 44326 46598 44360
rect 46024 44236 46058 44270
rect 46114 44236 46148 44270
rect 46204 44236 46238 44270
rect 46294 44236 46328 44270
rect 46384 44236 46418 44270
rect 46474 44236 46508 44270
rect 46564 44236 46598 44270
rect 46024 44146 46058 44180
rect 46114 44146 46148 44180
rect 46204 44146 46238 44180
rect 46294 44146 46328 44180
rect 46384 44146 46418 44180
rect 46474 44146 46508 44180
rect 46564 44146 46598 44180
rect 46024 44056 46058 44090
rect 46114 44056 46148 44090
rect 46204 44056 46238 44090
rect 46294 44056 46328 44090
rect 46384 44056 46418 44090
rect 46474 44056 46508 44090
rect 46564 44056 46598 44090
rect 46024 43966 46058 44000
rect 46114 43966 46148 44000
rect 46204 43966 46238 44000
rect 46294 43966 46328 44000
rect 46384 43966 46418 44000
rect 46474 43966 46508 44000
rect 46564 43966 46598 44000
rect 47364 44506 47398 44540
rect 47454 44506 47488 44540
rect 47544 44506 47578 44540
rect 47634 44506 47668 44540
rect 47724 44506 47758 44540
rect 47814 44506 47848 44540
rect 47904 44506 47938 44540
rect 47364 44416 47398 44450
rect 47454 44416 47488 44450
rect 47544 44416 47578 44450
rect 47634 44416 47668 44450
rect 47724 44416 47758 44450
rect 47814 44416 47848 44450
rect 47904 44416 47938 44450
rect 47364 44326 47398 44360
rect 47454 44326 47488 44360
rect 47544 44326 47578 44360
rect 47634 44326 47668 44360
rect 47724 44326 47758 44360
rect 47814 44326 47848 44360
rect 47904 44326 47938 44360
rect 47364 44236 47398 44270
rect 47454 44236 47488 44270
rect 47544 44236 47578 44270
rect 47634 44236 47668 44270
rect 47724 44236 47758 44270
rect 47814 44236 47848 44270
rect 47904 44236 47938 44270
rect 47364 44146 47398 44180
rect 47454 44146 47488 44180
rect 47544 44146 47578 44180
rect 47634 44146 47668 44180
rect 47724 44146 47758 44180
rect 47814 44146 47848 44180
rect 47904 44146 47938 44180
rect 47364 44056 47398 44090
rect 47454 44056 47488 44090
rect 47544 44056 47578 44090
rect 47634 44056 47668 44090
rect 47724 44056 47758 44090
rect 47814 44056 47848 44090
rect 47904 44056 47938 44090
rect 47364 43966 47398 44000
rect 47454 43966 47488 44000
rect 47544 43966 47578 44000
rect 47634 43966 47668 44000
rect 47724 43966 47758 44000
rect 47814 43966 47848 44000
rect 47904 43966 47938 44000
rect 48704 44506 48738 44540
rect 48794 44506 48828 44540
rect 48884 44506 48918 44540
rect 48974 44506 49008 44540
rect 49064 44506 49098 44540
rect 49154 44506 49188 44540
rect 49244 44506 49278 44540
rect 48704 44416 48738 44450
rect 48794 44416 48828 44450
rect 48884 44416 48918 44450
rect 48974 44416 49008 44450
rect 49064 44416 49098 44450
rect 49154 44416 49188 44450
rect 49244 44416 49278 44450
rect 48704 44326 48738 44360
rect 48794 44326 48828 44360
rect 48884 44326 48918 44360
rect 48974 44326 49008 44360
rect 49064 44326 49098 44360
rect 49154 44326 49188 44360
rect 49244 44326 49278 44360
rect 48704 44236 48738 44270
rect 48794 44236 48828 44270
rect 48884 44236 48918 44270
rect 48974 44236 49008 44270
rect 49064 44236 49098 44270
rect 49154 44236 49188 44270
rect 49244 44236 49278 44270
rect 48704 44146 48738 44180
rect 48794 44146 48828 44180
rect 48884 44146 48918 44180
rect 48974 44146 49008 44180
rect 49064 44146 49098 44180
rect 49154 44146 49188 44180
rect 49244 44146 49278 44180
rect 48704 44056 48738 44090
rect 48794 44056 48828 44090
rect 48884 44056 48918 44090
rect 48974 44056 49008 44090
rect 49064 44056 49098 44090
rect 49154 44056 49188 44090
rect 49244 44056 49278 44090
rect 48704 43966 48738 44000
rect 48794 43966 48828 44000
rect 48884 43966 48918 44000
rect 48974 43966 49008 44000
rect 49064 43966 49098 44000
rect 49154 43966 49188 44000
rect 49244 43966 49278 44000
rect 50044 44506 50078 44540
rect 50134 44506 50168 44540
rect 50224 44506 50258 44540
rect 50314 44506 50348 44540
rect 50404 44506 50438 44540
rect 50494 44506 50528 44540
rect 50584 44506 50618 44540
rect 50044 44416 50078 44450
rect 50134 44416 50168 44450
rect 50224 44416 50258 44450
rect 50314 44416 50348 44450
rect 50404 44416 50438 44450
rect 50494 44416 50528 44450
rect 50584 44416 50618 44450
rect 50044 44326 50078 44360
rect 50134 44326 50168 44360
rect 50224 44326 50258 44360
rect 50314 44326 50348 44360
rect 50404 44326 50438 44360
rect 50494 44326 50528 44360
rect 50584 44326 50618 44360
rect 50044 44236 50078 44270
rect 50134 44236 50168 44270
rect 50224 44236 50258 44270
rect 50314 44236 50348 44270
rect 50404 44236 50438 44270
rect 50494 44236 50528 44270
rect 50584 44236 50618 44270
rect 50044 44146 50078 44180
rect 50134 44146 50168 44180
rect 50224 44146 50258 44180
rect 50314 44146 50348 44180
rect 50404 44146 50438 44180
rect 50494 44146 50528 44180
rect 50584 44146 50618 44180
rect 50044 44056 50078 44090
rect 50134 44056 50168 44090
rect 50224 44056 50258 44090
rect 50314 44056 50348 44090
rect 50404 44056 50438 44090
rect 50494 44056 50528 44090
rect 50584 44056 50618 44090
rect 50044 43966 50078 44000
rect 50134 43966 50168 44000
rect 50224 43966 50258 44000
rect 50314 43966 50348 44000
rect 50404 43966 50438 44000
rect 50494 43966 50528 44000
rect 50584 43966 50618 44000
rect 51384 44506 51418 44540
rect 51474 44506 51508 44540
rect 51564 44506 51598 44540
rect 51654 44506 51688 44540
rect 51744 44506 51778 44540
rect 51834 44506 51868 44540
rect 51924 44506 51958 44540
rect 51384 44416 51418 44450
rect 51474 44416 51508 44450
rect 51564 44416 51598 44450
rect 51654 44416 51688 44450
rect 51744 44416 51778 44450
rect 51834 44416 51868 44450
rect 51924 44416 51958 44450
rect 51384 44326 51418 44360
rect 51474 44326 51508 44360
rect 51564 44326 51598 44360
rect 51654 44326 51688 44360
rect 51744 44326 51778 44360
rect 51834 44326 51868 44360
rect 51924 44326 51958 44360
rect 51384 44236 51418 44270
rect 51474 44236 51508 44270
rect 51564 44236 51598 44270
rect 51654 44236 51688 44270
rect 51744 44236 51778 44270
rect 51834 44236 51868 44270
rect 51924 44236 51958 44270
rect 51384 44146 51418 44180
rect 51474 44146 51508 44180
rect 51564 44146 51598 44180
rect 51654 44146 51688 44180
rect 51744 44146 51778 44180
rect 51834 44146 51868 44180
rect 51924 44146 51958 44180
rect 51384 44056 51418 44090
rect 51474 44056 51508 44090
rect 51564 44056 51598 44090
rect 51654 44056 51688 44090
rect 51744 44056 51778 44090
rect 51834 44056 51868 44090
rect 51924 44056 51958 44090
rect 51384 43966 51418 44000
rect 51474 43966 51508 44000
rect 51564 43966 51598 44000
rect 51654 43966 51688 44000
rect 51744 43966 51778 44000
rect 51834 43966 51868 44000
rect 51924 43966 51958 44000
rect 22721 41147 22755 41181
rect 22721 41079 22755 41113
rect 22721 41011 22755 41045
rect 22721 40943 22755 40977
rect 22721 40875 22755 40909
rect 22721 40807 22755 40841
rect 22721 40739 22755 40773
rect 22721 40671 22755 40705
rect 22721 40603 22755 40637
rect 22721 40535 22755 40569
rect 22721 40467 22755 40501
rect 22721 40399 22755 40433
rect 22721 40331 22755 40365
rect 22721 40263 22755 40297
rect 22721 40195 22755 40229
rect 22721 40127 22755 40161
rect 22721 40059 22755 40093
rect 22721 39991 22755 40025
rect 22721 39923 22755 39957
rect 23179 41147 23213 41181
rect 23179 41079 23213 41113
rect 23179 41011 23213 41045
rect 23179 40943 23213 40977
rect 23179 40875 23213 40909
rect 23179 40807 23213 40841
rect 23179 40739 23213 40773
rect 23179 40671 23213 40705
rect 23179 40603 23213 40637
rect 23179 40535 23213 40569
rect 23179 40467 23213 40501
rect 23179 40399 23213 40433
rect 23179 40331 23213 40365
rect 23179 40263 23213 40297
rect 23179 40195 23213 40229
rect 23179 40127 23213 40161
rect 23179 40059 23213 40093
rect 23179 39991 23213 40025
rect 23179 39923 23213 39957
rect 23637 41147 23671 41181
rect 23637 41079 23671 41113
rect 23637 41011 23671 41045
rect 23637 40943 23671 40977
rect 23637 40875 23671 40909
rect 23637 40807 23671 40841
rect 23637 40739 23671 40773
rect 23637 40671 23671 40705
rect 23637 40603 23671 40637
rect 23637 40535 23671 40569
rect 23637 40467 23671 40501
rect 23637 40399 23671 40433
rect 23637 40331 23671 40365
rect 23637 40263 23671 40297
rect 23637 40195 23671 40229
rect 23637 40127 23671 40161
rect 23637 40059 23671 40093
rect 23637 39991 23671 40025
rect 23637 39923 23671 39957
rect 24095 41147 24129 41181
rect 24095 41079 24129 41113
rect 24095 41011 24129 41045
rect 24095 40943 24129 40977
rect 24095 40875 24129 40909
rect 24095 40807 24129 40841
rect 24095 40739 24129 40773
rect 24095 40671 24129 40705
rect 24095 40603 24129 40637
rect 24095 40535 24129 40569
rect 24095 40467 24129 40501
rect 24095 40399 24129 40433
rect 24095 40331 24129 40365
rect 24095 40263 24129 40297
rect 24095 40195 24129 40229
rect 24095 40127 24129 40161
rect 24095 40059 24129 40093
rect 24095 39991 24129 40025
rect 24095 39923 24129 39957
rect 24553 41147 24587 41181
rect 24553 41079 24587 41113
rect 24553 41011 24587 41045
rect 24553 40943 24587 40977
rect 24553 40875 24587 40909
rect 24553 40807 24587 40841
rect 24553 40739 24587 40773
rect 24553 40671 24587 40705
rect 24553 40603 24587 40637
rect 24553 40535 24587 40569
rect 24553 40467 24587 40501
rect 24553 40399 24587 40433
rect 24553 40331 24587 40365
rect 24553 40263 24587 40297
rect 24553 40195 24587 40229
rect 24553 40127 24587 40161
rect 24553 40059 24587 40093
rect 24553 39991 24587 40025
rect 24553 39923 24587 39957
rect 25011 41147 25045 41181
rect 25011 41079 25045 41113
rect 25011 41011 25045 41045
rect 25011 40943 25045 40977
rect 25011 40875 25045 40909
rect 25011 40807 25045 40841
rect 25011 40739 25045 40773
rect 25011 40671 25045 40705
rect 25011 40603 25045 40637
rect 25011 40535 25045 40569
rect 25011 40467 25045 40501
rect 25011 40399 25045 40433
rect 25011 40331 25045 40365
rect 25011 40263 25045 40297
rect 25011 40195 25045 40229
rect 25011 40127 25045 40161
rect 25011 40059 25045 40093
rect 25011 39991 25045 40025
rect 25011 39923 25045 39957
rect 25469 41147 25503 41181
rect 25469 41079 25503 41113
rect 25469 41011 25503 41045
rect 25469 40943 25503 40977
rect 25469 40875 25503 40909
rect 25469 40807 25503 40841
rect 25469 40739 25503 40773
rect 25469 40671 25503 40705
rect 25469 40603 25503 40637
rect 25469 40535 25503 40569
rect 25469 40467 25503 40501
rect 25469 40399 25503 40433
rect 25469 40331 25503 40365
rect 25469 40263 25503 40297
rect 25469 40195 25503 40229
rect 25469 40127 25503 40161
rect 25469 40059 25503 40093
rect 25469 39991 25503 40025
rect 25469 39923 25503 39957
rect 25927 41147 25961 41181
rect 25927 41079 25961 41113
rect 25927 41011 25961 41045
rect 25927 40943 25961 40977
rect 25927 40875 25961 40909
rect 25927 40807 25961 40841
rect 25927 40739 25961 40773
rect 25927 40671 25961 40705
rect 25927 40603 25961 40637
rect 25927 40535 25961 40569
rect 25927 40467 25961 40501
rect 25927 40399 25961 40433
rect 25927 40331 25961 40365
rect 25927 40263 25961 40297
rect 25927 40195 25961 40229
rect 25927 40127 25961 40161
rect 25927 40059 25961 40093
rect 25927 39991 25961 40025
rect 25927 39923 25961 39957
rect 26385 41147 26419 41181
rect 26385 41079 26419 41113
rect 26385 41011 26419 41045
rect 26385 40943 26419 40977
rect 26385 40875 26419 40909
rect 26385 40807 26419 40841
rect 26385 40739 26419 40773
rect 26385 40671 26419 40705
rect 26385 40603 26419 40637
rect 26385 40535 26419 40569
rect 26385 40467 26419 40501
rect 26385 40399 26419 40433
rect 26385 40331 26419 40365
rect 26385 40263 26419 40297
rect 26385 40195 26419 40229
rect 26385 40127 26419 40161
rect 26385 40059 26419 40093
rect 26385 39991 26419 40025
rect 26385 39923 26419 39957
rect 26843 41147 26877 41181
rect 26843 41079 26877 41113
rect 26843 41011 26877 41045
rect 26843 40943 26877 40977
rect 26843 40875 26877 40909
rect 26843 40807 26877 40841
rect 26843 40739 26877 40773
rect 26843 40671 26877 40705
rect 26843 40603 26877 40637
rect 26843 40535 26877 40569
rect 26843 40467 26877 40501
rect 26843 40399 26877 40433
rect 26843 40331 26877 40365
rect 26843 40263 26877 40297
rect 26843 40195 26877 40229
rect 26843 40127 26877 40161
rect 26843 40059 26877 40093
rect 26843 39991 26877 40025
rect 26843 39923 26877 39957
rect 27301 41147 27335 41181
rect 27301 41079 27335 41113
rect 27301 41011 27335 41045
rect 27301 40943 27335 40977
rect 27301 40875 27335 40909
rect 27301 40807 27335 40841
rect 27301 40739 27335 40773
rect 27301 40671 27335 40705
rect 27301 40603 27335 40637
rect 27301 40535 27335 40569
rect 27301 40467 27335 40501
rect 27301 40399 27335 40433
rect 27301 40331 27335 40365
rect 27301 40263 27335 40297
rect 27301 40195 27335 40229
rect 27301 40127 27335 40161
rect 27301 40059 27335 40093
rect 27301 39991 27335 40025
rect 27301 39923 27335 39957
rect 27759 41147 27793 41181
rect 27759 41079 27793 41113
rect 27759 41011 27793 41045
rect 27759 40943 27793 40977
rect 27759 40875 27793 40909
rect 27759 40807 27793 40841
rect 27759 40739 27793 40773
rect 27759 40671 27793 40705
rect 27759 40603 27793 40637
rect 27759 40535 27793 40569
rect 27759 40467 27793 40501
rect 27759 40399 27793 40433
rect 27759 40331 27793 40365
rect 27759 40263 27793 40297
rect 27759 40195 27793 40229
rect 27759 40127 27793 40161
rect 27759 40059 27793 40093
rect 27759 39991 27793 40025
rect 27759 39923 27793 39957
rect 28217 41147 28251 41181
rect 28217 41079 28251 41113
rect 28217 41011 28251 41045
rect 28217 40943 28251 40977
rect 28217 40875 28251 40909
rect 28217 40807 28251 40841
rect 28217 40739 28251 40773
rect 28217 40671 28251 40705
rect 28217 40603 28251 40637
rect 28217 40535 28251 40569
rect 28217 40467 28251 40501
rect 28217 40399 28251 40433
rect 28217 40331 28251 40365
rect 28217 40263 28251 40297
rect 28217 40195 28251 40229
rect 28217 40127 28251 40161
rect 28217 40059 28251 40093
rect 28217 39991 28251 40025
rect 28217 39923 28251 39957
rect 29385 41147 29419 41181
rect 29385 41079 29419 41113
rect 29385 41011 29419 41045
rect 29385 40943 29419 40977
rect 29385 40875 29419 40909
rect 29385 40807 29419 40841
rect 29385 40739 29419 40773
rect 29385 40671 29419 40705
rect 29385 40603 29419 40637
rect 29385 40535 29419 40569
rect 29385 40467 29419 40501
rect 29385 40399 29419 40433
rect 29385 40331 29419 40365
rect 29385 40263 29419 40297
rect 29385 40195 29419 40229
rect 29385 40127 29419 40161
rect 29385 40059 29419 40093
rect 29385 39991 29419 40025
rect 29385 39923 29419 39957
rect 29843 41147 29877 41181
rect 29843 41079 29877 41113
rect 29843 41011 29877 41045
rect 29843 40943 29877 40977
rect 29843 40875 29877 40909
rect 29843 40807 29877 40841
rect 29843 40739 29877 40773
rect 29843 40671 29877 40705
rect 29843 40603 29877 40637
rect 29843 40535 29877 40569
rect 29843 40467 29877 40501
rect 29843 40399 29877 40433
rect 29843 40331 29877 40365
rect 29843 40263 29877 40297
rect 29843 40195 29877 40229
rect 29843 40127 29877 40161
rect 29843 40059 29877 40093
rect 29843 39991 29877 40025
rect 29843 39923 29877 39957
rect 30301 41147 30335 41181
rect 30301 41079 30335 41113
rect 30301 41011 30335 41045
rect 30301 40943 30335 40977
rect 30301 40875 30335 40909
rect 30301 40807 30335 40841
rect 30301 40739 30335 40773
rect 30301 40671 30335 40705
rect 30301 40603 30335 40637
rect 30301 40535 30335 40569
rect 30301 40467 30335 40501
rect 30301 40399 30335 40433
rect 30301 40331 30335 40365
rect 30301 40263 30335 40297
rect 30301 40195 30335 40229
rect 30301 40127 30335 40161
rect 30301 40059 30335 40093
rect 30301 39991 30335 40025
rect 30301 39923 30335 39957
rect 30759 41147 30793 41181
rect 30759 41079 30793 41113
rect 30759 41011 30793 41045
rect 30759 40943 30793 40977
rect 30759 40875 30793 40909
rect 30759 40807 30793 40841
rect 30759 40739 30793 40773
rect 30759 40671 30793 40705
rect 30759 40603 30793 40637
rect 30759 40535 30793 40569
rect 30759 40467 30793 40501
rect 30759 40399 30793 40433
rect 30759 40331 30793 40365
rect 30759 40263 30793 40297
rect 30759 40195 30793 40229
rect 30759 40127 30793 40161
rect 30759 40059 30793 40093
rect 30759 39991 30793 40025
rect 30759 39923 30793 39957
rect 31217 41147 31251 41181
rect 31217 41079 31251 41113
rect 31217 41011 31251 41045
rect 31217 40943 31251 40977
rect 31217 40875 31251 40909
rect 31217 40807 31251 40841
rect 31217 40739 31251 40773
rect 31217 40671 31251 40705
rect 31217 40603 31251 40637
rect 31217 40535 31251 40569
rect 31217 40467 31251 40501
rect 31217 40399 31251 40433
rect 31217 40331 31251 40365
rect 31217 40263 31251 40297
rect 31217 40195 31251 40229
rect 31217 40127 31251 40161
rect 31217 40059 31251 40093
rect 31217 39991 31251 40025
rect 31217 39923 31251 39957
rect 31675 41147 31709 41181
rect 31675 41079 31709 41113
rect 31675 41011 31709 41045
rect 31675 40943 31709 40977
rect 31675 40875 31709 40909
rect 31675 40807 31709 40841
rect 31675 40739 31709 40773
rect 31675 40671 31709 40705
rect 31675 40603 31709 40637
rect 31675 40535 31709 40569
rect 31675 40467 31709 40501
rect 31675 40399 31709 40433
rect 31675 40331 31709 40365
rect 31675 40263 31709 40297
rect 31675 40195 31709 40229
rect 31675 40127 31709 40161
rect 31675 40059 31709 40093
rect 31675 39991 31709 40025
rect 31675 39923 31709 39957
rect 32133 41147 32167 41181
rect 32133 41079 32167 41113
rect 32133 41011 32167 41045
rect 32133 40943 32167 40977
rect 32133 40875 32167 40909
rect 32133 40807 32167 40841
rect 32133 40739 32167 40773
rect 32133 40671 32167 40705
rect 32133 40603 32167 40637
rect 32133 40535 32167 40569
rect 32133 40467 32167 40501
rect 32133 40399 32167 40433
rect 32133 40331 32167 40365
rect 32133 40263 32167 40297
rect 32133 40195 32167 40229
rect 32133 40127 32167 40161
rect 32133 40059 32167 40093
rect 32133 39991 32167 40025
rect 32133 39923 32167 39957
rect 32591 41147 32625 41181
rect 32591 41079 32625 41113
rect 32591 41011 32625 41045
rect 32591 40943 32625 40977
rect 32591 40875 32625 40909
rect 32591 40807 32625 40841
rect 32591 40739 32625 40773
rect 32591 40671 32625 40705
rect 32591 40603 32625 40637
rect 32591 40535 32625 40569
rect 32591 40467 32625 40501
rect 32591 40399 32625 40433
rect 32591 40331 32625 40365
rect 32591 40263 32625 40297
rect 32591 40195 32625 40229
rect 32591 40127 32625 40161
rect 32591 40059 32625 40093
rect 32591 39991 32625 40025
rect 32591 39923 32625 39957
rect 33049 41147 33083 41181
rect 33049 41079 33083 41113
rect 33049 41011 33083 41045
rect 33049 40943 33083 40977
rect 33049 40875 33083 40909
rect 33049 40807 33083 40841
rect 33049 40739 33083 40773
rect 33049 40671 33083 40705
rect 33049 40603 33083 40637
rect 33049 40535 33083 40569
rect 33049 40467 33083 40501
rect 33049 40399 33083 40433
rect 33049 40331 33083 40365
rect 33049 40263 33083 40297
rect 33049 40195 33083 40229
rect 33049 40127 33083 40161
rect 33049 40059 33083 40093
rect 33049 39991 33083 40025
rect 33049 39923 33083 39957
rect 33507 41147 33541 41181
rect 33507 41079 33541 41113
rect 33507 41011 33541 41045
rect 33507 40943 33541 40977
rect 33507 40875 33541 40909
rect 33507 40807 33541 40841
rect 33507 40739 33541 40773
rect 33507 40671 33541 40705
rect 33507 40603 33541 40637
rect 33507 40535 33541 40569
rect 33507 40467 33541 40501
rect 33507 40399 33541 40433
rect 33507 40331 33541 40365
rect 33507 40263 33541 40297
rect 33507 40195 33541 40229
rect 33507 40127 33541 40161
rect 33507 40059 33541 40093
rect 33507 39991 33541 40025
rect 33507 39923 33541 39957
rect 33965 41147 33999 41181
rect 33965 41079 33999 41113
rect 33965 41011 33999 41045
rect 33965 40943 33999 40977
rect 33965 40875 33999 40909
rect 33965 40807 33999 40841
rect 33965 40739 33999 40773
rect 33965 40671 33999 40705
rect 33965 40603 33999 40637
rect 33965 40535 33999 40569
rect 33965 40467 33999 40501
rect 33965 40399 33999 40433
rect 33965 40331 33999 40365
rect 33965 40263 33999 40297
rect 33965 40195 33999 40229
rect 33965 40127 33999 40161
rect 33965 40059 33999 40093
rect 33965 39991 33999 40025
rect 33965 39923 33999 39957
rect 34423 41147 34457 41181
rect 34423 41079 34457 41113
rect 34423 41011 34457 41045
rect 34423 40943 34457 40977
rect 34423 40875 34457 40909
rect 34423 40807 34457 40841
rect 34423 40739 34457 40773
rect 34423 40671 34457 40705
rect 34423 40603 34457 40637
rect 34423 40535 34457 40569
rect 34423 40467 34457 40501
rect 34423 40399 34457 40433
rect 34423 40331 34457 40365
rect 34423 40263 34457 40297
rect 34423 40195 34457 40229
rect 34423 40127 34457 40161
rect 34423 40059 34457 40093
rect 34423 39991 34457 40025
rect 34423 39923 34457 39957
rect 34881 41147 34915 41181
rect 34881 41079 34915 41113
rect 34881 41011 34915 41045
rect 34881 40943 34915 40977
rect 34881 40875 34915 40909
rect 34881 40807 34915 40841
rect 34881 40739 34915 40773
rect 34881 40671 34915 40705
rect 34881 40603 34915 40637
rect 34881 40535 34915 40569
rect 34881 40467 34915 40501
rect 34881 40399 34915 40433
rect 34881 40331 34915 40365
rect 34881 40263 34915 40297
rect 34881 40195 34915 40229
rect 34881 40127 34915 40161
rect 34881 40059 34915 40093
rect 34881 39991 34915 40025
rect 34881 39923 34915 39957
rect 42168 40746 42202 40780
rect 42258 40746 42292 40780
rect 42348 40746 42382 40780
rect 42438 40746 42472 40780
rect 42528 40746 42562 40780
rect 42618 40746 42652 40780
rect 42708 40746 42742 40780
rect 42168 40656 42202 40690
rect 42258 40656 42292 40690
rect 42348 40656 42382 40690
rect 42438 40656 42472 40690
rect 42528 40656 42562 40690
rect 42618 40656 42652 40690
rect 42708 40656 42742 40690
rect 42168 40566 42202 40600
rect 42258 40566 42292 40600
rect 42348 40566 42382 40600
rect 42438 40566 42472 40600
rect 42528 40566 42562 40600
rect 42618 40566 42652 40600
rect 42708 40566 42742 40600
rect 42168 40476 42202 40510
rect 42258 40476 42292 40510
rect 42348 40476 42382 40510
rect 42438 40476 42472 40510
rect 42528 40476 42562 40510
rect 42618 40476 42652 40510
rect 42708 40476 42742 40510
rect 42168 40386 42202 40420
rect 42258 40386 42292 40420
rect 42348 40386 42382 40420
rect 42438 40386 42472 40420
rect 42528 40386 42562 40420
rect 42618 40386 42652 40420
rect 42708 40386 42742 40420
rect 42168 40296 42202 40330
rect 42258 40296 42292 40330
rect 42348 40296 42382 40330
rect 42438 40296 42472 40330
rect 42528 40296 42562 40330
rect 42618 40296 42652 40330
rect 42708 40296 42742 40330
rect 42168 40206 42202 40240
rect 42258 40206 42292 40240
rect 42348 40206 42382 40240
rect 42438 40206 42472 40240
rect 42528 40206 42562 40240
rect 42618 40206 42652 40240
rect 42708 40206 42742 40240
rect 43508 40746 43542 40780
rect 43598 40746 43632 40780
rect 43688 40746 43722 40780
rect 43778 40746 43812 40780
rect 43868 40746 43902 40780
rect 43958 40746 43992 40780
rect 44048 40746 44082 40780
rect 43508 40656 43542 40690
rect 43598 40656 43632 40690
rect 43688 40656 43722 40690
rect 43778 40656 43812 40690
rect 43868 40656 43902 40690
rect 43958 40656 43992 40690
rect 44048 40656 44082 40690
rect 43508 40566 43542 40600
rect 43598 40566 43632 40600
rect 43688 40566 43722 40600
rect 43778 40566 43812 40600
rect 43868 40566 43902 40600
rect 43958 40566 43992 40600
rect 44048 40566 44082 40600
rect 43508 40476 43542 40510
rect 43598 40476 43632 40510
rect 43688 40476 43722 40510
rect 43778 40476 43812 40510
rect 43868 40476 43902 40510
rect 43958 40476 43992 40510
rect 44048 40476 44082 40510
rect 43508 40386 43542 40420
rect 43598 40386 43632 40420
rect 43688 40386 43722 40420
rect 43778 40386 43812 40420
rect 43868 40386 43902 40420
rect 43958 40386 43992 40420
rect 44048 40386 44082 40420
rect 43508 40296 43542 40330
rect 43598 40296 43632 40330
rect 43688 40296 43722 40330
rect 43778 40296 43812 40330
rect 43868 40296 43902 40330
rect 43958 40296 43992 40330
rect 44048 40296 44082 40330
rect 43508 40206 43542 40240
rect 43598 40206 43632 40240
rect 43688 40206 43722 40240
rect 43778 40206 43812 40240
rect 43868 40206 43902 40240
rect 43958 40206 43992 40240
rect 44048 40206 44082 40240
rect 44848 40746 44882 40780
rect 44938 40746 44972 40780
rect 45028 40746 45062 40780
rect 45118 40746 45152 40780
rect 45208 40746 45242 40780
rect 45298 40746 45332 40780
rect 45388 40746 45422 40780
rect 44848 40656 44882 40690
rect 44938 40656 44972 40690
rect 45028 40656 45062 40690
rect 45118 40656 45152 40690
rect 45208 40656 45242 40690
rect 45298 40656 45332 40690
rect 45388 40656 45422 40690
rect 44848 40566 44882 40600
rect 44938 40566 44972 40600
rect 45028 40566 45062 40600
rect 45118 40566 45152 40600
rect 45208 40566 45242 40600
rect 45298 40566 45332 40600
rect 45388 40566 45422 40600
rect 44848 40476 44882 40510
rect 44938 40476 44972 40510
rect 45028 40476 45062 40510
rect 45118 40476 45152 40510
rect 45208 40476 45242 40510
rect 45298 40476 45332 40510
rect 45388 40476 45422 40510
rect 44848 40386 44882 40420
rect 44938 40386 44972 40420
rect 45028 40386 45062 40420
rect 45118 40386 45152 40420
rect 45208 40386 45242 40420
rect 45298 40386 45332 40420
rect 45388 40386 45422 40420
rect 44848 40296 44882 40330
rect 44938 40296 44972 40330
rect 45028 40296 45062 40330
rect 45118 40296 45152 40330
rect 45208 40296 45242 40330
rect 45298 40296 45332 40330
rect 45388 40296 45422 40330
rect 44848 40206 44882 40240
rect 44938 40206 44972 40240
rect 45028 40206 45062 40240
rect 45118 40206 45152 40240
rect 45208 40206 45242 40240
rect 45298 40206 45332 40240
rect 45388 40206 45422 40240
rect 46188 40746 46222 40780
rect 46278 40746 46312 40780
rect 46368 40746 46402 40780
rect 46458 40746 46492 40780
rect 46548 40746 46582 40780
rect 46638 40746 46672 40780
rect 46728 40746 46762 40780
rect 46188 40656 46222 40690
rect 46278 40656 46312 40690
rect 46368 40656 46402 40690
rect 46458 40656 46492 40690
rect 46548 40656 46582 40690
rect 46638 40656 46672 40690
rect 46728 40656 46762 40690
rect 46188 40566 46222 40600
rect 46278 40566 46312 40600
rect 46368 40566 46402 40600
rect 46458 40566 46492 40600
rect 46548 40566 46582 40600
rect 46638 40566 46672 40600
rect 46728 40566 46762 40600
rect 46188 40476 46222 40510
rect 46278 40476 46312 40510
rect 46368 40476 46402 40510
rect 46458 40476 46492 40510
rect 46548 40476 46582 40510
rect 46638 40476 46672 40510
rect 46728 40476 46762 40510
rect 46188 40386 46222 40420
rect 46278 40386 46312 40420
rect 46368 40386 46402 40420
rect 46458 40386 46492 40420
rect 46548 40386 46582 40420
rect 46638 40386 46672 40420
rect 46728 40386 46762 40420
rect 46188 40296 46222 40330
rect 46278 40296 46312 40330
rect 46368 40296 46402 40330
rect 46458 40296 46492 40330
rect 46548 40296 46582 40330
rect 46638 40296 46672 40330
rect 46728 40296 46762 40330
rect 46188 40206 46222 40240
rect 46278 40206 46312 40240
rect 46368 40206 46402 40240
rect 46458 40206 46492 40240
rect 46548 40206 46582 40240
rect 46638 40206 46672 40240
rect 46728 40206 46762 40240
rect 47528 40746 47562 40780
rect 47618 40746 47652 40780
rect 47708 40746 47742 40780
rect 47798 40746 47832 40780
rect 47888 40746 47922 40780
rect 47978 40746 48012 40780
rect 48068 40746 48102 40780
rect 47528 40656 47562 40690
rect 47618 40656 47652 40690
rect 47708 40656 47742 40690
rect 47798 40656 47832 40690
rect 47888 40656 47922 40690
rect 47978 40656 48012 40690
rect 48068 40656 48102 40690
rect 47528 40566 47562 40600
rect 47618 40566 47652 40600
rect 47708 40566 47742 40600
rect 47798 40566 47832 40600
rect 47888 40566 47922 40600
rect 47978 40566 48012 40600
rect 48068 40566 48102 40600
rect 47528 40476 47562 40510
rect 47618 40476 47652 40510
rect 47708 40476 47742 40510
rect 47798 40476 47832 40510
rect 47888 40476 47922 40510
rect 47978 40476 48012 40510
rect 48068 40476 48102 40510
rect 47528 40386 47562 40420
rect 47618 40386 47652 40420
rect 47708 40386 47742 40420
rect 47798 40386 47832 40420
rect 47888 40386 47922 40420
rect 47978 40386 48012 40420
rect 48068 40386 48102 40420
rect 47528 40296 47562 40330
rect 47618 40296 47652 40330
rect 47708 40296 47742 40330
rect 47798 40296 47832 40330
rect 47888 40296 47922 40330
rect 47978 40296 48012 40330
rect 48068 40296 48102 40330
rect 47528 40206 47562 40240
rect 47618 40206 47652 40240
rect 47708 40206 47742 40240
rect 47798 40206 47832 40240
rect 47888 40206 47922 40240
rect 47978 40206 48012 40240
rect 48068 40206 48102 40240
rect 48868 40746 48902 40780
rect 48958 40746 48992 40780
rect 49048 40746 49082 40780
rect 49138 40746 49172 40780
rect 49228 40746 49262 40780
rect 49318 40746 49352 40780
rect 49408 40746 49442 40780
rect 48868 40656 48902 40690
rect 48958 40656 48992 40690
rect 49048 40656 49082 40690
rect 49138 40656 49172 40690
rect 49228 40656 49262 40690
rect 49318 40656 49352 40690
rect 49408 40656 49442 40690
rect 48868 40566 48902 40600
rect 48958 40566 48992 40600
rect 49048 40566 49082 40600
rect 49138 40566 49172 40600
rect 49228 40566 49262 40600
rect 49318 40566 49352 40600
rect 49408 40566 49442 40600
rect 48868 40476 48902 40510
rect 48958 40476 48992 40510
rect 49048 40476 49082 40510
rect 49138 40476 49172 40510
rect 49228 40476 49262 40510
rect 49318 40476 49352 40510
rect 49408 40476 49442 40510
rect 48868 40386 48902 40420
rect 48958 40386 48992 40420
rect 49048 40386 49082 40420
rect 49138 40386 49172 40420
rect 49228 40386 49262 40420
rect 49318 40386 49352 40420
rect 49408 40386 49442 40420
rect 48868 40296 48902 40330
rect 48958 40296 48992 40330
rect 49048 40296 49082 40330
rect 49138 40296 49172 40330
rect 49228 40296 49262 40330
rect 49318 40296 49352 40330
rect 49408 40296 49442 40330
rect 48868 40206 48902 40240
rect 48958 40206 48992 40240
rect 49048 40206 49082 40240
rect 49138 40206 49172 40240
rect 49228 40206 49262 40240
rect 49318 40206 49352 40240
rect 49408 40206 49442 40240
rect 50208 40746 50242 40780
rect 50298 40746 50332 40780
rect 50388 40746 50422 40780
rect 50478 40746 50512 40780
rect 50568 40746 50602 40780
rect 50658 40746 50692 40780
rect 50748 40746 50782 40780
rect 50208 40656 50242 40690
rect 50298 40656 50332 40690
rect 50388 40656 50422 40690
rect 50478 40656 50512 40690
rect 50568 40656 50602 40690
rect 50658 40656 50692 40690
rect 50748 40656 50782 40690
rect 50208 40566 50242 40600
rect 50298 40566 50332 40600
rect 50388 40566 50422 40600
rect 50478 40566 50512 40600
rect 50568 40566 50602 40600
rect 50658 40566 50692 40600
rect 50748 40566 50782 40600
rect 50208 40476 50242 40510
rect 50298 40476 50332 40510
rect 50388 40476 50422 40510
rect 50478 40476 50512 40510
rect 50568 40476 50602 40510
rect 50658 40476 50692 40510
rect 50748 40476 50782 40510
rect 50208 40386 50242 40420
rect 50298 40386 50332 40420
rect 50388 40386 50422 40420
rect 50478 40386 50512 40420
rect 50568 40386 50602 40420
rect 50658 40386 50692 40420
rect 50748 40386 50782 40420
rect 50208 40296 50242 40330
rect 50298 40296 50332 40330
rect 50388 40296 50422 40330
rect 50478 40296 50512 40330
rect 50568 40296 50602 40330
rect 50658 40296 50692 40330
rect 50748 40296 50782 40330
rect 50208 40206 50242 40240
rect 50298 40206 50332 40240
rect 50388 40206 50422 40240
rect 50478 40206 50512 40240
rect 50568 40206 50602 40240
rect 50658 40206 50692 40240
rect 50748 40206 50782 40240
rect 51548 40746 51582 40780
rect 51638 40746 51672 40780
rect 51728 40746 51762 40780
rect 51818 40746 51852 40780
rect 51908 40746 51942 40780
rect 51998 40746 52032 40780
rect 52088 40746 52122 40780
rect 51548 40656 51582 40690
rect 51638 40656 51672 40690
rect 51728 40656 51762 40690
rect 51818 40656 51852 40690
rect 51908 40656 51942 40690
rect 51998 40656 52032 40690
rect 52088 40656 52122 40690
rect 51548 40566 51582 40600
rect 51638 40566 51672 40600
rect 51728 40566 51762 40600
rect 51818 40566 51852 40600
rect 51908 40566 51942 40600
rect 51998 40566 52032 40600
rect 52088 40566 52122 40600
rect 51548 40476 51582 40510
rect 51638 40476 51672 40510
rect 51728 40476 51762 40510
rect 51818 40476 51852 40510
rect 51908 40476 51942 40510
rect 51998 40476 52032 40510
rect 52088 40476 52122 40510
rect 51548 40386 51582 40420
rect 51638 40386 51672 40420
rect 51728 40386 51762 40420
rect 51818 40386 51852 40420
rect 51908 40386 51942 40420
rect 51998 40386 52032 40420
rect 52088 40386 52122 40420
rect 51548 40296 51582 40330
rect 51638 40296 51672 40330
rect 51728 40296 51762 40330
rect 51818 40296 51852 40330
rect 51908 40296 51942 40330
rect 51998 40296 52032 40330
rect 52088 40296 52122 40330
rect 51548 40206 51582 40240
rect 51638 40206 51672 40240
rect 51728 40206 51762 40240
rect 51818 40206 51852 40240
rect 51908 40206 51942 40240
rect 51998 40206 52032 40240
rect 52088 40206 52122 40240
rect 12376 36986 12410 37020
rect 12466 36986 12500 37020
rect 12556 36986 12590 37020
rect 12646 36986 12680 37020
rect 12736 36986 12770 37020
rect 12826 36986 12860 37020
rect 12916 36986 12950 37020
rect 12376 36896 12410 36930
rect 12466 36896 12500 36930
rect 12556 36896 12590 36930
rect 12646 36896 12680 36930
rect 12736 36896 12770 36930
rect 12826 36896 12860 36930
rect 12916 36896 12950 36930
rect 12376 36806 12410 36840
rect 12466 36806 12500 36840
rect 12556 36806 12590 36840
rect 12646 36806 12680 36840
rect 12736 36806 12770 36840
rect 12826 36806 12860 36840
rect 12916 36806 12950 36840
rect 12376 36716 12410 36750
rect 12466 36716 12500 36750
rect 12556 36716 12590 36750
rect 12646 36716 12680 36750
rect 12736 36716 12770 36750
rect 12826 36716 12860 36750
rect 12916 36716 12950 36750
rect 12376 36626 12410 36660
rect 12466 36626 12500 36660
rect 12556 36626 12590 36660
rect 12646 36626 12680 36660
rect 12736 36626 12770 36660
rect 12826 36626 12860 36660
rect 12916 36626 12950 36660
rect 12376 36536 12410 36570
rect 12466 36536 12500 36570
rect 12556 36536 12590 36570
rect 12646 36536 12680 36570
rect 12736 36536 12770 36570
rect 12826 36536 12860 36570
rect 12916 36536 12950 36570
rect 12376 36446 12410 36480
rect 12466 36446 12500 36480
rect 12556 36446 12590 36480
rect 12646 36446 12680 36480
rect 12736 36446 12770 36480
rect 12826 36446 12860 36480
rect 12916 36446 12950 36480
rect 37519 37387 37553 37421
rect 37519 37319 37553 37353
rect 37519 37251 37553 37285
rect 37519 37183 37553 37217
rect 37519 37115 37553 37149
rect 37519 37047 37553 37081
rect 37519 36979 37553 37013
rect 37519 36911 37553 36945
rect 37519 36843 37553 36877
rect 37519 36775 37553 36809
rect 37519 36707 37553 36741
rect 37519 36639 37553 36673
rect 37519 36571 37553 36605
rect 37519 36503 37553 36537
rect 37519 36435 37553 36469
rect 37519 36367 37553 36401
rect 37519 36299 37553 36333
rect 37519 36231 37553 36265
rect 37519 36163 37553 36197
rect 37977 37387 38011 37421
rect 37977 37319 38011 37353
rect 37977 37251 38011 37285
rect 37977 37183 38011 37217
rect 37977 37115 38011 37149
rect 37977 37047 38011 37081
rect 37977 36979 38011 37013
rect 37977 36911 38011 36945
rect 37977 36843 38011 36877
rect 37977 36775 38011 36809
rect 37977 36707 38011 36741
rect 37977 36639 38011 36673
rect 37977 36571 38011 36605
rect 37977 36503 38011 36537
rect 37977 36435 38011 36469
rect 37977 36367 38011 36401
rect 37977 36299 38011 36333
rect 37977 36231 38011 36265
rect 37977 36163 38011 36197
rect 38435 37387 38469 37421
rect 38435 37319 38469 37353
rect 38435 37251 38469 37285
rect 38435 37183 38469 37217
rect 38435 37115 38469 37149
rect 38435 37047 38469 37081
rect 38435 36979 38469 37013
rect 38435 36911 38469 36945
rect 38435 36843 38469 36877
rect 38435 36775 38469 36809
rect 38435 36707 38469 36741
rect 38435 36639 38469 36673
rect 38435 36571 38469 36605
rect 38435 36503 38469 36537
rect 38435 36435 38469 36469
rect 38435 36367 38469 36401
rect 38435 36299 38469 36333
rect 38435 36231 38469 36265
rect 38435 36163 38469 36197
rect 38893 37387 38927 37421
rect 38893 37319 38927 37353
rect 38893 37251 38927 37285
rect 38893 37183 38927 37217
rect 38893 37115 38927 37149
rect 38893 37047 38927 37081
rect 38893 36979 38927 37013
rect 38893 36911 38927 36945
rect 38893 36843 38927 36877
rect 38893 36775 38927 36809
rect 38893 36707 38927 36741
rect 38893 36639 38927 36673
rect 38893 36571 38927 36605
rect 38893 36503 38927 36537
rect 38893 36435 38927 36469
rect 38893 36367 38927 36401
rect 38893 36299 38927 36333
rect 38893 36231 38927 36265
rect 38893 36163 38927 36197
rect 39351 37387 39385 37421
rect 39351 37319 39385 37353
rect 39351 37251 39385 37285
rect 39351 37183 39385 37217
rect 39351 37115 39385 37149
rect 39351 37047 39385 37081
rect 39351 36979 39385 37013
rect 39351 36911 39385 36945
rect 39351 36843 39385 36877
rect 39351 36775 39385 36809
rect 39351 36707 39385 36741
rect 39351 36639 39385 36673
rect 39351 36571 39385 36605
rect 39351 36503 39385 36537
rect 39351 36435 39385 36469
rect 39351 36367 39385 36401
rect 39351 36299 39385 36333
rect 39351 36231 39385 36265
rect 39351 36163 39385 36197
rect 39809 37387 39843 37421
rect 39809 37319 39843 37353
rect 39809 37251 39843 37285
rect 39809 37183 39843 37217
rect 39809 37115 39843 37149
rect 39809 37047 39843 37081
rect 39809 36979 39843 37013
rect 39809 36911 39843 36945
rect 39809 36843 39843 36877
rect 39809 36775 39843 36809
rect 39809 36707 39843 36741
rect 39809 36639 39843 36673
rect 39809 36571 39843 36605
rect 39809 36503 39843 36537
rect 39809 36435 39843 36469
rect 39809 36367 39843 36401
rect 39809 36299 39843 36333
rect 39809 36231 39843 36265
rect 39809 36163 39843 36197
rect 40267 37387 40301 37421
rect 40267 37319 40301 37353
rect 40267 37251 40301 37285
rect 40267 37183 40301 37217
rect 40267 37115 40301 37149
rect 40267 37047 40301 37081
rect 40267 36979 40301 37013
rect 40267 36911 40301 36945
rect 40267 36843 40301 36877
rect 40267 36775 40301 36809
rect 40267 36707 40301 36741
rect 40267 36639 40301 36673
rect 40267 36571 40301 36605
rect 40267 36503 40301 36537
rect 40267 36435 40301 36469
rect 40267 36367 40301 36401
rect 40267 36299 40301 36333
rect 40267 36231 40301 36265
rect 40267 36163 40301 36197
rect 42168 36986 42202 37020
rect 42258 36986 42292 37020
rect 42348 36986 42382 37020
rect 42438 36986 42472 37020
rect 42528 36986 42562 37020
rect 42618 36986 42652 37020
rect 42708 36986 42742 37020
rect 42168 36896 42202 36930
rect 42258 36896 42292 36930
rect 42348 36896 42382 36930
rect 42438 36896 42472 36930
rect 42528 36896 42562 36930
rect 42618 36896 42652 36930
rect 42708 36896 42742 36930
rect 42168 36806 42202 36840
rect 42258 36806 42292 36840
rect 42348 36806 42382 36840
rect 42438 36806 42472 36840
rect 42528 36806 42562 36840
rect 42618 36806 42652 36840
rect 42708 36806 42742 36840
rect 42168 36716 42202 36750
rect 42258 36716 42292 36750
rect 42348 36716 42382 36750
rect 42438 36716 42472 36750
rect 42528 36716 42562 36750
rect 42618 36716 42652 36750
rect 42708 36716 42742 36750
rect 42168 36626 42202 36660
rect 42258 36626 42292 36660
rect 42348 36626 42382 36660
rect 42438 36626 42472 36660
rect 42528 36626 42562 36660
rect 42618 36626 42652 36660
rect 42708 36626 42742 36660
rect 42168 36536 42202 36570
rect 42258 36536 42292 36570
rect 42348 36536 42382 36570
rect 42438 36536 42472 36570
rect 42528 36536 42562 36570
rect 42618 36536 42652 36570
rect 42708 36536 42742 36570
rect 42168 36446 42202 36480
rect 42258 36446 42292 36480
rect 42348 36446 42382 36480
rect 42438 36446 42472 36480
rect 42528 36446 42562 36480
rect 42618 36446 42652 36480
rect 42708 36446 42742 36480
rect 43508 36986 43542 37020
rect 43598 36986 43632 37020
rect 43688 36986 43722 37020
rect 43778 36986 43812 37020
rect 43868 36986 43902 37020
rect 43958 36986 43992 37020
rect 44048 36986 44082 37020
rect 43508 36896 43542 36930
rect 43598 36896 43632 36930
rect 43688 36896 43722 36930
rect 43778 36896 43812 36930
rect 43868 36896 43902 36930
rect 43958 36896 43992 36930
rect 44048 36896 44082 36930
rect 43508 36806 43542 36840
rect 43598 36806 43632 36840
rect 43688 36806 43722 36840
rect 43778 36806 43812 36840
rect 43868 36806 43902 36840
rect 43958 36806 43992 36840
rect 44048 36806 44082 36840
rect 43508 36716 43542 36750
rect 43598 36716 43632 36750
rect 43688 36716 43722 36750
rect 43778 36716 43812 36750
rect 43868 36716 43902 36750
rect 43958 36716 43992 36750
rect 44048 36716 44082 36750
rect 43508 36626 43542 36660
rect 43598 36626 43632 36660
rect 43688 36626 43722 36660
rect 43778 36626 43812 36660
rect 43868 36626 43902 36660
rect 43958 36626 43992 36660
rect 44048 36626 44082 36660
rect 43508 36536 43542 36570
rect 43598 36536 43632 36570
rect 43688 36536 43722 36570
rect 43778 36536 43812 36570
rect 43868 36536 43902 36570
rect 43958 36536 43992 36570
rect 44048 36536 44082 36570
rect 43508 36446 43542 36480
rect 43598 36446 43632 36480
rect 43688 36446 43722 36480
rect 43778 36446 43812 36480
rect 43868 36446 43902 36480
rect 43958 36446 43992 36480
rect 44048 36446 44082 36480
rect 44848 36986 44882 37020
rect 44938 36986 44972 37020
rect 45028 36986 45062 37020
rect 45118 36986 45152 37020
rect 45208 36986 45242 37020
rect 45298 36986 45332 37020
rect 45388 36986 45422 37020
rect 44848 36896 44882 36930
rect 44938 36896 44972 36930
rect 45028 36896 45062 36930
rect 45118 36896 45152 36930
rect 45208 36896 45242 36930
rect 45298 36896 45332 36930
rect 45388 36896 45422 36930
rect 44848 36806 44882 36840
rect 44938 36806 44972 36840
rect 45028 36806 45062 36840
rect 45118 36806 45152 36840
rect 45208 36806 45242 36840
rect 45298 36806 45332 36840
rect 45388 36806 45422 36840
rect 44848 36716 44882 36750
rect 44938 36716 44972 36750
rect 45028 36716 45062 36750
rect 45118 36716 45152 36750
rect 45208 36716 45242 36750
rect 45298 36716 45332 36750
rect 45388 36716 45422 36750
rect 44848 36626 44882 36660
rect 44938 36626 44972 36660
rect 45028 36626 45062 36660
rect 45118 36626 45152 36660
rect 45208 36626 45242 36660
rect 45298 36626 45332 36660
rect 45388 36626 45422 36660
rect 44848 36536 44882 36570
rect 44938 36536 44972 36570
rect 45028 36536 45062 36570
rect 45118 36536 45152 36570
rect 45208 36536 45242 36570
rect 45298 36536 45332 36570
rect 45388 36536 45422 36570
rect 44848 36446 44882 36480
rect 44938 36446 44972 36480
rect 45028 36446 45062 36480
rect 45118 36446 45152 36480
rect 45208 36446 45242 36480
rect 45298 36446 45332 36480
rect 45388 36446 45422 36480
rect 46188 36986 46222 37020
rect 46278 36986 46312 37020
rect 46368 36986 46402 37020
rect 46458 36986 46492 37020
rect 46548 36986 46582 37020
rect 46638 36986 46672 37020
rect 46728 36986 46762 37020
rect 46188 36896 46222 36930
rect 46278 36896 46312 36930
rect 46368 36896 46402 36930
rect 46458 36896 46492 36930
rect 46548 36896 46582 36930
rect 46638 36896 46672 36930
rect 46728 36896 46762 36930
rect 46188 36806 46222 36840
rect 46278 36806 46312 36840
rect 46368 36806 46402 36840
rect 46458 36806 46492 36840
rect 46548 36806 46582 36840
rect 46638 36806 46672 36840
rect 46728 36806 46762 36840
rect 46188 36716 46222 36750
rect 46278 36716 46312 36750
rect 46368 36716 46402 36750
rect 46458 36716 46492 36750
rect 46548 36716 46582 36750
rect 46638 36716 46672 36750
rect 46728 36716 46762 36750
rect 46188 36626 46222 36660
rect 46278 36626 46312 36660
rect 46368 36626 46402 36660
rect 46458 36626 46492 36660
rect 46548 36626 46582 36660
rect 46638 36626 46672 36660
rect 46728 36626 46762 36660
rect 46188 36536 46222 36570
rect 46278 36536 46312 36570
rect 46368 36536 46402 36570
rect 46458 36536 46492 36570
rect 46548 36536 46582 36570
rect 46638 36536 46672 36570
rect 46728 36536 46762 36570
rect 46188 36446 46222 36480
rect 46278 36446 46312 36480
rect 46368 36446 46402 36480
rect 46458 36446 46492 36480
rect 46548 36446 46582 36480
rect 46638 36446 46672 36480
rect 46728 36446 46762 36480
rect 47528 36986 47562 37020
rect 47618 36986 47652 37020
rect 47708 36986 47742 37020
rect 47798 36986 47832 37020
rect 47888 36986 47922 37020
rect 47978 36986 48012 37020
rect 48068 36986 48102 37020
rect 47528 36896 47562 36930
rect 47618 36896 47652 36930
rect 47708 36896 47742 36930
rect 47798 36896 47832 36930
rect 47888 36896 47922 36930
rect 47978 36896 48012 36930
rect 48068 36896 48102 36930
rect 47528 36806 47562 36840
rect 47618 36806 47652 36840
rect 47708 36806 47742 36840
rect 47798 36806 47832 36840
rect 47888 36806 47922 36840
rect 47978 36806 48012 36840
rect 48068 36806 48102 36840
rect 47528 36716 47562 36750
rect 47618 36716 47652 36750
rect 47708 36716 47742 36750
rect 47798 36716 47832 36750
rect 47888 36716 47922 36750
rect 47978 36716 48012 36750
rect 48068 36716 48102 36750
rect 47528 36626 47562 36660
rect 47618 36626 47652 36660
rect 47708 36626 47742 36660
rect 47798 36626 47832 36660
rect 47888 36626 47922 36660
rect 47978 36626 48012 36660
rect 48068 36626 48102 36660
rect 47528 36536 47562 36570
rect 47618 36536 47652 36570
rect 47708 36536 47742 36570
rect 47798 36536 47832 36570
rect 47888 36536 47922 36570
rect 47978 36536 48012 36570
rect 48068 36536 48102 36570
rect 47528 36446 47562 36480
rect 47618 36446 47652 36480
rect 47708 36446 47742 36480
rect 47798 36446 47832 36480
rect 47888 36446 47922 36480
rect 47978 36446 48012 36480
rect 48068 36446 48102 36480
rect 48868 36986 48902 37020
rect 48958 36986 48992 37020
rect 49048 36986 49082 37020
rect 49138 36986 49172 37020
rect 49228 36986 49262 37020
rect 49318 36986 49352 37020
rect 49408 36986 49442 37020
rect 48868 36896 48902 36930
rect 48958 36896 48992 36930
rect 49048 36896 49082 36930
rect 49138 36896 49172 36930
rect 49228 36896 49262 36930
rect 49318 36896 49352 36930
rect 49408 36896 49442 36930
rect 48868 36806 48902 36840
rect 48958 36806 48992 36840
rect 49048 36806 49082 36840
rect 49138 36806 49172 36840
rect 49228 36806 49262 36840
rect 49318 36806 49352 36840
rect 49408 36806 49442 36840
rect 48868 36716 48902 36750
rect 48958 36716 48992 36750
rect 49048 36716 49082 36750
rect 49138 36716 49172 36750
rect 49228 36716 49262 36750
rect 49318 36716 49352 36750
rect 49408 36716 49442 36750
rect 48868 36626 48902 36660
rect 48958 36626 48992 36660
rect 49048 36626 49082 36660
rect 49138 36626 49172 36660
rect 49228 36626 49262 36660
rect 49318 36626 49352 36660
rect 49408 36626 49442 36660
rect 48868 36536 48902 36570
rect 48958 36536 48992 36570
rect 49048 36536 49082 36570
rect 49138 36536 49172 36570
rect 49228 36536 49262 36570
rect 49318 36536 49352 36570
rect 49408 36536 49442 36570
rect 48868 36446 48902 36480
rect 48958 36446 48992 36480
rect 49048 36446 49082 36480
rect 49138 36446 49172 36480
rect 49228 36446 49262 36480
rect 49318 36446 49352 36480
rect 49408 36446 49442 36480
rect 50208 36986 50242 37020
rect 50298 36986 50332 37020
rect 50388 36986 50422 37020
rect 50478 36986 50512 37020
rect 50568 36986 50602 37020
rect 50658 36986 50692 37020
rect 50748 36986 50782 37020
rect 50208 36896 50242 36930
rect 50298 36896 50332 36930
rect 50388 36896 50422 36930
rect 50478 36896 50512 36930
rect 50568 36896 50602 36930
rect 50658 36896 50692 36930
rect 50748 36896 50782 36930
rect 50208 36806 50242 36840
rect 50298 36806 50332 36840
rect 50388 36806 50422 36840
rect 50478 36806 50512 36840
rect 50568 36806 50602 36840
rect 50658 36806 50692 36840
rect 50748 36806 50782 36840
rect 50208 36716 50242 36750
rect 50298 36716 50332 36750
rect 50388 36716 50422 36750
rect 50478 36716 50512 36750
rect 50568 36716 50602 36750
rect 50658 36716 50692 36750
rect 50748 36716 50782 36750
rect 50208 36626 50242 36660
rect 50298 36626 50332 36660
rect 50388 36626 50422 36660
rect 50478 36626 50512 36660
rect 50568 36626 50602 36660
rect 50658 36626 50692 36660
rect 50748 36626 50782 36660
rect 50208 36536 50242 36570
rect 50298 36536 50332 36570
rect 50388 36536 50422 36570
rect 50478 36536 50512 36570
rect 50568 36536 50602 36570
rect 50658 36536 50692 36570
rect 50748 36536 50782 36570
rect 50208 36446 50242 36480
rect 50298 36446 50332 36480
rect 50388 36446 50422 36480
rect 50478 36446 50512 36480
rect 50568 36446 50602 36480
rect 50658 36446 50692 36480
rect 50748 36446 50782 36480
rect 51548 36986 51582 37020
rect 51638 36986 51672 37020
rect 51728 36986 51762 37020
rect 51818 36986 51852 37020
rect 51908 36986 51942 37020
rect 51998 36986 52032 37020
rect 52088 36986 52122 37020
rect 51548 36896 51582 36930
rect 51638 36896 51672 36930
rect 51728 36896 51762 36930
rect 51818 36896 51852 36930
rect 51908 36896 51942 36930
rect 51998 36896 52032 36930
rect 52088 36896 52122 36930
rect 51548 36806 51582 36840
rect 51638 36806 51672 36840
rect 51728 36806 51762 36840
rect 51818 36806 51852 36840
rect 51908 36806 51942 36840
rect 51998 36806 52032 36840
rect 52088 36806 52122 36840
rect 51548 36716 51582 36750
rect 51638 36716 51672 36750
rect 51728 36716 51762 36750
rect 51818 36716 51852 36750
rect 51908 36716 51942 36750
rect 51998 36716 52032 36750
rect 52088 36716 52122 36750
rect 51548 36626 51582 36660
rect 51638 36626 51672 36660
rect 51728 36626 51762 36660
rect 51818 36626 51852 36660
rect 51908 36626 51942 36660
rect 51998 36626 52032 36660
rect 52088 36626 52122 36660
rect 51548 36536 51582 36570
rect 51638 36536 51672 36570
rect 51728 36536 51762 36570
rect 51818 36536 51852 36570
rect 51908 36536 51942 36570
rect 51998 36536 52032 36570
rect 52088 36536 52122 36570
rect 51548 36446 51582 36480
rect 51638 36446 51672 36480
rect 51728 36446 51762 36480
rect 51818 36446 51852 36480
rect 51908 36446 51942 36480
rect 51998 36446 52032 36480
rect 52088 36446 52122 36480
rect 42168 33226 42202 33260
rect 42258 33226 42292 33260
rect 42348 33226 42382 33260
rect 42438 33226 42472 33260
rect 42528 33226 42562 33260
rect 42618 33226 42652 33260
rect 42708 33226 42742 33260
rect 42168 33136 42202 33170
rect 42258 33136 42292 33170
rect 42348 33136 42382 33170
rect 42438 33136 42472 33170
rect 42528 33136 42562 33170
rect 42618 33136 42652 33170
rect 42708 33136 42742 33170
rect 42168 33046 42202 33080
rect 42258 33046 42292 33080
rect 42348 33046 42382 33080
rect 42438 33046 42472 33080
rect 42528 33046 42562 33080
rect 42618 33046 42652 33080
rect 42708 33046 42742 33080
rect 42168 32956 42202 32990
rect 42258 32956 42292 32990
rect 42348 32956 42382 32990
rect 42438 32956 42472 32990
rect 42528 32956 42562 32990
rect 42618 32956 42652 32990
rect 42708 32956 42742 32990
rect 42168 32866 42202 32900
rect 42258 32866 42292 32900
rect 42348 32866 42382 32900
rect 42438 32866 42472 32900
rect 42528 32866 42562 32900
rect 42618 32866 42652 32900
rect 42708 32866 42742 32900
rect 42168 32776 42202 32810
rect 42258 32776 42292 32810
rect 42348 32776 42382 32810
rect 42438 32776 42472 32810
rect 42528 32776 42562 32810
rect 42618 32776 42652 32810
rect 42708 32776 42742 32810
rect 42168 32686 42202 32720
rect 42258 32686 42292 32720
rect 42348 32686 42382 32720
rect 42438 32686 42472 32720
rect 42528 32686 42562 32720
rect 42618 32686 42652 32720
rect 42708 32686 42742 32720
rect 43508 33226 43542 33260
rect 43598 33226 43632 33260
rect 43688 33226 43722 33260
rect 43778 33226 43812 33260
rect 43868 33226 43902 33260
rect 43958 33226 43992 33260
rect 44048 33226 44082 33260
rect 43508 33136 43542 33170
rect 43598 33136 43632 33170
rect 43688 33136 43722 33170
rect 43778 33136 43812 33170
rect 43868 33136 43902 33170
rect 43958 33136 43992 33170
rect 44048 33136 44082 33170
rect 43508 33046 43542 33080
rect 43598 33046 43632 33080
rect 43688 33046 43722 33080
rect 43778 33046 43812 33080
rect 43868 33046 43902 33080
rect 43958 33046 43992 33080
rect 44048 33046 44082 33080
rect 43508 32956 43542 32990
rect 43598 32956 43632 32990
rect 43688 32956 43722 32990
rect 43778 32956 43812 32990
rect 43868 32956 43902 32990
rect 43958 32956 43992 32990
rect 44048 32956 44082 32990
rect 43508 32866 43542 32900
rect 43598 32866 43632 32900
rect 43688 32866 43722 32900
rect 43778 32866 43812 32900
rect 43868 32866 43902 32900
rect 43958 32866 43992 32900
rect 44048 32866 44082 32900
rect 43508 32776 43542 32810
rect 43598 32776 43632 32810
rect 43688 32776 43722 32810
rect 43778 32776 43812 32810
rect 43868 32776 43902 32810
rect 43958 32776 43992 32810
rect 44048 32776 44082 32810
rect 43508 32686 43542 32720
rect 43598 32686 43632 32720
rect 43688 32686 43722 32720
rect 43778 32686 43812 32720
rect 43868 32686 43902 32720
rect 43958 32686 43992 32720
rect 44048 32686 44082 32720
rect 44848 33226 44882 33260
rect 44938 33226 44972 33260
rect 45028 33226 45062 33260
rect 45118 33226 45152 33260
rect 45208 33226 45242 33260
rect 45298 33226 45332 33260
rect 45388 33226 45422 33260
rect 44848 33136 44882 33170
rect 44938 33136 44972 33170
rect 45028 33136 45062 33170
rect 45118 33136 45152 33170
rect 45208 33136 45242 33170
rect 45298 33136 45332 33170
rect 45388 33136 45422 33170
rect 44848 33046 44882 33080
rect 44938 33046 44972 33080
rect 45028 33046 45062 33080
rect 45118 33046 45152 33080
rect 45208 33046 45242 33080
rect 45298 33046 45332 33080
rect 45388 33046 45422 33080
rect 44848 32956 44882 32990
rect 44938 32956 44972 32990
rect 45028 32956 45062 32990
rect 45118 32956 45152 32990
rect 45208 32956 45242 32990
rect 45298 32956 45332 32990
rect 45388 32956 45422 32990
rect 44848 32866 44882 32900
rect 44938 32866 44972 32900
rect 45028 32866 45062 32900
rect 45118 32866 45152 32900
rect 45208 32866 45242 32900
rect 45298 32866 45332 32900
rect 45388 32866 45422 32900
rect 44848 32776 44882 32810
rect 44938 32776 44972 32810
rect 45028 32776 45062 32810
rect 45118 32776 45152 32810
rect 45208 32776 45242 32810
rect 45298 32776 45332 32810
rect 45388 32776 45422 32810
rect 44848 32686 44882 32720
rect 44938 32686 44972 32720
rect 45028 32686 45062 32720
rect 45118 32686 45152 32720
rect 45208 32686 45242 32720
rect 45298 32686 45332 32720
rect 45388 32686 45422 32720
rect 46188 33226 46222 33260
rect 46278 33226 46312 33260
rect 46368 33226 46402 33260
rect 46458 33226 46492 33260
rect 46548 33226 46582 33260
rect 46638 33226 46672 33260
rect 46728 33226 46762 33260
rect 46188 33136 46222 33170
rect 46278 33136 46312 33170
rect 46368 33136 46402 33170
rect 46458 33136 46492 33170
rect 46548 33136 46582 33170
rect 46638 33136 46672 33170
rect 46728 33136 46762 33170
rect 46188 33046 46222 33080
rect 46278 33046 46312 33080
rect 46368 33046 46402 33080
rect 46458 33046 46492 33080
rect 46548 33046 46582 33080
rect 46638 33046 46672 33080
rect 46728 33046 46762 33080
rect 46188 32956 46222 32990
rect 46278 32956 46312 32990
rect 46368 32956 46402 32990
rect 46458 32956 46492 32990
rect 46548 32956 46582 32990
rect 46638 32956 46672 32990
rect 46728 32956 46762 32990
rect 46188 32866 46222 32900
rect 46278 32866 46312 32900
rect 46368 32866 46402 32900
rect 46458 32866 46492 32900
rect 46548 32866 46582 32900
rect 46638 32866 46672 32900
rect 46728 32866 46762 32900
rect 46188 32776 46222 32810
rect 46278 32776 46312 32810
rect 46368 32776 46402 32810
rect 46458 32776 46492 32810
rect 46548 32776 46582 32810
rect 46638 32776 46672 32810
rect 46728 32776 46762 32810
rect 46188 32686 46222 32720
rect 46278 32686 46312 32720
rect 46368 32686 46402 32720
rect 46458 32686 46492 32720
rect 46548 32686 46582 32720
rect 46638 32686 46672 32720
rect 46728 32686 46762 32720
rect 47528 33226 47562 33260
rect 47618 33226 47652 33260
rect 47708 33226 47742 33260
rect 47798 33226 47832 33260
rect 47888 33226 47922 33260
rect 47978 33226 48012 33260
rect 48068 33226 48102 33260
rect 47528 33136 47562 33170
rect 47618 33136 47652 33170
rect 47708 33136 47742 33170
rect 47798 33136 47832 33170
rect 47888 33136 47922 33170
rect 47978 33136 48012 33170
rect 48068 33136 48102 33170
rect 47528 33046 47562 33080
rect 47618 33046 47652 33080
rect 47708 33046 47742 33080
rect 47798 33046 47832 33080
rect 47888 33046 47922 33080
rect 47978 33046 48012 33080
rect 48068 33046 48102 33080
rect 47528 32956 47562 32990
rect 47618 32956 47652 32990
rect 47708 32956 47742 32990
rect 47798 32956 47832 32990
rect 47888 32956 47922 32990
rect 47978 32956 48012 32990
rect 48068 32956 48102 32990
rect 47528 32866 47562 32900
rect 47618 32866 47652 32900
rect 47708 32866 47742 32900
rect 47798 32866 47832 32900
rect 47888 32866 47922 32900
rect 47978 32866 48012 32900
rect 48068 32866 48102 32900
rect 47528 32776 47562 32810
rect 47618 32776 47652 32810
rect 47708 32776 47742 32810
rect 47798 32776 47832 32810
rect 47888 32776 47922 32810
rect 47978 32776 48012 32810
rect 48068 32776 48102 32810
rect 47528 32686 47562 32720
rect 47618 32686 47652 32720
rect 47708 32686 47742 32720
rect 47798 32686 47832 32720
rect 47888 32686 47922 32720
rect 47978 32686 48012 32720
rect 48068 32686 48102 32720
rect 48868 33226 48902 33260
rect 48958 33226 48992 33260
rect 49048 33226 49082 33260
rect 49138 33226 49172 33260
rect 49228 33226 49262 33260
rect 49318 33226 49352 33260
rect 49408 33226 49442 33260
rect 48868 33136 48902 33170
rect 48958 33136 48992 33170
rect 49048 33136 49082 33170
rect 49138 33136 49172 33170
rect 49228 33136 49262 33170
rect 49318 33136 49352 33170
rect 49408 33136 49442 33170
rect 48868 33046 48902 33080
rect 48958 33046 48992 33080
rect 49048 33046 49082 33080
rect 49138 33046 49172 33080
rect 49228 33046 49262 33080
rect 49318 33046 49352 33080
rect 49408 33046 49442 33080
rect 48868 32956 48902 32990
rect 48958 32956 48992 32990
rect 49048 32956 49082 32990
rect 49138 32956 49172 32990
rect 49228 32956 49262 32990
rect 49318 32956 49352 32990
rect 49408 32956 49442 32990
rect 48868 32866 48902 32900
rect 48958 32866 48992 32900
rect 49048 32866 49082 32900
rect 49138 32866 49172 32900
rect 49228 32866 49262 32900
rect 49318 32866 49352 32900
rect 49408 32866 49442 32900
rect 48868 32776 48902 32810
rect 48958 32776 48992 32810
rect 49048 32776 49082 32810
rect 49138 32776 49172 32810
rect 49228 32776 49262 32810
rect 49318 32776 49352 32810
rect 49408 32776 49442 32810
rect 48868 32686 48902 32720
rect 48958 32686 48992 32720
rect 49048 32686 49082 32720
rect 49138 32686 49172 32720
rect 49228 32686 49262 32720
rect 49318 32686 49352 32720
rect 49408 32686 49442 32720
rect 50208 33226 50242 33260
rect 50298 33226 50332 33260
rect 50388 33226 50422 33260
rect 50478 33226 50512 33260
rect 50568 33226 50602 33260
rect 50658 33226 50692 33260
rect 50748 33226 50782 33260
rect 50208 33136 50242 33170
rect 50298 33136 50332 33170
rect 50388 33136 50422 33170
rect 50478 33136 50512 33170
rect 50568 33136 50602 33170
rect 50658 33136 50692 33170
rect 50748 33136 50782 33170
rect 50208 33046 50242 33080
rect 50298 33046 50332 33080
rect 50388 33046 50422 33080
rect 50478 33046 50512 33080
rect 50568 33046 50602 33080
rect 50658 33046 50692 33080
rect 50748 33046 50782 33080
rect 50208 32956 50242 32990
rect 50298 32956 50332 32990
rect 50388 32956 50422 32990
rect 50478 32956 50512 32990
rect 50568 32956 50602 32990
rect 50658 32956 50692 32990
rect 50748 32956 50782 32990
rect 50208 32866 50242 32900
rect 50298 32866 50332 32900
rect 50388 32866 50422 32900
rect 50478 32866 50512 32900
rect 50568 32866 50602 32900
rect 50658 32866 50692 32900
rect 50748 32866 50782 32900
rect 50208 32776 50242 32810
rect 50298 32776 50332 32810
rect 50388 32776 50422 32810
rect 50478 32776 50512 32810
rect 50568 32776 50602 32810
rect 50658 32776 50692 32810
rect 50748 32776 50782 32810
rect 50208 32686 50242 32720
rect 50298 32686 50332 32720
rect 50388 32686 50422 32720
rect 50478 32686 50512 32720
rect 50568 32686 50602 32720
rect 50658 32686 50692 32720
rect 50748 32686 50782 32720
rect 51548 33226 51582 33260
rect 51638 33226 51672 33260
rect 51728 33226 51762 33260
rect 51818 33226 51852 33260
rect 51908 33226 51942 33260
rect 51998 33226 52032 33260
rect 52088 33226 52122 33260
rect 51548 33136 51582 33170
rect 51638 33136 51672 33170
rect 51728 33136 51762 33170
rect 51818 33136 51852 33170
rect 51908 33136 51942 33170
rect 51998 33136 52032 33170
rect 52088 33136 52122 33170
rect 51548 33046 51582 33080
rect 51638 33046 51672 33080
rect 51728 33046 51762 33080
rect 51818 33046 51852 33080
rect 51908 33046 51942 33080
rect 51998 33046 52032 33080
rect 52088 33046 52122 33080
rect 51548 32956 51582 32990
rect 51638 32956 51672 32990
rect 51728 32956 51762 32990
rect 51818 32956 51852 32990
rect 51908 32956 51942 32990
rect 51998 32956 52032 32990
rect 52088 32956 52122 32990
rect 51548 32866 51582 32900
rect 51638 32866 51672 32900
rect 51728 32866 51762 32900
rect 51818 32866 51852 32900
rect 51908 32866 51942 32900
rect 51998 32866 52032 32900
rect 52088 32866 52122 32900
rect 51548 32776 51582 32810
rect 51638 32776 51672 32810
rect 51728 32776 51762 32810
rect 51818 32776 51852 32810
rect 51908 32776 51942 32810
rect 51998 32776 52032 32810
rect 52088 32776 52122 32810
rect 51548 32686 51582 32720
rect 51638 32686 51672 32720
rect 51728 32686 51762 32720
rect 51818 32686 51852 32720
rect 51908 32686 51942 32720
rect 51998 32686 52032 32720
rect 52088 32686 52122 32720
rect 37519 29867 37553 29901
rect 37519 29799 37553 29833
rect 37519 29731 37553 29765
rect 37519 29663 37553 29697
rect 37519 29595 37553 29629
rect 37519 29527 37553 29561
rect 37519 29459 37553 29493
rect 37519 29391 37553 29425
rect 37519 29323 37553 29357
rect 37519 29255 37553 29289
rect 37519 29187 37553 29221
rect 37519 29119 37553 29153
rect 37519 29051 37553 29085
rect 37519 28983 37553 29017
rect 37519 28915 37553 28949
rect 37519 28847 37553 28881
rect 37519 28779 37553 28813
rect 37519 28711 37553 28745
rect 37519 28643 37553 28677
rect 37977 29867 38011 29901
rect 37977 29799 38011 29833
rect 37977 29731 38011 29765
rect 37977 29663 38011 29697
rect 37977 29595 38011 29629
rect 37977 29527 38011 29561
rect 37977 29459 38011 29493
rect 37977 29391 38011 29425
rect 37977 29323 38011 29357
rect 37977 29255 38011 29289
rect 37977 29187 38011 29221
rect 37977 29119 38011 29153
rect 37977 29051 38011 29085
rect 37977 28983 38011 29017
rect 37977 28915 38011 28949
rect 37977 28847 38011 28881
rect 37977 28779 38011 28813
rect 37977 28711 38011 28745
rect 37977 28643 38011 28677
rect 38435 29867 38469 29901
rect 38435 29799 38469 29833
rect 38435 29731 38469 29765
rect 38435 29663 38469 29697
rect 38435 29595 38469 29629
rect 38435 29527 38469 29561
rect 38435 29459 38469 29493
rect 38435 29391 38469 29425
rect 38435 29323 38469 29357
rect 38435 29255 38469 29289
rect 38435 29187 38469 29221
rect 38435 29119 38469 29153
rect 38435 29051 38469 29085
rect 38435 28983 38469 29017
rect 38435 28915 38469 28949
rect 38435 28847 38469 28881
rect 38435 28779 38469 28813
rect 38435 28711 38469 28745
rect 38435 28643 38469 28677
rect 38893 29867 38927 29901
rect 38893 29799 38927 29833
rect 38893 29731 38927 29765
rect 38893 29663 38927 29697
rect 38893 29595 38927 29629
rect 38893 29527 38927 29561
rect 38893 29459 38927 29493
rect 38893 29391 38927 29425
rect 38893 29323 38927 29357
rect 38893 29255 38927 29289
rect 38893 29187 38927 29221
rect 38893 29119 38927 29153
rect 38893 29051 38927 29085
rect 38893 28983 38927 29017
rect 38893 28915 38927 28949
rect 38893 28847 38927 28881
rect 38893 28779 38927 28813
rect 38893 28711 38927 28745
rect 38893 28643 38927 28677
rect 39351 29867 39385 29901
rect 39351 29799 39385 29833
rect 39351 29731 39385 29765
rect 39351 29663 39385 29697
rect 39351 29595 39385 29629
rect 39351 29527 39385 29561
rect 39351 29459 39385 29493
rect 39351 29391 39385 29425
rect 39351 29323 39385 29357
rect 39351 29255 39385 29289
rect 39351 29187 39385 29221
rect 39351 29119 39385 29153
rect 39351 29051 39385 29085
rect 39351 28983 39385 29017
rect 39351 28915 39385 28949
rect 39351 28847 39385 28881
rect 39351 28779 39385 28813
rect 39351 28711 39385 28745
rect 39351 28643 39385 28677
rect 39809 29867 39843 29901
rect 39809 29799 39843 29833
rect 39809 29731 39843 29765
rect 39809 29663 39843 29697
rect 39809 29595 39843 29629
rect 39809 29527 39843 29561
rect 39809 29459 39843 29493
rect 39809 29391 39843 29425
rect 39809 29323 39843 29357
rect 39809 29255 39843 29289
rect 39809 29187 39843 29221
rect 39809 29119 39843 29153
rect 39809 29051 39843 29085
rect 39809 28983 39843 29017
rect 39809 28915 39843 28949
rect 39809 28847 39843 28881
rect 39809 28779 39843 28813
rect 39809 28711 39843 28745
rect 39809 28643 39843 28677
rect 40267 29867 40301 29901
rect 40267 29799 40301 29833
rect 40267 29731 40301 29765
rect 40267 29663 40301 29697
rect 40267 29595 40301 29629
rect 40267 29527 40301 29561
rect 40267 29459 40301 29493
rect 40267 29391 40301 29425
rect 40267 29323 40301 29357
rect 40267 29255 40301 29289
rect 40267 29187 40301 29221
rect 40267 29119 40301 29153
rect 40267 29051 40301 29085
rect 40267 28983 40301 29017
rect 40267 28915 40301 28949
rect 40267 28847 40301 28881
rect 40267 28779 40301 28813
rect 40267 28711 40301 28745
rect 40267 28643 40301 28677
rect 42168 29466 42202 29500
rect 42258 29466 42292 29500
rect 42348 29466 42382 29500
rect 42438 29466 42472 29500
rect 42528 29466 42562 29500
rect 42618 29466 42652 29500
rect 42708 29466 42742 29500
rect 42168 29376 42202 29410
rect 42258 29376 42292 29410
rect 42348 29376 42382 29410
rect 42438 29376 42472 29410
rect 42528 29376 42562 29410
rect 42618 29376 42652 29410
rect 42708 29376 42742 29410
rect 42168 29286 42202 29320
rect 42258 29286 42292 29320
rect 42348 29286 42382 29320
rect 42438 29286 42472 29320
rect 42528 29286 42562 29320
rect 42618 29286 42652 29320
rect 42708 29286 42742 29320
rect 42168 29196 42202 29230
rect 42258 29196 42292 29230
rect 42348 29196 42382 29230
rect 42438 29196 42472 29230
rect 42528 29196 42562 29230
rect 42618 29196 42652 29230
rect 42708 29196 42742 29230
rect 42168 29106 42202 29140
rect 42258 29106 42292 29140
rect 42348 29106 42382 29140
rect 42438 29106 42472 29140
rect 42528 29106 42562 29140
rect 42618 29106 42652 29140
rect 42708 29106 42742 29140
rect 42168 29016 42202 29050
rect 42258 29016 42292 29050
rect 42348 29016 42382 29050
rect 42438 29016 42472 29050
rect 42528 29016 42562 29050
rect 42618 29016 42652 29050
rect 42708 29016 42742 29050
rect 42168 28926 42202 28960
rect 42258 28926 42292 28960
rect 42348 28926 42382 28960
rect 42438 28926 42472 28960
rect 42528 28926 42562 28960
rect 42618 28926 42652 28960
rect 42708 28926 42742 28960
rect 43508 29466 43542 29500
rect 43598 29466 43632 29500
rect 43688 29466 43722 29500
rect 43778 29466 43812 29500
rect 43868 29466 43902 29500
rect 43958 29466 43992 29500
rect 44048 29466 44082 29500
rect 43508 29376 43542 29410
rect 43598 29376 43632 29410
rect 43688 29376 43722 29410
rect 43778 29376 43812 29410
rect 43868 29376 43902 29410
rect 43958 29376 43992 29410
rect 44048 29376 44082 29410
rect 43508 29286 43542 29320
rect 43598 29286 43632 29320
rect 43688 29286 43722 29320
rect 43778 29286 43812 29320
rect 43868 29286 43902 29320
rect 43958 29286 43992 29320
rect 44048 29286 44082 29320
rect 43508 29196 43542 29230
rect 43598 29196 43632 29230
rect 43688 29196 43722 29230
rect 43778 29196 43812 29230
rect 43868 29196 43902 29230
rect 43958 29196 43992 29230
rect 44048 29196 44082 29230
rect 43508 29106 43542 29140
rect 43598 29106 43632 29140
rect 43688 29106 43722 29140
rect 43778 29106 43812 29140
rect 43868 29106 43902 29140
rect 43958 29106 43992 29140
rect 44048 29106 44082 29140
rect 43508 29016 43542 29050
rect 43598 29016 43632 29050
rect 43688 29016 43722 29050
rect 43778 29016 43812 29050
rect 43868 29016 43902 29050
rect 43958 29016 43992 29050
rect 44048 29016 44082 29050
rect 43508 28926 43542 28960
rect 43598 28926 43632 28960
rect 43688 28926 43722 28960
rect 43778 28926 43812 28960
rect 43868 28926 43902 28960
rect 43958 28926 43992 28960
rect 44048 28926 44082 28960
rect 44848 29466 44882 29500
rect 44938 29466 44972 29500
rect 45028 29466 45062 29500
rect 45118 29466 45152 29500
rect 45208 29466 45242 29500
rect 45298 29466 45332 29500
rect 45388 29466 45422 29500
rect 44848 29376 44882 29410
rect 44938 29376 44972 29410
rect 45028 29376 45062 29410
rect 45118 29376 45152 29410
rect 45208 29376 45242 29410
rect 45298 29376 45332 29410
rect 45388 29376 45422 29410
rect 44848 29286 44882 29320
rect 44938 29286 44972 29320
rect 45028 29286 45062 29320
rect 45118 29286 45152 29320
rect 45208 29286 45242 29320
rect 45298 29286 45332 29320
rect 45388 29286 45422 29320
rect 44848 29196 44882 29230
rect 44938 29196 44972 29230
rect 45028 29196 45062 29230
rect 45118 29196 45152 29230
rect 45208 29196 45242 29230
rect 45298 29196 45332 29230
rect 45388 29196 45422 29230
rect 44848 29106 44882 29140
rect 44938 29106 44972 29140
rect 45028 29106 45062 29140
rect 45118 29106 45152 29140
rect 45208 29106 45242 29140
rect 45298 29106 45332 29140
rect 45388 29106 45422 29140
rect 44848 29016 44882 29050
rect 44938 29016 44972 29050
rect 45028 29016 45062 29050
rect 45118 29016 45152 29050
rect 45208 29016 45242 29050
rect 45298 29016 45332 29050
rect 45388 29016 45422 29050
rect 44848 28926 44882 28960
rect 44938 28926 44972 28960
rect 45028 28926 45062 28960
rect 45118 28926 45152 28960
rect 45208 28926 45242 28960
rect 45298 28926 45332 28960
rect 45388 28926 45422 28960
rect 46188 29466 46222 29500
rect 46278 29466 46312 29500
rect 46368 29466 46402 29500
rect 46458 29466 46492 29500
rect 46548 29466 46582 29500
rect 46638 29466 46672 29500
rect 46728 29466 46762 29500
rect 46188 29376 46222 29410
rect 46278 29376 46312 29410
rect 46368 29376 46402 29410
rect 46458 29376 46492 29410
rect 46548 29376 46582 29410
rect 46638 29376 46672 29410
rect 46728 29376 46762 29410
rect 46188 29286 46222 29320
rect 46278 29286 46312 29320
rect 46368 29286 46402 29320
rect 46458 29286 46492 29320
rect 46548 29286 46582 29320
rect 46638 29286 46672 29320
rect 46728 29286 46762 29320
rect 46188 29196 46222 29230
rect 46278 29196 46312 29230
rect 46368 29196 46402 29230
rect 46458 29196 46492 29230
rect 46548 29196 46582 29230
rect 46638 29196 46672 29230
rect 46728 29196 46762 29230
rect 46188 29106 46222 29140
rect 46278 29106 46312 29140
rect 46368 29106 46402 29140
rect 46458 29106 46492 29140
rect 46548 29106 46582 29140
rect 46638 29106 46672 29140
rect 46728 29106 46762 29140
rect 46188 29016 46222 29050
rect 46278 29016 46312 29050
rect 46368 29016 46402 29050
rect 46458 29016 46492 29050
rect 46548 29016 46582 29050
rect 46638 29016 46672 29050
rect 46728 29016 46762 29050
rect 46188 28926 46222 28960
rect 46278 28926 46312 28960
rect 46368 28926 46402 28960
rect 46458 28926 46492 28960
rect 46548 28926 46582 28960
rect 46638 28926 46672 28960
rect 46728 28926 46762 28960
rect 47528 29466 47562 29500
rect 47618 29466 47652 29500
rect 47708 29466 47742 29500
rect 47798 29466 47832 29500
rect 47888 29466 47922 29500
rect 47978 29466 48012 29500
rect 48068 29466 48102 29500
rect 47528 29376 47562 29410
rect 47618 29376 47652 29410
rect 47708 29376 47742 29410
rect 47798 29376 47832 29410
rect 47888 29376 47922 29410
rect 47978 29376 48012 29410
rect 48068 29376 48102 29410
rect 47528 29286 47562 29320
rect 47618 29286 47652 29320
rect 47708 29286 47742 29320
rect 47798 29286 47832 29320
rect 47888 29286 47922 29320
rect 47978 29286 48012 29320
rect 48068 29286 48102 29320
rect 47528 29196 47562 29230
rect 47618 29196 47652 29230
rect 47708 29196 47742 29230
rect 47798 29196 47832 29230
rect 47888 29196 47922 29230
rect 47978 29196 48012 29230
rect 48068 29196 48102 29230
rect 47528 29106 47562 29140
rect 47618 29106 47652 29140
rect 47708 29106 47742 29140
rect 47798 29106 47832 29140
rect 47888 29106 47922 29140
rect 47978 29106 48012 29140
rect 48068 29106 48102 29140
rect 47528 29016 47562 29050
rect 47618 29016 47652 29050
rect 47708 29016 47742 29050
rect 47798 29016 47832 29050
rect 47888 29016 47922 29050
rect 47978 29016 48012 29050
rect 48068 29016 48102 29050
rect 47528 28926 47562 28960
rect 47618 28926 47652 28960
rect 47708 28926 47742 28960
rect 47798 28926 47832 28960
rect 47888 28926 47922 28960
rect 47978 28926 48012 28960
rect 48068 28926 48102 28960
rect 48868 29466 48902 29500
rect 48958 29466 48992 29500
rect 49048 29466 49082 29500
rect 49138 29466 49172 29500
rect 49228 29466 49262 29500
rect 49318 29466 49352 29500
rect 49408 29466 49442 29500
rect 48868 29376 48902 29410
rect 48958 29376 48992 29410
rect 49048 29376 49082 29410
rect 49138 29376 49172 29410
rect 49228 29376 49262 29410
rect 49318 29376 49352 29410
rect 49408 29376 49442 29410
rect 48868 29286 48902 29320
rect 48958 29286 48992 29320
rect 49048 29286 49082 29320
rect 49138 29286 49172 29320
rect 49228 29286 49262 29320
rect 49318 29286 49352 29320
rect 49408 29286 49442 29320
rect 48868 29196 48902 29230
rect 48958 29196 48992 29230
rect 49048 29196 49082 29230
rect 49138 29196 49172 29230
rect 49228 29196 49262 29230
rect 49318 29196 49352 29230
rect 49408 29196 49442 29230
rect 48868 29106 48902 29140
rect 48958 29106 48992 29140
rect 49048 29106 49082 29140
rect 49138 29106 49172 29140
rect 49228 29106 49262 29140
rect 49318 29106 49352 29140
rect 49408 29106 49442 29140
rect 48868 29016 48902 29050
rect 48958 29016 48992 29050
rect 49048 29016 49082 29050
rect 49138 29016 49172 29050
rect 49228 29016 49262 29050
rect 49318 29016 49352 29050
rect 49408 29016 49442 29050
rect 48868 28926 48902 28960
rect 48958 28926 48992 28960
rect 49048 28926 49082 28960
rect 49138 28926 49172 28960
rect 49228 28926 49262 28960
rect 49318 28926 49352 28960
rect 49408 28926 49442 28960
rect 50208 29466 50242 29500
rect 50298 29466 50332 29500
rect 50388 29466 50422 29500
rect 50478 29466 50512 29500
rect 50568 29466 50602 29500
rect 50658 29466 50692 29500
rect 50748 29466 50782 29500
rect 50208 29376 50242 29410
rect 50298 29376 50332 29410
rect 50388 29376 50422 29410
rect 50478 29376 50512 29410
rect 50568 29376 50602 29410
rect 50658 29376 50692 29410
rect 50748 29376 50782 29410
rect 50208 29286 50242 29320
rect 50298 29286 50332 29320
rect 50388 29286 50422 29320
rect 50478 29286 50512 29320
rect 50568 29286 50602 29320
rect 50658 29286 50692 29320
rect 50748 29286 50782 29320
rect 50208 29196 50242 29230
rect 50298 29196 50332 29230
rect 50388 29196 50422 29230
rect 50478 29196 50512 29230
rect 50568 29196 50602 29230
rect 50658 29196 50692 29230
rect 50748 29196 50782 29230
rect 50208 29106 50242 29140
rect 50298 29106 50332 29140
rect 50388 29106 50422 29140
rect 50478 29106 50512 29140
rect 50568 29106 50602 29140
rect 50658 29106 50692 29140
rect 50748 29106 50782 29140
rect 50208 29016 50242 29050
rect 50298 29016 50332 29050
rect 50388 29016 50422 29050
rect 50478 29016 50512 29050
rect 50568 29016 50602 29050
rect 50658 29016 50692 29050
rect 50748 29016 50782 29050
rect 50208 28926 50242 28960
rect 50298 28926 50332 28960
rect 50388 28926 50422 28960
rect 50478 28926 50512 28960
rect 50568 28926 50602 28960
rect 50658 28926 50692 28960
rect 50748 28926 50782 28960
rect 51548 29466 51582 29500
rect 51638 29466 51672 29500
rect 51728 29466 51762 29500
rect 51818 29466 51852 29500
rect 51908 29466 51942 29500
rect 51998 29466 52032 29500
rect 52088 29466 52122 29500
rect 51548 29376 51582 29410
rect 51638 29376 51672 29410
rect 51728 29376 51762 29410
rect 51818 29376 51852 29410
rect 51908 29376 51942 29410
rect 51998 29376 52032 29410
rect 52088 29376 52122 29410
rect 51548 29286 51582 29320
rect 51638 29286 51672 29320
rect 51728 29286 51762 29320
rect 51818 29286 51852 29320
rect 51908 29286 51942 29320
rect 51998 29286 52032 29320
rect 52088 29286 52122 29320
rect 51548 29196 51582 29230
rect 51638 29196 51672 29230
rect 51728 29196 51762 29230
rect 51818 29196 51852 29230
rect 51908 29196 51942 29230
rect 51998 29196 52032 29230
rect 52088 29196 52122 29230
rect 51548 29106 51582 29140
rect 51638 29106 51672 29140
rect 51728 29106 51762 29140
rect 51818 29106 51852 29140
rect 51908 29106 51942 29140
rect 51998 29106 52032 29140
rect 52088 29106 52122 29140
rect 51548 29016 51582 29050
rect 51638 29016 51672 29050
rect 51728 29016 51762 29050
rect 51818 29016 51852 29050
rect 51908 29016 51942 29050
rect 51998 29016 52032 29050
rect 52088 29016 52122 29050
rect 51548 28926 51582 28960
rect 51638 28926 51672 28960
rect 51728 28926 51762 28960
rect 51818 28926 51852 28960
rect 51908 28926 51942 28960
rect 51998 28926 52032 28960
rect 52088 28926 52122 28960
rect 24877 18587 24911 18621
rect 24877 18519 24911 18553
rect 24877 18451 24911 18485
rect 24877 18383 24911 18417
rect 24877 18315 24911 18349
rect 24877 18247 24911 18281
rect 24877 18179 24911 18213
rect 24877 18111 24911 18145
rect 24877 18043 24911 18077
rect 24877 17975 24911 18009
rect 24877 17907 24911 17941
rect 24877 17839 24911 17873
rect 24877 17771 24911 17805
rect 24877 17703 24911 17737
rect 24877 17635 24911 17669
rect 24877 17567 24911 17601
rect 24877 17499 24911 17533
rect 24877 17431 24911 17465
rect 24877 17363 24911 17397
rect 25335 18587 25369 18621
rect 25335 18519 25369 18553
rect 25335 18451 25369 18485
rect 25335 18383 25369 18417
rect 25335 18315 25369 18349
rect 25335 18247 25369 18281
rect 25335 18179 25369 18213
rect 25335 18111 25369 18145
rect 25335 18043 25369 18077
rect 25335 17975 25369 18009
rect 25335 17907 25369 17941
rect 25335 17839 25369 17873
rect 25335 17771 25369 17805
rect 25335 17703 25369 17737
rect 25335 17635 25369 17669
rect 25335 17567 25369 17601
rect 25335 17499 25369 17533
rect 25335 17431 25369 17465
rect 25335 17363 25369 17397
rect 25793 18587 25827 18621
rect 25793 18519 25827 18553
rect 25793 18451 25827 18485
rect 25793 18383 25827 18417
rect 25793 18315 25827 18349
rect 25793 18247 25827 18281
rect 25793 18179 25827 18213
rect 25793 18111 25827 18145
rect 25793 18043 25827 18077
rect 25793 17975 25827 18009
rect 25793 17907 25827 17941
rect 25793 17839 25827 17873
rect 25793 17771 25827 17805
rect 25793 17703 25827 17737
rect 25793 17635 25827 17669
rect 25793 17567 25827 17601
rect 25793 17499 25827 17533
rect 25793 17431 25827 17465
rect 25793 17363 25827 17397
rect 26251 18587 26285 18621
rect 26251 18519 26285 18553
rect 26251 18451 26285 18485
rect 26251 18383 26285 18417
rect 26251 18315 26285 18349
rect 26251 18247 26285 18281
rect 26251 18179 26285 18213
rect 26251 18111 26285 18145
rect 26251 18043 26285 18077
rect 26251 17975 26285 18009
rect 26251 17907 26285 17941
rect 26251 17839 26285 17873
rect 26251 17771 26285 17805
rect 26251 17703 26285 17737
rect 26251 17635 26285 17669
rect 26251 17567 26285 17601
rect 26251 17499 26285 17533
rect 26251 17431 26285 17465
rect 26251 17363 26285 17397
rect 26709 18587 26743 18621
rect 26709 18519 26743 18553
rect 26709 18451 26743 18485
rect 26709 18383 26743 18417
rect 26709 18315 26743 18349
rect 26709 18247 26743 18281
rect 26709 18179 26743 18213
rect 26709 18111 26743 18145
rect 26709 18043 26743 18077
rect 26709 17975 26743 18009
rect 26709 17907 26743 17941
rect 26709 17839 26743 17873
rect 26709 17771 26743 17805
rect 26709 17703 26743 17737
rect 26709 17635 26743 17669
rect 26709 17567 26743 17601
rect 26709 17499 26743 17533
rect 26709 17431 26743 17465
rect 26709 17363 26743 17397
rect 27167 18587 27201 18621
rect 27167 18519 27201 18553
rect 27167 18451 27201 18485
rect 27167 18383 27201 18417
rect 27167 18315 27201 18349
rect 27167 18247 27201 18281
rect 27167 18179 27201 18213
rect 27167 18111 27201 18145
rect 27167 18043 27201 18077
rect 27167 17975 27201 18009
rect 27167 17907 27201 17941
rect 27167 17839 27201 17873
rect 27167 17771 27201 17805
rect 27167 17703 27201 17737
rect 27167 17635 27201 17669
rect 27167 17567 27201 17601
rect 27167 17499 27201 17533
rect 27167 17431 27201 17465
rect 27167 17363 27201 17397
rect 27625 18587 27659 18621
rect 27625 18519 27659 18553
rect 27625 18451 27659 18485
rect 27625 18383 27659 18417
rect 27625 18315 27659 18349
rect 27625 18247 27659 18281
rect 27625 18179 27659 18213
rect 27625 18111 27659 18145
rect 27625 18043 27659 18077
rect 27625 17975 27659 18009
rect 27625 17907 27659 17941
rect 27625 17839 27659 17873
rect 27625 17771 27659 17805
rect 27625 17703 27659 17737
rect 27625 17635 27659 17669
rect 27625 17567 27659 17601
rect 27625 17499 27659 17533
rect 27625 17431 27659 17465
rect 27625 17363 27659 17397
rect 28083 18587 28117 18621
rect 28083 18519 28117 18553
rect 28083 18451 28117 18485
rect 28083 18383 28117 18417
rect 28083 18315 28117 18349
rect 28083 18247 28117 18281
rect 28083 18179 28117 18213
rect 28083 18111 28117 18145
rect 28083 18043 28117 18077
rect 28083 17975 28117 18009
rect 28083 17907 28117 17941
rect 28083 17839 28117 17873
rect 28083 17771 28117 17805
rect 28083 17703 28117 17737
rect 28083 17635 28117 17669
rect 28083 17567 28117 17601
rect 28083 17499 28117 17533
rect 28083 17431 28117 17465
rect 28083 17363 28117 17397
rect 28541 18587 28575 18621
rect 28541 18519 28575 18553
rect 28541 18451 28575 18485
rect 28541 18383 28575 18417
rect 28541 18315 28575 18349
rect 28541 18247 28575 18281
rect 28541 18179 28575 18213
rect 28541 18111 28575 18145
rect 28541 18043 28575 18077
rect 28541 17975 28575 18009
rect 28541 17907 28575 17941
rect 28541 17839 28575 17873
rect 28541 17771 28575 17805
rect 28541 17703 28575 17737
rect 28541 17635 28575 17669
rect 28541 17567 28575 17601
rect 28541 17499 28575 17533
rect 28541 17431 28575 17465
rect 28541 17363 28575 17397
rect 28999 18587 29033 18621
rect 28999 18519 29033 18553
rect 28999 18451 29033 18485
rect 28999 18383 29033 18417
rect 28999 18315 29033 18349
rect 28999 18247 29033 18281
rect 28999 18179 29033 18213
rect 28999 18111 29033 18145
rect 28999 18043 29033 18077
rect 28999 17975 29033 18009
rect 28999 17907 29033 17941
rect 28999 17839 29033 17873
rect 28999 17771 29033 17805
rect 28999 17703 29033 17737
rect 28999 17635 29033 17669
rect 28999 17567 29033 17601
rect 28999 17499 29033 17533
rect 28999 17431 29033 17465
rect 28999 17363 29033 17397
rect 29457 18587 29491 18621
rect 29457 18519 29491 18553
rect 29457 18451 29491 18485
rect 29457 18383 29491 18417
rect 29457 18315 29491 18349
rect 29457 18247 29491 18281
rect 29457 18179 29491 18213
rect 29457 18111 29491 18145
rect 29457 18043 29491 18077
rect 29457 17975 29491 18009
rect 29457 17907 29491 17941
rect 29457 17839 29491 17873
rect 29457 17771 29491 17805
rect 29457 17703 29491 17737
rect 29457 17635 29491 17669
rect 29457 17567 29491 17601
rect 29457 17499 29491 17533
rect 29457 17431 29491 17465
rect 29457 17363 29491 17397
rect 29915 18587 29949 18621
rect 29915 18519 29949 18553
rect 29915 18451 29949 18485
rect 29915 18383 29949 18417
rect 29915 18315 29949 18349
rect 29915 18247 29949 18281
rect 29915 18179 29949 18213
rect 29915 18111 29949 18145
rect 29915 18043 29949 18077
rect 29915 17975 29949 18009
rect 29915 17907 29949 17941
rect 29915 17839 29949 17873
rect 29915 17771 29949 17805
rect 29915 17703 29949 17737
rect 29915 17635 29949 17669
rect 29915 17567 29949 17601
rect 29915 17499 29949 17533
rect 29915 17431 29949 17465
rect 29915 17363 29949 17397
rect 30373 18587 30407 18621
rect 30373 18519 30407 18553
rect 30373 18451 30407 18485
rect 30373 18383 30407 18417
rect 30373 18315 30407 18349
rect 30373 18247 30407 18281
rect 30373 18179 30407 18213
rect 30373 18111 30407 18145
rect 30373 18043 30407 18077
rect 30373 17975 30407 18009
rect 30373 17907 30407 17941
rect 30373 17839 30407 17873
rect 30373 17771 30407 17805
rect 30373 17703 30407 17737
rect 30373 17635 30407 17669
rect 30373 17567 30407 17601
rect 30373 17499 30407 17533
rect 30373 17431 30407 17465
rect 30373 17363 30407 17397
rect 30831 18587 30865 18621
rect 30831 18519 30865 18553
rect 30831 18451 30865 18485
rect 30831 18383 30865 18417
rect 30831 18315 30865 18349
rect 30831 18247 30865 18281
rect 30831 18179 30865 18213
rect 30831 18111 30865 18145
rect 30831 18043 30865 18077
rect 30831 17975 30865 18009
rect 30831 17907 30865 17941
rect 30831 17839 30865 17873
rect 30831 17771 30865 17805
rect 30831 17703 30865 17737
rect 30831 17635 30865 17669
rect 30831 17567 30865 17601
rect 30831 17499 30865 17533
rect 30831 17431 30865 17465
rect 30831 17363 30865 17397
rect 31289 18587 31323 18621
rect 31289 18519 31323 18553
rect 31289 18451 31323 18485
rect 31289 18383 31323 18417
rect 31289 18315 31323 18349
rect 31289 18247 31323 18281
rect 31289 18179 31323 18213
rect 31289 18111 31323 18145
rect 31289 18043 31323 18077
rect 31289 17975 31323 18009
rect 31289 17907 31323 17941
rect 31289 17839 31323 17873
rect 31289 17771 31323 17805
rect 31289 17703 31323 17737
rect 31289 17635 31323 17669
rect 31289 17567 31323 17601
rect 31289 17499 31323 17533
rect 31289 17431 31323 17465
rect 31289 17363 31323 17397
rect 31747 18587 31781 18621
rect 31747 18519 31781 18553
rect 31747 18451 31781 18485
rect 31747 18383 31781 18417
rect 31747 18315 31781 18349
rect 31747 18247 31781 18281
rect 31747 18179 31781 18213
rect 31747 18111 31781 18145
rect 31747 18043 31781 18077
rect 31747 17975 31781 18009
rect 31747 17907 31781 17941
rect 31747 17839 31781 17873
rect 31747 17771 31781 17805
rect 31747 17703 31781 17737
rect 31747 17635 31781 17669
rect 31747 17567 31781 17601
rect 31747 17499 31781 17533
rect 31747 17431 31781 17465
rect 31747 17363 31781 17397
rect 32205 18587 32239 18621
rect 32205 18519 32239 18553
rect 32205 18451 32239 18485
rect 32205 18383 32239 18417
rect 32205 18315 32239 18349
rect 32205 18247 32239 18281
rect 32205 18179 32239 18213
rect 32205 18111 32239 18145
rect 32205 18043 32239 18077
rect 32205 17975 32239 18009
rect 32205 17907 32239 17941
rect 32205 17839 32239 17873
rect 32205 17771 32239 17805
rect 32205 17703 32239 17737
rect 32205 17635 32239 17669
rect 32205 17567 32239 17601
rect 32205 17499 32239 17533
rect 32205 17431 32239 17465
rect 32205 17363 32239 17397
rect 32663 18587 32697 18621
rect 32663 18519 32697 18553
rect 32663 18451 32697 18485
rect 32663 18383 32697 18417
rect 32663 18315 32697 18349
rect 32663 18247 32697 18281
rect 32663 18179 32697 18213
rect 32663 18111 32697 18145
rect 32663 18043 32697 18077
rect 32663 17975 32697 18009
rect 32663 17907 32697 17941
rect 32663 17839 32697 17873
rect 32663 17771 32697 17805
rect 32663 17703 32697 17737
rect 32663 17635 32697 17669
rect 32663 17567 32697 17601
rect 32663 17499 32697 17533
rect 32663 17431 32697 17465
rect 32663 17363 32697 17397
rect 33121 18587 33155 18621
rect 33121 18519 33155 18553
rect 33121 18451 33155 18485
rect 33121 18383 33155 18417
rect 33121 18315 33155 18349
rect 33121 18247 33155 18281
rect 33121 18179 33155 18213
rect 33121 18111 33155 18145
rect 33121 18043 33155 18077
rect 33121 17975 33155 18009
rect 33121 17907 33155 17941
rect 33121 17839 33155 17873
rect 33121 17771 33155 17805
rect 33121 17703 33155 17737
rect 33121 17635 33155 17669
rect 33121 17567 33155 17601
rect 33121 17499 33155 17533
rect 33121 17431 33155 17465
rect 33121 17363 33155 17397
rect 33579 18587 33613 18621
rect 33579 18519 33613 18553
rect 33579 18451 33613 18485
rect 33579 18383 33613 18417
rect 33579 18315 33613 18349
rect 33579 18247 33613 18281
rect 33579 18179 33613 18213
rect 33579 18111 33613 18145
rect 33579 18043 33613 18077
rect 33579 17975 33613 18009
rect 33579 17907 33613 17941
rect 33579 17839 33613 17873
rect 33579 17771 33613 17805
rect 33579 17703 33613 17737
rect 33579 17635 33613 17669
rect 33579 17567 33613 17601
rect 33579 17499 33613 17533
rect 33579 17431 33613 17465
rect 33579 17363 33613 17397
rect 34037 18587 34071 18621
rect 34037 18519 34071 18553
rect 34037 18451 34071 18485
rect 34037 18383 34071 18417
rect 34037 18315 34071 18349
rect 34037 18247 34071 18281
rect 34037 18179 34071 18213
rect 34037 18111 34071 18145
rect 34037 18043 34071 18077
rect 34037 17975 34071 18009
rect 34037 17907 34071 17941
rect 34037 17839 34071 17873
rect 34037 17771 34071 17805
rect 34037 17703 34071 17737
rect 34037 17635 34071 17669
rect 34037 17567 34071 17601
rect 34037 17499 34071 17533
rect 34037 17431 34071 17465
rect 34037 17363 34071 17397
rect 34495 18587 34529 18621
rect 34495 18519 34529 18553
rect 34495 18451 34529 18485
rect 34495 18383 34529 18417
rect 34495 18315 34529 18349
rect 34495 18247 34529 18281
rect 34495 18179 34529 18213
rect 34495 18111 34529 18145
rect 34495 18043 34529 18077
rect 34495 17975 34529 18009
rect 34495 17907 34529 17941
rect 34495 17839 34529 17873
rect 34495 17771 34529 17805
rect 34495 17703 34529 17737
rect 34495 17635 34529 17669
rect 34495 17567 34529 17601
rect 34495 17499 34529 17533
rect 34495 17431 34529 17465
rect 34495 17363 34529 17397
rect 34953 18587 34987 18621
rect 34953 18519 34987 18553
rect 34953 18451 34987 18485
rect 34953 18383 34987 18417
rect 34953 18315 34987 18349
rect 34953 18247 34987 18281
rect 34953 18179 34987 18213
rect 34953 18111 34987 18145
rect 34953 18043 34987 18077
rect 34953 17975 34987 18009
rect 34953 17907 34987 17941
rect 34953 17839 34987 17873
rect 34953 17771 34987 17805
rect 34953 17703 34987 17737
rect 34953 17635 34987 17669
rect 34953 17567 34987 17601
rect 34953 17499 34987 17533
rect 34953 17431 34987 17465
rect 34953 17363 34987 17397
rect 35411 18587 35445 18621
rect 35411 18519 35445 18553
rect 35411 18451 35445 18485
rect 35411 18383 35445 18417
rect 35411 18315 35445 18349
rect 35411 18247 35445 18281
rect 35411 18179 35445 18213
rect 35411 18111 35445 18145
rect 35411 18043 35445 18077
rect 35411 17975 35445 18009
rect 35411 17907 35445 17941
rect 35411 17839 35445 17873
rect 35411 17771 35445 17805
rect 35411 17703 35445 17737
rect 35411 17635 35445 17669
rect 35411 17567 35445 17601
rect 35411 17499 35445 17533
rect 35411 17431 35445 17465
rect 35411 17363 35445 17397
rect 35869 18587 35903 18621
rect 35869 18519 35903 18553
rect 35869 18451 35903 18485
rect 35869 18383 35903 18417
rect 35869 18315 35903 18349
rect 35869 18247 35903 18281
rect 35869 18179 35903 18213
rect 35869 18111 35903 18145
rect 35869 18043 35903 18077
rect 35869 17975 35903 18009
rect 35869 17907 35903 17941
rect 35869 17839 35903 17873
rect 35869 17771 35903 17805
rect 35869 17703 35903 17737
rect 35869 17635 35903 17669
rect 35869 17567 35903 17601
rect 35869 17499 35903 17533
rect 35869 17431 35903 17465
rect 35869 17363 35903 17397
rect 36327 18587 36361 18621
rect 36327 18519 36361 18553
rect 36327 18451 36361 18485
rect 36327 18383 36361 18417
rect 36327 18315 36361 18349
rect 36327 18247 36361 18281
rect 36327 18179 36361 18213
rect 36327 18111 36361 18145
rect 36327 18043 36361 18077
rect 36327 17975 36361 18009
rect 36327 17907 36361 17941
rect 36327 17839 36361 17873
rect 36327 17771 36361 17805
rect 36327 17703 36361 17737
rect 36327 17635 36361 17669
rect 36327 17567 36361 17601
rect 36327 17499 36361 17533
rect 36327 17431 36361 17465
rect 36327 17363 36361 17397
rect 36785 18587 36819 18621
rect 36785 18519 36819 18553
rect 36785 18451 36819 18485
rect 36785 18383 36819 18417
rect 36785 18315 36819 18349
rect 36785 18247 36819 18281
rect 36785 18179 36819 18213
rect 36785 18111 36819 18145
rect 36785 18043 36819 18077
rect 36785 17975 36819 18009
rect 36785 17907 36819 17941
rect 36785 17839 36819 17873
rect 36785 17771 36819 17805
rect 36785 17703 36819 17737
rect 36785 17635 36819 17669
rect 36785 17567 36819 17601
rect 36785 17499 36819 17533
rect 36785 17431 36819 17465
rect 36785 17363 36819 17397
rect 37243 18587 37277 18621
rect 37243 18519 37277 18553
rect 37243 18451 37277 18485
rect 37243 18383 37277 18417
rect 37243 18315 37277 18349
rect 37243 18247 37277 18281
rect 37243 18179 37277 18213
rect 37243 18111 37277 18145
rect 37243 18043 37277 18077
rect 37243 17975 37277 18009
rect 37243 17907 37277 17941
rect 37243 17839 37277 17873
rect 37243 17771 37277 17805
rect 37243 17703 37277 17737
rect 37243 17635 37277 17669
rect 37243 17567 37277 17601
rect 37243 17499 37277 17533
rect 37243 17431 37277 17465
rect 37243 17363 37277 17397
rect 37701 18587 37735 18621
rect 37701 18519 37735 18553
rect 37701 18451 37735 18485
rect 37701 18383 37735 18417
rect 37701 18315 37735 18349
rect 37701 18247 37735 18281
rect 37701 18179 37735 18213
rect 37701 18111 37735 18145
rect 37701 18043 37735 18077
rect 37701 17975 37735 18009
rect 37701 17907 37735 17941
rect 37701 17839 37735 17873
rect 37701 17771 37735 17805
rect 37701 17703 37735 17737
rect 37701 17635 37735 17669
rect 37701 17567 37735 17601
rect 37701 17499 37735 17533
rect 37701 17431 37735 17465
rect 37701 17363 37735 17397
rect 38159 18587 38193 18621
rect 38159 18519 38193 18553
rect 38159 18451 38193 18485
rect 38159 18383 38193 18417
rect 38159 18315 38193 18349
rect 38159 18247 38193 18281
rect 38159 18179 38193 18213
rect 38159 18111 38193 18145
rect 38159 18043 38193 18077
rect 38159 17975 38193 18009
rect 38159 17907 38193 17941
rect 38159 17839 38193 17873
rect 38159 17771 38193 17805
rect 38159 17703 38193 17737
rect 38159 17635 38193 17669
rect 38159 17567 38193 17601
rect 38159 17499 38193 17533
rect 38159 17431 38193 17465
rect 38159 17363 38193 17397
rect 38617 18587 38651 18621
rect 38617 18519 38651 18553
rect 38617 18451 38651 18485
rect 38617 18383 38651 18417
rect 38617 18315 38651 18349
rect 38617 18247 38651 18281
rect 38617 18179 38651 18213
rect 38617 18111 38651 18145
rect 38617 18043 38651 18077
rect 38617 17975 38651 18009
rect 38617 17907 38651 17941
rect 38617 17839 38651 17873
rect 38617 17771 38651 17805
rect 38617 17703 38651 17737
rect 38617 17635 38651 17669
rect 38617 17567 38651 17601
rect 38617 17499 38651 17533
rect 38617 17431 38651 17465
rect 38617 17363 38651 17397
rect 39075 18587 39109 18621
rect 39075 18519 39109 18553
rect 39075 18451 39109 18485
rect 39075 18383 39109 18417
rect 39075 18315 39109 18349
rect 39075 18247 39109 18281
rect 39075 18179 39109 18213
rect 39075 18111 39109 18145
rect 39075 18043 39109 18077
rect 39075 17975 39109 18009
rect 39075 17907 39109 17941
rect 39075 17839 39109 17873
rect 39075 17771 39109 17805
rect 39075 17703 39109 17737
rect 39075 17635 39109 17669
rect 39075 17567 39109 17601
rect 39075 17499 39109 17533
rect 39075 17431 39109 17465
rect 39075 17363 39109 17397
rect 39533 18587 39567 18621
rect 39533 18519 39567 18553
rect 39533 18451 39567 18485
rect 39533 18383 39567 18417
rect 39533 18315 39567 18349
rect 39533 18247 39567 18281
rect 39533 18179 39567 18213
rect 39533 18111 39567 18145
rect 39533 18043 39567 18077
rect 39533 17975 39567 18009
rect 39533 17907 39567 17941
rect 39533 17839 39567 17873
rect 39533 17771 39567 17805
rect 39533 17703 39567 17737
rect 39533 17635 39567 17669
rect 39533 17567 39567 17601
rect 39533 17499 39567 17533
rect 39533 17431 39567 17465
rect 39533 17363 39567 17397
rect 39991 18587 40025 18621
rect 39991 18519 40025 18553
rect 39991 18451 40025 18485
rect 39991 18383 40025 18417
rect 39991 18315 40025 18349
rect 39991 18247 40025 18281
rect 39991 18179 40025 18213
rect 39991 18111 40025 18145
rect 39991 18043 40025 18077
rect 39991 17975 40025 18009
rect 39991 17907 40025 17941
rect 39991 17839 40025 17873
rect 39991 17771 40025 17805
rect 39991 17703 40025 17737
rect 39991 17635 40025 17669
rect 39991 17567 40025 17601
rect 39991 17499 40025 17533
rect 39991 17431 40025 17465
rect 39991 17363 40025 17397
rect 40449 18587 40483 18621
rect 40449 18519 40483 18553
rect 40449 18451 40483 18485
rect 40449 18383 40483 18417
rect 40449 18315 40483 18349
rect 40449 18247 40483 18281
rect 40449 18179 40483 18213
rect 40449 18111 40483 18145
rect 40449 18043 40483 18077
rect 40449 17975 40483 18009
rect 40449 17907 40483 17941
rect 40449 17839 40483 17873
rect 40449 17771 40483 17805
rect 40449 17703 40483 17737
rect 40449 17635 40483 17669
rect 40449 17567 40483 17601
rect 40449 17499 40483 17533
rect 40449 17431 40483 17465
rect 40449 17363 40483 17397
rect 40907 18587 40941 18621
rect 40907 18519 40941 18553
rect 40907 18451 40941 18485
rect 40907 18383 40941 18417
rect 40907 18315 40941 18349
rect 40907 18247 40941 18281
rect 40907 18179 40941 18213
rect 40907 18111 40941 18145
rect 40907 18043 40941 18077
rect 40907 17975 40941 18009
rect 40907 17907 40941 17941
rect 40907 17839 40941 17873
rect 40907 17771 40941 17805
rect 40907 17703 40941 17737
rect 40907 17635 40941 17669
rect 40907 17567 40941 17601
rect 40907 17499 40941 17533
rect 40907 17431 40941 17465
rect 40907 17363 40941 17397
rect 41365 18587 41399 18621
rect 41365 18519 41399 18553
rect 41365 18451 41399 18485
rect 41365 18383 41399 18417
rect 41365 18315 41399 18349
rect 41365 18247 41399 18281
rect 41365 18179 41399 18213
rect 41365 18111 41399 18145
rect 41365 18043 41399 18077
rect 41365 17975 41399 18009
rect 41365 17907 41399 17941
rect 41365 17839 41399 17873
rect 41365 17771 41399 17805
rect 41365 17703 41399 17737
rect 41365 17635 41399 17669
rect 41365 17567 41399 17601
rect 41365 17499 41399 17533
rect 41365 17431 41399 17465
rect 41365 17363 41399 17397
rect 41823 18587 41857 18621
rect 41823 18519 41857 18553
rect 41823 18451 41857 18485
rect 41823 18383 41857 18417
rect 41823 18315 41857 18349
rect 41823 18247 41857 18281
rect 41823 18179 41857 18213
rect 41823 18111 41857 18145
rect 41823 18043 41857 18077
rect 41823 17975 41857 18009
rect 41823 17907 41857 17941
rect 41823 17839 41857 17873
rect 41823 17771 41857 17805
rect 41823 17703 41857 17737
rect 41823 17635 41857 17669
rect 41823 17567 41857 17601
rect 41823 17499 41857 17533
rect 41823 17431 41857 17465
rect 41823 17363 41857 17397
rect 42281 18587 42315 18621
rect 42281 18519 42315 18553
rect 42281 18451 42315 18485
rect 42281 18383 42315 18417
rect 42281 18315 42315 18349
rect 42281 18247 42315 18281
rect 42281 18179 42315 18213
rect 42281 18111 42315 18145
rect 42281 18043 42315 18077
rect 42281 17975 42315 18009
rect 42281 17907 42315 17941
rect 42281 17839 42315 17873
rect 42281 17771 42315 17805
rect 42281 17703 42315 17737
rect 42281 17635 42315 17669
rect 42281 17567 42315 17601
rect 42281 17499 42315 17533
rect 42281 17431 42315 17465
rect 42281 17363 42315 17397
rect 42739 18587 42773 18621
rect 42739 18519 42773 18553
rect 42739 18451 42773 18485
rect 42739 18383 42773 18417
rect 42739 18315 42773 18349
rect 42739 18247 42773 18281
rect 42739 18179 42773 18213
rect 42739 18111 42773 18145
rect 42739 18043 42773 18077
rect 42739 17975 42773 18009
rect 42739 17907 42773 17941
rect 42739 17839 42773 17873
rect 42739 17771 42773 17805
rect 42739 17703 42773 17737
rect 42739 17635 42773 17669
rect 42739 17567 42773 17601
rect 42739 17499 42773 17533
rect 42739 17431 42773 17465
rect 42739 17363 42773 17397
rect 43197 18587 43231 18621
rect 43197 18519 43231 18553
rect 43197 18451 43231 18485
rect 43197 18383 43231 18417
rect 43197 18315 43231 18349
rect 43197 18247 43231 18281
rect 43197 18179 43231 18213
rect 43197 18111 43231 18145
rect 43197 18043 43231 18077
rect 43197 17975 43231 18009
rect 43197 17907 43231 17941
rect 43197 17839 43231 17873
rect 43197 17771 43231 17805
rect 43197 17703 43231 17737
rect 43197 17635 43231 17669
rect 43197 17567 43231 17601
rect 43197 17499 43231 17533
rect 43197 17431 43231 17465
rect 43197 17363 43231 17397
rect 43655 18587 43689 18621
rect 43655 18519 43689 18553
rect 43655 18451 43689 18485
rect 43655 18383 43689 18417
rect 43655 18315 43689 18349
rect 43655 18247 43689 18281
rect 43655 18179 43689 18213
rect 43655 18111 43689 18145
rect 43655 18043 43689 18077
rect 43655 17975 43689 18009
rect 43655 17907 43689 17941
rect 43655 17839 43689 17873
rect 43655 17771 43689 17805
rect 43655 17703 43689 17737
rect 43655 17635 43689 17669
rect 43655 17567 43689 17601
rect 43655 17499 43689 17533
rect 43655 17431 43689 17465
rect 43655 17363 43689 17397
rect 44113 18587 44147 18621
rect 44113 18519 44147 18553
rect 44113 18451 44147 18485
rect 44113 18383 44147 18417
rect 44113 18315 44147 18349
rect 44113 18247 44147 18281
rect 44113 18179 44147 18213
rect 44113 18111 44147 18145
rect 44113 18043 44147 18077
rect 44113 17975 44147 18009
rect 44113 17907 44147 17941
rect 44113 17839 44147 17873
rect 44113 17771 44147 17805
rect 44113 17703 44147 17737
rect 44113 17635 44147 17669
rect 44113 17567 44147 17601
rect 44113 17499 44147 17533
rect 44113 17431 44147 17465
rect 44113 17363 44147 17397
rect 44571 18587 44605 18621
rect 44571 18519 44605 18553
rect 44571 18451 44605 18485
rect 44571 18383 44605 18417
rect 44571 18315 44605 18349
rect 44571 18247 44605 18281
rect 44571 18179 44605 18213
rect 44571 18111 44605 18145
rect 44571 18043 44605 18077
rect 44571 17975 44605 18009
rect 44571 17907 44605 17941
rect 44571 17839 44605 17873
rect 44571 17771 44605 17805
rect 44571 17703 44605 17737
rect 44571 17635 44605 17669
rect 44571 17567 44605 17601
rect 44571 17499 44605 17533
rect 44571 17431 44605 17465
rect 44571 17363 44605 17397
rect 45029 18587 45063 18621
rect 45029 18519 45063 18553
rect 45029 18451 45063 18485
rect 45029 18383 45063 18417
rect 45029 18315 45063 18349
rect 45029 18247 45063 18281
rect 45029 18179 45063 18213
rect 45029 18111 45063 18145
rect 45029 18043 45063 18077
rect 45029 17975 45063 18009
rect 45029 17907 45063 17941
rect 45029 17839 45063 17873
rect 45029 17771 45063 17805
rect 45029 17703 45063 17737
rect 45029 17635 45063 17669
rect 45029 17567 45063 17601
rect 45029 17499 45063 17533
rect 45029 17431 45063 17465
rect 45029 17363 45063 17397
rect 45487 18587 45521 18621
rect 45487 18519 45521 18553
rect 45487 18451 45521 18485
rect 45487 18383 45521 18417
rect 45487 18315 45521 18349
rect 45487 18247 45521 18281
rect 45487 18179 45521 18213
rect 45487 18111 45521 18145
rect 45487 18043 45521 18077
rect 45487 17975 45521 18009
rect 45487 17907 45521 17941
rect 45487 17839 45521 17873
rect 45487 17771 45521 17805
rect 45487 17703 45521 17737
rect 45487 17635 45521 17669
rect 45487 17567 45521 17601
rect 45487 17499 45521 17533
rect 45487 17431 45521 17465
rect 45487 17363 45521 17397
rect 45945 18587 45979 18621
rect 45945 18519 45979 18553
rect 45945 18451 45979 18485
rect 45945 18383 45979 18417
rect 45945 18315 45979 18349
rect 45945 18247 45979 18281
rect 45945 18179 45979 18213
rect 45945 18111 45979 18145
rect 45945 18043 45979 18077
rect 45945 17975 45979 18009
rect 45945 17907 45979 17941
rect 45945 17839 45979 17873
rect 45945 17771 45979 17805
rect 45945 17703 45979 17737
rect 45945 17635 45979 17669
rect 45945 17567 45979 17601
rect 45945 17499 45979 17533
rect 45945 17431 45979 17465
rect 45945 17363 45979 17397
rect 46403 18587 46437 18621
rect 46403 18519 46437 18553
rect 46403 18451 46437 18485
rect 46403 18383 46437 18417
rect 46403 18315 46437 18349
rect 46403 18247 46437 18281
rect 46403 18179 46437 18213
rect 46403 18111 46437 18145
rect 46403 18043 46437 18077
rect 46403 17975 46437 18009
rect 46403 17907 46437 17941
rect 46403 17839 46437 17873
rect 46403 17771 46437 17805
rect 46403 17703 46437 17737
rect 46403 17635 46437 17669
rect 46403 17567 46437 17601
rect 46403 17499 46437 17533
rect 46403 17431 46437 17465
rect 46403 17363 46437 17397
rect 46861 18587 46895 18621
rect 46861 18519 46895 18553
rect 46861 18451 46895 18485
rect 46861 18383 46895 18417
rect 46861 18315 46895 18349
rect 46861 18247 46895 18281
rect 46861 18179 46895 18213
rect 46861 18111 46895 18145
rect 46861 18043 46895 18077
rect 46861 17975 46895 18009
rect 46861 17907 46895 17941
rect 46861 17839 46895 17873
rect 46861 17771 46895 17805
rect 46861 17703 46895 17737
rect 46861 17635 46895 17669
rect 46861 17567 46895 17601
rect 46861 17499 46895 17533
rect 46861 17431 46895 17465
rect 46861 17363 46895 17397
rect 47319 18587 47353 18621
rect 47319 18519 47353 18553
rect 47319 18451 47353 18485
rect 47319 18383 47353 18417
rect 47319 18315 47353 18349
rect 47319 18247 47353 18281
rect 47319 18179 47353 18213
rect 47319 18111 47353 18145
rect 47319 18043 47353 18077
rect 47319 17975 47353 18009
rect 47319 17907 47353 17941
rect 47319 17839 47353 17873
rect 47319 17771 47353 17805
rect 47319 17703 47353 17737
rect 47319 17635 47353 17669
rect 47319 17567 47353 17601
rect 47319 17499 47353 17533
rect 47319 17431 47353 17465
rect 47319 17363 47353 17397
rect 47777 18587 47811 18621
rect 47777 18519 47811 18553
rect 47777 18451 47811 18485
rect 47777 18383 47811 18417
rect 47777 18315 47811 18349
rect 47777 18247 47811 18281
rect 47777 18179 47811 18213
rect 47777 18111 47811 18145
rect 47777 18043 47811 18077
rect 47777 17975 47811 18009
rect 47777 17907 47811 17941
rect 47777 17839 47811 17873
rect 47777 17771 47811 17805
rect 47777 17703 47811 17737
rect 47777 17635 47811 17669
rect 47777 17567 47811 17601
rect 47777 17499 47811 17533
rect 47777 17431 47811 17465
rect 47777 17363 47811 17397
rect 48235 18587 48269 18621
rect 48235 18519 48269 18553
rect 48235 18451 48269 18485
rect 48235 18383 48269 18417
rect 48235 18315 48269 18349
rect 48235 18247 48269 18281
rect 48235 18179 48269 18213
rect 48235 18111 48269 18145
rect 48235 18043 48269 18077
rect 48235 17975 48269 18009
rect 48235 17907 48269 17941
rect 48235 17839 48269 17873
rect 48235 17771 48269 17805
rect 48235 17703 48269 17737
rect 48235 17635 48269 17669
rect 48235 17567 48269 17601
rect 48235 17499 48269 17533
rect 48235 17431 48269 17465
rect 48235 17363 48269 17397
rect 48693 18587 48727 18621
rect 48693 18519 48727 18553
rect 48693 18451 48727 18485
rect 48693 18383 48727 18417
rect 48693 18315 48727 18349
rect 48693 18247 48727 18281
rect 48693 18179 48727 18213
rect 48693 18111 48727 18145
rect 48693 18043 48727 18077
rect 48693 17975 48727 18009
rect 48693 17907 48727 17941
rect 48693 17839 48727 17873
rect 48693 17771 48727 17805
rect 48693 17703 48727 17737
rect 48693 17635 48727 17669
rect 48693 17567 48727 17601
rect 48693 17499 48727 17533
rect 48693 17431 48727 17465
rect 48693 17363 48727 17397
rect 49151 18587 49185 18621
rect 49151 18519 49185 18553
rect 49151 18451 49185 18485
rect 49151 18383 49185 18417
rect 49151 18315 49185 18349
rect 49151 18247 49185 18281
rect 49151 18179 49185 18213
rect 49151 18111 49185 18145
rect 49151 18043 49185 18077
rect 49151 17975 49185 18009
rect 49151 17907 49185 17941
rect 49151 17839 49185 17873
rect 49151 17771 49185 17805
rect 49151 17703 49185 17737
rect 49151 17635 49185 17669
rect 49151 17567 49185 17601
rect 49151 17499 49185 17533
rect 49151 17431 49185 17465
rect 49151 17363 49185 17397
rect 49609 18587 49643 18621
rect 49609 18519 49643 18553
rect 49609 18451 49643 18485
rect 49609 18383 49643 18417
rect 49609 18315 49643 18349
rect 49609 18247 49643 18281
rect 49609 18179 49643 18213
rect 49609 18111 49643 18145
rect 49609 18043 49643 18077
rect 49609 17975 49643 18009
rect 49609 17907 49643 17941
rect 49609 17839 49643 17873
rect 49609 17771 49643 17805
rect 49609 17703 49643 17737
rect 49609 17635 49643 17669
rect 49609 17567 49643 17601
rect 49609 17499 49643 17533
rect 49609 17431 49643 17465
rect 49609 17363 49643 17397
rect 50067 18587 50101 18621
rect 50067 18519 50101 18553
rect 50067 18451 50101 18485
rect 50067 18383 50101 18417
rect 50067 18315 50101 18349
rect 50067 18247 50101 18281
rect 50067 18179 50101 18213
rect 50067 18111 50101 18145
rect 50067 18043 50101 18077
rect 50067 17975 50101 18009
rect 50067 17907 50101 17941
rect 50067 17839 50101 17873
rect 50067 17771 50101 17805
rect 50067 17703 50101 17737
rect 50067 17635 50101 17669
rect 50067 17567 50101 17601
rect 50067 17499 50101 17533
rect 50067 17431 50101 17465
rect 50067 17363 50101 17397
rect 50525 18587 50559 18621
rect 50525 18519 50559 18553
rect 50525 18451 50559 18485
rect 50525 18383 50559 18417
rect 50525 18315 50559 18349
rect 50525 18247 50559 18281
rect 50525 18179 50559 18213
rect 50525 18111 50559 18145
rect 50525 18043 50559 18077
rect 50525 17975 50559 18009
rect 50525 17907 50559 17941
rect 50525 17839 50559 17873
rect 50525 17771 50559 17805
rect 50525 17703 50559 17737
rect 50525 17635 50559 17669
rect 50525 17567 50559 17601
rect 50525 17499 50559 17533
rect 50525 17431 50559 17465
rect 50525 17363 50559 17397
rect 50983 18587 51017 18621
rect 50983 18519 51017 18553
rect 50983 18451 51017 18485
rect 50983 18383 51017 18417
rect 50983 18315 51017 18349
rect 50983 18247 51017 18281
rect 50983 18179 51017 18213
rect 50983 18111 51017 18145
rect 50983 18043 51017 18077
rect 50983 17975 51017 18009
rect 50983 17907 51017 17941
rect 50983 17839 51017 17873
rect 50983 17771 51017 17805
rect 50983 17703 51017 17737
rect 50983 17635 51017 17669
rect 50983 17567 51017 17601
rect 50983 17499 51017 17533
rect 50983 17431 51017 17465
rect 50983 17363 51017 17397
rect 51441 18587 51475 18621
rect 51441 18519 51475 18553
rect 51441 18451 51475 18485
rect 51441 18383 51475 18417
rect 51441 18315 51475 18349
rect 51441 18247 51475 18281
rect 51441 18179 51475 18213
rect 51441 18111 51475 18145
rect 51441 18043 51475 18077
rect 51441 17975 51475 18009
rect 51441 17907 51475 17941
rect 51441 17839 51475 17873
rect 51441 17771 51475 17805
rect 51441 17703 51475 17737
rect 51441 17635 51475 17669
rect 51441 17567 51475 17601
rect 51441 17499 51475 17533
rect 51441 17431 51475 17465
rect 51441 17363 51475 17397
rect 51899 18587 51933 18621
rect 51899 18519 51933 18553
rect 51899 18451 51933 18485
rect 51899 18383 51933 18417
rect 51899 18315 51933 18349
rect 51899 18247 51933 18281
rect 51899 18179 51933 18213
rect 51899 18111 51933 18145
rect 51899 18043 51933 18077
rect 51899 17975 51933 18009
rect 51899 17907 51933 17941
rect 51899 17839 51933 17873
rect 51899 17771 51933 17805
rect 51899 17703 51933 17737
rect 51899 17635 51933 17669
rect 51899 17567 51933 17601
rect 51899 17499 51933 17533
rect 51899 17431 51933 17465
rect 51899 17363 51933 17397
rect 52357 18587 52391 18621
rect 52357 18519 52391 18553
rect 52357 18451 52391 18485
rect 52357 18383 52391 18417
rect 52357 18315 52391 18349
rect 52357 18247 52391 18281
rect 52357 18179 52391 18213
rect 52357 18111 52391 18145
rect 52357 18043 52391 18077
rect 52357 17975 52391 18009
rect 52357 17907 52391 17941
rect 52357 17839 52391 17873
rect 52357 17771 52391 17805
rect 52357 17703 52391 17737
rect 52357 17635 52391 17669
rect 52357 17567 52391 17601
rect 52357 17499 52391 17533
rect 52357 17431 52391 17465
rect 52357 17363 52391 17397
<< psubdiff >>
rect 21744 48003 22360 48042
rect 21744 47901 21831 48003
rect 22273 47901 22360 48003
rect 21744 47862 22360 47901
rect 23858 47229 23898 47272
rect 23858 47195 23861 47229
rect 23895 47195 23898 47229
rect 23858 47152 23898 47195
rect 42986 44861 52314 44896
rect 42986 44838 43116 44861
rect 42986 44804 43020 44838
rect 43054 44827 43116 44838
rect 43150 44827 43206 44861
rect 43240 44827 43296 44861
rect 43330 44827 43386 44861
rect 43420 44827 43476 44861
rect 43510 44827 43566 44861
rect 43600 44827 43656 44861
rect 43690 44827 43746 44861
rect 43780 44827 43836 44861
rect 43870 44827 43926 44861
rect 43960 44827 44016 44861
rect 44050 44827 44106 44861
rect 44140 44838 44456 44861
rect 44140 44827 44207 44838
rect 43054 44804 44207 44827
rect 44241 44804 44360 44838
rect 44394 44827 44456 44838
rect 44490 44827 44546 44861
rect 44580 44827 44636 44861
rect 44670 44827 44726 44861
rect 44760 44827 44816 44861
rect 44850 44827 44906 44861
rect 44940 44827 44996 44861
rect 45030 44827 45086 44861
rect 45120 44827 45176 44861
rect 45210 44827 45266 44861
rect 45300 44827 45356 44861
rect 45390 44827 45446 44861
rect 45480 44838 45796 44861
rect 45480 44827 45547 44838
rect 44394 44804 45547 44827
rect 45581 44804 45700 44838
rect 45734 44827 45796 44838
rect 45830 44827 45886 44861
rect 45920 44827 45976 44861
rect 46010 44827 46066 44861
rect 46100 44827 46156 44861
rect 46190 44827 46246 44861
rect 46280 44827 46336 44861
rect 46370 44827 46426 44861
rect 46460 44827 46516 44861
rect 46550 44827 46606 44861
rect 46640 44827 46696 44861
rect 46730 44827 46786 44861
rect 46820 44838 47136 44861
rect 46820 44827 46887 44838
rect 45734 44804 46887 44827
rect 46921 44804 47040 44838
rect 47074 44827 47136 44838
rect 47170 44827 47226 44861
rect 47260 44827 47316 44861
rect 47350 44827 47406 44861
rect 47440 44827 47496 44861
rect 47530 44827 47586 44861
rect 47620 44827 47676 44861
rect 47710 44827 47766 44861
rect 47800 44827 47856 44861
rect 47890 44827 47946 44861
rect 47980 44827 48036 44861
rect 48070 44827 48126 44861
rect 48160 44838 48476 44861
rect 48160 44827 48227 44838
rect 47074 44804 48227 44827
rect 48261 44804 48380 44838
rect 48414 44827 48476 44838
rect 48510 44827 48566 44861
rect 48600 44827 48656 44861
rect 48690 44827 48746 44861
rect 48780 44827 48836 44861
rect 48870 44827 48926 44861
rect 48960 44827 49016 44861
rect 49050 44827 49106 44861
rect 49140 44827 49196 44861
rect 49230 44827 49286 44861
rect 49320 44827 49376 44861
rect 49410 44827 49466 44861
rect 49500 44838 49816 44861
rect 49500 44827 49567 44838
rect 48414 44804 49567 44827
rect 49601 44804 49720 44838
rect 49754 44827 49816 44838
rect 49850 44827 49906 44861
rect 49940 44827 49996 44861
rect 50030 44827 50086 44861
rect 50120 44827 50176 44861
rect 50210 44827 50266 44861
rect 50300 44827 50356 44861
rect 50390 44827 50446 44861
rect 50480 44827 50536 44861
rect 50570 44827 50626 44861
rect 50660 44827 50716 44861
rect 50750 44827 50806 44861
rect 50840 44838 51156 44861
rect 50840 44827 50907 44838
rect 49754 44804 50907 44827
rect 50941 44804 51060 44838
rect 51094 44827 51156 44838
rect 51190 44827 51246 44861
rect 51280 44827 51336 44861
rect 51370 44827 51426 44861
rect 51460 44827 51516 44861
rect 51550 44827 51606 44861
rect 51640 44827 51696 44861
rect 51730 44827 51786 44861
rect 51820 44827 51876 44861
rect 51910 44827 51966 44861
rect 52000 44827 52056 44861
rect 52090 44827 52146 44861
rect 52180 44838 52314 44861
rect 52180 44827 52247 44838
rect 51094 44804 52247 44827
rect 52281 44804 52314 44838
rect 42986 44795 52314 44804
rect 42986 44748 43087 44795
rect 42986 44714 43020 44748
rect 43054 44714 43087 44748
rect 44173 44748 44427 44795
rect 42986 44658 43087 44714
rect 42986 44624 43020 44658
rect 43054 44624 43087 44658
rect 42986 44568 43087 44624
rect 42986 44534 43020 44568
rect 43054 44534 43087 44568
rect 42986 44478 43087 44534
rect 42986 44444 43020 44478
rect 43054 44444 43087 44478
rect 42986 44388 43087 44444
rect 42986 44354 43020 44388
rect 43054 44354 43087 44388
rect 42986 44298 43087 44354
rect 42986 44264 43020 44298
rect 43054 44264 43087 44298
rect 42986 44208 43087 44264
rect 42986 44174 43020 44208
rect 43054 44174 43087 44208
rect 42986 44118 43087 44174
rect 42986 44084 43020 44118
rect 43054 44084 43087 44118
rect 42986 44028 43087 44084
rect 42986 43994 43020 44028
rect 43054 43994 43087 44028
rect 42986 43938 43087 43994
rect 42986 43904 43020 43938
rect 43054 43904 43087 43938
rect 42986 43848 43087 43904
rect 42986 43814 43020 43848
rect 43054 43814 43087 43848
rect 42986 43758 43087 43814
rect 44173 44714 44207 44748
rect 44241 44714 44360 44748
rect 44394 44714 44427 44748
rect 45513 44748 45767 44795
rect 44173 44658 44427 44714
rect 44173 44624 44207 44658
rect 44241 44624 44360 44658
rect 44394 44624 44427 44658
rect 44173 44568 44427 44624
rect 44173 44534 44207 44568
rect 44241 44534 44360 44568
rect 44394 44534 44427 44568
rect 44173 44478 44427 44534
rect 44173 44444 44207 44478
rect 44241 44444 44360 44478
rect 44394 44444 44427 44478
rect 44173 44388 44427 44444
rect 44173 44354 44207 44388
rect 44241 44354 44360 44388
rect 44394 44354 44427 44388
rect 44173 44298 44427 44354
rect 44173 44264 44207 44298
rect 44241 44264 44360 44298
rect 44394 44264 44427 44298
rect 44173 44208 44427 44264
rect 44173 44174 44207 44208
rect 44241 44174 44360 44208
rect 44394 44174 44427 44208
rect 44173 44118 44427 44174
rect 44173 44084 44207 44118
rect 44241 44084 44360 44118
rect 44394 44084 44427 44118
rect 44173 44028 44427 44084
rect 44173 43994 44207 44028
rect 44241 43994 44360 44028
rect 44394 43994 44427 44028
rect 44173 43938 44427 43994
rect 44173 43904 44207 43938
rect 44241 43904 44360 43938
rect 44394 43904 44427 43938
rect 44173 43848 44427 43904
rect 44173 43814 44207 43848
rect 44241 43814 44360 43848
rect 44394 43814 44427 43848
rect 42986 43724 43020 43758
rect 43054 43724 43087 43758
rect 42986 43709 43087 43724
rect 44173 43758 44427 43814
rect 45513 44714 45547 44748
rect 45581 44714 45700 44748
rect 45734 44714 45767 44748
rect 46853 44748 47107 44795
rect 45513 44658 45767 44714
rect 45513 44624 45547 44658
rect 45581 44624 45700 44658
rect 45734 44624 45767 44658
rect 45513 44568 45767 44624
rect 45513 44534 45547 44568
rect 45581 44534 45700 44568
rect 45734 44534 45767 44568
rect 45513 44478 45767 44534
rect 45513 44444 45547 44478
rect 45581 44444 45700 44478
rect 45734 44444 45767 44478
rect 45513 44388 45767 44444
rect 45513 44354 45547 44388
rect 45581 44354 45700 44388
rect 45734 44354 45767 44388
rect 45513 44298 45767 44354
rect 45513 44264 45547 44298
rect 45581 44264 45700 44298
rect 45734 44264 45767 44298
rect 45513 44208 45767 44264
rect 45513 44174 45547 44208
rect 45581 44174 45700 44208
rect 45734 44174 45767 44208
rect 45513 44118 45767 44174
rect 45513 44084 45547 44118
rect 45581 44084 45700 44118
rect 45734 44084 45767 44118
rect 45513 44028 45767 44084
rect 45513 43994 45547 44028
rect 45581 43994 45700 44028
rect 45734 43994 45767 44028
rect 45513 43938 45767 43994
rect 45513 43904 45547 43938
rect 45581 43904 45700 43938
rect 45734 43904 45767 43938
rect 45513 43848 45767 43904
rect 45513 43814 45547 43848
rect 45581 43814 45700 43848
rect 45734 43814 45767 43848
rect 44173 43724 44207 43758
rect 44241 43724 44360 43758
rect 44394 43724 44427 43758
rect 44173 43709 44427 43724
rect 45513 43758 45767 43814
rect 46853 44714 46887 44748
rect 46921 44714 47040 44748
rect 47074 44714 47107 44748
rect 48193 44748 48447 44795
rect 46853 44658 47107 44714
rect 46853 44624 46887 44658
rect 46921 44624 47040 44658
rect 47074 44624 47107 44658
rect 46853 44568 47107 44624
rect 46853 44534 46887 44568
rect 46921 44534 47040 44568
rect 47074 44534 47107 44568
rect 46853 44478 47107 44534
rect 46853 44444 46887 44478
rect 46921 44444 47040 44478
rect 47074 44444 47107 44478
rect 46853 44388 47107 44444
rect 46853 44354 46887 44388
rect 46921 44354 47040 44388
rect 47074 44354 47107 44388
rect 46853 44298 47107 44354
rect 46853 44264 46887 44298
rect 46921 44264 47040 44298
rect 47074 44264 47107 44298
rect 46853 44208 47107 44264
rect 46853 44174 46887 44208
rect 46921 44174 47040 44208
rect 47074 44174 47107 44208
rect 46853 44118 47107 44174
rect 46853 44084 46887 44118
rect 46921 44084 47040 44118
rect 47074 44084 47107 44118
rect 46853 44028 47107 44084
rect 46853 43994 46887 44028
rect 46921 43994 47040 44028
rect 47074 43994 47107 44028
rect 46853 43938 47107 43994
rect 46853 43904 46887 43938
rect 46921 43904 47040 43938
rect 47074 43904 47107 43938
rect 46853 43848 47107 43904
rect 46853 43814 46887 43848
rect 46921 43814 47040 43848
rect 47074 43814 47107 43848
rect 45513 43724 45547 43758
rect 45581 43724 45700 43758
rect 45734 43724 45767 43758
rect 45513 43709 45767 43724
rect 46853 43758 47107 43814
rect 48193 44714 48227 44748
rect 48261 44714 48380 44748
rect 48414 44714 48447 44748
rect 49533 44748 49787 44795
rect 48193 44658 48447 44714
rect 48193 44624 48227 44658
rect 48261 44624 48380 44658
rect 48414 44624 48447 44658
rect 48193 44568 48447 44624
rect 48193 44534 48227 44568
rect 48261 44534 48380 44568
rect 48414 44534 48447 44568
rect 48193 44478 48447 44534
rect 48193 44444 48227 44478
rect 48261 44444 48380 44478
rect 48414 44444 48447 44478
rect 48193 44388 48447 44444
rect 48193 44354 48227 44388
rect 48261 44354 48380 44388
rect 48414 44354 48447 44388
rect 48193 44298 48447 44354
rect 48193 44264 48227 44298
rect 48261 44264 48380 44298
rect 48414 44264 48447 44298
rect 48193 44208 48447 44264
rect 48193 44174 48227 44208
rect 48261 44174 48380 44208
rect 48414 44174 48447 44208
rect 48193 44118 48447 44174
rect 48193 44084 48227 44118
rect 48261 44084 48380 44118
rect 48414 44084 48447 44118
rect 48193 44028 48447 44084
rect 48193 43994 48227 44028
rect 48261 43994 48380 44028
rect 48414 43994 48447 44028
rect 48193 43938 48447 43994
rect 48193 43904 48227 43938
rect 48261 43904 48380 43938
rect 48414 43904 48447 43938
rect 48193 43848 48447 43904
rect 48193 43814 48227 43848
rect 48261 43814 48380 43848
rect 48414 43814 48447 43848
rect 46853 43724 46887 43758
rect 46921 43724 47040 43758
rect 47074 43724 47107 43758
rect 46853 43709 47107 43724
rect 48193 43758 48447 43814
rect 49533 44714 49567 44748
rect 49601 44714 49720 44748
rect 49754 44714 49787 44748
rect 50873 44748 51127 44795
rect 49533 44658 49787 44714
rect 49533 44624 49567 44658
rect 49601 44624 49720 44658
rect 49754 44624 49787 44658
rect 49533 44568 49787 44624
rect 49533 44534 49567 44568
rect 49601 44534 49720 44568
rect 49754 44534 49787 44568
rect 49533 44478 49787 44534
rect 49533 44444 49567 44478
rect 49601 44444 49720 44478
rect 49754 44444 49787 44478
rect 49533 44388 49787 44444
rect 49533 44354 49567 44388
rect 49601 44354 49720 44388
rect 49754 44354 49787 44388
rect 49533 44298 49787 44354
rect 49533 44264 49567 44298
rect 49601 44264 49720 44298
rect 49754 44264 49787 44298
rect 49533 44208 49787 44264
rect 49533 44174 49567 44208
rect 49601 44174 49720 44208
rect 49754 44174 49787 44208
rect 49533 44118 49787 44174
rect 49533 44084 49567 44118
rect 49601 44084 49720 44118
rect 49754 44084 49787 44118
rect 49533 44028 49787 44084
rect 49533 43994 49567 44028
rect 49601 43994 49720 44028
rect 49754 43994 49787 44028
rect 49533 43938 49787 43994
rect 49533 43904 49567 43938
rect 49601 43904 49720 43938
rect 49754 43904 49787 43938
rect 49533 43848 49787 43904
rect 49533 43814 49567 43848
rect 49601 43814 49720 43848
rect 49754 43814 49787 43848
rect 48193 43724 48227 43758
rect 48261 43724 48380 43758
rect 48414 43724 48447 43758
rect 48193 43709 48447 43724
rect 49533 43758 49787 43814
rect 50873 44714 50907 44748
rect 50941 44714 51060 44748
rect 51094 44714 51127 44748
rect 52213 44748 52314 44795
rect 50873 44658 51127 44714
rect 50873 44624 50907 44658
rect 50941 44624 51060 44658
rect 51094 44624 51127 44658
rect 50873 44568 51127 44624
rect 50873 44534 50907 44568
rect 50941 44534 51060 44568
rect 51094 44534 51127 44568
rect 50873 44478 51127 44534
rect 50873 44444 50907 44478
rect 50941 44444 51060 44478
rect 51094 44444 51127 44478
rect 50873 44388 51127 44444
rect 50873 44354 50907 44388
rect 50941 44354 51060 44388
rect 51094 44354 51127 44388
rect 50873 44298 51127 44354
rect 50873 44264 50907 44298
rect 50941 44264 51060 44298
rect 51094 44264 51127 44298
rect 50873 44208 51127 44264
rect 50873 44174 50907 44208
rect 50941 44174 51060 44208
rect 51094 44174 51127 44208
rect 50873 44118 51127 44174
rect 50873 44084 50907 44118
rect 50941 44084 51060 44118
rect 51094 44084 51127 44118
rect 50873 44028 51127 44084
rect 50873 43994 50907 44028
rect 50941 43994 51060 44028
rect 51094 43994 51127 44028
rect 50873 43938 51127 43994
rect 50873 43904 50907 43938
rect 50941 43904 51060 43938
rect 51094 43904 51127 43938
rect 50873 43848 51127 43904
rect 50873 43814 50907 43848
rect 50941 43814 51060 43848
rect 51094 43814 51127 43848
rect 49533 43724 49567 43758
rect 49601 43724 49720 43758
rect 49754 43724 49787 43758
rect 49533 43709 49787 43724
rect 50873 43758 51127 43814
rect 52213 44714 52247 44748
rect 52281 44714 52314 44748
rect 52213 44658 52314 44714
rect 52213 44624 52247 44658
rect 52281 44624 52314 44658
rect 52213 44568 52314 44624
rect 52213 44534 52247 44568
rect 52281 44534 52314 44568
rect 52213 44478 52314 44534
rect 52213 44444 52247 44478
rect 52281 44444 52314 44478
rect 52213 44388 52314 44444
rect 52213 44354 52247 44388
rect 52281 44354 52314 44388
rect 52213 44298 52314 44354
rect 52213 44264 52247 44298
rect 52281 44264 52314 44298
rect 52213 44208 52314 44264
rect 52213 44174 52247 44208
rect 52281 44174 52314 44208
rect 52213 44118 52314 44174
rect 52213 44084 52247 44118
rect 52281 44084 52314 44118
rect 52213 44028 52314 44084
rect 52213 43994 52247 44028
rect 52281 43994 52314 44028
rect 52213 43938 52314 43994
rect 52213 43904 52247 43938
rect 52281 43904 52314 43938
rect 52213 43848 52314 43904
rect 52213 43814 52247 43848
rect 52281 43814 52314 43848
rect 50873 43724 50907 43758
rect 50941 43724 51060 43758
rect 51094 43724 51127 43758
rect 50873 43709 51127 43724
rect 52213 43758 52314 43814
rect 52213 43724 52247 43758
rect 52281 43724 52314 43758
rect 52213 43709 52314 43724
rect 42986 43674 52314 43709
rect 14058 43469 14098 43512
rect 14058 43435 14061 43469
rect 14095 43435 14098 43469
rect 42986 43640 43116 43674
rect 43150 43640 43206 43674
rect 43240 43640 43296 43674
rect 43330 43640 43386 43674
rect 43420 43640 43476 43674
rect 43510 43640 43566 43674
rect 43600 43640 43656 43674
rect 43690 43640 43746 43674
rect 43780 43640 43836 43674
rect 43870 43640 43926 43674
rect 43960 43640 44016 43674
rect 44050 43640 44106 43674
rect 44140 43640 44456 43674
rect 44490 43640 44546 43674
rect 44580 43640 44636 43674
rect 44670 43640 44726 43674
rect 44760 43640 44816 43674
rect 44850 43640 44906 43674
rect 44940 43640 44996 43674
rect 45030 43640 45086 43674
rect 45120 43640 45176 43674
rect 45210 43640 45266 43674
rect 45300 43640 45356 43674
rect 45390 43640 45446 43674
rect 45480 43640 45796 43674
rect 45830 43640 45886 43674
rect 45920 43640 45976 43674
rect 46010 43640 46066 43674
rect 46100 43640 46156 43674
rect 46190 43640 46246 43674
rect 46280 43640 46336 43674
rect 46370 43640 46426 43674
rect 46460 43640 46516 43674
rect 46550 43640 46606 43674
rect 46640 43640 46696 43674
rect 46730 43640 46786 43674
rect 46820 43640 47136 43674
rect 47170 43640 47226 43674
rect 47260 43640 47316 43674
rect 47350 43640 47406 43674
rect 47440 43640 47496 43674
rect 47530 43640 47586 43674
rect 47620 43640 47676 43674
rect 47710 43640 47766 43674
rect 47800 43640 47856 43674
rect 47890 43640 47946 43674
rect 47980 43640 48036 43674
rect 48070 43640 48126 43674
rect 48160 43640 48476 43674
rect 48510 43640 48566 43674
rect 48600 43640 48656 43674
rect 48690 43640 48746 43674
rect 48780 43640 48836 43674
rect 48870 43640 48926 43674
rect 48960 43640 49016 43674
rect 49050 43640 49106 43674
rect 49140 43640 49196 43674
rect 49230 43640 49286 43674
rect 49320 43640 49376 43674
rect 49410 43640 49466 43674
rect 49500 43640 49816 43674
rect 49850 43640 49906 43674
rect 49940 43640 49996 43674
rect 50030 43640 50086 43674
rect 50120 43640 50176 43674
rect 50210 43640 50266 43674
rect 50300 43640 50356 43674
rect 50390 43640 50446 43674
rect 50480 43640 50536 43674
rect 50570 43640 50626 43674
rect 50660 43640 50716 43674
rect 50750 43640 50806 43674
rect 50840 43640 51156 43674
rect 51190 43640 51246 43674
rect 51280 43640 51336 43674
rect 51370 43640 51426 43674
rect 51460 43640 51516 43674
rect 51550 43640 51606 43674
rect 51640 43640 51696 43674
rect 51730 43640 51786 43674
rect 51820 43640 51876 43674
rect 51910 43640 51966 43674
rect 52000 43640 52056 43674
rect 52090 43640 52146 43674
rect 52180 43640 52314 43674
rect 42986 43608 52314 43640
rect 14058 43392 14098 43435
rect 41810 41101 52478 41136
rect 41810 41078 41940 41101
rect 41810 41044 41844 41078
rect 41878 41067 41940 41078
rect 41974 41067 42030 41101
rect 42064 41067 42120 41101
rect 42154 41067 42210 41101
rect 42244 41067 42300 41101
rect 42334 41067 42390 41101
rect 42424 41067 42480 41101
rect 42514 41067 42570 41101
rect 42604 41067 42660 41101
rect 42694 41067 42750 41101
rect 42784 41067 42840 41101
rect 42874 41067 42930 41101
rect 42964 41078 43280 41101
rect 42964 41067 43031 41078
rect 41878 41044 43031 41067
rect 43065 41044 43184 41078
rect 43218 41067 43280 41078
rect 43314 41067 43370 41101
rect 43404 41067 43460 41101
rect 43494 41067 43550 41101
rect 43584 41067 43640 41101
rect 43674 41067 43730 41101
rect 43764 41067 43820 41101
rect 43854 41067 43910 41101
rect 43944 41067 44000 41101
rect 44034 41067 44090 41101
rect 44124 41067 44180 41101
rect 44214 41067 44270 41101
rect 44304 41078 44620 41101
rect 44304 41067 44371 41078
rect 43218 41044 44371 41067
rect 44405 41044 44524 41078
rect 44558 41067 44620 41078
rect 44654 41067 44710 41101
rect 44744 41067 44800 41101
rect 44834 41067 44890 41101
rect 44924 41067 44980 41101
rect 45014 41067 45070 41101
rect 45104 41067 45160 41101
rect 45194 41067 45250 41101
rect 45284 41067 45340 41101
rect 45374 41067 45430 41101
rect 45464 41067 45520 41101
rect 45554 41067 45610 41101
rect 45644 41078 45960 41101
rect 45644 41067 45711 41078
rect 44558 41044 45711 41067
rect 45745 41044 45864 41078
rect 45898 41067 45960 41078
rect 45994 41067 46050 41101
rect 46084 41067 46140 41101
rect 46174 41067 46230 41101
rect 46264 41067 46320 41101
rect 46354 41067 46410 41101
rect 46444 41067 46500 41101
rect 46534 41067 46590 41101
rect 46624 41067 46680 41101
rect 46714 41067 46770 41101
rect 46804 41067 46860 41101
rect 46894 41067 46950 41101
rect 46984 41078 47300 41101
rect 46984 41067 47051 41078
rect 45898 41044 47051 41067
rect 47085 41044 47204 41078
rect 47238 41067 47300 41078
rect 47334 41067 47390 41101
rect 47424 41067 47480 41101
rect 47514 41067 47570 41101
rect 47604 41067 47660 41101
rect 47694 41067 47750 41101
rect 47784 41067 47840 41101
rect 47874 41067 47930 41101
rect 47964 41067 48020 41101
rect 48054 41067 48110 41101
rect 48144 41067 48200 41101
rect 48234 41067 48290 41101
rect 48324 41078 48640 41101
rect 48324 41067 48391 41078
rect 47238 41044 48391 41067
rect 48425 41044 48544 41078
rect 48578 41067 48640 41078
rect 48674 41067 48730 41101
rect 48764 41067 48820 41101
rect 48854 41067 48910 41101
rect 48944 41067 49000 41101
rect 49034 41067 49090 41101
rect 49124 41067 49180 41101
rect 49214 41067 49270 41101
rect 49304 41067 49360 41101
rect 49394 41067 49450 41101
rect 49484 41067 49540 41101
rect 49574 41067 49630 41101
rect 49664 41078 49980 41101
rect 49664 41067 49731 41078
rect 48578 41044 49731 41067
rect 49765 41044 49884 41078
rect 49918 41067 49980 41078
rect 50014 41067 50070 41101
rect 50104 41067 50160 41101
rect 50194 41067 50250 41101
rect 50284 41067 50340 41101
rect 50374 41067 50430 41101
rect 50464 41067 50520 41101
rect 50554 41067 50610 41101
rect 50644 41067 50700 41101
rect 50734 41067 50790 41101
rect 50824 41067 50880 41101
rect 50914 41067 50970 41101
rect 51004 41078 51320 41101
rect 51004 41067 51071 41078
rect 49918 41044 51071 41067
rect 51105 41044 51224 41078
rect 51258 41067 51320 41078
rect 51354 41067 51410 41101
rect 51444 41067 51500 41101
rect 51534 41067 51590 41101
rect 51624 41067 51680 41101
rect 51714 41067 51770 41101
rect 51804 41067 51860 41101
rect 51894 41067 51950 41101
rect 51984 41067 52040 41101
rect 52074 41067 52130 41101
rect 52164 41067 52220 41101
rect 52254 41067 52310 41101
rect 52344 41078 52478 41101
rect 52344 41067 52411 41078
rect 51258 41044 52411 41067
rect 52445 41044 52478 41078
rect 41810 41035 52478 41044
rect 41810 40988 41911 41035
rect 41810 40954 41844 40988
rect 41878 40954 41911 40988
rect 42997 40988 43251 41035
rect 41810 40898 41911 40954
rect 41810 40864 41844 40898
rect 41878 40864 41911 40898
rect 41810 40808 41911 40864
rect 41810 40774 41844 40808
rect 41878 40774 41911 40808
rect 41810 40718 41911 40774
rect 41810 40684 41844 40718
rect 41878 40684 41911 40718
rect 41810 40628 41911 40684
rect 41810 40594 41844 40628
rect 41878 40594 41911 40628
rect 41810 40538 41911 40594
rect 41810 40504 41844 40538
rect 41878 40504 41911 40538
rect 41810 40448 41911 40504
rect 41810 40414 41844 40448
rect 41878 40414 41911 40448
rect 41810 40358 41911 40414
rect 41810 40324 41844 40358
rect 41878 40324 41911 40358
rect 41810 40268 41911 40324
rect 41810 40234 41844 40268
rect 41878 40234 41911 40268
rect 41810 40178 41911 40234
rect 41810 40144 41844 40178
rect 41878 40144 41911 40178
rect 41810 40088 41911 40144
rect 41810 40054 41844 40088
rect 41878 40054 41911 40088
rect 41810 39998 41911 40054
rect 42997 40954 43031 40988
rect 43065 40954 43184 40988
rect 43218 40954 43251 40988
rect 44337 40988 44591 41035
rect 42997 40898 43251 40954
rect 42997 40864 43031 40898
rect 43065 40864 43184 40898
rect 43218 40864 43251 40898
rect 42997 40808 43251 40864
rect 42997 40774 43031 40808
rect 43065 40774 43184 40808
rect 43218 40774 43251 40808
rect 42997 40718 43251 40774
rect 42997 40684 43031 40718
rect 43065 40684 43184 40718
rect 43218 40684 43251 40718
rect 42997 40628 43251 40684
rect 42997 40594 43031 40628
rect 43065 40594 43184 40628
rect 43218 40594 43251 40628
rect 42997 40538 43251 40594
rect 42997 40504 43031 40538
rect 43065 40504 43184 40538
rect 43218 40504 43251 40538
rect 42997 40448 43251 40504
rect 42997 40414 43031 40448
rect 43065 40414 43184 40448
rect 43218 40414 43251 40448
rect 42997 40358 43251 40414
rect 42997 40324 43031 40358
rect 43065 40324 43184 40358
rect 43218 40324 43251 40358
rect 42997 40268 43251 40324
rect 42997 40234 43031 40268
rect 43065 40234 43184 40268
rect 43218 40234 43251 40268
rect 42997 40178 43251 40234
rect 42997 40144 43031 40178
rect 43065 40144 43184 40178
rect 43218 40144 43251 40178
rect 42997 40088 43251 40144
rect 42997 40054 43031 40088
rect 43065 40054 43184 40088
rect 43218 40054 43251 40088
rect 41810 39964 41844 39998
rect 41878 39964 41911 39998
rect 41810 39949 41911 39964
rect 42997 39998 43251 40054
rect 44337 40954 44371 40988
rect 44405 40954 44524 40988
rect 44558 40954 44591 40988
rect 45677 40988 45931 41035
rect 44337 40898 44591 40954
rect 44337 40864 44371 40898
rect 44405 40864 44524 40898
rect 44558 40864 44591 40898
rect 44337 40808 44591 40864
rect 44337 40774 44371 40808
rect 44405 40774 44524 40808
rect 44558 40774 44591 40808
rect 44337 40718 44591 40774
rect 44337 40684 44371 40718
rect 44405 40684 44524 40718
rect 44558 40684 44591 40718
rect 44337 40628 44591 40684
rect 44337 40594 44371 40628
rect 44405 40594 44524 40628
rect 44558 40594 44591 40628
rect 44337 40538 44591 40594
rect 44337 40504 44371 40538
rect 44405 40504 44524 40538
rect 44558 40504 44591 40538
rect 44337 40448 44591 40504
rect 44337 40414 44371 40448
rect 44405 40414 44524 40448
rect 44558 40414 44591 40448
rect 44337 40358 44591 40414
rect 44337 40324 44371 40358
rect 44405 40324 44524 40358
rect 44558 40324 44591 40358
rect 44337 40268 44591 40324
rect 44337 40234 44371 40268
rect 44405 40234 44524 40268
rect 44558 40234 44591 40268
rect 44337 40178 44591 40234
rect 44337 40144 44371 40178
rect 44405 40144 44524 40178
rect 44558 40144 44591 40178
rect 44337 40088 44591 40144
rect 44337 40054 44371 40088
rect 44405 40054 44524 40088
rect 44558 40054 44591 40088
rect 42997 39964 43031 39998
rect 43065 39964 43184 39998
rect 43218 39964 43251 39998
rect 42997 39949 43251 39964
rect 44337 39998 44591 40054
rect 45677 40954 45711 40988
rect 45745 40954 45864 40988
rect 45898 40954 45931 40988
rect 47017 40988 47271 41035
rect 45677 40898 45931 40954
rect 45677 40864 45711 40898
rect 45745 40864 45864 40898
rect 45898 40864 45931 40898
rect 45677 40808 45931 40864
rect 45677 40774 45711 40808
rect 45745 40774 45864 40808
rect 45898 40774 45931 40808
rect 45677 40718 45931 40774
rect 45677 40684 45711 40718
rect 45745 40684 45864 40718
rect 45898 40684 45931 40718
rect 45677 40628 45931 40684
rect 45677 40594 45711 40628
rect 45745 40594 45864 40628
rect 45898 40594 45931 40628
rect 45677 40538 45931 40594
rect 45677 40504 45711 40538
rect 45745 40504 45864 40538
rect 45898 40504 45931 40538
rect 45677 40448 45931 40504
rect 45677 40414 45711 40448
rect 45745 40414 45864 40448
rect 45898 40414 45931 40448
rect 45677 40358 45931 40414
rect 45677 40324 45711 40358
rect 45745 40324 45864 40358
rect 45898 40324 45931 40358
rect 45677 40268 45931 40324
rect 45677 40234 45711 40268
rect 45745 40234 45864 40268
rect 45898 40234 45931 40268
rect 45677 40178 45931 40234
rect 45677 40144 45711 40178
rect 45745 40144 45864 40178
rect 45898 40144 45931 40178
rect 45677 40088 45931 40144
rect 45677 40054 45711 40088
rect 45745 40054 45864 40088
rect 45898 40054 45931 40088
rect 44337 39964 44371 39998
rect 44405 39964 44524 39998
rect 44558 39964 44591 39998
rect 44337 39949 44591 39964
rect 45677 39998 45931 40054
rect 47017 40954 47051 40988
rect 47085 40954 47204 40988
rect 47238 40954 47271 40988
rect 48357 40988 48611 41035
rect 47017 40898 47271 40954
rect 47017 40864 47051 40898
rect 47085 40864 47204 40898
rect 47238 40864 47271 40898
rect 47017 40808 47271 40864
rect 47017 40774 47051 40808
rect 47085 40774 47204 40808
rect 47238 40774 47271 40808
rect 47017 40718 47271 40774
rect 47017 40684 47051 40718
rect 47085 40684 47204 40718
rect 47238 40684 47271 40718
rect 47017 40628 47271 40684
rect 47017 40594 47051 40628
rect 47085 40594 47204 40628
rect 47238 40594 47271 40628
rect 47017 40538 47271 40594
rect 47017 40504 47051 40538
rect 47085 40504 47204 40538
rect 47238 40504 47271 40538
rect 47017 40448 47271 40504
rect 47017 40414 47051 40448
rect 47085 40414 47204 40448
rect 47238 40414 47271 40448
rect 47017 40358 47271 40414
rect 47017 40324 47051 40358
rect 47085 40324 47204 40358
rect 47238 40324 47271 40358
rect 47017 40268 47271 40324
rect 47017 40234 47051 40268
rect 47085 40234 47204 40268
rect 47238 40234 47271 40268
rect 47017 40178 47271 40234
rect 47017 40144 47051 40178
rect 47085 40144 47204 40178
rect 47238 40144 47271 40178
rect 47017 40088 47271 40144
rect 47017 40054 47051 40088
rect 47085 40054 47204 40088
rect 47238 40054 47271 40088
rect 45677 39964 45711 39998
rect 45745 39964 45864 39998
rect 45898 39964 45931 39998
rect 45677 39949 45931 39964
rect 47017 39998 47271 40054
rect 48357 40954 48391 40988
rect 48425 40954 48544 40988
rect 48578 40954 48611 40988
rect 49697 40988 49951 41035
rect 48357 40898 48611 40954
rect 48357 40864 48391 40898
rect 48425 40864 48544 40898
rect 48578 40864 48611 40898
rect 48357 40808 48611 40864
rect 48357 40774 48391 40808
rect 48425 40774 48544 40808
rect 48578 40774 48611 40808
rect 48357 40718 48611 40774
rect 48357 40684 48391 40718
rect 48425 40684 48544 40718
rect 48578 40684 48611 40718
rect 48357 40628 48611 40684
rect 48357 40594 48391 40628
rect 48425 40594 48544 40628
rect 48578 40594 48611 40628
rect 48357 40538 48611 40594
rect 48357 40504 48391 40538
rect 48425 40504 48544 40538
rect 48578 40504 48611 40538
rect 48357 40448 48611 40504
rect 48357 40414 48391 40448
rect 48425 40414 48544 40448
rect 48578 40414 48611 40448
rect 48357 40358 48611 40414
rect 48357 40324 48391 40358
rect 48425 40324 48544 40358
rect 48578 40324 48611 40358
rect 48357 40268 48611 40324
rect 48357 40234 48391 40268
rect 48425 40234 48544 40268
rect 48578 40234 48611 40268
rect 48357 40178 48611 40234
rect 48357 40144 48391 40178
rect 48425 40144 48544 40178
rect 48578 40144 48611 40178
rect 48357 40088 48611 40144
rect 48357 40054 48391 40088
rect 48425 40054 48544 40088
rect 48578 40054 48611 40088
rect 47017 39964 47051 39998
rect 47085 39964 47204 39998
rect 47238 39964 47271 39998
rect 47017 39949 47271 39964
rect 48357 39998 48611 40054
rect 49697 40954 49731 40988
rect 49765 40954 49884 40988
rect 49918 40954 49951 40988
rect 51037 40988 51291 41035
rect 49697 40898 49951 40954
rect 49697 40864 49731 40898
rect 49765 40864 49884 40898
rect 49918 40864 49951 40898
rect 49697 40808 49951 40864
rect 49697 40774 49731 40808
rect 49765 40774 49884 40808
rect 49918 40774 49951 40808
rect 49697 40718 49951 40774
rect 49697 40684 49731 40718
rect 49765 40684 49884 40718
rect 49918 40684 49951 40718
rect 49697 40628 49951 40684
rect 49697 40594 49731 40628
rect 49765 40594 49884 40628
rect 49918 40594 49951 40628
rect 49697 40538 49951 40594
rect 49697 40504 49731 40538
rect 49765 40504 49884 40538
rect 49918 40504 49951 40538
rect 49697 40448 49951 40504
rect 49697 40414 49731 40448
rect 49765 40414 49884 40448
rect 49918 40414 49951 40448
rect 49697 40358 49951 40414
rect 49697 40324 49731 40358
rect 49765 40324 49884 40358
rect 49918 40324 49951 40358
rect 49697 40268 49951 40324
rect 49697 40234 49731 40268
rect 49765 40234 49884 40268
rect 49918 40234 49951 40268
rect 49697 40178 49951 40234
rect 49697 40144 49731 40178
rect 49765 40144 49884 40178
rect 49918 40144 49951 40178
rect 49697 40088 49951 40144
rect 49697 40054 49731 40088
rect 49765 40054 49884 40088
rect 49918 40054 49951 40088
rect 48357 39964 48391 39998
rect 48425 39964 48544 39998
rect 48578 39964 48611 39998
rect 48357 39949 48611 39964
rect 49697 39998 49951 40054
rect 51037 40954 51071 40988
rect 51105 40954 51224 40988
rect 51258 40954 51291 40988
rect 52377 40988 52478 41035
rect 51037 40898 51291 40954
rect 51037 40864 51071 40898
rect 51105 40864 51224 40898
rect 51258 40864 51291 40898
rect 51037 40808 51291 40864
rect 51037 40774 51071 40808
rect 51105 40774 51224 40808
rect 51258 40774 51291 40808
rect 51037 40718 51291 40774
rect 51037 40684 51071 40718
rect 51105 40684 51224 40718
rect 51258 40684 51291 40718
rect 51037 40628 51291 40684
rect 51037 40594 51071 40628
rect 51105 40594 51224 40628
rect 51258 40594 51291 40628
rect 51037 40538 51291 40594
rect 51037 40504 51071 40538
rect 51105 40504 51224 40538
rect 51258 40504 51291 40538
rect 51037 40448 51291 40504
rect 51037 40414 51071 40448
rect 51105 40414 51224 40448
rect 51258 40414 51291 40448
rect 51037 40358 51291 40414
rect 51037 40324 51071 40358
rect 51105 40324 51224 40358
rect 51258 40324 51291 40358
rect 51037 40268 51291 40324
rect 51037 40234 51071 40268
rect 51105 40234 51224 40268
rect 51258 40234 51291 40268
rect 51037 40178 51291 40234
rect 51037 40144 51071 40178
rect 51105 40144 51224 40178
rect 51258 40144 51291 40178
rect 51037 40088 51291 40144
rect 51037 40054 51071 40088
rect 51105 40054 51224 40088
rect 51258 40054 51291 40088
rect 49697 39964 49731 39998
rect 49765 39964 49884 39998
rect 49918 39964 49951 39998
rect 49697 39949 49951 39964
rect 51037 39998 51291 40054
rect 52377 40954 52411 40988
rect 52445 40954 52478 40988
rect 52377 40898 52478 40954
rect 52377 40864 52411 40898
rect 52445 40864 52478 40898
rect 52377 40808 52478 40864
rect 52377 40774 52411 40808
rect 52445 40774 52478 40808
rect 52377 40718 52478 40774
rect 52377 40684 52411 40718
rect 52445 40684 52478 40718
rect 52377 40628 52478 40684
rect 52377 40594 52411 40628
rect 52445 40594 52478 40628
rect 52377 40538 52478 40594
rect 52377 40504 52411 40538
rect 52445 40504 52478 40538
rect 52377 40448 52478 40504
rect 52377 40414 52411 40448
rect 52445 40414 52478 40448
rect 52377 40358 52478 40414
rect 52377 40324 52411 40358
rect 52445 40324 52478 40358
rect 52377 40268 52478 40324
rect 52377 40234 52411 40268
rect 52445 40234 52478 40268
rect 52377 40178 52478 40234
rect 52377 40144 52411 40178
rect 52445 40144 52478 40178
rect 52377 40088 52478 40144
rect 52377 40054 52411 40088
rect 52445 40054 52478 40088
rect 51037 39964 51071 39998
rect 51105 39964 51224 39998
rect 51258 39964 51291 39998
rect 51037 39949 51291 39964
rect 52377 39998 52478 40054
rect 52377 39964 52411 39998
rect 52445 39964 52478 39998
rect 52377 39949 52478 39964
rect 41810 39914 52478 39949
rect 41810 39880 41940 39914
rect 41974 39880 42030 39914
rect 42064 39880 42120 39914
rect 42154 39880 42210 39914
rect 42244 39880 42300 39914
rect 42334 39880 42390 39914
rect 42424 39880 42480 39914
rect 42514 39880 42570 39914
rect 42604 39880 42660 39914
rect 42694 39880 42750 39914
rect 42784 39880 42840 39914
rect 42874 39880 42930 39914
rect 42964 39880 43280 39914
rect 43314 39880 43370 39914
rect 43404 39880 43460 39914
rect 43494 39880 43550 39914
rect 43584 39880 43640 39914
rect 43674 39880 43730 39914
rect 43764 39880 43820 39914
rect 43854 39880 43910 39914
rect 43944 39880 44000 39914
rect 44034 39880 44090 39914
rect 44124 39880 44180 39914
rect 44214 39880 44270 39914
rect 44304 39880 44620 39914
rect 44654 39880 44710 39914
rect 44744 39880 44800 39914
rect 44834 39880 44890 39914
rect 44924 39880 44980 39914
rect 45014 39880 45070 39914
rect 45104 39880 45160 39914
rect 45194 39880 45250 39914
rect 45284 39880 45340 39914
rect 45374 39880 45430 39914
rect 45464 39880 45520 39914
rect 45554 39880 45610 39914
rect 45644 39880 45960 39914
rect 45994 39880 46050 39914
rect 46084 39880 46140 39914
rect 46174 39880 46230 39914
rect 46264 39880 46320 39914
rect 46354 39880 46410 39914
rect 46444 39880 46500 39914
rect 46534 39880 46590 39914
rect 46624 39880 46680 39914
rect 46714 39880 46770 39914
rect 46804 39880 46860 39914
rect 46894 39880 46950 39914
rect 46984 39880 47300 39914
rect 47334 39880 47390 39914
rect 47424 39880 47480 39914
rect 47514 39880 47570 39914
rect 47604 39880 47660 39914
rect 47694 39880 47750 39914
rect 47784 39880 47840 39914
rect 47874 39880 47930 39914
rect 47964 39880 48020 39914
rect 48054 39880 48110 39914
rect 48144 39880 48200 39914
rect 48234 39880 48290 39914
rect 48324 39880 48640 39914
rect 48674 39880 48730 39914
rect 48764 39880 48820 39914
rect 48854 39880 48910 39914
rect 48944 39880 49000 39914
rect 49034 39880 49090 39914
rect 49124 39880 49180 39914
rect 49214 39880 49270 39914
rect 49304 39880 49360 39914
rect 49394 39880 49450 39914
rect 49484 39880 49540 39914
rect 49574 39880 49630 39914
rect 49664 39880 49980 39914
rect 50014 39880 50070 39914
rect 50104 39880 50160 39914
rect 50194 39880 50250 39914
rect 50284 39880 50340 39914
rect 50374 39880 50430 39914
rect 50464 39880 50520 39914
rect 50554 39880 50610 39914
rect 50644 39880 50700 39914
rect 50734 39880 50790 39914
rect 50824 39880 50880 39914
rect 50914 39880 50970 39914
rect 51004 39880 51320 39914
rect 51354 39880 51410 39914
rect 51444 39880 51500 39914
rect 51534 39880 51590 39914
rect 51624 39880 51680 39914
rect 51714 39880 51770 39914
rect 51804 39880 51860 39914
rect 51894 39880 51950 39914
rect 51984 39880 52040 39914
rect 52074 39880 52130 39914
rect 52164 39880 52220 39914
rect 52254 39880 52310 39914
rect 52344 39880 52478 39914
rect 41810 39848 52478 39880
rect 37216 39709 37256 39752
rect 37216 39675 37219 39709
rect 37253 39675 37256 39709
rect 37216 39632 37256 39675
rect 38276 39679 38396 39682
rect 38276 39645 38321 39679
rect 38355 39645 38396 39679
rect 38276 39632 38396 39645
rect 39576 39679 39696 39682
rect 39576 39645 39621 39679
rect 39655 39645 39696 39679
rect 39576 39632 39696 39645
rect 12018 37341 13306 37376
rect 12018 37318 12148 37341
rect 12018 37284 12052 37318
rect 12086 37307 12148 37318
rect 12182 37307 12238 37341
rect 12272 37307 12328 37341
rect 12362 37307 12418 37341
rect 12452 37307 12508 37341
rect 12542 37307 12598 37341
rect 12632 37307 12688 37341
rect 12722 37307 12778 37341
rect 12812 37307 12868 37341
rect 12902 37307 12958 37341
rect 12992 37307 13048 37341
rect 13082 37307 13138 37341
rect 13172 37318 13306 37341
rect 13172 37307 13239 37318
rect 12086 37284 13239 37307
rect 13273 37284 13306 37318
rect 12018 37275 13306 37284
rect 12018 37228 12119 37275
rect 12018 37194 12052 37228
rect 12086 37194 12119 37228
rect 13205 37228 13306 37275
rect 12018 37138 12119 37194
rect 12018 37104 12052 37138
rect 12086 37104 12119 37138
rect 12018 37048 12119 37104
rect 12018 37014 12052 37048
rect 12086 37014 12119 37048
rect 12018 36958 12119 37014
rect 12018 36924 12052 36958
rect 12086 36924 12119 36958
rect 12018 36868 12119 36924
rect 12018 36834 12052 36868
rect 12086 36834 12119 36868
rect 12018 36778 12119 36834
rect 12018 36744 12052 36778
rect 12086 36744 12119 36778
rect 12018 36688 12119 36744
rect 12018 36654 12052 36688
rect 12086 36654 12119 36688
rect 12018 36598 12119 36654
rect 12018 36564 12052 36598
rect 12086 36564 12119 36598
rect 12018 36508 12119 36564
rect 12018 36474 12052 36508
rect 12086 36474 12119 36508
rect 12018 36418 12119 36474
rect 12018 36384 12052 36418
rect 12086 36384 12119 36418
rect 12018 36328 12119 36384
rect 12018 36294 12052 36328
rect 12086 36294 12119 36328
rect 12018 36238 12119 36294
rect 13205 37194 13239 37228
rect 13273 37194 13306 37228
rect 13205 37138 13306 37194
rect 13205 37104 13239 37138
rect 13273 37104 13306 37138
rect 13205 37048 13306 37104
rect 13205 37014 13239 37048
rect 13273 37014 13306 37048
rect 13205 36958 13306 37014
rect 13205 36924 13239 36958
rect 13273 36924 13306 36958
rect 13205 36868 13306 36924
rect 13205 36834 13239 36868
rect 13273 36834 13306 36868
rect 13205 36778 13306 36834
rect 13205 36744 13239 36778
rect 13273 36744 13306 36778
rect 13205 36688 13306 36744
rect 13205 36654 13239 36688
rect 13273 36654 13306 36688
rect 13205 36598 13306 36654
rect 13205 36564 13239 36598
rect 13273 36564 13306 36598
rect 14590 36723 15206 36762
rect 14590 36621 14677 36723
rect 15119 36621 15206 36723
rect 14590 36582 15206 36621
rect 17334 36723 17950 36762
rect 17334 36621 17421 36723
rect 17863 36621 17950 36723
rect 17334 36582 17950 36621
rect 20366 36723 20982 36762
rect 20366 36621 20453 36723
rect 20895 36621 20982 36723
rect 20366 36582 20982 36621
rect 23410 36723 24026 36762
rect 23410 36621 23497 36723
rect 23939 36621 24026 36723
rect 23410 36582 24026 36621
rect 13205 36508 13306 36564
rect 13205 36474 13239 36508
rect 13273 36474 13306 36508
rect 13205 36418 13306 36474
rect 13205 36384 13239 36418
rect 13273 36384 13306 36418
rect 13205 36328 13306 36384
rect 13205 36294 13239 36328
rect 13273 36294 13306 36328
rect 12018 36204 12052 36238
rect 12086 36204 12119 36238
rect 12018 36189 12119 36204
rect 13205 36238 13306 36294
rect 13205 36204 13239 36238
rect 13273 36204 13306 36238
rect 13205 36189 13306 36204
rect 12018 36154 13306 36189
rect 12018 36120 12148 36154
rect 12182 36120 12238 36154
rect 12272 36120 12328 36154
rect 12362 36120 12418 36154
rect 12452 36120 12508 36154
rect 12542 36120 12598 36154
rect 12632 36120 12688 36154
rect 12722 36120 12778 36154
rect 12812 36120 12868 36154
rect 12902 36120 12958 36154
rect 12992 36120 13048 36154
rect 13082 36120 13138 36154
rect 13172 36120 13306 36154
rect 12018 36088 13306 36120
rect 41810 37341 52478 37376
rect 41810 37318 41940 37341
rect 41810 37284 41844 37318
rect 41878 37307 41940 37318
rect 41974 37307 42030 37341
rect 42064 37307 42120 37341
rect 42154 37307 42210 37341
rect 42244 37307 42300 37341
rect 42334 37307 42390 37341
rect 42424 37307 42480 37341
rect 42514 37307 42570 37341
rect 42604 37307 42660 37341
rect 42694 37307 42750 37341
rect 42784 37307 42840 37341
rect 42874 37307 42930 37341
rect 42964 37318 43280 37341
rect 42964 37307 43031 37318
rect 41878 37284 43031 37307
rect 43065 37284 43184 37318
rect 43218 37307 43280 37318
rect 43314 37307 43370 37341
rect 43404 37307 43460 37341
rect 43494 37307 43550 37341
rect 43584 37307 43640 37341
rect 43674 37307 43730 37341
rect 43764 37307 43820 37341
rect 43854 37307 43910 37341
rect 43944 37307 44000 37341
rect 44034 37307 44090 37341
rect 44124 37307 44180 37341
rect 44214 37307 44270 37341
rect 44304 37318 44620 37341
rect 44304 37307 44371 37318
rect 43218 37284 44371 37307
rect 44405 37284 44524 37318
rect 44558 37307 44620 37318
rect 44654 37307 44710 37341
rect 44744 37307 44800 37341
rect 44834 37307 44890 37341
rect 44924 37307 44980 37341
rect 45014 37307 45070 37341
rect 45104 37307 45160 37341
rect 45194 37307 45250 37341
rect 45284 37307 45340 37341
rect 45374 37307 45430 37341
rect 45464 37307 45520 37341
rect 45554 37307 45610 37341
rect 45644 37318 45960 37341
rect 45644 37307 45711 37318
rect 44558 37284 45711 37307
rect 45745 37284 45864 37318
rect 45898 37307 45960 37318
rect 45994 37307 46050 37341
rect 46084 37307 46140 37341
rect 46174 37307 46230 37341
rect 46264 37307 46320 37341
rect 46354 37307 46410 37341
rect 46444 37307 46500 37341
rect 46534 37307 46590 37341
rect 46624 37307 46680 37341
rect 46714 37307 46770 37341
rect 46804 37307 46860 37341
rect 46894 37307 46950 37341
rect 46984 37318 47300 37341
rect 46984 37307 47051 37318
rect 45898 37284 47051 37307
rect 47085 37284 47204 37318
rect 47238 37307 47300 37318
rect 47334 37307 47390 37341
rect 47424 37307 47480 37341
rect 47514 37307 47570 37341
rect 47604 37307 47660 37341
rect 47694 37307 47750 37341
rect 47784 37307 47840 37341
rect 47874 37307 47930 37341
rect 47964 37307 48020 37341
rect 48054 37307 48110 37341
rect 48144 37307 48200 37341
rect 48234 37307 48290 37341
rect 48324 37318 48640 37341
rect 48324 37307 48391 37318
rect 47238 37284 48391 37307
rect 48425 37284 48544 37318
rect 48578 37307 48640 37318
rect 48674 37307 48730 37341
rect 48764 37307 48820 37341
rect 48854 37307 48910 37341
rect 48944 37307 49000 37341
rect 49034 37307 49090 37341
rect 49124 37307 49180 37341
rect 49214 37307 49270 37341
rect 49304 37307 49360 37341
rect 49394 37307 49450 37341
rect 49484 37307 49540 37341
rect 49574 37307 49630 37341
rect 49664 37318 49980 37341
rect 49664 37307 49731 37318
rect 48578 37284 49731 37307
rect 49765 37284 49884 37318
rect 49918 37307 49980 37318
rect 50014 37307 50070 37341
rect 50104 37307 50160 37341
rect 50194 37307 50250 37341
rect 50284 37307 50340 37341
rect 50374 37307 50430 37341
rect 50464 37307 50520 37341
rect 50554 37307 50610 37341
rect 50644 37307 50700 37341
rect 50734 37307 50790 37341
rect 50824 37307 50880 37341
rect 50914 37307 50970 37341
rect 51004 37318 51320 37341
rect 51004 37307 51071 37318
rect 49918 37284 51071 37307
rect 51105 37284 51224 37318
rect 51258 37307 51320 37318
rect 51354 37307 51410 37341
rect 51444 37307 51500 37341
rect 51534 37307 51590 37341
rect 51624 37307 51680 37341
rect 51714 37307 51770 37341
rect 51804 37307 51860 37341
rect 51894 37307 51950 37341
rect 51984 37307 52040 37341
rect 52074 37307 52130 37341
rect 52164 37307 52220 37341
rect 52254 37307 52310 37341
rect 52344 37318 52478 37341
rect 52344 37307 52411 37318
rect 51258 37284 52411 37307
rect 52445 37284 52478 37318
rect 41810 37275 52478 37284
rect 41810 37228 41911 37275
rect 41810 37194 41844 37228
rect 41878 37194 41911 37228
rect 42997 37228 43251 37275
rect 41810 37138 41911 37194
rect 41810 37104 41844 37138
rect 41878 37104 41911 37138
rect 41810 37048 41911 37104
rect 41810 37014 41844 37048
rect 41878 37014 41911 37048
rect 41810 36958 41911 37014
rect 41810 36924 41844 36958
rect 41878 36924 41911 36958
rect 41810 36868 41911 36924
rect 41810 36834 41844 36868
rect 41878 36834 41911 36868
rect 41810 36778 41911 36834
rect 41810 36744 41844 36778
rect 41878 36744 41911 36778
rect 41810 36688 41911 36744
rect 41810 36654 41844 36688
rect 41878 36654 41911 36688
rect 41810 36598 41911 36654
rect 41810 36564 41844 36598
rect 41878 36564 41911 36598
rect 41810 36508 41911 36564
rect 41810 36474 41844 36508
rect 41878 36474 41911 36508
rect 41810 36418 41911 36474
rect 41810 36384 41844 36418
rect 41878 36384 41911 36418
rect 41810 36328 41911 36384
rect 41810 36294 41844 36328
rect 41878 36294 41911 36328
rect 41810 36238 41911 36294
rect 42997 37194 43031 37228
rect 43065 37194 43184 37228
rect 43218 37194 43251 37228
rect 44337 37228 44591 37275
rect 42997 37138 43251 37194
rect 42997 37104 43031 37138
rect 43065 37104 43184 37138
rect 43218 37104 43251 37138
rect 42997 37048 43251 37104
rect 42997 37014 43031 37048
rect 43065 37014 43184 37048
rect 43218 37014 43251 37048
rect 42997 36958 43251 37014
rect 42997 36924 43031 36958
rect 43065 36924 43184 36958
rect 43218 36924 43251 36958
rect 42997 36868 43251 36924
rect 42997 36834 43031 36868
rect 43065 36834 43184 36868
rect 43218 36834 43251 36868
rect 42997 36778 43251 36834
rect 42997 36744 43031 36778
rect 43065 36744 43184 36778
rect 43218 36744 43251 36778
rect 42997 36688 43251 36744
rect 42997 36654 43031 36688
rect 43065 36654 43184 36688
rect 43218 36654 43251 36688
rect 42997 36598 43251 36654
rect 42997 36564 43031 36598
rect 43065 36564 43184 36598
rect 43218 36564 43251 36598
rect 42997 36508 43251 36564
rect 42997 36474 43031 36508
rect 43065 36474 43184 36508
rect 43218 36474 43251 36508
rect 42997 36418 43251 36474
rect 42997 36384 43031 36418
rect 43065 36384 43184 36418
rect 43218 36384 43251 36418
rect 42997 36328 43251 36384
rect 42997 36294 43031 36328
rect 43065 36294 43184 36328
rect 43218 36294 43251 36328
rect 41810 36204 41844 36238
rect 41878 36204 41911 36238
rect 41810 36189 41911 36204
rect 42997 36238 43251 36294
rect 44337 37194 44371 37228
rect 44405 37194 44524 37228
rect 44558 37194 44591 37228
rect 45677 37228 45931 37275
rect 44337 37138 44591 37194
rect 44337 37104 44371 37138
rect 44405 37104 44524 37138
rect 44558 37104 44591 37138
rect 44337 37048 44591 37104
rect 44337 37014 44371 37048
rect 44405 37014 44524 37048
rect 44558 37014 44591 37048
rect 44337 36958 44591 37014
rect 44337 36924 44371 36958
rect 44405 36924 44524 36958
rect 44558 36924 44591 36958
rect 44337 36868 44591 36924
rect 44337 36834 44371 36868
rect 44405 36834 44524 36868
rect 44558 36834 44591 36868
rect 44337 36778 44591 36834
rect 44337 36744 44371 36778
rect 44405 36744 44524 36778
rect 44558 36744 44591 36778
rect 44337 36688 44591 36744
rect 44337 36654 44371 36688
rect 44405 36654 44524 36688
rect 44558 36654 44591 36688
rect 44337 36598 44591 36654
rect 44337 36564 44371 36598
rect 44405 36564 44524 36598
rect 44558 36564 44591 36598
rect 44337 36508 44591 36564
rect 44337 36474 44371 36508
rect 44405 36474 44524 36508
rect 44558 36474 44591 36508
rect 44337 36418 44591 36474
rect 44337 36384 44371 36418
rect 44405 36384 44524 36418
rect 44558 36384 44591 36418
rect 44337 36328 44591 36384
rect 44337 36294 44371 36328
rect 44405 36294 44524 36328
rect 44558 36294 44591 36328
rect 42997 36204 43031 36238
rect 43065 36204 43184 36238
rect 43218 36204 43251 36238
rect 42997 36189 43251 36204
rect 44337 36238 44591 36294
rect 45677 37194 45711 37228
rect 45745 37194 45864 37228
rect 45898 37194 45931 37228
rect 47017 37228 47271 37275
rect 45677 37138 45931 37194
rect 45677 37104 45711 37138
rect 45745 37104 45864 37138
rect 45898 37104 45931 37138
rect 45677 37048 45931 37104
rect 45677 37014 45711 37048
rect 45745 37014 45864 37048
rect 45898 37014 45931 37048
rect 45677 36958 45931 37014
rect 45677 36924 45711 36958
rect 45745 36924 45864 36958
rect 45898 36924 45931 36958
rect 45677 36868 45931 36924
rect 45677 36834 45711 36868
rect 45745 36834 45864 36868
rect 45898 36834 45931 36868
rect 45677 36778 45931 36834
rect 45677 36744 45711 36778
rect 45745 36744 45864 36778
rect 45898 36744 45931 36778
rect 45677 36688 45931 36744
rect 45677 36654 45711 36688
rect 45745 36654 45864 36688
rect 45898 36654 45931 36688
rect 45677 36598 45931 36654
rect 45677 36564 45711 36598
rect 45745 36564 45864 36598
rect 45898 36564 45931 36598
rect 45677 36508 45931 36564
rect 45677 36474 45711 36508
rect 45745 36474 45864 36508
rect 45898 36474 45931 36508
rect 45677 36418 45931 36474
rect 45677 36384 45711 36418
rect 45745 36384 45864 36418
rect 45898 36384 45931 36418
rect 45677 36328 45931 36384
rect 45677 36294 45711 36328
rect 45745 36294 45864 36328
rect 45898 36294 45931 36328
rect 44337 36204 44371 36238
rect 44405 36204 44524 36238
rect 44558 36204 44591 36238
rect 44337 36189 44591 36204
rect 45677 36238 45931 36294
rect 47017 37194 47051 37228
rect 47085 37194 47204 37228
rect 47238 37194 47271 37228
rect 48357 37228 48611 37275
rect 47017 37138 47271 37194
rect 47017 37104 47051 37138
rect 47085 37104 47204 37138
rect 47238 37104 47271 37138
rect 47017 37048 47271 37104
rect 47017 37014 47051 37048
rect 47085 37014 47204 37048
rect 47238 37014 47271 37048
rect 47017 36958 47271 37014
rect 47017 36924 47051 36958
rect 47085 36924 47204 36958
rect 47238 36924 47271 36958
rect 47017 36868 47271 36924
rect 47017 36834 47051 36868
rect 47085 36834 47204 36868
rect 47238 36834 47271 36868
rect 47017 36778 47271 36834
rect 47017 36744 47051 36778
rect 47085 36744 47204 36778
rect 47238 36744 47271 36778
rect 47017 36688 47271 36744
rect 47017 36654 47051 36688
rect 47085 36654 47204 36688
rect 47238 36654 47271 36688
rect 47017 36598 47271 36654
rect 47017 36564 47051 36598
rect 47085 36564 47204 36598
rect 47238 36564 47271 36598
rect 47017 36508 47271 36564
rect 47017 36474 47051 36508
rect 47085 36474 47204 36508
rect 47238 36474 47271 36508
rect 47017 36418 47271 36474
rect 47017 36384 47051 36418
rect 47085 36384 47204 36418
rect 47238 36384 47271 36418
rect 47017 36328 47271 36384
rect 47017 36294 47051 36328
rect 47085 36294 47204 36328
rect 47238 36294 47271 36328
rect 45677 36204 45711 36238
rect 45745 36204 45864 36238
rect 45898 36204 45931 36238
rect 45677 36189 45931 36204
rect 47017 36238 47271 36294
rect 48357 37194 48391 37228
rect 48425 37194 48544 37228
rect 48578 37194 48611 37228
rect 49697 37228 49951 37275
rect 48357 37138 48611 37194
rect 48357 37104 48391 37138
rect 48425 37104 48544 37138
rect 48578 37104 48611 37138
rect 48357 37048 48611 37104
rect 48357 37014 48391 37048
rect 48425 37014 48544 37048
rect 48578 37014 48611 37048
rect 48357 36958 48611 37014
rect 48357 36924 48391 36958
rect 48425 36924 48544 36958
rect 48578 36924 48611 36958
rect 48357 36868 48611 36924
rect 48357 36834 48391 36868
rect 48425 36834 48544 36868
rect 48578 36834 48611 36868
rect 48357 36778 48611 36834
rect 48357 36744 48391 36778
rect 48425 36744 48544 36778
rect 48578 36744 48611 36778
rect 48357 36688 48611 36744
rect 48357 36654 48391 36688
rect 48425 36654 48544 36688
rect 48578 36654 48611 36688
rect 48357 36598 48611 36654
rect 48357 36564 48391 36598
rect 48425 36564 48544 36598
rect 48578 36564 48611 36598
rect 48357 36508 48611 36564
rect 48357 36474 48391 36508
rect 48425 36474 48544 36508
rect 48578 36474 48611 36508
rect 48357 36418 48611 36474
rect 48357 36384 48391 36418
rect 48425 36384 48544 36418
rect 48578 36384 48611 36418
rect 48357 36328 48611 36384
rect 48357 36294 48391 36328
rect 48425 36294 48544 36328
rect 48578 36294 48611 36328
rect 47017 36204 47051 36238
rect 47085 36204 47204 36238
rect 47238 36204 47271 36238
rect 47017 36189 47271 36204
rect 48357 36238 48611 36294
rect 49697 37194 49731 37228
rect 49765 37194 49884 37228
rect 49918 37194 49951 37228
rect 51037 37228 51291 37275
rect 49697 37138 49951 37194
rect 49697 37104 49731 37138
rect 49765 37104 49884 37138
rect 49918 37104 49951 37138
rect 49697 37048 49951 37104
rect 49697 37014 49731 37048
rect 49765 37014 49884 37048
rect 49918 37014 49951 37048
rect 49697 36958 49951 37014
rect 49697 36924 49731 36958
rect 49765 36924 49884 36958
rect 49918 36924 49951 36958
rect 49697 36868 49951 36924
rect 49697 36834 49731 36868
rect 49765 36834 49884 36868
rect 49918 36834 49951 36868
rect 49697 36778 49951 36834
rect 49697 36744 49731 36778
rect 49765 36744 49884 36778
rect 49918 36744 49951 36778
rect 49697 36688 49951 36744
rect 49697 36654 49731 36688
rect 49765 36654 49884 36688
rect 49918 36654 49951 36688
rect 49697 36598 49951 36654
rect 49697 36564 49731 36598
rect 49765 36564 49884 36598
rect 49918 36564 49951 36598
rect 49697 36508 49951 36564
rect 49697 36474 49731 36508
rect 49765 36474 49884 36508
rect 49918 36474 49951 36508
rect 49697 36418 49951 36474
rect 49697 36384 49731 36418
rect 49765 36384 49884 36418
rect 49918 36384 49951 36418
rect 49697 36328 49951 36384
rect 49697 36294 49731 36328
rect 49765 36294 49884 36328
rect 49918 36294 49951 36328
rect 48357 36204 48391 36238
rect 48425 36204 48544 36238
rect 48578 36204 48611 36238
rect 48357 36189 48611 36204
rect 49697 36238 49951 36294
rect 51037 37194 51071 37228
rect 51105 37194 51224 37228
rect 51258 37194 51291 37228
rect 52377 37228 52478 37275
rect 51037 37138 51291 37194
rect 51037 37104 51071 37138
rect 51105 37104 51224 37138
rect 51258 37104 51291 37138
rect 51037 37048 51291 37104
rect 51037 37014 51071 37048
rect 51105 37014 51224 37048
rect 51258 37014 51291 37048
rect 51037 36958 51291 37014
rect 51037 36924 51071 36958
rect 51105 36924 51224 36958
rect 51258 36924 51291 36958
rect 51037 36868 51291 36924
rect 51037 36834 51071 36868
rect 51105 36834 51224 36868
rect 51258 36834 51291 36868
rect 51037 36778 51291 36834
rect 51037 36744 51071 36778
rect 51105 36744 51224 36778
rect 51258 36744 51291 36778
rect 51037 36688 51291 36744
rect 51037 36654 51071 36688
rect 51105 36654 51224 36688
rect 51258 36654 51291 36688
rect 51037 36598 51291 36654
rect 51037 36564 51071 36598
rect 51105 36564 51224 36598
rect 51258 36564 51291 36598
rect 51037 36508 51291 36564
rect 51037 36474 51071 36508
rect 51105 36474 51224 36508
rect 51258 36474 51291 36508
rect 51037 36418 51291 36474
rect 51037 36384 51071 36418
rect 51105 36384 51224 36418
rect 51258 36384 51291 36418
rect 51037 36328 51291 36384
rect 51037 36294 51071 36328
rect 51105 36294 51224 36328
rect 51258 36294 51291 36328
rect 49697 36204 49731 36238
rect 49765 36204 49884 36238
rect 49918 36204 49951 36238
rect 49697 36189 49951 36204
rect 51037 36238 51291 36294
rect 52377 37194 52411 37228
rect 52445 37194 52478 37228
rect 52377 37138 52478 37194
rect 52377 37104 52411 37138
rect 52445 37104 52478 37138
rect 52377 37048 52478 37104
rect 52377 37014 52411 37048
rect 52445 37014 52478 37048
rect 52377 36958 52478 37014
rect 52377 36924 52411 36958
rect 52445 36924 52478 36958
rect 52377 36868 52478 36924
rect 52377 36834 52411 36868
rect 52445 36834 52478 36868
rect 52377 36778 52478 36834
rect 52377 36744 52411 36778
rect 52445 36744 52478 36778
rect 52377 36688 52478 36744
rect 52377 36654 52411 36688
rect 52445 36654 52478 36688
rect 52377 36598 52478 36654
rect 52377 36564 52411 36598
rect 52445 36564 52478 36598
rect 52377 36508 52478 36564
rect 52377 36474 52411 36508
rect 52445 36474 52478 36508
rect 52377 36418 52478 36474
rect 52377 36384 52411 36418
rect 52445 36384 52478 36418
rect 52377 36328 52478 36384
rect 52377 36294 52411 36328
rect 52445 36294 52478 36328
rect 51037 36204 51071 36238
rect 51105 36204 51224 36238
rect 51258 36204 51291 36238
rect 51037 36189 51291 36204
rect 52377 36238 52478 36294
rect 52377 36204 52411 36238
rect 52445 36204 52478 36238
rect 52377 36189 52478 36204
rect 41810 36154 52478 36189
rect 25358 35949 25398 35992
rect 41810 36120 41940 36154
rect 41974 36120 42030 36154
rect 42064 36120 42120 36154
rect 42154 36120 42210 36154
rect 42244 36120 42300 36154
rect 42334 36120 42390 36154
rect 42424 36120 42480 36154
rect 42514 36120 42570 36154
rect 42604 36120 42660 36154
rect 42694 36120 42750 36154
rect 42784 36120 42840 36154
rect 42874 36120 42930 36154
rect 42964 36120 43280 36154
rect 43314 36120 43370 36154
rect 43404 36120 43460 36154
rect 43494 36120 43550 36154
rect 43584 36120 43640 36154
rect 43674 36120 43730 36154
rect 43764 36120 43820 36154
rect 43854 36120 43910 36154
rect 43944 36120 44000 36154
rect 44034 36120 44090 36154
rect 44124 36120 44180 36154
rect 44214 36120 44270 36154
rect 44304 36120 44620 36154
rect 44654 36120 44710 36154
rect 44744 36120 44800 36154
rect 44834 36120 44890 36154
rect 44924 36120 44980 36154
rect 45014 36120 45070 36154
rect 45104 36120 45160 36154
rect 45194 36120 45250 36154
rect 45284 36120 45340 36154
rect 45374 36120 45430 36154
rect 45464 36120 45520 36154
rect 45554 36120 45610 36154
rect 45644 36120 45960 36154
rect 45994 36120 46050 36154
rect 46084 36120 46140 36154
rect 46174 36120 46230 36154
rect 46264 36120 46320 36154
rect 46354 36120 46410 36154
rect 46444 36120 46500 36154
rect 46534 36120 46590 36154
rect 46624 36120 46680 36154
rect 46714 36120 46770 36154
rect 46804 36120 46860 36154
rect 46894 36120 46950 36154
rect 46984 36120 47300 36154
rect 47334 36120 47390 36154
rect 47424 36120 47480 36154
rect 47514 36120 47570 36154
rect 47604 36120 47660 36154
rect 47694 36120 47750 36154
rect 47784 36120 47840 36154
rect 47874 36120 47930 36154
rect 47964 36120 48020 36154
rect 48054 36120 48110 36154
rect 48144 36120 48200 36154
rect 48234 36120 48290 36154
rect 48324 36120 48640 36154
rect 48674 36120 48730 36154
rect 48764 36120 48820 36154
rect 48854 36120 48910 36154
rect 48944 36120 49000 36154
rect 49034 36120 49090 36154
rect 49124 36120 49180 36154
rect 49214 36120 49270 36154
rect 49304 36120 49360 36154
rect 49394 36120 49450 36154
rect 49484 36120 49540 36154
rect 49574 36120 49630 36154
rect 49664 36120 49980 36154
rect 50014 36120 50070 36154
rect 50104 36120 50160 36154
rect 50194 36120 50250 36154
rect 50284 36120 50340 36154
rect 50374 36120 50430 36154
rect 50464 36120 50520 36154
rect 50554 36120 50610 36154
rect 50644 36120 50700 36154
rect 50734 36120 50790 36154
rect 50824 36120 50880 36154
rect 50914 36120 50970 36154
rect 51004 36120 51320 36154
rect 51354 36120 51410 36154
rect 51444 36120 51500 36154
rect 51534 36120 51590 36154
rect 51624 36120 51680 36154
rect 51714 36120 51770 36154
rect 51804 36120 51860 36154
rect 51894 36120 51950 36154
rect 51984 36120 52040 36154
rect 52074 36120 52130 36154
rect 52164 36120 52220 36154
rect 52254 36120 52310 36154
rect 52344 36120 52478 36154
rect 41810 36088 52478 36120
rect 25358 35915 25361 35949
rect 25395 35915 25398 35949
rect 25358 35872 25398 35915
rect 26418 35919 26538 35922
rect 26418 35885 26463 35919
rect 26497 35885 26538 35919
rect 26418 35872 26538 35885
rect 27718 35919 27838 35922
rect 27718 35885 27763 35919
rect 27797 35885 27838 35919
rect 27718 35872 27838 35885
rect 41810 33581 52478 33616
rect 41810 33558 41940 33581
rect 41810 33524 41844 33558
rect 41878 33547 41940 33558
rect 41974 33547 42030 33581
rect 42064 33547 42120 33581
rect 42154 33547 42210 33581
rect 42244 33547 42300 33581
rect 42334 33547 42390 33581
rect 42424 33547 42480 33581
rect 42514 33547 42570 33581
rect 42604 33547 42660 33581
rect 42694 33547 42750 33581
rect 42784 33547 42840 33581
rect 42874 33547 42930 33581
rect 42964 33558 43280 33581
rect 42964 33547 43031 33558
rect 41878 33524 43031 33547
rect 43065 33524 43184 33558
rect 43218 33547 43280 33558
rect 43314 33547 43370 33581
rect 43404 33547 43460 33581
rect 43494 33547 43550 33581
rect 43584 33547 43640 33581
rect 43674 33547 43730 33581
rect 43764 33547 43820 33581
rect 43854 33547 43910 33581
rect 43944 33547 44000 33581
rect 44034 33547 44090 33581
rect 44124 33547 44180 33581
rect 44214 33547 44270 33581
rect 44304 33558 44620 33581
rect 44304 33547 44371 33558
rect 43218 33524 44371 33547
rect 44405 33524 44524 33558
rect 44558 33547 44620 33558
rect 44654 33547 44710 33581
rect 44744 33547 44800 33581
rect 44834 33547 44890 33581
rect 44924 33547 44980 33581
rect 45014 33547 45070 33581
rect 45104 33547 45160 33581
rect 45194 33547 45250 33581
rect 45284 33547 45340 33581
rect 45374 33547 45430 33581
rect 45464 33547 45520 33581
rect 45554 33547 45610 33581
rect 45644 33558 45960 33581
rect 45644 33547 45711 33558
rect 44558 33524 45711 33547
rect 45745 33524 45864 33558
rect 45898 33547 45960 33558
rect 45994 33547 46050 33581
rect 46084 33547 46140 33581
rect 46174 33547 46230 33581
rect 46264 33547 46320 33581
rect 46354 33547 46410 33581
rect 46444 33547 46500 33581
rect 46534 33547 46590 33581
rect 46624 33547 46680 33581
rect 46714 33547 46770 33581
rect 46804 33547 46860 33581
rect 46894 33547 46950 33581
rect 46984 33558 47300 33581
rect 46984 33547 47051 33558
rect 45898 33524 47051 33547
rect 47085 33524 47204 33558
rect 47238 33547 47300 33558
rect 47334 33547 47390 33581
rect 47424 33547 47480 33581
rect 47514 33547 47570 33581
rect 47604 33547 47660 33581
rect 47694 33547 47750 33581
rect 47784 33547 47840 33581
rect 47874 33547 47930 33581
rect 47964 33547 48020 33581
rect 48054 33547 48110 33581
rect 48144 33547 48200 33581
rect 48234 33547 48290 33581
rect 48324 33558 48640 33581
rect 48324 33547 48391 33558
rect 47238 33524 48391 33547
rect 48425 33524 48544 33558
rect 48578 33547 48640 33558
rect 48674 33547 48730 33581
rect 48764 33547 48820 33581
rect 48854 33547 48910 33581
rect 48944 33547 49000 33581
rect 49034 33547 49090 33581
rect 49124 33547 49180 33581
rect 49214 33547 49270 33581
rect 49304 33547 49360 33581
rect 49394 33547 49450 33581
rect 49484 33547 49540 33581
rect 49574 33547 49630 33581
rect 49664 33558 49980 33581
rect 49664 33547 49731 33558
rect 48578 33524 49731 33547
rect 49765 33524 49884 33558
rect 49918 33547 49980 33558
rect 50014 33547 50070 33581
rect 50104 33547 50160 33581
rect 50194 33547 50250 33581
rect 50284 33547 50340 33581
rect 50374 33547 50430 33581
rect 50464 33547 50520 33581
rect 50554 33547 50610 33581
rect 50644 33547 50700 33581
rect 50734 33547 50790 33581
rect 50824 33547 50880 33581
rect 50914 33547 50970 33581
rect 51004 33558 51320 33581
rect 51004 33547 51071 33558
rect 49918 33524 51071 33547
rect 51105 33524 51224 33558
rect 51258 33547 51320 33558
rect 51354 33547 51410 33581
rect 51444 33547 51500 33581
rect 51534 33547 51590 33581
rect 51624 33547 51680 33581
rect 51714 33547 51770 33581
rect 51804 33547 51860 33581
rect 51894 33547 51950 33581
rect 51984 33547 52040 33581
rect 52074 33547 52130 33581
rect 52164 33547 52220 33581
rect 52254 33547 52310 33581
rect 52344 33558 52478 33581
rect 52344 33547 52411 33558
rect 51258 33524 52411 33547
rect 52445 33524 52478 33558
rect 41810 33515 52478 33524
rect 41810 33468 41911 33515
rect 41810 33434 41844 33468
rect 41878 33434 41911 33468
rect 42997 33468 43251 33515
rect 41810 33378 41911 33434
rect 41810 33344 41844 33378
rect 41878 33344 41911 33378
rect 41810 33288 41911 33344
rect 41810 33254 41844 33288
rect 41878 33254 41911 33288
rect 41810 33198 41911 33254
rect 41810 33164 41844 33198
rect 41878 33164 41911 33198
rect 41810 33108 41911 33164
rect 41810 33074 41844 33108
rect 41878 33074 41911 33108
rect 41810 33018 41911 33074
rect 20176 32963 20792 33002
rect 20176 32861 20263 32963
rect 20705 32861 20792 32963
rect 20176 32822 20792 32861
rect 23208 32963 23824 33002
rect 23208 32861 23295 32963
rect 23737 32861 23824 32963
rect 23208 32822 23824 32861
rect 41810 32984 41844 33018
rect 41878 32984 41911 33018
rect 41810 32928 41911 32984
rect 41810 32894 41844 32928
rect 41878 32894 41911 32928
rect 41810 32838 41911 32894
rect 41810 32804 41844 32838
rect 41878 32804 41911 32838
rect 41810 32748 41911 32804
rect 41810 32714 41844 32748
rect 41878 32714 41911 32748
rect 41810 32658 41911 32714
rect 41810 32624 41844 32658
rect 41878 32624 41911 32658
rect 41810 32568 41911 32624
rect 41810 32534 41844 32568
rect 41878 32534 41911 32568
rect 41810 32478 41911 32534
rect 42997 33434 43031 33468
rect 43065 33434 43184 33468
rect 43218 33434 43251 33468
rect 44337 33468 44591 33515
rect 42997 33378 43251 33434
rect 42997 33344 43031 33378
rect 43065 33344 43184 33378
rect 43218 33344 43251 33378
rect 42997 33288 43251 33344
rect 42997 33254 43031 33288
rect 43065 33254 43184 33288
rect 43218 33254 43251 33288
rect 42997 33198 43251 33254
rect 42997 33164 43031 33198
rect 43065 33164 43184 33198
rect 43218 33164 43251 33198
rect 42997 33108 43251 33164
rect 42997 33074 43031 33108
rect 43065 33074 43184 33108
rect 43218 33074 43251 33108
rect 42997 33018 43251 33074
rect 42997 32984 43031 33018
rect 43065 32984 43184 33018
rect 43218 32984 43251 33018
rect 42997 32928 43251 32984
rect 42997 32894 43031 32928
rect 43065 32894 43184 32928
rect 43218 32894 43251 32928
rect 42997 32838 43251 32894
rect 42997 32804 43031 32838
rect 43065 32804 43184 32838
rect 43218 32804 43251 32838
rect 42997 32748 43251 32804
rect 42997 32714 43031 32748
rect 43065 32714 43184 32748
rect 43218 32714 43251 32748
rect 42997 32658 43251 32714
rect 42997 32624 43031 32658
rect 43065 32624 43184 32658
rect 43218 32624 43251 32658
rect 42997 32568 43251 32624
rect 42997 32534 43031 32568
rect 43065 32534 43184 32568
rect 43218 32534 43251 32568
rect 41810 32444 41844 32478
rect 41878 32444 41911 32478
rect 41810 32429 41911 32444
rect 42997 32478 43251 32534
rect 44337 33434 44371 33468
rect 44405 33434 44524 33468
rect 44558 33434 44591 33468
rect 45677 33468 45931 33515
rect 44337 33378 44591 33434
rect 44337 33344 44371 33378
rect 44405 33344 44524 33378
rect 44558 33344 44591 33378
rect 44337 33288 44591 33344
rect 44337 33254 44371 33288
rect 44405 33254 44524 33288
rect 44558 33254 44591 33288
rect 44337 33198 44591 33254
rect 44337 33164 44371 33198
rect 44405 33164 44524 33198
rect 44558 33164 44591 33198
rect 44337 33108 44591 33164
rect 44337 33074 44371 33108
rect 44405 33074 44524 33108
rect 44558 33074 44591 33108
rect 44337 33018 44591 33074
rect 44337 32984 44371 33018
rect 44405 32984 44524 33018
rect 44558 32984 44591 33018
rect 44337 32928 44591 32984
rect 44337 32894 44371 32928
rect 44405 32894 44524 32928
rect 44558 32894 44591 32928
rect 44337 32838 44591 32894
rect 44337 32804 44371 32838
rect 44405 32804 44524 32838
rect 44558 32804 44591 32838
rect 44337 32748 44591 32804
rect 44337 32714 44371 32748
rect 44405 32714 44524 32748
rect 44558 32714 44591 32748
rect 44337 32658 44591 32714
rect 44337 32624 44371 32658
rect 44405 32624 44524 32658
rect 44558 32624 44591 32658
rect 44337 32568 44591 32624
rect 44337 32534 44371 32568
rect 44405 32534 44524 32568
rect 44558 32534 44591 32568
rect 42997 32444 43031 32478
rect 43065 32444 43184 32478
rect 43218 32444 43251 32478
rect 42997 32429 43251 32444
rect 44337 32478 44591 32534
rect 45677 33434 45711 33468
rect 45745 33434 45864 33468
rect 45898 33434 45931 33468
rect 47017 33468 47271 33515
rect 45677 33378 45931 33434
rect 45677 33344 45711 33378
rect 45745 33344 45864 33378
rect 45898 33344 45931 33378
rect 45677 33288 45931 33344
rect 45677 33254 45711 33288
rect 45745 33254 45864 33288
rect 45898 33254 45931 33288
rect 45677 33198 45931 33254
rect 45677 33164 45711 33198
rect 45745 33164 45864 33198
rect 45898 33164 45931 33198
rect 45677 33108 45931 33164
rect 45677 33074 45711 33108
rect 45745 33074 45864 33108
rect 45898 33074 45931 33108
rect 45677 33018 45931 33074
rect 45677 32984 45711 33018
rect 45745 32984 45864 33018
rect 45898 32984 45931 33018
rect 45677 32928 45931 32984
rect 45677 32894 45711 32928
rect 45745 32894 45864 32928
rect 45898 32894 45931 32928
rect 45677 32838 45931 32894
rect 45677 32804 45711 32838
rect 45745 32804 45864 32838
rect 45898 32804 45931 32838
rect 45677 32748 45931 32804
rect 45677 32714 45711 32748
rect 45745 32714 45864 32748
rect 45898 32714 45931 32748
rect 45677 32658 45931 32714
rect 45677 32624 45711 32658
rect 45745 32624 45864 32658
rect 45898 32624 45931 32658
rect 45677 32568 45931 32624
rect 45677 32534 45711 32568
rect 45745 32534 45864 32568
rect 45898 32534 45931 32568
rect 44337 32444 44371 32478
rect 44405 32444 44524 32478
rect 44558 32444 44591 32478
rect 44337 32429 44591 32444
rect 45677 32478 45931 32534
rect 47017 33434 47051 33468
rect 47085 33434 47204 33468
rect 47238 33434 47271 33468
rect 48357 33468 48611 33515
rect 47017 33378 47271 33434
rect 47017 33344 47051 33378
rect 47085 33344 47204 33378
rect 47238 33344 47271 33378
rect 47017 33288 47271 33344
rect 47017 33254 47051 33288
rect 47085 33254 47204 33288
rect 47238 33254 47271 33288
rect 47017 33198 47271 33254
rect 47017 33164 47051 33198
rect 47085 33164 47204 33198
rect 47238 33164 47271 33198
rect 47017 33108 47271 33164
rect 47017 33074 47051 33108
rect 47085 33074 47204 33108
rect 47238 33074 47271 33108
rect 47017 33018 47271 33074
rect 47017 32984 47051 33018
rect 47085 32984 47204 33018
rect 47238 32984 47271 33018
rect 47017 32928 47271 32984
rect 47017 32894 47051 32928
rect 47085 32894 47204 32928
rect 47238 32894 47271 32928
rect 47017 32838 47271 32894
rect 47017 32804 47051 32838
rect 47085 32804 47204 32838
rect 47238 32804 47271 32838
rect 47017 32748 47271 32804
rect 47017 32714 47051 32748
rect 47085 32714 47204 32748
rect 47238 32714 47271 32748
rect 47017 32658 47271 32714
rect 47017 32624 47051 32658
rect 47085 32624 47204 32658
rect 47238 32624 47271 32658
rect 47017 32568 47271 32624
rect 47017 32534 47051 32568
rect 47085 32534 47204 32568
rect 47238 32534 47271 32568
rect 45677 32444 45711 32478
rect 45745 32444 45864 32478
rect 45898 32444 45931 32478
rect 45677 32429 45931 32444
rect 47017 32478 47271 32534
rect 48357 33434 48391 33468
rect 48425 33434 48544 33468
rect 48578 33434 48611 33468
rect 49697 33468 49951 33515
rect 48357 33378 48611 33434
rect 48357 33344 48391 33378
rect 48425 33344 48544 33378
rect 48578 33344 48611 33378
rect 48357 33288 48611 33344
rect 48357 33254 48391 33288
rect 48425 33254 48544 33288
rect 48578 33254 48611 33288
rect 48357 33198 48611 33254
rect 48357 33164 48391 33198
rect 48425 33164 48544 33198
rect 48578 33164 48611 33198
rect 48357 33108 48611 33164
rect 48357 33074 48391 33108
rect 48425 33074 48544 33108
rect 48578 33074 48611 33108
rect 48357 33018 48611 33074
rect 48357 32984 48391 33018
rect 48425 32984 48544 33018
rect 48578 32984 48611 33018
rect 48357 32928 48611 32984
rect 48357 32894 48391 32928
rect 48425 32894 48544 32928
rect 48578 32894 48611 32928
rect 48357 32838 48611 32894
rect 48357 32804 48391 32838
rect 48425 32804 48544 32838
rect 48578 32804 48611 32838
rect 48357 32748 48611 32804
rect 48357 32714 48391 32748
rect 48425 32714 48544 32748
rect 48578 32714 48611 32748
rect 48357 32658 48611 32714
rect 48357 32624 48391 32658
rect 48425 32624 48544 32658
rect 48578 32624 48611 32658
rect 48357 32568 48611 32624
rect 48357 32534 48391 32568
rect 48425 32534 48544 32568
rect 48578 32534 48611 32568
rect 47017 32444 47051 32478
rect 47085 32444 47204 32478
rect 47238 32444 47271 32478
rect 47017 32429 47271 32444
rect 48357 32478 48611 32534
rect 49697 33434 49731 33468
rect 49765 33434 49884 33468
rect 49918 33434 49951 33468
rect 51037 33468 51291 33515
rect 49697 33378 49951 33434
rect 49697 33344 49731 33378
rect 49765 33344 49884 33378
rect 49918 33344 49951 33378
rect 49697 33288 49951 33344
rect 49697 33254 49731 33288
rect 49765 33254 49884 33288
rect 49918 33254 49951 33288
rect 49697 33198 49951 33254
rect 49697 33164 49731 33198
rect 49765 33164 49884 33198
rect 49918 33164 49951 33198
rect 49697 33108 49951 33164
rect 49697 33074 49731 33108
rect 49765 33074 49884 33108
rect 49918 33074 49951 33108
rect 49697 33018 49951 33074
rect 49697 32984 49731 33018
rect 49765 32984 49884 33018
rect 49918 32984 49951 33018
rect 49697 32928 49951 32984
rect 49697 32894 49731 32928
rect 49765 32894 49884 32928
rect 49918 32894 49951 32928
rect 49697 32838 49951 32894
rect 49697 32804 49731 32838
rect 49765 32804 49884 32838
rect 49918 32804 49951 32838
rect 49697 32748 49951 32804
rect 49697 32714 49731 32748
rect 49765 32714 49884 32748
rect 49918 32714 49951 32748
rect 49697 32658 49951 32714
rect 49697 32624 49731 32658
rect 49765 32624 49884 32658
rect 49918 32624 49951 32658
rect 49697 32568 49951 32624
rect 49697 32534 49731 32568
rect 49765 32534 49884 32568
rect 49918 32534 49951 32568
rect 48357 32444 48391 32478
rect 48425 32444 48544 32478
rect 48578 32444 48611 32478
rect 48357 32429 48611 32444
rect 49697 32478 49951 32534
rect 51037 33434 51071 33468
rect 51105 33434 51224 33468
rect 51258 33434 51291 33468
rect 52377 33468 52478 33515
rect 51037 33378 51291 33434
rect 51037 33344 51071 33378
rect 51105 33344 51224 33378
rect 51258 33344 51291 33378
rect 51037 33288 51291 33344
rect 51037 33254 51071 33288
rect 51105 33254 51224 33288
rect 51258 33254 51291 33288
rect 51037 33198 51291 33254
rect 51037 33164 51071 33198
rect 51105 33164 51224 33198
rect 51258 33164 51291 33198
rect 51037 33108 51291 33164
rect 51037 33074 51071 33108
rect 51105 33074 51224 33108
rect 51258 33074 51291 33108
rect 51037 33018 51291 33074
rect 51037 32984 51071 33018
rect 51105 32984 51224 33018
rect 51258 32984 51291 33018
rect 51037 32928 51291 32984
rect 51037 32894 51071 32928
rect 51105 32894 51224 32928
rect 51258 32894 51291 32928
rect 51037 32838 51291 32894
rect 51037 32804 51071 32838
rect 51105 32804 51224 32838
rect 51258 32804 51291 32838
rect 51037 32748 51291 32804
rect 51037 32714 51071 32748
rect 51105 32714 51224 32748
rect 51258 32714 51291 32748
rect 51037 32658 51291 32714
rect 51037 32624 51071 32658
rect 51105 32624 51224 32658
rect 51258 32624 51291 32658
rect 51037 32568 51291 32624
rect 51037 32534 51071 32568
rect 51105 32534 51224 32568
rect 51258 32534 51291 32568
rect 49697 32444 49731 32478
rect 49765 32444 49884 32478
rect 49918 32444 49951 32478
rect 49697 32429 49951 32444
rect 51037 32478 51291 32534
rect 52377 33434 52411 33468
rect 52445 33434 52478 33468
rect 52377 33378 52478 33434
rect 52377 33344 52411 33378
rect 52445 33344 52478 33378
rect 52377 33288 52478 33344
rect 52377 33254 52411 33288
rect 52445 33254 52478 33288
rect 52377 33198 52478 33254
rect 52377 33164 52411 33198
rect 52445 33164 52478 33198
rect 52377 33108 52478 33164
rect 52377 33074 52411 33108
rect 52445 33074 52478 33108
rect 52377 33018 52478 33074
rect 52377 32984 52411 33018
rect 52445 32984 52478 33018
rect 52377 32928 52478 32984
rect 52377 32894 52411 32928
rect 52445 32894 52478 32928
rect 52377 32838 52478 32894
rect 52377 32804 52411 32838
rect 52445 32804 52478 32838
rect 52377 32748 52478 32804
rect 52377 32714 52411 32748
rect 52445 32714 52478 32748
rect 52377 32658 52478 32714
rect 52377 32624 52411 32658
rect 52445 32624 52478 32658
rect 52377 32568 52478 32624
rect 52377 32534 52411 32568
rect 52445 32534 52478 32568
rect 51037 32444 51071 32478
rect 51105 32444 51224 32478
rect 51258 32444 51291 32478
rect 51037 32429 51291 32444
rect 52377 32478 52478 32534
rect 52377 32444 52411 32478
rect 52445 32444 52478 32478
rect 52377 32429 52478 32444
rect 41810 32394 52478 32429
rect 41810 32360 41940 32394
rect 41974 32360 42030 32394
rect 42064 32360 42120 32394
rect 42154 32360 42210 32394
rect 42244 32360 42300 32394
rect 42334 32360 42390 32394
rect 42424 32360 42480 32394
rect 42514 32360 42570 32394
rect 42604 32360 42660 32394
rect 42694 32360 42750 32394
rect 42784 32360 42840 32394
rect 42874 32360 42930 32394
rect 42964 32360 43280 32394
rect 43314 32360 43370 32394
rect 43404 32360 43460 32394
rect 43494 32360 43550 32394
rect 43584 32360 43640 32394
rect 43674 32360 43730 32394
rect 43764 32360 43820 32394
rect 43854 32360 43910 32394
rect 43944 32360 44000 32394
rect 44034 32360 44090 32394
rect 44124 32360 44180 32394
rect 44214 32360 44270 32394
rect 44304 32360 44620 32394
rect 44654 32360 44710 32394
rect 44744 32360 44800 32394
rect 44834 32360 44890 32394
rect 44924 32360 44980 32394
rect 45014 32360 45070 32394
rect 45104 32360 45160 32394
rect 45194 32360 45250 32394
rect 45284 32360 45340 32394
rect 45374 32360 45430 32394
rect 45464 32360 45520 32394
rect 45554 32360 45610 32394
rect 45644 32360 45960 32394
rect 45994 32360 46050 32394
rect 46084 32360 46140 32394
rect 46174 32360 46230 32394
rect 46264 32360 46320 32394
rect 46354 32360 46410 32394
rect 46444 32360 46500 32394
rect 46534 32360 46590 32394
rect 46624 32360 46680 32394
rect 46714 32360 46770 32394
rect 46804 32360 46860 32394
rect 46894 32360 46950 32394
rect 46984 32360 47300 32394
rect 47334 32360 47390 32394
rect 47424 32360 47480 32394
rect 47514 32360 47570 32394
rect 47604 32360 47660 32394
rect 47694 32360 47750 32394
rect 47784 32360 47840 32394
rect 47874 32360 47930 32394
rect 47964 32360 48020 32394
rect 48054 32360 48110 32394
rect 48144 32360 48200 32394
rect 48234 32360 48290 32394
rect 48324 32360 48640 32394
rect 48674 32360 48730 32394
rect 48764 32360 48820 32394
rect 48854 32360 48910 32394
rect 48944 32360 49000 32394
rect 49034 32360 49090 32394
rect 49124 32360 49180 32394
rect 49214 32360 49270 32394
rect 49304 32360 49360 32394
rect 49394 32360 49450 32394
rect 49484 32360 49540 32394
rect 49574 32360 49630 32394
rect 49664 32360 49980 32394
rect 50014 32360 50070 32394
rect 50104 32360 50160 32394
rect 50194 32360 50250 32394
rect 50284 32360 50340 32394
rect 50374 32360 50430 32394
rect 50464 32360 50520 32394
rect 50554 32360 50610 32394
rect 50644 32360 50700 32394
rect 50734 32360 50790 32394
rect 50824 32360 50880 32394
rect 50914 32360 50970 32394
rect 51004 32360 51320 32394
rect 51354 32360 51410 32394
rect 51444 32360 51500 32394
rect 51534 32360 51590 32394
rect 51624 32360 51680 32394
rect 51714 32360 51770 32394
rect 51804 32360 51860 32394
rect 51894 32360 51950 32394
rect 51984 32360 52040 32394
rect 52074 32360 52130 32394
rect 52164 32360 52220 32394
rect 52254 32360 52310 32394
rect 52344 32360 52478 32394
rect 41810 32328 52478 32360
rect 17432 29203 18048 29242
rect 17432 29101 17519 29203
rect 17961 29101 18048 29203
rect 17432 29062 18048 29101
rect 20176 29203 20792 29242
rect 20176 29101 20263 29203
rect 20705 29101 20792 29203
rect 20176 29062 20792 29101
rect 22920 29203 23536 29242
rect 22920 29101 23007 29203
rect 23449 29101 23536 29203
rect 22920 29062 23536 29101
rect 28114 29203 28730 29242
rect 28114 29101 28201 29203
rect 28643 29101 28730 29203
rect 28114 29062 28730 29101
rect 41810 29821 52478 29856
rect 41810 29798 41940 29821
rect 41810 29764 41844 29798
rect 41878 29787 41940 29798
rect 41974 29787 42030 29821
rect 42064 29787 42120 29821
rect 42154 29787 42210 29821
rect 42244 29787 42300 29821
rect 42334 29787 42390 29821
rect 42424 29787 42480 29821
rect 42514 29787 42570 29821
rect 42604 29787 42660 29821
rect 42694 29787 42750 29821
rect 42784 29787 42840 29821
rect 42874 29787 42930 29821
rect 42964 29798 43280 29821
rect 42964 29787 43031 29798
rect 41878 29764 43031 29787
rect 43065 29764 43184 29798
rect 43218 29787 43280 29798
rect 43314 29787 43370 29821
rect 43404 29787 43460 29821
rect 43494 29787 43550 29821
rect 43584 29787 43640 29821
rect 43674 29787 43730 29821
rect 43764 29787 43820 29821
rect 43854 29787 43910 29821
rect 43944 29787 44000 29821
rect 44034 29787 44090 29821
rect 44124 29787 44180 29821
rect 44214 29787 44270 29821
rect 44304 29798 44620 29821
rect 44304 29787 44371 29798
rect 43218 29764 44371 29787
rect 44405 29764 44524 29798
rect 44558 29787 44620 29798
rect 44654 29787 44710 29821
rect 44744 29787 44800 29821
rect 44834 29787 44890 29821
rect 44924 29787 44980 29821
rect 45014 29787 45070 29821
rect 45104 29787 45160 29821
rect 45194 29787 45250 29821
rect 45284 29787 45340 29821
rect 45374 29787 45430 29821
rect 45464 29787 45520 29821
rect 45554 29787 45610 29821
rect 45644 29798 45960 29821
rect 45644 29787 45711 29798
rect 44558 29764 45711 29787
rect 45745 29764 45864 29798
rect 45898 29787 45960 29798
rect 45994 29787 46050 29821
rect 46084 29787 46140 29821
rect 46174 29787 46230 29821
rect 46264 29787 46320 29821
rect 46354 29787 46410 29821
rect 46444 29787 46500 29821
rect 46534 29787 46590 29821
rect 46624 29787 46680 29821
rect 46714 29787 46770 29821
rect 46804 29787 46860 29821
rect 46894 29787 46950 29821
rect 46984 29798 47300 29821
rect 46984 29787 47051 29798
rect 45898 29764 47051 29787
rect 47085 29764 47204 29798
rect 47238 29787 47300 29798
rect 47334 29787 47390 29821
rect 47424 29787 47480 29821
rect 47514 29787 47570 29821
rect 47604 29787 47660 29821
rect 47694 29787 47750 29821
rect 47784 29787 47840 29821
rect 47874 29787 47930 29821
rect 47964 29787 48020 29821
rect 48054 29787 48110 29821
rect 48144 29787 48200 29821
rect 48234 29787 48290 29821
rect 48324 29798 48640 29821
rect 48324 29787 48391 29798
rect 47238 29764 48391 29787
rect 48425 29764 48544 29798
rect 48578 29787 48640 29798
rect 48674 29787 48730 29821
rect 48764 29787 48820 29821
rect 48854 29787 48910 29821
rect 48944 29787 49000 29821
rect 49034 29787 49090 29821
rect 49124 29787 49180 29821
rect 49214 29787 49270 29821
rect 49304 29787 49360 29821
rect 49394 29787 49450 29821
rect 49484 29787 49540 29821
rect 49574 29787 49630 29821
rect 49664 29798 49980 29821
rect 49664 29787 49731 29798
rect 48578 29764 49731 29787
rect 49765 29764 49884 29798
rect 49918 29787 49980 29798
rect 50014 29787 50070 29821
rect 50104 29787 50160 29821
rect 50194 29787 50250 29821
rect 50284 29787 50340 29821
rect 50374 29787 50430 29821
rect 50464 29787 50520 29821
rect 50554 29787 50610 29821
rect 50644 29787 50700 29821
rect 50734 29787 50790 29821
rect 50824 29787 50880 29821
rect 50914 29787 50970 29821
rect 51004 29798 51320 29821
rect 51004 29787 51071 29798
rect 49918 29764 51071 29787
rect 51105 29764 51224 29798
rect 51258 29787 51320 29798
rect 51354 29787 51410 29821
rect 51444 29787 51500 29821
rect 51534 29787 51590 29821
rect 51624 29787 51680 29821
rect 51714 29787 51770 29821
rect 51804 29787 51860 29821
rect 51894 29787 51950 29821
rect 51984 29787 52040 29821
rect 52074 29787 52130 29821
rect 52164 29787 52220 29821
rect 52254 29787 52310 29821
rect 52344 29798 52478 29821
rect 52344 29787 52411 29798
rect 51258 29764 52411 29787
rect 52445 29764 52478 29798
rect 41810 29755 52478 29764
rect 41810 29708 41911 29755
rect 41810 29674 41844 29708
rect 41878 29674 41911 29708
rect 42997 29708 43251 29755
rect 41810 29618 41911 29674
rect 41810 29584 41844 29618
rect 41878 29584 41911 29618
rect 41810 29528 41911 29584
rect 41810 29494 41844 29528
rect 41878 29494 41911 29528
rect 41810 29438 41911 29494
rect 41810 29404 41844 29438
rect 41878 29404 41911 29438
rect 41810 29348 41911 29404
rect 41810 29314 41844 29348
rect 41878 29314 41911 29348
rect 41810 29258 41911 29314
rect 41810 29224 41844 29258
rect 41878 29224 41911 29258
rect 41810 29168 41911 29224
rect 41810 29134 41844 29168
rect 41878 29134 41911 29168
rect 41810 29078 41911 29134
rect 41810 29044 41844 29078
rect 41878 29044 41911 29078
rect 41810 28988 41911 29044
rect 41810 28954 41844 28988
rect 41878 28954 41911 28988
rect 41810 28898 41911 28954
rect 41810 28864 41844 28898
rect 41878 28864 41911 28898
rect 41810 28808 41911 28864
rect 41810 28774 41844 28808
rect 41878 28774 41911 28808
rect 41810 28718 41911 28774
rect 42997 29674 43031 29708
rect 43065 29674 43184 29708
rect 43218 29674 43251 29708
rect 44337 29708 44591 29755
rect 42997 29618 43251 29674
rect 42997 29584 43031 29618
rect 43065 29584 43184 29618
rect 43218 29584 43251 29618
rect 42997 29528 43251 29584
rect 42997 29494 43031 29528
rect 43065 29494 43184 29528
rect 43218 29494 43251 29528
rect 42997 29438 43251 29494
rect 42997 29404 43031 29438
rect 43065 29404 43184 29438
rect 43218 29404 43251 29438
rect 42997 29348 43251 29404
rect 42997 29314 43031 29348
rect 43065 29314 43184 29348
rect 43218 29314 43251 29348
rect 42997 29258 43251 29314
rect 42997 29224 43031 29258
rect 43065 29224 43184 29258
rect 43218 29224 43251 29258
rect 42997 29168 43251 29224
rect 42997 29134 43031 29168
rect 43065 29134 43184 29168
rect 43218 29134 43251 29168
rect 42997 29078 43251 29134
rect 42997 29044 43031 29078
rect 43065 29044 43184 29078
rect 43218 29044 43251 29078
rect 42997 28988 43251 29044
rect 42997 28954 43031 28988
rect 43065 28954 43184 28988
rect 43218 28954 43251 28988
rect 42997 28898 43251 28954
rect 42997 28864 43031 28898
rect 43065 28864 43184 28898
rect 43218 28864 43251 28898
rect 42997 28808 43251 28864
rect 42997 28774 43031 28808
rect 43065 28774 43184 28808
rect 43218 28774 43251 28808
rect 41810 28684 41844 28718
rect 41878 28684 41911 28718
rect 41810 28669 41911 28684
rect 42997 28718 43251 28774
rect 44337 29674 44371 29708
rect 44405 29674 44524 29708
rect 44558 29674 44591 29708
rect 45677 29708 45931 29755
rect 44337 29618 44591 29674
rect 44337 29584 44371 29618
rect 44405 29584 44524 29618
rect 44558 29584 44591 29618
rect 44337 29528 44591 29584
rect 44337 29494 44371 29528
rect 44405 29494 44524 29528
rect 44558 29494 44591 29528
rect 44337 29438 44591 29494
rect 44337 29404 44371 29438
rect 44405 29404 44524 29438
rect 44558 29404 44591 29438
rect 44337 29348 44591 29404
rect 44337 29314 44371 29348
rect 44405 29314 44524 29348
rect 44558 29314 44591 29348
rect 44337 29258 44591 29314
rect 44337 29224 44371 29258
rect 44405 29224 44524 29258
rect 44558 29224 44591 29258
rect 44337 29168 44591 29224
rect 44337 29134 44371 29168
rect 44405 29134 44524 29168
rect 44558 29134 44591 29168
rect 44337 29078 44591 29134
rect 44337 29044 44371 29078
rect 44405 29044 44524 29078
rect 44558 29044 44591 29078
rect 44337 28988 44591 29044
rect 44337 28954 44371 28988
rect 44405 28954 44524 28988
rect 44558 28954 44591 28988
rect 44337 28898 44591 28954
rect 44337 28864 44371 28898
rect 44405 28864 44524 28898
rect 44558 28864 44591 28898
rect 44337 28808 44591 28864
rect 44337 28774 44371 28808
rect 44405 28774 44524 28808
rect 44558 28774 44591 28808
rect 42997 28684 43031 28718
rect 43065 28684 43184 28718
rect 43218 28684 43251 28718
rect 42997 28669 43251 28684
rect 44337 28718 44591 28774
rect 45677 29674 45711 29708
rect 45745 29674 45864 29708
rect 45898 29674 45931 29708
rect 47017 29708 47271 29755
rect 45677 29618 45931 29674
rect 45677 29584 45711 29618
rect 45745 29584 45864 29618
rect 45898 29584 45931 29618
rect 45677 29528 45931 29584
rect 45677 29494 45711 29528
rect 45745 29494 45864 29528
rect 45898 29494 45931 29528
rect 45677 29438 45931 29494
rect 45677 29404 45711 29438
rect 45745 29404 45864 29438
rect 45898 29404 45931 29438
rect 45677 29348 45931 29404
rect 45677 29314 45711 29348
rect 45745 29314 45864 29348
rect 45898 29314 45931 29348
rect 45677 29258 45931 29314
rect 45677 29224 45711 29258
rect 45745 29224 45864 29258
rect 45898 29224 45931 29258
rect 45677 29168 45931 29224
rect 45677 29134 45711 29168
rect 45745 29134 45864 29168
rect 45898 29134 45931 29168
rect 45677 29078 45931 29134
rect 45677 29044 45711 29078
rect 45745 29044 45864 29078
rect 45898 29044 45931 29078
rect 45677 28988 45931 29044
rect 45677 28954 45711 28988
rect 45745 28954 45864 28988
rect 45898 28954 45931 28988
rect 45677 28898 45931 28954
rect 45677 28864 45711 28898
rect 45745 28864 45864 28898
rect 45898 28864 45931 28898
rect 45677 28808 45931 28864
rect 45677 28774 45711 28808
rect 45745 28774 45864 28808
rect 45898 28774 45931 28808
rect 44337 28684 44371 28718
rect 44405 28684 44524 28718
rect 44558 28684 44591 28718
rect 44337 28669 44591 28684
rect 45677 28718 45931 28774
rect 47017 29674 47051 29708
rect 47085 29674 47204 29708
rect 47238 29674 47271 29708
rect 48357 29708 48611 29755
rect 47017 29618 47271 29674
rect 47017 29584 47051 29618
rect 47085 29584 47204 29618
rect 47238 29584 47271 29618
rect 47017 29528 47271 29584
rect 47017 29494 47051 29528
rect 47085 29494 47204 29528
rect 47238 29494 47271 29528
rect 47017 29438 47271 29494
rect 47017 29404 47051 29438
rect 47085 29404 47204 29438
rect 47238 29404 47271 29438
rect 47017 29348 47271 29404
rect 47017 29314 47051 29348
rect 47085 29314 47204 29348
rect 47238 29314 47271 29348
rect 47017 29258 47271 29314
rect 47017 29224 47051 29258
rect 47085 29224 47204 29258
rect 47238 29224 47271 29258
rect 47017 29168 47271 29224
rect 47017 29134 47051 29168
rect 47085 29134 47204 29168
rect 47238 29134 47271 29168
rect 47017 29078 47271 29134
rect 47017 29044 47051 29078
rect 47085 29044 47204 29078
rect 47238 29044 47271 29078
rect 47017 28988 47271 29044
rect 47017 28954 47051 28988
rect 47085 28954 47204 28988
rect 47238 28954 47271 28988
rect 47017 28898 47271 28954
rect 47017 28864 47051 28898
rect 47085 28864 47204 28898
rect 47238 28864 47271 28898
rect 47017 28808 47271 28864
rect 47017 28774 47051 28808
rect 47085 28774 47204 28808
rect 47238 28774 47271 28808
rect 45677 28684 45711 28718
rect 45745 28684 45864 28718
rect 45898 28684 45931 28718
rect 45677 28669 45931 28684
rect 47017 28718 47271 28774
rect 48357 29674 48391 29708
rect 48425 29674 48544 29708
rect 48578 29674 48611 29708
rect 49697 29708 49951 29755
rect 48357 29618 48611 29674
rect 48357 29584 48391 29618
rect 48425 29584 48544 29618
rect 48578 29584 48611 29618
rect 48357 29528 48611 29584
rect 48357 29494 48391 29528
rect 48425 29494 48544 29528
rect 48578 29494 48611 29528
rect 48357 29438 48611 29494
rect 48357 29404 48391 29438
rect 48425 29404 48544 29438
rect 48578 29404 48611 29438
rect 48357 29348 48611 29404
rect 48357 29314 48391 29348
rect 48425 29314 48544 29348
rect 48578 29314 48611 29348
rect 48357 29258 48611 29314
rect 48357 29224 48391 29258
rect 48425 29224 48544 29258
rect 48578 29224 48611 29258
rect 48357 29168 48611 29224
rect 48357 29134 48391 29168
rect 48425 29134 48544 29168
rect 48578 29134 48611 29168
rect 48357 29078 48611 29134
rect 48357 29044 48391 29078
rect 48425 29044 48544 29078
rect 48578 29044 48611 29078
rect 48357 28988 48611 29044
rect 48357 28954 48391 28988
rect 48425 28954 48544 28988
rect 48578 28954 48611 28988
rect 48357 28898 48611 28954
rect 48357 28864 48391 28898
rect 48425 28864 48544 28898
rect 48578 28864 48611 28898
rect 48357 28808 48611 28864
rect 48357 28774 48391 28808
rect 48425 28774 48544 28808
rect 48578 28774 48611 28808
rect 47017 28684 47051 28718
rect 47085 28684 47204 28718
rect 47238 28684 47271 28718
rect 47017 28669 47271 28684
rect 48357 28718 48611 28774
rect 49697 29674 49731 29708
rect 49765 29674 49884 29708
rect 49918 29674 49951 29708
rect 51037 29708 51291 29755
rect 49697 29618 49951 29674
rect 49697 29584 49731 29618
rect 49765 29584 49884 29618
rect 49918 29584 49951 29618
rect 49697 29528 49951 29584
rect 49697 29494 49731 29528
rect 49765 29494 49884 29528
rect 49918 29494 49951 29528
rect 49697 29438 49951 29494
rect 49697 29404 49731 29438
rect 49765 29404 49884 29438
rect 49918 29404 49951 29438
rect 49697 29348 49951 29404
rect 49697 29314 49731 29348
rect 49765 29314 49884 29348
rect 49918 29314 49951 29348
rect 49697 29258 49951 29314
rect 49697 29224 49731 29258
rect 49765 29224 49884 29258
rect 49918 29224 49951 29258
rect 49697 29168 49951 29224
rect 49697 29134 49731 29168
rect 49765 29134 49884 29168
rect 49918 29134 49951 29168
rect 49697 29078 49951 29134
rect 49697 29044 49731 29078
rect 49765 29044 49884 29078
rect 49918 29044 49951 29078
rect 49697 28988 49951 29044
rect 49697 28954 49731 28988
rect 49765 28954 49884 28988
rect 49918 28954 49951 28988
rect 49697 28898 49951 28954
rect 49697 28864 49731 28898
rect 49765 28864 49884 28898
rect 49918 28864 49951 28898
rect 49697 28808 49951 28864
rect 49697 28774 49731 28808
rect 49765 28774 49884 28808
rect 49918 28774 49951 28808
rect 48357 28684 48391 28718
rect 48425 28684 48544 28718
rect 48578 28684 48611 28718
rect 48357 28669 48611 28684
rect 49697 28718 49951 28774
rect 51037 29674 51071 29708
rect 51105 29674 51224 29708
rect 51258 29674 51291 29708
rect 52377 29708 52478 29755
rect 51037 29618 51291 29674
rect 51037 29584 51071 29618
rect 51105 29584 51224 29618
rect 51258 29584 51291 29618
rect 51037 29528 51291 29584
rect 51037 29494 51071 29528
rect 51105 29494 51224 29528
rect 51258 29494 51291 29528
rect 51037 29438 51291 29494
rect 51037 29404 51071 29438
rect 51105 29404 51224 29438
rect 51258 29404 51291 29438
rect 51037 29348 51291 29404
rect 51037 29314 51071 29348
rect 51105 29314 51224 29348
rect 51258 29314 51291 29348
rect 51037 29258 51291 29314
rect 51037 29224 51071 29258
rect 51105 29224 51224 29258
rect 51258 29224 51291 29258
rect 51037 29168 51291 29224
rect 51037 29134 51071 29168
rect 51105 29134 51224 29168
rect 51258 29134 51291 29168
rect 51037 29078 51291 29134
rect 51037 29044 51071 29078
rect 51105 29044 51224 29078
rect 51258 29044 51291 29078
rect 51037 28988 51291 29044
rect 51037 28954 51071 28988
rect 51105 28954 51224 28988
rect 51258 28954 51291 28988
rect 51037 28898 51291 28954
rect 51037 28864 51071 28898
rect 51105 28864 51224 28898
rect 51258 28864 51291 28898
rect 51037 28808 51291 28864
rect 51037 28774 51071 28808
rect 51105 28774 51224 28808
rect 51258 28774 51291 28808
rect 49697 28684 49731 28718
rect 49765 28684 49884 28718
rect 49918 28684 49951 28718
rect 49697 28669 49951 28684
rect 51037 28718 51291 28774
rect 52377 29674 52411 29708
rect 52445 29674 52478 29708
rect 52377 29618 52478 29674
rect 52377 29584 52411 29618
rect 52445 29584 52478 29618
rect 52377 29528 52478 29584
rect 52377 29494 52411 29528
rect 52445 29494 52478 29528
rect 52377 29438 52478 29494
rect 52377 29404 52411 29438
rect 52445 29404 52478 29438
rect 52377 29348 52478 29404
rect 52377 29314 52411 29348
rect 52445 29314 52478 29348
rect 52377 29258 52478 29314
rect 52377 29224 52411 29258
rect 52445 29224 52478 29258
rect 52377 29168 52478 29224
rect 52377 29134 52411 29168
rect 52445 29134 52478 29168
rect 52377 29078 52478 29134
rect 52377 29044 52411 29078
rect 52445 29044 52478 29078
rect 52377 28988 52478 29044
rect 52377 28954 52411 28988
rect 52445 28954 52478 28988
rect 52377 28898 52478 28954
rect 52377 28864 52411 28898
rect 52445 28864 52478 28898
rect 52377 28808 52478 28864
rect 52377 28774 52411 28808
rect 52445 28774 52478 28808
rect 51037 28684 51071 28718
rect 51105 28684 51224 28718
rect 51258 28684 51291 28718
rect 51037 28669 51291 28684
rect 52377 28718 52478 28774
rect 52377 28684 52411 28718
rect 52445 28684 52478 28718
rect 52377 28669 52478 28684
rect 41810 28634 52478 28669
rect 41810 28600 41940 28634
rect 41974 28600 42030 28634
rect 42064 28600 42120 28634
rect 42154 28600 42210 28634
rect 42244 28600 42300 28634
rect 42334 28600 42390 28634
rect 42424 28600 42480 28634
rect 42514 28600 42570 28634
rect 42604 28600 42660 28634
rect 42694 28600 42750 28634
rect 42784 28600 42840 28634
rect 42874 28600 42930 28634
rect 42964 28600 43280 28634
rect 43314 28600 43370 28634
rect 43404 28600 43460 28634
rect 43494 28600 43550 28634
rect 43584 28600 43640 28634
rect 43674 28600 43730 28634
rect 43764 28600 43820 28634
rect 43854 28600 43910 28634
rect 43944 28600 44000 28634
rect 44034 28600 44090 28634
rect 44124 28600 44180 28634
rect 44214 28600 44270 28634
rect 44304 28600 44620 28634
rect 44654 28600 44710 28634
rect 44744 28600 44800 28634
rect 44834 28600 44890 28634
rect 44924 28600 44980 28634
rect 45014 28600 45070 28634
rect 45104 28600 45160 28634
rect 45194 28600 45250 28634
rect 45284 28600 45340 28634
rect 45374 28600 45430 28634
rect 45464 28600 45520 28634
rect 45554 28600 45610 28634
rect 45644 28600 45960 28634
rect 45994 28600 46050 28634
rect 46084 28600 46140 28634
rect 46174 28600 46230 28634
rect 46264 28600 46320 28634
rect 46354 28600 46410 28634
rect 46444 28600 46500 28634
rect 46534 28600 46590 28634
rect 46624 28600 46680 28634
rect 46714 28600 46770 28634
rect 46804 28600 46860 28634
rect 46894 28600 46950 28634
rect 46984 28600 47300 28634
rect 47334 28600 47390 28634
rect 47424 28600 47480 28634
rect 47514 28600 47570 28634
rect 47604 28600 47660 28634
rect 47694 28600 47750 28634
rect 47784 28600 47840 28634
rect 47874 28600 47930 28634
rect 47964 28600 48020 28634
rect 48054 28600 48110 28634
rect 48144 28600 48200 28634
rect 48234 28600 48290 28634
rect 48324 28600 48640 28634
rect 48674 28600 48730 28634
rect 48764 28600 48820 28634
rect 48854 28600 48910 28634
rect 48944 28600 49000 28634
rect 49034 28600 49090 28634
rect 49124 28600 49180 28634
rect 49214 28600 49270 28634
rect 49304 28600 49360 28634
rect 49394 28600 49450 28634
rect 49484 28600 49540 28634
rect 49574 28600 49630 28634
rect 49664 28600 49980 28634
rect 50014 28600 50070 28634
rect 50104 28600 50160 28634
rect 50194 28600 50250 28634
rect 50284 28600 50340 28634
rect 50374 28600 50430 28634
rect 50464 28600 50520 28634
rect 50554 28600 50610 28634
rect 50644 28600 50700 28634
rect 50734 28600 50790 28634
rect 50824 28600 50880 28634
rect 50914 28600 50970 28634
rect 51004 28600 51320 28634
rect 51354 28600 51410 28634
rect 51444 28600 51500 28634
rect 51534 28600 51590 28634
rect 51624 28600 51680 28634
rect 51714 28600 51770 28634
rect 51804 28600 51860 28634
rect 51894 28600 51950 28634
rect 51984 28600 52040 28634
rect 52074 28600 52130 28634
rect 52164 28600 52220 28634
rect 52254 28600 52310 28634
rect 52344 28600 52478 28634
rect 41810 28568 52478 28600
rect 23312 25443 23928 25482
rect 23312 25341 23399 25443
rect 23841 25341 23928 25443
rect 23312 25302 23928 25341
rect 38306 25443 38922 25482
rect 38306 25341 38393 25443
rect 38835 25341 38922 25443
rect 38306 25302 38922 25341
rect 41050 25443 41666 25482
rect 41050 25341 41137 25443
rect 41579 25341 41666 25443
rect 41050 25302 41666 25341
rect 43794 25443 44410 25482
rect 43794 25341 43881 25443
rect 44323 25341 44410 25443
rect 43794 25302 44410 25341
rect 46538 25443 47154 25482
rect 46538 25341 46625 25443
rect 47067 25341 47154 25443
rect 46538 25302 47154 25341
rect 49282 25443 49898 25482
rect 49282 25341 49369 25443
rect 49811 25341 49898 25443
rect 49282 25302 49898 25341
rect 25358 24669 25398 24712
rect 25358 24635 25361 24669
rect 25395 24635 25398 24669
rect 25358 24592 25398 24635
rect 26418 24639 26538 24642
rect 26418 24605 26463 24639
rect 26497 24605 26538 24639
rect 26418 24592 26538 24605
rect 27718 24639 27838 24642
rect 27718 24605 27763 24639
rect 27797 24605 27838 24639
rect 27718 24592 27838 24605
rect 24782 21683 25398 21722
rect 24782 21581 24869 21683
rect 25311 21581 25398 21683
rect 24782 21542 25398 21581
rect 28114 21683 28730 21722
rect 28114 21581 28201 21683
rect 28643 21581 28730 21683
rect 28114 21542 28730 21581
rect 30858 21683 31474 21722
rect 30858 21581 30945 21683
rect 31387 21581 31474 21683
rect 30858 21542 31474 21581
rect 34092 21683 34708 21722
rect 34092 21581 34179 21683
rect 34621 21581 34708 21683
rect 34092 21542 34708 21581
rect 38306 21683 38922 21722
rect 38306 21581 38393 21683
rect 38835 21581 38922 21683
rect 38306 21542 38922 21581
rect 41050 21683 41666 21722
rect 41050 21581 41137 21683
rect 41579 21581 41666 21683
rect 41050 21542 41666 21581
rect 49282 21683 49898 21722
rect 49282 21581 49369 21683
rect 49811 21581 49898 21683
rect 49282 21542 49898 21581
rect 44774 14163 45390 14202
rect 44774 14061 44861 14163
rect 45303 14061 45390 14163
rect 44774 14022 45390 14061
rect 47518 14163 48134 14202
rect 47518 14061 47605 14163
rect 48047 14061 48134 14163
rect 47518 14022 48134 14061
rect 50262 14163 50878 14202
rect 50262 14061 50349 14163
rect 50791 14061 50878 14163
rect 50262 14022 50878 14061
rect 44676 10403 45292 10442
rect 44676 10301 44763 10403
rect 45205 10301 45292 10403
rect 44676 10262 45292 10301
rect 47420 10403 48036 10442
rect 47420 10301 47507 10403
rect 47949 10301 48036 10403
rect 47420 10262 48036 10301
rect 50164 10403 50780 10442
rect 50164 10301 50251 10403
rect 50693 10301 50780 10403
rect 50164 10262 50780 10301
rect 45460 6643 46076 6682
rect 45460 6541 45547 6643
rect 45989 6541 46076 6643
rect 45460 6502 46076 6541
rect 48204 6643 48820 6682
rect 48204 6541 48291 6643
rect 48733 6541 48820 6643
rect 48204 6502 48820 6541
rect 50948 6643 51564 6682
rect 50948 6541 51035 6643
rect 51477 6541 51564 6643
rect 50948 6502 51564 6541
<< nsubdiff >>
rect 25828 48879 25948 48882
rect 24770 48829 24810 48872
rect 25828 48845 25873 48879
rect 25907 48845 25948 48879
rect 25828 48842 25948 48845
rect 27128 48879 27248 48882
rect 27128 48845 27173 48879
rect 27207 48845 27248 48879
rect 27128 48842 27248 48845
rect 28428 48879 28548 48882
rect 28428 48845 28473 48879
rect 28507 48845 28548 48879
rect 28428 48842 28548 48845
rect 29728 48879 29848 48882
rect 29728 48845 29773 48879
rect 29807 48845 29848 48879
rect 29728 48842 29848 48845
rect 31028 48879 31148 48882
rect 31028 48845 31073 48879
rect 31107 48845 31148 48879
rect 31028 48842 31148 48845
rect 32328 48879 32448 48882
rect 32328 48845 32373 48879
rect 32407 48845 32448 48879
rect 32328 48842 32448 48845
rect 33628 48879 33748 48882
rect 33628 48845 33673 48879
rect 33707 48845 33748 48879
rect 33628 48842 33748 48845
rect 34928 48879 35048 48882
rect 34928 48845 34973 48879
rect 35007 48845 35048 48879
rect 34928 48842 35048 48845
rect 36228 48879 36348 48882
rect 36228 48845 36273 48879
rect 36307 48845 36348 48879
rect 36228 48842 36348 48845
rect 37528 48879 37648 48882
rect 37528 48845 37573 48879
rect 37607 48845 37648 48879
rect 37528 48842 37648 48845
rect 38828 48879 38948 48882
rect 38828 48845 38873 48879
rect 38907 48845 38948 48879
rect 38828 48842 38948 48845
rect 40128 48879 40248 48882
rect 40128 48845 40173 48879
rect 40207 48845 40248 48879
rect 40128 48842 40248 48845
rect 41428 48879 41548 48882
rect 41428 48845 41473 48879
rect 41507 48845 41548 48879
rect 41428 48842 41548 48845
rect 42728 48879 42848 48882
rect 42728 48845 42773 48879
rect 42807 48845 42848 48879
rect 42728 48842 42848 48845
rect 44028 48879 44148 48882
rect 44028 48845 44073 48879
rect 44107 48845 44148 48879
rect 44028 48842 44148 48845
rect 45328 48879 45448 48882
rect 45328 48845 45373 48879
rect 45407 48845 45448 48879
rect 45328 48842 45448 48845
rect 46628 48879 46748 48882
rect 46628 48845 46673 48879
rect 46707 48845 46748 48879
rect 46628 48842 46748 48845
rect 47928 48879 48048 48882
rect 47928 48845 47973 48879
rect 48007 48845 48048 48879
rect 47928 48842 48048 48845
rect 49228 48879 49348 48882
rect 49228 48845 49273 48879
rect 49307 48845 49348 48879
rect 49228 48842 49348 48845
rect 50528 48879 50648 48882
rect 50528 48845 50573 48879
rect 50607 48845 50648 48879
rect 50528 48842 50648 48845
rect 24770 48795 24773 48829
rect 24807 48795 24810 48829
rect 24770 48752 24810 48795
rect 16028 45119 16148 45122
rect 14970 45069 15010 45112
rect 16028 45085 16073 45119
rect 16107 45085 16148 45119
rect 16028 45082 16148 45085
rect 17328 45119 17448 45122
rect 17328 45085 17373 45119
rect 17407 45085 17448 45119
rect 17328 45082 17448 45085
rect 18628 45119 18748 45122
rect 18628 45085 18673 45119
rect 18707 45085 18748 45119
rect 18628 45082 18748 45085
rect 19928 45119 20048 45122
rect 19928 45085 19973 45119
rect 20007 45085 20048 45119
rect 19928 45082 20048 45085
rect 21228 45119 21348 45122
rect 21228 45085 21273 45119
rect 21307 45085 21348 45119
rect 21228 45082 21348 45085
rect 22528 45119 22648 45122
rect 22528 45085 22573 45119
rect 22607 45085 22648 45119
rect 22528 45082 22648 45085
rect 23828 45119 23948 45122
rect 23828 45085 23873 45119
rect 23907 45085 23948 45119
rect 23828 45082 23948 45085
rect 25128 45119 25248 45122
rect 25128 45085 25173 45119
rect 25207 45085 25248 45119
rect 25128 45082 25248 45085
rect 26428 45119 26548 45122
rect 26428 45085 26473 45119
rect 26507 45085 26548 45119
rect 26428 45082 26548 45085
rect 27728 45119 27848 45122
rect 27728 45085 27773 45119
rect 27807 45085 27848 45119
rect 27728 45082 27848 45085
rect 29028 45119 29148 45122
rect 29028 45085 29073 45119
rect 29107 45085 29148 45119
rect 29028 45082 29148 45085
rect 30328 45119 30448 45122
rect 30328 45085 30373 45119
rect 30407 45085 30448 45119
rect 30328 45082 30448 45085
rect 31628 45119 31748 45122
rect 31628 45085 31673 45119
rect 31707 45085 31748 45119
rect 31628 45082 31748 45085
rect 32928 45119 33048 45122
rect 32928 45085 32973 45119
rect 33007 45085 33048 45119
rect 32928 45082 33048 45085
rect 34228 45119 34348 45122
rect 34228 45085 34273 45119
rect 34307 45085 34348 45119
rect 34228 45082 34348 45085
rect 35528 45119 35648 45122
rect 35528 45085 35573 45119
rect 35607 45085 35648 45119
rect 35528 45082 35648 45085
rect 36828 45119 36948 45122
rect 36828 45085 36873 45119
rect 36907 45085 36948 45119
rect 36828 45082 36948 45085
rect 38128 45119 38248 45122
rect 38128 45085 38173 45119
rect 38207 45085 38248 45119
rect 38128 45082 38248 45085
rect 39428 45119 39548 45122
rect 39428 45085 39473 45119
rect 39507 45085 39548 45119
rect 39428 45082 39548 45085
rect 40728 45119 40848 45122
rect 40728 45085 40773 45119
rect 40807 45085 40848 45119
rect 40728 45082 40848 45085
rect 14970 45035 14973 45069
rect 15007 45035 15010 45069
rect 14970 44992 15010 45035
rect 43149 44714 44111 44733
rect 43149 44680 43280 44714
rect 43314 44680 43370 44714
rect 43404 44680 43460 44714
rect 43494 44680 43550 44714
rect 43584 44680 43640 44714
rect 43674 44680 43730 44714
rect 43764 44680 43820 44714
rect 43854 44680 43910 44714
rect 43944 44680 44000 44714
rect 44034 44680 44111 44714
rect 43149 44661 44111 44680
rect 43149 44657 43221 44661
rect 43149 44623 43168 44657
rect 43202 44623 43221 44657
rect 43149 44567 43221 44623
rect 44039 44638 44111 44661
rect 44039 44604 44058 44638
rect 44092 44604 44111 44638
rect 43149 44533 43168 44567
rect 43202 44533 43221 44567
rect 43149 44477 43221 44533
rect 43149 44443 43168 44477
rect 43202 44443 43221 44477
rect 43149 44387 43221 44443
rect 43149 44353 43168 44387
rect 43202 44353 43221 44387
rect 43149 44297 43221 44353
rect 43149 44263 43168 44297
rect 43202 44263 43221 44297
rect 43149 44207 43221 44263
rect 43149 44173 43168 44207
rect 43202 44173 43221 44207
rect 43149 44117 43221 44173
rect 43149 44083 43168 44117
rect 43202 44083 43221 44117
rect 43149 44027 43221 44083
rect 43149 43993 43168 44027
rect 43202 43993 43221 44027
rect 43149 43937 43221 43993
rect 43149 43903 43168 43937
rect 43202 43903 43221 43937
rect 44039 44548 44111 44604
rect 44039 44514 44058 44548
rect 44092 44514 44111 44548
rect 44039 44458 44111 44514
rect 44039 44424 44058 44458
rect 44092 44424 44111 44458
rect 44039 44368 44111 44424
rect 44039 44334 44058 44368
rect 44092 44334 44111 44368
rect 44039 44278 44111 44334
rect 44039 44244 44058 44278
rect 44092 44244 44111 44278
rect 44039 44188 44111 44244
rect 44039 44154 44058 44188
rect 44092 44154 44111 44188
rect 44039 44098 44111 44154
rect 44039 44064 44058 44098
rect 44092 44064 44111 44098
rect 44039 44008 44111 44064
rect 44039 43974 44058 44008
rect 44092 43974 44111 44008
rect 44039 43918 44111 43974
rect 43149 43843 43221 43903
rect 44039 43884 44058 43918
rect 44092 43884 44111 43918
rect 44039 43843 44111 43884
rect 43149 43824 44111 43843
rect 43149 43790 43246 43824
rect 43280 43790 43336 43824
rect 43370 43790 43426 43824
rect 43460 43790 43516 43824
rect 43550 43790 43606 43824
rect 43640 43790 43696 43824
rect 43730 43790 43786 43824
rect 43820 43790 43876 43824
rect 43910 43790 43966 43824
rect 44000 43790 44111 43824
rect 43149 43771 44111 43790
rect 44489 44714 45451 44733
rect 44489 44680 44620 44714
rect 44654 44680 44710 44714
rect 44744 44680 44800 44714
rect 44834 44680 44890 44714
rect 44924 44680 44980 44714
rect 45014 44680 45070 44714
rect 45104 44680 45160 44714
rect 45194 44680 45250 44714
rect 45284 44680 45340 44714
rect 45374 44680 45451 44714
rect 44489 44661 45451 44680
rect 44489 44657 44561 44661
rect 44489 44623 44508 44657
rect 44542 44623 44561 44657
rect 44489 44567 44561 44623
rect 45379 44638 45451 44661
rect 45379 44604 45398 44638
rect 45432 44604 45451 44638
rect 44489 44533 44508 44567
rect 44542 44533 44561 44567
rect 44489 44477 44561 44533
rect 44489 44443 44508 44477
rect 44542 44443 44561 44477
rect 44489 44387 44561 44443
rect 44489 44353 44508 44387
rect 44542 44353 44561 44387
rect 44489 44297 44561 44353
rect 44489 44263 44508 44297
rect 44542 44263 44561 44297
rect 44489 44207 44561 44263
rect 44489 44173 44508 44207
rect 44542 44173 44561 44207
rect 44489 44117 44561 44173
rect 44489 44083 44508 44117
rect 44542 44083 44561 44117
rect 44489 44027 44561 44083
rect 44489 43993 44508 44027
rect 44542 43993 44561 44027
rect 44489 43937 44561 43993
rect 44489 43903 44508 43937
rect 44542 43903 44561 43937
rect 45379 44548 45451 44604
rect 45379 44514 45398 44548
rect 45432 44514 45451 44548
rect 45379 44458 45451 44514
rect 45379 44424 45398 44458
rect 45432 44424 45451 44458
rect 45379 44368 45451 44424
rect 45379 44334 45398 44368
rect 45432 44334 45451 44368
rect 45379 44278 45451 44334
rect 45379 44244 45398 44278
rect 45432 44244 45451 44278
rect 45379 44188 45451 44244
rect 45379 44154 45398 44188
rect 45432 44154 45451 44188
rect 45379 44098 45451 44154
rect 45379 44064 45398 44098
rect 45432 44064 45451 44098
rect 45379 44008 45451 44064
rect 45379 43974 45398 44008
rect 45432 43974 45451 44008
rect 45379 43918 45451 43974
rect 44489 43843 44561 43903
rect 45379 43884 45398 43918
rect 45432 43884 45451 43918
rect 45379 43843 45451 43884
rect 44489 43824 45451 43843
rect 44489 43790 44586 43824
rect 44620 43790 44676 43824
rect 44710 43790 44766 43824
rect 44800 43790 44856 43824
rect 44890 43790 44946 43824
rect 44980 43790 45036 43824
rect 45070 43790 45126 43824
rect 45160 43790 45216 43824
rect 45250 43790 45306 43824
rect 45340 43790 45451 43824
rect 44489 43771 45451 43790
rect 45829 44714 46791 44733
rect 45829 44680 45960 44714
rect 45994 44680 46050 44714
rect 46084 44680 46140 44714
rect 46174 44680 46230 44714
rect 46264 44680 46320 44714
rect 46354 44680 46410 44714
rect 46444 44680 46500 44714
rect 46534 44680 46590 44714
rect 46624 44680 46680 44714
rect 46714 44680 46791 44714
rect 45829 44661 46791 44680
rect 45829 44657 45901 44661
rect 45829 44623 45848 44657
rect 45882 44623 45901 44657
rect 45829 44567 45901 44623
rect 46719 44638 46791 44661
rect 46719 44604 46738 44638
rect 46772 44604 46791 44638
rect 45829 44533 45848 44567
rect 45882 44533 45901 44567
rect 45829 44477 45901 44533
rect 45829 44443 45848 44477
rect 45882 44443 45901 44477
rect 45829 44387 45901 44443
rect 45829 44353 45848 44387
rect 45882 44353 45901 44387
rect 45829 44297 45901 44353
rect 45829 44263 45848 44297
rect 45882 44263 45901 44297
rect 45829 44207 45901 44263
rect 45829 44173 45848 44207
rect 45882 44173 45901 44207
rect 45829 44117 45901 44173
rect 45829 44083 45848 44117
rect 45882 44083 45901 44117
rect 45829 44027 45901 44083
rect 45829 43993 45848 44027
rect 45882 43993 45901 44027
rect 45829 43937 45901 43993
rect 45829 43903 45848 43937
rect 45882 43903 45901 43937
rect 46719 44548 46791 44604
rect 46719 44514 46738 44548
rect 46772 44514 46791 44548
rect 46719 44458 46791 44514
rect 46719 44424 46738 44458
rect 46772 44424 46791 44458
rect 46719 44368 46791 44424
rect 46719 44334 46738 44368
rect 46772 44334 46791 44368
rect 46719 44278 46791 44334
rect 46719 44244 46738 44278
rect 46772 44244 46791 44278
rect 46719 44188 46791 44244
rect 46719 44154 46738 44188
rect 46772 44154 46791 44188
rect 46719 44098 46791 44154
rect 46719 44064 46738 44098
rect 46772 44064 46791 44098
rect 46719 44008 46791 44064
rect 46719 43974 46738 44008
rect 46772 43974 46791 44008
rect 46719 43918 46791 43974
rect 45829 43843 45901 43903
rect 46719 43884 46738 43918
rect 46772 43884 46791 43918
rect 46719 43843 46791 43884
rect 45829 43824 46791 43843
rect 45829 43790 45926 43824
rect 45960 43790 46016 43824
rect 46050 43790 46106 43824
rect 46140 43790 46196 43824
rect 46230 43790 46286 43824
rect 46320 43790 46376 43824
rect 46410 43790 46466 43824
rect 46500 43790 46556 43824
rect 46590 43790 46646 43824
rect 46680 43790 46791 43824
rect 45829 43771 46791 43790
rect 47169 44714 48131 44733
rect 47169 44680 47300 44714
rect 47334 44680 47390 44714
rect 47424 44680 47480 44714
rect 47514 44680 47570 44714
rect 47604 44680 47660 44714
rect 47694 44680 47750 44714
rect 47784 44680 47840 44714
rect 47874 44680 47930 44714
rect 47964 44680 48020 44714
rect 48054 44680 48131 44714
rect 47169 44661 48131 44680
rect 47169 44657 47241 44661
rect 47169 44623 47188 44657
rect 47222 44623 47241 44657
rect 47169 44567 47241 44623
rect 48059 44638 48131 44661
rect 48059 44604 48078 44638
rect 48112 44604 48131 44638
rect 47169 44533 47188 44567
rect 47222 44533 47241 44567
rect 47169 44477 47241 44533
rect 47169 44443 47188 44477
rect 47222 44443 47241 44477
rect 47169 44387 47241 44443
rect 47169 44353 47188 44387
rect 47222 44353 47241 44387
rect 47169 44297 47241 44353
rect 47169 44263 47188 44297
rect 47222 44263 47241 44297
rect 47169 44207 47241 44263
rect 47169 44173 47188 44207
rect 47222 44173 47241 44207
rect 47169 44117 47241 44173
rect 47169 44083 47188 44117
rect 47222 44083 47241 44117
rect 47169 44027 47241 44083
rect 47169 43993 47188 44027
rect 47222 43993 47241 44027
rect 47169 43937 47241 43993
rect 47169 43903 47188 43937
rect 47222 43903 47241 43937
rect 48059 44548 48131 44604
rect 48059 44514 48078 44548
rect 48112 44514 48131 44548
rect 48059 44458 48131 44514
rect 48059 44424 48078 44458
rect 48112 44424 48131 44458
rect 48059 44368 48131 44424
rect 48059 44334 48078 44368
rect 48112 44334 48131 44368
rect 48059 44278 48131 44334
rect 48059 44244 48078 44278
rect 48112 44244 48131 44278
rect 48059 44188 48131 44244
rect 48059 44154 48078 44188
rect 48112 44154 48131 44188
rect 48059 44098 48131 44154
rect 48059 44064 48078 44098
rect 48112 44064 48131 44098
rect 48059 44008 48131 44064
rect 48059 43974 48078 44008
rect 48112 43974 48131 44008
rect 48059 43918 48131 43974
rect 47169 43843 47241 43903
rect 48059 43884 48078 43918
rect 48112 43884 48131 43918
rect 48059 43843 48131 43884
rect 47169 43824 48131 43843
rect 47169 43790 47266 43824
rect 47300 43790 47356 43824
rect 47390 43790 47446 43824
rect 47480 43790 47536 43824
rect 47570 43790 47626 43824
rect 47660 43790 47716 43824
rect 47750 43790 47806 43824
rect 47840 43790 47896 43824
rect 47930 43790 47986 43824
rect 48020 43790 48131 43824
rect 47169 43771 48131 43790
rect 48509 44714 49471 44733
rect 48509 44680 48640 44714
rect 48674 44680 48730 44714
rect 48764 44680 48820 44714
rect 48854 44680 48910 44714
rect 48944 44680 49000 44714
rect 49034 44680 49090 44714
rect 49124 44680 49180 44714
rect 49214 44680 49270 44714
rect 49304 44680 49360 44714
rect 49394 44680 49471 44714
rect 48509 44661 49471 44680
rect 48509 44657 48581 44661
rect 48509 44623 48528 44657
rect 48562 44623 48581 44657
rect 48509 44567 48581 44623
rect 49399 44638 49471 44661
rect 49399 44604 49418 44638
rect 49452 44604 49471 44638
rect 48509 44533 48528 44567
rect 48562 44533 48581 44567
rect 48509 44477 48581 44533
rect 48509 44443 48528 44477
rect 48562 44443 48581 44477
rect 48509 44387 48581 44443
rect 48509 44353 48528 44387
rect 48562 44353 48581 44387
rect 48509 44297 48581 44353
rect 48509 44263 48528 44297
rect 48562 44263 48581 44297
rect 48509 44207 48581 44263
rect 48509 44173 48528 44207
rect 48562 44173 48581 44207
rect 48509 44117 48581 44173
rect 48509 44083 48528 44117
rect 48562 44083 48581 44117
rect 48509 44027 48581 44083
rect 48509 43993 48528 44027
rect 48562 43993 48581 44027
rect 48509 43937 48581 43993
rect 48509 43903 48528 43937
rect 48562 43903 48581 43937
rect 49399 44548 49471 44604
rect 49399 44514 49418 44548
rect 49452 44514 49471 44548
rect 49399 44458 49471 44514
rect 49399 44424 49418 44458
rect 49452 44424 49471 44458
rect 49399 44368 49471 44424
rect 49399 44334 49418 44368
rect 49452 44334 49471 44368
rect 49399 44278 49471 44334
rect 49399 44244 49418 44278
rect 49452 44244 49471 44278
rect 49399 44188 49471 44244
rect 49399 44154 49418 44188
rect 49452 44154 49471 44188
rect 49399 44098 49471 44154
rect 49399 44064 49418 44098
rect 49452 44064 49471 44098
rect 49399 44008 49471 44064
rect 49399 43974 49418 44008
rect 49452 43974 49471 44008
rect 49399 43918 49471 43974
rect 48509 43843 48581 43903
rect 49399 43884 49418 43918
rect 49452 43884 49471 43918
rect 49399 43843 49471 43884
rect 48509 43824 49471 43843
rect 48509 43790 48606 43824
rect 48640 43790 48696 43824
rect 48730 43790 48786 43824
rect 48820 43790 48876 43824
rect 48910 43790 48966 43824
rect 49000 43790 49056 43824
rect 49090 43790 49146 43824
rect 49180 43790 49236 43824
rect 49270 43790 49326 43824
rect 49360 43790 49471 43824
rect 48509 43771 49471 43790
rect 49849 44714 50811 44733
rect 49849 44680 49980 44714
rect 50014 44680 50070 44714
rect 50104 44680 50160 44714
rect 50194 44680 50250 44714
rect 50284 44680 50340 44714
rect 50374 44680 50430 44714
rect 50464 44680 50520 44714
rect 50554 44680 50610 44714
rect 50644 44680 50700 44714
rect 50734 44680 50811 44714
rect 49849 44661 50811 44680
rect 49849 44657 49921 44661
rect 49849 44623 49868 44657
rect 49902 44623 49921 44657
rect 49849 44567 49921 44623
rect 50739 44638 50811 44661
rect 50739 44604 50758 44638
rect 50792 44604 50811 44638
rect 49849 44533 49868 44567
rect 49902 44533 49921 44567
rect 49849 44477 49921 44533
rect 49849 44443 49868 44477
rect 49902 44443 49921 44477
rect 49849 44387 49921 44443
rect 49849 44353 49868 44387
rect 49902 44353 49921 44387
rect 49849 44297 49921 44353
rect 49849 44263 49868 44297
rect 49902 44263 49921 44297
rect 49849 44207 49921 44263
rect 49849 44173 49868 44207
rect 49902 44173 49921 44207
rect 49849 44117 49921 44173
rect 49849 44083 49868 44117
rect 49902 44083 49921 44117
rect 49849 44027 49921 44083
rect 49849 43993 49868 44027
rect 49902 43993 49921 44027
rect 49849 43937 49921 43993
rect 49849 43903 49868 43937
rect 49902 43903 49921 43937
rect 50739 44548 50811 44604
rect 50739 44514 50758 44548
rect 50792 44514 50811 44548
rect 50739 44458 50811 44514
rect 50739 44424 50758 44458
rect 50792 44424 50811 44458
rect 50739 44368 50811 44424
rect 50739 44334 50758 44368
rect 50792 44334 50811 44368
rect 50739 44278 50811 44334
rect 50739 44244 50758 44278
rect 50792 44244 50811 44278
rect 50739 44188 50811 44244
rect 50739 44154 50758 44188
rect 50792 44154 50811 44188
rect 50739 44098 50811 44154
rect 50739 44064 50758 44098
rect 50792 44064 50811 44098
rect 50739 44008 50811 44064
rect 50739 43974 50758 44008
rect 50792 43974 50811 44008
rect 50739 43918 50811 43974
rect 49849 43843 49921 43903
rect 50739 43884 50758 43918
rect 50792 43884 50811 43918
rect 50739 43843 50811 43884
rect 49849 43824 50811 43843
rect 49849 43790 49946 43824
rect 49980 43790 50036 43824
rect 50070 43790 50126 43824
rect 50160 43790 50216 43824
rect 50250 43790 50306 43824
rect 50340 43790 50396 43824
rect 50430 43790 50486 43824
rect 50520 43790 50576 43824
rect 50610 43790 50666 43824
rect 50700 43790 50811 43824
rect 49849 43771 50811 43790
rect 51189 44714 52151 44733
rect 51189 44680 51320 44714
rect 51354 44680 51410 44714
rect 51444 44680 51500 44714
rect 51534 44680 51590 44714
rect 51624 44680 51680 44714
rect 51714 44680 51770 44714
rect 51804 44680 51860 44714
rect 51894 44680 51950 44714
rect 51984 44680 52040 44714
rect 52074 44680 52151 44714
rect 51189 44661 52151 44680
rect 51189 44657 51261 44661
rect 51189 44623 51208 44657
rect 51242 44623 51261 44657
rect 51189 44567 51261 44623
rect 52079 44638 52151 44661
rect 52079 44604 52098 44638
rect 52132 44604 52151 44638
rect 51189 44533 51208 44567
rect 51242 44533 51261 44567
rect 51189 44477 51261 44533
rect 51189 44443 51208 44477
rect 51242 44443 51261 44477
rect 51189 44387 51261 44443
rect 51189 44353 51208 44387
rect 51242 44353 51261 44387
rect 51189 44297 51261 44353
rect 51189 44263 51208 44297
rect 51242 44263 51261 44297
rect 51189 44207 51261 44263
rect 51189 44173 51208 44207
rect 51242 44173 51261 44207
rect 51189 44117 51261 44173
rect 51189 44083 51208 44117
rect 51242 44083 51261 44117
rect 51189 44027 51261 44083
rect 51189 43993 51208 44027
rect 51242 43993 51261 44027
rect 51189 43937 51261 43993
rect 51189 43903 51208 43937
rect 51242 43903 51261 43937
rect 52079 44548 52151 44604
rect 52079 44514 52098 44548
rect 52132 44514 52151 44548
rect 52079 44458 52151 44514
rect 52079 44424 52098 44458
rect 52132 44424 52151 44458
rect 52079 44368 52151 44424
rect 52079 44334 52098 44368
rect 52132 44334 52151 44368
rect 52079 44278 52151 44334
rect 52079 44244 52098 44278
rect 52132 44244 52151 44278
rect 52079 44188 52151 44244
rect 52079 44154 52098 44188
rect 52132 44154 52151 44188
rect 52079 44098 52151 44154
rect 52079 44064 52098 44098
rect 52132 44064 52151 44098
rect 52079 44008 52151 44064
rect 52079 43974 52098 44008
rect 52132 43974 52151 44008
rect 52079 43918 52151 43974
rect 51189 43843 51261 43903
rect 52079 43884 52098 43918
rect 52132 43884 52151 43918
rect 52079 43843 52151 43884
rect 51189 43824 52151 43843
rect 51189 43790 51286 43824
rect 51320 43790 51376 43824
rect 51410 43790 51466 43824
rect 51500 43790 51556 43824
rect 51590 43790 51646 43824
rect 51680 43790 51736 43824
rect 51770 43790 51826 43824
rect 51860 43790 51916 43824
rect 51950 43790 52006 43824
rect 52040 43790 52151 43824
rect 51189 43771 52151 43790
rect 23672 41359 23792 41362
rect 22614 41309 22654 41352
rect 23672 41325 23717 41359
rect 23751 41325 23792 41359
rect 23672 41322 23792 41325
rect 24972 41359 25092 41362
rect 24972 41325 25017 41359
rect 25051 41325 25092 41359
rect 24972 41322 25092 41325
rect 26272 41359 26392 41362
rect 26272 41325 26317 41359
rect 26351 41325 26392 41359
rect 30336 41359 30456 41362
rect 26272 41322 26392 41325
rect 22614 41275 22617 41309
rect 22651 41275 22654 41309
rect 22614 41232 22654 41275
rect 29278 41309 29318 41352
rect 30336 41325 30381 41359
rect 30415 41325 30456 41359
rect 30336 41322 30456 41325
rect 31636 41359 31756 41362
rect 31636 41325 31681 41359
rect 31715 41325 31756 41359
rect 31636 41322 31756 41325
rect 32936 41359 33056 41362
rect 32936 41325 32981 41359
rect 33015 41325 33056 41359
rect 32936 41322 33056 41325
rect 29278 41275 29281 41309
rect 29315 41275 29318 41309
rect 29278 41232 29318 41275
rect 41973 40954 42935 40973
rect 41973 40920 42104 40954
rect 42138 40920 42194 40954
rect 42228 40920 42284 40954
rect 42318 40920 42374 40954
rect 42408 40920 42464 40954
rect 42498 40920 42554 40954
rect 42588 40920 42644 40954
rect 42678 40920 42734 40954
rect 42768 40920 42824 40954
rect 42858 40920 42935 40954
rect 41973 40901 42935 40920
rect 41973 40897 42045 40901
rect 41973 40863 41992 40897
rect 42026 40863 42045 40897
rect 41973 40807 42045 40863
rect 42863 40878 42935 40901
rect 42863 40844 42882 40878
rect 42916 40844 42935 40878
rect 41973 40773 41992 40807
rect 42026 40773 42045 40807
rect 41973 40717 42045 40773
rect 41973 40683 41992 40717
rect 42026 40683 42045 40717
rect 41973 40627 42045 40683
rect 41973 40593 41992 40627
rect 42026 40593 42045 40627
rect 41973 40537 42045 40593
rect 41973 40503 41992 40537
rect 42026 40503 42045 40537
rect 41973 40447 42045 40503
rect 41973 40413 41992 40447
rect 42026 40413 42045 40447
rect 41973 40357 42045 40413
rect 41973 40323 41992 40357
rect 42026 40323 42045 40357
rect 41973 40267 42045 40323
rect 41973 40233 41992 40267
rect 42026 40233 42045 40267
rect 41973 40177 42045 40233
rect 41973 40143 41992 40177
rect 42026 40143 42045 40177
rect 42863 40788 42935 40844
rect 42863 40754 42882 40788
rect 42916 40754 42935 40788
rect 42863 40698 42935 40754
rect 42863 40664 42882 40698
rect 42916 40664 42935 40698
rect 42863 40608 42935 40664
rect 42863 40574 42882 40608
rect 42916 40574 42935 40608
rect 42863 40518 42935 40574
rect 42863 40484 42882 40518
rect 42916 40484 42935 40518
rect 42863 40428 42935 40484
rect 42863 40394 42882 40428
rect 42916 40394 42935 40428
rect 42863 40338 42935 40394
rect 42863 40304 42882 40338
rect 42916 40304 42935 40338
rect 42863 40248 42935 40304
rect 42863 40214 42882 40248
rect 42916 40214 42935 40248
rect 42863 40158 42935 40214
rect 41973 40083 42045 40143
rect 42863 40124 42882 40158
rect 42916 40124 42935 40158
rect 42863 40083 42935 40124
rect 41973 40064 42935 40083
rect 41973 40030 42070 40064
rect 42104 40030 42160 40064
rect 42194 40030 42250 40064
rect 42284 40030 42340 40064
rect 42374 40030 42430 40064
rect 42464 40030 42520 40064
rect 42554 40030 42610 40064
rect 42644 40030 42700 40064
rect 42734 40030 42790 40064
rect 42824 40030 42935 40064
rect 41973 40011 42935 40030
rect 43313 40954 44275 40973
rect 43313 40920 43444 40954
rect 43478 40920 43534 40954
rect 43568 40920 43624 40954
rect 43658 40920 43714 40954
rect 43748 40920 43804 40954
rect 43838 40920 43894 40954
rect 43928 40920 43984 40954
rect 44018 40920 44074 40954
rect 44108 40920 44164 40954
rect 44198 40920 44275 40954
rect 43313 40901 44275 40920
rect 43313 40897 43385 40901
rect 43313 40863 43332 40897
rect 43366 40863 43385 40897
rect 43313 40807 43385 40863
rect 44203 40878 44275 40901
rect 44203 40844 44222 40878
rect 44256 40844 44275 40878
rect 43313 40773 43332 40807
rect 43366 40773 43385 40807
rect 43313 40717 43385 40773
rect 43313 40683 43332 40717
rect 43366 40683 43385 40717
rect 43313 40627 43385 40683
rect 43313 40593 43332 40627
rect 43366 40593 43385 40627
rect 43313 40537 43385 40593
rect 43313 40503 43332 40537
rect 43366 40503 43385 40537
rect 43313 40447 43385 40503
rect 43313 40413 43332 40447
rect 43366 40413 43385 40447
rect 43313 40357 43385 40413
rect 43313 40323 43332 40357
rect 43366 40323 43385 40357
rect 43313 40267 43385 40323
rect 43313 40233 43332 40267
rect 43366 40233 43385 40267
rect 43313 40177 43385 40233
rect 43313 40143 43332 40177
rect 43366 40143 43385 40177
rect 44203 40788 44275 40844
rect 44203 40754 44222 40788
rect 44256 40754 44275 40788
rect 44203 40698 44275 40754
rect 44203 40664 44222 40698
rect 44256 40664 44275 40698
rect 44203 40608 44275 40664
rect 44203 40574 44222 40608
rect 44256 40574 44275 40608
rect 44203 40518 44275 40574
rect 44203 40484 44222 40518
rect 44256 40484 44275 40518
rect 44203 40428 44275 40484
rect 44203 40394 44222 40428
rect 44256 40394 44275 40428
rect 44203 40338 44275 40394
rect 44203 40304 44222 40338
rect 44256 40304 44275 40338
rect 44203 40248 44275 40304
rect 44203 40214 44222 40248
rect 44256 40214 44275 40248
rect 44203 40158 44275 40214
rect 43313 40083 43385 40143
rect 44203 40124 44222 40158
rect 44256 40124 44275 40158
rect 44203 40083 44275 40124
rect 43313 40064 44275 40083
rect 43313 40030 43410 40064
rect 43444 40030 43500 40064
rect 43534 40030 43590 40064
rect 43624 40030 43680 40064
rect 43714 40030 43770 40064
rect 43804 40030 43860 40064
rect 43894 40030 43950 40064
rect 43984 40030 44040 40064
rect 44074 40030 44130 40064
rect 44164 40030 44275 40064
rect 43313 40011 44275 40030
rect 44653 40954 45615 40973
rect 44653 40920 44784 40954
rect 44818 40920 44874 40954
rect 44908 40920 44964 40954
rect 44998 40920 45054 40954
rect 45088 40920 45144 40954
rect 45178 40920 45234 40954
rect 45268 40920 45324 40954
rect 45358 40920 45414 40954
rect 45448 40920 45504 40954
rect 45538 40920 45615 40954
rect 44653 40901 45615 40920
rect 44653 40897 44725 40901
rect 44653 40863 44672 40897
rect 44706 40863 44725 40897
rect 44653 40807 44725 40863
rect 45543 40878 45615 40901
rect 45543 40844 45562 40878
rect 45596 40844 45615 40878
rect 44653 40773 44672 40807
rect 44706 40773 44725 40807
rect 44653 40717 44725 40773
rect 44653 40683 44672 40717
rect 44706 40683 44725 40717
rect 44653 40627 44725 40683
rect 44653 40593 44672 40627
rect 44706 40593 44725 40627
rect 44653 40537 44725 40593
rect 44653 40503 44672 40537
rect 44706 40503 44725 40537
rect 44653 40447 44725 40503
rect 44653 40413 44672 40447
rect 44706 40413 44725 40447
rect 44653 40357 44725 40413
rect 44653 40323 44672 40357
rect 44706 40323 44725 40357
rect 44653 40267 44725 40323
rect 44653 40233 44672 40267
rect 44706 40233 44725 40267
rect 44653 40177 44725 40233
rect 44653 40143 44672 40177
rect 44706 40143 44725 40177
rect 45543 40788 45615 40844
rect 45543 40754 45562 40788
rect 45596 40754 45615 40788
rect 45543 40698 45615 40754
rect 45543 40664 45562 40698
rect 45596 40664 45615 40698
rect 45543 40608 45615 40664
rect 45543 40574 45562 40608
rect 45596 40574 45615 40608
rect 45543 40518 45615 40574
rect 45543 40484 45562 40518
rect 45596 40484 45615 40518
rect 45543 40428 45615 40484
rect 45543 40394 45562 40428
rect 45596 40394 45615 40428
rect 45543 40338 45615 40394
rect 45543 40304 45562 40338
rect 45596 40304 45615 40338
rect 45543 40248 45615 40304
rect 45543 40214 45562 40248
rect 45596 40214 45615 40248
rect 45543 40158 45615 40214
rect 44653 40083 44725 40143
rect 45543 40124 45562 40158
rect 45596 40124 45615 40158
rect 45543 40083 45615 40124
rect 44653 40064 45615 40083
rect 44653 40030 44750 40064
rect 44784 40030 44840 40064
rect 44874 40030 44930 40064
rect 44964 40030 45020 40064
rect 45054 40030 45110 40064
rect 45144 40030 45200 40064
rect 45234 40030 45290 40064
rect 45324 40030 45380 40064
rect 45414 40030 45470 40064
rect 45504 40030 45615 40064
rect 44653 40011 45615 40030
rect 45993 40954 46955 40973
rect 45993 40920 46124 40954
rect 46158 40920 46214 40954
rect 46248 40920 46304 40954
rect 46338 40920 46394 40954
rect 46428 40920 46484 40954
rect 46518 40920 46574 40954
rect 46608 40920 46664 40954
rect 46698 40920 46754 40954
rect 46788 40920 46844 40954
rect 46878 40920 46955 40954
rect 45993 40901 46955 40920
rect 45993 40897 46065 40901
rect 45993 40863 46012 40897
rect 46046 40863 46065 40897
rect 45993 40807 46065 40863
rect 46883 40878 46955 40901
rect 46883 40844 46902 40878
rect 46936 40844 46955 40878
rect 45993 40773 46012 40807
rect 46046 40773 46065 40807
rect 45993 40717 46065 40773
rect 45993 40683 46012 40717
rect 46046 40683 46065 40717
rect 45993 40627 46065 40683
rect 45993 40593 46012 40627
rect 46046 40593 46065 40627
rect 45993 40537 46065 40593
rect 45993 40503 46012 40537
rect 46046 40503 46065 40537
rect 45993 40447 46065 40503
rect 45993 40413 46012 40447
rect 46046 40413 46065 40447
rect 45993 40357 46065 40413
rect 45993 40323 46012 40357
rect 46046 40323 46065 40357
rect 45993 40267 46065 40323
rect 45993 40233 46012 40267
rect 46046 40233 46065 40267
rect 45993 40177 46065 40233
rect 45993 40143 46012 40177
rect 46046 40143 46065 40177
rect 46883 40788 46955 40844
rect 46883 40754 46902 40788
rect 46936 40754 46955 40788
rect 46883 40698 46955 40754
rect 46883 40664 46902 40698
rect 46936 40664 46955 40698
rect 46883 40608 46955 40664
rect 46883 40574 46902 40608
rect 46936 40574 46955 40608
rect 46883 40518 46955 40574
rect 46883 40484 46902 40518
rect 46936 40484 46955 40518
rect 46883 40428 46955 40484
rect 46883 40394 46902 40428
rect 46936 40394 46955 40428
rect 46883 40338 46955 40394
rect 46883 40304 46902 40338
rect 46936 40304 46955 40338
rect 46883 40248 46955 40304
rect 46883 40214 46902 40248
rect 46936 40214 46955 40248
rect 46883 40158 46955 40214
rect 45993 40083 46065 40143
rect 46883 40124 46902 40158
rect 46936 40124 46955 40158
rect 46883 40083 46955 40124
rect 45993 40064 46955 40083
rect 45993 40030 46090 40064
rect 46124 40030 46180 40064
rect 46214 40030 46270 40064
rect 46304 40030 46360 40064
rect 46394 40030 46450 40064
rect 46484 40030 46540 40064
rect 46574 40030 46630 40064
rect 46664 40030 46720 40064
rect 46754 40030 46810 40064
rect 46844 40030 46955 40064
rect 45993 40011 46955 40030
rect 47333 40954 48295 40973
rect 47333 40920 47464 40954
rect 47498 40920 47554 40954
rect 47588 40920 47644 40954
rect 47678 40920 47734 40954
rect 47768 40920 47824 40954
rect 47858 40920 47914 40954
rect 47948 40920 48004 40954
rect 48038 40920 48094 40954
rect 48128 40920 48184 40954
rect 48218 40920 48295 40954
rect 47333 40901 48295 40920
rect 47333 40897 47405 40901
rect 47333 40863 47352 40897
rect 47386 40863 47405 40897
rect 47333 40807 47405 40863
rect 48223 40878 48295 40901
rect 48223 40844 48242 40878
rect 48276 40844 48295 40878
rect 47333 40773 47352 40807
rect 47386 40773 47405 40807
rect 47333 40717 47405 40773
rect 47333 40683 47352 40717
rect 47386 40683 47405 40717
rect 47333 40627 47405 40683
rect 47333 40593 47352 40627
rect 47386 40593 47405 40627
rect 47333 40537 47405 40593
rect 47333 40503 47352 40537
rect 47386 40503 47405 40537
rect 47333 40447 47405 40503
rect 47333 40413 47352 40447
rect 47386 40413 47405 40447
rect 47333 40357 47405 40413
rect 47333 40323 47352 40357
rect 47386 40323 47405 40357
rect 47333 40267 47405 40323
rect 47333 40233 47352 40267
rect 47386 40233 47405 40267
rect 47333 40177 47405 40233
rect 47333 40143 47352 40177
rect 47386 40143 47405 40177
rect 48223 40788 48295 40844
rect 48223 40754 48242 40788
rect 48276 40754 48295 40788
rect 48223 40698 48295 40754
rect 48223 40664 48242 40698
rect 48276 40664 48295 40698
rect 48223 40608 48295 40664
rect 48223 40574 48242 40608
rect 48276 40574 48295 40608
rect 48223 40518 48295 40574
rect 48223 40484 48242 40518
rect 48276 40484 48295 40518
rect 48223 40428 48295 40484
rect 48223 40394 48242 40428
rect 48276 40394 48295 40428
rect 48223 40338 48295 40394
rect 48223 40304 48242 40338
rect 48276 40304 48295 40338
rect 48223 40248 48295 40304
rect 48223 40214 48242 40248
rect 48276 40214 48295 40248
rect 48223 40158 48295 40214
rect 47333 40083 47405 40143
rect 48223 40124 48242 40158
rect 48276 40124 48295 40158
rect 48223 40083 48295 40124
rect 47333 40064 48295 40083
rect 47333 40030 47430 40064
rect 47464 40030 47520 40064
rect 47554 40030 47610 40064
rect 47644 40030 47700 40064
rect 47734 40030 47790 40064
rect 47824 40030 47880 40064
rect 47914 40030 47970 40064
rect 48004 40030 48060 40064
rect 48094 40030 48150 40064
rect 48184 40030 48295 40064
rect 47333 40011 48295 40030
rect 48673 40954 49635 40973
rect 48673 40920 48804 40954
rect 48838 40920 48894 40954
rect 48928 40920 48984 40954
rect 49018 40920 49074 40954
rect 49108 40920 49164 40954
rect 49198 40920 49254 40954
rect 49288 40920 49344 40954
rect 49378 40920 49434 40954
rect 49468 40920 49524 40954
rect 49558 40920 49635 40954
rect 48673 40901 49635 40920
rect 48673 40897 48745 40901
rect 48673 40863 48692 40897
rect 48726 40863 48745 40897
rect 48673 40807 48745 40863
rect 49563 40878 49635 40901
rect 49563 40844 49582 40878
rect 49616 40844 49635 40878
rect 48673 40773 48692 40807
rect 48726 40773 48745 40807
rect 48673 40717 48745 40773
rect 48673 40683 48692 40717
rect 48726 40683 48745 40717
rect 48673 40627 48745 40683
rect 48673 40593 48692 40627
rect 48726 40593 48745 40627
rect 48673 40537 48745 40593
rect 48673 40503 48692 40537
rect 48726 40503 48745 40537
rect 48673 40447 48745 40503
rect 48673 40413 48692 40447
rect 48726 40413 48745 40447
rect 48673 40357 48745 40413
rect 48673 40323 48692 40357
rect 48726 40323 48745 40357
rect 48673 40267 48745 40323
rect 48673 40233 48692 40267
rect 48726 40233 48745 40267
rect 48673 40177 48745 40233
rect 48673 40143 48692 40177
rect 48726 40143 48745 40177
rect 49563 40788 49635 40844
rect 49563 40754 49582 40788
rect 49616 40754 49635 40788
rect 49563 40698 49635 40754
rect 49563 40664 49582 40698
rect 49616 40664 49635 40698
rect 49563 40608 49635 40664
rect 49563 40574 49582 40608
rect 49616 40574 49635 40608
rect 49563 40518 49635 40574
rect 49563 40484 49582 40518
rect 49616 40484 49635 40518
rect 49563 40428 49635 40484
rect 49563 40394 49582 40428
rect 49616 40394 49635 40428
rect 49563 40338 49635 40394
rect 49563 40304 49582 40338
rect 49616 40304 49635 40338
rect 49563 40248 49635 40304
rect 49563 40214 49582 40248
rect 49616 40214 49635 40248
rect 49563 40158 49635 40214
rect 48673 40083 48745 40143
rect 49563 40124 49582 40158
rect 49616 40124 49635 40158
rect 49563 40083 49635 40124
rect 48673 40064 49635 40083
rect 48673 40030 48770 40064
rect 48804 40030 48860 40064
rect 48894 40030 48950 40064
rect 48984 40030 49040 40064
rect 49074 40030 49130 40064
rect 49164 40030 49220 40064
rect 49254 40030 49310 40064
rect 49344 40030 49400 40064
rect 49434 40030 49490 40064
rect 49524 40030 49635 40064
rect 48673 40011 49635 40030
rect 50013 40954 50975 40973
rect 50013 40920 50144 40954
rect 50178 40920 50234 40954
rect 50268 40920 50324 40954
rect 50358 40920 50414 40954
rect 50448 40920 50504 40954
rect 50538 40920 50594 40954
rect 50628 40920 50684 40954
rect 50718 40920 50774 40954
rect 50808 40920 50864 40954
rect 50898 40920 50975 40954
rect 50013 40901 50975 40920
rect 50013 40897 50085 40901
rect 50013 40863 50032 40897
rect 50066 40863 50085 40897
rect 50013 40807 50085 40863
rect 50903 40878 50975 40901
rect 50903 40844 50922 40878
rect 50956 40844 50975 40878
rect 50013 40773 50032 40807
rect 50066 40773 50085 40807
rect 50013 40717 50085 40773
rect 50013 40683 50032 40717
rect 50066 40683 50085 40717
rect 50013 40627 50085 40683
rect 50013 40593 50032 40627
rect 50066 40593 50085 40627
rect 50013 40537 50085 40593
rect 50013 40503 50032 40537
rect 50066 40503 50085 40537
rect 50013 40447 50085 40503
rect 50013 40413 50032 40447
rect 50066 40413 50085 40447
rect 50013 40357 50085 40413
rect 50013 40323 50032 40357
rect 50066 40323 50085 40357
rect 50013 40267 50085 40323
rect 50013 40233 50032 40267
rect 50066 40233 50085 40267
rect 50013 40177 50085 40233
rect 50013 40143 50032 40177
rect 50066 40143 50085 40177
rect 50903 40788 50975 40844
rect 50903 40754 50922 40788
rect 50956 40754 50975 40788
rect 50903 40698 50975 40754
rect 50903 40664 50922 40698
rect 50956 40664 50975 40698
rect 50903 40608 50975 40664
rect 50903 40574 50922 40608
rect 50956 40574 50975 40608
rect 50903 40518 50975 40574
rect 50903 40484 50922 40518
rect 50956 40484 50975 40518
rect 50903 40428 50975 40484
rect 50903 40394 50922 40428
rect 50956 40394 50975 40428
rect 50903 40338 50975 40394
rect 50903 40304 50922 40338
rect 50956 40304 50975 40338
rect 50903 40248 50975 40304
rect 50903 40214 50922 40248
rect 50956 40214 50975 40248
rect 50903 40158 50975 40214
rect 50013 40083 50085 40143
rect 50903 40124 50922 40158
rect 50956 40124 50975 40158
rect 50903 40083 50975 40124
rect 50013 40064 50975 40083
rect 50013 40030 50110 40064
rect 50144 40030 50200 40064
rect 50234 40030 50290 40064
rect 50324 40030 50380 40064
rect 50414 40030 50470 40064
rect 50504 40030 50560 40064
rect 50594 40030 50650 40064
rect 50684 40030 50740 40064
rect 50774 40030 50830 40064
rect 50864 40030 50975 40064
rect 50013 40011 50975 40030
rect 51353 40954 52315 40973
rect 51353 40920 51484 40954
rect 51518 40920 51574 40954
rect 51608 40920 51664 40954
rect 51698 40920 51754 40954
rect 51788 40920 51844 40954
rect 51878 40920 51934 40954
rect 51968 40920 52024 40954
rect 52058 40920 52114 40954
rect 52148 40920 52204 40954
rect 52238 40920 52315 40954
rect 51353 40901 52315 40920
rect 51353 40897 51425 40901
rect 51353 40863 51372 40897
rect 51406 40863 51425 40897
rect 51353 40807 51425 40863
rect 52243 40878 52315 40901
rect 52243 40844 52262 40878
rect 52296 40844 52315 40878
rect 51353 40773 51372 40807
rect 51406 40773 51425 40807
rect 51353 40717 51425 40773
rect 51353 40683 51372 40717
rect 51406 40683 51425 40717
rect 51353 40627 51425 40683
rect 51353 40593 51372 40627
rect 51406 40593 51425 40627
rect 51353 40537 51425 40593
rect 51353 40503 51372 40537
rect 51406 40503 51425 40537
rect 51353 40447 51425 40503
rect 51353 40413 51372 40447
rect 51406 40413 51425 40447
rect 51353 40357 51425 40413
rect 51353 40323 51372 40357
rect 51406 40323 51425 40357
rect 51353 40267 51425 40323
rect 51353 40233 51372 40267
rect 51406 40233 51425 40267
rect 51353 40177 51425 40233
rect 51353 40143 51372 40177
rect 51406 40143 51425 40177
rect 52243 40788 52315 40844
rect 52243 40754 52262 40788
rect 52296 40754 52315 40788
rect 52243 40698 52315 40754
rect 52243 40664 52262 40698
rect 52296 40664 52315 40698
rect 52243 40608 52315 40664
rect 52243 40574 52262 40608
rect 52296 40574 52315 40608
rect 52243 40518 52315 40574
rect 52243 40484 52262 40518
rect 52296 40484 52315 40518
rect 52243 40428 52315 40484
rect 52243 40394 52262 40428
rect 52296 40394 52315 40428
rect 52243 40338 52315 40394
rect 52243 40304 52262 40338
rect 52296 40304 52315 40338
rect 52243 40248 52315 40304
rect 52243 40214 52262 40248
rect 52296 40214 52315 40248
rect 52243 40158 52315 40214
rect 51353 40083 51425 40143
rect 52243 40124 52262 40158
rect 52296 40124 52315 40158
rect 52243 40083 52315 40124
rect 51353 40064 52315 40083
rect 51353 40030 51450 40064
rect 51484 40030 51540 40064
rect 51574 40030 51630 40064
rect 51664 40030 51720 40064
rect 51754 40030 51810 40064
rect 51844 40030 51900 40064
rect 51934 40030 51990 40064
rect 52024 40030 52080 40064
rect 52114 40030 52170 40064
rect 52204 40030 52315 40064
rect 51353 40011 52315 40030
rect 38470 37599 38590 37602
rect 37412 37549 37452 37592
rect 38470 37565 38515 37599
rect 38549 37565 38590 37599
rect 38470 37562 38590 37565
rect 37412 37515 37415 37549
rect 37449 37515 37452 37549
rect 37412 37472 37452 37515
rect 12181 37194 13143 37213
rect 12181 37160 12312 37194
rect 12346 37160 12402 37194
rect 12436 37160 12492 37194
rect 12526 37160 12582 37194
rect 12616 37160 12672 37194
rect 12706 37160 12762 37194
rect 12796 37160 12852 37194
rect 12886 37160 12942 37194
rect 12976 37160 13032 37194
rect 13066 37160 13143 37194
rect 12181 37141 13143 37160
rect 12181 37137 12253 37141
rect 12181 37103 12200 37137
rect 12234 37103 12253 37137
rect 12181 37047 12253 37103
rect 13071 37118 13143 37141
rect 13071 37084 13090 37118
rect 13124 37084 13143 37118
rect 12181 37013 12200 37047
rect 12234 37013 12253 37047
rect 12181 36957 12253 37013
rect 12181 36923 12200 36957
rect 12234 36923 12253 36957
rect 12181 36867 12253 36923
rect 12181 36833 12200 36867
rect 12234 36833 12253 36867
rect 12181 36777 12253 36833
rect 12181 36743 12200 36777
rect 12234 36743 12253 36777
rect 12181 36687 12253 36743
rect 12181 36653 12200 36687
rect 12234 36653 12253 36687
rect 12181 36597 12253 36653
rect 12181 36563 12200 36597
rect 12234 36563 12253 36597
rect 12181 36507 12253 36563
rect 12181 36473 12200 36507
rect 12234 36473 12253 36507
rect 12181 36417 12253 36473
rect 12181 36383 12200 36417
rect 12234 36383 12253 36417
rect 13071 37028 13143 37084
rect 13071 36994 13090 37028
rect 13124 36994 13143 37028
rect 13071 36938 13143 36994
rect 13071 36904 13090 36938
rect 13124 36904 13143 36938
rect 13071 36848 13143 36904
rect 13071 36814 13090 36848
rect 13124 36814 13143 36848
rect 13071 36758 13143 36814
rect 13071 36724 13090 36758
rect 13124 36724 13143 36758
rect 13071 36668 13143 36724
rect 13071 36634 13090 36668
rect 13124 36634 13143 36668
rect 13071 36578 13143 36634
rect 13071 36544 13090 36578
rect 13124 36544 13143 36578
rect 13071 36488 13143 36544
rect 13071 36454 13090 36488
rect 13124 36454 13143 36488
rect 13071 36398 13143 36454
rect 12181 36323 12253 36383
rect 13071 36364 13090 36398
rect 13124 36364 13143 36398
rect 13071 36323 13143 36364
rect 12181 36304 13143 36323
rect 12181 36270 12278 36304
rect 12312 36270 12368 36304
rect 12402 36270 12458 36304
rect 12492 36270 12548 36304
rect 12582 36270 12638 36304
rect 12672 36270 12728 36304
rect 12762 36270 12818 36304
rect 12852 36270 12908 36304
rect 12942 36270 12998 36304
rect 13032 36270 13143 36304
rect 12181 36251 13143 36270
rect 41973 37194 42935 37213
rect 41973 37160 42104 37194
rect 42138 37160 42194 37194
rect 42228 37160 42284 37194
rect 42318 37160 42374 37194
rect 42408 37160 42464 37194
rect 42498 37160 42554 37194
rect 42588 37160 42644 37194
rect 42678 37160 42734 37194
rect 42768 37160 42824 37194
rect 42858 37160 42935 37194
rect 41973 37141 42935 37160
rect 41973 37137 42045 37141
rect 41973 37103 41992 37137
rect 42026 37103 42045 37137
rect 41973 37047 42045 37103
rect 42863 37118 42935 37141
rect 42863 37084 42882 37118
rect 42916 37084 42935 37118
rect 41973 37013 41992 37047
rect 42026 37013 42045 37047
rect 41973 36957 42045 37013
rect 41973 36923 41992 36957
rect 42026 36923 42045 36957
rect 41973 36867 42045 36923
rect 41973 36833 41992 36867
rect 42026 36833 42045 36867
rect 41973 36777 42045 36833
rect 41973 36743 41992 36777
rect 42026 36743 42045 36777
rect 41973 36687 42045 36743
rect 41973 36653 41992 36687
rect 42026 36653 42045 36687
rect 41973 36597 42045 36653
rect 41973 36563 41992 36597
rect 42026 36563 42045 36597
rect 41973 36507 42045 36563
rect 41973 36473 41992 36507
rect 42026 36473 42045 36507
rect 41973 36417 42045 36473
rect 41973 36383 41992 36417
rect 42026 36383 42045 36417
rect 42863 37028 42935 37084
rect 42863 36994 42882 37028
rect 42916 36994 42935 37028
rect 42863 36938 42935 36994
rect 42863 36904 42882 36938
rect 42916 36904 42935 36938
rect 42863 36848 42935 36904
rect 42863 36814 42882 36848
rect 42916 36814 42935 36848
rect 42863 36758 42935 36814
rect 42863 36724 42882 36758
rect 42916 36724 42935 36758
rect 42863 36668 42935 36724
rect 42863 36634 42882 36668
rect 42916 36634 42935 36668
rect 42863 36578 42935 36634
rect 42863 36544 42882 36578
rect 42916 36544 42935 36578
rect 42863 36488 42935 36544
rect 42863 36454 42882 36488
rect 42916 36454 42935 36488
rect 42863 36398 42935 36454
rect 41973 36323 42045 36383
rect 42863 36364 42882 36398
rect 42916 36364 42935 36398
rect 42863 36323 42935 36364
rect 41973 36304 42935 36323
rect 41973 36270 42070 36304
rect 42104 36270 42160 36304
rect 42194 36270 42250 36304
rect 42284 36270 42340 36304
rect 42374 36270 42430 36304
rect 42464 36270 42520 36304
rect 42554 36270 42610 36304
rect 42644 36270 42700 36304
rect 42734 36270 42790 36304
rect 42824 36270 42935 36304
rect 41973 36251 42935 36270
rect 43313 37194 44275 37213
rect 43313 37160 43444 37194
rect 43478 37160 43534 37194
rect 43568 37160 43624 37194
rect 43658 37160 43714 37194
rect 43748 37160 43804 37194
rect 43838 37160 43894 37194
rect 43928 37160 43984 37194
rect 44018 37160 44074 37194
rect 44108 37160 44164 37194
rect 44198 37160 44275 37194
rect 43313 37141 44275 37160
rect 43313 37137 43385 37141
rect 43313 37103 43332 37137
rect 43366 37103 43385 37137
rect 43313 37047 43385 37103
rect 44203 37118 44275 37141
rect 44203 37084 44222 37118
rect 44256 37084 44275 37118
rect 43313 37013 43332 37047
rect 43366 37013 43385 37047
rect 43313 36957 43385 37013
rect 43313 36923 43332 36957
rect 43366 36923 43385 36957
rect 43313 36867 43385 36923
rect 43313 36833 43332 36867
rect 43366 36833 43385 36867
rect 43313 36777 43385 36833
rect 43313 36743 43332 36777
rect 43366 36743 43385 36777
rect 43313 36687 43385 36743
rect 43313 36653 43332 36687
rect 43366 36653 43385 36687
rect 43313 36597 43385 36653
rect 43313 36563 43332 36597
rect 43366 36563 43385 36597
rect 43313 36507 43385 36563
rect 43313 36473 43332 36507
rect 43366 36473 43385 36507
rect 43313 36417 43385 36473
rect 43313 36383 43332 36417
rect 43366 36383 43385 36417
rect 44203 37028 44275 37084
rect 44203 36994 44222 37028
rect 44256 36994 44275 37028
rect 44203 36938 44275 36994
rect 44203 36904 44222 36938
rect 44256 36904 44275 36938
rect 44203 36848 44275 36904
rect 44203 36814 44222 36848
rect 44256 36814 44275 36848
rect 44203 36758 44275 36814
rect 44203 36724 44222 36758
rect 44256 36724 44275 36758
rect 44203 36668 44275 36724
rect 44203 36634 44222 36668
rect 44256 36634 44275 36668
rect 44203 36578 44275 36634
rect 44203 36544 44222 36578
rect 44256 36544 44275 36578
rect 44203 36488 44275 36544
rect 44203 36454 44222 36488
rect 44256 36454 44275 36488
rect 44203 36398 44275 36454
rect 43313 36323 43385 36383
rect 44203 36364 44222 36398
rect 44256 36364 44275 36398
rect 44203 36323 44275 36364
rect 43313 36304 44275 36323
rect 43313 36270 43410 36304
rect 43444 36270 43500 36304
rect 43534 36270 43590 36304
rect 43624 36270 43680 36304
rect 43714 36270 43770 36304
rect 43804 36270 43860 36304
rect 43894 36270 43950 36304
rect 43984 36270 44040 36304
rect 44074 36270 44130 36304
rect 44164 36270 44275 36304
rect 43313 36251 44275 36270
rect 44653 37194 45615 37213
rect 44653 37160 44784 37194
rect 44818 37160 44874 37194
rect 44908 37160 44964 37194
rect 44998 37160 45054 37194
rect 45088 37160 45144 37194
rect 45178 37160 45234 37194
rect 45268 37160 45324 37194
rect 45358 37160 45414 37194
rect 45448 37160 45504 37194
rect 45538 37160 45615 37194
rect 44653 37141 45615 37160
rect 44653 37137 44725 37141
rect 44653 37103 44672 37137
rect 44706 37103 44725 37137
rect 44653 37047 44725 37103
rect 45543 37118 45615 37141
rect 45543 37084 45562 37118
rect 45596 37084 45615 37118
rect 44653 37013 44672 37047
rect 44706 37013 44725 37047
rect 44653 36957 44725 37013
rect 44653 36923 44672 36957
rect 44706 36923 44725 36957
rect 44653 36867 44725 36923
rect 44653 36833 44672 36867
rect 44706 36833 44725 36867
rect 44653 36777 44725 36833
rect 44653 36743 44672 36777
rect 44706 36743 44725 36777
rect 44653 36687 44725 36743
rect 44653 36653 44672 36687
rect 44706 36653 44725 36687
rect 44653 36597 44725 36653
rect 44653 36563 44672 36597
rect 44706 36563 44725 36597
rect 44653 36507 44725 36563
rect 44653 36473 44672 36507
rect 44706 36473 44725 36507
rect 44653 36417 44725 36473
rect 44653 36383 44672 36417
rect 44706 36383 44725 36417
rect 45543 37028 45615 37084
rect 45543 36994 45562 37028
rect 45596 36994 45615 37028
rect 45543 36938 45615 36994
rect 45543 36904 45562 36938
rect 45596 36904 45615 36938
rect 45543 36848 45615 36904
rect 45543 36814 45562 36848
rect 45596 36814 45615 36848
rect 45543 36758 45615 36814
rect 45543 36724 45562 36758
rect 45596 36724 45615 36758
rect 45543 36668 45615 36724
rect 45543 36634 45562 36668
rect 45596 36634 45615 36668
rect 45543 36578 45615 36634
rect 45543 36544 45562 36578
rect 45596 36544 45615 36578
rect 45543 36488 45615 36544
rect 45543 36454 45562 36488
rect 45596 36454 45615 36488
rect 45543 36398 45615 36454
rect 44653 36323 44725 36383
rect 45543 36364 45562 36398
rect 45596 36364 45615 36398
rect 45543 36323 45615 36364
rect 44653 36304 45615 36323
rect 44653 36270 44750 36304
rect 44784 36270 44840 36304
rect 44874 36270 44930 36304
rect 44964 36270 45020 36304
rect 45054 36270 45110 36304
rect 45144 36270 45200 36304
rect 45234 36270 45290 36304
rect 45324 36270 45380 36304
rect 45414 36270 45470 36304
rect 45504 36270 45615 36304
rect 44653 36251 45615 36270
rect 45993 37194 46955 37213
rect 45993 37160 46124 37194
rect 46158 37160 46214 37194
rect 46248 37160 46304 37194
rect 46338 37160 46394 37194
rect 46428 37160 46484 37194
rect 46518 37160 46574 37194
rect 46608 37160 46664 37194
rect 46698 37160 46754 37194
rect 46788 37160 46844 37194
rect 46878 37160 46955 37194
rect 45993 37141 46955 37160
rect 45993 37137 46065 37141
rect 45993 37103 46012 37137
rect 46046 37103 46065 37137
rect 45993 37047 46065 37103
rect 46883 37118 46955 37141
rect 46883 37084 46902 37118
rect 46936 37084 46955 37118
rect 45993 37013 46012 37047
rect 46046 37013 46065 37047
rect 45993 36957 46065 37013
rect 45993 36923 46012 36957
rect 46046 36923 46065 36957
rect 45993 36867 46065 36923
rect 45993 36833 46012 36867
rect 46046 36833 46065 36867
rect 45993 36777 46065 36833
rect 45993 36743 46012 36777
rect 46046 36743 46065 36777
rect 45993 36687 46065 36743
rect 45993 36653 46012 36687
rect 46046 36653 46065 36687
rect 45993 36597 46065 36653
rect 45993 36563 46012 36597
rect 46046 36563 46065 36597
rect 45993 36507 46065 36563
rect 45993 36473 46012 36507
rect 46046 36473 46065 36507
rect 45993 36417 46065 36473
rect 45993 36383 46012 36417
rect 46046 36383 46065 36417
rect 46883 37028 46955 37084
rect 46883 36994 46902 37028
rect 46936 36994 46955 37028
rect 46883 36938 46955 36994
rect 46883 36904 46902 36938
rect 46936 36904 46955 36938
rect 46883 36848 46955 36904
rect 46883 36814 46902 36848
rect 46936 36814 46955 36848
rect 46883 36758 46955 36814
rect 46883 36724 46902 36758
rect 46936 36724 46955 36758
rect 46883 36668 46955 36724
rect 46883 36634 46902 36668
rect 46936 36634 46955 36668
rect 46883 36578 46955 36634
rect 46883 36544 46902 36578
rect 46936 36544 46955 36578
rect 46883 36488 46955 36544
rect 46883 36454 46902 36488
rect 46936 36454 46955 36488
rect 46883 36398 46955 36454
rect 45993 36323 46065 36383
rect 46883 36364 46902 36398
rect 46936 36364 46955 36398
rect 46883 36323 46955 36364
rect 45993 36304 46955 36323
rect 45993 36270 46090 36304
rect 46124 36270 46180 36304
rect 46214 36270 46270 36304
rect 46304 36270 46360 36304
rect 46394 36270 46450 36304
rect 46484 36270 46540 36304
rect 46574 36270 46630 36304
rect 46664 36270 46720 36304
rect 46754 36270 46810 36304
rect 46844 36270 46955 36304
rect 45993 36251 46955 36270
rect 47333 37194 48295 37213
rect 47333 37160 47464 37194
rect 47498 37160 47554 37194
rect 47588 37160 47644 37194
rect 47678 37160 47734 37194
rect 47768 37160 47824 37194
rect 47858 37160 47914 37194
rect 47948 37160 48004 37194
rect 48038 37160 48094 37194
rect 48128 37160 48184 37194
rect 48218 37160 48295 37194
rect 47333 37141 48295 37160
rect 47333 37137 47405 37141
rect 47333 37103 47352 37137
rect 47386 37103 47405 37137
rect 47333 37047 47405 37103
rect 48223 37118 48295 37141
rect 48223 37084 48242 37118
rect 48276 37084 48295 37118
rect 47333 37013 47352 37047
rect 47386 37013 47405 37047
rect 47333 36957 47405 37013
rect 47333 36923 47352 36957
rect 47386 36923 47405 36957
rect 47333 36867 47405 36923
rect 47333 36833 47352 36867
rect 47386 36833 47405 36867
rect 47333 36777 47405 36833
rect 47333 36743 47352 36777
rect 47386 36743 47405 36777
rect 47333 36687 47405 36743
rect 47333 36653 47352 36687
rect 47386 36653 47405 36687
rect 47333 36597 47405 36653
rect 47333 36563 47352 36597
rect 47386 36563 47405 36597
rect 47333 36507 47405 36563
rect 47333 36473 47352 36507
rect 47386 36473 47405 36507
rect 47333 36417 47405 36473
rect 47333 36383 47352 36417
rect 47386 36383 47405 36417
rect 48223 37028 48295 37084
rect 48223 36994 48242 37028
rect 48276 36994 48295 37028
rect 48223 36938 48295 36994
rect 48223 36904 48242 36938
rect 48276 36904 48295 36938
rect 48223 36848 48295 36904
rect 48223 36814 48242 36848
rect 48276 36814 48295 36848
rect 48223 36758 48295 36814
rect 48223 36724 48242 36758
rect 48276 36724 48295 36758
rect 48223 36668 48295 36724
rect 48223 36634 48242 36668
rect 48276 36634 48295 36668
rect 48223 36578 48295 36634
rect 48223 36544 48242 36578
rect 48276 36544 48295 36578
rect 48223 36488 48295 36544
rect 48223 36454 48242 36488
rect 48276 36454 48295 36488
rect 48223 36398 48295 36454
rect 47333 36323 47405 36383
rect 48223 36364 48242 36398
rect 48276 36364 48295 36398
rect 48223 36323 48295 36364
rect 47333 36304 48295 36323
rect 47333 36270 47430 36304
rect 47464 36270 47520 36304
rect 47554 36270 47610 36304
rect 47644 36270 47700 36304
rect 47734 36270 47790 36304
rect 47824 36270 47880 36304
rect 47914 36270 47970 36304
rect 48004 36270 48060 36304
rect 48094 36270 48150 36304
rect 48184 36270 48295 36304
rect 47333 36251 48295 36270
rect 48673 37194 49635 37213
rect 48673 37160 48804 37194
rect 48838 37160 48894 37194
rect 48928 37160 48984 37194
rect 49018 37160 49074 37194
rect 49108 37160 49164 37194
rect 49198 37160 49254 37194
rect 49288 37160 49344 37194
rect 49378 37160 49434 37194
rect 49468 37160 49524 37194
rect 49558 37160 49635 37194
rect 48673 37141 49635 37160
rect 48673 37137 48745 37141
rect 48673 37103 48692 37137
rect 48726 37103 48745 37137
rect 48673 37047 48745 37103
rect 49563 37118 49635 37141
rect 49563 37084 49582 37118
rect 49616 37084 49635 37118
rect 48673 37013 48692 37047
rect 48726 37013 48745 37047
rect 48673 36957 48745 37013
rect 48673 36923 48692 36957
rect 48726 36923 48745 36957
rect 48673 36867 48745 36923
rect 48673 36833 48692 36867
rect 48726 36833 48745 36867
rect 48673 36777 48745 36833
rect 48673 36743 48692 36777
rect 48726 36743 48745 36777
rect 48673 36687 48745 36743
rect 48673 36653 48692 36687
rect 48726 36653 48745 36687
rect 48673 36597 48745 36653
rect 48673 36563 48692 36597
rect 48726 36563 48745 36597
rect 48673 36507 48745 36563
rect 48673 36473 48692 36507
rect 48726 36473 48745 36507
rect 48673 36417 48745 36473
rect 48673 36383 48692 36417
rect 48726 36383 48745 36417
rect 49563 37028 49635 37084
rect 49563 36994 49582 37028
rect 49616 36994 49635 37028
rect 49563 36938 49635 36994
rect 49563 36904 49582 36938
rect 49616 36904 49635 36938
rect 49563 36848 49635 36904
rect 49563 36814 49582 36848
rect 49616 36814 49635 36848
rect 49563 36758 49635 36814
rect 49563 36724 49582 36758
rect 49616 36724 49635 36758
rect 49563 36668 49635 36724
rect 49563 36634 49582 36668
rect 49616 36634 49635 36668
rect 49563 36578 49635 36634
rect 49563 36544 49582 36578
rect 49616 36544 49635 36578
rect 49563 36488 49635 36544
rect 49563 36454 49582 36488
rect 49616 36454 49635 36488
rect 49563 36398 49635 36454
rect 48673 36323 48745 36383
rect 49563 36364 49582 36398
rect 49616 36364 49635 36398
rect 49563 36323 49635 36364
rect 48673 36304 49635 36323
rect 48673 36270 48770 36304
rect 48804 36270 48860 36304
rect 48894 36270 48950 36304
rect 48984 36270 49040 36304
rect 49074 36270 49130 36304
rect 49164 36270 49220 36304
rect 49254 36270 49310 36304
rect 49344 36270 49400 36304
rect 49434 36270 49490 36304
rect 49524 36270 49635 36304
rect 48673 36251 49635 36270
rect 50013 37194 50975 37213
rect 50013 37160 50144 37194
rect 50178 37160 50234 37194
rect 50268 37160 50324 37194
rect 50358 37160 50414 37194
rect 50448 37160 50504 37194
rect 50538 37160 50594 37194
rect 50628 37160 50684 37194
rect 50718 37160 50774 37194
rect 50808 37160 50864 37194
rect 50898 37160 50975 37194
rect 50013 37141 50975 37160
rect 50013 37137 50085 37141
rect 50013 37103 50032 37137
rect 50066 37103 50085 37137
rect 50013 37047 50085 37103
rect 50903 37118 50975 37141
rect 50903 37084 50922 37118
rect 50956 37084 50975 37118
rect 50013 37013 50032 37047
rect 50066 37013 50085 37047
rect 50013 36957 50085 37013
rect 50013 36923 50032 36957
rect 50066 36923 50085 36957
rect 50013 36867 50085 36923
rect 50013 36833 50032 36867
rect 50066 36833 50085 36867
rect 50013 36777 50085 36833
rect 50013 36743 50032 36777
rect 50066 36743 50085 36777
rect 50013 36687 50085 36743
rect 50013 36653 50032 36687
rect 50066 36653 50085 36687
rect 50013 36597 50085 36653
rect 50013 36563 50032 36597
rect 50066 36563 50085 36597
rect 50013 36507 50085 36563
rect 50013 36473 50032 36507
rect 50066 36473 50085 36507
rect 50013 36417 50085 36473
rect 50013 36383 50032 36417
rect 50066 36383 50085 36417
rect 50903 37028 50975 37084
rect 50903 36994 50922 37028
rect 50956 36994 50975 37028
rect 50903 36938 50975 36994
rect 50903 36904 50922 36938
rect 50956 36904 50975 36938
rect 50903 36848 50975 36904
rect 50903 36814 50922 36848
rect 50956 36814 50975 36848
rect 50903 36758 50975 36814
rect 50903 36724 50922 36758
rect 50956 36724 50975 36758
rect 50903 36668 50975 36724
rect 50903 36634 50922 36668
rect 50956 36634 50975 36668
rect 50903 36578 50975 36634
rect 50903 36544 50922 36578
rect 50956 36544 50975 36578
rect 50903 36488 50975 36544
rect 50903 36454 50922 36488
rect 50956 36454 50975 36488
rect 50903 36398 50975 36454
rect 50013 36323 50085 36383
rect 50903 36364 50922 36398
rect 50956 36364 50975 36398
rect 50903 36323 50975 36364
rect 50013 36304 50975 36323
rect 50013 36270 50110 36304
rect 50144 36270 50200 36304
rect 50234 36270 50290 36304
rect 50324 36270 50380 36304
rect 50414 36270 50470 36304
rect 50504 36270 50560 36304
rect 50594 36270 50650 36304
rect 50684 36270 50740 36304
rect 50774 36270 50830 36304
rect 50864 36270 50975 36304
rect 50013 36251 50975 36270
rect 51353 37194 52315 37213
rect 51353 37160 51484 37194
rect 51518 37160 51574 37194
rect 51608 37160 51664 37194
rect 51698 37160 51754 37194
rect 51788 37160 51844 37194
rect 51878 37160 51934 37194
rect 51968 37160 52024 37194
rect 52058 37160 52114 37194
rect 52148 37160 52204 37194
rect 52238 37160 52315 37194
rect 51353 37141 52315 37160
rect 51353 37137 51425 37141
rect 51353 37103 51372 37137
rect 51406 37103 51425 37137
rect 51353 37047 51425 37103
rect 52243 37118 52315 37141
rect 52243 37084 52262 37118
rect 52296 37084 52315 37118
rect 51353 37013 51372 37047
rect 51406 37013 51425 37047
rect 51353 36957 51425 37013
rect 51353 36923 51372 36957
rect 51406 36923 51425 36957
rect 51353 36867 51425 36923
rect 51353 36833 51372 36867
rect 51406 36833 51425 36867
rect 51353 36777 51425 36833
rect 51353 36743 51372 36777
rect 51406 36743 51425 36777
rect 51353 36687 51425 36743
rect 51353 36653 51372 36687
rect 51406 36653 51425 36687
rect 51353 36597 51425 36653
rect 51353 36563 51372 36597
rect 51406 36563 51425 36597
rect 51353 36507 51425 36563
rect 51353 36473 51372 36507
rect 51406 36473 51425 36507
rect 51353 36417 51425 36473
rect 51353 36383 51372 36417
rect 51406 36383 51425 36417
rect 52243 37028 52315 37084
rect 52243 36994 52262 37028
rect 52296 36994 52315 37028
rect 52243 36938 52315 36994
rect 52243 36904 52262 36938
rect 52296 36904 52315 36938
rect 52243 36848 52315 36904
rect 52243 36814 52262 36848
rect 52296 36814 52315 36848
rect 52243 36758 52315 36814
rect 52243 36724 52262 36758
rect 52296 36724 52315 36758
rect 52243 36668 52315 36724
rect 52243 36634 52262 36668
rect 52296 36634 52315 36668
rect 52243 36578 52315 36634
rect 52243 36544 52262 36578
rect 52296 36544 52315 36578
rect 52243 36488 52315 36544
rect 52243 36454 52262 36488
rect 52296 36454 52315 36488
rect 52243 36398 52315 36454
rect 51353 36323 51425 36383
rect 52243 36364 52262 36398
rect 52296 36364 52315 36398
rect 52243 36323 52315 36364
rect 51353 36304 52315 36323
rect 51353 36270 51450 36304
rect 51484 36270 51540 36304
rect 51574 36270 51630 36304
rect 51664 36270 51720 36304
rect 51754 36270 51810 36304
rect 51844 36270 51900 36304
rect 51934 36270 51990 36304
rect 52024 36270 52080 36304
rect 52114 36270 52170 36304
rect 52204 36270 52315 36304
rect 51353 36251 52315 36270
rect 41973 33434 42935 33453
rect 41973 33400 42104 33434
rect 42138 33400 42194 33434
rect 42228 33400 42284 33434
rect 42318 33400 42374 33434
rect 42408 33400 42464 33434
rect 42498 33400 42554 33434
rect 42588 33400 42644 33434
rect 42678 33400 42734 33434
rect 42768 33400 42824 33434
rect 42858 33400 42935 33434
rect 41973 33381 42935 33400
rect 41973 33377 42045 33381
rect 41973 33343 41992 33377
rect 42026 33343 42045 33377
rect 41973 33287 42045 33343
rect 42863 33358 42935 33381
rect 42863 33324 42882 33358
rect 42916 33324 42935 33358
rect 41973 33253 41992 33287
rect 42026 33253 42045 33287
rect 41973 33197 42045 33253
rect 41973 33163 41992 33197
rect 42026 33163 42045 33197
rect 41973 33107 42045 33163
rect 41973 33073 41992 33107
rect 42026 33073 42045 33107
rect 41973 33017 42045 33073
rect 41973 32983 41992 33017
rect 42026 32983 42045 33017
rect 41973 32927 42045 32983
rect 41973 32893 41992 32927
rect 42026 32893 42045 32927
rect 41973 32837 42045 32893
rect 41973 32803 41992 32837
rect 42026 32803 42045 32837
rect 41973 32747 42045 32803
rect 41973 32713 41992 32747
rect 42026 32713 42045 32747
rect 41973 32657 42045 32713
rect 41973 32623 41992 32657
rect 42026 32623 42045 32657
rect 42863 33268 42935 33324
rect 42863 33234 42882 33268
rect 42916 33234 42935 33268
rect 42863 33178 42935 33234
rect 42863 33144 42882 33178
rect 42916 33144 42935 33178
rect 42863 33088 42935 33144
rect 42863 33054 42882 33088
rect 42916 33054 42935 33088
rect 42863 32998 42935 33054
rect 42863 32964 42882 32998
rect 42916 32964 42935 32998
rect 42863 32908 42935 32964
rect 42863 32874 42882 32908
rect 42916 32874 42935 32908
rect 42863 32818 42935 32874
rect 42863 32784 42882 32818
rect 42916 32784 42935 32818
rect 42863 32728 42935 32784
rect 42863 32694 42882 32728
rect 42916 32694 42935 32728
rect 42863 32638 42935 32694
rect 41973 32563 42045 32623
rect 42863 32604 42882 32638
rect 42916 32604 42935 32638
rect 42863 32563 42935 32604
rect 41973 32544 42935 32563
rect 41973 32510 42070 32544
rect 42104 32510 42160 32544
rect 42194 32510 42250 32544
rect 42284 32510 42340 32544
rect 42374 32510 42430 32544
rect 42464 32510 42520 32544
rect 42554 32510 42610 32544
rect 42644 32510 42700 32544
rect 42734 32510 42790 32544
rect 42824 32510 42935 32544
rect 41973 32491 42935 32510
rect 43313 33434 44275 33453
rect 43313 33400 43444 33434
rect 43478 33400 43534 33434
rect 43568 33400 43624 33434
rect 43658 33400 43714 33434
rect 43748 33400 43804 33434
rect 43838 33400 43894 33434
rect 43928 33400 43984 33434
rect 44018 33400 44074 33434
rect 44108 33400 44164 33434
rect 44198 33400 44275 33434
rect 43313 33381 44275 33400
rect 43313 33377 43385 33381
rect 43313 33343 43332 33377
rect 43366 33343 43385 33377
rect 43313 33287 43385 33343
rect 44203 33358 44275 33381
rect 44203 33324 44222 33358
rect 44256 33324 44275 33358
rect 43313 33253 43332 33287
rect 43366 33253 43385 33287
rect 43313 33197 43385 33253
rect 43313 33163 43332 33197
rect 43366 33163 43385 33197
rect 43313 33107 43385 33163
rect 43313 33073 43332 33107
rect 43366 33073 43385 33107
rect 43313 33017 43385 33073
rect 43313 32983 43332 33017
rect 43366 32983 43385 33017
rect 43313 32927 43385 32983
rect 43313 32893 43332 32927
rect 43366 32893 43385 32927
rect 43313 32837 43385 32893
rect 43313 32803 43332 32837
rect 43366 32803 43385 32837
rect 43313 32747 43385 32803
rect 43313 32713 43332 32747
rect 43366 32713 43385 32747
rect 43313 32657 43385 32713
rect 43313 32623 43332 32657
rect 43366 32623 43385 32657
rect 44203 33268 44275 33324
rect 44203 33234 44222 33268
rect 44256 33234 44275 33268
rect 44203 33178 44275 33234
rect 44203 33144 44222 33178
rect 44256 33144 44275 33178
rect 44203 33088 44275 33144
rect 44203 33054 44222 33088
rect 44256 33054 44275 33088
rect 44203 32998 44275 33054
rect 44203 32964 44222 32998
rect 44256 32964 44275 32998
rect 44203 32908 44275 32964
rect 44203 32874 44222 32908
rect 44256 32874 44275 32908
rect 44203 32818 44275 32874
rect 44203 32784 44222 32818
rect 44256 32784 44275 32818
rect 44203 32728 44275 32784
rect 44203 32694 44222 32728
rect 44256 32694 44275 32728
rect 44203 32638 44275 32694
rect 43313 32563 43385 32623
rect 44203 32604 44222 32638
rect 44256 32604 44275 32638
rect 44203 32563 44275 32604
rect 43313 32544 44275 32563
rect 43313 32510 43410 32544
rect 43444 32510 43500 32544
rect 43534 32510 43590 32544
rect 43624 32510 43680 32544
rect 43714 32510 43770 32544
rect 43804 32510 43860 32544
rect 43894 32510 43950 32544
rect 43984 32510 44040 32544
rect 44074 32510 44130 32544
rect 44164 32510 44275 32544
rect 43313 32491 44275 32510
rect 44653 33434 45615 33453
rect 44653 33400 44784 33434
rect 44818 33400 44874 33434
rect 44908 33400 44964 33434
rect 44998 33400 45054 33434
rect 45088 33400 45144 33434
rect 45178 33400 45234 33434
rect 45268 33400 45324 33434
rect 45358 33400 45414 33434
rect 45448 33400 45504 33434
rect 45538 33400 45615 33434
rect 44653 33381 45615 33400
rect 44653 33377 44725 33381
rect 44653 33343 44672 33377
rect 44706 33343 44725 33377
rect 44653 33287 44725 33343
rect 45543 33358 45615 33381
rect 45543 33324 45562 33358
rect 45596 33324 45615 33358
rect 44653 33253 44672 33287
rect 44706 33253 44725 33287
rect 44653 33197 44725 33253
rect 44653 33163 44672 33197
rect 44706 33163 44725 33197
rect 44653 33107 44725 33163
rect 44653 33073 44672 33107
rect 44706 33073 44725 33107
rect 44653 33017 44725 33073
rect 44653 32983 44672 33017
rect 44706 32983 44725 33017
rect 44653 32927 44725 32983
rect 44653 32893 44672 32927
rect 44706 32893 44725 32927
rect 44653 32837 44725 32893
rect 44653 32803 44672 32837
rect 44706 32803 44725 32837
rect 44653 32747 44725 32803
rect 44653 32713 44672 32747
rect 44706 32713 44725 32747
rect 44653 32657 44725 32713
rect 44653 32623 44672 32657
rect 44706 32623 44725 32657
rect 45543 33268 45615 33324
rect 45543 33234 45562 33268
rect 45596 33234 45615 33268
rect 45543 33178 45615 33234
rect 45543 33144 45562 33178
rect 45596 33144 45615 33178
rect 45543 33088 45615 33144
rect 45543 33054 45562 33088
rect 45596 33054 45615 33088
rect 45543 32998 45615 33054
rect 45543 32964 45562 32998
rect 45596 32964 45615 32998
rect 45543 32908 45615 32964
rect 45543 32874 45562 32908
rect 45596 32874 45615 32908
rect 45543 32818 45615 32874
rect 45543 32784 45562 32818
rect 45596 32784 45615 32818
rect 45543 32728 45615 32784
rect 45543 32694 45562 32728
rect 45596 32694 45615 32728
rect 45543 32638 45615 32694
rect 44653 32563 44725 32623
rect 45543 32604 45562 32638
rect 45596 32604 45615 32638
rect 45543 32563 45615 32604
rect 44653 32544 45615 32563
rect 44653 32510 44750 32544
rect 44784 32510 44840 32544
rect 44874 32510 44930 32544
rect 44964 32510 45020 32544
rect 45054 32510 45110 32544
rect 45144 32510 45200 32544
rect 45234 32510 45290 32544
rect 45324 32510 45380 32544
rect 45414 32510 45470 32544
rect 45504 32510 45615 32544
rect 44653 32491 45615 32510
rect 45993 33434 46955 33453
rect 45993 33400 46124 33434
rect 46158 33400 46214 33434
rect 46248 33400 46304 33434
rect 46338 33400 46394 33434
rect 46428 33400 46484 33434
rect 46518 33400 46574 33434
rect 46608 33400 46664 33434
rect 46698 33400 46754 33434
rect 46788 33400 46844 33434
rect 46878 33400 46955 33434
rect 45993 33381 46955 33400
rect 45993 33377 46065 33381
rect 45993 33343 46012 33377
rect 46046 33343 46065 33377
rect 45993 33287 46065 33343
rect 46883 33358 46955 33381
rect 46883 33324 46902 33358
rect 46936 33324 46955 33358
rect 45993 33253 46012 33287
rect 46046 33253 46065 33287
rect 45993 33197 46065 33253
rect 45993 33163 46012 33197
rect 46046 33163 46065 33197
rect 45993 33107 46065 33163
rect 45993 33073 46012 33107
rect 46046 33073 46065 33107
rect 45993 33017 46065 33073
rect 45993 32983 46012 33017
rect 46046 32983 46065 33017
rect 45993 32927 46065 32983
rect 45993 32893 46012 32927
rect 46046 32893 46065 32927
rect 45993 32837 46065 32893
rect 45993 32803 46012 32837
rect 46046 32803 46065 32837
rect 45993 32747 46065 32803
rect 45993 32713 46012 32747
rect 46046 32713 46065 32747
rect 45993 32657 46065 32713
rect 45993 32623 46012 32657
rect 46046 32623 46065 32657
rect 46883 33268 46955 33324
rect 46883 33234 46902 33268
rect 46936 33234 46955 33268
rect 46883 33178 46955 33234
rect 46883 33144 46902 33178
rect 46936 33144 46955 33178
rect 46883 33088 46955 33144
rect 46883 33054 46902 33088
rect 46936 33054 46955 33088
rect 46883 32998 46955 33054
rect 46883 32964 46902 32998
rect 46936 32964 46955 32998
rect 46883 32908 46955 32964
rect 46883 32874 46902 32908
rect 46936 32874 46955 32908
rect 46883 32818 46955 32874
rect 46883 32784 46902 32818
rect 46936 32784 46955 32818
rect 46883 32728 46955 32784
rect 46883 32694 46902 32728
rect 46936 32694 46955 32728
rect 46883 32638 46955 32694
rect 45993 32563 46065 32623
rect 46883 32604 46902 32638
rect 46936 32604 46955 32638
rect 46883 32563 46955 32604
rect 45993 32544 46955 32563
rect 45993 32510 46090 32544
rect 46124 32510 46180 32544
rect 46214 32510 46270 32544
rect 46304 32510 46360 32544
rect 46394 32510 46450 32544
rect 46484 32510 46540 32544
rect 46574 32510 46630 32544
rect 46664 32510 46720 32544
rect 46754 32510 46810 32544
rect 46844 32510 46955 32544
rect 45993 32491 46955 32510
rect 47333 33434 48295 33453
rect 47333 33400 47464 33434
rect 47498 33400 47554 33434
rect 47588 33400 47644 33434
rect 47678 33400 47734 33434
rect 47768 33400 47824 33434
rect 47858 33400 47914 33434
rect 47948 33400 48004 33434
rect 48038 33400 48094 33434
rect 48128 33400 48184 33434
rect 48218 33400 48295 33434
rect 47333 33381 48295 33400
rect 47333 33377 47405 33381
rect 47333 33343 47352 33377
rect 47386 33343 47405 33377
rect 47333 33287 47405 33343
rect 48223 33358 48295 33381
rect 48223 33324 48242 33358
rect 48276 33324 48295 33358
rect 47333 33253 47352 33287
rect 47386 33253 47405 33287
rect 47333 33197 47405 33253
rect 47333 33163 47352 33197
rect 47386 33163 47405 33197
rect 47333 33107 47405 33163
rect 47333 33073 47352 33107
rect 47386 33073 47405 33107
rect 47333 33017 47405 33073
rect 47333 32983 47352 33017
rect 47386 32983 47405 33017
rect 47333 32927 47405 32983
rect 47333 32893 47352 32927
rect 47386 32893 47405 32927
rect 47333 32837 47405 32893
rect 47333 32803 47352 32837
rect 47386 32803 47405 32837
rect 47333 32747 47405 32803
rect 47333 32713 47352 32747
rect 47386 32713 47405 32747
rect 47333 32657 47405 32713
rect 47333 32623 47352 32657
rect 47386 32623 47405 32657
rect 48223 33268 48295 33324
rect 48223 33234 48242 33268
rect 48276 33234 48295 33268
rect 48223 33178 48295 33234
rect 48223 33144 48242 33178
rect 48276 33144 48295 33178
rect 48223 33088 48295 33144
rect 48223 33054 48242 33088
rect 48276 33054 48295 33088
rect 48223 32998 48295 33054
rect 48223 32964 48242 32998
rect 48276 32964 48295 32998
rect 48223 32908 48295 32964
rect 48223 32874 48242 32908
rect 48276 32874 48295 32908
rect 48223 32818 48295 32874
rect 48223 32784 48242 32818
rect 48276 32784 48295 32818
rect 48223 32728 48295 32784
rect 48223 32694 48242 32728
rect 48276 32694 48295 32728
rect 48223 32638 48295 32694
rect 47333 32563 47405 32623
rect 48223 32604 48242 32638
rect 48276 32604 48295 32638
rect 48223 32563 48295 32604
rect 47333 32544 48295 32563
rect 47333 32510 47430 32544
rect 47464 32510 47520 32544
rect 47554 32510 47610 32544
rect 47644 32510 47700 32544
rect 47734 32510 47790 32544
rect 47824 32510 47880 32544
rect 47914 32510 47970 32544
rect 48004 32510 48060 32544
rect 48094 32510 48150 32544
rect 48184 32510 48295 32544
rect 47333 32491 48295 32510
rect 48673 33434 49635 33453
rect 48673 33400 48804 33434
rect 48838 33400 48894 33434
rect 48928 33400 48984 33434
rect 49018 33400 49074 33434
rect 49108 33400 49164 33434
rect 49198 33400 49254 33434
rect 49288 33400 49344 33434
rect 49378 33400 49434 33434
rect 49468 33400 49524 33434
rect 49558 33400 49635 33434
rect 48673 33381 49635 33400
rect 48673 33377 48745 33381
rect 48673 33343 48692 33377
rect 48726 33343 48745 33377
rect 48673 33287 48745 33343
rect 49563 33358 49635 33381
rect 49563 33324 49582 33358
rect 49616 33324 49635 33358
rect 48673 33253 48692 33287
rect 48726 33253 48745 33287
rect 48673 33197 48745 33253
rect 48673 33163 48692 33197
rect 48726 33163 48745 33197
rect 48673 33107 48745 33163
rect 48673 33073 48692 33107
rect 48726 33073 48745 33107
rect 48673 33017 48745 33073
rect 48673 32983 48692 33017
rect 48726 32983 48745 33017
rect 48673 32927 48745 32983
rect 48673 32893 48692 32927
rect 48726 32893 48745 32927
rect 48673 32837 48745 32893
rect 48673 32803 48692 32837
rect 48726 32803 48745 32837
rect 48673 32747 48745 32803
rect 48673 32713 48692 32747
rect 48726 32713 48745 32747
rect 48673 32657 48745 32713
rect 48673 32623 48692 32657
rect 48726 32623 48745 32657
rect 49563 33268 49635 33324
rect 49563 33234 49582 33268
rect 49616 33234 49635 33268
rect 49563 33178 49635 33234
rect 49563 33144 49582 33178
rect 49616 33144 49635 33178
rect 49563 33088 49635 33144
rect 49563 33054 49582 33088
rect 49616 33054 49635 33088
rect 49563 32998 49635 33054
rect 49563 32964 49582 32998
rect 49616 32964 49635 32998
rect 49563 32908 49635 32964
rect 49563 32874 49582 32908
rect 49616 32874 49635 32908
rect 49563 32818 49635 32874
rect 49563 32784 49582 32818
rect 49616 32784 49635 32818
rect 49563 32728 49635 32784
rect 49563 32694 49582 32728
rect 49616 32694 49635 32728
rect 49563 32638 49635 32694
rect 48673 32563 48745 32623
rect 49563 32604 49582 32638
rect 49616 32604 49635 32638
rect 49563 32563 49635 32604
rect 48673 32544 49635 32563
rect 48673 32510 48770 32544
rect 48804 32510 48860 32544
rect 48894 32510 48950 32544
rect 48984 32510 49040 32544
rect 49074 32510 49130 32544
rect 49164 32510 49220 32544
rect 49254 32510 49310 32544
rect 49344 32510 49400 32544
rect 49434 32510 49490 32544
rect 49524 32510 49635 32544
rect 48673 32491 49635 32510
rect 50013 33434 50975 33453
rect 50013 33400 50144 33434
rect 50178 33400 50234 33434
rect 50268 33400 50324 33434
rect 50358 33400 50414 33434
rect 50448 33400 50504 33434
rect 50538 33400 50594 33434
rect 50628 33400 50684 33434
rect 50718 33400 50774 33434
rect 50808 33400 50864 33434
rect 50898 33400 50975 33434
rect 50013 33381 50975 33400
rect 50013 33377 50085 33381
rect 50013 33343 50032 33377
rect 50066 33343 50085 33377
rect 50013 33287 50085 33343
rect 50903 33358 50975 33381
rect 50903 33324 50922 33358
rect 50956 33324 50975 33358
rect 50013 33253 50032 33287
rect 50066 33253 50085 33287
rect 50013 33197 50085 33253
rect 50013 33163 50032 33197
rect 50066 33163 50085 33197
rect 50013 33107 50085 33163
rect 50013 33073 50032 33107
rect 50066 33073 50085 33107
rect 50013 33017 50085 33073
rect 50013 32983 50032 33017
rect 50066 32983 50085 33017
rect 50013 32927 50085 32983
rect 50013 32893 50032 32927
rect 50066 32893 50085 32927
rect 50013 32837 50085 32893
rect 50013 32803 50032 32837
rect 50066 32803 50085 32837
rect 50013 32747 50085 32803
rect 50013 32713 50032 32747
rect 50066 32713 50085 32747
rect 50013 32657 50085 32713
rect 50013 32623 50032 32657
rect 50066 32623 50085 32657
rect 50903 33268 50975 33324
rect 50903 33234 50922 33268
rect 50956 33234 50975 33268
rect 50903 33178 50975 33234
rect 50903 33144 50922 33178
rect 50956 33144 50975 33178
rect 50903 33088 50975 33144
rect 50903 33054 50922 33088
rect 50956 33054 50975 33088
rect 50903 32998 50975 33054
rect 50903 32964 50922 32998
rect 50956 32964 50975 32998
rect 50903 32908 50975 32964
rect 50903 32874 50922 32908
rect 50956 32874 50975 32908
rect 50903 32818 50975 32874
rect 50903 32784 50922 32818
rect 50956 32784 50975 32818
rect 50903 32728 50975 32784
rect 50903 32694 50922 32728
rect 50956 32694 50975 32728
rect 50903 32638 50975 32694
rect 50013 32563 50085 32623
rect 50903 32604 50922 32638
rect 50956 32604 50975 32638
rect 50903 32563 50975 32604
rect 50013 32544 50975 32563
rect 50013 32510 50110 32544
rect 50144 32510 50200 32544
rect 50234 32510 50290 32544
rect 50324 32510 50380 32544
rect 50414 32510 50470 32544
rect 50504 32510 50560 32544
rect 50594 32510 50650 32544
rect 50684 32510 50740 32544
rect 50774 32510 50830 32544
rect 50864 32510 50975 32544
rect 50013 32491 50975 32510
rect 51353 33434 52315 33453
rect 51353 33400 51484 33434
rect 51518 33400 51574 33434
rect 51608 33400 51664 33434
rect 51698 33400 51754 33434
rect 51788 33400 51844 33434
rect 51878 33400 51934 33434
rect 51968 33400 52024 33434
rect 52058 33400 52114 33434
rect 52148 33400 52204 33434
rect 52238 33400 52315 33434
rect 51353 33381 52315 33400
rect 51353 33377 51425 33381
rect 51353 33343 51372 33377
rect 51406 33343 51425 33377
rect 51353 33287 51425 33343
rect 52243 33358 52315 33381
rect 52243 33324 52262 33358
rect 52296 33324 52315 33358
rect 51353 33253 51372 33287
rect 51406 33253 51425 33287
rect 51353 33197 51425 33253
rect 51353 33163 51372 33197
rect 51406 33163 51425 33197
rect 51353 33107 51425 33163
rect 51353 33073 51372 33107
rect 51406 33073 51425 33107
rect 51353 33017 51425 33073
rect 51353 32983 51372 33017
rect 51406 32983 51425 33017
rect 51353 32927 51425 32983
rect 51353 32893 51372 32927
rect 51406 32893 51425 32927
rect 51353 32837 51425 32893
rect 51353 32803 51372 32837
rect 51406 32803 51425 32837
rect 51353 32747 51425 32803
rect 51353 32713 51372 32747
rect 51406 32713 51425 32747
rect 51353 32657 51425 32713
rect 51353 32623 51372 32657
rect 51406 32623 51425 32657
rect 52243 33268 52315 33324
rect 52243 33234 52262 33268
rect 52296 33234 52315 33268
rect 52243 33178 52315 33234
rect 52243 33144 52262 33178
rect 52296 33144 52315 33178
rect 52243 33088 52315 33144
rect 52243 33054 52262 33088
rect 52296 33054 52315 33088
rect 52243 32998 52315 33054
rect 52243 32964 52262 32998
rect 52296 32964 52315 32998
rect 52243 32908 52315 32964
rect 52243 32874 52262 32908
rect 52296 32874 52315 32908
rect 52243 32818 52315 32874
rect 52243 32784 52262 32818
rect 52296 32784 52315 32818
rect 52243 32728 52315 32784
rect 52243 32694 52262 32728
rect 52296 32694 52315 32728
rect 52243 32638 52315 32694
rect 51353 32563 51425 32623
rect 52243 32604 52262 32638
rect 52296 32604 52315 32638
rect 52243 32563 52315 32604
rect 51353 32544 52315 32563
rect 51353 32510 51450 32544
rect 51484 32510 51540 32544
rect 51574 32510 51630 32544
rect 51664 32510 51720 32544
rect 51754 32510 51810 32544
rect 51844 32510 51900 32544
rect 51934 32510 51990 32544
rect 52024 32510 52080 32544
rect 52114 32510 52170 32544
rect 52204 32510 52315 32544
rect 51353 32491 52315 32510
rect 38470 30079 38590 30082
rect 37412 30029 37452 30072
rect 38470 30045 38515 30079
rect 38549 30045 38590 30079
rect 38470 30042 38590 30045
rect 37412 29995 37415 30029
rect 37449 29995 37452 30029
rect 37412 29952 37452 29995
rect 41973 29674 42935 29693
rect 41973 29640 42104 29674
rect 42138 29640 42194 29674
rect 42228 29640 42284 29674
rect 42318 29640 42374 29674
rect 42408 29640 42464 29674
rect 42498 29640 42554 29674
rect 42588 29640 42644 29674
rect 42678 29640 42734 29674
rect 42768 29640 42824 29674
rect 42858 29640 42935 29674
rect 41973 29621 42935 29640
rect 41973 29617 42045 29621
rect 41973 29583 41992 29617
rect 42026 29583 42045 29617
rect 41973 29527 42045 29583
rect 42863 29598 42935 29621
rect 42863 29564 42882 29598
rect 42916 29564 42935 29598
rect 41973 29493 41992 29527
rect 42026 29493 42045 29527
rect 41973 29437 42045 29493
rect 41973 29403 41992 29437
rect 42026 29403 42045 29437
rect 41973 29347 42045 29403
rect 41973 29313 41992 29347
rect 42026 29313 42045 29347
rect 41973 29257 42045 29313
rect 41973 29223 41992 29257
rect 42026 29223 42045 29257
rect 41973 29167 42045 29223
rect 41973 29133 41992 29167
rect 42026 29133 42045 29167
rect 41973 29077 42045 29133
rect 41973 29043 41992 29077
rect 42026 29043 42045 29077
rect 41973 28987 42045 29043
rect 41973 28953 41992 28987
rect 42026 28953 42045 28987
rect 41973 28897 42045 28953
rect 41973 28863 41992 28897
rect 42026 28863 42045 28897
rect 42863 29508 42935 29564
rect 42863 29474 42882 29508
rect 42916 29474 42935 29508
rect 42863 29418 42935 29474
rect 42863 29384 42882 29418
rect 42916 29384 42935 29418
rect 42863 29328 42935 29384
rect 42863 29294 42882 29328
rect 42916 29294 42935 29328
rect 42863 29238 42935 29294
rect 42863 29204 42882 29238
rect 42916 29204 42935 29238
rect 42863 29148 42935 29204
rect 42863 29114 42882 29148
rect 42916 29114 42935 29148
rect 42863 29058 42935 29114
rect 42863 29024 42882 29058
rect 42916 29024 42935 29058
rect 42863 28968 42935 29024
rect 42863 28934 42882 28968
rect 42916 28934 42935 28968
rect 42863 28878 42935 28934
rect 41973 28803 42045 28863
rect 42863 28844 42882 28878
rect 42916 28844 42935 28878
rect 42863 28803 42935 28844
rect 41973 28784 42935 28803
rect 41973 28750 42070 28784
rect 42104 28750 42160 28784
rect 42194 28750 42250 28784
rect 42284 28750 42340 28784
rect 42374 28750 42430 28784
rect 42464 28750 42520 28784
rect 42554 28750 42610 28784
rect 42644 28750 42700 28784
rect 42734 28750 42790 28784
rect 42824 28750 42935 28784
rect 41973 28731 42935 28750
rect 43313 29674 44275 29693
rect 43313 29640 43444 29674
rect 43478 29640 43534 29674
rect 43568 29640 43624 29674
rect 43658 29640 43714 29674
rect 43748 29640 43804 29674
rect 43838 29640 43894 29674
rect 43928 29640 43984 29674
rect 44018 29640 44074 29674
rect 44108 29640 44164 29674
rect 44198 29640 44275 29674
rect 43313 29621 44275 29640
rect 43313 29617 43385 29621
rect 43313 29583 43332 29617
rect 43366 29583 43385 29617
rect 43313 29527 43385 29583
rect 44203 29598 44275 29621
rect 44203 29564 44222 29598
rect 44256 29564 44275 29598
rect 43313 29493 43332 29527
rect 43366 29493 43385 29527
rect 43313 29437 43385 29493
rect 43313 29403 43332 29437
rect 43366 29403 43385 29437
rect 43313 29347 43385 29403
rect 43313 29313 43332 29347
rect 43366 29313 43385 29347
rect 43313 29257 43385 29313
rect 43313 29223 43332 29257
rect 43366 29223 43385 29257
rect 43313 29167 43385 29223
rect 43313 29133 43332 29167
rect 43366 29133 43385 29167
rect 43313 29077 43385 29133
rect 43313 29043 43332 29077
rect 43366 29043 43385 29077
rect 43313 28987 43385 29043
rect 43313 28953 43332 28987
rect 43366 28953 43385 28987
rect 43313 28897 43385 28953
rect 43313 28863 43332 28897
rect 43366 28863 43385 28897
rect 44203 29508 44275 29564
rect 44203 29474 44222 29508
rect 44256 29474 44275 29508
rect 44203 29418 44275 29474
rect 44203 29384 44222 29418
rect 44256 29384 44275 29418
rect 44203 29328 44275 29384
rect 44203 29294 44222 29328
rect 44256 29294 44275 29328
rect 44203 29238 44275 29294
rect 44203 29204 44222 29238
rect 44256 29204 44275 29238
rect 44203 29148 44275 29204
rect 44203 29114 44222 29148
rect 44256 29114 44275 29148
rect 44203 29058 44275 29114
rect 44203 29024 44222 29058
rect 44256 29024 44275 29058
rect 44203 28968 44275 29024
rect 44203 28934 44222 28968
rect 44256 28934 44275 28968
rect 44203 28878 44275 28934
rect 43313 28803 43385 28863
rect 44203 28844 44222 28878
rect 44256 28844 44275 28878
rect 44203 28803 44275 28844
rect 43313 28784 44275 28803
rect 43313 28750 43410 28784
rect 43444 28750 43500 28784
rect 43534 28750 43590 28784
rect 43624 28750 43680 28784
rect 43714 28750 43770 28784
rect 43804 28750 43860 28784
rect 43894 28750 43950 28784
rect 43984 28750 44040 28784
rect 44074 28750 44130 28784
rect 44164 28750 44275 28784
rect 43313 28731 44275 28750
rect 44653 29674 45615 29693
rect 44653 29640 44784 29674
rect 44818 29640 44874 29674
rect 44908 29640 44964 29674
rect 44998 29640 45054 29674
rect 45088 29640 45144 29674
rect 45178 29640 45234 29674
rect 45268 29640 45324 29674
rect 45358 29640 45414 29674
rect 45448 29640 45504 29674
rect 45538 29640 45615 29674
rect 44653 29621 45615 29640
rect 44653 29617 44725 29621
rect 44653 29583 44672 29617
rect 44706 29583 44725 29617
rect 44653 29527 44725 29583
rect 45543 29598 45615 29621
rect 45543 29564 45562 29598
rect 45596 29564 45615 29598
rect 44653 29493 44672 29527
rect 44706 29493 44725 29527
rect 44653 29437 44725 29493
rect 44653 29403 44672 29437
rect 44706 29403 44725 29437
rect 44653 29347 44725 29403
rect 44653 29313 44672 29347
rect 44706 29313 44725 29347
rect 44653 29257 44725 29313
rect 44653 29223 44672 29257
rect 44706 29223 44725 29257
rect 44653 29167 44725 29223
rect 44653 29133 44672 29167
rect 44706 29133 44725 29167
rect 44653 29077 44725 29133
rect 44653 29043 44672 29077
rect 44706 29043 44725 29077
rect 44653 28987 44725 29043
rect 44653 28953 44672 28987
rect 44706 28953 44725 28987
rect 44653 28897 44725 28953
rect 44653 28863 44672 28897
rect 44706 28863 44725 28897
rect 45543 29508 45615 29564
rect 45543 29474 45562 29508
rect 45596 29474 45615 29508
rect 45543 29418 45615 29474
rect 45543 29384 45562 29418
rect 45596 29384 45615 29418
rect 45543 29328 45615 29384
rect 45543 29294 45562 29328
rect 45596 29294 45615 29328
rect 45543 29238 45615 29294
rect 45543 29204 45562 29238
rect 45596 29204 45615 29238
rect 45543 29148 45615 29204
rect 45543 29114 45562 29148
rect 45596 29114 45615 29148
rect 45543 29058 45615 29114
rect 45543 29024 45562 29058
rect 45596 29024 45615 29058
rect 45543 28968 45615 29024
rect 45543 28934 45562 28968
rect 45596 28934 45615 28968
rect 45543 28878 45615 28934
rect 44653 28803 44725 28863
rect 45543 28844 45562 28878
rect 45596 28844 45615 28878
rect 45543 28803 45615 28844
rect 44653 28784 45615 28803
rect 44653 28750 44750 28784
rect 44784 28750 44840 28784
rect 44874 28750 44930 28784
rect 44964 28750 45020 28784
rect 45054 28750 45110 28784
rect 45144 28750 45200 28784
rect 45234 28750 45290 28784
rect 45324 28750 45380 28784
rect 45414 28750 45470 28784
rect 45504 28750 45615 28784
rect 44653 28731 45615 28750
rect 45993 29674 46955 29693
rect 45993 29640 46124 29674
rect 46158 29640 46214 29674
rect 46248 29640 46304 29674
rect 46338 29640 46394 29674
rect 46428 29640 46484 29674
rect 46518 29640 46574 29674
rect 46608 29640 46664 29674
rect 46698 29640 46754 29674
rect 46788 29640 46844 29674
rect 46878 29640 46955 29674
rect 45993 29621 46955 29640
rect 45993 29617 46065 29621
rect 45993 29583 46012 29617
rect 46046 29583 46065 29617
rect 45993 29527 46065 29583
rect 46883 29598 46955 29621
rect 46883 29564 46902 29598
rect 46936 29564 46955 29598
rect 45993 29493 46012 29527
rect 46046 29493 46065 29527
rect 45993 29437 46065 29493
rect 45993 29403 46012 29437
rect 46046 29403 46065 29437
rect 45993 29347 46065 29403
rect 45993 29313 46012 29347
rect 46046 29313 46065 29347
rect 45993 29257 46065 29313
rect 45993 29223 46012 29257
rect 46046 29223 46065 29257
rect 45993 29167 46065 29223
rect 45993 29133 46012 29167
rect 46046 29133 46065 29167
rect 45993 29077 46065 29133
rect 45993 29043 46012 29077
rect 46046 29043 46065 29077
rect 45993 28987 46065 29043
rect 45993 28953 46012 28987
rect 46046 28953 46065 28987
rect 45993 28897 46065 28953
rect 45993 28863 46012 28897
rect 46046 28863 46065 28897
rect 46883 29508 46955 29564
rect 46883 29474 46902 29508
rect 46936 29474 46955 29508
rect 46883 29418 46955 29474
rect 46883 29384 46902 29418
rect 46936 29384 46955 29418
rect 46883 29328 46955 29384
rect 46883 29294 46902 29328
rect 46936 29294 46955 29328
rect 46883 29238 46955 29294
rect 46883 29204 46902 29238
rect 46936 29204 46955 29238
rect 46883 29148 46955 29204
rect 46883 29114 46902 29148
rect 46936 29114 46955 29148
rect 46883 29058 46955 29114
rect 46883 29024 46902 29058
rect 46936 29024 46955 29058
rect 46883 28968 46955 29024
rect 46883 28934 46902 28968
rect 46936 28934 46955 28968
rect 46883 28878 46955 28934
rect 45993 28803 46065 28863
rect 46883 28844 46902 28878
rect 46936 28844 46955 28878
rect 46883 28803 46955 28844
rect 45993 28784 46955 28803
rect 45993 28750 46090 28784
rect 46124 28750 46180 28784
rect 46214 28750 46270 28784
rect 46304 28750 46360 28784
rect 46394 28750 46450 28784
rect 46484 28750 46540 28784
rect 46574 28750 46630 28784
rect 46664 28750 46720 28784
rect 46754 28750 46810 28784
rect 46844 28750 46955 28784
rect 45993 28731 46955 28750
rect 47333 29674 48295 29693
rect 47333 29640 47464 29674
rect 47498 29640 47554 29674
rect 47588 29640 47644 29674
rect 47678 29640 47734 29674
rect 47768 29640 47824 29674
rect 47858 29640 47914 29674
rect 47948 29640 48004 29674
rect 48038 29640 48094 29674
rect 48128 29640 48184 29674
rect 48218 29640 48295 29674
rect 47333 29621 48295 29640
rect 47333 29617 47405 29621
rect 47333 29583 47352 29617
rect 47386 29583 47405 29617
rect 47333 29527 47405 29583
rect 48223 29598 48295 29621
rect 48223 29564 48242 29598
rect 48276 29564 48295 29598
rect 47333 29493 47352 29527
rect 47386 29493 47405 29527
rect 47333 29437 47405 29493
rect 47333 29403 47352 29437
rect 47386 29403 47405 29437
rect 47333 29347 47405 29403
rect 47333 29313 47352 29347
rect 47386 29313 47405 29347
rect 47333 29257 47405 29313
rect 47333 29223 47352 29257
rect 47386 29223 47405 29257
rect 47333 29167 47405 29223
rect 47333 29133 47352 29167
rect 47386 29133 47405 29167
rect 47333 29077 47405 29133
rect 47333 29043 47352 29077
rect 47386 29043 47405 29077
rect 47333 28987 47405 29043
rect 47333 28953 47352 28987
rect 47386 28953 47405 28987
rect 47333 28897 47405 28953
rect 47333 28863 47352 28897
rect 47386 28863 47405 28897
rect 48223 29508 48295 29564
rect 48223 29474 48242 29508
rect 48276 29474 48295 29508
rect 48223 29418 48295 29474
rect 48223 29384 48242 29418
rect 48276 29384 48295 29418
rect 48223 29328 48295 29384
rect 48223 29294 48242 29328
rect 48276 29294 48295 29328
rect 48223 29238 48295 29294
rect 48223 29204 48242 29238
rect 48276 29204 48295 29238
rect 48223 29148 48295 29204
rect 48223 29114 48242 29148
rect 48276 29114 48295 29148
rect 48223 29058 48295 29114
rect 48223 29024 48242 29058
rect 48276 29024 48295 29058
rect 48223 28968 48295 29024
rect 48223 28934 48242 28968
rect 48276 28934 48295 28968
rect 48223 28878 48295 28934
rect 47333 28803 47405 28863
rect 48223 28844 48242 28878
rect 48276 28844 48295 28878
rect 48223 28803 48295 28844
rect 47333 28784 48295 28803
rect 47333 28750 47430 28784
rect 47464 28750 47520 28784
rect 47554 28750 47610 28784
rect 47644 28750 47700 28784
rect 47734 28750 47790 28784
rect 47824 28750 47880 28784
rect 47914 28750 47970 28784
rect 48004 28750 48060 28784
rect 48094 28750 48150 28784
rect 48184 28750 48295 28784
rect 47333 28731 48295 28750
rect 48673 29674 49635 29693
rect 48673 29640 48804 29674
rect 48838 29640 48894 29674
rect 48928 29640 48984 29674
rect 49018 29640 49074 29674
rect 49108 29640 49164 29674
rect 49198 29640 49254 29674
rect 49288 29640 49344 29674
rect 49378 29640 49434 29674
rect 49468 29640 49524 29674
rect 49558 29640 49635 29674
rect 48673 29621 49635 29640
rect 48673 29617 48745 29621
rect 48673 29583 48692 29617
rect 48726 29583 48745 29617
rect 48673 29527 48745 29583
rect 49563 29598 49635 29621
rect 49563 29564 49582 29598
rect 49616 29564 49635 29598
rect 48673 29493 48692 29527
rect 48726 29493 48745 29527
rect 48673 29437 48745 29493
rect 48673 29403 48692 29437
rect 48726 29403 48745 29437
rect 48673 29347 48745 29403
rect 48673 29313 48692 29347
rect 48726 29313 48745 29347
rect 48673 29257 48745 29313
rect 48673 29223 48692 29257
rect 48726 29223 48745 29257
rect 48673 29167 48745 29223
rect 48673 29133 48692 29167
rect 48726 29133 48745 29167
rect 48673 29077 48745 29133
rect 48673 29043 48692 29077
rect 48726 29043 48745 29077
rect 48673 28987 48745 29043
rect 48673 28953 48692 28987
rect 48726 28953 48745 28987
rect 48673 28897 48745 28953
rect 48673 28863 48692 28897
rect 48726 28863 48745 28897
rect 49563 29508 49635 29564
rect 49563 29474 49582 29508
rect 49616 29474 49635 29508
rect 49563 29418 49635 29474
rect 49563 29384 49582 29418
rect 49616 29384 49635 29418
rect 49563 29328 49635 29384
rect 49563 29294 49582 29328
rect 49616 29294 49635 29328
rect 49563 29238 49635 29294
rect 49563 29204 49582 29238
rect 49616 29204 49635 29238
rect 49563 29148 49635 29204
rect 49563 29114 49582 29148
rect 49616 29114 49635 29148
rect 49563 29058 49635 29114
rect 49563 29024 49582 29058
rect 49616 29024 49635 29058
rect 49563 28968 49635 29024
rect 49563 28934 49582 28968
rect 49616 28934 49635 28968
rect 49563 28878 49635 28934
rect 48673 28803 48745 28863
rect 49563 28844 49582 28878
rect 49616 28844 49635 28878
rect 49563 28803 49635 28844
rect 48673 28784 49635 28803
rect 48673 28750 48770 28784
rect 48804 28750 48860 28784
rect 48894 28750 48950 28784
rect 48984 28750 49040 28784
rect 49074 28750 49130 28784
rect 49164 28750 49220 28784
rect 49254 28750 49310 28784
rect 49344 28750 49400 28784
rect 49434 28750 49490 28784
rect 49524 28750 49635 28784
rect 48673 28731 49635 28750
rect 50013 29674 50975 29693
rect 50013 29640 50144 29674
rect 50178 29640 50234 29674
rect 50268 29640 50324 29674
rect 50358 29640 50414 29674
rect 50448 29640 50504 29674
rect 50538 29640 50594 29674
rect 50628 29640 50684 29674
rect 50718 29640 50774 29674
rect 50808 29640 50864 29674
rect 50898 29640 50975 29674
rect 50013 29621 50975 29640
rect 50013 29617 50085 29621
rect 50013 29583 50032 29617
rect 50066 29583 50085 29617
rect 50013 29527 50085 29583
rect 50903 29598 50975 29621
rect 50903 29564 50922 29598
rect 50956 29564 50975 29598
rect 50013 29493 50032 29527
rect 50066 29493 50085 29527
rect 50013 29437 50085 29493
rect 50013 29403 50032 29437
rect 50066 29403 50085 29437
rect 50013 29347 50085 29403
rect 50013 29313 50032 29347
rect 50066 29313 50085 29347
rect 50013 29257 50085 29313
rect 50013 29223 50032 29257
rect 50066 29223 50085 29257
rect 50013 29167 50085 29223
rect 50013 29133 50032 29167
rect 50066 29133 50085 29167
rect 50013 29077 50085 29133
rect 50013 29043 50032 29077
rect 50066 29043 50085 29077
rect 50013 28987 50085 29043
rect 50013 28953 50032 28987
rect 50066 28953 50085 28987
rect 50013 28897 50085 28953
rect 50013 28863 50032 28897
rect 50066 28863 50085 28897
rect 50903 29508 50975 29564
rect 50903 29474 50922 29508
rect 50956 29474 50975 29508
rect 50903 29418 50975 29474
rect 50903 29384 50922 29418
rect 50956 29384 50975 29418
rect 50903 29328 50975 29384
rect 50903 29294 50922 29328
rect 50956 29294 50975 29328
rect 50903 29238 50975 29294
rect 50903 29204 50922 29238
rect 50956 29204 50975 29238
rect 50903 29148 50975 29204
rect 50903 29114 50922 29148
rect 50956 29114 50975 29148
rect 50903 29058 50975 29114
rect 50903 29024 50922 29058
rect 50956 29024 50975 29058
rect 50903 28968 50975 29024
rect 50903 28934 50922 28968
rect 50956 28934 50975 28968
rect 50903 28878 50975 28934
rect 50013 28803 50085 28863
rect 50903 28844 50922 28878
rect 50956 28844 50975 28878
rect 50903 28803 50975 28844
rect 50013 28784 50975 28803
rect 50013 28750 50110 28784
rect 50144 28750 50200 28784
rect 50234 28750 50290 28784
rect 50324 28750 50380 28784
rect 50414 28750 50470 28784
rect 50504 28750 50560 28784
rect 50594 28750 50650 28784
rect 50684 28750 50740 28784
rect 50774 28750 50830 28784
rect 50864 28750 50975 28784
rect 50013 28731 50975 28750
rect 51353 29674 52315 29693
rect 51353 29640 51484 29674
rect 51518 29640 51574 29674
rect 51608 29640 51664 29674
rect 51698 29640 51754 29674
rect 51788 29640 51844 29674
rect 51878 29640 51934 29674
rect 51968 29640 52024 29674
rect 52058 29640 52114 29674
rect 52148 29640 52204 29674
rect 52238 29640 52315 29674
rect 51353 29621 52315 29640
rect 51353 29617 51425 29621
rect 51353 29583 51372 29617
rect 51406 29583 51425 29617
rect 51353 29527 51425 29583
rect 52243 29598 52315 29621
rect 52243 29564 52262 29598
rect 52296 29564 52315 29598
rect 51353 29493 51372 29527
rect 51406 29493 51425 29527
rect 51353 29437 51425 29493
rect 51353 29403 51372 29437
rect 51406 29403 51425 29437
rect 51353 29347 51425 29403
rect 51353 29313 51372 29347
rect 51406 29313 51425 29347
rect 51353 29257 51425 29313
rect 51353 29223 51372 29257
rect 51406 29223 51425 29257
rect 51353 29167 51425 29223
rect 51353 29133 51372 29167
rect 51406 29133 51425 29167
rect 51353 29077 51425 29133
rect 51353 29043 51372 29077
rect 51406 29043 51425 29077
rect 51353 28987 51425 29043
rect 51353 28953 51372 28987
rect 51406 28953 51425 28987
rect 51353 28897 51425 28953
rect 51353 28863 51372 28897
rect 51406 28863 51425 28897
rect 52243 29508 52315 29564
rect 52243 29474 52262 29508
rect 52296 29474 52315 29508
rect 52243 29418 52315 29474
rect 52243 29384 52262 29418
rect 52296 29384 52315 29418
rect 52243 29328 52315 29384
rect 52243 29294 52262 29328
rect 52296 29294 52315 29328
rect 52243 29238 52315 29294
rect 52243 29204 52262 29238
rect 52296 29204 52315 29238
rect 52243 29148 52315 29204
rect 52243 29114 52262 29148
rect 52296 29114 52315 29148
rect 52243 29058 52315 29114
rect 52243 29024 52262 29058
rect 52296 29024 52315 29058
rect 52243 28968 52315 29024
rect 52243 28934 52262 28968
rect 52296 28934 52315 28968
rect 52243 28878 52315 28934
rect 51353 28803 51425 28863
rect 52243 28844 52262 28878
rect 52296 28844 52315 28878
rect 52243 28803 52315 28844
rect 51353 28784 52315 28803
rect 51353 28750 51450 28784
rect 51484 28750 51540 28784
rect 51574 28750 51630 28784
rect 51664 28750 51720 28784
rect 51754 28750 51810 28784
rect 51844 28750 51900 28784
rect 51934 28750 51990 28784
rect 52024 28750 52080 28784
rect 52114 28750 52170 28784
rect 52204 28750 52315 28784
rect 51353 28731 52315 28750
rect 25828 18799 25948 18802
rect 24770 18749 24810 18792
rect 25828 18765 25873 18799
rect 25907 18765 25948 18799
rect 25828 18762 25948 18765
rect 27128 18799 27248 18802
rect 27128 18765 27173 18799
rect 27207 18765 27248 18799
rect 27128 18762 27248 18765
rect 28428 18799 28548 18802
rect 28428 18765 28473 18799
rect 28507 18765 28548 18799
rect 28428 18762 28548 18765
rect 29728 18799 29848 18802
rect 29728 18765 29773 18799
rect 29807 18765 29848 18799
rect 29728 18762 29848 18765
rect 31028 18799 31148 18802
rect 31028 18765 31073 18799
rect 31107 18765 31148 18799
rect 31028 18762 31148 18765
rect 32328 18799 32448 18802
rect 32328 18765 32373 18799
rect 32407 18765 32448 18799
rect 32328 18762 32448 18765
rect 33628 18799 33748 18802
rect 33628 18765 33673 18799
rect 33707 18765 33748 18799
rect 33628 18762 33748 18765
rect 34928 18799 35048 18802
rect 34928 18765 34973 18799
rect 35007 18765 35048 18799
rect 34928 18762 35048 18765
rect 36228 18799 36348 18802
rect 36228 18765 36273 18799
rect 36307 18765 36348 18799
rect 36228 18762 36348 18765
rect 37528 18799 37648 18802
rect 37528 18765 37573 18799
rect 37607 18765 37648 18799
rect 37528 18762 37648 18765
rect 38828 18799 38948 18802
rect 38828 18765 38873 18799
rect 38907 18765 38948 18799
rect 38828 18762 38948 18765
rect 40128 18799 40248 18802
rect 40128 18765 40173 18799
rect 40207 18765 40248 18799
rect 40128 18762 40248 18765
rect 41428 18799 41548 18802
rect 41428 18765 41473 18799
rect 41507 18765 41548 18799
rect 41428 18762 41548 18765
rect 42728 18799 42848 18802
rect 42728 18765 42773 18799
rect 42807 18765 42848 18799
rect 42728 18762 42848 18765
rect 44028 18799 44148 18802
rect 44028 18765 44073 18799
rect 44107 18765 44148 18799
rect 44028 18762 44148 18765
rect 45328 18799 45448 18802
rect 45328 18765 45373 18799
rect 45407 18765 45448 18799
rect 45328 18762 45448 18765
rect 46628 18799 46748 18802
rect 46628 18765 46673 18799
rect 46707 18765 46748 18799
rect 46628 18762 46748 18765
rect 47928 18799 48048 18802
rect 47928 18765 47973 18799
rect 48007 18765 48048 18799
rect 47928 18762 48048 18765
rect 49228 18799 49348 18802
rect 49228 18765 49273 18799
rect 49307 18765 49348 18799
rect 49228 18762 49348 18765
rect 50528 18799 50648 18802
rect 50528 18765 50573 18799
rect 50607 18765 50648 18799
rect 50528 18762 50648 18765
rect 24770 18715 24773 18749
rect 24807 18715 24810 18749
rect 24770 18672 24810 18715
<< psubdiffcont >>
rect 21831 47901 22273 48003
rect 23861 47195 23895 47229
rect 43020 44804 43054 44838
rect 43116 44827 43150 44861
rect 43206 44827 43240 44861
rect 43296 44827 43330 44861
rect 43386 44827 43420 44861
rect 43476 44827 43510 44861
rect 43566 44827 43600 44861
rect 43656 44827 43690 44861
rect 43746 44827 43780 44861
rect 43836 44827 43870 44861
rect 43926 44827 43960 44861
rect 44016 44827 44050 44861
rect 44106 44827 44140 44861
rect 44207 44804 44241 44838
rect 44360 44804 44394 44838
rect 44456 44827 44490 44861
rect 44546 44827 44580 44861
rect 44636 44827 44670 44861
rect 44726 44827 44760 44861
rect 44816 44827 44850 44861
rect 44906 44827 44940 44861
rect 44996 44827 45030 44861
rect 45086 44827 45120 44861
rect 45176 44827 45210 44861
rect 45266 44827 45300 44861
rect 45356 44827 45390 44861
rect 45446 44827 45480 44861
rect 45547 44804 45581 44838
rect 45700 44804 45734 44838
rect 45796 44827 45830 44861
rect 45886 44827 45920 44861
rect 45976 44827 46010 44861
rect 46066 44827 46100 44861
rect 46156 44827 46190 44861
rect 46246 44827 46280 44861
rect 46336 44827 46370 44861
rect 46426 44827 46460 44861
rect 46516 44827 46550 44861
rect 46606 44827 46640 44861
rect 46696 44827 46730 44861
rect 46786 44827 46820 44861
rect 46887 44804 46921 44838
rect 47040 44804 47074 44838
rect 47136 44827 47170 44861
rect 47226 44827 47260 44861
rect 47316 44827 47350 44861
rect 47406 44827 47440 44861
rect 47496 44827 47530 44861
rect 47586 44827 47620 44861
rect 47676 44827 47710 44861
rect 47766 44827 47800 44861
rect 47856 44827 47890 44861
rect 47946 44827 47980 44861
rect 48036 44827 48070 44861
rect 48126 44827 48160 44861
rect 48227 44804 48261 44838
rect 48380 44804 48414 44838
rect 48476 44827 48510 44861
rect 48566 44827 48600 44861
rect 48656 44827 48690 44861
rect 48746 44827 48780 44861
rect 48836 44827 48870 44861
rect 48926 44827 48960 44861
rect 49016 44827 49050 44861
rect 49106 44827 49140 44861
rect 49196 44827 49230 44861
rect 49286 44827 49320 44861
rect 49376 44827 49410 44861
rect 49466 44827 49500 44861
rect 49567 44804 49601 44838
rect 49720 44804 49754 44838
rect 49816 44827 49850 44861
rect 49906 44827 49940 44861
rect 49996 44827 50030 44861
rect 50086 44827 50120 44861
rect 50176 44827 50210 44861
rect 50266 44827 50300 44861
rect 50356 44827 50390 44861
rect 50446 44827 50480 44861
rect 50536 44827 50570 44861
rect 50626 44827 50660 44861
rect 50716 44827 50750 44861
rect 50806 44827 50840 44861
rect 50907 44804 50941 44838
rect 51060 44804 51094 44838
rect 51156 44827 51190 44861
rect 51246 44827 51280 44861
rect 51336 44827 51370 44861
rect 51426 44827 51460 44861
rect 51516 44827 51550 44861
rect 51606 44827 51640 44861
rect 51696 44827 51730 44861
rect 51786 44827 51820 44861
rect 51876 44827 51910 44861
rect 51966 44827 52000 44861
rect 52056 44827 52090 44861
rect 52146 44827 52180 44861
rect 52247 44804 52281 44838
rect 43020 44714 43054 44748
rect 43020 44624 43054 44658
rect 43020 44534 43054 44568
rect 43020 44444 43054 44478
rect 43020 44354 43054 44388
rect 43020 44264 43054 44298
rect 43020 44174 43054 44208
rect 43020 44084 43054 44118
rect 43020 43994 43054 44028
rect 43020 43904 43054 43938
rect 43020 43814 43054 43848
rect 44207 44714 44241 44748
rect 44360 44714 44394 44748
rect 44207 44624 44241 44658
rect 44360 44624 44394 44658
rect 44207 44534 44241 44568
rect 44360 44534 44394 44568
rect 44207 44444 44241 44478
rect 44360 44444 44394 44478
rect 44207 44354 44241 44388
rect 44360 44354 44394 44388
rect 44207 44264 44241 44298
rect 44360 44264 44394 44298
rect 44207 44174 44241 44208
rect 44360 44174 44394 44208
rect 44207 44084 44241 44118
rect 44360 44084 44394 44118
rect 44207 43994 44241 44028
rect 44360 43994 44394 44028
rect 44207 43904 44241 43938
rect 44360 43904 44394 43938
rect 44207 43814 44241 43848
rect 44360 43814 44394 43848
rect 43020 43724 43054 43758
rect 45547 44714 45581 44748
rect 45700 44714 45734 44748
rect 45547 44624 45581 44658
rect 45700 44624 45734 44658
rect 45547 44534 45581 44568
rect 45700 44534 45734 44568
rect 45547 44444 45581 44478
rect 45700 44444 45734 44478
rect 45547 44354 45581 44388
rect 45700 44354 45734 44388
rect 45547 44264 45581 44298
rect 45700 44264 45734 44298
rect 45547 44174 45581 44208
rect 45700 44174 45734 44208
rect 45547 44084 45581 44118
rect 45700 44084 45734 44118
rect 45547 43994 45581 44028
rect 45700 43994 45734 44028
rect 45547 43904 45581 43938
rect 45700 43904 45734 43938
rect 45547 43814 45581 43848
rect 45700 43814 45734 43848
rect 44207 43724 44241 43758
rect 44360 43724 44394 43758
rect 46887 44714 46921 44748
rect 47040 44714 47074 44748
rect 46887 44624 46921 44658
rect 47040 44624 47074 44658
rect 46887 44534 46921 44568
rect 47040 44534 47074 44568
rect 46887 44444 46921 44478
rect 47040 44444 47074 44478
rect 46887 44354 46921 44388
rect 47040 44354 47074 44388
rect 46887 44264 46921 44298
rect 47040 44264 47074 44298
rect 46887 44174 46921 44208
rect 47040 44174 47074 44208
rect 46887 44084 46921 44118
rect 47040 44084 47074 44118
rect 46887 43994 46921 44028
rect 47040 43994 47074 44028
rect 46887 43904 46921 43938
rect 47040 43904 47074 43938
rect 46887 43814 46921 43848
rect 47040 43814 47074 43848
rect 45547 43724 45581 43758
rect 45700 43724 45734 43758
rect 48227 44714 48261 44748
rect 48380 44714 48414 44748
rect 48227 44624 48261 44658
rect 48380 44624 48414 44658
rect 48227 44534 48261 44568
rect 48380 44534 48414 44568
rect 48227 44444 48261 44478
rect 48380 44444 48414 44478
rect 48227 44354 48261 44388
rect 48380 44354 48414 44388
rect 48227 44264 48261 44298
rect 48380 44264 48414 44298
rect 48227 44174 48261 44208
rect 48380 44174 48414 44208
rect 48227 44084 48261 44118
rect 48380 44084 48414 44118
rect 48227 43994 48261 44028
rect 48380 43994 48414 44028
rect 48227 43904 48261 43938
rect 48380 43904 48414 43938
rect 48227 43814 48261 43848
rect 48380 43814 48414 43848
rect 46887 43724 46921 43758
rect 47040 43724 47074 43758
rect 49567 44714 49601 44748
rect 49720 44714 49754 44748
rect 49567 44624 49601 44658
rect 49720 44624 49754 44658
rect 49567 44534 49601 44568
rect 49720 44534 49754 44568
rect 49567 44444 49601 44478
rect 49720 44444 49754 44478
rect 49567 44354 49601 44388
rect 49720 44354 49754 44388
rect 49567 44264 49601 44298
rect 49720 44264 49754 44298
rect 49567 44174 49601 44208
rect 49720 44174 49754 44208
rect 49567 44084 49601 44118
rect 49720 44084 49754 44118
rect 49567 43994 49601 44028
rect 49720 43994 49754 44028
rect 49567 43904 49601 43938
rect 49720 43904 49754 43938
rect 49567 43814 49601 43848
rect 49720 43814 49754 43848
rect 48227 43724 48261 43758
rect 48380 43724 48414 43758
rect 50907 44714 50941 44748
rect 51060 44714 51094 44748
rect 50907 44624 50941 44658
rect 51060 44624 51094 44658
rect 50907 44534 50941 44568
rect 51060 44534 51094 44568
rect 50907 44444 50941 44478
rect 51060 44444 51094 44478
rect 50907 44354 50941 44388
rect 51060 44354 51094 44388
rect 50907 44264 50941 44298
rect 51060 44264 51094 44298
rect 50907 44174 50941 44208
rect 51060 44174 51094 44208
rect 50907 44084 50941 44118
rect 51060 44084 51094 44118
rect 50907 43994 50941 44028
rect 51060 43994 51094 44028
rect 50907 43904 50941 43938
rect 51060 43904 51094 43938
rect 50907 43814 50941 43848
rect 51060 43814 51094 43848
rect 49567 43724 49601 43758
rect 49720 43724 49754 43758
rect 52247 44714 52281 44748
rect 52247 44624 52281 44658
rect 52247 44534 52281 44568
rect 52247 44444 52281 44478
rect 52247 44354 52281 44388
rect 52247 44264 52281 44298
rect 52247 44174 52281 44208
rect 52247 44084 52281 44118
rect 52247 43994 52281 44028
rect 52247 43904 52281 43938
rect 52247 43814 52281 43848
rect 50907 43724 50941 43758
rect 51060 43724 51094 43758
rect 52247 43724 52281 43758
rect 14061 43435 14095 43469
rect 43116 43640 43150 43674
rect 43206 43640 43240 43674
rect 43296 43640 43330 43674
rect 43386 43640 43420 43674
rect 43476 43640 43510 43674
rect 43566 43640 43600 43674
rect 43656 43640 43690 43674
rect 43746 43640 43780 43674
rect 43836 43640 43870 43674
rect 43926 43640 43960 43674
rect 44016 43640 44050 43674
rect 44106 43640 44140 43674
rect 44456 43640 44490 43674
rect 44546 43640 44580 43674
rect 44636 43640 44670 43674
rect 44726 43640 44760 43674
rect 44816 43640 44850 43674
rect 44906 43640 44940 43674
rect 44996 43640 45030 43674
rect 45086 43640 45120 43674
rect 45176 43640 45210 43674
rect 45266 43640 45300 43674
rect 45356 43640 45390 43674
rect 45446 43640 45480 43674
rect 45796 43640 45830 43674
rect 45886 43640 45920 43674
rect 45976 43640 46010 43674
rect 46066 43640 46100 43674
rect 46156 43640 46190 43674
rect 46246 43640 46280 43674
rect 46336 43640 46370 43674
rect 46426 43640 46460 43674
rect 46516 43640 46550 43674
rect 46606 43640 46640 43674
rect 46696 43640 46730 43674
rect 46786 43640 46820 43674
rect 47136 43640 47170 43674
rect 47226 43640 47260 43674
rect 47316 43640 47350 43674
rect 47406 43640 47440 43674
rect 47496 43640 47530 43674
rect 47586 43640 47620 43674
rect 47676 43640 47710 43674
rect 47766 43640 47800 43674
rect 47856 43640 47890 43674
rect 47946 43640 47980 43674
rect 48036 43640 48070 43674
rect 48126 43640 48160 43674
rect 48476 43640 48510 43674
rect 48566 43640 48600 43674
rect 48656 43640 48690 43674
rect 48746 43640 48780 43674
rect 48836 43640 48870 43674
rect 48926 43640 48960 43674
rect 49016 43640 49050 43674
rect 49106 43640 49140 43674
rect 49196 43640 49230 43674
rect 49286 43640 49320 43674
rect 49376 43640 49410 43674
rect 49466 43640 49500 43674
rect 49816 43640 49850 43674
rect 49906 43640 49940 43674
rect 49996 43640 50030 43674
rect 50086 43640 50120 43674
rect 50176 43640 50210 43674
rect 50266 43640 50300 43674
rect 50356 43640 50390 43674
rect 50446 43640 50480 43674
rect 50536 43640 50570 43674
rect 50626 43640 50660 43674
rect 50716 43640 50750 43674
rect 50806 43640 50840 43674
rect 51156 43640 51190 43674
rect 51246 43640 51280 43674
rect 51336 43640 51370 43674
rect 51426 43640 51460 43674
rect 51516 43640 51550 43674
rect 51606 43640 51640 43674
rect 51696 43640 51730 43674
rect 51786 43640 51820 43674
rect 51876 43640 51910 43674
rect 51966 43640 52000 43674
rect 52056 43640 52090 43674
rect 52146 43640 52180 43674
rect 41844 41044 41878 41078
rect 41940 41067 41974 41101
rect 42030 41067 42064 41101
rect 42120 41067 42154 41101
rect 42210 41067 42244 41101
rect 42300 41067 42334 41101
rect 42390 41067 42424 41101
rect 42480 41067 42514 41101
rect 42570 41067 42604 41101
rect 42660 41067 42694 41101
rect 42750 41067 42784 41101
rect 42840 41067 42874 41101
rect 42930 41067 42964 41101
rect 43031 41044 43065 41078
rect 43184 41044 43218 41078
rect 43280 41067 43314 41101
rect 43370 41067 43404 41101
rect 43460 41067 43494 41101
rect 43550 41067 43584 41101
rect 43640 41067 43674 41101
rect 43730 41067 43764 41101
rect 43820 41067 43854 41101
rect 43910 41067 43944 41101
rect 44000 41067 44034 41101
rect 44090 41067 44124 41101
rect 44180 41067 44214 41101
rect 44270 41067 44304 41101
rect 44371 41044 44405 41078
rect 44524 41044 44558 41078
rect 44620 41067 44654 41101
rect 44710 41067 44744 41101
rect 44800 41067 44834 41101
rect 44890 41067 44924 41101
rect 44980 41067 45014 41101
rect 45070 41067 45104 41101
rect 45160 41067 45194 41101
rect 45250 41067 45284 41101
rect 45340 41067 45374 41101
rect 45430 41067 45464 41101
rect 45520 41067 45554 41101
rect 45610 41067 45644 41101
rect 45711 41044 45745 41078
rect 45864 41044 45898 41078
rect 45960 41067 45994 41101
rect 46050 41067 46084 41101
rect 46140 41067 46174 41101
rect 46230 41067 46264 41101
rect 46320 41067 46354 41101
rect 46410 41067 46444 41101
rect 46500 41067 46534 41101
rect 46590 41067 46624 41101
rect 46680 41067 46714 41101
rect 46770 41067 46804 41101
rect 46860 41067 46894 41101
rect 46950 41067 46984 41101
rect 47051 41044 47085 41078
rect 47204 41044 47238 41078
rect 47300 41067 47334 41101
rect 47390 41067 47424 41101
rect 47480 41067 47514 41101
rect 47570 41067 47604 41101
rect 47660 41067 47694 41101
rect 47750 41067 47784 41101
rect 47840 41067 47874 41101
rect 47930 41067 47964 41101
rect 48020 41067 48054 41101
rect 48110 41067 48144 41101
rect 48200 41067 48234 41101
rect 48290 41067 48324 41101
rect 48391 41044 48425 41078
rect 48544 41044 48578 41078
rect 48640 41067 48674 41101
rect 48730 41067 48764 41101
rect 48820 41067 48854 41101
rect 48910 41067 48944 41101
rect 49000 41067 49034 41101
rect 49090 41067 49124 41101
rect 49180 41067 49214 41101
rect 49270 41067 49304 41101
rect 49360 41067 49394 41101
rect 49450 41067 49484 41101
rect 49540 41067 49574 41101
rect 49630 41067 49664 41101
rect 49731 41044 49765 41078
rect 49884 41044 49918 41078
rect 49980 41067 50014 41101
rect 50070 41067 50104 41101
rect 50160 41067 50194 41101
rect 50250 41067 50284 41101
rect 50340 41067 50374 41101
rect 50430 41067 50464 41101
rect 50520 41067 50554 41101
rect 50610 41067 50644 41101
rect 50700 41067 50734 41101
rect 50790 41067 50824 41101
rect 50880 41067 50914 41101
rect 50970 41067 51004 41101
rect 51071 41044 51105 41078
rect 51224 41044 51258 41078
rect 51320 41067 51354 41101
rect 51410 41067 51444 41101
rect 51500 41067 51534 41101
rect 51590 41067 51624 41101
rect 51680 41067 51714 41101
rect 51770 41067 51804 41101
rect 51860 41067 51894 41101
rect 51950 41067 51984 41101
rect 52040 41067 52074 41101
rect 52130 41067 52164 41101
rect 52220 41067 52254 41101
rect 52310 41067 52344 41101
rect 52411 41044 52445 41078
rect 41844 40954 41878 40988
rect 41844 40864 41878 40898
rect 41844 40774 41878 40808
rect 41844 40684 41878 40718
rect 41844 40594 41878 40628
rect 41844 40504 41878 40538
rect 41844 40414 41878 40448
rect 41844 40324 41878 40358
rect 41844 40234 41878 40268
rect 41844 40144 41878 40178
rect 41844 40054 41878 40088
rect 43031 40954 43065 40988
rect 43184 40954 43218 40988
rect 43031 40864 43065 40898
rect 43184 40864 43218 40898
rect 43031 40774 43065 40808
rect 43184 40774 43218 40808
rect 43031 40684 43065 40718
rect 43184 40684 43218 40718
rect 43031 40594 43065 40628
rect 43184 40594 43218 40628
rect 43031 40504 43065 40538
rect 43184 40504 43218 40538
rect 43031 40414 43065 40448
rect 43184 40414 43218 40448
rect 43031 40324 43065 40358
rect 43184 40324 43218 40358
rect 43031 40234 43065 40268
rect 43184 40234 43218 40268
rect 43031 40144 43065 40178
rect 43184 40144 43218 40178
rect 43031 40054 43065 40088
rect 43184 40054 43218 40088
rect 41844 39964 41878 39998
rect 44371 40954 44405 40988
rect 44524 40954 44558 40988
rect 44371 40864 44405 40898
rect 44524 40864 44558 40898
rect 44371 40774 44405 40808
rect 44524 40774 44558 40808
rect 44371 40684 44405 40718
rect 44524 40684 44558 40718
rect 44371 40594 44405 40628
rect 44524 40594 44558 40628
rect 44371 40504 44405 40538
rect 44524 40504 44558 40538
rect 44371 40414 44405 40448
rect 44524 40414 44558 40448
rect 44371 40324 44405 40358
rect 44524 40324 44558 40358
rect 44371 40234 44405 40268
rect 44524 40234 44558 40268
rect 44371 40144 44405 40178
rect 44524 40144 44558 40178
rect 44371 40054 44405 40088
rect 44524 40054 44558 40088
rect 43031 39964 43065 39998
rect 43184 39964 43218 39998
rect 45711 40954 45745 40988
rect 45864 40954 45898 40988
rect 45711 40864 45745 40898
rect 45864 40864 45898 40898
rect 45711 40774 45745 40808
rect 45864 40774 45898 40808
rect 45711 40684 45745 40718
rect 45864 40684 45898 40718
rect 45711 40594 45745 40628
rect 45864 40594 45898 40628
rect 45711 40504 45745 40538
rect 45864 40504 45898 40538
rect 45711 40414 45745 40448
rect 45864 40414 45898 40448
rect 45711 40324 45745 40358
rect 45864 40324 45898 40358
rect 45711 40234 45745 40268
rect 45864 40234 45898 40268
rect 45711 40144 45745 40178
rect 45864 40144 45898 40178
rect 45711 40054 45745 40088
rect 45864 40054 45898 40088
rect 44371 39964 44405 39998
rect 44524 39964 44558 39998
rect 47051 40954 47085 40988
rect 47204 40954 47238 40988
rect 47051 40864 47085 40898
rect 47204 40864 47238 40898
rect 47051 40774 47085 40808
rect 47204 40774 47238 40808
rect 47051 40684 47085 40718
rect 47204 40684 47238 40718
rect 47051 40594 47085 40628
rect 47204 40594 47238 40628
rect 47051 40504 47085 40538
rect 47204 40504 47238 40538
rect 47051 40414 47085 40448
rect 47204 40414 47238 40448
rect 47051 40324 47085 40358
rect 47204 40324 47238 40358
rect 47051 40234 47085 40268
rect 47204 40234 47238 40268
rect 47051 40144 47085 40178
rect 47204 40144 47238 40178
rect 47051 40054 47085 40088
rect 47204 40054 47238 40088
rect 45711 39964 45745 39998
rect 45864 39964 45898 39998
rect 48391 40954 48425 40988
rect 48544 40954 48578 40988
rect 48391 40864 48425 40898
rect 48544 40864 48578 40898
rect 48391 40774 48425 40808
rect 48544 40774 48578 40808
rect 48391 40684 48425 40718
rect 48544 40684 48578 40718
rect 48391 40594 48425 40628
rect 48544 40594 48578 40628
rect 48391 40504 48425 40538
rect 48544 40504 48578 40538
rect 48391 40414 48425 40448
rect 48544 40414 48578 40448
rect 48391 40324 48425 40358
rect 48544 40324 48578 40358
rect 48391 40234 48425 40268
rect 48544 40234 48578 40268
rect 48391 40144 48425 40178
rect 48544 40144 48578 40178
rect 48391 40054 48425 40088
rect 48544 40054 48578 40088
rect 47051 39964 47085 39998
rect 47204 39964 47238 39998
rect 49731 40954 49765 40988
rect 49884 40954 49918 40988
rect 49731 40864 49765 40898
rect 49884 40864 49918 40898
rect 49731 40774 49765 40808
rect 49884 40774 49918 40808
rect 49731 40684 49765 40718
rect 49884 40684 49918 40718
rect 49731 40594 49765 40628
rect 49884 40594 49918 40628
rect 49731 40504 49765 40538
rect 49884 40504 49918 40538
rect 49731 40414 49765 40448
rect 49884 40414 49918 40448
rect 49731 40324 49765 40358
rect 49884 40324 49918 40358
rect 49731 40234 49765 40268
rect 49884 40234 49918 40268
rect 49731 40144 49765 40178
rect 49884 40144 49918 40178
rect 49731 40054 49765 40088
rect 49884 40054 49918 40088
rect 48391 39964 48425 39998
rect 48544 39964 48578 39998
rect 51071 40954 51105 40988
rect 51224 40954 51258 40988
rect 51071 40864 51105 40898
rect 51224 40864 51258 40898
rect 51071 40774 51105 40808
rect 51224 40774 51258 40808
rect 51071 40684 51105 40718
rect 51224 40684 51258 40718
rect 51071 40594 51105 40628
rect 51224 40594 51258 40628
rect 51071 40504 51105 40538
rect 51224 40504 51258 40538
rect 51071 40414 51105 40448
rect 51224 40414 51258 40448
rect 51071 40324 51105 40358
rect 51224 40324 51258 40358
rect 51071 40234 51105 40268
rect 51224 40234 51258 40268
rect 51071 40144 51105 40178
rect 51224 40144 51258 40178
rect 51071 40054 51105 40088
rect 51224 40054 51258 40088
rect 49731 39964 49765 39998
rect 49884 39964 49918 39998
rect 52411 40954 52445 40988
rect 52411 40864 52445 40898
rect 52411 40774 52445 40808
rect 52411 40684 52445 40718
rect 52411 40594 52445 40628
rect 52411 40504 52445 40538
rect 52411 40414 52445 40448
rect 52411 40324 52445 40358
rect 52411 40234 52445 40268
rect 52411 40144 52445 40178
rect 52411 40054 52445 40088
rect 51071 39964 51105 39998
rect 51224 39964 51258 39998
rect 52411 39964 52445 39998
rect 41940 39880 41974 39914
rect 42030 39880 42064 39914
rect 42120 39880 42154 39914
rect 42210 39880 42244 39914
rect 42300 39880 42334 39914
rect 42390 39880 42424 39914
rect 42480 39880 42514 39914
rect 42570 39880 42604 39914
rect 42660 39880 42694 39914
rect 42750 39880 42784 39914
rect 42840 39880 42874 39914
rect 42930 39880 42964 39914
rect 43280 39880 43314 39914
rect 43370 39880 43404 39914
rect 43460 39880 43494 39914
rect 43550 39880 43584 39914
rect 43640 39880 43674 39914
rect 43730 39880 43764 39914
rect 43820 39880 43854 39914
rect 43910 39880 43944 39914
rect 44000 39880 44034 39914
rect 44090 39880 44124 39914
rect 44180 39880 44214 39914
rect 44270 39880 44304 39914
rect 44620 39880 44654 39914
rect 44710 39880 44744 39914
rect 44800 39880 44834 39914
rect 44890 39880 44924 39914
rect 44980 39880 45014 39914
rect 45070 39880 45104 39914
rect 45160 39880 45194 39914
rect 45250 39880 45284 39914
rect 45340 39880 45374 39914
rect 45430 39880 45464 39914
rect 45520 39880 45554 39914
rect 45610 39880 45644 39914
rect 45960 39880 45994 39914
rect 46050 39880 46084 39914
rect 46140 39880 46174 39914
rect 46230 39880 46264 39914
rect 46320 39880 46354 39914
rect 46410 39880 46444 39914
rect 46500 39880 46534 39914
rect 46590 39880 46624 39914
rect 46680 39880 46714 39914
rect 46770 39880 46804 39914
rect 46860 39880 46894 39914
rect 46950 39880 46984 39914
rect 47300 39880 47334 39914
rect 47390 39880 47424 39914
rect 47480 39880 47514 39914
rect 47570 39880 47604 39914
rect 47660 39880 47694 39914
rect 47750 39880 47784 39914
rect 47840 39880 47874 39914
rect 47930 39880 47964 39914
rect 48020 39880 48054 39914
rect 48110 39880 48144 39914
rect 48200 39880 48234 39914
rect 48290 39880 48324 39914
rect 48640 39880 48674 39914
rect 48730 39880 48764 39914
rect 48820 39880 48854 39914
rect 48910 39880 48944 39914
rect 49000 39880 49034 39914
rect 49090 39880 49124 39914
rect 49180 39880 49214 39914
rect 49270 39880 49304 39914
rect 49360 39880 49394 39914
rect 49450 39880 49484 39914
rect 49540 39880 49574 39914
rect 49630 39880 49664 39914
rect 49980 39880 50014 39914
rect 50070 39880 50104 39914
rect 50160 39880 50194 39914
rect 50250 39880 50284 39914
rect 50340 39880 50374 39914
rect 50430 39880 50464 39914
rect 50520 39880 50554 39914
rect 50610 39880 50644 39914
rect 50700 39880 50734 39914
rect 50790 39880 50824 39914
rect 50880 39880 50914 39914
rect 50970 39880 51004 39914
rect 51320 39880 51354 39914
rect 51410 39880 51444 39914
rect 51500 39880 51534 39914
rect 51590 39880 51624 39914
rect 51680 39880 51714 39914
rect 51770 39880 51804 39914
rect 51860 39880 51894 39914
rect 51950 39880 51984 39914
rect 52040 39880 52074 39914
rect 52130 39880 52164 39914
rect 52220 39880 52254 39914
rect 52310 39880 52344 39914
rect 37219 39675 37253 39709
rect 38321 39645 38355 39679
rect 39621 39645 39655 39679
rect 12052 37284 12086 37318
rect 12148 37307 12182 37341
rect 12238 37307 12272 37341
rect 12328 37307 12362 37341
rect 12418 37307 12452 37341
rect 12508 37307 12542 37341
rect 12598 37307 12632 37341
rect 12688 37307 12722 37341
rect 12778 37307 12812 37341
rect 12868 37307 12902 37341
rect 12958 37307 12992 37341
rect 13048 37307 13082 37341
rect 13138 37307 13172 37341
rect 13239 37284 13273 37318
rect 12052 37194 12086 37228
rect 12052 37104 12086 37138
rect 12052 37014 12086 37048
rect 12052 36924 12086 36958
rect 12052 36834 12086 36868
rect 12052 36744 12086 36778
rect 12052 36654 12086 36688
rect 12052 36564 12086 36598
rect 12052 36474 12086 36508
rect 12052 36384 12086 36418
rect 12052 36294 12086 36328
rect 13239 37194 13273 37228
rect 13239 37104 13273 37138
rect 13239 37014 13273 37048
rect 13239 36924 13273 36958
rect 13239 36834 13273 36868
rect 13239 36744 13273 36778
rect 13239 36654 13273 36688
rect 13239 36564 13273 36598
rect 14677 36621 15119 36723
rect 17421 36621 17863 36723
rect 20453 36621 20895 36723
rect 23497 36621 23939 36723
rect 13239 36474 13273 36508
rect 13239 36384 13273 36418
rect 13239 36294 13273 36328
rect 12052 36204 12086 36238
rect 13239 36204 13273 36238
rect 12148 36120 12182 36154
rect 12238 36120 12272 36154
rect 12328 36120 12362 36154
rect 12418 36120 12452 36154
rect 12508 36120 12542 36154
rect 12598 36120 12632 36154
rect 12688 36120 12722 36154
rect 12778 36120 12812 36154
rect 12868 36120 12902 36154
rect 12958 36120 12992 36154
rect 13048 36120 13082 36154
rect 13138 36120 13172 36154
rect 41844 37284 41878 37318
rect 41940 37307 41974 37341
rect 42030 37307 42064 37341
rect 42120 37307 42154 37341
rect 42210 37307 42244 37341
rect 42300 37307 42334 37341
rect 42390 37307 42424 37341
rect 42480 37307 42514 37341
rect 42570 37307 42604 37341
rect 42660 37307 42694 37341
rect 42750 37307 42784 37341
rect 42840 37307 42874 37341
rect 42930 37307 42964 37341
rect 43031 37284 43065 37318
rect 43184 37284 43218 37318
rect 43280 37307 43314 37341
rect 43370 37307 43404 37341
rect 43460 37307 43494 37341
rect 43550 37307 43584 37341
rect 43640 37307 43674 37341
rect 43730 37307 43764 37341
rect 43820 37307 43854 37341
rect 43910 37307 43944 37341
rect 44000 37307 44034 37341
rect 44090 37307 44124 37341
rect 44180 37307 44214 37341
rect 44270 37307 44304 37341
rect 44371 37284 44405 37318
rect 44524 37284 44558 37318
rect 44620 37307 44654 37341
rect 44710 37307 44744 37341
rect 44800 37307 44834 37341
rect 44890 37307 44924 37341
rect 44980 37307 45014 37341
rect 45070 37307 45104 37341
rect 45160 37307 45194 37341
rect 45250 37307 45284 37341
rect 45340 37307 45374 37341
rect 45430 37307 45464 37341
rect 45520 37307 45554 37341
rect 45610 37307 45644 37341
rect 45711 37284 45745 37318
rect 45864 37284 45898 37318
rect 45960 37307 45994 37341
rect 46050 37307 46084 37341
rect 46140 37307 46174 37341
rect 46230 37307 46264 37341
rect 46320 37307 46354 37341
rect 46410 37307 46444 37341
rect 46500 37307 46534 37341
rect 46590 37307 46624 37341
rect 46680 37307 46714 37341
rect 46770 37307 46804 37341
rect 46860 37307 46894 37341
rect 46950 37307 46984 37341
rect 47051 37284 47085 37318
rect 47204 37284 47238 37318
rect 47300 37307 47334 37341
rect 47390 37307 47424 37341
rect 47480 37307 47514 37341
rect 47570 37307 47604 37341
rect 47660 37307 47694 37341
rect 47750 37307 47784 37341
rect 47840 37307 47874 37341
rect 47930 37307 47964 37341
rect 48020 37307 48054 37341
rect 48110 37307 48144 37341
rect 48200 37307 48234 37341
rect 48290 37307 48324 37341
rect 48391 37284 48425 37318
rect 48544 37284 48578 37318
rect 48640 37307 48674 37341
rect 48730 37307 48764 37341
rect 48820 37307 48854 37341
rect 48910 37307 48944 37341
rect 49000 37307 49034 37341
rect 49090 37307 49124 37341
rect 49180 37307 49214 37341
rect 49270 37307 49304 37341
rect 49360 37307 49394 37341
rect 49450 37307 49484 37341
rect 49540 37307 49574 37341
rect 49630 37307 49664 37341
rect 49731 37284 49765 37318
rect 49884 37284 49918 37318
rect 49980 37307 50014 37341
rect 50070 37307 50104 37341
rect 50160 37307 50194 37341
rect 50250 37307 50284 37341
rect 50340 37307 50374 37341
rect 50430 37307 50464 37341
rect 50520 37307 50554 37341
rect 50610 37307 50644 37341
rect 50700 37307 50734 37341
rect 50790 37307 50824 37341
rect 50880 37307 50914 37341
rect 50970 37307 51004 37341
rect 51071 37284 51105 37318
rect 51224 37284 51258 37318
rect 51320 37307 51354 37341
rect 51410 37307 51444 37341
rect 51500 37307 51534 37341
rect 51590 37307 51624 37341
rect 51680 37307 51714 37341
rect 51770 37307 51804 37341
rect 51860 37307 51894 37341
rect 51950 37307 51984 37341
rect 52040 37307 52074 37341
rect 52130 37307 52164 37341
rect 52220 37307 52254 37341
rect 52310 37307 52344 37341
rect 52411 37284 52445 37318
rect 41844 37194 41878 37228
rect 41844 37104 41878 37138
rect 41844 37014 41878 37048
rect 41844 36924 41878 36958
rect 41844 36834 41878 36868
rect 41844 36744 41878 36778
rect 41844 36654 41878 36688
rect 41844 36564 41878 36598
rect 41844 36474 41878 36508
rect 41844 36384 41878 36418
rect 41844 36294 41878 36328
rect 43031 37194 43065 37228
rect 43184 37194 43218 37228
rect 43031 37104 43065 37138
rect 43184 37104 43218 37138
rect 43031 37014 43065 37048
rect 43184 37014 43218 37048
rect 43031 36924 43065 36958
rect 43184 36924 43218 36958
rect 43031 36834 43065 36868
rect 43184 36834 43218 36868
rect 43031 36744 43065 36778
rect 43184 36744 43218 36778
rect 43031 36654 43065 36688
rect 43184 36654 43218 36688
rect 43031 36564 43065 36598
rect 43184 36564 43218 36598
rect 43031 36474 43065 36508
rect 43184 36474 43218 36508
rect 43031 36384 43065 36418
rect 43184 36384 43218 36418
rect 43031 36294 43065 36328
rect 43184 36294 43218 36328
rect 41844 36204 41878 36238
rect 44371 37194 44405 37228
rect 44524 37194 44558 37228
rect 44371 37104 44405 37138
rect 44524 37104 44558 37138
rect 44371 37014 44405 37048
rect 44524 37014 44558 37048
rect 44371 36924 44405 36958
rect 44524 36924 44558 36958
rect 44371 36834 44405 36868
rect 44524 36834 44558 36868
rect 44371 36744 44405 36778
rect 44524 36744 44558 36778
rect 44371 36654 44405 36688
rect 44524 36654 44558 36688
rect 44371 36564 44405 36598
rect 44524 36564 44558 36598
rect 44371 36474 44405 36508
rect 44524 36474 44558 36508
rect 44371 36384 44405 36418
rect 44524 36384 44558 36418
rect 44371 36294 44405 36328
rect 44524 36294 44558 36328
rect 43031 36204 43065 36238
rect 43184 36204 43218 36238
rect 45711 37194 45745 37228
rect 45864 37194 45898 37228
rect 45711 37104 45745 37138
rect 45864 37104 45898 37138
rect 45711 37014 45745 37048
rect 45864 37014 45898 37048
rect 45711 36924 45745 36958
rect 45864 36924 45898 36958
rect 45711 36834 45745 36868
rect 45864 36834 45898 36868
rect 45711 36744 45745 36778
rect 45864 36744 45898 36778
rect 45711 36654 45745 36688
rect 45864 36654 45898 36688
rect 45711 36564 45745 36598
rect 45864 36564 45898 36598
rect 45711 36474 45745 36508
rect 45864 36474 45898 36508
rect 45711 36384 45745 36418
rect 45864 36384 45898 36418
rect 45711 36294 45745 36328
rect 45864 36294 45898 36328
rect 44371 36204 44405 36238
rect 44524 36204 44558 36238
rect 47051 37194 47085 37228
rect 47204 37194 47238 37228
rect 47051 37104 47085 37138
rect 47204 37104 47238 37138
rect 47051 37014 47085 37048
rect 47204 37014 47238 37048
rect 47051 36924 47085 36958
rect 47204 36924 47238 36958
rect 47051 36834 47085 36868
rect 47204 36834 47238 36868
rect 47051 36744 47085 36778
rect 47204 36744 47238 36778
rect 47051 36654 47085 36688
rect 47204 36654 47238 36688
rect 47051 36564 47085 36598
rect 47204 36564 47238 36598
rect 47051 36474 47085 36508
rect 47204 36474 47238 36508
rect 47051 36384 47085 36418
rect 47204 36384 47238 36418
rect 47051 36294 47085 36328
rect 47204 36294 47238 36328
rect 45711 36204 45745 36238
rect 45864 36204 45898 36238
rect 48391 37194 48425 37228
rect 48544 37194 48578 37228
rect 48391 37104 48425 37138
rect 48544 37104 48578 37138
rect 48391 37014 48425 37048
rect 48544 37014 48578 37048
rect 48391 36924 48425 36958
rect 48544 36924 48578 36958
rect 48391 36834 48425 36868
rect 48544 36834 48578 36868
rect 48391 36744 48425 36778
rect 48544 36744 48578 36778
rect 48391 36654 48425 36688
rect 48544 36654 48578 36688
rect 48391 36564 48425 36598
rect 48544 36564 48578 36598
rect 48391 36474 48425 36508
rect 48544 36474 48578 36508
rect 48391 36384 48425 36418
rect 48544 36384 48578 36418
rect 48391 36294 48425 36328
rect 48544 36294 48578 36328
rect 47051 36204 47085 36238
rect 47204 36204 47238 36238
rect 49731 37194 49765 37228
rect 49884 37194 49918 37228
rect 49731 37104 49765 37138
rect 49884 37104 49918 37138
rect 49731 37014 49765 37048
rect 49884 37014 49918 37048
rect 49731 36924 49765 36958
rect 49884 36924 49918 36958
rect 49731 36834 49765 36868
rect 49884 36834 49918 36868
rect 49731 36744 49765 36778
rect 49884 36744 49918 36778
rect 49731 36654 49765 36688
rect 49884 36654 49918 36688
rect 49731 36564 49765 36598
rect 49884 36564 49918 36598
rect 49731 36474 49765 36508
rect 49884 36474 49918 36508
rect 49731 36384 49765 36418
rect 49884 36384 49918 36418
rect 49731 36294 49765 36328
rect 49884 36294 49918 36328
rect 48391 36204 48425 36238
rect 48544 36204 48578 36238
rect 51071 37194 51105 37228
rect 51224 37194 51258 37228
rect 51071 37104 51105 37138
rect 51224 37104 51258 37138
rect 51071 37014 51105 37048
rect 51224 37014 51258 37048
rect 51071 36924 51105 36958
rect 51224 36924 51258 36958
rect 51071 36834 51105 36868
rect 51224 36834 51258 36868
rect 51071 36744 51105 36778
rect 51224 36744 51258 36778
rect 51071 36654 51105 36688
rect 51224 36654 51258 36688
rect 51071 36564 51105 36598
rect 51224 36564 51258 36598
rect 51071 36474 51105 36508
rect 51224 36474 51258 36508
rect 51071 36384 51105 36418
rect 51224 36384 51258 36418
rect 51071 36294 51105 36328
rect 51224 36294 51258 36328
rect 49731 36204 49765 36238
rect 49884 36204 49918 36238
rect 52411 37194 52445 37228
rect 52411 37104 52445 37138
rect 52411 37014 52445 37048
rect 52411 36924 52445 36958
rect 52411 36834 52445 36868
rect 52411 36744 52445 36778
rect 52411 36654 52445 36688
rect 52411 36564 52445 36598
rect 52411 36474 52445 36508
rect 52411 36384 52445 36418
rect 52411 36294 52445 36328
rect 51071 36204 51105 36238
rect 51224 36204 51258 36238
rect 52411 36204 52445 36238
rect 41940 36120 41974 36154
rect 42030 36120 42064 36154
rect 42120 36120 42154 36154
rect 42210 36120 42244 36154
rect 42300 36120 42334 36154
rect 42390 36120 42424 36154
rect 42480 36120 42514 36154
rect 42570 36120 42604 36154
rect 42660 36120 42694 36154
rect 42750 36120 42784 36154
rect 42840 36120 42874 36154
rect 42930 36120 42964 36154
rect 43280 36120 43314 36154
rect 43370 36120 43404 36154
rect 43460 36120 43494 36154
rect 43550 36120 43584 36154
rect 43640 36120 43674 36154
rect 43730 36120 43764 36154
rect 43820 36120 43854 36154
rect 43910 36120 43944 36154
rect 44000 36120 44034 36154
rect 44090 36120 44124 36154
rect 44180 36120 44214 36154
rect 44270 36120 44304 36154
rect 44620 36120 44654 36154
rect 44710 36120 44744 36154
rect 44800 36120 44834 36154
rect 44890 36120 44924 36154
rect 44980 36120 45014 36154
rect 45070 36120 45104 36154
rect 45160 36120 45194 36154
rect 45250 36120 45284 36154
rect 45340 36120 45374 36154
rect 45430 36120 45464 36154
rect 45520 36120 45554 36154
rect 45610 36120 45644 36154
rect 45960 36120 45994 36154
rect 46050 36120 46084 36154
rect 46140 36120 46174 36154
rect 46230 36120 46264 36154
rect 46320 36120 46354 36154
rect 46410 36120 46444 36154
rect 46500 36120 46534 36154
rect 46590 36120 46624 36154
rect 46680 36120 46714 36154
rect 46770 36120 46804 36154
rect 46860 36120 46894 36154
rect 46950 36120 46984 36154
rect 47300 36120 47334 36154
rect 47390 36120 47424 36154
rect 47480 36120 47514 36154
rect 47570 36120 47604 36154
rect 47660 36120 47694 36154
rect 47750 36120 47784 36154
rect 47840 36120 47874 36154
rect 47930 36120 47964 36154
rect 48020 36120 48054 36154
rect 48110 36120 48144 36154
rect 48200 36120 48234 36154
rect 48290 36120 48324 36154
rect 48640 36120 48674 36154
rect 48730 36120 48764 36154
rect 48820 36120 48854 36154
rect 48910 36120 48944 36154
rect 49000 36120 49034 36154
rect 49090 36120 49124 36154
rect 49180 36120 49214 36154
rect 49270 36120 49304 36154
rect 49360 36120 49394 36154
rect 49450 36120 49484 36154
rect 49540 36120 49574 36154
rect 49630 36120 49664 36154
rect 49980 36120 50014 36154
rect 50070 36120 50104 36154
rect 50160 36120 50194 36154
rect 50250 36120 50284 36154
rect 50340 36120 50374 36154
rect 50430 36120 50464 36154
rect 50520 36120 50554 36154
rect 50610 36120 50644 36154
rect 50700 36120 50734 36154
rect 50790 36120 50824 36154
rect 50880 36120 50914 36154
rect 50970 36120 51004 36154
rect 51320 36120 51354 36154
rect 51410 36120 51444 36154
rect 51500 36120 51534 36154
rect 51590 36120 51624 36154
rect 51680 36120 51714 36154
rect 51770 36120 51804 36154
rect 51860 36120 51894 36154
rect 51950 36120 51984 36154
rect 52040 36120 52074 36154
rect 52130 36120 52164 36154
rect 52220 36120 52254 36154
rect 52310 36120 52344 36154
rect 25361 35915 25395 35949
rect 26463 35885 26497 35919
rect 27763 35885 27797 35919
rect 41844 33524 41878 33558
rect 41940 33547 41974 33581
rect 42030 33547 42064 33581
rect 42120 33547 42154 33581
rect 42210 33547 42244 33581
rect 42300 33547 42334 33581
rect 42390 33547 42424 33581
rect 42480 33547 42514 33581
rect 42570 33547 42604 33581
rect 42660 33547 42694 33581
rect 42750 33547 42784 33581
rect 42840 33547 42874 33581
rect 42930 33547 42964 33581
rect 43031 33524 43065 33558
rect 43184 33524 43218 33558
rect 43280 33547 43314 33581
rect 43370 33547 43404 33581
rect 43460 33547 43494 33581
rect 43550 33547 43584 33581
rect 43640 33547 43674 33581
rect 43730 33547 43764 33581
rect 43820 33547 43854 33581
rect 43910 33547 43944 33581
rect 44000 33547 44034 33581
rect 44090 33547 44124 33581
rect 44180 33547 44214 33581
rect 44270 33547 44304 33581
rect 44371 33524 44405 33558
rect 44524 33524 44558 33558
rect 44620 33547 44654 33581
rect 44710 33547 44744 33581
rect 44800 33547 44834 33581
rect 44890 33547 44924 33581
rect 44980 33547 45014 33581
rect 45070 33547 45104 33581
rect 45160 33547 45194 33581
rect 45250 33547 45284 33581
rect 45340 33547 45374 33581
rect 45430 33547 45464 33581
rect 45520 33547 45554 33581
rect 45610 33547 45644 33581
rect 45711 33524 45745 33558
rect 45864 33524 45898 33558
rect 45960 33547 45994 33581
rect 46050 33547 46084 33581
rect 46140 33547 46174 33581
rect 46230 33547 46264 33581
rect 46320 33547 46354 33581
rect 46410 33547 46444 33581
rect 46500 33547 46534 33581
rect 46590 33547 46624 33581
rect 46680 33547 46714 33581
rect 46770 33547 46804 33581
rect 46860 33547 46894 33581
rect 46950 33547 46984 33581
rect 47051 33524 47085 33558
rect 47204 33524 47238 33558
rect 47300 33547 47334 33581
rect 47390 33547 47424 33581
rect 47480 33547 47514 33581
rect 47570 33547 47604 33581
rect 47660 33547 47694 33581
rect 47750 33547 47784 33581
rect 47840 33547 47874 33581
rect 47930 33547 47964 33581
rect 48020 33547 48054 33581
rect 48110 33547 48144 33581
rect 48200 33547 48234 33581
rect 48290 33547 48324 33581
rect 48391 33524 48425 33558
rect 48544 33524 48578 33558
rect 48640 33547 48674 33581
rect 48730 33547 48764 33581
rect 48820 33547 48854 33581
rect 48910 33547 48944 33581
rect 49000 33547 49034 33581
rect 49090 33547 49124 33581
rect 49180 33547 49214 33581
rect 49270 33547 49304 33581
rect 49360 33547 49394 33581
rect 49450 33547 49484 33581
rect 49540 33547 49574 33581
rect 49630 33547 49664 33581
rect 49731 33524 49765 33558
rect 49884 33524 49918 33558
rect 49980 33547 50014 33581
rect 50070 33547 50104 33581
rect 50160 33547 50194 33581
rect 50250 33547 50284 33581
rect 50340 33547 50374 33581
rect 50430 33547 50464 33581
rect 50520 33547 50554 33581
rect 50610 33547 50644 33581
rect 50700 33547 50734 33581
rect 50790 33547 50824 33581
rect 50880 33547 50914 33581
rect 50970 33547 51004 33581
rect 51071 33524 51105 33558
rect 51224 33524 51258 33558
rect 51320 33547 51354 33581
rect 51410 33547 51444 33581
rect 51500 33547 51534 33581
rect 51590 33547 51624 33581
rect 51680 33547 51714 33581
rect 51770 33547 51804 33581
rect 51860 33547 51894 33581
rect 51950 33547 51984 33581
rect 52040 33547 52074 33581
rect 52130 33547 52164 33581
rect 52220 33547 52254 33581
rect 52310 33547 52344 33581
rect 52411 33524 52445 33558
rect 41844 33434 41878 33468
rect 41844 33344 41878 33378
rect 41844 33254 41878 33288
rect 41844 33164 41878 33198
rect 41844 33074 41878 33108
rect 20263 32861 20705 32963
rect 23295 32861 23737 32963
rect 41844 32984 41878 33018
rect 41844 32894 41878 32928
rect 41844 32804 41878 32838
rect 41844 32714 41878 32748
rect 41844 32624 41878 32658
rect 41844 32534 41878 32568
rect 43031 33434 43065 33468
rect 43184 33434 43218 33468
rect 43031 33344 43065 33378
rect 43184 33344 43218 33378
rect 43031 33254 43065 33288
rect 43184 33254 43218 33288
rect 43031 33164 43065 33198
rect 43184 33164 43218 33198
rect 43031 33074 43065 33108
rect 43184 33074 43218 33108
rect 43031 32984 43065 33018
rect 43184 32984 43218 33018
rect 43031 32894 43065 32928
rect 43184 32894 43218 32928
rect 43031 32804 43065 32838
rect 43184 32804 43218 32838
rect 43031 32714 43065 32748
rect 43184 32714 43218 32748
rect 43031 32624 43065 32658
rect 43184 32624 43218 32658
rect 43031 32534 43065 32568
rect 43184 32534 43218 32568
rect 41844 32444 41878 32478
rect 44371 33434 44405 33468
rect 44524 33434 44558 33468
rect 44371 33344 44405 33378
rect 44524 33344 44558 33378
rect 44371 33254 44405 33288
rect 44524 33254 44558 33288
rect 44371 33164 44405 33198
rect 44524 33164 44558 33198
rect 44371 33074 44405 33108
rect 44524 33074 44558 33108
rect 44371 32984 44405 33018
rect 44524 32984 44558 33018
rect 44371 32894 44405 32928
rect 44524 32894 44558 32928
rect 44371 32804 44405 32838
rect 44524 32804 44558 32838
rect 44371 32714 44405 32748
rect 44524 32714 44558 32748
rect 44371 32624 44405 32658
rect 44524 32624 44558 32658
rect 44371 32534 44405 32568
rect 44524 32534 44558 32568
rect 43031 32444 43065 32478
rect 43184 32444 43218 32478
rect 45711 33434 45745 33468
rect 45864 33434 45898 33468
rect 45711 33344 45745 33378
rect 45864 33344 45898 33378
rect 45711 33254 45745 33288
rect 45864 33254 45898 33288
rect 45711 33164 45745 33198
rect 45864 33164 45898 33198
rect 45711 33074 45745 33108
rect 45864 33074 45898 33108
rect 45711 32984 45745 33018
rect 45864 32984 45898 33018
rect 45711 32894 45745 32928
rect 45864 32894 45898 32928
rect 45711 32804 45745 32838
rect 45864 32804 45898 32838
rect 45711 32714 45745 32748
rect 45864 32714 45898 32748
rect 45711 32624 45745 32658
rect 45864 32624 45898 32658
rect 45711 32534 45745 32568
rect 45864 32534 45898 32568
rect 44371 32444 44405 32478
rect 44524 32444 44558 32478
rect 47051 33434 47085 33468
rect 47204 33434 47238 33468
rect 47051 33344 47085 33378
rect 47204 33344 47238 33378
rect 47051 33254 47085 33288
rect 47204 33254 47238 33288
rect 47051 33164 47085 33198
rect 47204 33164 47238 33198
rect 47051 33074 47085 33108
rect 47204 33074 47238 33108
rect 47051 32984 47085 33018
rect 47204 32984 47238 33018
rect 47051 32894 47085 32928
rect 47204 32894 47238 32928
rect 47051 32804 47085 32838
rect 47204 32804 47238 32838
rect 47051 32714 47085 32748
rect 47204 32714 47238 32748
rect 47051 32624 47085 32658
rect 47204 32624 47238 32658
rect 47051 32534 47085 32568
rect 47204 32534 47238 32568
rect 45711 32444 45745 32478
rect 45864 32444 45898 32478
rect 48391 33434 48425 33468
rect 48544 33434 48578 33468
rect 48391 33344 48425 33378
rect 48544 33344 48578 33378
rect 48391 33254 48425 33288
rect 48544 33254 48578 33288
rect 48391 33164 48425 33198
rect 48544 33164 48578 33198
rect 48391 33074 48425 33108
rect 48544 33074 48578 33108
rect 48391 32984 48425 33018
rect 48544 32984 48578 33018
rect 48391 32894 48425 32928
rect 48544 32894 48578 32928
rect 48391 32804 48425 32838
rect 48544 32804 48578 32838
rect 48391 32714 48425 32748
rect 48544 32714 48578 32748
rect 48391 32624 48425 32658
rect 48544 32624 48578 32658
rect 48391 32534 48425 32568
rect 48544 32534 48578 32568
rect 47051 32444 47085 32478
rect 47204 32444 47238 32478
rect 49731 33434 49765 33468
rect 49884 33434 49918 33468
rect 49731 33344 49765 33378
rect 49884 33344 49918 33378
rect 49731 33254 49765 33288
rect 49884 33254 49918 33288
rect 49731 33164 49765 33198
rect 49884 33164 49918 33198
rect 49731 33074 49765 33108
rect 49884 33074 49918 33108
rect 49731 32984 49765 33018
rect 49884 32984 49918 33018
rect 49731 32894 49765 32928
rect 49884 32894 49918 32928
rect 49731 32804 49765 32838
rect 49884 32804 49918 32838
rect 49731 32714 49765 32748
rect 49884 32714 49918 32748
rect 49731 32624 49765 32658
rect 49884 32624 49918 32658
rect 49731 32534 49765 32568
rect 49884 32534 49918 32568
rect 48391 32444 48425 32478
rect 48544 32444 48578 32478
rect 51071 33434 51105 33468
rect 51224 33434 51258 33468
rect 51071 33344 51105 33378
rect 51224 33344 51258 33378
rect 51071 33254 51105 33288
rect 51224 33254 51258 33288
rect 51071 33164 51105 33198
rect 51224 33164 51258 33198
rect 51071 33074 51105 33108
rect 51224 33074 51258 33108
rect 51071 32984 51105 33018
rect 51224 32984 51258 33018
rect 51071 32894 51105 32928
rect 51224 32894 51258 32928
rect 51071 32804 51105 32838
rect 51224 32804 51258 32838
rect 51071 32714 51105 32748
rect 51224 32714 51258 32748
rect 51071 32624 51105 32658
rect 51224 32624 51258 32658
rect 51071 32534 51105 32568
rect 51224 32534 51258 32568
rect 49731 32444 49765 32478
rect 49884 32444 49918 32478
rect 52411 33434 52445 33468
rect 52411 33344 52445 33378
rect 52411 33254 52445 33288
rect 52411 33164 52445 33198
rect 52411 33074 52445 33108
rect 52411 32984 52445 33018
rect 52411 32894 52445 32928
rect 52411 32804 52445 32838
rect 52411 32714 52445 32748
rect 52411 32624 52445 32658
rect 52411 32534 52445 32568
rect 51071 32444 51105 32478
rect 51224 32444 51258 32478
rect 52411 32444 52445 32478
rect 41940 32360 41974 32394
rect 42030 32360 42064 32394
rect 42120 32360 42154 32394
rect 42210 32360 42244 32394
rect 42300 32360 42334 32394
rect 42390 32360 42424 32394
rect 42480 32360 42514 32394
rect 42570 32360 42604 32394
rect 42660 32360 42694 32394
rect 42750 32360 42784 32394
rect 42840 32360 42874 32394
rect 42930 32360 42964 32394
rect 43280 32360 43314 32394
rect 43370 32360 43404 32394
rect 43460 32360 43494 32394
rect 43550 32360 43584 32394
rect 43640 32360 43674 32394
rect 43730 32360 43764 32394
rect 43820 32360 43854 32394
rect 43910 32360 43944 32394
rect 44000 32360 44034 32394
rect 44090 32360 44124 32394
rect 44180 32360 44214 32394
rect 44270 32360 44304 32394
rect 44620 32360 44654 32394
rect 44710 32360 44744 32394
rect 44800 32360 44834 32394
rect 44890 32360 44924 32394
rect 44980 32360 45014 32394
rect 45070 32360 45104 32394
rect 45160 32360 45194 32394
rect 45250 32360 45284 32394
rect 45340 32360 45374 32394
rect 45430 32360 45464 32394
rect 45520 32360 45554 32394
rect 45610 32360 45644 32394
rect 45960 32360 45994 32394
rect 46050 32360 46084 32394
rect 46140 32360 46174 32394
rect 46230 32360 46264 32394
rect 46320 32360 46354 32394
rect 46410 32360 46444 32394
rect 46500 32360 46534 32394
rect 46590 32360 46624 32394
rect 46680 32360 46714 32394
rect 46770 32360 46804 32394
rect 46860 32360 46894 32394
rect 46950 32360 46984 32394
rect 47300 32360 47334 32394
rect 47390 32360 47424 32394
rect 47480 32360 47514 32394
rect 47570 32360 47604 32394
rect 47660 32360 47694 32394
rect 47750 32360 47784 32394
rect 47840 32360 47874 32394
rect 47930 32360 47964 32394
rect 48020 32360 48054 32394
rect 48110 32360 48144 32394
rect 48200 32360 48234 32394
rect 48290 32360 48324 32394
rect 48640 32360 48674 32394
rect 48730 32360 48764 32394
rect 48820 32360 48854 32394
rect 48910 32360 48944 32394
rect 49000 32360 49034 32394
rect 49090 32360 49124 32394
rect 49180 32360 49214 32394
rect 49270 32360 49304 32394
rect 49360 32360 49394 32394
rect 49450 32360 49484 32394
rect 49540 32360 49574 32394
rect 49630 32360 49664 32394
rect 49980 32360 50014 32394
rect 50070 32360 50104 32394
rect 50160 32360 50194 32394
rect 50250 32360 50284 32394
rect 50340 32360 50374 32394
rect 50430 32360 50464 32394
rect 50520 32360 50554 32394
rect 50610 32360 50644 32394
rect 50700 32360 50734 32394
rect 50790 32360 50824 32394
rect 50880 32360 50914 32394
rect 50970 32360 51004 32394
rect 51320 32360 51354 32394
rect 51410 32360 51444 32394
rect 51500 32360 51534 32394
rect 51590 32360 51624 32394
rect 51680 32360 51714 32394
rect 51770 32360 51804 32394
rect 51860 32360 51894 32394
rect 51950 32360 51984 32394
rect 52040 32360 52074 32394
rect 52130 32360 52164 32394
rect 52220 32360 52254 32394
rect 52310 32360 52344 32394
rect 17519 29101 17961 29203
rect 20263 29101 20705 29203
rect 23007 29101 23449 29203
rect 28201 29101 28643 29203
rect 41844 29764 41878 29798
rect 41940 29787 41974 29821
rect 42030 29787 42064 29821
rect 42120 29787 42154 29821
rect 42210 29787 42244 29821
rect 42300 29787 42334 29821
rect 42390 29787 42424 29821
rect 42480 29787 42514 29821
rect 42570 29787 42604 29821
rect 42660 29787 42694 29821
rect 42750 29787 42784 29821
rect 42840 29787 42874 29821
rect 42930 29787 42964 29821
rect 43031 29764 43065 29798
rect 43184 29764 43218 29798
rect 43280 29787 43314 29821
rect 43370 29787 43404 29821
rect 43460 29787 43494 29821
rect 43550 29787 43584 29821
rect 43640 29787 43674 29821
rect 43730 29787 43764 29821
rect 43820 29787 43854 29821
rect 43910 29787 43944 29821
rect 44000 29787 44034 29821
rect 44090 29787 44124 29821
rect 44180 29787 44214 29821
rect 44270 29787 44304 29821
rect 44371 29764 44405 29798
rect 44524 29764 44558 29798
rect 44620 29787 44654 29821
rect 44710 29787 44744 29821
rect 44800 29787 44834 29821
rect 44890 29787 44924 29821
rect 44980 29787 45014 29821
rect 45070 29787 45104 29821
rect 45160 29787 45194 29821
rect 45250 29787 45284 29821
rect 45340 29787 45374 29821
rect 45430 29787 45464 29821
rect 45520 29787 45554 29821
rect 45610 29787 45644 29821
rect 45711 29764 45745 29798
rect 45864 29764 45898 29798
rect 45960 29787 45994 29821
rect 46050 29787 46084 29821
rect 46140 29787 46174 29821
rect 46230 29787 46264 29821
rect 46320 29787 46354 29821
rect 46410 29787 46444 29821
rect 46500 29787 46534 29821
rect 46590 29787 46624 29821
rect 46680 29787 46714 29821
rect 46770 29787 46804 29821
rect 46860 29787 46894 29821
rect 46950 29787 46984 29821
rect 47051 29764 47085 29798
rect 47204 29764 47238 29798
rect 47300 29787 47334 29821
rect 47390 29787 47424 29821
rect 47480 29787 47514 29821
rect 47570 29787 47604 29821
rect 47660 29787 47694 29821
rect 47750 29787 47784 29821
rect 47840 29787 47874 29821
rect 47930 29787 47964 29821
rect 48020 29787 48054 29821
rect 48110 29787 48144 29821
rect 48200 29787 48234 29821
rect 48290 29787 48324 29821
rect 48391 29764 48425 29798
rect 48544 29764 48578 29798
rect 48640 29787 48674 29821
rect 48730 29787 48764 29821
rect 48820 29787 48854 29821
rect 48910 29787 48944 29821
rect 49000 29787 49034 29821
rect 49090 29787 49124 29821
rect 49180 29787 49214 29821
rect 49270 29787 49304 29821
rect 49360 29787 49394 29821
rect 49450 29787 49484 29821
rect 49540 29787 49574 29821
rect 49630 29787 49664 29821
rect 49731 29764 49765 29798
rect 49884 29764 49918 29798
rect 49980 29787 50014 29821
rect 50070 29787 50104 29821
rect 50160 29787 50194 29821
rect 50250 29787 50284 29821
rect 50340 29787 50374 29821
rect 50430 29787 50464 29821
rect 50520 29787 50554 29821
rect 50610 29787 50644 29821
rect 50700 29787 50734 29821
rect 50790 29787 50824 29821
rect 50880 29787 50914 29821
rect 50970 29787 51004 29821
rect 51071 29764 51105 29798
rect 51224 29764 51258 29798
rect 51320 29787 51354 29821
rect 51410 29787 51444 29821
rect 51500 29787 51534 29821
rect 51590 29787 51624 29821
rect 51680 29787 51714 29821
rect 51770 29787 51804 29821
rect 51860 29787 51894 29821
rect 51950 29787 51984 29821
rect 52040 29787 52074 29821
rect 52130 29787 52164 29821
rect 52220 29787 52254 29821
rect 52310 29787 52344 29821
rect 52411 29764 52445 29798
rect 41844 29674 41878 29708
rect 41844 29584 41878 29618
rect 41844 29494 41878 29528
rect 41844 29404 41878 29438
rect 41844 29314 41878 29348
rect 41844 29224 41878 29258
rect 41844 29134 41878 29168
rect 41844 29044 41878 29078
rect 41844 28954 41878 28988
rect 41844 28864 41878 28898
rect 41844 28774 41878 28808
rect 43031 29674 43065 29708
rect 43184 29674 43218 29708
rect 43031 29584 43065 29618
rect 43184 29584 43218 29618
rect 43031 29494 43065 29528
rect 43184 29494 43218 29528
rect 43031 29404 43065 29438
rect 43184 29404 43218 29438
rect 43031 29314 43065 29348
rect 43184 29314 43218 29348
rect 43031 29224 43065 29258
rect 43184 29224 43218 29258
rect 43031 29134 43065 29168
rect 43184 29134 43218 29168
rect 43031 29044 43065 29078
rect 43184 29044 43218 29078
rect 43031 28954 43065 28988
rect 43184 28954 43218 28988
rect 43031 28864 43065 28898
rect 43184 28864 43218 28898
rect 43031 28774 43065 28808
rect 43184 28774 43218 28808
rect 41844 28684 41878 28718
rect 44371 29674 44405 29708
rect 44524 29674 44558 29708
rect 44371 29584 44405 29618
rect 44524 29584 44558 29618
rect 44371 29494 44405 29528
rect 44524 29494 44558 29528
rect 44371 29404 44405 29438
rect 44524 29404 44558 29438
rect 44371 29314 44405 29348
rect 44524 29314 44558 29348
rect 44371 29224 44405 29258
rect 44524 29224 44558 29258
rect 44371 29134 44405 29168
rect 44524 29134 44558 29168
rect 44371 29044 44405 29078
rect 44524 29044 44558 29078
rect 44371 28954 44405 28988
rect 44524 28954 44558 28988
rect 44371 28864 44405 28898
rect 44524 28864 44558 28898
rect 44371 28774 44405 28808
rect 44524 28774 44558 28808
rect 43031 28684 43065 28718
rect 43184 28684 43218 28718
rect 45711 29674 45745 29708
rect 45864 29674 45898 29708
rect 45711 29584 45745 29618
rect 45864 29584 45898 29618
rect 45711 29494 45745 29528
rect 45864 29494 45898 29528
rect 45711 29404 45745 29438
rect 45864 29404 45898 29438
rect 45711 29314 45745 29348
rect 45864 29314 45898 29348
rect 45711 29224 45745 29258
rect 45864 29224 45898 29258
rect 45711 29134 45745 29168
rect 45864 29134 45898 29168
rect 45711 29044 45745 29078
rect 45864 29044 45898 29078
rect 45711 28954 45745 28988
rect 45864 28954 45898 28988
rect 45711 28864 45745 28898
rect 45864 28864 45898 28898
rect 45711 28774 45745 28808
rect 45864 28774 45898 28808
rect 44371 28684 44405 28718
rect 44524 28684 44558 28718
rect 47051 29674 47085 29708
rect 47204 29674 47238 29708
rect 47051 29584 47085 29618
rect 47204 29584 47238 29618
rect 47051 29494 47085 29528
rect 47204 29494 47238 29528
rect 47051 29404 47085 29438
rect 47204 29404 47238 29438
rect 47051 29314 47085 29348
rect 47204 29314 47238 29348
rect 47051 29224 47085 29258
rect 47204 29224 47238 29258
rect 47051 29134 47085 29168
rect 47204 29134 47238 29168
rect 47051 29044 47085 29078
rect 47204 29044 47238 29078
rect 47051 28954 47085 28988
rect 47204 28954 47238 28988
rect 47051 28864 47085 28898
rect 47204 28864 47238 28898
rect 47051 28774 47085 28808
rect 47204 28774 47238 28808
rect 45711 28684 45745 28718
rect 45864 28684 45898 28718
rect 48391 29674 48425 29708
rect 48544 29674 48578 29708
rect 48391 29584 48425 29618
rect 48544 29584 48578 29618
rect 48391 29494 48425 29528
rect 48544 29494 48578 29528
rect 48391 29404 48425 29438
rect 48544 29404 48578 29438
rect 48391 29314 48425 29348
rect 48544 29314 48578 29348
rect 48391 29224 48425 29258
rect 48544 29224 48578 29258
rect 48391 29134 48425 29168
rect 48544 29134 48578 29168
rect 48391 29044 48425 29078
rect 48544 29044 48578 29078
rect 48391 28954 48425 28988
rect 48544 28954 48578 28988
rect 48391 28864 48425 28898
rect 48544 28864 48578 28898
rect 48391 28774 48425 28808
rect 48544 28774 48578 28808
rect 47051 28684 47085 28718
rect 47204 28684 47238 28718
rect 49731 29674 49765 29708
rect 49884 29674 49918 29708
rect 49731 29584 49765 29618
rect 49884 29584 49918 29618
rect 49731 29494 49765 29528
rect 49884 29494 49918 29528
rect 49731 29404 49765 29438
rect 49884 29404 49918 29438
rect 49731 29314 49765 29348
rect 49884 29314 49918 29348
rect 49731 29224 49765 29258
rect 49884 29224 49918 29258
rect 49731 29134 49765 29168
rect 49884 29134 49918 29168
rect 49731 29044 49765 29078
rect 49884 29044 49918 29078
rect 49731 28954 49765 28988
rect 49884 28954 49918 28988
rect 49731 28864 49765 28898
rect 49884 28864 49918 28898
rect 49731 28774 49765 28808
rect 49884 28774 49918 28808
rect 48391 28684 48425 28718
rect 48544 28684 48578 28718
rect 51071 29674 51105 29708
rect 51224 29674 51258 29708
rect 51071 29584 51105 29618
rect 51224 29584 51258 29618
rect 51071 29494 51105 29528
rect 51224 29494 51258 29528
rect 51071 29404 51105 29438
rect 51224 29404 51258 29438
rect 51071 29314 51105 29348
rect 51224 29314 51258 29348
rect 51071 29224 51105 29258
rect 51224 29224 51258 29258
rect 51071 29134 51105 29168
rect 51224 29134 51258 29168
rect 51071 29044 51105 29078
rect 51224 29044 51258 29078
rect 51071 28954 51105 28988
rect 51224 28954 51258 28988
rect 51071 28864 51105 28898
rect 51224 28864 51258 28898
rect 51071 28774 51105 28808
rect 51224 28774 51258 28808
rect 49731 28684 49765 28718
rect 49884 28684 49918 28718
rect 52411 29674 52445 29708
rect 52411 29584 52445 29618
rect 52411 29494 52445 29528
rect 52411 29404 52445 29438
rect 52411 29314 52445 29348
rect 52411 29224 52445 29258
rect 52411 29134 52445 29168
rect 52411 29044 52445 29078
rect 52411 28954 52445 28988
rect 52411 28864 52445 28898
rect 52411 28774 52445 28808
rect 51071 28684 51105 28718
rect 51224 28684 51258 28718
rect 52411 28684 52445 28718
rect 41940 28600 41974 28634
rect 42030 28600 42064 28634
rect 42120 28600 42154 28634
rect 42210 28600 42244 28634
rect 42300 28600 42334 28634
rect 42390 28600 42424 28634
rect 42480 28600 42514 28634
rect 42570 28600 42604 28634
rect 42660 28600 42694 28634
rect 42750 28600 42784 28634
rect 42840 28600 42874 28634
rect 42930 28600 42964 28634
rect 43280 28600 43314 28634
rect 43370 28600 43404 28634
rect 43460 28600 43494 28634
rect 43550 28600 43584 28634
rect 43640 28600 43674 28634
rect 43730 28600 43764 28634
rect 43820 28600 43854 28634
rect 43910 28600 43944 28634
rect 44000 28600 44034 28634
rect 44090 28600 44124 28634
rect 44180 28600 44214 28634
rect 44270 28600 44304 28634
rect 44620 28600 44654 28634
rect 44710 28600 44744 28634
rect 44800 28600 44834 28634
rect 44890 28600 44924 28634
rect 44980 28600 45014 28634
rect 45070 28600 45104 28634
rect 45160 28600 45194 28634
rect 45250 28600 45284 28634
rect 45340 28600 45374 28634
rect 45430 28600 45464 28634
rect 45520 28600 45554 28634
rect 45610 28600 45644 28634
rect 45960 28600 45994 28634
rect 46050 28600 46084 28634
rect 46140 28600 46174 28634
rect 46230 28600 46264 28634
rect 46320 28600 46354 28634
rect 46410 28600 46444 28634
rect 46500 28600 46534 28634
rect 46590 28600 46624 28634
rect 46680 28600 46714 28634
rect 46770 28600 46804 28634
rect 46860 28600 46894 28634
rect 46950 28600 46984 28634
rect 47300 28600 47334 28634
rect 47390 28600 47424 28634
rect 47480 28600 47514 28634
rect 47570 28600 47604 28634
rect 47660 28600 47694 28634
rect 47750 28600 47784 28634
rect 47840 28600 47874 28634
rect 47930 28600 47964 28634
rect 48020 28600 48054 28634
rect 48110 28600 48144 28634
rect 48200 28600 48234 28634
rect 48290 28600 48324 28634
rect 48640 28600 48674 28634
rect 48730 28600 48764 28634
rect 48820 28600 48854 28634
rect 48910 28600 48944 28634
rect 49000 28600 49034 28634
rect 49090 28600 49124 28634
rect 49180 28600 49214 28634
rect 49270 28600 49304 28634
rect 49360 28600 49394 28634
rect 49450 28600 49484 28634
rect 49540 28600 49574 28634
rect 49630 28600 49664 28634
rect 49980 28600 50014 28634
rect 50070 28600 50104 28634
rect 50160 28600 50194 28634
rect 50250 28600 50284 28634
rect 50340 28600 50374 28634
rect 50430 28600 50464 28634
rect 50520 28600 50554 28634
rect 50610 28600 50644 28634
rect 50700 28600 50734 28634
rect 50790 28600 50824 28634
rect 50880 28600 50914 28634
rect 50970 28600 51004 28634
rect 51320 28600 51354 28634
rect 51410 28600 51444 28634
rect 51500 28600 51534 28634
rect 51590 28600 51624 28634
rect 51680 28600 51714 28634
rect 51770 28600 51804 28634
rect 51860 28600 51894 28634
rect 51950 28600 51984 28634
rect 52040 28600 52074 28634
rect 52130 28600 52164 28634
rect 52220 28600 52254 28634
rect 52310 28600 52344 28634
rect 23399 25341 23841 25443
rect 38393 25341 38835 25443
rect 41137 25341 41579 25443
rect 43881 25341 44323 25443
rect 46625 25341 47067 25443
rect 49369 25341 49811 25443
rect 25361 24635 25395 24669
rect 26463 24605 26497 24639
rect 27763 24605 27797 24639
rect 24869 21581 25311 21683
rect 28201 21581 28643 21683
rect 30945 21581 31387 21683
rect 34179 21581 34621 21683
rect 38393 21581 38835 21683
rect 41137 21581 41579 21683
rect 49369 21581 49811 21683
rect 44861 14061 45303 14163
rect 47605 14061 48047 14163
rect 50349 14061 50791 14163
rect 44763 10301 45205 10403
rect 47507 10301 47949 10403
rect 50251 10301 50693 10403
rect 45547 6541 45989 6643
rect 48291 6541 48733 6643
rect 51035 6541 51477 6643
<< nsubdiffcont >>
rect 25873 48845 25907 48879
rect 27173 48845 27207 48879
rect 28473 48845 28507 48879
rect 29773 48845 29807 48879
rect 31073 48845 31107 48879
rect 32373 48845 32407 48879
rect 33673 48845 33707 48879
rect 34973 48845 35007 48879
rect 36273 48845 36307 48879
rect 37573 48845 37607 48879
rect 38873 48845 38907 48879
rect 40173 48845 40207 48879
rect 41473 48845 41507 48879
rect 42773 48845 42807 48879
rect 44073 48845 44107 48879
rect 45373 48845 45407 48879
rect 46673 48845 46707 48879
rect 47973 48845 48007 48879
rect 49273 48845 49307 48879
rect 50573 48845 50607 48879
rect 24773 48795 24807 48829
rect 16073 45085 16107 45119
rect 17373 45085 17407 45119
rect 18673 45085 18707 45119
rect 19973 45085 20007 45119
rect 21273 45085 21307 45119
rect 22573 45085 22607 45119
rect 23873 45085 23907 45119
rect 25173 45085 25207 45119
rect 26473 45085 26507 45119
rect 27773 45085 27807 45119
rect 29073 45085 29107 45119
rect 30373 45085 30407 45119
rect 31673 45085 31707 45119
rect 32973 45085 33007 45119
rect 34273 45085 34307 45119
rect 35573 45085 35607 45119
rect 36873 45085 36907 45119
rect 38173 45085 38207 45119
rect 39473 45085 39507 45119
rect 40773 45085 40807 45119
rect 14973 45035 15007 45069
rect 43280 44680 43314 44714
rect 43370 44680 43404 44714
rect 43460 44680 43494 44714
rect 43550 44680 43584 44714
rect 43640 44680 43674 44714
rect 43730 44680 43764 44714
rect 43820 44680 43854 44714
rect 43910 44680 43944 44714
rect 44000 44680 44034 44714
rect 43168 44623 43202 44657
rect 44058 44604 44092 44638
rect 43168 44533 43202 44567
rect 43168 44443 43202 44477
rect 43168 44353 43202 44387
rect 43168 44263 43202 44297
rect 43168 44173 43202 44207
rect 43168 44083 43202 44117
rect 43168 43993 43202 44027
rect 43168 43903 43202 43937
rect 44058 44514 44092 44548
rect 44058 44424 44092 44458
rect 44058 44334 44092 44368
rect 44058 44244 44092 44278
rect 44058 44154 44092 44188
rect 44058 44064 44092 44098
rect 44058 43974 44092 44008
rect 44058 43884 44092 43918
rect 43246 43790 43280 43824
rect 43336 43790 43370 43824
rect 43426 43790 43460 43824
rect 43516 43790 43550 43824
rect 43606 43790 43640 43824
rect 43696 43790 43730 43824
rect 43786 43790 43820 43824
rect 43876 43790 43910 43824
rect 43966 43790 44000 43824
rect 44620 44680 44654 44714
rect 44710 44680 44744 44714
rect 44800 44680 44834 44714
rect 44890 44680 44924 44714
rect 44980 44680 45014 44714
rect 45070 44680 45104 44714
rect 45160 44680 45194 44714
rect 45250 44680 45284 44714
rect 45340 44680 45374 44714
rect 44508 44623 44542 44657
rect 45398 44604 45432 44638
rect 44508 44533 44542 44567
rect 44508 44443 44542 44477
rect 44508 44353 44542 44387
rect 44508 44263 44542 44297
rect 44508 44173 44542 44207
rect 44508 44083 44542 44117
rect 44508 43993 44542 44027
rect 44508 43903 44542 43937
rect 45398 44514 45432 44548
rect 45398 44424 45432 44458
rect 45398 44334 45432 44368
rect 45398 44244 45432 44278
rect 45398 44154 45432 44188
rect 45398 44064 45432 44098
rect 45398 43974 45432 44008
rect 45398 43884 45432 43918
rect 44586 43790 44620 43824
rect 44676 43790 44710 43824
rect 44766 43790 44800 43824
rect 44856 43790 44890 43824
rect 44946 43790 44980 43824
rect 45036 43790 45070 43824
rect 45126 43790 45160 43824
rect 45216 43790 45250 43824
rect 45306 43790 45340 43824
rect 45960 44680 45994 44714
rect 46050 44680 46084 44714
rect 46140 44680 46174 44714
rect 46230 44680 46264 44714
rect 46320 44680 46354 44714
rect 46410 44680 46444 44714
rect 46500 44680 46534 44714
rect 46590 44680 46624 44714
rect 46680 44680 46714 44714
rect 45848 44623 45882 44657
rect 46738 44604 46772 44638
rect 45848 44533 45882 44567
rect 45848 44443 45882 44477
rect 45848 44353 45882 44387
rect 45848 44263 45882 44297
rect 45848 44173 45882 44207
rect 45848 44083 45882 44117
rect 45848 43993 45882 44027
rect 45848 43903 45882 43937
rect 46738 44514 46772 44548
rect 46738 44424 46772 44458
rect 46738 44334 46772 44368
rect 46738 44244 46772 44278
rect 46738 44154 46772 44188
rect 46738 44064 46772 44098
rect 46738 43974 46772 44008
rect 46738 43884 46772 43918
rect 45926 43790 45960 43824
rect 46016 43790 46050 43824
rect 46106 43790 46140 43824
rect 46196 43790 46230 43824
rect 46286 43790 46320 43824
rect 46376 43790 46410 43824
rect 46466 43790 46500 43824
rect 46556 43790 46590 43824
rect 46646 43790 46680 43824
rect 47300 44680 47334 44714
rect 47390 44680 47424 44714
rect 47480 44680 47514 44714
rect 47570 44680 47604 44714
rect 47660 44680 47694 44714
rect 47750 44680 47784 44714
rect 47840 44680 47874 44714
rect 47930 44680 47964 44714
rect 48020 44680 48054 44714
rect 47188 44623 47222 44657
rect 48078 44604 48112 44638
rect 47188 44533 47222 44567
rect 47188 44443 47222 44477
rect 47188 44353 47222 44387
rect 47188 44263 47222 44297
rect 47188 44173 47222 44207
rect 47188 44083 47222 44117
rect 47188 43993 47222 44027
rect 47188 43903 47222 43937
rect 48078 44514 48112 44548
rect 48078 44424 48112 44458
rect 48078 44334 48112 44368
rect 48078 44244 48112 44278
rect 48078 44154 48112 44188
rect 48078 44064 48112 44098
rect 48078 43974 48112 44008
rect 48078 43884 48112 43918
rect 47266 43790 47300 43824
rect 47356 43790 47390 43824
rect 47446 43790 47480 43824
rect 47536 43790 47570 43824
rect 47626 43790 47660 43824
rect 47716 43790 47750 43824
rect 47806 43790 47840 43824
rect 47896 43790 47930 43824
rect 47986 43790 48020 43824
rect 48640 44680 48674 44714
rect 48730 44680 48764 44714
rect 48820 44680 48854 44714
rect 48910 44680 48944 44714
rect 49000 44680 49034 44714
rect 49090 44680 49124 44714
rect 49180 44680 49214 44714
rect 49270 44680 49304 44714
rect 49360 44680 49394 44714
rect 48528 44623 48562 44657
rect 49418 44604 49452 44638
rect 48528 44533 48562 44567
rect 48528 44443 48562 44477
rect 48528 44353 48562 44387
rect 48528 44263 48562 44297
rect 48528 44173 48562 44207
rect 48528 44083 48562 44117
rect 48528 43993 48562 44027
rect 48528 43903 48562 43937
rect 49418 44514 49452 44548
rect 49418 44424 49452 44458
rect 49418 44334 49452 44368
rect 49418 44244 49452 44278
rect 49418 44154 49452 44188
rect 49418 44064 49452 44098
rect 49418 43974 49452 44008
rect 49418 43884 49452 43918
rect 48606 43790 48640 43824
rect 48696 43790 48730 43824
rect 48786 43790 48820 43824
rect 48876 43790 48910 43824
rect 48966 43790 49000 43824
rect 49056 43790 49090 43824
rect 49146 43790 49180 43824
rect 49236 43790 49270 43824
rect 49326 43790 49360 43824
rect 49980 44680 50014 44714
rect 50070 44680 50104 44714
rect 50160 44680 50194 44714
rect 50250 44680 50284 44714
rect 50340 44680 50374 44714
rect 50430 44680 50464 44714
rect 50520 44680 50554 44714
rect 50610 44680 50644 44714
rect 50700 44680 50734 44714
rect 49868 44623 49902 44657
rect 50758 44604 50792 44638
rect 49868 44533 49902 44567
rect 49868 44443 49902 44477
rect 49868 44353 49902 44387
rect 49868 44263 49902 44297
rect 49868 44173 49902 44207
rect 49868 44083 49902 44117
rect 49868 43993 49902 44027
rect 49868 43903 49902 43937
rect 50758 44514 50792 44548
rect 50758 44424 50792 44458
rect 50758 44334 50792 44368
rect 50758 44244 50792 44278
rect 50758 44154 50792 44188
rect 50758 44064 50792 44098
rect 50758 43974 50792 44008
rect 50758 43884 50792 43918
rect 49946 43790 49980 43824
rect 50036 43790 50070 43824
rect 50126 43790 50160 43824
rect 50216 43790 50250 43824
rect 50306 43790 50340 43824
rect 50396 43790 50430 43824
rect 50486 43790 50520 43824
rect 50576 43790 50610 43824
rect 50666 43790 50700 43824
rect 51320 44680 51354 44714
rect 51410 44680 51444 44714
rect 51500 44680 51534 44714
rect 51590 44680 51624 44714
rect 51680 44680 51714 44714
rect 51770 44680 51804 44714
rect 51860 44680 51894 44714
rect 51950 44680 51984 44714
rect 52040 44680 52074 44714
rect 51208 44623 51242 44657
rect 52098 44604 52132 44638
rect 51208 44533 51242 44567
rect 51208 44443 51242 44477
rect 51208 44353 51242 44387
rect 51208 44263 51242 44297
rect 51208 44173 51242 44207
rect 51208 44083 51242 44117
rect 51208 43993 51242 44027
rect 51208 43903 51242 43937
rect 52098 44514 52132 44548
rect 52098 44424 52132 44458
rect 52098 44334 52132 44368
rect 52098 44244 52132 44278
rect 52098 44154 52132 44188
rect 52098 44064 52132 44098
rect 52098 43974 52132 44008
rect 52098 43884 52132 43918
rect 51286 43790 51320 43824
rect 51376 43790 51410 43824
rect 51466 43790 51500 43824
rect 51556 43790 51590 43824
rect 51646 43790 51680 43824
rect 51736 43790 51770 43824
rect 51826 43790 51860 43824
rect 51916 43790 51950 43824
rect 52006 43790 52040 43824
rect 23717 41325 23751 41359
rect 25017 41325 25051 41359
rect 26317 41325 26351 41359
rect 22617 41275 22651 41309
rect 30381 41325 30415 41359
rect 31681 41325 31715 41359
rect 32981 41325 33015 41359
rect 29281 41275 29315 41309
rect 42104 40920 42138 40954
rect 42194 40920 42228 40954
rect 42284 40920 42318 40954
rect 42374 40920 42408 40954
rect 42464 40920 42498 40954
rect 42554 40920 42588 40954
rect 42644 40920 42678 40954
rect 42734 40920 42768 40954
rect 42824 40920 42858 40954
rect 41992 40863 42026 40897
rect 42882 40844 42916 40878
rect 41992 40773 42026 40807
rect 41992 40683 42026 40717
rect 41992 40593 42026 40627
rect 41992 40503 42026 40537
rect 41992 40413 42026 40447
rect 41992 40323 42026 40357
rect 41992 40233 42026 40267
rect 41992 40143 42026 40177
rect 42882 40754 42916 40788
rect 42882 40664 42916 40698
rect 42882 40574 42916 40608
rect 42882 40484 42916 40518
rect 42882 40394 42916 40428
rect 42882 40304 42916 40338
rect 42882 40214 42916 40248
rect 42882 40124 42916 40158
rect 42070 40030 42104 40064
rect 42160 40030 42194 40064
rect 42250 40030 42284 40064
rect 42340 40030 42374 40064
rect 42430 40030 42464 40064
rect 42520 40030 42554 40064
rect 42610 40030 42644 40064
rect 42700 40030 42734 40064
rect 42790 40030 42824 40064
rect 43444 40920 43478 40954
rect 43534 40920 43568 40954
rect 43624 40920 43658 40954
rect 43714 40920 43748 40954
rect 43804 40920 43838 40954
rect 43894 40920 43928 40954
rect 43984 40920 44018 40954
rect 44074 40920 44108 40954
rect 44164 40920 44198 40954
rect 43332 40863 43366 40897
rect 44222 40844 44256 40878
rect 43332 40773 43366 40807
rect 43332 40683 43366 40717
rect 43332 40593 43366 40627
rect 43332 40503 43366 40537
rect 43332 40413 43366 40447
rect 43332 40323 43366 40357
rect 43332 40233 43366 40267
rect 43332 40143 43366 40177
rect 44222 40754 44256 40788
rect 44222 40664 44256 40698
rect 44222 40574 44256 40608
rect 44222 40484 44256 40518
rect 44222 40394 44256 40428
rect 44222 40304 44256 40338
rect 44222 40214 44256 40248
rect 44222 40124 44256 40158
rect 43410 40030 43444 40064
rect 43500 40030 43534 40064
rect 43590 40030 43624 40064
rect 43680 40030 43714 40064
rect 43770 40030 43804 40064
rect 43860 40030 43894 40064
rect 43950 40030 43984 40064
rect 44040 40030 44074 40064
rect 44130 40030 44164 40064
rect 44784 40920 44818 40954
rect 44874 40920 44908 40954
rect 44964 40920 44998 40954
rect 45054 40920 45088 40954
rect 45144 40920 45178 40954
rect 45234 40920 45268 40954
rect 45324 40920 45358 40954
rect 45414 40920 45448 40954
rect 45504 40920 45538 40954
rect 44672 40863 44706 40897
rect 45562 40844 45596 40878
rect 44672 40773 44706 40807
rect 44672 40683 44706 40717
rect 44672 40593 44706 40627
rect 44672 40503 44706 40537
rect 44672 40413 44706 40447
rect 44672 40323 44706 40357
rect 44672 40233 44706 40267
rect 44672 40143 44706 40177
rect 45562 40754 45596 40788
rect 45562 40664 45596 40698
rect 45562 40574 45596 40608
rect 45562 40484 45596 40518
rect 45562 40394 45596 40428
rect 45562 40304 45596 40338
rect 45562 40214 45596 40248
rect 45562 40124 45596 40158
rect 44750 40030 44784 40064
rect 44840 40030 44874 40064
rect 44930 40030 44964 40064
rect 45020 40030 45054 40064
rect 45110 40030 45144 40064
rect 45200 40030 45234 40064
rect 45290 40030 45324 40064
rect 45380 40030 45414 40064
rect 45470 40030 45504 40064
rect 46124 40920 46158 40954
rect 46214 40920 46248 40954
rect 46304 40920 46338 40954
rect 46394 40920 46428 40954
rect 46484 40920 46518 40954
rect 46574 40920 46608 40954
rect 46664 40920 46698 40954
rect 46754 40920 46788 40954
rect 46844 40920 46878 40954
rect 46012 40863 46046 40897
rect 46902 40844 46936 40878
rect 46012 40773 46046 40807
rect 46012 40683 46046 40717
rect 46012 40593 46046 40627
rect 46012 40503 46046 40537
rect 46012 40413 46046 40447
rect 46012 40323 46046 40357
rect 46012 40233 46046 40267
rect 46012 40143 46046 40177
rect 46902 40754 46936 40788
rect 46902 40664 46936 40698
rect 46902 40574 46936 40608
rect 46902 40484 46936 40518
rect 46902 40394 46936 40428
rect 46902 40304 46936 40338
rect 46902 40214 46936 40248
rect 46902 40124 46936 40158
rect 46090 40030 46124 40064
rect 46180 40030 46214 40064
rect 46270 40030 46304 40064
rect 46360 40030 46394 40064
rect 46450 40030 46484 40064
rect 46540 40030 46574 40064
rect 46630 40030 46664 40064
rect 46720 40030 46754 40064
rect 46810 40030 46844 40064
rect 47464 40920 47498 40954
rect 47554 40920 47588 40954
rect 47644 40920 47678 40954
rect 47734 40920 47768 40954
rect 47824 40920 47858 40954
rect 47914 40920 47948 40954
rect 48004 40920 48038 40954
rect 48094 40920 48128 40954
rect 48184 40920 48218 40954
rect 47352 40863 47386 40897
rect 48242 40844 48276 40878
rect 47352 40773 47386 40807
rect 47352 40683 47386 40717
rect 47352 40593 47386 40627
rect 47352 40503 47386 40537
rect 47352 40413 47386 40447
rect 47352 40323 47386 40357
rect 47352 40233 47386 40267
rect 47352 40143 47386 40177
rect 48242 40754 48276 40788
rect 48242 40664 48276 40698
rect 48242 40574 48276 40608
rect 48242 40484 48276 40518
rect 48242 40394 48276 40428
rect 48242 40304 48276 40338
rect 48242 40214 48276 40248
rect 48242 40124 48276 40158
rect 47430 40030 47464 40064
rect 47520 40030 47554 40064
rect 47610 40030 47644 40064
rect 47700 40030 47734 40064
rect 47790 40030 47824 40064
rect 47880 40030 47914 40064
rect 47970 40030 48004 40064
rect 48060 40030 48094 40064
rect 48150 40030 48184 40064
rect 48804 40920 48838 40954
rect 48894 40920 48928 40954
rect 48984 40920 49018 40954
rect 49074 40920 49108 40954
rect 49164 40920 49198 40954
rect 49254 40920 49288 40954
rect 49344 40920 49378 40954
rect 49434 40920 49468 40954
rect 49524 40920 49558 40954
rect 48692 40863 48726 40897
rect 49582 40844 49616 40878
rect 48692 40773 48726 40807
rect 48692 40683 48726 40717
rect 48692 40593 48726 40627
rect 48692 40503 48726 40537
rect 48692 40413 48726 40447
rect 48692 40323 48726 40357
rect 48692 40233 48726 40267
rect 48692 40143 48726 40177
rect 49582 40754 49616 40788
rect 49582 40664 49616 40698
rect 49582 40574 49616 40608
rect 49582 40484 49616 40518
rect 49582 40394 49616 40428
rect 49582 40304 49616 40338
rect 49582 40214 49616 40248
rect 49582 40124 49616 40158
rect 48770 40030 48804 40064
rect 48860 40030 48894 40064
rect 48950 40030 48984 40064
rect 49040 40030 49074 40064
rect 49130 40030 49164 40064
rect 49220 40030 49254 40064
rect 49310 40030 49344 40064
rect 49400 40030 49434 40064
rect 49490 40030 49524 40064
rect 50144 40920 50178 40954
rect 50234 40920 50268 40954
rect 50324 40920 50358 40954
rect 50414 40920 50448 40954
rect 50504 40920 50538 40954
rect 50594 40920 50628 40954
rect 50684 40920 50718 40954
rect 50774 40920 50808 40954
rect 50864 40920 50898 40954
rect 50032 40863 50066 40897
rect 50922 40844 50956 40878
rect 50032 40773 50066 40807
rect 50032 40683 50066 40717
rect 50032 40593 50066 40627
rect 50032 40503 50066 40537
rect 50032 40413 50066 40447
rect 50032 40323 50066 40357
rect 50032 40233 50066 40267
rect 50032 40143 50066 40177
rect 50922 40754 50956 40788
rect 50922 40664 50956 40698
rect 50922 40574 50956 40608
rect 50922 40484 50956 40518
rect 50922 40394 50956 40428
rect 50922 40304 50956 40338
rect 50922 40214 50956 40248
rect 50922 40124 50956 40158
rect 50110 40030 50144 40064
rect 50200 40030 50234 40064
rect 50290 40030 50324 40064
rect 50380 40030 50414 40064
rect 50470 40030 50504 40064
rect 50560 40030 50594 40064
rect 50650 40030 50684 40064
rect 50740 40030 50774 40064
rect 50830 40030 50864 40064
rect 51484 40920 51518 40954
rect 51574 40920 51608 40954
rect 51664 40920 51698 40954
rect 51754 40920 51788 40954
rect 51844 40920 51878 40954
rect 51934 40920 51968 40954
rect 52024 40920 52058 40954
rect 52114 40920 52148 40954
rect 52204 40920 52238 40954
rect 51372 40863 51406 40897
rect 52262 40844 52296 40878
rect 51372 40773 51406 40807
rect 51372 40683 51406 40717
rect 51372 40593 51406 40627
rect 51372 40503 51406 40537
rect 51372 40413 51406 40447
rect 51372 40323 51406 40357
rect 51372 40233 51406 40267
rect 51372 40143 51406 40177
rect 52262 40754 52296 40788
rect 52262 40664 52296 40698
rect 52262 40574 52296 40608
rect 52262 40484 52296 40518
rect 52262 40394 52296 40428
rect 52262 40304 52296 40338
rect 52262 40214 52296 40248
rect 52262 40124 52296 40158
rect 51450 40030 51484 40064
rect 51540 40030 51574 40064
rect 51630 40030 51664 40064
rect 51720 40030 51754 40064
rect 51810 40030 51844 40064
rect 51900 40030 51934 40064
rect 51990 40030 52024 40064
rect 52080 40030 52114 40064
rect 52170 40030 52204 40064
rect 38515 37565 38549 37599
rect 37415 37515 37449 37549
rect 12312 37160 12346 37194
rect 12402 37160 12436 37194
rect 12492 37160 12526 37194
rect 12582 37160 12616 37194
rect 12672 37160 12706 37194
rect 12762 37160 12796 37194
rect 12852 37160 12886 37194
rect 12942 37160 12976 37194
rect 13032 37160 13066 37194
rect 12200 37103 12234 37137
rect 13090 37084 13124 37118
rect 12200 37013 12234 37047
rect 12200 36923 12234 36957
rect 12200 36833 12234 36867
rect 12200 36743 12234 36777
rect 12200 36653 12234 36687
rect 12200 36563 12234 36597
rect 12200 36473 12234 36507
rect 12200 36383 12234 36417
rect 13090 36994 13124 37028
rect 13090 36904 13124 36938
rect 13090 36814 13124 36848
rect 13090 36724 13124 36758
rect 13090 36634 13124 36668
rect 13090 36544 13124 36578
rect 13090 36454 13124 36488
rect 13090 36364 13124 36398
rect 12278 36270 12312 36304
rect 12368 36270 12402 36304
rect 12458 36270 12492 36304
rect 12548 36270 12582 36304
rect 12638 36270 12672 36304
rect 12728 36270 12762 36304
rect 12818 36270 12852 36304
rect 12908 36270 12942 36304
rect 12998 36270 13032 36304
rect 42104 37160 42138 37194
rect 42194 37160 42228 37194
rect 42284 37160 42318 37194
rect 42374 37160 42408 37194
rect 42464 37160 42498 37194
rect 42554 37160 42588 37194
rect 42644 37160 42678 37194
rect 42734 37160 42768 37194
rect 42824 37160 42858 37194
rect 41992 37103 42026 37137
rect 42882 37084 42916 37118
rect 41992 37013 42026 37047
rect 41992 36923 42026 36957
rect 41992 36833 42026 36867
rect 41992 36743 42026 36777
rect 41992 36653 42026 36687
rect 41992 36563 42026 36597
rect 41992 36473 42026 36507
rect 41992 36383 42026 36417
rect 42882 36994 42916 37028
rect 42882 36904 42916 36938
rect 42882 36814 42916 36848
rect 42882 36724 42916 36758
rect 42882 36634 42916 36668
rect 42882 36544 42916 36578
rect 42882 36454 42916 36488
rect 42882 36364 42916 36398
rect 42070 36270 42104 36304
rect 42160 36270 42194 36304
rect 42250 36270 42284 36304
rect 42340 36270 42374 36304
rect 42430 36270 42464 36304
rect 42520 36270 42554 36304
rect 42610 36270 42644 36304
rect 42700 36270 42734 36304
rect 42790 36270 42824 36304
rect 43444 37160 43478 37194
rect 43534 37160 43568 37194
rect 43624 37160 43658 37194
rect 43714 37160 43748 37194
rect 43804 37160 43838 37194
rect 43894 37160 43928 37194
rect 43984 37160 44018 37194
rect 44074 37160 44108 37194
rect 44164 37160 44198 37194
rect 43332 37103 43366 37137
rect 44222 37084 44256 37118
rect 43332 37013 43366 37047
rect 43332 36923 43366 36957
rect 43332 36833 43366 36867
rect 43332 36743 43366 36777
rect 43332 36653 43366 36687
rect 43332 36563 43366 36597
rect 43332 36473 43366 36507
rect 43332 36383 43366 36417
rect 44222 36994 44256 37028
rect 44222 36904 44256 36938
rect 44222 36814 44256 36848
rect 44222 36724 44256 36758
rect 44222 36634 44256 36668
rect 44222 36544 44256 36578
rect 44222 36454 44256 36488
rect 44222 36364 44256 36398
rect 43410 36270 43444 36304
rect 43500 36270 43534 36304
rect 43590 36270 43624 36304
rect 43680 36270 43714 36304
rect 43770 36270 43804 36304
rect 43860 36270 43894 36304
rect 43950 36270 43984 36304
rect 44040 36270 44074 36304
rect 44130 36270 44164 36304
rect 44784 37160 44818 37194
rect 44874 37160 44908 37194
rect 44964 37160 44998 37194
rect 45054 37160 45088 37194
rect 45144 37160 45178 37194
rect 45234 37160 45268 37194
rect 45324 37160 45358 37194
rect 45414 37160 45448 37194
rect 45504 37160 45538 37194
rect 44672 37103 44706 37137
rect 45562 37084 45596 37118
rect 44672 37013 44706 37047
rect 44672 36923 44706 36957
rect 44672 36833 44706 36867
rect 44672 36743 44706 36777
rect 44672 36653 44706 36687
rect 44672 36563 44706 36597
rect 44672 36473 44706 36507
rect 44672 36383 44706 36417
rect 45562 36994 45596 37028
rect 45562 36904 45596 36938
rect 45562 36814 45596 36848
rect 45562 36724 45596 36758
rect 45562 36634 45596 36668
rect 45562 36544 45596 36578
rect 45562 36454 45596 36488
rect 45562 36364 45596 36398
rect 44750 36270 44784 36304
rect 44840 36270 44874 36304
rect 44930 36270 44964 36304
rect 45020 36270 45054 36304
rect 45110 36270 45144 36304
rect 45200 36270 45234 36304
rect 45290 36270 45324 36304
rect 45380 36270 45414 36304
rect 45470 36270 45504 36304
rect 46124 37160 46158 37194
rect 46214 37160 46248 37194
rect 46304 37160 46338 37194
rect 46394 37160 46428 37194
rect 46484 37160 46518 37194
rect 46574 37160 46608 37194
rect 46664 37160 46698 37194
rect 46754 37160 46788 37194
rect 46844 37160 46878 37194
rect 46012 37103 46046 37137
rect 46902 37084 46936 37118
rect 46012 37013 46046 37047
rect 46012 36923 46046 36957
rect 46012 36833 46046 36867
rect 46012 36743 46046 36777
rect 46012 36653 46046 36687
rect 46012 36563 46046 36597
rect 46012 36473 46046 36507
rect 46012 36383 46046 36417
rect 46902 36994 46936 37028
rect 46902 36904 46936 36938
rect 46902 36814 46936 36848
rect 46902 36724 46936 36758
rect 46902 36634 46936 36668
rect 46902 36544 46936 36578
rect 46902 36454 46936 36488
rect 46902 36364 46936 36398
rect 46090 36270 46124 36304
rect 46180 36270 46214 36304
rect 46270 36270 46304 36304
rect 46360 36270 46394 36304
rect 46450 36270 46484 36304
rect 46540 36270 46574 36304
rect 46630 36270 46664 36304
rect 46720 36270 46754 36304
rect 46810 36270 46844 36304
rect 47464 37160 47498 37194
rect 47554 37160 47588 37194
rect 47644 37160 47678 37194
rect 47734 37160 47768 37194
rect 47824 37160 47858 37194
rect 47914 37160 47948 37194
rect 48004 37160 48038 37194
rect 48094 37160 48128 37194
rect 48184 37160 48218 37194
rect 47352 37103 47386 37137
rect 48242 37084 48276 37118
rect 47352 37013 47386 37047
rect 47352 36923 47386 36957
rect 47352 36833 47386 36867
rect 47352 36743 47386 36777
rect 47352 36653 47386 36687
rect 47352 36563 47386 36597
rect 47352 36473 47386 36507
rect 47352 36383 47386 36417
rect 48242 36994 48276 37028
rect 48242 36904 48276 36938
rect 48242 36814 48276 36848
rect 48242 36724 48276 36758
rect 48242 36634 48276 36668
rect 48242 36544 48276 36578
rect 48242 36454 48276 36488
rect 48242 36364 48276 36398
rect 47430 36270 47464 36304
rect 47520 36270 47554 36304
rect 47610 36270 47644 36304
rect 47700 36270 47734 36304
rect 47790 36270 47824 36304
rect 47880 36270 47914 36304
rect 47970 36270 48004 36304
rect 48060 36270 48094 36304
rect 48150 36270 48184 36304
rect 48804 37160 48838 37194
rect 48894 37160 48928 37194
rect 48984 37160 49018 37194
rect 49074 37160 49108 37194
rect 49164 37160 49198 37194
rect 49254 37160 49288 37194
rect 49344 37160 49378 37194
rect 49434 37160 49468 37194
rect 49524 37160 49558 37194
rect 48692 37103 48726 37137
rect 49582 37084 49616 37118
rect 48692 37013 48726 37047
rect 48692 36923 48726 36957
rect 48692 36833 48726 36867
rect 48692 36743 48726 36777
rect 48692 36653 48726 36687
rect 48692 36563 48726 36597
rect 48692 36473 48726 36507
rect 48692 36383 48726 36417
rect 49582 36994 49616 37028
rect 49582 36904 49616 36938
rect 49582 36814 49616 36848
rect 49582 36724 49616 36758
rect 49582 36634 49616 36668
rect 49582 36544 49616 36578
rect 49582 36454 49616 36488
rect 49582 36364 49616 36398
rect 48770 36270 48804 36304
rect 48860 36270 48894 36304
rect 48950 36270 48984 36304
rect 49040 36270 49074 36304
rect 49130 36270 49164 36304
rect 49220 36270 49254 36304
rect 49310 36270 49344 36304
rect 49400 36270 49434 36304
rect 49490 36270 49524 36304
rect 50144 37160 50178 37194
rect 50234 37160 50268 37194
rect 50324 37160 50358 37194
rect 50414 37160 50448 37194
rect 50504 37160 50538 37194
rect 50594 37160 50628 37194
rect 50684 37160 50718 37194
rect 50774 37160 50808 37194
rect 50864 37160 50898 37194
rect 50032 37103 50066 37137
rect 50922 37084 50956 37118
rect 50032 37013 50066 37047
rect 50032 36923 50066 36957
rect 50032 36833 50066 36867
rect 50032 36743 50066 36777
rect 50032 36653 50066 36687
rect 50032 36563 50066 36597
rect 50032 36473 50066 36507
rect 50032 36383 50066 36417
rect 50922 36994 50956 37028
rect 50922 36904 50956 36938
rect 50922 36814 50956 36848
rect 50922 36724 50956 36758
rect 50922 36634 50956 36668
rect 50922 36544 50956 36578
rect 50922 36454 50956 36488
rect 50922 36364 50956 36398
rect 50110 36270 50144 36304
rect 50200 36270 50234 36304
rect 50290 36270 50324 36304
rect 50380 36270 50414 36304
rect 50470 36270 50504 36304
rect 50560 36270 50594 36304
rect 50650 36270 50684 36304
rect 50740 36270 50774 36304
rect 50830 36270 50864 36304
rect 51484 37160 51518 37194
rect 51574 37160 51608 37194
rect 51664 37160 51698 37194
rect 51754 37160 51788 37194
rect 51844 37160 51878 37194
rect 51934 37160 51968 37194
rect 52024 37160 52058 37194
rect 52114 37160 52148 37194
rect 52204 37160 52238 37194
rect 51372 37103 51406 37137
rect 52262 37084 52296 37118
rect 51372 37013 51406 37047
rect 51372 36923 51406 36957
rect 51372 36833 51406 36867
rect 51372 36743 51406 36777
rect 51372 36653 51406 36687
rect 51372 36563 51406 36597
rect 51372 36473 51406 36507
rect 51372 36383 51406 36417
rect 52262 36994 52296 37028
rect 52262 36904 52296 36938
rect 52262 36814 52296 36848
rect 52262 36724 52296 36758
rect 52262 36634 52296 36668
rect 52262 36544 52296 36578
rect 52262 36454 52296 36488
rect 52262 36364 52296 36398
rect 51450 36270 51484 36304
rect 51540 36270 51574 36304
rect 51630 36270 51664 36304
rect 51720 36270 51754 36304
rect 51810 36270 51844 36304
rect 51900 36270 51934 36304
rect 51990 36270 52024 36304
rect 52080 36270 52114 36304
rect 52170 36270 52204 36304
rect 42104 33400 42138 33434
rect 42194 33400 42228 33434
rect 42284 33400 42318 33434
rect 42374 33400 42408 33434
rect 42464 33400 42498 33434
rect 42554 33400 42588 33434
rect 42644 33400 42678 33434
rect 42734 33400 42768 33434
rect 42824 33400 42858 33434
rect 41992 33343 42026 33377
rect 42882 33324 42916 33358
rect 41992 33253 42026 33287
rect 41992 33163 42026 33197
rect 41992 33073 42026 33107
rect 41992 32983 42026 33017
rect 41992 32893 42026 32927
rect 41992 32803 42026 32837
rect 41992 32713 42026 32747
rect 41992 32623 42026 32657
rect 42882 33234 42916 33268
rect 42882 33144 42916 33178
rect 42882 33054 42916 33088
rect 42882 32964 42916 32998
rect 42882 32874 42916 32908
rect 42882 32784 42916 32818
rect 42882 32694 42916 32728
rect 42882 32604 42916 32638
rect 42070 32510 42104 32544
rect 42160 32510 42194 32544
rect 42250 32510 42284 32544
rect 42340 32510 42374 32544
rect 42430 32510 42464 32544
rect 42520 32510 42554 32544
rect 42610 32510 42644 32544
rect 42700 32510 42734 32544
rect 42790 32510 42824 32544
rect 43444 33400 43478 33434
rect 43534 33400 43568 33434
rect 43624 33400 43658 33434
rect 43714 33400 43748 33434
rect 43804 33400 43838 33434
rect 43894 33400 43928 33434
rect 43984 33400 44018 33434
rect 44074 33400 44108 33434
rect 44164 33400 44198 33434
rect 43332 33343 43366 33377
rect 44222 33324 44256 33358
rect 43332 33253 43366 33287
rect 43332 33163 43366 33197
rect 43332 33073 43366 33107
rect 43332 32983 43366 33017
rect 43332 32893 43366 32927
rect 43332 32803 43366 32837
rect 43332 32713 43366 32747
rect 43332 32623 43366 32657
rect 44222 33234 44256 33268
rect 44222 33144 44256 33178
rect 44222 33054 44256 33088
rect 44222 32964 44256 32998
rect 44222 32874 44256 32908
rect 44222 32784 44256 32818
rect 44222 32694 44256 32728
rect 44222 32604 44256 32638
rect 43410 32510 43444 32544
rect 43500 32510 43534 32544
rect 43590 32510 43624 32544
rect 43680 32510 43714 32544
rect 43770 32510 43804 32544
rect 43860 32510 43894 32544
rect 43950 32510 43984 32544
rect 44040 32510 44074 32544
rect 44130 32510 44164 32544
rect 44784 33400 44818 33434
rect 44874 33400 44908 33434
rect 44964 33400 44998 33434
rect 45054 33400 45088 33434
rect 45144 33400 45178 33434
rect 45234 33400 45268 33434
rect 45324 33400 45358 33434
rect 45414 33400 45448 33434
rect 45504 33400 45538 33434
rect 44672 33343 44706 33377
rect 45562 33324 45596 33358
rect 44672 33253 44706 33287
rect 44672 33163 44706 33197
rect 44672 33073 44706 33107
rect 44672 32983 44706 33017
rect 44672 32893 44706 32927
rect 44672 32803 44706 32837
rect 44672 32713 44706 32747
rect 44672 32623 44706 32657
rect 45562 33234 45596 33268
rect 45562 33144 45596 33178
rect 45562 33054 45596 33088
rect 45562 32964 45596 32998
rect 45562 32874 45596 32908
rect 45562 32784 45596 32818
rect 45562 32694 45596 32728
rect 45562 32604 45596 32638
rect 44750 32510 44784 32544
rect 44840 32510 44874 32544
rect 44930 32510 44964 32544
rect 45020 32510 45054 32544
rect 45110 32510 45144 32544
rect 45200 32510 45234 32544
rect 45290 32510 45324 32544
rect 45380 32510 45414 32544
rect 45470 32510 45504 32544
rect 46124 33400 46158 33434
rect 46214 33400 46248 33434
rect 46304 33400 46338 33434
rect 46394 33400 46428 33434
rect 46484 33400 46518 33434
rect 46574 33400 46608 33434
rect 46664 33400 46698 33434
rect 46754 33400 46788 33434
rect 46844 33400 46878 33434
rect 46012 33343 46046 33377
rect 46902 33324 46936 33358
rect 46012 33253 46046 33287
rect 46012 33163 46046 33197
rect 46012 33073 46046 33107
rect 46012 32983 46046 33017
rect 46012 32893 46046 32927
rect 46012 32803 46046 32837
rect 46012 32713 46046 32747
rect 46012 32623 46046 32657
rect 46902 33234 46936 33268
rect 46902 33144 46936 33178
rect 46902 33054 46936 33088
rect 46902 32964 46936 32998
rect 46902 32874 46936 32908
rect 46902 32784 46936 32818
rect 46902 32694 46936 32728
rect 46902 32604 46936 32638
rect 46090 32510 46124 32544
rect 46180 32510 46214 32544
rect 46270 32510 46304 32544
rect 46360 32510 46394 32544
rect 46450 32510 46484 32544
rect 46540 32510 46574 32544
rect 46630 32510 46664 32544
rect 46720 32510 46754 32544
rect 46810 32510 46844 32544
rect 47464 33400 47498 33434
rect 47554 33400 47588 33434
rect 47644 33400 47678 33434
rect 47734 33400 47768 33434
rect 47824 33400 47858 33434
rect 47914 33400 47948 33434
rect 48004 33400 48038 33434
rect 48094 33400 48128 33434
rect 48184 33400 48218 33434
rect 47352 33343 47386 33377
rect 48242 33324 48276 33358
rect 47352 33253 47386 33287
rect 47352 33163 47386 33197
rect 47352 33073 47386 33107
rect 47352 32983 47386 33017
rect 47352 32893 47386 32927
rect 47352 32803 47386 32837
rect 47352 32713 47386 32747
rect 47352 32623 47386 32657
rect 48242 33234 48276 33268
rect 48242 33144 48276 33178
rect 48242 33054 48276 33088
rect 48242 32964 48276 32998
rect 48242 32874 48276 32908
rect 48242 32784 48276 32818
rect 48242 32694 48276 32728
rect 48242 32604 48276 32638
rect 47430 32510 47464 32544
rect 47520 32510 47554 32544
rect 47610 32510 47644 32544
rect 47700 32510 47734 32544
rect 47790 32510 47824 32544
rect 47880 32510 47914 32544
rect 47970 32510 48004 32544
rect 48060 32510 48094 32544
rect 48150 32510 48184 32544
rect 48804 33400 48838 33434
rect 48894 33400 48928 33434
rect 48984 33400 49018 33434
rect 49074 33400 49108 33434
rect 49164 33400 49198 33434
rect 49254 33400 49288 33434
rect 49344 33400 49378 33434
rect 49434 33400 49468 33434
rect 49524 33400 49558 33434
rect 48692 33343 48726 33377
rect 49582 33324 49616 33358
rect 48692 33253 48726 33287
rect 48692 33163 48726 33197
rect 48692 33073 48726 33107
rect 48692 32983 48726 33017
rect 48692 32893 48726 32927
rect 48692 32803 48726 32837
rect 48692 32713 48726 32747
rect 48692 32623 48726 32657
rect 49582 33234 49616 33268
rect 49582 33144 49616 33178
rect 49582 33054 49616 33088
rect 49582 32964 49616 32998
rect 49582 32874 49616 32908
rect 49582 32784 49616 32818
rect 49582 32694 49616 32728
rect 49582 32604 49616 32638
rect 48770 32510 48804 32544
rect 48860 32510 48894 32544
rect 48950 32510 48984 32544
rect 49040 32510 49074 32544
rect 49130 32510 49164 32544
rect 49220 32510 49254 32544
rect 49310 32510 49344 32544
rect 49400 32510 49434 32544
rect 49490 32510 49524 32544
rect 50144 33400 50178 33434
rect 50234 33400 50268 33434
rect 50324 33400 50358 33434
rect 50414 33400 50448 33434
rect 50504 33400 50538 33434
rect 50594 33400 50628 33434
rect 50684 33400 50718 33434
rect 50774 33400 50808 33434
rect 50864 33400 50898 33434
rect 50032 33343 50066 33377
rect 50922 33324 50956 33358
rect 50032 33253 50066 33287
rect 50032 33163 50066 33197
rect 50032 33073 50066 33107
rect 50032 32983 50066 33017
rect 50032 32893 50066 32927
rect 50032 32803 50066 32837
rect 50032 32713 50066 32747
rect 50032 32623 50066 32657
rect 50922 33234 50956 33268
rect 50922 33144 50956 33178
rect 50922 33054 50956 33088
rect 50922 32964 50956 32998
rect 50922 32874 50956 32908
rect 50922 32784 50956 32818
rect 50922 32694 50956 32728
rect 50922 32604 50956 32638
rect 50110 32510 50144 32544
rect 50200 32510 50234 32544
rect 50290 32510 50324 32544
rect 50380 32510 50414 32544
rect 50470 32510 50504 32544
rect 50560 32510 50594 32544
rect 50650 32510 50684 32544
rect 50740 32510 50774 32544
rect 50830 32510 50864 32544
rect 51484 33400 51518 33434
rect 51574 33400 51608 33434
rect 51664 33400 51698 33434
rect 51754 33400 51788 33434
rect 51844 33400 51878 33434
rect 51934 33400 51968 33434
rect 52024 33400 52058 33434
rect 52114 33400 52148 33434
rect 52204 33400 52238 33434
rect 51372 33343 51406 33377
rect 52262 33324 52296 33358
rect 51372 33253 51406 33287
rect 51372 33163 51406 33197
rect 51372 33073 51406 33107
rect 51372 32983 51406 33017
rect 51372 32893 51406 32927
rect 51372 32803 51406 32837
rect 51372 32713 51406 32747
rect 51372 32623 51406 32657
rect 52262 33234 52296 33268
rect 52262 33144 52296 33178
rect 52262 33054 52296 33088
rect 52262 32964 52296 32998
rect 52262 32874 52296 32908
rect 52262 32784 52296 32818
rect 52262 32694 52296 32728
rect 52262 32604 52296 32638
rect 51450 32510 51484 32544
rect 51540 32510 51574 32544
rect 51630 32510 51664 32544
rect 51720 32510 51754 32544
rect 51810 32510 51844 32544
rect 51900 32510 51934 32544
rect 51990 32510 52024 32544
rect 52080 32510 52114 32544
rect 52170 32510 52204 32544
rect 38515 30045 38549 30079
rect 37415 29995 37449 30029
rect 42104 29640 42138 29674
rect 42194 29640 42228 29674
rect 42284 29640 42318 29674
rect 42374 29640 42408 29674
rect 42464 29640 42498 29674
rect 42554 29640 42588 29674
rect 42644 29640 42678 29674
rect 42734 29640 42768 29674
rect 42824 29640 42858 29674
rect 41992 29583 42026 29617
rect 42882 29564 42916 29598
rect 41992 29493 42026 29527
rect 41992 29403 42026 29437
rect 41992 29313 42026 29347
rect 41992 29223 42026 29257
rect 41992 29133 42026 29167
rect 41992 29043 42026 29077
rect 41992 28953 42026 28987
rect 41992 28863 42026 28897
rect 42882 29474 42916 29508
rect 42882 29384 42916 29418
rect 42882 29294 42916 29328
rect 42882 29204 42916 29238
rect 42882 29114 42916 29148
rect 42882 29024 42916 29058
rect 42882 28934 42916 28968
rect 42882 28844 42916 28878
rect 42070 28750 42104 28784
rect 42160 28750 42194 28784
rect 42250 28750 42284 28784
rect 42340 28750 42374 28784
rect 42430 28750 42464 28784
rect 42520 28750 42554 28784
rect 42610 28750 42644 28784
rect 42700 28750 42734 28784
rect 42790 28750 42824 28784
rect 43444 29640 43478 29674
rect 43534 29640 43568 29674
rect 43624 29640 43658 29674
rect 43714 29640 43748 29674
rect 43804 29640 43838 29674
rect 43894 29640 43928 29674
rect 43984 29640 44018 29674
rect 44074 29640 44108 29674
rect 44164 29640 44198 29674
rect 43332 29583 43366 29617
rect 44222 29564 44256 29598
rect 43332 29493 43366 29527
rect 43332 29403 43366 29437
rect 43332 29313 43366 29347
rect 43332 29223 43366 29257
rect 43332 29133 43366 29167
rect 43332 29043 43366 29077
rect 43332 28953 43366 28987
rect 43332 28863 43366 28897
rect 44222 29474 44256 29508
rect 44222 29384 44256 29418
rect 44222 29294 44256 29328
rect 44222 29204 44256 29238
rect 44222 29114 44256 29148
rect 44222 29024 44256 29058
rect 44222 28934 44256 28968
rect 44222 28844 44256 28878
rect 43410 28750 43444 28784
rect 43500 28750 43534 28784
rect 43590 28750 43624 28784
rect 43680 28750 43714 28784
rect 43770 28750 43804 28784
rect 43860 28750 43894 28784
rect 43950 28750 43984 28784
rect 44040 28750 44074 28784
rect 44130 28750 44164 28784
rect 44784 29640 44818 29674
rect 44874 29640 44908 29674
rect 44964 29640 44998 29674
rect 45054 29640 45088 29674
rect 45144 29640 45178 29674
rect 45234 29640 45268 29674
rect 45324 29640 45358 29674
rect 45414 29640 45448 29674
rect 45504 29640 45538 29674
rect 44672 29583 44706 29617
rect 45562 29564 45596 29598
rect 44672 29493 44706 29527
rect 44672 29403 44706 29437
rect 44672 29313 44706 29347
rect 44672 29223 44706 29257
rect 44672 29133 44706 29167
rect 44672 29043 44706 29077
rect 44672 28953 44706 28987
rect 44672 28863 44706 28897
rect 45562 29474 45596 29508
rect 45562 29384 45596 29418
rect 45562 29294 45596 29328
rect 45562 29204 45596 29238
rect 45562 29114 45596 29148
rect 45562 29024 45596 29058
rect 45562 28934 45596 28968
rect 45562 28844 45596 28878
rect 44750 28750 44784 28784
rect 44840 28750 44874 28784
rect 44930 28750 44964 28784
rect 45020 28750 45054 28784
rect 45110 28750 45144 28784
rect 45200 28750 45234 28784
rect 45290 28750 45324 28784
rect 45380 28750 45414 28784
rect 45470 28750 45504 28784
rect 46124 29640 46158 29674
rect 46214 29640 46248 29674
rect 46304 29640 46338 29674
rect 46394 29640 46428 29674
rect 46484 29640 46518 29674
rect 46574 29640 46608 29674
rect 46664 29640 46698 29674
rect 46754 29640 46788 29674
rect 46844 29640 46878 29674
rect 46012 29583 46046 29617
rect 46902 29564 46936 29598
rect 46012 29493 46046 29527
rect 46012 29403 46046 29437
rect 46012 29313 46046 29347
rect 46012 29223 46046 29257
rect 46012 29133 46046 29167
rect 46012 29043 46046 29077
rect 46012 28953 46046 28987
rect 46012 28863 46046 28897
rect 46902 29474 46936 29508
rect 46902 29384 46936 29418
rect 46902 29294 46936 29328
rect 46902 29204 46936 29238
rect 46902 29114 46936 29148
rect 46902 29024 46936 29058
rect 46902 28934 46936 28968
rect 46902 28844 46936 28878
rect 46090 28750 46124 28784
rect 46180 28750 46214 28784
rect 46270 28750 46304 28784
rect 46360 28750 46394 28784
rect 46450 28750 46484 28784
rect 46540 28750 46574 28784
rect 46630 28750 46664 28784
rect 46720 28750 46754 28784
rect 46810 28750 46844 28784
rect 47464 29640 47498 29674
rect 47554 29640 47588 29674
rect 47644 29640 47678 29674
rect 47734 29640 47768 29674
rect 47824 29640 47858 29674
rect 47914 29640 47948 29674
rect 48004 29640 48038 29674
rect 48094 29640 48128 29674
rect 48184 29640 48218 29674
rect 47352 29583 47386 29617
rect 48242 29564 48276 29598
rect 47352 29493 47386 29527
rect 47352 29403 47386 29437
rect 47352 29313 47386 29347
rect 47352 29223 47386 29257
rect 47352 29133 47386 29167
rect 47352 29043 47386 29077
rect 47352 28953 47386 28987
rect 47352 28863 47386 28897
rect 48242 29474 48276 29508
rect 48242 29384 48276 29418
rect 48242 29294 48276 29328
rect 48242 29204 48276 29238
rect 48242 29114 48276 29148
rect 48242 29024 48276 29058
rect 48242 28934 48276 28968
rect 48242 28844 48276 28878
rect 47430 28750 47464 28784
rect 47520 28750 47554 28784
rect 47610 28750 47644 28784
rect 47700 28750 47734 28784
rect 47790 28750 47824 28784
rect 47880 28750 47914 28784
rect 47970 28750 48004 28784
rect 48060 28750 48094 28784
rect 48150 28750 48184 28784
rect 48804 29640 48838 29674
rect 48894 29640 48928 29674
rect 48984 29640 49018 29674
rect 49074 29640 49108 29674
rect 49164 29640 49198 29674
rect 49254 29640 49288 29674
rect 49344 29640 49378 29674
rect 49434 29640 49468 29674
rect 49524 29640 49558 29674
rect 48692 29583 48726 29617
rect 49582 29564 49616 29598
rect 48692 29493 48726 29527
rect 48692 29403 48726 29437
rect 48692 29313 48726 29347
rect 48692 29223 48726 29257
rect 48692 29133 48726 29167
rect 48692 29043 48726 29077
rect 48692 28953 48726 28987
rect 48692 28863 48726 28897
rect 49582 29474 49616 29508
rect 49582 29384 49616 29418
rect 49582 29294 49616 29328
rect 49582 29204 49616 29238
rect 49582 29114 49616 29148
rect 49582 29024 49616 29058
rect 49582 28934 49616 28968
rect 49582 28844 49616 28878
rect 48770 28750 48804 28784
rect 48860 28750 48894 28784
rect 48950 28750 48984 28784
rect 49040 28750 49074 28784
rect 49130 28750 49164 28784
rect 49220 28750 49254 28784
rect 49310 28750 49344 28784
rect 49400 28750 49434 28784
rect 49490 28750 49524 28784
rect 50144 29640 50178 29674
rect 50234 29640 50268 29674
rect 50324 29640 50358 29674
rect 50414 29640 50448 29674
rect 50504 29640 50538 29674
rect 50594 29640 50628 29674
rect 50684 29640 50718 29674
rect 50774 29640 50808 29674
rect 50864 29640 50898 29674
rect 50032 29583 50066 29617
rect 50922 29564 50956 29598
rect 50032 29493 50066 29527
rect 50032 29403 50066 29437
rect 50032 29313 50066 29347
rect 50032 29223 50066 29257
rect 50032 29133 50066 29167
rect 50032 29043 50066 29077
rect 50032 28953 50066 28987
rect 50032 28863 50066 28897
rect 50922 29474 50956 29508
rect 50922 29384 50956 29418
rect 50922 29294 50956 29328
rect 50922 29204 50956 29238
rect 50922 29114 50956 29148
rect 50922 29024 50956 29058
rect 50922 28934 50956 28968
rect 50922 28844 50956 28878
rect 50110 28750 50144 28784
rect 50200 28750 50234 28784
rect 50290 28750 50324 28784
rect 50380 28750 50414 28784
rect 50470 28750 50504 28784
rect 50560 28750 50594 28784
rect 50650 28750 50684 28784
rect 50740 28750 50774 28784
rect 50830 28750 50864 28784
rect 51484 29640 51518 29674
rect 51574 29640 51608 29674
rect 51664 29640 51698 29674
rect 51754 29640 51788 29674
rect 51844 29640 51878 29674
rect 51934 29640 51968 29674
rect 52024 29640 52058 29674
rect 52114 29640 52148 29674
rect 52204 29640 52238 29674
rect 51372 29583 51406 29617
rect 52262 29564 52296 29598
rect 51372 29493 51406 29527
rect 51372 29403 51406 29437
rect 51372 29313 51406 29347
rect 51372 29223 51406 29257
rect 51372 29133 51406 29167
rect 51372 29043 51406 29077
rect 51372 28953 51406 28987
rect 51372 28863 51406 28897
rect 52262 29474 52296 29508
rect 52262 29384 52296 29418
rect 52262 29294 52296 29328
rect 52262 29204 52296 29238
rect 52262 29114 52296 29148
rect 52262 29024 52296 29058
rect 52262 28934 52296 28968
rect 52262 28844 52296 28878
rect 51450 28750 51484 28784
rect 51540 28750 51574 28784
rect 51630 28750 51664 28784
rect 51720 28750 51754 28784
rect 51810 28750 51844 28784
rect 51900 28750 51934 28784
rect 51990 28750 52024 28784
rect 52080 28750 52114 28784
rect 52170 28750 52204 28784
rect 25873 18765 25907 18799
rect 27173 18765 27207 18799
rect 28473 18765 28507 18799
rect 29773 18765 29807 18799
rect 31073 18765 31107 18799
rect 32373 18765 32407 18799
rect 33673 18765 33707 18799
rect 34973 18765 35007 18799
rect 36273 18765 36307 18799
rect 37573 18765 37607 18799
rect 38873 18765 38907 18799
rect 40173 18765 40207 18799
rect 41473 18765 41507 18799
rect 42773 18765 42807 18799
rect 44073 18765 44107 18799
rect 45373 18765 45407 18799
rect 46673 18765 46707 18799
rect 47973 18765 48007 18799
rect 49273 18765 49307 18799
rect 50573 18765 50607 18799
rect 24773 18715 24807 18749
<< poly >>
rect 24923 48717 25323 48743
rect 25381 48717 25781 48743
rect 25839 48717 26239 48743
rect 26297 48717 26697 48743
rect 26755 48717 27155 48743
rect 27213 48717 27613 48743
rect 27671 48717 28071 48743
rect 28129 48717 28529 48743
rect 28587 48717 28987 48743
rect 29045 48717 29445 48743
rect 29503 48717 29903 48743
rect 29961 48717 30361 48743
rect 30419 48717 30819 48743
rect 30877 48717 31277 48743
rect 31335 48717 31735 48743
rect 31793 48717 32193 48743
rect 32251 48717 32651 48743
rect 32709 48717 33109 48743
rect 33167 48717 33567 48743
rect 33625 48717 34025 48743
rect 34083 48717 34483 48743
rect 34541 48717 34941 48743
rect 34999 48717 35399 48743
rect 35457 48717 35857 48743
rect 35915 48717 36315 48743
rect 36373 48717 36773 48743
rect 36831 48717 37231 48743
rect 37289 48717 37689 48743
rect 37747 48717 38147 48743
rect 38205 48717 38605 48743
rect 38663 48717 39063 48743
rect 39121 48717 39521 48743
rect 39579 48717 39979 48743
rect 40037 48717 40437 48743
rect 40495 48717 40895 48743
rect 40953 48717 41353 48743
rect 41411 48717 41811 48743
rect 41869 48717 42269 48743
rect 42327 48717 42727 48743
rect 42785 48717 43185 48743
rect 43243 48717 43643 48743
rect 43701 48717 44101 48743
rect 44159 48717 44559 48743
rect 44617 48717 45017 48743
rect 45075 48717 45475 48743
rect 45533 48717 45933 48743
rect 45991 48717 46391 48743
rect 46449 48717 46849 48743
rect 46907 48717 47307 48743
rect 47365 48717 47765 48743
rect 47823 48717 48223 48743
rect 48281 48717 48681 48743
rect 48739 48717 49139 48743
rect 49197 48717 49597 48743
rect 49655 48717 50055 48743
rect 50113 48717 50513 48743
rect 50571 48717 50971 48743
rect 51029 48717 51429 48743
rect 51487 48717 51887 48743
rect 51945 48717 52345 48743
rect 23976 48472 24376 48498
rect 23976 47646 24376 47672
rect 24124 47296 24244 47646
rect 24923 47401 25323 47427
rect 25381 47401 25781 47427
rect 25839 47401 26239 47427
rect 26297 47401 26697 47427
rect 26755 47401 27155 47427
rect 27213 47401 27613 47427
rect 27671 47401 28071 47427
rect 28129 47401 28529 47427
rect 28587 47401 28987 47427
rect 29045 47401 29445 47427
rect 29503 47401 29903 47427
rect 29961 47401 30361 47427
rect 30419 47401 30819 47427
rect 30877 47401 31277 47427
rect 31335 47401 31735 47427
rect 31793 47401 32193 47427
rect 32251 47401 32651 47427
rect 32709 47401 33109 47427
rect 33167 47401 33567 47427
rect 33625 47401 34025 47427
rect 34083 47401 34483 47427
rect 34541 47401 34941 47427
rect 34999 47401 35399 47427
rect 35457 47401 35857 47427
rect 35915 47401 36315 47427
rect 36373 47401 36773 47427
rect 36831 47401 37231 47427
rect 37289 47401 37689 47427
rect 37747 47401 38147 47427
rect 38205 47401 38605 47427
rect 38663 47401 39063 47427
rect 39121 47401 39521 47427
rect 39579 47401 39979 47427
rect 40037 47401 40437 47427
rect 40495 47401 40895 47427
rect 40953 47401 41353 47427
rect 41411 47401 41811 47427
rect 41869 47401 42269 47427
rect 42327 47401 42727 47427
rect 42785 47401 43185 47427
rect 43243 47401 43643 47427
rect 43701 47401 44101 47427
rect 44159 47401 44559 47427
rect 44617 47401 45017 47427
rect 45075 47401 45475 47427
rect 45533 47401 45933 47427
rect 45991 47401 46391 47427
rect 46449 47401 46849 47427
rect 46907 47401 47307 47427
rect 47365 47401 47765 47427
rect 47823 47401 48223 47427
rect 48281 47401 48681 47427
rect 48739 47401 49139 47427
rect 49197 47401 49597 47427
rect 49655 47401 50055 47427
rect 50113 47401 50513 47427
rect 50571 47401 50971 47427
rect 51029 47401 51429 47427
rect 51487 47401 51887 47427
rect 51945 47401 52345 47427
rect 23998 47263 24434 47296
rect 23998 47229 24101 47263
rect 24135 47229 24434 47263
rect 25070 47256 25190 47401
rect 25526 47256 25646 47401
rect 25982 47256 26102 47401
rect 26438 47256 26558 47401
rect 26894 47256 27014 47401
rect 27350 47256 27470 47401
rect 27806 47256 27926 47401
rect 28262 47256 28382 47401
rect 28718 47256 28838 47401
rect 29174 47256 29294 47401
rect 29630 47256 29750 47401
rect 30086 47256 30206 47401
rect 30542 47256 30662 47401
rect 30998 47256 31118 47401
rect 31454 47256 31574 47401
rect 31910 47256 32030 47401
rect 32366 47256 32486 47401
rect 32822 47256 32942 47401
rect 33278 47256 33398 47401
rect 33734 47256 33854 47401
rect 34190 47256 34310 47401
rect 34646 47256 34766 47401
rect 35102 47256 35222 47401
rect 35558 47256 35678 47401
rect 36014 47256 36134 47401
rect 36470 47256 36590 47401
rect 36926 47256 37046 47401
rect 37382 47256 37502 47401
rect 37838 47256 37958 47401
rect 38294 47256 38414 47401
rect 38750 47256 38870 47401
rect 39206 47256 39326 47401
rect 39662 47256 39782 47401
rect 40118 47256 40238 47401
rect 40574 47256 40694 47401
rect 41030 47256 41150 47401
rect 41486 47256 41606 47401
rect 41942 47256 42062 47401
rect 42398 47256 42518 47401
rect 42854 47256 42974 47401
rect 43310 47256 43430 47401
rect 43766 47256 43886 47401
rect 44222 47256 44342 47401
rect 44678 47256 44798 47401
rect 45134 47256 45254 47401
rect 45590 47256 45710 47401
rect 46046 47256 46166 47401
rect 46502 47256 46622 47401
rect 46958 47256 47078 47401
rect 47414 47256 47534 47401
rect 47870 47256 47990 47401
rect 48326 47256 48446 47401
rect 48782 47256 48902 47401
rect 49238 47256 49358 47401
rect 49694 47256 49814 47401
rect 50150 47256 50270 47401
rect 50606 47256 50726 47401
rect 51062 47256 51182 47401
rect 51518 47256 51638 47401
rect 51974 47256 52094 47401
rect 23998 47196 24434 47229
rect 24830 47223 52438 47256
rect 24830 47189 25013 47223
rect 25047 47189 25413 47223
rect 25447 47189 25813 47223
rect 25847 47189 26213 47223
rect 26247 47189 26613 47223
rect 26647 47189 27013 47223
rect 27047 47189 27413 47223
rect 27447 47189 27813 47223
rect 27847 47189 28213 47223
rect 28247 47189 28613 47223
rect 28647 47189 29013 47223
rect 29047 47189 29413 47223
rect 29447 47189 29813 47223
rect 29847 47189 30213 47223
rect 30247 47189 30613 47223
rect 30647 47189 31013 47223
rect 31047 47189 31413 47223
rect 31447 47189 31813 47223
rect 31847 47189 32213 47223
rect 32247 47189 32613 47223
rect 32647 47189 33013 47223
rect 33047 47189 33413 47223
rect 33447 47189 33813 47223
rect 33847 47189 34213 47223
rect 34247 47189 34613 47223
rect 34647 47189 35013 47223
rect 35047 47189 35413 47223
rect 35447 47189 35813 47223
rect 35847 47189 36213 47223
rect 36247 47189 36613 47223
rect 36647 47189 37013 47223
rect 37047 47189 37413 47223
rect 37447 47189 37813 47223
rect 37847 47189 38213 47223
rect 38247 47189 38613 47223
rect 38647 47189 39013 47223
rect 39047 47189 39413 47223
rect 39447 47189 39813 47223
rect 39847 47189 40213 47223
rect 40247 47189 40613 47223
rect 40647 47189 41013 47223
rect 41047 47189 41413 47223
rect 41447 47189 41813 47223
rect 41847 47189 42213 47223
rect 42247 47189 42613 47223
rect 42647 47189 43013 47223
rect 43047 47189 43413 47223
rect 43447 47189 43813 47223
rect 43847 47189 44213 47223
rect 44247 47189 44613 47223
rect 44647 47189 45013 47223
rect 45047 47189 45413 47223
rect 45447 47189 45813 47223
rect 45847 47189 46213 47223
rect 46247 47189 46613 47223
rect 46647 47189 47013 47223
rect 47047 47189 47413 47223
rect 47447 47189 47813 47223
rect 47847 47189 48213 47223
rect 48247 47189 48613 47223
rect 48647 47189 49013 47223
rect 49047 47189 49413 47223
rect 49447 47189 49813 47223
rect 49847 47189 50213 47223
rect 50247 47189 50613 47223
rect 50647 47189 51013 47223
rect 51047 47189 51413 47223
rect 51447 47189 51813 47223
rect 51847 47189 52213 47223
rect 52247 47189 52438 47223
rect 24830 47156 52438 47189
rect 15123 44957 15523 44983
rect 15581 44957 15981 44983
rect 16039 44957 16439 44983
rect 16497 44957 16897 44983
rect 16955 44957 17355 44983
rect 17413 44957 17813 44983
rect 17871 44957 18271 44983
rect 18329 44957 18729 44983
rect 18787 44957 19187 44983
rect 19245 44957 19645 44983
rect 19703 44957 20103 44983
rect 20161 44957 20561 44983
rect 20619 44957 21019 44983
rect 21077 44957 21477 44983
rect 21535 44957 21935 44983
rect 21993 44957 22393 44983
rect 22451 44957 22851 44983
rect 22909 44957 23309 44983
rect 23367 44957 23767 44983
rect 23825 44957 24225 44983
rect 24283 44957 24683 44983
rect 24741 44957 25141 44983
rect 25199 44957 25599 44983
rect 25657 44957 26057 44983
rect 26115 44957 26515 44983
rect 26573 44957 26973 44983
rect 27031 44957 27431 44983
rect 27489 44957 27889 44983
rect 27947 44957 28347 44983
rect 28405 44957 28805 44983
rect 28863 44957 29263 44983
rect 29321 44957 29721 44983
rect 29779 44957 30179 44983
rect 30237 44957 30637 44983
rect 30695 44957 31095 44983
rect 31153 44957 31553 44983
rect 31611 44957 32011 44983
rect 32069 44957 32469 44983
rect 32527 44957 32927 44983
rect 32985 44957 33385 44983
rect 33443 44957 33843 44983
rect 33901 44957 34301 44983
rect 34359 44957 34759 44983
rect 34817 44957 35217 44983
rect 35275 44957 35675 44983
rect 35733 44957 36133 44983
rect 36191 44957 36591 44983
rect 36649 44957 37049 44983
rect 37107 44957 37507 44983
rect 37565 44957 37965 44983
rect 38023 44957 38423 44983
rect 38481 44957 38881 44983
rect 38939 44957 39339 44983
rect 39397 44957 39797 44983
rect 39855 44957 40255 44983
rect 40313 44957 40713 44983
rect 40771 44957 41171 44983
rect 41229 44957 41629 44983
rect 41687 44957 42087 44983
rect 42145 44957 42545 44983
rect 14176 44712 14576 44738
rect 14176 43886 14576 43912
rect 14324 43536 14444 43886
rect 15123 43641 15523 43667
rect 15581 43641 15981 43667
rect 16039 43641 16439 43667
rect 16497 43641 16897 43667
rect 16955 43641 17355 43667
rect 17413 43641 17813 43667
rect 17871 43641 18271 43667
rect 18329 43641 18729 43667
rect 18787 43641 19187 43667
rect 19245 43641 19645 43667
rect 19703 43641 20103 43667
rect 20161 43641 20561 43667
rect 20619 43641 21019 43667
rect 21077 43641 21477 43667
rect 21535 43641 21935 43667
rect 21993 43641 22393 43667
rect 22451 43641 22851 43667
rect 22909 43641 23309 43667
rect 23367 43641 23767 43667
rect 23825 43641 24225 43667
rect 24283 43641 24683 43667
rect 24741 43641 25141 43667
rect 25199 43641 25599 43667
rect 25657 43641 26057 43667
rect 26115 43641 26515 43667
rect 26573 43641 26973 43667
rect 27031 43641 27431 43667
rect 27489 43641 27889 43667
rect 27947 43641 28347 43667
rect 28405 43641 28805 43667
rect 28863 43641 29263 43667
rect 29321 43641 29721 43667
rect 29779 43641 30179 43667
rect 30237 43641 30637 43667
rect 30695 43641 31095 43667
rect 31153 43641 31553 43667
rect 31611 43641 32011 43667
rect 32069 43641 32469 43667
rect 32527 43641 32927 43667
rect 32985 43641 33385 43667
rect 33443 43641 33843 43667
rect 33901 43641 34301 43667
rect 34359 43641 34759 43667
rect 34817 43641 35217 43667
rect 35275 43641 35675 43667
rect 35733 43641 36133 43667
rect 36191 43641 36591 43667
rect 36649 43641 37049 43667
rect 37107 43641 37507 43667
rect 37565 43641 37965 43667
rect 38023 43641 38423 43667
rect 38481 43641 38881 43667
rect 38939 43641 39339 43667
rect 39397 43641 39797 43667
rect 39855 43641 40255 43667
rect 40313 43641 40713 43667
rect 40771 43641 41171 43667
rect 41229 43641 41629 43667
rect 41687 43641 42087 43667
rect 42145 43641 42545 43667
rect 14198 43503 14634 43536
rect 14198 43469 14301 43503
rect 14335 43469 14634 43503
rect 15270 43496 15390 43641
rect 15726 43496 15846 43641
rect 16182 43496 16302 43641
rect 16638 43496 16758 43641
rect 17094 43496 17214 43641
rect 17550 43496 17670 43641
rect 18006 43496 18126 43641
rect 18462 43496 18582 43641
rect 18918 43496 19038 43641
rect 19374 43496 19494 43641
rect 19830 43496 19950 43641
rect 20286 43496 20406 43641
rect 20742 43496 20862 43641
rect 21198 43496 21318 43641
rect 21654 43496 21774 43641
rect 22110 43496 22230 43641
rect 22566 43496 22686 43641
rect 23022 43496 23142 43641
rect 23478 43496 23598 43641
rect 23934 43496 24054 43641
rect 24390 43496 24510 43641
rect 24846 43496 24966 43641
rect 25302 43496 25422 43641
rect 25758 43496 25878 43641
rect 26214 43496 26334 43641
rect 26670 43496 26790 43641
rect 27126 43496 27246 43641
rect 27582 43496 27702 43641
rect 28038 43496 28158 43641
rect 28494 43496 28614 43641
rect 28950 43496 29070 43641
rect 29406 43496 29526 43641
rect 29862 43496 29982 43641
rect 30318 43496 30438 43641
rect 30774 43496 30894 43641
rect 31230 43496 31350 43641
rect 31686 43496 31806 43641
rect 32142 43496 32262 43641
rect 32598 43496 32718 43641
rect 33054 43496 33174 43641
rect 33510 43496 33630 43641
rect 33966 43496 34086 43641
rect 34422 43496 34542 43641
rect 34878 43496 34998 43641
rect 35334 43496 35454 43641
rect 35790 43496 35910 43641
rect 36246 43496 36366 43641
rect 36702 43496 36822 43641
rect 37158 43496 37278 43641
rect 37614 43496 37734 43641
rect 38070 43496 38190 43641
rect 38526 43496 38646 43641
rect 38982 43496 39102 43641
rect 39438 43496 39558 43641
rect 39894 43496 40014 43641
rect 40350 43496 40470 43641
rect 40806 43496 40926 43641
rect 41262 43496 41382 43641
rect 41718 43496 41838 43641
rect 42174 43496 42294 43641
rect 14198 43436 14634 43469
rect 15030 43463 42638 43496
rect 15030 43429 15213 43463
rect 15247 43429 15613 43463
rect 15647 43429 16013 43463
rect 16047 43429 16413 43463
rect 16447 43429 16813 43463
rect 16847 43429 17213 43463
rect 17247 43429 17613 43463
rect 17647 43429 18013 43463
rect 18047 43429 18413 43463
rect 18447 43429 18813 43463
rect 18847 43429 19213 43463
rect 19247 43429 19613 43463
rect 19647 43429 20013 43463
rect 20047 43429 20413 43463
rect 20447 43429 20813 43463
rect 20847 43429 21213 43463
rect 21247 43429 21613 43463
rect 21647 43429 22013 43463
rect 22047 43429 22413 43463
rect 22447 43429 22813 43463
rect 22847 43429 23213 43463
rect 23247 43429 23613 43463
rect 23647 43429 24013 43463
rect 24047 43429 24413 43463
rect 24447 43429 24813 43463
rect 24847 43429 25213 43463
rect 25247 43429 25613 43463
rect 25647 43429 26013 43463
rect 26047 43429 26413 43463
rect 26447 43429 26813 43463
rect 26847 43429 27213 43463
rect 27247 43429 27613 43463
rect 27647 43429 28013 43463
rect 28047 43429 28413 43463
rect 28447 43429 28813 43463
rect 28847 43429 29213 43463
rect 29247 43429 29613 43463
rect 29647 43429 30013 43463
rect 30047 43429 30413 43463
rect 30447 43429 30813 43463
rect 30847 43429 31213 43463
rect 31247 43429 31613 43463
rect 31647 43429 32013 43463
rect 32047 43429 32413 43463
rect 32447 43429 32813 43463
rect 32847 43429 33213 43463
rect 33247 43429 33613 43463
rect 33647 43429 34013 43463
rect 34047 43429 34413 43463
rect 34447 43429 34813 43463
rect 34847 43429 35213 43463
rect 35247 43429 35613 43463
rect 35647 43429 36013 43463
rect 36047 43429 36413 43463
rect 36447 43429 36813 43463
rect 36847 43429 37213 43463
rect 37247 43429 37613 43463
rect 37647 43429 38013 43463
rect 38047 43429 38413 43463
rect 38447 43429 38813 43463
rect 38847 43429 39213 43463
rect 39247 43429 39613 43463
rect 39647 43429 40013 43463
rect 40047 43429 40413 43463
rect 40447 43429 40813 43463
rect 40847 43429 41213 43463
rect 41247 43429 41613 43463
rect 41647 43429 42013 43463
rect 42047 43429 42413 43463
rect 42447 43429 42638 43463
rect 15030 43396 42638 43429
rect 22767 41197 23167 41223
rect 23225 41197 23625 41223
rect 23683 41197 24083 41223
rect 24141 41197 24541 41223
rect 24599 41197 24999 41223
rect 25057 41197 25457 41223
rect 25515 41197 25915 41223
rect 25973 41197 26373 41223
rect 26431 41197 26831 41223
rect 26889 41197 27289 41223
rect 27347 41197 27747 41223
rect 27805 41197 28205 41223
rect 29431 41197 29831 41223
rect 29889 41197 30289 41223
rect 30347 41197 30747 41223
rect 30805 41197 31205 41223
rect 31263 41197 31663 41223
rect 31721 41197 32121 41223
rect 32179 41197 32579 41223
rect 32637 41197 33037 41223
rect 33095 41197 33495 41223
rect 33553 41197 33953 41223
rect 34011 41197 34411 41223
rect 34469 41197 34869 41223
rect 37334 40952 37734 40978
rect 37792 40952 38192 40978
rect 38250 40952 38650 40978
rect 38708 40952 39108 40978
rect 39166 40952 39566 40978
rect 39624 40952 40024 40978
rect 40082 40952 40482 40978
rect 40540 40952 40940 40978
rect 40998 40952 41398 40978
rect 37334 40126 37734 40152
rect 37792 40126 38192 40152
rect 38250 40126 38650 40152
rect 38708 40126 39108 40152
rect 39166 40126 39566 40152
rect 39624 40126 40024 40152
rect 40082 40126 40482 40152
rect 40540 40126 40940 40152
rect 40998 40126 41398 40152
rect 37482 39936 37602 40126
rect 37938 39936 38058 40126
rect 38394 39936 38514 40126
rect 38850 39936 38970 40126
rect 39306 39936 39426 40126
rect 39762 39936 39882 40126
rect 40218 39936 40338 40126
rect 40674 39936 40794 40126
rect 41130 39936 41250 40126
rect 22767 39881 23167 39907
rect 23225 39881 23625 39907
rect 23683 39881 24083 39907
rect 24141 39881 24541 39907
rect 24599 39881 24999 39907
rect 25057 39881 25457 39907
rect 25515 39881 25915 39907
rect 25973 39881 26373 39907
rect 26431 39881 26831 39907
rect 26889 39881 27289 39907
rect 27347 39881 27747 39907
rect 27805 39881 28205 39907
rect 29431 39881 29831 39907
rect 29889 39881 30289 39907
rect 30347 39881 30747 39907
rect 30805 39881 31205 39907
rect 31263 39881 31663 39907
rect 31721 39881 32121 39907
rect 32179 39881 32579 39907
rect 32637 39881 33037 39907
rect 33095 39881 33495 39907
rect 33553 39881 33953 39907
rect 34011 39881 34411 39907
rect 34469 39881 34869 39907
rect 37356 39903 41456 39936
rect 22914 39736 23034 39881
rect 23370 39736 23490 39881
rect 23826 39736 23946 39881
rect 24282 39736 24402 39881
rect 24738 39736 24858 39881
rect 25194 39736 25314 39881
rect 25650 39736 25770 39881
rect 26106 39736 26226 39881
rect 26562 39736 26682 39881
rect 27018 39736 27138 39881
rect 27474 39736 27594 39881
rect 27930 39736 28050 39881
rect 29578 39736 29698 39881
rect 30034 39736 30154 39881
rect 30490 39736 30610 39881
rect 30946 39736 31066 39881
rect 31402 39736 31522 39881
rect 31858 39736 31978 39881
rect 32314 39736 32434 39881
rect 32770 39736 32890 39881
rect 33226 39736 33346 39881
rect 33682 39736 33802 39881
rect 34138 39736 34258 39881
rect 34594 39736 34714 39881
rect 37356 39869 37459 39903
rect 37493 39869 37859 39903
rect 37893 39869 38259 39903
rect 38293 39869 38659 39903
rect 38693 39869 39059 39903
rect 39093 39869 39459 39903
rect 39493 39869 39859 39903
rect 39893 39869 40259 39903
rect 40293 39869 40659 39903
rect 40693 39869 41059 39903
rect 41093 39869 41456 39903
rect 37356 39836 41456 39869
rect 22674 39703 28298 39736
rect 22674 39669 22857 39703
rect 22891 39669 23257 39703
rect 23291 39669 23657 39703
rect 23691 39669 24057 39703
rect 24091 39669 24457 39703
rect 24491 39669 24857 39703
rect 24891 39669 25257 39703
rect 25291 39669 25657 39703
rect 25691 39669 26057 39703
rect 26091 39669 26457 39703
rect 26491 39669 26857 39703
rect 26891 39669 27257 39703
rect 27291 39669 27657 39703
rect 27691 39669 28057 39703
rect 28091 39669 28298 39703
rect 22674 39636 28298 39669
rect 29338 39703 34962 39736
rect 29338 39669 29521 39703
rect 29555 39669 29921 39703
rect 29955 39669 30321 39703
rect 30355 39669 30721 39703
rect 30755 39669 31121 39703
rect 31155 39669 31521 39703
rect 31555 39669 31921 39703
rect 31955 39669 32321 39703
rect 32355 39669 32721 39703
rect 32755 39669 33121 39703
rect 33155 39669 33521 39703
rect 33555 39669 33921 39703
rect 33955 39669 34321 39703
rect 34355 39669 34721 39703
rect 34755 39669 34962 39703
rect 29338 39636 34962 39669
rect 37565 37437 37965 37463
rect 38023 37437 38423 37463
rect 38481 37437 38881 37463
rect 38939 37437 39339 37463
rect 39397 37437 39797 37463
rect 39855 37437 40255 37463
rect 25476 37192 25876 37218
rect 25934 37192 26334 37218
rect 26392 37192 26792 37218
rect 26850 37192 27250 37218
rect 27308 37192 27708 37218
rect 27766 37192 28166 37218
rect 28224 37192 28624 37218
rect 28682 37192 29082 37218
rect 29140 37192 29540 37218
rect 25476 36366 25876 36392
rect 25934 36366 26334 36392
rect 26392 36366 26792 36392
rect 26850 36366 27250 36392
rect 27308 36366 27708 36392
rect 27766 36366 28166 36392
rect 28224 36366 28624 36392
rect 28682 36366 29082 36392
rect 29140 36366 29540 36392
rect 25624 36176 25744 36366
rect 26080 36176 26200 36366
rect 26536 36176 26656 36366
rect 26992 36176 27112 36366
rect 27448 36176 27568 36366
rect 27904 36176 28024 36366
rect 28360 36176 28480 36366
rect 28816 36176 28936 36366
rect 29272 36176 29392 36366
rect 25498 36143 29598 36176
rect 25498 36109 25601 36143
rect 25635 36109 26001 36143
rect 26035 36109 26401 36143
rect 26435 36109 26801 36143
rect 26835 36109 27201 36143
rect 27235 36109 27601 36143
rect 27635 36109 28001 36143
rect 28035 36109 28401 36143
rect 28435 36109 28801 36143
rect 28835 36109 29201 36143
rect 29235 36109 29598 36143
rect 37565 36121 37965 36147
rect 38023 36121 38423 36147
rect 38481 36121 38881 36147
rect 38939 36121 39339 36147
rect 39397 36121 39797 36147
rect 39855 36121 40255 36147
rect 25498 36076 29598 36109
rect 37712 35976 37832 36121
rect 38168 35976 38288 36121
rect 38624 35976 38744 36121
rect 39080 35976 39200 36121
rect 39536 35976 39656 36121
rect 39992 35976 40112 36121
rect 37472 35943 40348 35976
rect 37472 35909 37655 35943
rect 37689 35909 38055 35943
rect 38089 35909 38455 35943
rect 38489 35909 38855 35943
rect 38889 35909 39255 35943
rect 39289 35909 39655 35943
rect 39689 35909 40055 35943
rect 40089 35909 40348 35943
rect 37472 35876 40348 35909
rect 37565 29917 37965 29943
rect 38023 29917 38423 29943
rect 38481 29917 38881 29943
rect 38939 29917 39339 29943
rect 39397 29917 39797 29943
rect 39855 29917 40255 29943
rect 37565 28601 37965 28627
rect 38023 28601 38423 28627
rect 38481 28601 38881 28627
rect 38939 28601 39339 28627
rect 39397 28601 39797 28627
rect 39855 28601 40255 28627
rect 37712 28456 37832 28601
rect 38168 28456 38288 28601
rect 38624 28456 38744 28601
rect 39080 28456 39200 28601
rect 39536 28456 39656 28601
rect 39992 28456 40112 28601
rect 37472 28423 40348 28456
rect 37472 28389 37655 28423
rect 37689 28389 38055 28423
rect 38089 28389 38455 28423
rect 38489 28389 38855 28423
rect 38889 28389 39255 28423
rect 39289 28389 39655 28423
rect 39689 28389 40055 28423
rect 40089 28389 40348 28423
rect 37472 28356 40348 28389
rect 25476 25912 25876 25938
rect 25934 25912 26334 25938
rect 26392 25912 26792 25938
rect 26850 25912 27250 25938
rect 27308 25912 27708 25938
rect 27766 25912 28166 25938
rect 28224 25912 28624 25938
rect 28682 25912 29082 25938
rect 29140 25912 29540 25938
rect 25476 25086 25876 25112
rect 25934 25086 26334 25112
rect 26392 25086 26792 25112
rect 26850 25086 27250 25112
rect 27308 25086 27708 25112
rect 27766 25086 28166 25112
rect 28224 25086 28624 25112
rect 28682 25086 29082 25112
rect 29140 25086 29540 25112
rect 25624 24896 25744 25086
rect 26080 24896 26200 25086
rect 26536 24896 26656 25086
rect 26992 24896 27112 25086
rect 27448 24896 27568 25086
rect 27904 24896 28024 25086
rect 28360 24896 28480 25086
rect 28816 24896 28936 25086
rect 29272 24896 29392 25086
rect 25498 24863 29598 24896
rect 25498 24829 25601 24863
rect 25635 24829 26001 24863
rect 26035 24829 26401 24863
rect 26435 24829 26801 24863
rect 26835 24829 27201 24863
rect 27235 24829 27601 24863
rect 27635 24829 28001 24863
rect 28035 24829 28401 24863
rect 28435 24829 28801 24863
rect 28835 24829 29201 24863
rect 29235 24829 29598 24863
rect 25498 24796 29598 24829
rect 24923 18637 25323 18663
rect 25381 18637 25781 18663
rect 25839 18637 26239 18663
rect 26297 18637 26697 18663
rect 26755 18637 27155 18663
rect 27213 18637 27613 18663
rect 27671 18637 28071 18663
rect 28129 18637 28529 18663
rect 28587 18637 28987 18663
rect 29045 18637 29445 18663
rect 29503 18637 29903 18663
rect 29961 18637 30361 18663
rect 30419 18637 30819 18663
rect 30877 18637 31277 18663
rect 31335 18637 31735 18663
rect 31793 18637 32193 18663
rect 32251 18637 32651 18663
rect 32709 18637 33109 18663
rect 33167 18637 33567 18663
rect 33625 18637 34025 18663
rect 34083 18637 34483 18663
rect 34541 18637 34941 18663
rect 34999 18637 35399 18663
rect 35457 18637 35857 18663
rect 35915 18637 36315 18663
rect 36373 18637 36773 18663
rect 36831 18637 37231 18663
rect 37289 18637 37689 18663
rect 37747 18637 38147 18663
rect 38205 18637 38605 18663
rect 38663 18637 39063 18663
rect 39121 18637 39521 18663
rect 39579 18637 39979 18663
rect 40037 18637 40437 18663
rect 40495 18637 40895 18663
rect 40953 18637 41353 18663
rect 41411 18637 41811 18663
rect 41869 18637 42269 18663
rect 42327 18637 42727 18663
rect 42785 18637 43185 18663
rect 43243 18637 43643 18663
rect 43701 18637 44101 18663
rect 44159 18637 44559 18663
rect 44617 18637 45017 18663
rect 45075 18637 45475 18663
rect 45533 18637 45933 18663
rect 45991 18637 46391 18663
rect 46449 18637 46849 18663
rect 46907 18637 47307 18663
rect 47365 18637 47765 18663
rect 47823 18637 48223 18663
rect 48281 18637 48681 18663
rect 48739 18637 49139 18663
rect 49197 18637 49597 18663
rect 49655 18637 50055 18663
rect 50113 18637 50513 18663
rect 50571 18637 50971 18663
rect 51029 18637 51429 18663
rect 51487 18637 51887 18663
rect 51945 18637 52345 18663
rect 24923 17321 25323 17347
rect 25381 17321 25781 17347
rect 25839 17321 26239 17347
rect 26297 17321 26697 17347
rect 26755 17321 27155 17347
rect 27213 17321 27613 17347
rect 27671 17321 28071 17347
rect 28129 17321 28529 17347
rect 28587 17321 28987 17347
rect 29045 17321 29445 17347
rect 29503 17321 29903 17347
rect 29961 17321 30361 17347
rect 30419 17321 30819 17347
rect 30877 17321 31277 17347
rect 31335 17321 31735 17347
rect 31793 17321 32193 17347
rect 32251 17321 32651 17347
rect 32709 17321 33109 17347
rect 33167 17321 33567 17347
rect 33625 17321 34025 17347
rect 34083 17321 34483 17347
rect 34541 17321 34941 17347
rect 34999 17321 35399 17347
rect 35457 17321 35857 17347
rect 35915 17321 36315 17347
rect 36373 17321 36773 17347
rect 36831 17321 37231 17347
rect 37289 17321 37689 17347
rect 37747 17321 38147 17347
rect 38205 17321 38605 17347
rect 38663 17321 39063 17347
rect 39121 17321 39521 17347
rect 39579 17321 39979 17347
rect 40037 17321 40437 17347
rect 40495 17321 40895 17347
rect 40953 17321 41353 17347
rect 41411 17321 41811 17347
rect 41869 17321 42269 17347
rect 42327 17321 42727 17347
rect 42785 17321 43185 17347
rect 43243 17321 43643 17347
rect 43701 17321 44101 17347
rect 44159 17321 44559 17347
rect 44617 17321 45017 17347
rect 45075 17321 45475 17347
rect 45533 17321 45933 17347
rect 45991 17321 46391 17347
rect 46449 17321 46849 17347
rect 46907 17321 47307 17347
rect 47365 17321 47765 17347
rect 47823 17321 48223 17347
rect 48281 17321 48681 17347
rect 48739 17321 49139 17347
rect 49197 17321 49597 17347
rect 49655 17321 50055 17347
rect 50113 17321 50513 17347
rect 50571 17321 50971 17347
rect 51029 17321 51429 17347
rect 51487 17321 51887 17347
rect 51945 17321 52345 17347
rect 25070 17176 25190 17321
rect 25526 17176 25646 17321
rect 25982 17176 26102 17321
rect 26438 17176 26558 17321
rect 26894 17176 27014 17321
rect 27350 17176 27470 17321
rect 27806 17176 27926 17321
rect 28262 17176 28382 17321
rect 28718 17176 28838 17321
rect 29174 17176 29294 17321
rect 29630 17176 29750 17321
rect 30086 17176 30206 17321
rect 30542 17176 30662 17321
rect 30998 17176 31118 17321
rect 31454 17176 31574 17321
rect 31910 17176 32030 17321
rect 32366 17176 32486 17321
rect 32822 17176 32942 17321
rect 33278 17176 33398 17321
rect 33734 17176 33854 17321
rect 34190 17176 34310 17321
rect 34646 17176 34766 17321
rect 35102 17176 35222 17321
rect 35558 17176 35678 17321
rect 36014 17176 36134 17321
rect 36470 17176 36590 17321
rect 36926 17176 37046 17321
rect 37382 17176 37502 17321
rect 37838 17176 37958 17321
rect 38294 17176 38414 17321
rect 38750 17176 38870 17321
rect 39206 17176 39326 17321
rect 39662 17176 39782 17321
rect 40118 17176 40238 17321
rect 40574 17176 40694 17321
rect 41030 17176 41150 17321
rect 41486 17176 41606 17321
rect 41942 17176 42062 17321
rect 42398 17176 42518 17321
rect 42854 17176 42974 17321
rect 43310 17176 43430 17321
rect 43766 17176 43886 17321
rect 44222 17176 44342 17321
rect 44678 17176 44798 17321
rect 45134 17176 45254 17321
rect 45590 17176 45710 17321
rect 46046 17176 46166 17321
rect 46502 17176 46622 17321
rect 46958 17176 47078 17321
rect 47414 17176 47534 17321
rect 47870 17176 47990 17321
rect 48326 17176 48446 17321
rect 48782 17176 48902 17321
rect 49238 17176 49358 17321
rect 49694 17176 49814 17321
rect 50150 17176 50270 17321
rect 50606 17176 50726 17321
rect 51062 17176 51182 17321
rect 51518 17176 51638 17321
rect 51974 17176 52094 17321
rect 24830 17143 52438 17176
rect 24830 17109 25013 17143
rect 25047 17109 25413 17143
rect 25447 17109 25813 17143
rect 25847 17109 26213 17143
rect 26247 17109 26613 17143
rect 26647 17109 27013 17143
rect 27047 17109 27413 17143
rect 27447 17109 27813 17143
rect 27847 17109 28213 17143
rect 28247 17109 28613 17143
rect 28647 17109 29013 17143
rect 29047 17109 29413 17143
rect 29447 17109 29813 17143
rect 29847 17109 30213 17143
rect 30247 17109 30613 17143
rect 30647 17109 31013 17143
rect 31047 17109 31413 17143
rect 31447 17109 31813 17143
rect 31847 17109 32213 17143
rect 32247 17109 32613 17143
rect 32647 17109 33013 17143
rect 33047 17109 33413 17143
rect 33447 17109 33813 17143
rect 33847 17109 34213 17143
rect 34247 17109 34613 17143
rect 34647 17109 35013 17143
rect 35047 17109 35413 17143
rect 35447 17109 35813 17143
rect 35847 17109 36213 17143
rect 36247 17109 36613 17143
rect 36647 17109 37013 17143
rect 37047 17109 37413 17143
rect 37447 17109 37813 17143
rect 37847 17109 38213 17143
rect 38247 17109 38613 17143
rect 38647 17109 39013 17143
rect 39047 17109 39413 17143
rect 39447 17109 39813 17143
rect 39847 17109 40213 17143
rect 40247 17109 40613 17143
rect 40647 17109 41013 17143
rect 41047 17109 41413 17143
rect 41447 17109 41813 17143
rect 41847 17109 42213 17143
rect 42247 17109 42613 17143
rect 42647 17109 43013 17143
rect 43047 17109 43413 17143
rect 43447 17109 43813 17143
rect 43847 17109 44213 17143
rect 44247 17109 44613 17143
rect 44647 17109 45013 17143
rect 45047 17109 45413 17143
rect 45447 17109 45813 17143
rect 45847 17109 46213 17143
rect 46247 17109 46613 17143
rect 46647 17109 47013 17143
rect 47047 17109 47413 17143
rect 47447 17109 47813 17143
rect 47847 17109 48213 17143
rect 48247 17109 48613 17143
rect 48647 17109 49013 17143
rect 49047 17109 49413 17143
rect 49447 17109 49813 17143
rect 49847 17109 50213 17143
rect 50247 17109 50613 17143
rect 50647 17109 51013 17143
rect 51047 17109 51413 17143
rect 51447 17109 51813 17143
rect 51847 17109 52213 17143
rect 52247 17109 52438 17143
rect 24830 17076 52438 17109
<< polycont >>
rect 24101 47229 24135 47263
rect 25013 47189 25047 47223
rect 25413 47189 25447 47223
rect 25813 47189 25847 47223
rect 26213 47189 26247 47223
rect 26613 47189 26647 47223
rect 27013 47189 27047 47223
rect 27413 47189 27447 47223
rect 27813 47189 27847 47223
rect 28213 47189 28247 47223
rect 28613 47189 28647 47223
rect 29013 47189 29047 47223
rect 29413 47189 29447 47223
rect 29813 47189 29847 47223
rect 30213 47189 30247 47223
rect 30613 47189 30647 47223
rect 31013 47189 31047 47223
rect 31413 47189 31447 47223
rect 31813 47189 31847 47223
rect 32213 47189 32247 47223
rect 32613 47189 32647 47223
rect 33013 47189 33047 47223
rect 33413 47189 33447 47223
rect 33813 47189 33847 47223
rect 34213 47189 34247 47223
rect 34613 47189 34647 47223
rect 35013 47189 35047 47223
rect 35413 47189 35447 47223
rect 35813 47189 35847 47223
rect 36213 47189 36247 47223
rect 36613 47189 36647 47223
rect 37013 47189 37047 47223
rect 37413 47189 37447 47223
rect 37813 47189 37847 47223
rect 38213 47189 38247 47223
rect 38613 47189 38647 47223
rect 39013 47189 39047 47223
rect 39413 47189 39447 47223
rect 39813 47189 39847 47223
rect 40213 47189 40247 47223
rect 40613 47189 40647 47223
rect 41013 47189 41047 47223
rect 41413 47189 41447 47223
rect 41813 47189 41847 47223
rect 42213 47189 42247 47223
rect 42613 47189 42647 47223
rect 43013 47189 43047 47223
rect 43413 47189 43447 47223
rect 43813 47189 43847 47223
rect 44213 47189 44247 47223
rect 44613 47189 44647 47223
rect 45013 47189 45047 47223
rect 45413 47189 45447 47223
rect 45813 47189 45847 47223
rect 46213 47189 46247 47223
rect 46613 47189 46647 47223
rect 47013 47189 47047 47223
rect 47413 47189 47447 47223
rect 47813 47189 47847 47223
rect 48213 47189 48247 47223
rect 48613 47189 48647 47223
rect 49013 47189 49047 47223
rect 49413 47189 49447 47223
rect 49813 47189 49847 47223
rect 50213 47189 50247 47223
rect 50613 47189 50647 47223
rect 51013 47189 51047 47223
rect 51413 47189 51447 47223
rect 51813 47189 51847 47223
rect 52213 47189 52247 47223
rect 14301 43469 14335 43503
rect 15213 43429 15247 43463
rect 15613 43429 15647 43463
rect 16013 43429 16047 43463
rect 16413 43429 16447 43463
rect 16813 43429 16847 43463
rect 17213 43429 17247 43463
rect 17613 43429 17647 43463
rect 18013 43429 18047 43463
rect 18413 43429 18447 43463
rect 18813 43429 18847 43463
rect 19213 43429 19247 43463
rect 19613 43429 19647 43463
rect 20013 43429 20047 43463
rect 20413 43429 20447 43463
rect 20813 43429 20847 43463
rect 21213 43429 21247 43463
rect 21613 43429 21647 43463
rect 22013 43429 22047 43463
rect 22413 43429 22447 43463
rect 22813 43429 22847 43463
rect 23213 43429 23247 43463
rect 23613 43429 23647 43463
rect 24013 43429 24047 43463
rect 24413 43429 24447 43463
rect 24813 43429 24847 43463
rect 25213 43429 25247 43463
rect 25613 43429 25647 43463
rect 26013 43429 26047 43463
rect 26413 43429 26447 43463
rect 26813 43429 26847 43463
rect 27213 43429 27247 43463
rect 27613 43429 27647 43463
rect 28013 43429 28047 43463
rect 28413 43429 28447 43463
rect 28813 43429 28847 43463
rect 29213 43429 29247 43463
rect 29613 43429 29647 43463
rect 30013 43429 30047 43463
rect 30413 43429 30447 43463
rect 30813 43429 30847 43463
rect 31213 43429 31247 43463
rect 31613 43429 31647 43463
rect 32013 43429 32047 43463
rect 32413 43429 32447 43463
rect 32813 43429 32847 43463
rect 33213 43429 33247 43463
rect 33613 43429 33647 43463
rect 34013 43429 34047 43463
rect 34413 43429 34447 43463
rect 34813 43429 34847 43463
rect 35213 43429 35247 43463
rect 35613 43429 35647 43463
rect 36013 43429 36047 43463
rect 36413 43429 36447 43463
rect 36813 43429 36847 43463
rect 37213 43429 37247 43463
rect 37613 43429 37647 43463
rect 38013 43429 38047 43463
rect 38413 43429 38447 43463
rect 38813 43429 38847 43463
rect 39213 43429 39247 43463
rect 39613 43429 39647 43463
rect 40013 43429 40047 43463
rect 40413 43429 40447 43463
rect 40813 43429 40847 43463
rect 41213 43429 41247 43463
rect 41613 43429 41647 43463
rect 42013 43429 42047 43463
rect 42413 43429 42447 43463
rect 37459 39869 37493 39903
rect 37859 39869 37893 39903
rect 38259 39869 38293 39903
rect 38659 39869 38693 39903
rect 39059 39869 39093 39903
rect 39459 39869 39493 39903
rect 39859 39869 39893 39903
rect 40259 39869 40293 39903
rect 40659 39869 40693 39903
rect 41059 39869 41093 39903
rect 22857 39669 22891 39703
rect 23257 39669 23291 39703
rect 23657 39669 23691 39703
rect 24057 39669 24091 39703
rect 24457 39669 24491 39703
rect 24857 39669 24891 39703
rect 25257 39669 25291 39703
rect 25657 39669 25691 39703
rect 26057 39669 26091 39703
rect 26457 39669 26491 39703
rect 26857 39669 26891 39703
rect 27257 39669 27291 39703
rect 27657 39669 27691 39703
rect 28057 39669 28091 39703
rect 29521 39669 29555 39703
rect 29921 39669 29955 39703
rect 30321 39669 30355 39703
rect 30721 39669 30755 39703
rect 31121 39669 31155 39703
rect 31521 39669 31555 39703
rect 31921 39669 31955 39703
rect 32321 39669 32355 39703
rect 32721 39669 32755 39703
rect 33121 39669 33155 39703
rect 33521 39669 33555 39703
rect 33921 39669 33955 39703
rect 34321 39669 34355 39703
rect 34721 39669 34755 39703
rect 25601 36109 25635 36143
rect 26001 36109 26035 36143
rect 26401 36109 26435 36143
rect 26801 36109 26835 36143
rect 27201 36109 27235 36143
rect 27601 36109 27635 36143
rect 28001 36109 28035 36143
rect 28401 36109 28435 36143
rect 28801 36109 28835 36143
rect 29201 36109 29235 36143
rect 37655 35909 37689 35943
rect 38055 35909 38089 35943
rect 38455 35909 38489 35943
rect 38855 35909 38889 35943
rect 39255 35909 39289 35943
rect 39655 35909 39689 35943
rect 40055 35909 40089 35943
rect 37655 28389 37689 28423
rect 38055 28389 38089 28423
rect 38455 28389 38489 28423
rect 38855 28389 38889 28423
rect 39255 28389 39289 28423
rect 39655 28389 39689 28423
rect 40055 28389 40089 28423
rect 25601 24829 25635 24863
rect 26001 24829 26035 24863
rect 26401 24829 26435 24863
rect 26801 24829 26835 24863
rect 27201 24829 27235 24863
rect 27601 24829 27635 24863
rect 28001 24829 28035 24863
rect 28401 24829 28435 24863
rect 28801 24829 28835 24863
rect 29201 24829 29235 24863
rect 25013 17109 25047 17143
rect 25413 17109 25447 17143
rect 25813 17109 25847 17143
rect 26213 17109 26247 17143
rect 26613 17109 26647 17143
rect 27013 17109 27047 17143
rect 27413 17109 27447 17143
rect 27813 17109 27847 17143
rect 28213 17109 28247 17143
rect 28613 17109 28647 17143
rect 29013 17109 29047 17143
rect 29413 17109 29447 17143
rect 29813 17109 29847 17143
rect 30213 17109 30247 17143
rect 30613 17109 30647 17143
rect 31013 17109 31047 17143
rect 31413 17109 31447 17143
rect 31813 17109 31847 17143
rect 32213 17109 32247 17143
rect 32613 17109 32647 17143
rect 33013 17109 33047 17143
rect 33413 17109 33447 17143
rect 33813 17109 33847 17143
rect 34213 17109 34247 17143
rect 34613 17109 34647 17143
rect 35013 17109 35047 17143
rect 35413 17109 35447 17143
rect 35813 17109 35847 17143
rect 36213 17109 36247 17143
rect 36613 17109 36647 17143
rect 37013 17109 37047 17143
rect 37413 17109 37447 17143
rect 37813 17109 37847 17143
rect 38213 17109 38247 17143
rect 38613 17109 38647 17143
rect 39013 17109 39047 17143
rect 39413 17109 39447 17143
rect 39813 17109 39847 17143
rect 40213 17109 40247 17143
rect 40613 17109 40647 17143
rect 41013 17109 41047 17143
rect 41413 17109 41447 17143
rect 41813 17109 41847 17143
rect 42213 17109 42247 17143
rect 42613 17109 42647 17143
rect 43013 17109 43047 17143
rect 43413 17109 43447 17143
rect 43813 17109 43847 17143
rect 44213 17109 44247 17143
rect 44613 17109 44647 17143
rect 45013 17109 45047 17143
rect 45413 17109 45447 17143
rect 45813 17109 45847 17143
rect 46213 17109 46247 17143
rect 46613 17109 46647 17143
rect 47013 17109 47047 17143
rect 47413 17109 47447 17143
rect 47813 17109 47847 17143
rect 48213 17109 48247 17143
rect 48613 17109 48647 17143
rect 49013 17109 49047 17143
rect 49413 17109 49447 17143
rect 49813 17109 49847 17143
rect 50213 17109 50247 17143
rect 50613 17109 50647 17143
rect 51013 17109 51047 17143
rect 51413 17109 51447 17143
rect 51813 17109 51847 17143
rect 52213 17109 52247 17143
<< xpolycontact >>
rect 20832 48147 21264 48717
rect 22840 48147 23272 48717
rect 20832 47187 21264 47757
rect 22840 47187 23272 47757
rect 13678 36867 14110 37437
rect 15686 36867 16118 37437
rect 16422 36867 16854 37437
rect 18430 36867 18862 37437
rect 19167 36867 19599 37437
rect 21749 36867 22181 37437
rect 22498 36867 22930 37437
rect 24506 36867 24938 37437
rect 13678 35907 14110 36477
rect 15686 35907 16118 36477
rect 16422 35907 16854 36477
rect 18430 35907 18862 36477
rect 19167 35907 19599 36477
rect 21749 35907 22181 36477
rect 22498 35907 22930 36477
rect 24506 35907 24938 36477
rect 19264 33107 19696 33677
rect 21272 33107 21704 33677
rect 22009 33107 22441 33677
rect 24591 33107 25023 33677
rect 19264 32147 19696 32717
rect 21272 32147 21704 32717
rect 22009 32147 22441 32717
rect 24591 32147 25023 32717
rect 16520 29347 16952 29917
rect 18528 29347 18960 29917
rect 19264 29347 19696 29917
rect 21272 29347 21704 29917
rect 22008 29347 22440 29917
rect 24016 29347 24448 29917
rect 27202 29347 27634 29917
rect 29210 29347 29642 29917
rect 16520 28387 16952 28957
rect 18528 28387 18960 28957
rect 19264 28387 19696 28957
rect 21272 28387 21704 28957
rect 22008 28387 22440 28957
rect 24016 28387 24448 28957
rect 27202 28387 27634 28957
rect 29210 28387 29642 28957
rect 22400 25587 22832 26157
rect 24408 25587 24840 26157
rect 22400 24627 22832 25197
rect 24408 24627 24840 25197
rect 37394 25587 37826 26157
rect 39402 25587 39834 26157
rect 40138 25587 40570 26157
rect 42146 25587 42578 26157
rect 42882 25587 43314 26157
rect 44890 25587 45322 26157
rect 45626 25587 46058 26157
rect 47634 25587 48066 26157
rect 48370 25587 48802 26157
rect 50378 25587 50810 26157
rect 37394 24627 37826 25197
rect 39402 24627 39834 25197
rect 40138 24627 40570 25197
rect 42146 24627 42578 25197
rect 42882 24627 43314 25197
rect 44890 24627 45322 25197
rect 45626 24627 46058 25197
rect 47634 24627 48066 25197
rect 48370 24627 48802 25197
rect 50378 24627 50810 25197
rect 23870 21827 24302 22397
rect 25878 21827 26310 22397
rect 27202 21827 27634 22397
rect 29210 21827 29642 22397
rect 29946 21827 30378 22397
rect 31954 21827 32386 22397
rect 33180 21827 33612 22397
rect 35188 21827 35620 22397
rect 37394 21827 37826 22397
rect 39402 21827 39834 22397
rect 40138 21827 40570 22397
rect 42146 21827 42578 22397
rect 48370 21827 48802 22397
rect 50378 21827 50810 22397
rect 23870 20867 24302 21437
rect 25878 20867 26310 21437
rect 27202 20867 27634 21437
rect 29210 20867 29642 21437
rect 29946 20867 30378 21437
rect 31954 20867 32386 21437
rect 33180 20867 33612 21437
rect 35188 20867 35620 21437
rect 37394 20867 37826 21437
rect 39402 20867 39834 21437
rect 40138 20867 40570 21437
rect 42146 20867 42578 21437
rect 48370 20867 48802 21437
rect 50378 20867 50810 21437
rect 43862 14307 44294 14877
rect 45870 14307 46302 14877
rect 46606 14307 47038 14877
rect 48614 14307 49046 14877
rect 49350 14307 49782 14877
rect 51358 14307 51790 14877
rect 43862 13347 44294 13917
rect 45870 13347 46302 13917
rect 46606 13347 47038 13917
rect 48614 13347 49046 13917
rect 49350 13347 49782 13917
rect 51358 13347 51790 13917
rect 43764 10547 44196 11117
rect 45772 10547 46204 11117
rect 46508 10547 46940 11117
rect 48516 10547 48948 11117
rect 49252 10547 49684 11117
rect 51260 10547 51692 11117
rect 43764 9587 44196 10157
rect 45772 9587 46204 10157
rect 46508 9587 46940 10157
rect 48516 9587 48948 10157
rect 49252 9587 49684 10157
rect 51260 9587 51692 10157
rect 44548 6787 44980 7357
rect 46556 6787 46988 7357
rect 47292 6787 47724 7357
rect 49300 6787 49732 7357
rect 50036 6787 50468 7357
rect 52044 6787 52476 7357
rect 44548 5827 44980 6397
rect 46556 5827 46988 6397
rect 47292 5827 47724 6397
rect 49300 5827 49732 6397
rect 50036 5827 50468 6397
rect 52044 5827 52476 6397
<< xpolyres >>
rect 21264 48147 22840 48717
rect 21264 47187 22840 47757
rect 14110 36867 15686 37437
rect 16854 36867 18430 37437
rect 19599 36867 21749 37437
rect 22930 36867 24506 37437
rect 14110 35907 15686 36477
rect 16854 35907 18430 36477
rect 19599 35907 21749 36477
rect 22930 35907 24506 36477
rect 19696 33107 21272 33677
rect 22441 33107 24591 33677
rect 19696 32147 21272 32717
rect 22441 32147 24591 32717
rect 16952 29347 18528 29917
rect 19696 29347 21272 29917
rect 22440 29347 24016 29917
rect 27634 29347 29210 29917
rect 16952 28387 18528 28957
rect 19696 28387 21272 28957
rect 22440 28387 24016 28957
rect 27634 28387 29210 28957
rect 22832 25587 24408 26157
rect 22832 24627 24408 25197
rect 37826 25587 39402 26157
rect 40570 25587 42146 26157
rect 43314 25587 44890 26157
rect 46058 25587 47634 26157
rect 48802 25587 50378 26157
rect 37826 24627 39402 25197
rect 40570 24627 42146 25197
rect 43314 24627 44890 25197
rect 46058 24627 47634 25197
rect 48802 24627 50378 25197
rect 24302 21827 25878 22397
rect 27634 21827 29210 22397
rect 30378 21827 31954 22397
rect 33612 21827 35188 22397
rect 37826 21827 39402 22397
rect 40570 21827 42146 22397
rect 48802 21827 50378 22397
rect 24302 20867 25878 21437
rect 27634 20867 29210 21437
rect 30378 20867 31954 21437
rect 33612 20867 35188 21437
rect 37826 20867 39402 21437
rect 40570 20867 42146 21437
rect 48802 20867 50378 21437
rect 44294 14307 45870 14877
rect 47038 14307 48614 14877
rect 49782 14307 51358 14877
rect 44294 13347 45870 13917
rect 47038 13347 48614 13917
rect 49782 13347 51358 13917
rect 44196 10547 45772 11117
rect 46940 10547 48516 11117
rect 49684 10547 51260 11117
rect 44196 9587 45772 10157
rect 46940 9587 48516 10157
rect 49684 9587 51260 10157
rect 44980 6787 46556 7357
rect 47724 6787 49300 7357
rect 50468 6787 52044 7357
rect 44980 5827 46556 6397
rect 47724 5827 49300 6397
rect 50468 5827 52044 6397
<< locali >>
rect 5918 48969 13086 48982
rect 5918 48935 6101 48969
rect 6135 48935 6501 48969
rect 6535 48935 6901 48969
rect 6935 48935 7301 48969
rect 7335 48935 7701 48969
rect 7735 48935 8101 48969
rect 8135 48935 8501 48969
rect 8535 48935 8901 48969
rect 8935 48935 9301 48969
rect 9335 48935 9701 48969
rect 9735 48935 10101 48969
rect 10135 48935 10501 48969
rect 10535 48935 10901 48969
rect 10935 48935 11301 48969
rect 11335 48935 11701 48969
rect 11735 48935 12101 48969
rect 12135 48935 12501 48969
rect 12535 48935 12901 48969
rect 12935 48935 13086 48969
rect 5918 48922 13086 48935
rect 13366 48969 20534 48982
rect 13366 48935 13549 48969
rect 13583 48935 13949 48969
rect 13983 48935 14349 48969
rect 14383 48935 14749 48969
rect 14783 48935 15149 48969
rect 15183 48935 15549 48969
rect 15583 48935 15949 48969
rect 15983 48935 16349 48969
rect 16383 48935 16749 48969
rect 16783 48935 17149 48969
rect 17183 48935 17549 48969
rect 17583 48935 17949 48969
rect 17983 48935 18349 48969
rect 18383 48935 18749 48969
rect 18783 48935 19149 48969
rect 19183 48935 19549 48969
rect 19583 48935 19949 48969
rect 19983 48935 20349 48969
rect 20383 48935 20534 48969
rect 13366 48922 20534 48935
rect 20832 48969 23272 48982
rect 20832 48935 21015 48969
rect 21049 48935 21215 48969
rect 21249 48935 21415 48969
rect 21449 48935 21615 48969
rect 21649 48935 21815 48969
rect 21849 48935 22015 48969
rect 22049 48935 22215 48969
rect 22249 48935 22415 48969
rect 22449 48935 22615 48969
rect 22649 48935 22815 48969
rect 22849 48935 23015 48969
rect 23049 48935 23272 48969
rect 20832 48922 23272 48935
rect 23820 48969 24434 48982
rect 23820 48935 24101 48969
rect 24135 48935 24434 48969
rect 23820 48922 24434 48935
rect 24732 48969 52438 48982
rect 24732 48935 25013 48969
rect 25047 48935 25413 48969
rect 25447 48935 25813 48969
rect 25847 48935 26213 48969
rect 26247 48935 26613 48969
rect 26647 48935 27013 48969
rect 27047 48935 27413 48969
rect 27447 48935 27813 48969
rect 27847 48935 28213 48969
rect 28247 48935 28613 48969
rect 28647 48935 29013 48969
rect 29047 48935 29413 48969
rect 29447 48935 29813 48969
rect 29847 48935 30213 48969
rect 30247 48935 30613 48969
rect 30647 48935 31013 48969
rect 31047 48935 31413 48969
rect 31447 48935 31813 48969
rect 31847 48935 32213 48969
rect 32247 48935 32613 48969
rect 32647 48935 33013 48969
rect 33047 48935 33413 48969
rect 33447 48935 33813 48969
rect 33847 48935 34213 48969
rect 34247 48935 34613 48969
rect 34647 48935 35013 48969
rect 35047 48935 35413 48969
rect 35447 48935 35813 48969
rect 35847 48935 36213 48969
rect 36247 48935 36613 48969
rect 36647 48935 37013 48969
rect 37047 48935 37413 48969
rect 37447 48935 37813 48969
rect 37847 48935 38213 48969
rect 38247 48935 38613 48969
rect 38647 48935 39013 48969
rect 39047 48935 39413 48969
rect 39447 48935 39813 48969
rect 39847 48935 40213 48969
rect 40247 48935 40613 48969
rect 40647 48935 41013 48969
rect 41047 48935 41413 48969
rect 41447 48935 41813 48969
rect 41847 48935 42213 48969
rect 42247 48935 42613 48969
rect 42647 48935 43013 48969
rect 43047 48935 43413 48969
rect 43447 48935 43813 48969
rect 43847 48935 44213 48969
rect 44247 48935 44613 48969
rect 44647 48935 45013 48969
rect 45047 48935 45413 48969
rect 45447 48935 45813 48969
rect 45847 48935 46213 48969
rect 46247 48935 46613 48969
rect 46647 48935 47013 48969
rect 47047 48935 47413 48969
rect 47447 48935 47813 48969
rect 47847 48935 48213 48969
rect 48247 48935 48613 48969
rect 48647 48935 49013 48969
rect 49047 48935 49413 48969
rect 49447 48935 49813 48969
rect 49847 48935 50213 48969
rect 50247 48935 50613 48969
rect 50647 48935 51013 48969
rect 51047 48935 51413 48969
rect 51447 48935 51813 48969
rect 51847 48935 52213 48969
rect 52247 48935 52438 48969
rect 24732 48922 52438 48935
rect 24760 48829 24820 48922
rect 25808 48879 25968 48922
rect 25808 48845 25873 48879
rect 25907 48845 25968 48879
rect 25808 48842 25968 48845
rect 27108 48879 27268 48922
rect 27108 48845 27173 48879
rect 27207 48845 27268 48879
rect 27108 48842 27268 48845
rect 28408 48879 28568 48922
rect 28408 48845 28473 48879
rect 28507 48845 28568 48879
rect 28408 48842 28568 48845
rect 29708 48879 29868 48922
rect 29708 48845 29773 48879
rect 29807 48845 29868 48879
rect 29708 48842 29868 48845
rect 31008 48879 31168 48922
rect 31008 48845 31073 48879
rect 31107 48845 31168 48879
rect 31008 48842 31168 48845
rect 32308 48879 32468 48922
rect 32308 48845 32373 48879
rect 32407 48845 32468 48879
rect 32308 48842 32468 48845
rect 33608 48879 33768 48922
rect 33608 48845 33673 48879
rect 33707 48845 33768 48879
rect 33608 48842 33768 48845
rect 34908 48879 35068 48922
rect 34908 48845 34973 48879
rect 35007 48845 35068 48879
rect 34908 48842 35068 48845
rect 36208 48879 36368 48922
rect 36208 48845 36273 48879
rect 36307 48845 36368 48879
rect 36208 48842 36368 48845
rect 37508 48879 37668 48922
rect 37508 48845 37573 48879
rect 37607 48845 37668 48879
rect 37508 48842 37668 48845
rect 38808 48879 38968 48922
rect 38808 48845 38873 48879
rect 38907 48845 38968 48879
rect 38808 48842 38968 48845
rect 40108 48879 40268 48922
rect 40108 48845 40173 48879
rect 40207 48845 40268 48879
rect 40108 48842 40268 48845
rect 41408 48879 41568 48922
rect 41408 48845 41473 48879
rect 41507 48845 41568 48879
rect 41408 48842 41568 48845
rect 42708 48879 42868 48922
rect 42708 48845 42773 48879
rect 42807 48845 42868 48879
rect 42708 48842 42868 48845
rect 44008 48879 44168 48922
rect 44008 48845 44073 48879
rect 44107 48845 44168 48879
rect 44008 48842 44168 48845
rect 45308 48879 45468 48922
rect 45308 48845 45373 48879
rect 45407 48845 45468 48879
rect 45308 48842 45468 48845
rect 46608 48879 46768 48922
rect 46608 48845 46673 48879
rect 46707 48845 46768 48879
rect 46608 48842 46768 48845
rect 47908 48879 48068 48922
rect 47908 48845 47973 48879
rect 48007 48845 48068 48879
rect 47908 48842 48068 48845
rect 49208 48879 49368 48922
rect 49208 48845 49273 48879
rect 49307 48845 49368 48879
rect 49208 48842 49368 48845
rect 50508 48879 50668 48922
rect 50508 48845 50573 48879
rect 50607 48845 50668 48879
rect 50508 48842 50668 48845
rect 23918 48762 24434 48822
rect 24760 48795 24773 48829
rect 24807 48795 24820 48829
rect 24387 48476 24421 48762
rect 24760 48712 24820 48795
rect 24890 48762 52438 48802
rect 24877 48701 24911 48721
rect 24877 48633 24911 48667
rect 24877 48565 24911 48595
rect 24877 48497 24911 48523
rect 21744 48003 22360 48042
rect 21744 47901 21831 48003
rect 22273 47901 22360 48003
rect 21744 47102 22360 47901
rect 22840 47757 23272 48147
rect 23930 48449 23964 48476
rect 24387 48458 24422 48476
rect 23930 48377 23964 48395
rect 23930 48305 23964 48327
rect 23930 48233 23964 48259
rect 23930 48161 23964 48191
rect 23930 48089 23964 48123
rect 23930 48021 23964 48055
rect 23930 47953 23964 47983
rect 23930 47885 23964 47911
rect 23930 47817 23964 47839
rect 23930 47749 23964 47767
rect 23929 47695 23930 47726
rect 23929 47668 23964 47695
rect 24388 48449 24422 48458
rect 24388 48377 24422 48395
rect 24388 48305 24422 48327
rect 24388 48233 24422 48259
rect 24388 48161 24422 48191
rect 24388 48089 24422 48123
rect 24388 48021 24422 48055
rect 24388 47953 24422 47983
rect 24388 47885 24422 47911
rect 24388 47817 24422 47839
rect 24388 47749 24422 47767
rect 24388 47668 24422 47695
rect 24877 48429 24911 48451
rect 24877 48361 24911 48379
rect 24877 48293 24911 48307
rect 24877 48225 24911 48235
rect 24877 48157 24911 48163
rect 24877 48089 24911 48091
rect 24877 48053 24911 48055
rect 24877 47981 24911 47987
rect 24877 47909 24911 47919
rect 24877 47837 24911 47851
rect 24877 47765 24911 47783
rect 24877 47693 24911 47715
rect 23929 47502 23963 47668
rect 24877 47621 24911 47647
rect 24877 47549 24911 47579
rect 23918 47442 24434 47502
rect 24877 47477 24911 47511
rect 24877 47342 24911 47443
rect 25335 48701 25369 48762
rect 25335 48633 25369 48667
rect 25335 48565 25369 48595
rect 25335 48497 25369 48523
rect 25335 48429 25369 48451
rect 25335 48361 25369 48379
rect 25335 48293 25369 48307
rect 25335 48225 25369 48235
rect 25335 48157 25369 48163
rect 25335 48089 25369 48091
rect 25335 48053 25369 48055
rect 25335 47981 25369 47987
rect 25335 47909 25369 47919
rect 25335 47837 25369 47851
rect 25335 47765 25369 47783
rect 25335 47693 25369 47715
rect 25335 47621 25369 47647
rect 25335 47549 25369 47579
rect 25335 47477 25369 47511
rect 25335 47423 25369 47443
rect 25793 48701 25827 48721
rect 25793 48633 25827 48667
rect 25793 48565 25827 48595
rect 25793 48497 25827 48523
rect 25793 48429 25827 48451
rect 25793 48361 25827 48379
rect 25793 48293 25827 48307
rect 25793 48225 25827 48235
rect 25793 48157 25827 48163
rect 25793 48089 25827 48091
rect 25793 48053 25827 48055
rect 25793 47981 25827 47987
rect 25793 47909 25827 47919
rect 25793 47837 25827 47851
rect 25793 47765 25827 47783
rect 25793 47693 25827 47715
rect 25793 47621 25827 47647
rect 25793 47549 25827 47579
rect 25793 47477 25827 47511
rect 25793 47342 25827 47443
rect 26251 48701 26285 48762
rect 26251 48633 26285 48667
rect 26251 48565 26285 48595
rect 26251 48497 26285 48523
rect 26251 48429 26285 48451
rect 26251 48361 26285 48379
rect 26251 48293 26285 48307
rect 26251 48225 26285 48235
rect 26251 48157 26285 48163
rect 26251 48089 26285 48091
rect 26251 48053 26285 48055
rect 26251 47981 26285 47987
rect 26251 47909 26285 47919
rect 26251 47837 26285 47851
rect 26251 47765 26285 47783
rect 26251 47693 26285 47715
rect 26251 47621 26285 47647
rect 26251 47549 26285 47579
rect 26251 47477 26285 47511
rect 26251 47423 26285 47443
rect 26709 48701 26743 48721
rect 26709 48633 26743 48667
rect 26709 48565 26743 48595
rect 26709 48497 26743 48523
rect 26709 48429 26743 48451
rect 26709 48361 26743 48379
rect 26709 48293 26743 48307
rect 26709 48225 26743 48235
rect 26709 48157 26743 48163
rect 26709 48089 26743 48091
rect 26709 48053 26743 48055
rect 26709 47981 26743 47987
rect 26709 47909 26743 47919
rect 26709 47837 26743 47851
rect 26709 47765 26743 47783
rect 26709 47693 26743 47715
rect 26709 47621 26743 47647
rect 26709 47549 26743 47579
rect 26709 47477 26743 47511
rect 26709 47342 26743 47443
rect 27167 48701 27201 48762
rect 27167 48633 27201 48667
rect 27167 48565 27201 48595
rect 27167 48497 27201 48523
rect 27167 48429 27201 48451
rect 27167 48361 27201 48379
rect 27167 48293 27201 48307
rect 27167 48225 27201 48235
rect 27167 48157 27201 48163
rect 27167 48089 27201 48091
rect 27167 48053 27201 48055
rect 27167 47981 27201 47987
rect 27167 47909 27201 47919
rect 27167 47837 27201 47851
rect 27167 47765 27201 47783
rect 27167 47693 27201 47715
rect 27167 47621 27201 47647
rect 27167 47549 27201 47579
rect 27167 47477 27201 47511
rect 27167 47423 27201 47443
rect 27625 48701 27659 48721
rect 27625 48633 27659 48667
rect 27625 48565 27659 48595
rect 27625 48497 27659 48523
rect 27625 48429 27659 48451
rect 27625 48361 27659 48379
rect 27625 48293 27659 48307
rect 27625 48225 27659 48235
rect 27625 48157 27659 48163
rect 27625 48089 27659 48091
rect 27625 48053 27659 48055
rect 27625 47981 27659 47987
rect 27625 47909 27659 47919
rect 27625 47837 27659 47851
rect 27625 47765 27659 47783
rect 27625 47693 27659 47715
rect 27625 47621 27659 47647
rect 27625 47549 27659 47579
rect 27625 47477 27659 47511
rect 27625 47342 27659 47443
rect 28083 48701 28117 48762
rect 28083 48633 28117 48667
rect 28083 48565 28117 48595
rect 28083 48497 28117 48523
rect 28083 48429 28117 48451
rect 28083 48361 28117 48379
rect 28083 48293 28117 48307
rect 28083 48225 28117 48235
rect 28083 48157 28117 48163
rect 28083 48089 28117 48091
rect 28083 48053 28117 48055
rect 28083 47981 28117 47987
rect 28083 47909 28117 47919
rect 28083 47837 28117 47851
rect 28083 47765 28117 47783
rect 28083 47693 28117 47715
rect 28083 47621 28117 47647
rect 28083 47549 28117 47579
rect 28083 47477 28117 47511
rect 28083 47423 28117 47443
rect 28541 48701 28575 48721
rect 28541 48633 28575 48667
rect 28541 48565 28575 48595
rect 28541 48497 28575 48523
rect 28541 48429 28575 48451
rect 28541 48361 28575 48379
rect 28541 48293 28575 48307
rect 28541 48225 28575 48235
rect 28541 48157 28575 48163
rect 28541 48089 28575 48091
rect 28541 48053 28575 48055
rect 28541 47981 28575 47987
rect 28541 47909 28575 47919
rect 28541 47837 28575 47851
rect 28541 47765 28575 47783
rect 28541 47693 28575 47715
rect 28541 47621 28575 47647
rect 28541 47549 28575 47579
rect 28541 47477 28575 47511
rect 28541 47342 28575 47443
rect 28999 48701 29033 48762
rect 28999 48633 29033 48667
rect 28999 48565 29033 48595
rect 28999 48497 29033 48523
rect 28999 48429 29033 48451
rect 28999 48361 29033 48379
rect 28999 48293 29033 48307
rect 28999 48225 29033 48235
rect 28999 48157 29033 48163
rect 28999 48089 29033 48091
rect 28999 48053 29033 48055
rect 28999 47981 29033 47987
rect 28999 47909 29033 47919
rect 28999 47837 29033 47851
rect 28999 47765 29033 47783
rect 28999 47693 29033 47715
rect 28999 47621 29033 47647
rect 28999 47549 29033 47579
rect 28999 47477 29033 47511
rect 28999 47423 29033 47443
rect 29457 48701 29491 48721
rect 29457 48633 29491 48667
rect 29457 48565 29491 48595
rect 29457 48497 29491 48523
rect 29457 48429 29491 48451
rect 29457 48361 29491 48379
rect 29457 48293 29491 48307
rect 29457 48225 29491 48235
rect 29457 48157 29491 48163
rect 29457 48089 29491 48091
rect 29457 48053 29491 48055
rect 29457 47981 29491 47987
rect 29457 47909 29491 47919
rect 29457 47837 29491 47851
rect 29457 47765 29491 47783
rect 29457 47693 29491 47715
rect 29457 47621 29491 47647
rect 29457 47549 29491 47579
rect 29457 47477 29491 47511
rect 29457 47342 29491 47443
rect 29915 48701 29949 48762
rect 29915 48633 29949 48667
rect 29915 48565 29949 48595
rect 29915 48497 29949 48523
rect 29915 48429 29949 48451
rect 29915 48361 29949 48379
rect 29915 48293 29949 48307
rect 29915 48225 29949 48235
rect 29915 48157 29949 48163
rect 29915 48089 29949 48091
rect 29915 48053 29949 48055
rect 29915 47981 29949 47987
rect 29915 47909 29949 47919
rect 29915 47837 29949 47851
rect 29915 47765 29949 47783
rect 29915 47693 29949 47715
rect 29915 47621 29949 47647
rect 29915 47549 29949 47579
rect 29915 47477 29949 47511
rect 29915 47423 29949 47443
rect 30373 48701 30407 48721
rect 30373 48633 30407 48667
rect 30373 48565 30407 48595
rect 30373 48497 30407 48523
rect 30373 48429 30407 48451
rect 30373 48361 30407 48379
rect 30373 48293 30407 48307
rect 30373 48225 30407 48235
rect 30373 48157 30407 48163
rect 30373 48089 30407 48091
rect 30373 48053 30407 48055
rect 30373 47981 30407 47987
rect 30373 47909 30407 47919
rect 30373 47837 30407 47851
rect 30373 47765 30407 47783
rect 30373 47693 30407 47715
rect 30373 47621 30407 47647
rect 30373 47549 30407 47579
rect 30373 47477 30407 47511
rect 30373 47342 30407 47443
rect 30831 48701 30865 48762
rect 30831 48633 30865 48667
rect 30831 48565 30865 48595
rect 30831 48497 30865 48523
rect 30831 48429 30865 48451
rect 30831 48361 30865 48379
rect 30831 48293 30865 48307
rect 30831 48225 30865 48235
rect 30831 48157 30865 48163
rect 30831 48089 30865 48091
rect 30831 48053 30865 48055
rect 30831 47981 30865 47987
rect 30831 47909 30865 47919
rect 30831 47837 30865 47851
rect 30831 47765 30865 47783
rect 30831 47693 30865 47715
rect 30831 47621 30865 47647
rect 30831 47549 30865 47579
rect 30831 47477 30865 47511
rect 30831 47423 30865 47443
rect 31289 48701 31323 48721
rect 31289 48633 31323 48667
rect 31289 48565 31323 48595
rect 31289 48497 31323 48523
rect 31289 48429 31323 48451
rect 31289 48361 31323 48379
rect 31289 48293 31323 48307
rect 31289 48225 31323 48235
rect 31289 48157 31323 48163
rect 31289 48089 31323 48091
rect 31289 48053 31323 48055
rect 31289 47981 31323 47987
rect 31289 47909 31323 47919
rect 31289 47837 31323 47851
rect 31289 47765 31323 47783
rect 31289 47693 31323 47715
rect 31289 47621 31323 47647
rect 31289 47549 31323 47579
rect 31289 47477 31323 47511
rect 31289 47342 31323 47443
rect 31747 48701 31781 48762
rect 31747 48633 31781 48667
rect 31747 48565 31781 48595
rect 31747 48497 31781 48523
rect 31747 48429 31781 48451
rect 31747 48361 31781 48379
rect 31747 48293 31781 48307
rect 31747 48225 31781 48235
rect 31747 48157 31781 48163
rect 31747 48089 31781 48091
rect 31747 48053 31781 48055
rect 31747 47981 31781 47987
rect 31747 47909 31781 47919
rect 31747 47837 31781 47851
rect 31747 47765 31781 47783
rect 31747 47693 31781 47715
rect 31747 47621 31781 47647
rect 31747 47549 31781 47579
rect 31747 47477 31781 47511
rect 31747 47423 31781 47443
rect 32205 48701 32239 48721
rect 32205 48633 32239 48667
rect 32205 48565 32239 48595
rect 32205 48497 32239 48523
rect 32205 48429 32239 48451
rect 32205 48361 32239 48379
rect 32205 48293 32239 48307
rect 32205 48225 32239 48235
rect 32205 48157 32239 48163
rect 32205 48089 32239 48091
rect 32205 48053 32239 48055
rect 32205 47981 32239 47987
rect 32205 47909 32239 47919
rect 32205 47837 32239 47851
rect 32205 47765 32239 47783
rect 32205 47693 32239 47715
rect 32205 47621 32239 47647
rect 32205 47549 32239 47579
rect 32205 47477 32239 47511
rect 32205 47342 32239 47443
rect 32663 48701 32697 48762
rect 32663 48633 32697 48667
rect 32663 48565 32697 48595
rect 32663 48497 32697 48523
rect 32663 48429 32697 48451
rect 32663 48361 32697 48379
rect 32663 48293 32697 48307
rect 32663 48225 32697 48235
rect 32663 48157 32697 48163
rect 32663 48089 32697 48091
rect 32663 48053 32697 48055
rect 32663 47981 32697 47987
rect 32663 47909 32697 47919
rect 32663 47837 32697 47851
rect 32663 47765 32697 47783
rect 32663 47693 32697 47715
rect 32663 47621 32697 47647
rect 32663 47549 32697 47579
rect 32663 47477 32697 47511
rect 32663 47423 32697 47443
rect 33121 48701 33155 48721
rect 33121 48633 33155 48667
rect 33121 48565 33155 48595
rect 33121 48497 33155 48523
rect 33121 48429 33155 48451
rect 33121 48361 33155 48379
rect 33121 48293 33155 48307
rect 33121 48225 33155 48235
rect 33121 48157 33155 48163
rect 33121 48089 33155 48091
rect 33121 48053 33155 48055
rect 33121 47981 33155 47987
rect 33121 47909 33155 47919
rect 33121 47837 33155 47851
rect 33121 47765 33155 47783
rect 33121 47693 33155 47715
rect 33121 47621 33155 47647
rect 33121 47549 33155 47579
rect 33121 47477 33155 47511
rect 33121 47342 33155 47443
rect 33579 48701 33613 48762
rect 33579 48633 33613 48667
rect 33579 48565 33613 48595
rect 33579 48497 33613 48523
rect 33579 48429 33613 48451
rect 33579 48361 33613 48379
rect 33579 48293 33613 48307
rect 33579 48225 33613 48235
rect 33579 48157 33613 48163
rect 33579 48089 33613 48091
rect 33579 48053 33613 48055
rect 33579 47981 33613 47987
rect 33579 47909 33613 47919
rect 33579 47837 33613 47851
rect 33579 47765 33613 47783
rect 33579 47693 33613 47715
rect 33579 47621 33613 47647
rect 33579 47549 33613 47579
rect 33579 47477 33613 47511
rect 33579 47423 33613 47443
rect 34037 48701 34071 48721
rect 34037 48633 34071 48667
rect 34037 48565 34071 48595
rect 34037 48497 34071 48523
rect 34037 48429 34071 48451
rect 34037 48361 34071 48379
rect 34037 48293 34071 48307
rect 34037 48225 34071 48235
rect 34037 48157 34071 48163
rect 34037 48089 34071 48091
rect 34037 48053 34071 48055
rect 34037 47981 34071 47987
rect 34037 47909 34071 47919
rect 34037 47837 34071 47851
rect 34037 47765 34071 47783
rect 34037 47693 34071 47715
rect 34037 47621 34071 47647
rect 34037 47549 34071 47579
rect 34037 47477 34071 47511
rect 34037 47342 34071 47443
rect 34495 48701 34529 48762
rect 34495 48633 34529 48667
rect 34495 48565 34529 48595
rect 34495 48497 34529 48523
rect 34495 48429 34529 48451
rect 34495 48361 34529 48379
rect 34495 48293 34529 48307
rect 34495 48225 34529 48235
rect 34495 48157 34529 48163
rect 34495 48089 34529 48091
rect 34495 48053 34529 48055
rect 34495 47981 34529 47987
rect 34495 47909 34529 47919
rect 34495 47837 34529 47851
rect 34495 47765 34529 47783
rect 34495 47693 34529 47715
rect 34495 47621 34529 47647
rect 34495 47549 34529 47579
rect 34495 47477 34529 47511
rect 34495 47423 34529 47443
rect 34953 48701 34987 48721
rect 34953 48633 34987 48667
rect 34953 48565 34987 48595
rect 34953 48497 34987 48523
rect 34953 48429 34987 48451
rect 34953 48361 34987 48379
rect 34953 48293 34987 48307
rect 34953 48225 34987 48235
rect 34953 48157 34987 48163
rect 34953 48089 34987 48091
rect 34953 48053 34987 48055
rect 34953 47981 34987 47987
rect 34953 47909 34987 47919
rect 34953 47837 34987 47851
rect 34953 47765 34987 47783
rect 34953 47693 34987 47715
rect 34953 47621 34987 47647
rect 34953 47549 34987 47579
rect 34953 47477 34987 47511
rect 34953 47342 34987 47443
rect 35411 48701 35445 48762
rect 35411 48633 35445 48667
rect 35411 48565 35445 48595
rect 35411 48497 35445 48523
rect 35411 48429 35445 48451
rect 35411 48361 35445 48379
rect 35411 48293 35445 48307
rect 35411 48225 35445 48235
rect 35411 48157 35445 48163
rect 35411 48089 35445 48091
rect 35411 48053 35445 48055
rect 35411 47981 35445 47987
rect 35411 47909 35445 47919
rect 35411 47837 35445 47851
rect 35411 47765 35445 47783
rect 35411 47693 35445 47715
rect 35411 47621 35445 47647
rect 35411 47549 35445 47579
rect 35411 47477 35445 47511
rect 35411 47423 35445 47443
rect 35869 48701 35903 48721
rect 35869 48633 35903 48667
rect 35869 48565 35903 48595
rect 35869 48497 35903 48523
rect 35869 48429 35903 48451
rect 35869 48361 35903 48379
rect 35869 48293 35903 48307
rect 35869 48225 35903 48235
rect 35869 48157 35903 48163
rect 35869 48089 35903 48091
rect 35869 48053 35903 48055
rect 35869 47981 35903 47987
rect 35869 47909 35903 47919
rect 35869 47837 35903 47851
rect 35869 47765 35903 47783
rect 35869 47693 35903 47715
rect 35869 47621 35903 47647
rect 35869 47549 35903 47579
rect 35869 47477 35903 47511
rect 35869 47342 35903 47443
rect 36327 48701 36361 48762
rect 36327 48633 36361 48667
rect 36327 48565 36361 48595
rect 36327 48497 36361 48523
rect 36327 48429 36361 48451
rect 36327 48361 36361 48379
rect 36327 48293 36361 48307
rect 36327 48225 36361 48235
rect 36327 48157 36361 48163
rect 36327 48089 36361 48091
rect 36327 48053 36361 48055
rect 36327 47981 36361 47987
rect 36327 47909 36361 47919
rect 36327 47837 36361 47851
rect 36327 47765 36361 47783
rect 36327 47693 36361 47715
rect 36327 47621 36361 47647
rect 36327 47549 36361 47579
rect 36327 47477 36361 47511
rect 36327 47423 36361 47443
rect 36785 48701 36819 48721
rect 36785 48633 36819 48667
rect 36785 48565 36819 48595
rect 36785 48497 36819 48523
rect 36785 48429 36819 48451
rect 36785 48361 36819 48379
rect 36785 48293 36819 48307
rect 36785 48225 36819 48235
rect 36785 48157 36819 48163
rect 36785 48089 36819 48091
rect 36785 48053 36819 48055
rect 36785 47981 36819 47987
rect 36785 47909 36819 47919
rect 36785 47837 36819 47851
rect 36785 47765 36819 47783
rect 36785 47693 36819 47715
rect 36785 47621 36819 47647
rect 36785 47549 36819 47579
rect 36785 47477 36819 47511
rect 36785 47342 36819 47443
rect 37243 48701 37277 48762
rect 37243 48633 37277 48667
rect 37243 48565 37277 48595
rect 37243 48497 37277 48523
rect 37243 48429 37277 48451
rect 37243 48361 37277 48379
rect 37243 48293 37277 48307
rect 37243 48225 37277 48235
rect 37243 48157 37277 48163
rect 37243 48089 37277 48091
rect 37243 48053 37277 48055
rect 37243 47981 37277 47987
rect 37243 47909 37277 47919
rect 37243 47837 37277 47851
rect 37243 47765 37277 47783
rect 37243 47693 37277 47715
rect 37243 47621 37277 47647
rect 37243 47549 37277 47579
rect 37243 47477 37277 47511
rect 37243 47423 37277 47443
rect 37701 48701 37735 48721
rect 37701 48633 37735 48667
rect 37701 48565 37735 48595
rect 37701 48497 37735 48523
rect 37701 48429 37735 48451
rect 37701 48361 37735 48379
rect 37701 48293 37735 48307
rect 37701 48225 37735 48235
rect 37701 48157 37735 48163
rect 37701 48089 37735 48091
rect 37701 48053 37735 48055
rect 37701 47981 37735 47987
rect 37701 47909 37735 47919
rect 37701 47837 37735 47851
rect 37701 47765 37735 47783
rect 37701 47693 37735 47715
rect 37701 47621 37735 47647
rect 37701 47549 37735 47579
rect 37701 47477 37735 47511
rect 37701 47342 37735 47443
rect 38159 48701 38193 48762
rect 38159 48633 38193 48667
rect 38159 48565 38193 48595
rect 38159 48497 38193 48523
rect 38159 48429 38193 48451
rect 38159 48361 38193 48379
rect 38159 48293 38193 48307
rect 38159 48225 38193 48235
rect 38159 48157 38193 48163
rect 38159 48089 38193 48091
rect 38159 48053 38193 48055
rect 38159 47981 38193 47987
rect 38159 47909 38193 47919
rect 38159 47837 38193 47851
rect 38159 47765 38193 47783
rect 38159 47693 38193 47715
rect 38159 47621 38193 47647
rect 38159 47549 38193 47579
rect 38159 47477 38193 47511
rect 38159 47423 38193 47443
rect 38617 48701 38651 48721
rect 38617 48633 38651 48667
rect 38617 48565 38651 48595
rect 38617 48497 38651 48523
rect 38617 48429 38651 48451
rect 38617 48361 38651 48379
rect 38617 48293 38651 48307
rect 38617 48225 38651 48235
rect 38617 48157 38651 48163
rect 38617 48089 38651 48091
rect 38617 48053 38651 48055
rect 38617 47981 38651 47987
rect 38617 47909 38651 47919
rect 38617 47837 38651 47851
rect 38617 47765 38651 47783
rect 38617 47693 38651 47715
rect 38617 47621 38651 47647
rect 38617 47549 38651 47579
rect 38617 47477 38651 47511
rect 38617 47342 38651 47443
rect 39075 48701 39109 48762
rect 39075 48633 39109 48667
rect 39075 48565 39109 48595
rect 39075 48497 39109 48523
rect 39075 48429 39109 48451
rect 39075 48361 39109 48379
rect 39075 48293 39109 48307
rect 39075 48225 39109 48235
rect 39075 48157 39109 48163
rect 39075 48089 39109 48091
rect 39075 48053 39109 48055
rect 39075 47981 39109 47987
rect 39075 47909 39109 47919
rect 39075 47837 39109 47851
rect 39075 47765 39109 47783
rect 39075 47693 39109 47715
rect 39075 47621 39109 47647
rect 39075 47549 39109 47579
rect 39075 47477 39109 47511
rect 39075 47423 39109 47443
rect 39533 48701 39567 48721
rect 39533 48633 39567 48667
rect 39533 48565 39567 48595
rect 39533 48497 39567 48523
rect 39533 48429 39567 48451
rect 39533 48361 39567 48379
rect 39533 48293 39567 48307
rect 39533 48225 39567 48235
rect 39533 48157 39567 48163
rect 39533 48089 39567 48091
rect 39533 48053 39567 48055
rect 39533 47981 39567 47987
rect 39533 47909 39567 47919
rect 39533 47837 39567 47851
rect 39533 47765 39567 47783
rect 39533 47693 39567 47715
rect 39533 47621 39567 47647
rect 39533 47549 39567 47579
rect 39533 47477 39567 47511
rect 39533 47342 39567 47443
rect 39991 48701 40025 48762
rect 39991 48633 40025 48667
rect 39991 48565 40025 48595
rect 39991 48497 40025 48523
rect 39991 48429 40025 48451
rect 39991 48361 40025 48379
rect 39991 48293 40025 48307
rect 39991 48225 40025 48235
rect 39991 48157 40025 48163
rect 39991 48089 40025 48091
rect 39991 48053 40025 48055
rect 39991 47981 40025 47987
rect 39991 47909 40025 47919
rect 39991 47837 40025 47851
rect 39991 47765 40025 47783
rect 39991 47693 40025 47715
rect 39991 47621 40025 47647
rect 39991 47549 40025 47579
rect 39991 47477 40025 47511
rect 39991 47423 40025 47443
rect 40449 48701 40483 48721
rect 40449 48633 40483 48667
rect 40449 48565 40483 48595
rect 40449 48497 40483 48523
rect 40449 48429 40483 48451
rect 40449 48361 40483 48379
rect 40449 48293 40483 48307
rect 40449 48225 40483 48235
rect 40449 48157 40483 48163
rect 40449 48089 40483 48091
rect 40449 48053 40483 48055
rect 40449 47981 40483 47987
rect 40449 47909 40483 47919
rect 40449 47837 40483 47851
rect 40449 47765 40483 47783
rect 40449 47693 40483 47715
rect 40449 47621 40483 47647
rect 40449 47549 40483 47579
rect 40449 47477 40483 47511
rect 40449 47342 40483 47443
rect 40907 48701 40941 48762
rect 40907 48633 40941 48667
rect 40907 48565 40941 48595
rect 40907 48497 40941 48523
rect 40907 48429 40941 48451
rect 40907 48361 40941 48379
rect 40907 48293 40941 48307
rect 40907 48225 40941 48235
rect 40907 48157 40941 48163
rect 40907 48089 40941 48091
rect 40907 48053 40941 48055
rect 40907 47981 40941 47987
rect 40907 47909 40941 47919
rect 40907 47837 40941 47851
rect 40907 47765 40941 47783
rect 40907 47693 40941 47715
rect 40907 47621 40941 47647
rect 40907 47549 40941 47579
rect 40907 47477 40941 47511
rect 40907 47423 40941 47443
rect 41365 48701 41399 48721
rect 41365 48633 41399 48667
rect 41365 48565 41399 48595
rect 41365 48497 41399 48523
rect 41365 48429 41399 48451
rect 41365 48361 41399 48379
rect 41365 48293 41399 48307
rect 41365 48225 41399 48235
rect 41365 48157 41399 48163
rect 41365 48089 41399 48091
rect 41365 48053 41399 48055
rect 41365 47981 41399 47987
rect 41365 47909 41399 47919
rect 41365 47837 41399 47851
rect 41365 47765 41399 47783
rect 41365 47693 41399 47715
rect 41365 47621 41399 47647
rect 41365 47549 41399 47579
rect 41365 47477 41399 47511
rect 41365 47342 41399 47443
rect 41823 48701 41857 48762
rect 41823 48633 41857 48667
rect 41823 48565 41857 48595
rect 41823 48497 41857 48523
rect 41823 48429 41857 48451
rect 41823 48361 41857 48379
rect 41823 48293 41857 48307
rect 41823 48225 41857 48235
rect 41823 48157 41857 48163
rect 41823 48089 41857 48091
rect 41823 48053 41857 48055
rect 41823 47981 41857 47987
rect 41823 47909 41857 47919
rect 41823 47837 41857 47851
rect 41823 47765 41857 47783
rect 41823 47693 41857 47715
rect 41823 47621 41857 47647
rect 41823 47549 41857 47579
rect 41823 47477 41857 47511
rect 41823 47423 41857 47443
rect 42281 48701 42315 48721
rect 42281 48633 42315 48667
rect 42281 48565 42315 48595
rect 42281 48497 42315 48523
rect 42281 48429 42315 48451
rect 42281 48361 42315 48379
rect 42281 48293 42315 48307
rect 42281 48225 42315 48235
rect 42281 48157 42315 48163
rect 42281 48089 42315 48091
rect 42281 48053 42315 48055
rect 42281 47981 42315 47987
rect 42281 47909 42315 47919
rect 42281 47837 42315 47851
rect 42281 47765 42315 47783
rect 42281 47693 42315 47715
rect 42281 47621 42315 47647
rect 42281 47549 42315 47579
rect 42281 47477 42315 47511
rect 42281 47342 42315 47443
rect 42739 48701 42773 48762
rect 42739 48633 42773 48667
rect 42739 48565 42773 48595
rect 42739 48497 42773 48523
rect 42739 48429 42773 48451
rect 42739 48361 42773 48379
rect 42739 48293 42773 48307
rect 42739 48225 42773 48235
rect 42739 48157 42773 48163
rect 42739 48089 42773 48091
rect 42739 48053 42773 48055
rect 42739 47981 42773 47987
rect 42739 47909 42773 47919
rect 42739 47837 42773 47851
rect 42739 47765 42773 47783
rect 42739 47693 42773 47715
rect 42739 47621 42773 47647
rect 42739 47549 42773 47579
rect 42739 47477 42773 47511
rect 42739 47423 42773 47443
rect 43197 48701 43231 48721
rect 43197 48633 43231 48667
rect 43197 48565 43231 48595
rect 43197 48497 43231 48523
rect 43197 48429 43231 48451
rect 43197 48361 43231 48379
rect 43197 48293 43231 48307
rect 43197 48225 43231 48235
rect 43197 48157 43231 48163
rect 43197 48089 43231 48091
rect 43197 48053 43231 48055
rect 43197 47981 43231 47987
rect 43197 47909 43231 47919
rect 43197 47837 43231 47851
rect 43197 47765 43231 47783
rect 43197 47693 43231 47715
rect 43197 47621 43231 47647
rect 43197 47549 43231 47579
rect 43197 47477 43231 47511
rect 43197 47342 43231 47443
rect 43655 48701 43689 48762
rect 43655 48633 43689 48667
rect 43655 48565 43689 48595
rect 43655 48497 43689 48523
rect 43655 48429 43689 48451
rect 43655 48361 43689 48379
rect 43655 48293 43689 48307
rect 43655 48225 43689 48235
rect 43655 48157 43689 48163
rect 43655 48089 43689 48091
rect 43655 48053 43689 48055
rect 43655 47981 43689 47987
rect 43655 47909 43689 47919
rect 43655 47837 43689 47851
rect 43655 47765 43689 47783
rect 43655 47693 43689 47715
rect 43655 47621 43689 47647
rect 43655 47549 43689 47579
rect 43655 47477 43689 47511
rect 43655 47423 43689 47443
rect 44113 48701 44147 48721
rect 44113 48633 44147 48667
rect 44113 48565 44147 48595
rect 44113 48497 44147 48523
rect 44113 48429 44147 48451
rect 44113 48361 44147 48379
rect 44113 48293 44147 48307
rect 44113 48225 44147 48235
rect 44113 48157 44147 48163
rect 44113 48089 44147 48091
rect 44113 48053 44147 48055
rect 44113 47981 44147 47987
rect 44113 47909 44147 47919
rect 44113 47837 44147 47851
rect 44113 47765 44147 47783
rect 44113 47693 44147 47715
rect 44113 47621 44147 47647
rect 44113 47549 44147 47579
rect 44113 47477 44147 47511
rect 44113 47342 44147 47443
rect 44571 48701 44605 48762
rect 44571 48633 44605 48667
rect 44571 48565 44605 48595
rect 44571 48497 44605 48523
rect 44571 48429 44605 48451
rect 44571 48361 44605 48379
rect 44571 48293 44605 48307
rect 44571 48225 44605 48235
rect 44571 48157 44605 48163
rect 44571 48089 44605 48091
rect 44571 48053 44605 48055
rect 44571 47981 44605 47987
rect 44571 47909 44605 47919
rect 44571 47837 44605 47851
rect 44571 47765 44605 47783
rect 44571 47693 44605 47715
rect 44571 47621 44605 47647
rect 44571 47549 44605 47579
rect 44571 47477 44605 47511
rect 44571 47423 44605 47443
rect 45029 48701 45063 48721
rect 45029 48633 45063 48667
rect 45029 48565 45063 48595
rect 45029 48497 45063 48523
rect 45029 48429 45063 48451
rect 45029 48361 45063 48379
rect 45029 48293 45063 48307
rect 45029 48225 45063 48235
rect 45029 48157 45063 48163
rect 45029 48089 45063 48091
rect 45029 48053 45063 48055
rect 45029 47981 45063 47987
rect 45029 47909 45063 47919
rect 45029 47837 45063 47851
rect 45029 47765 45063 47783
rect 45029 47693 45063 47715
rect 45029 47621 45063 47647
rect 45029 47549 45063 47579
rect 45029 47477 45063 47511
rect 45029 47342 45063 47443
rect 45487 48701 45521 48762
rect 45487 48633 45521 48667
rect 45487 48565 45521 48595
rect 45487 48497 45521 48523
rect 45487 48429 45521 48451
rect 45487 48361 45521 48379
rect 45487 48293 45521 48307
rect 45487 48225 45521 48235
rect 45487 48157 45521 48163
rect 45487 48089 45521 48091
rect 45487 48053 45521 48055
rect 45487 47981 45521 47987
rect 45487 47909 45521 47919
rect 45487 47837 45521 47851
rect 45487 47765 45521 47783
rect 45487 47693 45521 47715
rect 45487 47621 45521 47647
rect 45487 47549 45521 47579
rect 45487 47477 45521 47511
rect 45487 47423 45521 47443
rect 45945 48701 45979 48721
rect 45945 48633 45979 48667
rect 45945 48565 45979 48595
rect 45945 48497 45979 48523
rect 45945 48429 45979 48451
rect 45945 48361 45979 48379
rect 45945 48293 45979 48307
rect 45945 48225 45979 48235
rect 45945 48157 45979 48163
rect 45945 48089 45979 48091
rect 45945 48053 45979 48055
rect 45945 47981 45979 47987
rect 45945 47909 45979 47919
rect 45945 47837 45979 47851
rect 45945 47765 45979 47783
rect 45945 47693 45979 47715
rect 45945 47621 45979 47647
rect 45945 47549 45979 47579
rect 45945 47477 45979 47511
rect 45945 47342 45979 47443
rect 46403 48701 46437 48762
rect 46403 48633 46437 48667
rect 46403 48565 46437 48595
rect 46403 48497 46437 48523
rect 46403 48429 46437 48451
rect 46403 48361 46437 48379
rect 46403 48293 46437 48307
rect 46403 48225 46437 48235
rect 46403 48157 46437 48163
rect 46403 48089 46437 48091
rect 46403 48053 46437 48055
rect 46403 47981 46437 47987
rect 46403 47909 46437 47919
rect 46403 47837 46437 47851
rect 46403 47765 46437 47783
rect 46403 47693 46437 47715
rect 46403 47621 46437 47647
rect 46403 47549 46437 47579
rect 46403 47477 46437 47511
rect 46403 47423 46437 47443
rect 46861 48701 46895 48721
rect 46861 48633 46895 48667
rect 46861 48565 46895 48595
rect 46861 48497 46895 48523
rect 46861 48429 46895 48451
rect 46861 48361 46895 48379
rect 46861 48293 46895 48307
rect 46861 48225 46895 48235
rect 46861 48157 46895 48163
rect 46861 48089 46895 48091
rect 46861 48053 46895 48055
rect 46861 47981 46895 47987
rect 46861 47909 46895 47919
rect 46861 47837 46895 47851
rect 46861 47765 46895 47783
rect 46861 47693 46895 47715
rect 46861 47621 46895 47647
rect 46861 47549 46895 47579
rect 46861 47477 46895 47511
rect 46861 47342 46895 47443
rect 47319 48701 47353 48762
rect 47319 48633 47353 48667
rect 47319 48565 47353 48595
rect 47319 48497 47353 48523
rect 47319 48429 47353 48451
rect 47319 48361 47353 48379
rect 47319 48293 47353 48307
rect 47319 48225 47353 48235
rect 47319 48157 47353 48163
rect 47319 48089 47353 48091
rect 47319 48053 47353 48055
rect 47319 47981 47353 47987
rect 47319 47909 47353 47919
rect 47319 47837 47353 47851
rect 47319 47765 47353 47783
rect 47319 47693 47353 47715
rect 47319 47621 47353 47647
rect 47319 47549 47353 47579
rect 47319 47477 47353 47511
rect 47319 47423 47353 47443
rect 47777 48701 47811 48721
rect 47777 48633 47811 48667
rect 47777 48565 47811 48595
rect 47777 48497 47811 48523
rect 47777 48429 47811 48451
rect 47777 48361 47811 48379
rect 47777 48293 47811 48307
rect 47777 48225 47811 48235
rect 47777 48157 47811 48163
rect 47777 48089 47811 48091
rect 47777 48053 47811 48055
rect 47777 47981 47811 47987
rect 47777 47909 47811 47919
rect 47777 47837 47811 47851
rect 47777 47765 47811 47783
rect 47777 47693 47811 47715
rect 47777 47621 47811 47647
rect 47777 47549 47811 47579
rect 47777 47477 47811 47511
rect 47777 47342 47811 47443
rect 48235 48701 48269 48762
rect 48235 48633 48269 48667
rect 48235 48565 48269 48595
rect 48235 48497 48269 48523
rect 48235 48429 48269 48451
rect 48235 48361 48269 48379
rect 48235 48293 48269 48307
rect 48235 48225 48269 48235
rect 48235 48157 48269 48163
rect 48235 48089 48269 48091
rect 48235 48053 48269 48055
rect 48235 47981 48269 47987
rect 48235 47909 48269 47919
rect 48235 47837 48269 47851
rect 48235 47765 48269 47783
rect 48235 47693 48269 47715
rect 48235 47621 48269 47647
rect 48235 47549 48269 47579
rect 48235 47477 48269 47511
rect 48235 47423 48269 47443
rect 48693 48701 48727 48721
rect 48693 48633 48727 48667
rect 48693 48565 48727 48595
rect 48693 48497 48727 48523
rect 48693 48429 48727 48451
rect 48693 48361 48727 48379
rect 48693 48293 48727 48307
rect 48693 48225 48727 48235
rect 48693 48157 48727 48163
rect 48693 48089 48727 48091
rect 48693 48053 48727 48055
rect 48693 47981 48727 47987
rect 48693 47909 48727 47919
rect 48693 47837 48727 47851
rect 48693 47765 48727 47783
rect 48693 47693 48727 47715
rect 48693 47621 48727 47647
rect 48693 47549 48727 47579
rect 48693 47477 48727 47511
rect 48693 47342 48727 47443
rect 49151 48701 49185 48762
rect 49151 48633 49185 48667
rect 49151 48565 49185 48595
rect 49151 48497 49185 48523
rect 49151 48429 49185 48451
rect 49151 48361 49185 48379
rect 49151 48293 49185 48307
rect 49151 48225 49185 48235
rect 49151 48157 49185 48163
rect 49151 48089 49185 48091
rect 49151 48053 49185 48055
rect 49151 47981 49185 47987
rect 49151 47909 49185 47919
rect 49151 47837 49185 47851
rect 49151 47765 49185 47783
rect 49151 47693 49185 47715
rect 49151 47621 49185 47647
rect 49151 47549 49185 47579
rect 49151 47477 49185 47511
rect 49151 47423 49185 47443
rect 49609 48701 49643 48721
rect 49609 48633 49643 48667
rect 49609 48565 49643 48595
rect 49609 48497 49643 48523
rect 49609 48429 49643 48451
rect 49609 48361 49643 48379
rect 49609 48293 49643 48307
rect 49609 48225 49643 48235
rect 49609 48157 49643 48163
rect 49609 48089 49643 48091
rect 49609 48053 49643 48055
rect 49609 47981 49643 47987
rect 49609 47909 49643 47919
rect 49609 47837 49643 47851
rect 49609 47765 49643 47783
rect 49609 47693 49643 47715
rect 49609 47621 49643 47647
rect 49609 47549 49643 47579
rect 49609 47477 49643 47511
rect 49609 47342 49643 47443
rect 50067 48701 50101 48762
rect 50067 48633 50101 48667
rect 50067 48565 50101 48595
rect 50067 48497 50101 48523
rect 50067 48429 50101 48451
rect 50067 48361 50101 48379
rect 50067 48293 50101 48307
rect 50067 48225 50101 48235
rect 50067 48157 50101 48163
rect 50067 48089 50101 48091
rect 50067 48053 50101 48055
rect 50067 47981 50101 47987
rect 50067 47909 50101 47919
rect 50067 47837 50101 47851
rect 50067 47765 50101 47783
rect 50067 47693 50101 47715
rect 50067 47621 50101 47647
rect 50067 47549 50101 47579
rect 50067 47477 50101 47511
rect 50067 47423 50101 47443
rect 50525 48701 50559 48721
rect 50525 48633 50559 48667
rect 50525 48565 50559 48595
rect 50525 48497 50559 48523
rect 50525 48429 50559 48451
rect 50525 48361 50559 48379
rect 50525 48293 50559 48307
rect 50525 48225 50559 48235
rect 50525 48157 50559 48163
rect 50525 48089 50559 48091
rect 50525 48053 50559 48055
rect 50525 47981 50559 47987
rect 50525 47909 50559 47919
rect 50525 47837 50559 47851
rect 50525 47765 50559 47783
rect 50525 47693 50559 47715
rect 50525 47621 50559 47647
rect 50525 47549 50559 47579
rect 50525 47477 50559 47511
rect 50525 47342 50559 47443
rect 50983 48701 51017 48762
rect 50983 48633 51017 48667
rect 50983 48565 51017 48595
rect 50983 48497 51017 48523
rect 50983 48429 51017 48451
rect 50983 48361 51017 48379
rect 50983 48293 51017 48307
rect 50983 48225 51017 48235
rect 50983 48157 51017 48163
rect 50983 48089 51017 48091
rect 50983 48053 51017 48055
rect 50983 47981 51017 47987
rect 50983 47909 51017 47919
rect 50983 47837 51017 47851
rect 50983 47765 51017 47783
rect 50983 47693 51017 47715
rect 50983 47621 51017 47647
rect 50983 47549 51017 47579
rect 50983 47477 51017 47511
rect 50983 47423 51017 47443
rect 51441 48701 51475 48721
rect 51441 48633 51475 48667
rect 51441 48565 51475 48595
rect 51441 48497 51475 48523
rect 51441 48429 51475 48451
rect 51441 48361 51475 48379
rect 51441 48293 51475 48307
rect 51441 48225 51475 48235
rect 51441 48157 51475 48163
rect 51441 48089 51475 48091
rect 51441 48053 51475 48055
rect 51441 47981 51475 47987
rect 51441 47909 51475 47919
rect 51441 47837 51475 47851
rect 51441 47765 51475 47783
rect 51441 47693 51475 47715
rect 51441 47621 51475 47647
rect 51441 47549 51475 47579
rect 51441 47477 51475 47511
rect 51441 47342 51475 47443
rect 51899 48701 51933 48762
rect 51899 48633 51933 48667
rect 51899 48565 51933 48595
rect 51899 48497 51933 48523
rect 51899 48429 51933 48451
rect 51899 48361 51933 48379
rect 51899 48293 51933 48307
rect 51899 48225 51933 48235
rect 51899 48157 51933 48163
rect 51899 48089 51933 48091
rect 51899 48053 51933 48055
rect 51899 47981 51933 47987
rect 51899 47909 51933 47919
rect 51899 47837 51933 47851
rect 51899 47765 51933 47783
rect 51899 47693 51933 47715
rect 51899 47621 51933 47647
rect 51899 47549 51933 47579
rect 51899 47477 51933 47511
rect 51899 47423 51933 47443
rect 52357 48701 52391 48721
rect 52357 48633 52391 48667
rect 52357 48565 52391 48595
rect 52357 48497 52391 48523
rect 52357 48429 52391 48451
rect 52357 48361 52391 48379
rect 52357 48293 52391 48307
rect 52357 48225 52391 48235
rect 52357 48157 52391 48163
rect 52357 48089 52391 48091
rect 52357 48053 52391 48055
rect 52357 47981 52391 47987
rect 52357 47909 52391 47919
rect 52357 47837 52391 47851
rect 52357 47765 52391 47783
rect 52357 47693 52391 47715
rect 52357 47621 52391 47647
rect 52357 47549 52391 47579
rect 52357 47477 52391 47511
rect 52357 47342 52391 47443
rect 23848 47229 23908 47312
rect 24830 47282 52438 47342
rect 23848 47195 23861 47229
rect 23895 47195 23908 47229
rect 23998 47263 24434 47276
rect 23998 47243 24101 47263
rect 23998 47216 24041 47243
rect 24075 47229 24101 47243
rect 24135 47229 24434 47263
rect 24075 47216 24434 47229
rect 24830 47223 29469 47236
rect 23848 47102 23908 47195
rect 24830 47189 25013 47223
rect 25047 47189 25413 47223
rect 25447 47189 25813 47223
rect 25847 47189 26213 47223
rect 26247 47189 26613 47223
rect 26647 47189 27013 47223
rect 27047 47189 27413 47223
rect 27447 47189 27813 47223
rect 27847 47189 28213 47223
rect 28247 47189 28613 47223
rect 28647 47189 29013 47223
rect 29047 47189 29413 47223
rect 29447 47209 29469 47223
rect 29503 47223 52438 47236
rect 29503 47209 29813 47223
rect 29447 47189 29813 47209
rect 29847 47189 30213 47223
rect 30247 47189 30613 47223
rect 30647 47189 31013 47223
rect 31047 47189 31413 47223
rect 31447 47189 31813 47223
rect 31847 47189 32213 47223
rect 32247 47189 32613 47223
rect 32647 47189 33013 47223
rect 33047 47189 33413 47223
rect 33447 47189 33813 47223
rect 33847 47189 34213 47223
rect 34247 47189 34613 47223
rect 34647 47189 35013 47223
rect 35047 47189 35413 47223
rect 35447 47189 35813 47223
rect 35847 47189 36213 47223
rect 36247 47189 36613 47223
rect 36647 47189 37013 47223
rect 37047 47189 37413 47223
rect 37447 47189 37813 47223
rect 37847 47189 38213 47223
rect 38247 47189 38613 47223
rect 38647 47189 39013 47223
rect 39047 47189 39413 47223
rect 39447 47189 39813 47223
rect 39847 47189 40213 47223
rect 40247 47189 40613 47223
rect 40647 47189 41013 47223
rect 41047 47189 41413 47223
rect 41447 47189 41813 47223
rect 41847 47189 42213 47223
rect 42247 47189 42613 47223
rect 42647 47189 43013 47223
rect 43047 47189 43413 47223
rect 43447 47189 43813 47223
rect 43847 47189 44213 47223
rect 44247 47189 44613 47223
rect 44647 47189 45013 47223
rect 45047 47189 45413 47223
rect 45447 47189 45813 47223
rect 45847 47189 46213 47223
rect 46247 47189 46613 47223
rect 46647 47189 47013 47223
rect 47047 47189 47413 47223
rect 47447 47189 47813 47223
rect 47847 47189 48213 47223
rect 48247 47189 48613 47223
rect 48647 47189 49013 47223
rect 49047 47189 49413 47223
rect 49447 47189 49813 47223
rect 49847 47189 50213 47223
rect 50247 47189 50613 47223
rect 50647 47189 51013 47223
rect 51047 47189 51413 47223
rect 51447 47189 51813 47223
rect 51847 47189 52213 47223
rect 52247 47189 52438 47223
rect 24830 47176 52438 47189
rect 5918 47089 13086 47102
rect 5918 47055 6101 47089
rect 6135 47055 6501 47089
rect 6535 47055 6901 47089
rect 6935 47055 7301 47089
rect 7335 47055 7701 47089
rect 7735 47055 8101 47089
rect 8135 47055 8501 47089
rect 8535 47055 8901 47089
rect 8935 47055 9301 47089
rect 9335 47055 9701 47089
rect 9735 47055 10101 47089
rect 10135 47055 10501 47089
rect 10535 47055 10901 47089
rect 10935 47055 11301 47089
rect 11335 47055 11701 47089
rect 11735 47055 12101 47089
rect 12135 47055 12501 47089
rect 12535 47055 12901 47089
rect 12935 47055 13086 47089
rect 5918 47042 13086 47055
rect 13366 47089 20534 47102
rect 13366 47055 13549 47089
rect 13583 47055 13949 47089
rect 13983 47055 14349 47089
rect 14383 47055 14749 47089
rect 14783 47055 15149 47089
rect 15183 47055 15549 47089
rect 15583 47055 15949 47089
rect 15983 47055 16349 47089
rect 16383 47055 16749 47089
rect 16783 47055 17149 47089
rect 17183 47055 17549 47089
rect 17583 47055 17949 47089
rect 17983 47055 18349 47089
rect 18383 47055 18749 47089
rect 18783 47055 19149 47089
rect 19183 47055 19549 47089
rect 19583 47055 19949 47089
rect 19983 47055 20349 47089
rect 20383 47055 20534 47089
rect 13366 47042 20534 47055
rect 20832 47089 23272 47102
rect 20832 47055 21015 47089
rect 21049 47055 21215 47089
rect 21249 47055 21415 47089
rect 21449 47055 21615 47089
rect 21649 47055 21815 47089
rect 21849 47055 22015 47089
rect 22049 47055 22215 47089
rect 22249 47055 22415 47089
rect 22449 47055 22615 47089
rect 22649 47055 22815 47089
rect 22849 47055 23015 47089
rect 23049 47055 23272 47089
rect 20832 47042 23272 47055
rect 23820 47089 24434 47102
rect 23820 47055 24101 47089
rect 24135 47055 24434 47089
rect 23820 47042 24434 47055
rect 24732 47089 52438 47102
rect 24732 47055 25013 47089
rect 25047 47055 25413 47089
rect 25447 47055 25813 47089
rect 25847 47055 26213 47089
rect 26247 47055 26613 47089
rect 26647 47055 27013 47089
rect 27047 47055 27413 47089
rect 27447 47055 27813 47089
rect 27847 47055 28213 47089
rect 28247 47055 28613 47089
rect 28647 47055 29013 47089
rect 29047 47055 29413 47089
rect 29447 47055 29813 47089
rect 29847 47055 30213 47089
rect 30247 47055 30613 47089
rect 30647 47055 31013 47089
rect 31047 47055 31413 47089
rect 31447 47055 31813 47089
rect 31847 47055 32213 47089
rect 32247 47055 32613 47089
rect 32647 47055 33013 47089
rect 33047 47055 33413 47089
rect 33447 47055 33813 47089
rect 33847 47055 34213 47089
rect 34247 47055 34613 47089
rect 34647 47055 35013 47089
rect 35047 47055 35413 47089
rect 35447 47055 35813 47089
rect 35847 47055 36213 47089
rect 36247 47055 36613 47089
rect 36647 47055 37013 47089
rect 37047 47055 37413 47089
rect 37447 47055 37813 47089
rect 37847 47055 38213 47089
rect 38247 47055 38613 47089
rect 38647 47055 39013 47089
rect 39047 47055 39413 47089
rect 39447 47055 39813 47089
rect 39847 47055 40213 47089
rect 40247 47055 40613 47089
rect 40647 47055 41013 47089
rect 41047 47055 41413 47089
rect 41447 47055 41813 47089
rect 41847 47055 42213 47089
rect 42247 47055 42613 47089
rect 42647 47055 43013 47089
rect 43047 47055 43413 47089
rect 43447 47055 43813 47089
rect 43847 47055 44213 47089
rect 44247 47055 44613 47089
rect 44647 47055 45013 47089
rect 45047 47055 45413 47089
rect 45447 47055 45813 47089
rect 45847 47055 46213 47089
rect 46247 47055 46613 47089
rect 46647 47055 47013 47089
rect 47047 47055 47413 47089
rect 47447 47055 47813 47089
rect 47847 47055 48213 47089
rect 48247 47055 48613 47089
rect 48647 47055 49013 47089
rect 49047 47055 49413 47089
rect 49447 47055 49813 47089
rect 49847 47055 50213 47089
rect 50247 47055 50613 47089
rect 50647 47055 51013 47089
rect 51047 47055 51413 47089
rect 51447 47055 51813 47089
rect 51847 47055 52213 47089
rect 52247 47055 52438 47089
rect 24732 47042 52438 47055
rect 5918 45209 13086 45222
rect 5918 45175 6101 45209
rect 6135 45175 6501 45209
rect 6535 45175 6901 45209
rect 6935 45175 7301 45209
rect 7335 45175 7701 45209
rect 7735 45175 8101 45209
rect 8135 45175 8501 45209
rect 8535 45175 8901 45209
rect 8935 45175 9301 45209
rect 9335 45175 9701 45209
rect 9735 45175 10101 45209
rect 10135 45175 10501 45209
rect 10535 45175 10901 45209
rect 10935 45175 11301 45209
rect 11335 45175 11701 45209
rect 11735 45175 12101 45209
rect 12135 45175 12501 45209
rect 12535 45175 12901 45209
rect 12935 45175 13086 45209
rect 5918 45162 13086 45175
rect 14020 45209 14634 45222
rect 14020 45175 14301 45209
rect 14335 45175 14634 45209
rect 14020 45162 14634 45175
rect 14932 45209 42638 45222
rect 14932 45175 15213 45209
rect 15247 45175 15613 45209
rect 15647 45175 16013 45209
rect 16047 45175 16413 45209
rect 16447 45175 16813 45209
rect 16847 45175 17213 45209
rect 17247 45175 17613 45209
rect 17647 45175 18013 45209
rect 18047 45175 18413 45209
rect 18447 45175 18813 45209
rect 18847 45175 19213 45209
rect 19247 45175 19613 45209
rect 19647 45175 20013 45209
rect 20047 45175 20413 45209
rect 20447 45175 20813 45209
rect 20847 45175 21213 45209
rect 21247 45175 21613 45209
rect 21647 45175 22013 45209
rect 22047 45175 22413 45209
rect 22447 45175 22813 45209
rect 22847 45175 23213 45209
rect 23247 45175 23613 45209
rect 23647 45175 24013 45209
rect 24047 45175 24413 45209
rect 24447 45175 24813 45209
rect 24847 45175 25213 45209
rect 25247 45175 25613 45209
rect 25647 45175 26013 45209
rect 26047 45175 26413 45209
rect 26447 45175 26813 45209
rect 26847 45175 27213 45209
rect 27247 45175 27613 45209
rect 27647 45175 28013 45209
rect 28047 45175 28413 45209
rect 28447 45175 28813 45209
rect 28847 45175 29213 45209
rect 29247 45175 29613 45209
rect 29647 45175 30013 45209
rect 30047 45175 30413 45209
rect 30447 45175 30813 45209
rect 30847 45175 31213 45209
rect 31247 45175 31613 45209
rect 31647 45175 32013 45209
rect 32047 45175 32413 45209
rect 32447 45175 32813 45209
rect 32847 45175 33213 45209
rect 33247 45175 33613 45209
rect 33647 45175 34013 45209
rect 34047 45175 34413 45209
rect 34447 45175 34813 45209
rect 34847 45175 35213 45209
rect 35247 45175 35613 45209
rect 35647 45175 36013 45209
rect 36047 45175 36413 45209
rect 36447 45175 36813 45209
rect 36847 45175 37213 45209
rect 37247 45175 37613 45209
rect 37647 45175 38013 45209
rect 38047 45175 38413 45209
rect 38447 45175 38813 45209
rect 38847 45175 39213 45209
rect 39247 45175 39613 45209
rect 39647 45175 40013 45209
rect 40047 45175 40413 45209
rect 40447 45175 40813 45209
rect 40847 45175 41213 45209
rect 41247 45175 41613 45209
rect 41647 45175 42013 45209
rect 42047 45175 42413 45209
rect 42447 45175 42638 45209
rect 14932 45162 42638 45175
rect 42960 45209 52340 45222
rect 42960 45175 43143 45209
rect 43177 45175 43343 45209
rect 43377 45175 43543 45209
rect 43577 45175 43743 45209
rect 43777 45175 43943 45209
rect 43977 45175 44143 45209
rect 44177 45175 44343 45209
rect 44377 45175 44543 45209
rect 44577 45175 44743 45209
rect 44777 45175 44943 45209
rect 44977 45175 45143 45209
rect 45177 45175 45343 45209
rect 45377 45175 45543 45209
rect 45577 45175 45743 45209
rect 45777 45175 45943 45209
rect 45977 45175 46143 45209
rect 46177 45175 46343 45209
rect 46377 45175 46543 45209
rect 46577 45175 46743 45209
rect 46777 45175 46943 45209
rect 46977 45175 47143 45209
rect 47177 45175 47343 45209
rect 47377 45175 47543 45209
rect 47577 45175 47743 45209
rect 47777 45175 47943 45209
rect 47977 45175 48143 45209
rect 48177 45175 48343 45209
rect 48377 45175 48543 45209
rect 48577 45175 48743 45209
rect 48777 45175 48943 45209
rect 48977 45175 49143 45209
rect 49177 45175 49343 45209
rect 49377 45175 49543 45209
rect 49577 45175 49743 45209
rect 49777 45175 49943 45209
rect 49977 45175 50143 45209
rect 50177 45175 50343 45209
rect 50377 45175 50543 45209
rect 50577 45175 50743 45209
rect 50777 45175 50943 45209
rect 50977 45175 51143 45209
rect 51177 45175 51343 45209
rect 51377 45175 51543 45209
rect 51577 45175 51743 45209
rect 51777 45175 51943 45209
rect 51977 45175 52143 45209
rect 52177 45175 52340 45209
rect 42960 45162 52340 45175
rect 14960 45069 15020 45162
rect 16008 45119 16168 45162
rect 16008 45085 16073 45119
rect 16107 45085 16168 45119
rect 16008 45082 16168 45085
rect 17308 45119 17468 45162
rect 17308 45085 17373 45119
rect 17407 45085 17468 45119
rect 17308 45082 17468 45085
rect 18608 45119 18768 45162
rect 18608 45085 18673 45119
rect 18707 45085 18768 45119
rect 18608 45082 18768 45085
rect 19908 45119 20068 45162
rect 19908 45085 19973 45119
rect 20007 45085 20068 45119
rect 19908 45082 20068 45085
rect 21208 45119 21368 45162
rect 21208 45085 21273 45119
rect 21307 45085 21368 45119
rect 21208 45082 21368 45085
rect 22508 45119 22668 45162
rect 22508 45085 22573 45119
rect 22607 45085 22668 45119
rect 22508 45082 22668 45085
rect 23808 45119 23968 45162
rect 23808 45085 23873 45119
rect 23907 45085 23968 45119
rect 23808 45082 23968 45085
rect 25108 45119 25268 45162
rect 25108 45085 25173 45119
rect 25207 45085 25268 45119
rect 25108 45082 25268 45085
rect 26408 45119 26568 45162
rect 26408 45085 26473 45119
rect 26507 45085 26568 45119
rect 26408 45082 26568 45085
rect 27708 45119 27868 45162
rect 27708 45085 27773 45119
rect 27807 45085 27868 45119
rect 27708 45082 27868 45085
rect 29008 45119 29168 45162
rect 29008 45085 29073 45119
rect 29107 45085 29168 45119
rect 29008 45082 29168 45085
rect 30308 45119 30468 45162
rect 30308 45085 30373 45119
rect 30407 45085 30468 45119
rect 30308 45082 30468 45085
rect 31608 45119 31768 45162
rect 31608 45085 31673 45119
rect 31707 45085 31768 45119
rect 31608 45082 31768 45085
rect 32908 45119 33068 45162
rect 32908 45085 32973 45119
rect 33007 45085 33068 45119
rect 32908 45082 33068 45085
rect 34208 45119 34368 45162
rect 34208 45085 34273 45119
rect 34307 45085 34368 45119
rect 34208 45082 34368 45085
rect 35508 45119 35668 45162
rect 35508 45085 35573 45119
rect 35607 45085 35668 45119
rect 35508 45082 35668 45085
rect 36808 45119 36968 45162
rect 36808 45085 36873 45119
rect 36907 45085 36968 45119
rect 36808 45082 36968 45085
rect 38108 45119 38268 45162
rect 38108 45085 38173 45119
rect 38207 45085 38268 45119
rect 38108 45082 38268 45085
rect 39408 45119 39568 45162
rect 39408 45085 39473 45119
rect 39507 45085 39568 45119
rect 39408 45082 39568 45085
rect 40708 45119 40868 45162
rect 40708 45085 40773 45119
rect 40807 45085 40868 45119
rect 40708 45082 40868 45085
rect 14118 45002 14634 45062
rect 14960 45035 14973 45069
rect 15007 45035 15020 45069
rect 14587 44716 14621 45002
rect 14960 44952 15020 45035
rect 15090 45002 42638 45042
rect 15077 44941 15111 44961
rect 15077 44873 15111 44907
rect 15077 44805 15111 44835
rect 15077 44737 15111 44763
rect 14130 44689 14164 44716
rect 14587 44698 14622 44716
rect 14130 44617 14164 44635
rect 14130 44545 14164 44567
rect 14130 44473 14164 44499
rect 14130 44401 14164 44431
rect 14130 44329 14164 44363
rect 14130 44261 14164 44295
rect 14130 44193 14164 44223
rect 14130 44125 14164 44151
rect 14130 44057 14164 44079
rect 14130 43989 14164 44007
rect 14129 43935 14130 43966
rect 14129 43908 14164 43935
rect 14588 44689 14622 44698
rect 14588 44617 14622 44635
rect 14588 44545 14622 44567
rect 14588 44473 14622 44499
rect 14588 44401 14622 44431
rect 14588 44329 14622 44363
rect 14588 44261 14622 44295
rect 14588 44193 14622 44223
rect 14588 44125 14622 44151
rect 14588 44057 14622 44079
rect 14588 43989 14622 44007
rect 14588 43908 14622 43935
rect 15077 44669 15111 44691
rect 15077 44601 15111 44619
rect 15077 44533 15111 44547
rect 15077 44465 15111 44475
rect 15077 44397 15111 44403
rect 15077 44329 15111 44331
rect 15077 44293 15111 44295
rect 15077 44221 15111 44227
rect 15077 44149 15111 44159
rect 15077 44077 15111 44091
rect 15077 44005 15111 44023
rect 15077 43933 15111 43955
rect 14129 43742 14163 43908
rect 15077 43861 15111 43887
rect 15077 43789 15111 43819
rect 14118 43707 14634 43742
rect 14118 43682 14381 43707
rect 14415 43682 14634 43707
rect 15077 43717 15111 43751
rect 15077 43582 15111 43683
rect 15535 44941 15569 45002
rect 15535 44873 15569 44907
rect 15535 44805 15569 44835
rect 15535 44737 15569 44763
rect 15535 44669 15569 44691
rect 15535 44601 15569 44619
rect 15535 44533 15569 44547
rect 15535 44465 15569 44475
rect 15535 44397 15569 44403
rect 15535 44329 15569 44331
rect 15535 44293 15569 44295
rect 15535 44221 15569 44227
rect 15535 44149 15569 44159
rect 15535 44077 15569 44091
rect 15535 44005 15569 44023
rect 15535 43933 15569 43955
rect 15535 43861 15569 43887
rect 15535 43789 15569 43819
rect 15535 43717 15569 43751
rect 15535 43663 15569 43683
rect 15993 44941 16027 44961
rect 15993 44873 16027 44907
rect 15993 44805 16027 44835
rect 15993 44737 16027 44763
rect 15993 44669 16027 44691
rect 15993 44601 16027 44619
rect 15993 44533 16027 44547
rect 15993 44465 16027 44475
rect 15993 44397 16027 44403
rect 15993 44329 16027 44331
rect 15993 44293 16027 44295
rect 15993 44221 16027 44227
rect 15993 44149 16027 44159
rect 15993 44077 16027 44091
rect 15993 44005 16027 44023
rect 15993 43933 16027 43955
rect 15993 43861 16027 43887
rect 15993 43789 16027 43819
rect 15993 43717 16027 43751
rect 15993 43582 16027 43683
rect 16451 44941 16485 45002
rect 16451 44873 16485 44907
rect 16451 44805 16485 44835
rect 16451 44737 16485 44763
rect 16451 44669 16485 44691
rect 16451 44601 16485 44619
rect 16451 44533 16485 44547
rect 16451 44465 16485 44475
rect 16451 44397 16485 44403
rect 16451 44329 16485 44331
rect 16451 44293 16485 44295
rect 16451 44221 16485 44227
rect 16451 44149 16485 44159
rect 16451 44077 16485 44091
rect 16451 44005 16485 44023
rect 16451 43933 16485 43955
rect 16451 43861 16485 43887
rect 16451 43789 16485 43819
rect 16451 43717 16485 43751
rect 16451 43663 16485 43683
rect 16909 44941 16943 44961
rect 16909 44873 16943 44907
rect 16909 44805 16943 44835
rect 16909 44737 16943 44763
rect 16909 44669 16943 44691
rect 16909 44601 16943 44619
rect 16909 44533 16943 44547
rect 16909 44465 16943 44475
rect 16909 44397 16943 44403
rect 16909 44329 16943 44331
rect 16909 44293 16943 44295
rect 16909 44221 16943 44227
rect 16909 44149 16943 44159
rect 16909 44077 16943 44091
rect 16909 44005 16943 44023
rect 16909 43933 16943 43955
rect 16909 43861 16943 43887
rect 16909 43789 16943 43819
rect 16909 43717 16943 43751
rect 16909 43582 16943 43683
rect 17367 44941 17401 45002
rect 17367 44873 17401 44907
rect 17367 44805 17401 44835
rect 17367 44737 17401 44763
rect 17367 44669 17401 44691
rect 17367 44601 17401 44619
rect 17367 44533 17401 44547
rect 17367 44465 17401 44475
rect 17367 44397 17401 44403
rect 17367 44329 17401 44331
rect 17367 44293 17401 44295
rect 17367 44221 17401 44227
rect 17367 44149 17401 44159
rect 17367 44077 17401 44091
rect 17367 44005 17401 44023
rect 17367 43933 17401 43955
rect 17367 43861 17401 43887
rect 17367 43789 17401 43819
rect 17367 43717 17401 43751
rect 17367 43663 17401 43683
rect 17825 44941 17859 44961
rect 17825 44873 17859 44907
rect 17825 44805 17859 44835
rect 17825 44737 17859 44763
rect 17825 44669 17859 44691
rect 17825 44601 17859 44619
rect 17825 44533 17859 44547
rect 17825 44465 17859 44475
rect 17825 44397 17859 44403
rect 17825 44329 17859 44331
rect 17825 44293 17859 44295
rect 17825 44221 17859 44227
rect 17825 44149 17859 44159
rect 17825 44077 17859 44091
rect 17825 44005 17859 44023
rect 17825 43933 17859 43955
rect 17825 43861 17859 43887
rect 17825 43789 17859 43819
rect 17825 43717 17859 43751
rect 17825 43582 17859 43683
rect 18283 44941 18317 45002
rect 18283 44873 18317 44907
rect 18283 44805 18317 44835
rect 18283 44737 18317 44763
rect 18283 44669 18317 44691
rect 18283 44601 18317 44619
rect 18283 44533 18317 44547
rect 18283 44465 18317 44475
rect 18283 44397 18317 44403
rect 18283 44329 18317 44331
rect 18283 44293 18317 44295
rect 18283 44221 18317 44227
rect 18283 44149 18317 44159
rect 18283 44077 18317 44091
rect 18283 44005 18317 44023
rect 18283 43933 18317 43955
rect 18283 43861 18317 43887
rect 18283 43789 18317 43819
rect 18283 43717 18317 43751
rect 18283 43663 18317 43683
rect 18741 44941 18775 44961
rect 18741 44873 18775 44907
rect 18741 44805 18775 44835
rect 18741 44737 18775 44763
rect 18741 44669 18775 44691
rect 18741 44601 18775 44619
rect 18741 44533 18775 44547
rect 18741 44465 18775 44475
rect 18741 44397 18775 44403
rect 18741 44329 18775 44331
rect 18741 44293 18775 44295
rect 18741 44221 18775 44227
rect 18741 44149 18775 44159
rect 18741 44077 18775 44091
rect 18741 44005 18775 44023
rect 18741 43933 18775 43955
rect 18741 43861 18775 43887
rect 18741 43789 18775 43819
rect 18741 43717 18775 43751
rect 18741 43582 18775 43683
rect 19199 44941 19233 45002
rect 19199 44873 19233 44907
rect 19199 44805 19233 44835
rect 19199 44737 19233 44763
rect 19199 44669 19233 44691
rect 19199 44601 19233 44619
rect 19199 44533 19233 44547
rect 19199 44465 19233 44475
rect 19199 44397 19233 44403
rect 19199 44329 19233 44331
rect 19199 44293 19233 44295
rect 19199 44221 19233 44227
rect 19199 44149 19233 44159
rect 19199 44077 19233 44091
rect 19199 44005 19233 44023
rect 19199 43933 19233 43955
rect 19199 43861 19233 43887
rect 19199 43789 19233 43819
rect 19199 43717 19233 43751
rect 19199 43663 19233 43683
rect 19657 44941 19691 44961
rect 19657 44873 19691 44907
rect 19657 44805 19691 44835
rect 19657 44737 19691 44763
rect 19657 44669 19691 44691
rect 19657 44601 19691 44619
rect 19657 44533 19691 44547
rect 19657 44465 19691 44475
rect 19657 44397 19691 44403
rect 19657 44329 19691 44331
rect 19657 44293 19691 44295
rect 19657 44221 19691 44227
rect 19657 44149 19691 44159
rect 19657 44077 19691 44091
rect 19657 44005 19691 44023
rect 19657 43933 19691 43955
rect 19657 43861 19691 43887
rect 19657 43789 19691 43819
rect 19657 43717 19691 43751
rect 19657 43582 19691 43683
rect 20115 44941 20149 45002
rect 20115 44873 20149 44907
rect 20115 44805 20149 44835
rect 20115 44737 20149 44763
rect 20115 44669 20149 44691
rect 20115 44601 20149 44619
rect 20115 44533 20149 44547
rect 20115 44465 20149 44475
rect 20115 44397 20149 44403
rect 20115 44329 20149 44331
rect 20115 44293 20149 44295
rect 20115 44221 20149 44227
rect 20115 44149 20149 44159
rect 20115 44077 20149 44091
rect 20115 44005 20149 44023
rect 20115 43933 20149 43955
rect 20115 43861 20149 43887
rect 20115 43789 20149 43819
rect 20115 43717 20149 43751
rect 20115 43663 20149 43683
rect 20573 44941 20607 44961
rect 20573 44873 20607 44907
rect 20573 44805 20607 44835
rect 20573 44737 20607 44763
rect 20573 44669 20607 44691
rect 20573 44601 20607 44619
rect 20573 44533 20607 44547
rect 20573 44465 20607 44475
rect 20573 44397 20607 44403
rect 20573 44329 20607 44331
rect 20573 44293 20607 44295
rect 20573 44221 20607 44227
rect 20573 44149 20607 44159
rect 20573 44077 20607 44091
rect 20573 44005 20607 44023
rect 20573 43933 20607 43955
rect 20573 43861 20607 43887
rect 20573 43789 20607 43819
rect 20573 43717 20607 43751
rect 20573 43582 20607 43683
rect 21031 44941 21065 45002
rect 21031 44873 21065 44907
rect 21031 44805 21065 44835
rect 21031 44737 21065 44763
rect 21031 44669 21065 44691
rect 21031 44601 21065 44619
rect 21031 44533 21065 44547
rect 21031 44465 21065 44475
rect 21031 44397 21065 44403
rect 21031 44329 21065 44331
rect 21031 44293 21065 44295
rect 21031 44221 21065 44227
rect 21031 44149 21065 44159
rect 21031 44077 21065 44091
rect 21031 44005 21065 44023
rect 21031 43933 21065 43955
rect 21031 43861 21065 43887
rect 21031 43789 21065 43819
rect 21031 43717 21065 43751
rect 21031 43663 21065 43683
rect 21489 44941 21523 44961
rect 21489 44873 21523 44907
rect 21489 44805 21523 44835
rect 21489 44737 21523 44763
rect 21489 44669 21523 44691
rect 21489 44601 21523 44619
rect 21489 44533 21523 44547
rect 21489 44465 21523 44475
rect 21489 44397 21523 44403
rect 21489 44329 21523 44331
rect 21489 44293 21523 44295
rect 21489 44221 21523 44227
rect 21489 44149 21523 44159
rect 21489 44077 21523 44091
rect 21489 44005 21523 44023
rect 21489 43933 21523 43955
rect 21489 43861 21523 43887
rect 21489 43789 21523 43819
rect 21489 43717 21523 43751
rect 21489 43582 21523 43683
rect 21947 44941 21981 45002
rect 21947 44873 21981 44907
rect 21947 44805 21981 44835
rect 21947 44737 21981 44763
rect 21947 44669 21981 44691
rect 21947 44601 21981 44619
rect 21947 44533 21981 44547
rect 21947 44465 21981 44475
rect 21947 44397 21981 44403
rect 21947 44329 21981 44331
rect 21947 44293 21981 44295
rect 21947 44221 21981 44227
rect 21947 44149 21981 44159
rect 21947 44077 21981 44091
rect 21947 44005 21981 44023
rect 21947 43933 21981 43955
rect 21947 43861 21981 43887
rect 21947 43789 21981 43819
rect 21947 43717 21981 43751
rect 21947 43663 21981 43683
rect 22405 44941 22439 44961
rect 22405 44873 22439 44907
rect 22405 44805 22439 44835
rect 22405 44737 22439 44763
rect 22405 44669 22439 44691
rect 22405 44601 22439 44619
rect 22405 44533 22439 44547
rect 22405 44465 22439 44475
rect 22405 44397 22439 44403
rect 22405 44329 22439 44331
rect 22405 44293 22439 44295
rect 22405 44221 22439 44227
rect 22405 44149 22439 44159
rect 22405 44077 22439 44091
rect 22405 44005 22439 44023
rect 22405 43933 22439 43955
rect 22405 43861 22439 43887
rect 22405 43789 22439 43819
rect 22405 43717 22439 43751
rect 22405 43582 22439 43683
rect 22863 44941 22897 45002
rect 22863 44873 22897 44907
rect 22863 44805 22897 44835
rect 22863 44737 22897 44763
rect 22863 44669 22897 44691
rect 22863 44601 22897 44619
rect 22863 44533 22897 44547
rect 22863 44465 22897 44475
rect 22863 44397 22897 44403
rect 22863 44329 22897 44331
rect 22863 44293 22897 44295
rect 22863 44221 22897 44227
rect 22863 44149 22897 44159
rect 22863 44077 22897 44091
rect 22863 44005 22897 44023
rect 22863 43933 22897 43955
rect 22863 43861 22897 43887
rect 22863 43789 22897 43819
rect 22863 43717 22897 43751
rect 22863 43663 22897 43683
rect 23321 44941 23355 44961
rect 23321 44873 23355 44907
rect 23321 44805 23355 44835
rect 23321 44737 23355 44763
rect 23321 44669 23355 44691
rect 23321 44601 23355 44619
rect 23321 44533 23355 44547
rect 23321 44465 23355 44475
rect 23321 44397 23355 44403
rect 23321 44329 23355 44331
rect 23321 44293 23355 44295
rect 23321 44221 23355 44227
rect 23321 44149 23355 44159
rect 23321 44077 23355 44091
rect 23321 44005 23355 44023
rect 23321 43933 23355 43955
rect 23321 43861 23355 43887
rect 23321 43789 23355 43819
rect 23321 43717 23355 43751
rect 23321 43582 23355 43683
rect 23779 44941 23813 45002
rect 23779 44873 23813 44907
rect 23779 44805 23813 44835
rect 23779 44737 23813 44763
rect 23779 44669 23813 44691
rect 23779 44601 23813 44619
rect 23779 44533 23813 44547
rect 23779 44465 23813 44475
rect 23779 44397 23813 44403
rect 23779 44329 23813 44331
rect 23779 44293 23813 44295
rect 23779 44221 23813 44227
rect 23779 44149 23813 44159
rect 23779 44077 23813 44091
rect 23779 44005 23813 44023
rect 23779 43933 23813 43955
rect 23779 43861 23813 43887
rect 23779 43789 23813 43819
rect 23779 43717 23813 43751
rect 23779 43663 23813 43683
rect 24237 44941 24271 44961
rect 24237 44873 24271 44907
rect 24237 44805 24271 44835
rect 24237 44737 24271 44763
rect 24237 44669 24271 44691
rect 24237 44601 24271 44619
rect 24237 44533 24271 44547
rect 24237 44465 24271 44475
rect 24237 44397 24271 44403
rect 24237 44329 24271 44331
rect 24237 44293 24271 44295
rect 24237 44221 24271 44227
rect 24237 44149 24271 44159
rect 24237 44077 24271 44091
rect 24237 44005 24271 44023
rect 24237 43933 24271 43955
rect 24237 43861 24271 43887
rect 24237 43789 24271 43819
rect 24237 43717 24271 43751
rect 24237 43582 24271 43683
rect 24695 44941 24729 45002
rect 24695 44873 24729 44907
rect 24695 44805 24729 44835
rect 24695 44737 24729 44763
rect 24695 44669 24729 44691
rect 24695 44601 24729 44619
rect 24695 44533 24729 44547
rect 24695 44465 24729 44475
rect 24695 44397 24729 44403
rect 24695 44329 24729 44331
rect 24695 44293 24729 44295
rect 24695 44221 24729 44227
rect 24695 44149 24729 44159
rect 24695 44077 24729 44091
rect 24695 44005 24729 44023
rect 24695 43933 24729 43955
rect 24695 43861 24729 43887
rect 24695 43789 24729 43819
rect 24695 43717 24729 43751
rect 24695 43663 24729 43683
rect 25153 44941 25187 44961
rect 25153 44873 25187 44907
rect 25153 44805 25187 44835
rect 25153 44737 25187 44763
rect 25153 44669 25187 44691
rect 25153 44601 25187 44619
rect 25153 44533 25187 44547
rect 25153 44465 25187 44475
rect 25153 44397 25187 44403
rect 25153 44329 25187 44331
rect 25153 44293 25187 44295
rect 25153 44221 25187 44227
rect 25153 44149 25187 44159
rect 25153 44077 25187 44091
rect 25153 44005 25187 44023
rect 25153 43933 25187 43955
rect 25153 43861 25187 43887
rect 25153 43789 25187 43819
rect 25153 43717 25187 43751
rect 25153 43582 25187 43683
rect 25611 44941 25645 45002
rect 25611 44873 25645 44907
rect 25611 44805 25645 44835
rect 25611 44737 25645 44763
rect 25611 44669 25645 44691
rect 25611 44601 25645 44619
rect 25611 44533 25645 44547
rect 25611 44465 25645 44475
rect 25611 44397 25645 44403
rect 25611 44329 25645 44331
rect 25611 44293 25645 44295
rect 25611 44221 25645 44227
rect 25611 44149 25645 44159
rect 25611 44077 25645 44091
rect 25611 44005 25645 44023
rect 25611 43933 25645 43955
rect 25611 43861 25645 43887
rect 25611 43789 25645 43819
rect 25611 43717 25645 43751
rect 25611 43663 25645 43683
rect 26069 44941 26103 44961
rect 26069 44873 26103 44907
rect 26069 44805 26103 44835
rect 26069 44737 26103 44763
rect 26069 44669 26103 44691
rect 26069 44601 26103 44619
rect 26069 44533 26103 44547
rect 26069 44465 26103 44475
rect 26069 44397 26103 44403
rect 26069 44329 26103 44331
rect 26069 44293 26103 44295
rect 26069 44221 26103 44227
rect 26069 44149 26103 44159
rect 26069 44077 26103 44091
rect 26069 44005 26103 44023
rect 26069 43933 26103 43955
rect 26069 43861 26103 43887
rect 26069 43789 26103 43819
rect 26069 43717 26103 43751
rect 26069 43582 26103 43683
rect 26527 44941 26561 45002
rect 26527 44873 26561 44907
rect 26527 44805 26561 44835
rect 26527 44737 26561 44763
rect 26527 44669 26561 44691
rect 26527 44601 26561 44619
rect 26527 44533 26561 44547
rect 26527 44465 26561 44475
rect 26527 44397 26561 44403
rect 26527 44329 26561 44331
rect 26527 44293 26561 44295
rect 26527 44221 26561 44227
rect 26527 44149 26561 44159
rect 26527 44077 26561 44091
rect 26527 44005 26561 44023
rect 26527 43933 26561 43955
rect 26527 43861 26561 43887
rect 26527 43789 26561 43819
rect 26527 43717 26561 43751
rect 26527 43663 26561 43683
rect 26985 44941 27019 44961
rect 26985 44873 27019 44907
rect 26985 44805 27019 44835
rect 26985 44737 27019 44763
rect 26985 44669 27019 44691
rect 26985 44601 27019 44619
rect 26985 44533 27019 44547
rect 26985 44465 27019 44475
rect 26985 44397 27019 44403
rect 26985 44329 27019 44331
rect 26985 44293 27019 44295
rect 26985 44221 27019 44227
rect 26985 44149 27019 44159
rect 26985 44077 27019 44091
rect 26985 44005 27019 44023
rect 26985 43933 27019 43955
rect 26985 43861 27019 43887
rect 26985 43789 27019 43819
rect 26985 43717 27019 43751
rect 26985 43582 27019 43683
rect 27443 44941 27477 45002
rect 27443 44873 27477 44907
rect 27443 44805 27477 44835
rect 27443 44737 27477 44763
rect 27443 44669 27477 44691
rect 27443 44601 27477 44619
rect 27443 44533 27477 44547
rect 27443 44465 27477 44475
rect 27443 44397 27477 44403
rect 27443 44329 27477 44331
rect 27443 44293 27477 44295
rect 27443 44221 27477 44227
rect 27443 44149 27477 44159
rect 27443 44077 27477 44091
rect 27443 44005 27477 44023
rect 27443 43933 27477 43955
rect 27443 43861 27477 43887
rect 27443 43789 27477 43819
rect 27443 43717 27477 43751
rect 27443 43663 27477 43683
rect 27901 44941 27935 44961
rect 27901 44873 27935 44907
rect 27901 44805 27935 44835
rect 27901 44737 27935 44763
rect 27901 44669 27935 44691
rect 27901 44601 27935 44619
rect 27901 44533 27935 44547
rect 27901 44465 27935 44475
rect 27901 44397 27935 44403
rect 27901 44329 27935 44331
rect 27901 44293 27935 44295
rect 27901 44221 27935 44227
rect 27901 44149 27935 44159
rect 27901 44077 27935 44091
rect 27901 44005 27935 44023
rect 27901 43933 27935 43955
rect 27901 43861 27935 43887
rect 27901 43789 27935 43819
rect 27901 43717 27935 43751
rect 27901 43582 27935 43683
rect 28359 44941 28393 45002
rect 28359 44873 28393 44907
rect 28359 44805 28393 44835
rect 28359 44737 28393 44763
rect 28359 44669 28393 44691
rect 28359 44601 28393 44619
rect 28359 44533 28393 44547
rect 28359 44465 28393 44475
rect 28359 44397 28393 44403
rect 28359 44329 28393 44331
rect 28359 44293 28393 44295
rect 28359 44221 28393 44227
rect 28359 44149 28393 44159
rect 28359 44077 28393 44091
rect 28359 44005 28393 44023
rect 28359 43933 28393 43955
rect 28359 43861 28393 43887
rect 28359 43789 28393 43819
rect 28359 43717 28393 43751
rect 28359 43663 28393 43683
rect 28817 44941 28851 44961
rect 28817 44873 28851 44907
rect 28817 44805 28851 44835
rect 28817 44737 28851 44763
rect 28817 44669 28851 44691
rect 28817 44601 28851 44619
rect 28817 44533 28851 44547
rect 28817 44465 28851 44475
rect 28817 44397 28851 44403
rect 28817 44329 28851 44331
rect 28817 44293 28851 44295
rect 28817 44221 28851 44227
rect 28817 44149 28851 44159
rect 28817 44077 28851 44091
rect 28817 44005 28851 44023
rect 28817 43933 28851 43955
rect 28817 43861 28851 43887
rect 28817 43789 28851 43819
rect 28817 43717 28851 43751
rect 28817 43582 28851 43683
rect 29275 44941 29309 45002
rect 29275 44873 29309 44907
rect 29275 44805 29309 44835
rect 29275 44737 29309 44763
rect 29275 44669 29309 44691
rect 29275 44601 29309 44619
rect 29275 44533 29309 44547
rect 29275 44465 29309 44475
rect 29275 44397 29309 44403
rect 29275 44329 29309 44331
rect 29275 44293 29309 44295
rect 29275 44221 29309 44227
rect 29275 44149 29309 44159
rect 29275 44077 29309 44091
rect 29275 44005 29309 44023
rect 29275 43933 29309 43955
rect 29275 43861 29309 43887
rect 29275 43789 29309 43819
rect 29275 43717 29309 43751
rect 29275 43663 29309 43683
rect 29733 44941 29767 44961
rect 29733 44873 29767 44907
rect 29733 44805 29767 44835
rect 29733 44737 29767 44763
rect 29733 44669 29767 44691
rect 29733 44601 29767 44619
rect 29733 44533 29767 44547
rect 29733 44465 29767 44475
rect 29733 44397 29767 44403
rect 29733 44329 29767 44331
rect 29733 44293 29767 44295
rect 29733 44221 29767 44227
rect 29733 44149 29767 44159
rect 29733 44077 29767 44091
rect 29733 44005 29767 44023
rect 29733 43933 29767 43955
rect 29733 43861 29767 43887
rect 29733 43789 29767 43819
rect 29733 43717 29767 43751
rect 29733 43582 29767 43683
rect 30191 44941 30225 45002
rect 30191 44873 30225 44907
rect 30191 44805 30225 44835
rect 30191 44737 30225 44763
rect 30191 44669 30225 44691
rect 30191 44601 30225 44619
rect 30191 44533 30225 44547
rect 30191 44465 30225 44475
rect 30191 44397 30225 44403
rect 30191 44329 30225 44331
rect 30191 44293 30225 44295
rect 30191 44221 30225 44227
rect 30191 44149 30225 44159
rect 30191 44077 30225 44091
rect 30191 44005 30225 44023
rect 30191 43933 30225 43955
rect 30191 43861 30225 43887
rect 30191 43789 30225 43819
rect 30191 43717 30225 43751
rect 30191 43663 30225 43683
rect 30649 44941 30683 44961
rect 30649 44873 30683 44907
rect 30649 44805 30683 44835
rect 30649 44737 30683 44763
rect 30649 44669 30683 44691
rect 30649 44601 30683 44619
rect 30649 44533 30683 44547
rect 30649 44465 30683 44475
rect 30649 44397 30683 44403
rect 30649 44329 30683 44331
rect 30649 44293 30683 44295
rect 30649 44221 30683 44227
rect 30649 44149 30683 44159
rect 30649 44077 30683 44091
rect 30649 44005 30683 44023
rect 30649 43933 30683 43955
rect 30649 43861 30683 43887
rect 30649 43789 30683 43819
rect 30649 43717 30683 43751
rect 30649 43582 30683 43683
rect 31107 44941 31141 45002
rect 31107 44873 31141 44907
rect 31107 44805 31141 44835
rect 31107 44737 31141 44763
rect 31107 44669 31141 44691
rect 31107 44601 31141 44619
rect 31107 44533 31141 44547
rect 31107 44465 31141 44475
rect 31107 44397 31141 44403
rect 31107 44329 31141 44331
rect 31107 44293 31141 44295
rect 31107 44221 31141 44227
rect 31107 44149 31141 44159
rect 31107 44077 31141 44091
rect 31107 44005 31141 44023
rect 31107 43933 31141 43955
rect 31107 43861 31141 43887
rect 31107 43789 31141 43819
rect 31107 43717 31141 43751
rect 31107 43663 31141 43683
rect 31565 44941 31599 44961
rect 31565 44873 31599 44907
rect 31565 44805 31599 44835
rect 31565 44737 31599 44763
rect 31565 44669 31599 44691
rect 31565 44601 31599 44619
rect 31565 44533 31599 44547
rect 31565 44465 31599 44475
rect 31565 44397 31599 44403
rect 31565 44329 31599 44331
rect 31565 44293 31599 44295
rect 31565 44221 31599 44227
rect 31565 44149 31599 44159
rect 31565 44077 31599 44091
rect 31565 44005 31599 44023
rect 31565 43933 31599 43955
rect 31565 43861 31599 43887
rect 31565 43789 31599 43819
rect 31565 43717 31599 43751
rect 31565 43582 31599 43683
rect 32023 44941 32057 45002
rect 32023 44873 32057 44907
rect 32023 44805 32057 44835
rect 32023 44737 32057 44763
rect 32023 44669 32057 44691
rect 32023 44601 32057 44619
rect 32023 44533 32057 44547
rect 32023 44465 32057 44475
rect 32023 44397 32057 44403
rect 32023 44329 32057 44331
rect 32023 44293 32057 44295
rect 32023 44221 32057 44227
rect 32023 44149 32057 44159
rect 32023 44077 32057 44091
rect 32023 44005 32057 44023
rect 32023 43933 32057 43955
rect 32023 43861 32057 43887
rect 32023 43789 32057 43819
rect 32023 43717 32057 43751
rect 32023 43663 32057 43683
rect 32481 44941 32515 44961
rect 32481 44873 32515 44907
rect 32481 44805 32515 44835
rect 32481 44737 32515 44763
rect 32481 44669 32515 44691
rect 32481 44601 32515 44619
rect 32481 44533 32515 44547
rect 32481 44465 32515 44475
rect 32481 44397 32515 44403
rect 32481 44329 32515 44331
rect 32481 44293 32515 44295
rect 32481 44221 32515 44227
rect 32481 44149 32515 44159
rect 32481 44077 32515 44091
rect 32481 44005 32515 44023
rect 32481 43933 32515 43955
rect 32481 43861 32515 43887
rect 32481 43789 32515 43819
rect 32481 43717 32515 43751
rect 32481 43582 32515 43683
rect 32939 44941 32973 45002
rect 32939 44873 32973 44907
rect 32939 44805 32973 44835
rect 32939 44737 32973 44763
rect 32939 44669 32973 44691
rect 32939 44601 32973 44619
rect 32939 44533 32973 44547
rect 32939 44465 32973 44475
rect 32939 44397 32973 44403
rect 32939 44329 32973 44331
rect 32939 44293 32973 44295
rect 32939 44221 32973 44227
rect 32939 44149 32973 44159
rect 32939 44077 32973 44091
rect 32939 44005 32973 44023
rect 32939 43933 32973 43955
rect 32939 43861 32973 43887
rect 32939 43789 32973 43819
rect 32939 43717 32973 43751
rect 32939 43663 32973 43683
rect 33397 44941 33431 44961
rect 33397 44873 33431 44907
rect 33397 44805 33431 44835
rect 33397 44737 33431 44763
rect 33397 44669 33431 44691
rect 33397 44601 33431 44619
rect 33397 44533 33431 44547
rect 33397 44465 33431 44475
rect 33397 44397 33431 44403
rect 33397 44329 33431 44331
rect 33397 44293 33431 44295
rect 33397 44221 33431 44227
rect 33397 44149 33431 44159
rect 33397 44077 33431 44091
rect 33397 44005 33431 44023
rect 33397 43933 33431 43955
rect 33397 43861 33431 43887
rect 33397 43789 33431 43819
rect 33397 43717 33431 43751
rect 33397 43582 33431 43683
rect 33855 44941 33889 45002
rect 33855 44873 33889 44907
rect 33855 44805 33889 44835
rect 33855 44737 33889 44763
rect 33855 44669 33889 44691
rect 33855 44601 33889 44619
rect 33855 44533 33889 44547
rect 33855 44465 33889 44475
rect 33855 44397 33889 44403
rect 33855 44329 33889 44331
rect 33855 44293 33889 44295
rect 33855 44221 33889 44227
rect 33855 44149 33889 44159
rect 33855 44077 33889 44091
rect 33855 44005 33889 44023
rect 33855 43933 33889 43955
rect 33855 43861 33889 43887
rect 33855 43789 33889 43819
rect 33855 43717 33889 43751
rect 33855 43663 33889 43683
rect 34313 44941 34347 44961
rect 34313 44873 34347 44907
rect 34313 44805 34347 44835
rect 34313 44737 34347 44763
rect 34313 44669 34347 44691
rect 34313 44601 34347 44619
rect 34313 44533 34347 44547
rect 34313 44465 34347 44475
rect 34313 44397 34347 44403
rect 34313 44329 34347 44331
rect 34313 44293 34347 44295
rect 34313 44221 34347 44227
rect 34313 44149 34347 44159
rect 34313 44077 34347 44091
rect 34313 44005 34347 44023
rect 34313 43933 34347 43955
rect 34313 43861 34347 43887
rect 34313 43789 34347 43819
rect 34313 43717 34347 43751
rect 34313 43582 34347 43683
rect 34771 44941 34805 45002
rect 34771 44873 34805 44907
rect 34771 44805 34805 44835
rect 34771 44737 34805 44763
rect 34771 44669 34805 44691
rect 34771 44601 34805 44619
rect 34771 44533 34805 44547
rect 34771 44465 34805 44475
rect 34771 44397 34805 44403
rect 34771 44329 34805 44331
rect 34771 44293 34805 44295
rect 34771 44221 34805 44227
rect 34771 44149 34805 44159
rect 34771 44077 34805 44091
rect 34771 44005 34805 44023
rect 34771 43933 34805 43955
rect 34771 43861 34805 43887
rect 34771 43789 34805 43819
rect 34771 43717 34805 43751
rect 34771 43663 34805 43683
rect 35229 44941 35263 44961
rect 35229 44873 35263 44907
rect 35229 44805 35263 44835
rect 35229 44737 35263 44763
rect 35229 44669 35263 44691
rect 35229 44601 35263 44619
rect 35229 44533 35263 44547
rect 35229 44465 35263 44475
rect 35229 44397 35263 44403
rect 35229 44329 35263 44331
rect 35229 44293 35263 44295
rect 35229 44221 35263 44227
rect 35229 44149 35263 44159
rect 35229 44077 35263 44091
rect 35229 44005 35263 44023
rect 35229 43933 35263 43955
rect 35229 43861 35263 43887
rect 35229 43789 35263 43819
rect 35229 43717 35263 43751
rect 35229 43582 35263 43683
rect 35687 44941 35721 45002
rect 35687 44873 35721 44907
rect 35687 44805 35721 44835
rect 35687 44737 35721 44763
rect 35687 44669 35721 44691
rect 35687 44601 35721 44619
rect 35687 44533 35721 44547
rect 35687 44465 35721 44475
rect 35687 44397 35721 44403
rect 35687 44329 35721 44331
rect 35687 44293 35721 44295
rect 35687 44221 35721 44227
rect 35687 44149 35721 44159
rect 35687 44077 35721 44091
rect 35687 44005 35721 44023
rect 35687 43933 35721 43955
rect 35687 43861 35721 43887
rect 35687 43789 35721 43819
rect 35687 43717 35721 43751
rect 35687 43663 35721 43683
rect 36145 44941 36179 44961
rect 36145 44873 36179 44907
rect 36145 44805 36179 44835
rect 36145 44737 36179 44763
rect 36145 44669 36179 44691
rect 36145 44601 36179 44619
rect 36145 44533 36179 44547
rect 36145 44465 36179 44475
rect 36145 44397 36179 44403
rect 36145 44329 36179 44331
rect 36145 44293 36179 44295
rect 36145 44221 36179 44227
rect 36145 44149 36179 44159
rect 36145 44077 36179 44091
rect 36145 44005 36179 44023
rect 36145 43933 36179 43955
rect 36145 43861 36179 43887
rect 36145 43789 36179 43819
rect 36145 43717 36179 43751
rect 36145 43582 36179 43683
rect 36603 44941 36637 45002
rect 36603 44873 36637 44907
rect 36603 44805 36637 44835
rect 36603 44737 36637 44763
rect 36603 44669 36637 44691
rect 36603 44601 36637 44619
rect 36603 44533 36637 44547
rect 36603 44465 36637 44475
rect 36603 44397 36637 44403
rect 36603 44329 36637 44331
rect 36603 44293 36637 44295
rect 36603 44221 36637 44227
rect 36603 44149 36637 44159
rect 36603 44077 36637 44091
rect 36603 44005 36637 44023
rect 36603 43933 36637 43955
rect 36603 43861 36637 43887
rect 36603 43789 36637 43819
rect 36603 43717 36637 43751
rect 36603 43663 36637 43683
rect 37061 44941 37095 44961
rect 37061 44873 37095 44907
rect 37061 44805 37095 44835
rect 37061 44737 37095 44763
rect 37061 44669 37095 44691
rect 37061 44601 37095 44619
rect 37061 44533 37095 44547
rect 37061 44465 37095 44475
rect 37061 44397 37095 44403
rect 37061 44329 37095 44331
rect 37061 44293 37095 44295
rect 37061 44221 37095 44227
rect 37061 44149 37095 44159
rect 37061 44077 37095 44091
rect 37061 44005 37095 44023
rect 37061 43933 37095 43955
rect 37061 43861 37095 43887
rect 37061 43789 37095 43819
rect 37061 43717 37095 43751
rect 37061 43582 37095 43683
rect 37519 44941 37553 45002
rect 37519 44873 37553 44907
rect 37519 44805 37553 44835
rect 37519 44737 37553 44763
rect 37519 44669 37553 44691
rect 37519 44601 37553 44619
rect 37519 44533 37553 44547
rect 37519 44465 37553 44475
rect 37519 44397 37553 44403
rect 37519 44329 37553 44331
rect 37519 44293 37553 44295
rect 37519 44221 37553 44227
rect 37519 44149 37553 44159
rect 37519 44077 37553 44091
rect 37519 44005 37553 44023
rect 37519 43933 37553 43955
rect 37519 43861 37553 43887
rect 37519 43789 37553 43819
rect 37519 43717 37553 43751
rect 37519 43663 37553 43683
rect 37977 44941 38011 44961
rect 37977 44873 38011 44907
rect 37977 44805 38011 44835
rect 37977 44737 38011 44763
rect 37977 44669 38011 44691
rect 37977 44601 38011 44619
rect 37977 44533 38011 44547
rect 37977 44465 38011 44475
rect 37977 44397 38011 44403
rect 37977 44329 38011 44331
rect 37977 44293 38011 44295
rect 37977 44221 38011 44227
rect 37977 44149 38011 44159
rect 37977 44077 38011 44091
rect 37977 44005 38011 44023
rect 37977 43933 38011 43955
rect 37977 43861 38011 43887
rect 37977 43789 38011 43819
rect 37977 43717 38011 43751
rect 37977 43582 38011 43683
rect 38435 44941 38469 45002
rect 38435 44873 38469 44907
rect 38435 44805 38469 44835
rect 38435 44737 38469 44763
rect 38435 44669 38469 44691
rect 38435 44601 38469 44619
rect 38435 44533 38469 44547
rect 38435 44465 38469 44475
rect 38435 44397 38469 44403
rect 38435 44329 38469 44331
rect 38435 44293 38469 44295
rect 38435 44221 38469 44227
rect 38435 44149 38469 44159
rect 38435 44077 38469 44091
rect 38435 44005 38469 44023
rect 38435 43933 38469 43955
rect 38435 43861 38469 43887
rect 38435 43789 38469 43819
rect 38435 43717 38469 43751
rect 38435 43663 38469 43683
rect 38893 44941 38927 44961
rect 38893 44873 38927 44907
rect 38893 44805 38927 44835
rect 38893 44737 38927 44763
rect 38893 44669 38927 44691
rect 38893 44601 38927 44619
rect 38893 44533 38927 44547
rect 38893 44465 38927 44475
rect 38893 44397 38927 44403
rect 38893 44329 38927 44331
rect 38893 44293 38927 44295
rect 38893 44221 38927 44227
rect 38893 44149 38927 44159
rect 38893 44077 38927 44091
rect 38893 44005 38927 44023
rect 38893 43933 38927 43955
rect 38893 43861 38927 43887
rect 38893 43789 38927 43819
rect 38893 43717 38927 43751
rect 38893 43582 38927 43683
rect 39351 44941 39385 45002
rect 39351 44873 39385 44907
rect 39351 44805 39385 44835
rect 39351 44737 39385 44763
rect 39351 44669 39385 44691
rect 39351 44601 39385 44619
rect 39351 44533 39385 44547
rect 39351 44465 39385 44475
rect 39351 44397 39385 44403
rect 39351 44329 39385 44331
rect 39351 44293 39385 44295
rect 39351 44221 39385 44227
rect 39351 44149 39385 44159
rect 39351 44077 39385 44091
rect 39351 44005 39385 44023
rect 39351 43933 39385 43955
rect 39351 43861 39385 43887
rect 39351 43789 39385 43819
rect 39351 43717 39385 43751
rect 39351 43663 39385 43683
rect 39809 44941 39843 44961
rect 39809 44873 39843 44907
rect 39809 44805 39843 44835
rect 39809 44737 39843 44763
rect 39809 44669 39843 44691
rect 39809 44601 39843 44619
rect 39809 44533 39843 44547
rect 39809 44465 39843 44475
rect 39809 44397 39843 44403
rect 39809 44329 39843 44331
rect 39809 44293 39843 44295
rect 39809 44221 39843 44227
rect 39809 44149 39843 44159
rect 39809 44077 39843 44091
rect 39809 44005 39843 44023
rect 39809 43933 39843 43955
rect 39809 43861 39843 43887
rect 39809 43789 39843 43819
rect 39809 43717 39843 43751
rect 39809 43582 39843 43683
rect 40267 44941 40301 45002
rect 40267 44873 40301 44907
rect 40267 44805 40301 44835
rect 40267 44737 40301 44763
rect 40267 44669 40301 44691
rect 40267 44601 40301 44619
rect 40267 44533 40301 44547
rect 40267 44465 40301 44475
rect 40267 44397 40301 44403
rect 40267 44329 40301 44331
rect 40267 44293 40301 44295
rect 40267 44221 40301 44227
rect 40267 44149 40301 44159
rect 40267 44077 40301 44091
rect 40267 44005 40301 44023
rect 40267 43933 40301 43955
rect 40267 43861 40301 43887
rect 40267 43789 40301 43819
rect 40267 43717 40301 43751
rect 40267 43663 40301 43683
rect 40725 44941 40759 44961
rect 40725 44873 40759 44907
rect 40725 44805 40759 44835
rect 40725 44737 40759 44763
rect 40725 44669 40759 44691
rect 40725 44601 40759 44619
rect 40725 44533 40759 44547
rect 40725 44465 40759 44475
rect 40725 44397 40759 44403
rect 40725 44329 40759 44331
rect 40725 44293 40759 44295
rect 40725 44221 40759 44227
rect 40725 44149 40759 44159
rect 40725 44077 40759 44091
rect 40725 44005 40759 44023
rect 40725 43933 40759 43955
rect 40725 43861 40759 43887
rect 40725 43789 40759 43819
rect 40725 43717 40759 43751
rect 40725 43582 40759 43683
rect 41183 44941 41217 45002
rect 41183 44873 41217 44907
rect 41183 44805 41217 44835
rect 41183 44737 41217 44763
rect 41183 44669 41217 44691
rect 41183 44601 41217 44619
rect 41183 44533 41217 44547
rect 41183 44465 41217 44475
rect 41183 44397 41217 44403
rect 41183 44329 41217 44331
rect 41183 44293 41217 44295
rect 41183 44221 41217 44227
rect 41183 44149 41217 44159
rect 41183 44077 41217 44091
rect 41183 44005 41217 44023
rect 41183 43933 41217 43955
rect 41183 43861 41217 43887
rect 41183 43789 41217 43819
rect 41183 43717 41217 43751
rect 41183 43663 41217 43683
rect 41641 44941 41675 44961
rect 41641 44873 41675 44907
rect 41641 44805 41675 44835
rect 41641 44737 41675 44763
rect 41641 44669 41675 44691
rect 41641 44601 41675 44619
rect 41641 44533 41675 44547
rect 41641 44465 41675 44475
rect 41641 44397 41675 44403
rect 41641 44329 41675 44331
rect 41641 44293 41675 44295
rect 41641 44221 41675 44227
rect 41641 44149 41675 44159
rect 41641 44077 41675 44091
rect 41641 44005 41675 44023
rect 41641 43933 41675 43955
rect 41641 43861 41675 43887
rect 41641 43789 41675 43819
rect 41641 43717 41675 43751
rect 41641 43582 41675 43683
rect 42099 44941 42133 45002
rect 42099 44873 42133 44907
rect 42099 44805 42133 44835
rect 42099 44737 42133 44763
rect 42099 44669 42133 44691
rect 42099 44601 42133 44619
rect 42099 44533 42133 44547
rect 42099 44465 42133 44475
rect 42099 44397 42133 44403
rect 42099 44329 42133 44331
rect 42099 44293 42133 44295
rect 42099 44221 42133 44227
rect 42099 44149 42133 44159
rect 42099 44077 42133 44091
rect 42099 44005 42133 44023
rect 42099 43933 42133 43955
rect 42099 43861 42133 43887
rect 42099 43789 42133 43819
rect 42099 43717 42133 43751
rect 42099 43663 42133 43683
rect 42557 44941 42591 44961
rect 42557 44873 42591 44907
rect 42557 44805 42591 44835
rect 42557 44737 42591 44763
rect 42557 44669 42591 44691
rect 42557 44601 42591 44619
rect 42557 44533 42591 44547
rect 42557 44465 42591 44475
rect 42557 44397 42591 44403
rect 42557 44329 42591 44331
rect 42557 44293 42591 44295
rect 42557 44221 42591 44227
rect 42557 44149 42591 44159
rect 42557 44077 42591 44091
rect 42557 44005 42591 44023
rect 42557 43933 42591 43955
rect 42557 43861 42591 43887
rect 42557 43789 42591 43819
rect 42557 43717 42591 43751
rect 42557 43582 42591 43683
rect 42986 44876 52314 44896
rect 42986 44842 43006 44876
rect 43040 44842 43096 44876
rect 43130 44861 43186 44876
rect 43220 44861 43276 44876
rect 43310 44861 43366 44876
rect 43400 44861 43456 44876
rect 43490 44861 43546 44876
rect 43580 44861 43636 44876
rect 43670 44861 43726 44876
rect 43760 44861 43816 44876
rect 43850 44861 43906 44876
rect 43940 44861 43996 44876
rect 44030 44861 44086 44876
rect 44120 44861 44176 44876
rect 43150 44842 43186 44861
rect 43240 44842 43276 44861
rect 43330 44842 43366 44861
rect 43420 44842 43456 44861
rect 43510 44842 43546 44861
rect 43600 44842 43636 44861
rect 43690 44842 43726 44861
rect 43780 44842 43816 44861
rect 43870 44842 43906 44861
rect 43960 44842 43996 44861
rect 44050 44842 44086 44861
rect 44140 44842 44176 44861
rect 44210 44842 44346 44876
rect 44380 44842 44436 44876
rect 44470 44861 44526 44876
rect 44560 44861 44616 44876
rect 44650 44861 44706 44876
rect 44740 44861 44796 44876
rect 44830 44861 44886 44876
rect 44920 44861 44976 44876
rect 45010 44861 45066 44876
rect 45100 44861 45156 44876
rect 45190 44861 45246 44876
rect 45280 44861 45336 44876
rect 45370 44861 45426 44876
rect 45460 44861 45516 44876
rect 44490 44842 44526 44861
rect 44580 44842 44616 44861
rect 44670 44842 44706 44861
rect 44760 44842 44796 44861
rect 44850 44842 44886 44861
rect 44940 44842 44976 44861
rect 45030 44842 45066 44861
rect 45120 44842 45156 44861
rect 45210 44842 45246 44861
rect 45300 44842 45336 44861
rect 45390 44842 45426 44861
rect 45480 44842 45516 44861
rect 45550 44842 45686 44876
rect 45720 44842 45776 44876
rect 45810 44861 45866 44876
rect 45900 44861 45956 44876
rect 45990 44861 46046 44876
rect 46080 44861 46136 44876
rect 46170 44861 46226 44876
rect 46260 44861 46316 44876
rect 46350 44861 46406 44876
rect 46440 44861 46496 44876
rect 46530 44861 46586 44876
rect 46620 44861 46676 44876
rect 46710 44861 46766 44876
rect 46800 44861 46856 44876
rect 45830 44842 45866 44861
rect 45920 44842 45956 44861
rect 46010 44842 46046 44861
rect 46100 44842 46136 44861
rect 46190 44842 46226 44861
rect 46280 44842 46316 44861
rect 46370 44842 46406 44861
rect 46460 44842 46496 44861
rect 46550 44842 46586 44861
rect 46640 44842 46676 44861
rect 46730 44842 46766 44861
rect 46820 44842 46856 44861
rect 46890 44842 47026 44876
rect 47060 44842 47116 44876
rect 47150 44861 47206 44876
rect 47240 44861 47296 44876
rect 47330 44861 47386 44876
rect 47420 44861 47476 44876
rect 47510 44861 47566 44876
rect 47600 44861 47656 44876
rect 47690 44861 47746 44876
rect 47780 44861 47836 44876
rect 47870 44861 47926 44876
rect 47960 44861 48016 44876
rect 48050 44861 48106 44876
rect 48140 44861 48196 44876
rect 47170 44842 47206 44861
rect 47260 44842 47296 44861
rect 47350 44842 47386 44861
rect 47440 44842 47476 44861
rect 47530 44842 47566 44861
rect 47620 44842 47656 44861
rect 47710 44842 47746 44861
rect 47800 44842 47836 44861
rect 47890 44842 47926 44861
rect 47980 44842 48016 44861
rect 48070 44842 48106 44861
rect 48160 44842 48196 44861
rect 48230 44842 48366 44876
rect 48400 44842 48456 44876
rect 48490 44861 48546 44876
rect 48580 44861 48636 44876
rect 48670 44861 48726 44876
rect 48760 44861 48816 44876
rect 48850 44861 48906 44876
rect 48940 44861 48996 44876
rect 49030 44861 49086 44876
rect 49120 44861 49176 44876
rect 49210 44861 49266 44876
rect 49300 44861 49356 44876
rect 49390 44861 49446 44876
rect 49480 44861 49536 44876
rect 48510 44842 48546 44861
rect 48600 44842 48636 44861
rect 48690 44842 48726 44861
rect 48780 44842 48816 44861
rect 48870 44842 48906 44861
rect 48960 44842 48996 44861
rect 49050 44842 49086 44861
rect 49140 44842 49176 44861
rect 49230 44842 49266 44861
rect 49320 44842 49356 44861
rect 49410 44842 49446 44861
rect 49500 44842 49536 44861
rect 49570 44842 49706 44876
rect 49740 44842 49796 44876
rect 49830 44861 49886 44876
rect 49920 44861 49976 44876
rect 50010 44861 50066 44876
rect 50100 44861 50156 44876
rect 50190 44861 50246 44876
rect 50280 44861 50336 44876
rect 50370 44861 50426 44876
rect 50460 44861 50516 44876
rect 50550 44861 50606 44876
rect 50640 44861 50696 44876
rect 50730 44861 50786 44876
rect 50820 44861 50876 44876
rect 49850 44842 49886 44861
rect 49940 44842 49976 44861
rect 50030 44842 50066 44861
rect 50120 44842 50156 44861
rect 50210 44842 50246 44861
rect 50300 44842 50336 44861
rect 50390 44842 50426 44861
rect 50480 44842 50516 44861
rect 50570 44842 50606 44861
rect 50660 44842 50696 44861
rect 50750 44842 50786 44861
rect 50840 44842 50876 44861
rect 50910 44842 51046 44876
rect 51080 44842 51136 44876
rect 51170 44861 51226 44876
rect 51260 44861 51316 44876
rect 51350 44861 51406 44876
rect 51440 44861 51496 44876
rect 51530 44861 51586 44876
rect 51620 44861 51676 44876
rect 51710 44861 51766 44876
rect 51800 44861 51856 44876
rect 51890 44861 51946 44876
rect 51980 44861 52036 44876
rect 52070 44861 52126 44876
rect 52160 44861 52216 44876
rect 51190 44842 51226 44861
rect 51280 44842 51316 44861
rect 51370 44842 51406 44861
rect 51460 44842 51496 44861
rect 51550 44842 51586 44861
rect 51640 44842 51676 44861
rect 51730 44842 51766 44861
rect 51820 44842 51856 44861
rect 51910 44842 51946 44861
rect 52000 44842 52036 44861
rect 52090 44842 52126 44861
rect 52180 44842 52216 44861
rect 52250 44842 52314 44876
rect 42986 44838 43116 44842
rect 42986 44804 43020 44838
rect 43054 44827 43116 44838
rect 43150 44827 43206 44842
rect 43240 44827 43296 44842
rect 43330 44827 43386 44842
rect 43420 44827 43476 44842
rect 43510 44827 43566 44842
rect 43600 44827 43656 44842
rect 43690 44827 43746 44842
rect 43780 44827 43836 44842
rect 43870 44827 43926 44842
rect 43960 44827 44016 44842
rect 44050 44827 44106 44842
rect 44140 44838 44456 44842
rect 44140 44827 44207 44838
rect 43054 44804 44207 44827
rect 44241 44804 44360 44838
rect 44394 44827 44456 44838
rect 44490 44827 44546 44842
rect 44580 44827 44636 44842
rect 44670 44827 44726 44842
rect 44760 44827 44816 44842
rect 44850 44827 44906 44842
rect 44940 44827 44996 44842
rect 45030 44827 45086 44842
rect 45120 44827 45176 44842
rect 45210 44827 45266 44842
rect 45300 44827 45356 44842
rect 45390 44827 45446 44842
rect 45480 44838 45796 44842
rect 45480 44827 45547 44838
rect 44394 44804 45547 44827
rect 45581 44804 45700 44838
rect 45734 44827 45796 44838
rect 45830 44827 45886 44842
rect 45920 44827 45976 44842
rect 46010 44827 46066 44842
rect 46100 44827 46156 44842
rect 46190 44827 46246 44842
rect 46280 44827 46336 44842
rect 46370 44827 46426 44842
rect 46460 44827 46516 44842
rect 46550 44827 46606 44842
rect 46640 44827 46696 44842
rect 46730 44827 46786 44842
rect 46820 44838 47136 44842
rect 46820 44827 46887 44838
rect 45734 44804 46887 44827
rect 46921 44804 47040 44838
rect 47074 44827 47136 44838
rect 47170 44827 47226 44842
rect 47260 44827 47316 44842
rect 47350 44827 47406 44842
rect 47440 44827 47496 44842
rect 47530 44827 47586 44842
rect 47620 44827 47676 44842
rect 47710 44827 47766 44842
rect 47800 44827 47856 44842
rect 47890 44827 47946 44842
rect 47980 44827 48036 44842
rect 48070 44827 48126 44842
rect 48160 44838 48476 44842
rect 48160 44827 48227 44838
rect 47074 44804 48227 44827
rect 48261 44804 48380 44838
rect 48414 44827 48476 44838
rect 48510 44827 48566 44842
rect 48600 44827 48656 44842
rect 48690 44827 48746 44842
rect 48780 44827 48836 44842
rect 48870 44827 48926 44842
rect 48960 44827 49016 44842
rect 49050 44827 49106 44842
rect 49140 44827 49196 44842
rect 49230 44827 49286 44842
rect 49320 44827 49376 44842
rect 49410 44827 49466 44842
rect 49500 44838 49816 44842
rect 49500 44827 49567 44838
rect 48414 44804 49567 44827
rect 49601 44804 49720 44838
rect 49754 44827 49816 44838
rect 49850 44827 49906 44842
rect 49940 44827 49996 44842
rect 50030 44827 50086 44842
rect 50120 44827 50176 44842
rect 50210 44827 50266 44842
rect 50300 44827 50356 44842
rect 50390 44827 50446 44842
rect 50480 44827 50536 44842
rect 50570 44827 50626 44842
rect 50660 44827 50716 44842
rect 50750 44827 50806 44842
rect 50840 44838 51156 44842
rect 50840 44827 50907 44838
rect 49754 44804 50907 44827
rect 50941 44804 51060 44838
rect 51094 44827 51156 44838
rect 51190 44827 51246 44842
rect 51280 44827 51336 44842
rect 51370 44827 51426 44842
rect 51460 44827 51516 44842
rect 51550 44827 51606 44842
rect 51640 44827 51696 44842
rect 51730 44827 51786 44842
rect 51820 44827 51876 44842
rect 51910 44827 51966 44842
rect 52000 44827 52056 44842
rect 52090 44827 52146 44842
rect 52180 44838 52314 44842
rect 52180 44827 52247 44838
rect 51094 44804 52247 44827
rect 52281 44804 52314 44838
rect 42986 44797 52314 44804
rect 42986 44748 43085 44797
rect 42986 44714 43020 44748
rect 43054 44714 43085 44748
rect 44175 44748 44425 44797
rect 42986 44658 43085 44714
rect 42986 44624 43020 44658
rect 43054 44624 43085 44658
rect 42986 44568 43085 44624
rect 42986 44534 43020 44568
rect 43054 44534 43085 44568
rect 42986 44478 43085 44534
rect 42986 44444 43020 44478
rect 43054 44444 43085 44478
rect 42986 44388 43085 44444
rect 42986 44354 43020 44388
rect 43054 44354 43085 44388
rect 42986 44298 43085 44354
rect 42986 44264 43020 44298
rect 43054 44264 43085 44298
rect 42986 44208 43085 44264
rect 42986 44174 43020 44208
rect 43054 44174 43085 44208
rect 42986 44118 43085 44174
rect 42986 44084 43020 44118
rect 43054 44084 43085 44118
rect 42986 44028 43085 44084
rect 42986 43994 43020 44028
rect 43054 43994 43085 44028
rect 42986 43938 43085 43994
rect 42986 43904 43020 43938
rect 43054 43904 43085 43938
rect 42986 43848 43085 43904
rect 42986 43814 43020 43848
rect 43054 43814 43085 43848
rect 42986 43758 43085 43814
rect 43149 44716 44111 44733
rect 43149 44682 43170 44716
rect 43204 44682 43260 44716
rect 43294 44714 43350 44716
rect 43384 44714 43440 44716
rect 43474 44714 43530 44716
rect 43564 44714 43620 44716
rect 43654 44714 43710 44716
rect 43744 44714 43800 44716
rect 43834 44714 43890 44716
rect 43924 44714 43980 44716
rect 44014 44714 44070 44716
rect 43314 44682 43350 44714
rect 43404 44682 43440 44714
rect 43494 44682 43530 44714
rect 43584 44682 43620 44714
rect 43674 44682 43710 44714
rect 43764 44682 43800 44714
rect 43854 44682 43890 44714
rect 43944 44682 43980 44714
rect 44034 44682 44070 44714
rect 44104 44682 44111 44716
rect 43149 44680 43280 44682
rect 43314 44680 43370 44682
rect 43404 44680 43460 44682
rect 43494 44680 43550 44682
rect 43584 44680 43640 44682
rect 43674 44680 43730 44682
rect 43764 44680 43820 44682
rect 43854 44680 43910 44682
rect 43944 44680 44000 44682
rect 44034 44680 44111 44682
rect 43149 44661 44111 44680
rect 43149 44657 43221 44661
rect 43149 44623 43168 44657
rect 43202 44623 43221 44657
rect 43149 44567 43221 44623
rect 44039 44638 44111 44661
rect 44039 44604 44058 44638
rect 44092 44604 44111 44638
rect 43149 44533 43168 44567
rect 43202 44533 43221 44567
rect 43149 44477 43221 44533
rect 43149 44443 43168 44477
rect 43202 44443 43221 44477
rect 43149 44387 43221 44443
rect 43149 44353 43168 44387
rect 43202 44353 43221 44387
rect 43149 44297 43221 44353
rect 43149 44263 43168 44297
rect 43202 44263 43221 44297
rect 43149 44207 43221 44263
rect 43149 44173 43168 44207
rect 43202 44173 43221 44207
rect 43149 44117 43221 44173
rect 43149 44083 43168 44117
rect 43202 44083 43221 44117
rect 43149 44027 43221 44083
rect 43149 43993 43168 44027
rect 43202 43993 43221 44027
rect 43149 43937 43221 43993
rect 43149 43903 43168 43937
rect 43202 43903 43221 43937
rect 43283 44540 43977 44599
rect 43283 44506 43344 44540
rect 43378 44512 43434 44540
rect 43468 44512 43524 44540
rect 43558 44512 43614 44540
rect 43390 44506 43434 44512
rect 43490 44506 43524 44512
rect 43590 44506 43614 44512
rect 43648 44512 43704 44540
rect 43648 44506 43656 44512
rect 43283 44478 43356 44506
rect 43390 44478 43456 44506
rect 43490 44478 43556 44506
rect 43590 44478 43656 44506
rect 43690 44506 43704 44512
rect 43738 44512 43794 44540
rect 43738 44506 43756 44512
rect 43690 44478 43756 44506
rect 43790 44506 43794 44512
rect 43828 44512 43884 44540
rect 43828 44506 43856 44512
rect 43918 44506 43977 44540
rect 43790 44478 43856 44506
rect 43890 44478 43977 44506
rect 43283 44450 43977 44478
rect 43283 44416 43344 44450
rect 43378 44416 43434 44450
rect 43468 44416 43524 44450
rect 43558 44416 43614 44450
rect 43648 44416 43704 44450
rect 43738 44416 43794 44450
rect 43828 44416 43884 44450
rect 43918 44416 43977 44450
rect 43283 44412 43977 44416
rect 43283 44378 43356 44412
rect 43390 44378 43456 44412
rect 43490 44378 43556 44412
rect 43590 44378 43656 44412
rect 43690 44378 43756 44412
rect 43790 44378 43856 44412
rect 43890 44378 43977 44412
rect 43283 44360 43977 44378
rect 43283 44326 43344 44360
rect 43378 44326 43434 44360
rect 43468 44326 43524 44360
rect 43558 44326 43614 44360
rect 43648 44326 43704 44360
rect 43738 44326 43794 44360
rect 43828 44326 43884 44360
rect 43918 44326 43977 44360
rect 43283 44312 43977 44326
rect 43283 44278 43356 44312
rect 43390 44278 43456 44312
rect 43490 44278 43556 44312
rect 43590 44278 43656 44312
rect 43690 44278 43756 44312
rect 43790 44278 43856 44312
rect 43890 44278 43977 44312
rect 43283 44270 43977 44278
rect 43283 44236 43344 44270
rect 43378 44236 43434 44270
rect 43468 44236 43524 44270
rect 43558 44236 43614 44270
rect 43648 44236 43704 44270
rect 43738 44236 43794 44270
rect 43828 44236 43884 44270
rect 43918 44236 43977 44270
rect 43283 44212 43977 44236
rect 43283 44180 43356 44212
rect 43390 44180 43456 44212
rect 43490 44180 43556 44212
rect 43590 44180 43656 44212
rect 43283 44146 43344 44180
rect 43390 44178 43434 44180
rect 43490 44178 43524 44180
rect 43590 44178 43614 44180
rect 43378 44146 43434 44178
rect 43468 44146 43524 44178
rect 43558 44146 43614 44178
rect 43648 44178 43656 44180
rect 43690 44180 43756 44212
rect 43690 44178 43704 44180
rect 43648 44146 43704 44178
rect 43738 44178 43756 44180
rect 43790 44180 43856 44212
rect 43890 44180 43977 44212
rect 43790 44178 43794 44180
rect 43738 44146 43794 44178
rect 43828 44178 43856 44180
rect 43828 44146 43884 44178
rect 43918 44146 43977 44180
rect 43283 44112 43977 44146
rect 43283 44090 43356 44112
rect 43390 44090 43456 44112
rect 43490 44090 43556 44112
rect 43590 44090 43656 44112
rect 43283 44056 43344 44090
rect 43390 44078 43434 44090
rect 43490 44078 43524 44090
rect 43590 44078 43614 44090
rect 43378 44056 43434 44078
rect 43468 44056 43524 44078
rect 43558 44056 43614 44078
rect 43648 44078 43656 44090
rect 43690 44090 43756 44112
rect 43690 44078 43704 44090
rect 43648 44056 43704 44078
rect 43738 44078 43756 44090
rect 43790 44090 43856 44112
rect 43890 44090 43977 44112
rect 43790 44078 43794 44090
rect 43738 44056 43794 44078
rect 43828 44078 43856 44090
rect 43828 44056 43884 44078
rect 43918 44056 43977 44090
rect 43283 44012 43977 44056
rect 43283 44000 43356 44012
rect 43390 44000 43456 44012
rect 43490 44000 43556 44012
rect 43590 44000 43656 44012
rect 43283 43966 43344 44000
rect 43390 43978 43434 44000
rect 43490 43978 43524 44000
rect 43590 43978 43614 44000
rect 43378 43966 43434 43978
rect 43468 43966 43524 43978
rect 43558 43966 43614 43978
rect 43648 43978 43656 44000
rect 43690 44000 43756 44012
rect 43690 43978 43704 44000
rect 43648 43966 43704 43978
rect 43738 43978 43756 44000
rect 43790 44000 43856 44012
rect 43890 44000 43977 44012
rect 43790 43978 43794 44000
rect 43738 43966 43794 43978
rect 43828 43978 43856 44000
rect 43828 43966 43884 43978
rect 43918 43966 43977 44000
rect 43283 43905 43977 43966
rect 44039 44548 44111 44604
rect 44039 44514 44058 44548
rect 44092 44514 44111 44548
rect 44039 44458 44111 44514
rect 44039 44424 44058 44458
rect 44092 44424 44111 44458
rect 44039 44368 44111 44424
rect 44039 44334 44058 44368
rect 44092 44334 44111 44368
rect 44039 44278 44111 44334
rect 44039 44244 44058 44278
rect 44092 44244 44111 44278
rect 44039 44188 44111 44244
rect 44039 44154 44058 44188
rect 44092 44154 44111 44188
rect 44039 44098 44111 44154
rect 44039 44064 44058 44098
rect 44092 44064 44111 44098
rect 44039 44008 44111 44064
rect 44039 43974 44058 44008
rect 44092 43974 44111 44008
rect 44039 43918 44111 43974
rect 43149 43843 43221 43903
rect 44039 43884 44058 43918
rect 44092 43884 44111 43918
rect 44039 43843 44111 43884
rect 43149 43824 44111 43843
rect 43149 43790 43246 43824
rect 43280 43790 43336 43824
rect 43370 43790 43426 43824
rect 43460 43790 43516 43824
rect 43550 43790 43606 43824
rect 43640 43790 43696 43824
rect 43730 43790 43786 43824
rect 43820 43790 43876 43824
rect 43910 43790 43966 43824
rect 44000 43790 44111 43824
rect 43149 43771 44111 43790
rect 44175 44714 44207 44748
rect 44241 44714 44360 44748
rect 44394 44714 44425 44748
rect 45515 44748 45765 44797
rect 44175 44658 44425 44714
rect 44175 44624 44207 44658
rect 44241 44624 44360 44658
rect 44394 44624 44425 44658
rect 44175 44568 44425 44624
rect 44175 44534 44207 44568
rect 44241 44534 44360 44568
rect 44394 44534 44425 44568
rect 44175 44478 44425 44534
rect 44175 44444 44207 44478
rect 44241 44444 44360 44478
rect 44394 44444 44425 44478
rect 44175 44388 44425 44444
rect 44175 44354 44207 44388
rect 44241 44354 44360 44388
rect 44394 44354 44425 44388
rect 44175 44298 44425 44354
rect 44175 44264 44207 44298
rect 44241 44264 44360 44298
rect 44394 44264 44425 44298
rect 44175 44208 44425 44264
rect 44175 44174 44207 44208
rect 44241 44174 44360 44208
rect 44394 44174 44425 44208
rect 44175 44118 44425 44174
rect 44175 44084 44207 44118
rect 44241 44084 44360 44118
rect 44394 44084 44425 44118
rect 44175 44028 44425 44084
rect 44175 43994 44207 44028
rect 44241 43994 44360 44028
rect 44394 43994 44425 44028
rect 44175 43938 44425 43994
rect 44175 43904 44207 43938
rect 44241 43904 44360 43938
rect 44394 43904 44425 43938
rect 44175 43848 44425 43904
rect 44175 43814 44207 43848
rect 44241 43814 44360 43848
rect 44394 43814 44425 43848
rect 42986 43724 43020 43758
rect 43054 43724 43085 43758
rect 42986 43707 43085 43724
rect 44175 43758 44425 43814
rect 44489 44716 45451 44733
rect 44489 44682 44510 44716
rect 44544 44682 44600 44716
rect 44634 44714 44690 44716
rect 44724 44714 44780 44716
rect 44814 44714 44870 44716
rect 44904 44714 44960 44716
rect 44994 44714 45050 44716
rect 45084 44714 45140 44716
rect 45174 44714 45230 44716
rect 45264 44714 45320 44716
rect 45354 44714 45410 44716
rect 44654 44682 44690 44714
rect 44744 44682 44780 44714
rect 44834 44682 44870 44714
rect 44924 44682 44960 44714
rect 45014 44682 45050 44714
rect 45104 44682 45140 44714
rect 45194 44682 45230 44714
rect 45284 44682 45320 44714
rect 45374 44682 45410 44714
rect 45444 44682 45451 44716
rect 44489 44680 44620 44682
rect 44654 44680 44710 44682
rect 44744 44680 44800 44682
rect 44834 44680 44890 44682
rect 44924 44680 44980 44682
rect 45014 44680 45070 44682
rect 45104 44680 45160 44682
rect 45194 44680 45250 44682
rect 45284 44680 45340 44682
rect 45374 44680 45451 44682
rect 44489 44661 45451 44680
rect 44489 44657 44561 44661
rect 44489 44623 44508 44657
rect 44542 44623 44561 44657
rect 44489 44567 44561 44623
rect 45379 44638 45451 44661
rect 45379 44604 45398 44638
rect 45432 44604 45451 44638
rect 44489 44533 44508 44567
rect 44542 44533 44561 44567
rect 44489 44477 44561 44533
rect 44489 44443 44508 44477
rect 44542 44443 44561 44477
rect 44489 44387 44561 44443
rect 44489 44353 44508 44387
rect 44542 44353 44561 44387
rect 44489 44297 44561 44353
rect 44489 44263 44508 44297
rect 44542 44263 44561 44297
rect 44489 44207 44561 44263
rect 44489 44173 44508 44207
rect 44542 44173 44561 44207
rect 44489 44117 44561 44173
rect 44489 44083 44508 44117
rect 44542 44083 44561 44117
rect 44489 44027 44561 44083
rect 44489 43993 44508 44027
rect 44542 43993 44561 44027
rect 44489 43937 44561 43993
rect 44489 43903 44508 43937
rect 44542 43903 44561 43937
rect 44623 44540 45317 44599
rect 44623 44506 44684 44540
rect 44718 44512 44774 44540
rect 44808 44512 44864 44540
rect 44898 44512 44954 44540
rect 44730 44506 44774 44512
rect 44830 44506 44864 44512
rect 44930 44506 44954 44512
rect 44988 44512 45044 44540
rect 44988 44506 44996 44512
rect 44623 44478 44696 44506
rect 44730 44478 44796 44506
rect 44830 44478 44896 44506
rect 44930 44478 44996 44506
rect 45030 44506 45044 44512
rect 45078 44512 45134 44540
rect 45078 44506 45096 44512
rect 45030 44478 45096 44506
rect 45130 44506 45134 44512
rect 45168 44512 45224 44540
rect 45168 44506 45196 44512
rect 45258 44506 45317 44540
rect 45130 44478 45196 44506
rect 45230 44478 45317 44506
rect 44623 44450 45317 44478
rect 44623 44416 44684 44450
rect 44718 44416 44774 44450
rect 44808 44416 44864 44450
rect 44898 44416 44954 44450
rect 44988 44416 45044 44450
rect 45078 44416 45134 44450
rect 45168 44416 45224 44450
rect 45258 44416 45317 44450
rect 44623 44412 45317 44416
rect 44623 44378 44696 44412
rect 44730 44378 44796 44412
rect 44830 44378 44896 44412
rect 44930 44378 44996 44412
rect 45030 44378 45096 44412
rect 45130 44378 45196 44412
rect 45230 44378 45317 44412
rect 44623 44360 45317 44378
rect 44623 44326 44684 44360
rect 44718 44326 44774 44360
rect 44808 44326 44864 44360
rect 44898 44326 44954 44360
rect 44988 44326 45044 44360
rect 45078 44326 45134 44360
rect 45168 44326 45224 44360
rect 45258 44326 45317 44360
rect 44623 44312 45317 44326
rect 44623 44278 44696 44312
rect 44730 44278 44796 44312
rect 44830 44278 44896 44312
rect 44930 44278 44996 44312
rect 45030 44278 45096 44312
rect 45130 44278 45196 44312
rect 45230 44278 45317 44312
rect 44623 44270 45317 44278
rect 44623 44236 44684 44270
rect 44718 44236 44774 44270
rect 44808 44236 44864 44270
rect 44898 44236 44954 44270
rect 44988 44236 45044 44270
rect 45078 44236 45134 44270
rect 45168 44236 45224 44270
rect 45258 44236 45317 44270
rect 44623 44212 45317 44236
rect 44623 44180 44696 44212
rect 44730 44180 44796 44212
rect 44830 44180 44896 44212
rect 44930 44180 44996 44212
rect 44623 44146 44684 44180
rect 44730 44178 44774 44180
rect 44830 44178 44864 44180
rect 44930 44178 44954 44180
rect 44718 44146 44774 44178
rect 44808 44146 44864 44178
rect 44898 44146 44954 44178
rect 44988 44178 44996 44180
rect 45030 44180 45096 44212
rect 45030 44178 45044 44180
rect 44988 44146 45044 44178
rect 45078 44178 45096 44180
rect 45130 44180 45196 44212
rect 45230 44180 45317 44212
rect 45130 44178 45134 44180
rect 45078 44146 45134 44178
rect 45168 44178 45196 44180
rect 45168 44146 45224 44178
rect 45258 44146 45317 44180
rect 44623 44112 45317 44146
rect 44623 44090 44696 44112
rect 44730 44090 44796 44112
rect 44830 44090 44896 44112
rect 44930 44090 44996 44112
rect 44623 44056 44684 44090
rect 44730 44078 44774 44090
rect 44830 44078 44864 44090
rect 44930 44078 44954 44090
rect 44718 44056 44774 44078
rect 44808 44056 44864 44078
rect 44898 44056 44954 44078
rect 44988 44078 44996 44090
rect 45030 44090 45096 44112
rect 45030 44078 45044 44090
rect 44988 44056 45044 44078
rect 45078 44078 45096 44090
rect 45130 44090 45196 44112
rect 45230 44090 45317 44112
rect 45130 44078 45134 44090
rect 45078 44056 45134 44078
rect 45168 44078 45196 44090
rect 45168 44056 45224 44078
rect 45258 44056 45317 44090
rect 44623 44012 45317 44056
rect 44623 44000 44696 44012
rect 44730 44000 44796 44012
rect 44830 44000 44896 44012
rect 44930 44000 44996 44012
rect 44623 43966 44684 44000
rect 44730 43978 44774 44000
rect 44830 43978 44864 44000
rect 44930 43978 44954 44000
rect 44718 43966 44774 43978
rect 44808 43966 44864 43978
rect 44898 43966 44954 43978
rect 44988 43978 44996 44000
rect 45030 44000 45096 44012
rect 45030 43978 45044 44000
rect 44988 43966 45044 43978
rect 45078 43978 45096 44000
rect 45130 44000 45196 44012
rect 45230 44000 45317 44012
rect 45130 43978 45134 44000
rect 45078 43966 45134 43978
rect 45168 43978 45196 44000
rect 45168 43966 45224 43978
rect 45258 43966 45317 44000
rect 44623 43905 45317 43966
rect 45379 44548 45451 44604
rect 45379 44514 45398 44548
rect 45432 44514 45451 44548
rect 45379 44458 45451 44514
rect 45379 44424 45398 44458
rect 45432 44424 45451 44458
rect 45379 44368 45451 44424
rect 45379 44334 45398 44368
rect 45432 44334 45451 44368
rect 45379 44278 45451 44334
rect 45379 44244 45398 44278
rect 45432 44244 45451 44278
rect 45379 44188 45451 44244
rect 45379 44154 45398 44188
rect 45432 44154 45451 44188
rect 45379 44098 45451 44154
rect 45379 44064 45398 44098
rect 45432 44064 45451 44098
rect 45379 44008 45451 44064
rect 45379 43974 45398 44008
rect 45432 43974 45451 44008
rect 45379 43918 45451 43974
rect 44489 43843 44561 43903
rect 45379 43884 45398 43918
rect 45432 43884 45451 43918
rect 45379 43843 45451 43884
rect 44489 43824 45451 43843
rect 44489 43790 44586 43824
rect 44620 43790 44676 43824
rect 44710 43790 44766 43824
rect 44800 43790 44856 43824
rect 44890 43790 44946 43824
rect 44980 43790 45036 43824
rect 45070 43790 45126 43824
rect 45160 43790 45216 43824
rect 45250 43790 45306 43824
rect 45340 43790 45451 43824
rect 44489 43771 45451 43790
rect 45515 44714 45547 44748
rect 45581 44714 45700 44748
rect 45734 44714 45765 44748
rect 46855 44748 47105 44797
rect 45515 44658 45765 44714
rect 45515 44624 45547 44658
rect 45581 44624 45700 44658
rect 45734 44624 45765 44658
rect 45515 44568 45765 44624
rect 45515 44534 45547 44568
rect 45581 44534 45700 44568
rect 45734 44534 45765 44568
rect 45515 44478 45765 44534
rect 45515 44444 45547 44478
rect 45581 44444 45700 44478
rect 45734 44444 45765 44478
rect 45515 44388 45765 44444
rect 45515 44354 45547 44388
rect 45581 44354 45700 44388
rect 45734 44354 45765 44388
rect 45515 44298 45765 44354
rect 45515 44264 45547 44298
rect 45581 44264 45700 44298
rect 45734 44264 45765 44298
rect 45515 44208 45765 44264
rect 45515 44174 45547 44208
rect 45581 44174 45700 44208
rect 45734 44174 45765 44208
rect 45515 44118 45765 44174
rect 45515 44084 45547 44118
rect 45581 44084 45700 44118
rect 45734 44084 45765 44118
rect 45515 44028 45765 44084
rect 45515 43994 45547 44028
rect 45581 43994 45700 44028
rect 45734 43994 45765 44028
rect 45515 43938 45765 43994
rect 45515 43904 45547 43938
rect 45581 43904 45700 43938
rect 45734 43904 45765 43938
rect 45515 43848 45765 43904
rect 45515 43814 45547 43848
rect 45581 43814 45700 43848
rect 45734 43814 45765 43848
rect 44175 43724 44207 43758
rect 44241 43724 44360 43758
rect 44394 43724 44425 43758
rect 44175 43707 44425 43724
rect 45515 43758 45765 43814
rect 45829 44716 46791 44733
rect 45829 44682 45850 44716
rect 45884 44682 45940 44716
rect 45974 44714 46030 44716
rect 46064 44714 46120 44716
rect 46154 44714 46210 44716
rect 46244 44714 46300 44716
rect 46334 44714 46390 44716
rect 46424 44714 46480 44716
rect 46514 44714 46570 44716
rect 46604 44714 46660 44716
rect 46694 44714 46750 44716
rect 45994 44682 46030 44714
rect 46084 44682 46120 44714
rect 46174 44682 46210 44714
rect 46264 44682 46300 44714
rect 46354 44682 46390 44714
rect 46444 44682 46480 44714
rect 46534 44682 46570 44714
rect 46624 44682 46660 44714
rect 46714 44682 46750 44714
rect 46784 44682 46791 44716
rect 45829 44680 45960 44682
rect 45994 44680 46050 44682
rect 46084 44680 46140 44682
rect 46174 44680 46230 44682
rect 46264 44680 46320 44682
rect 46354 44680 46410 44682
rect 46444 44680 46500 44682
rect 46534 44680 46590 44682
rect 46624 44680 46680 44682
rect 46714 44680 46791 44682
rect 45829 44661 46791 44680
rect 45829 44657 45901 44661
rect 45829 44623 45848 44657
rect 45882 44623 45901 44657
rect 45829 44567 45901 44623
rect 46719 44638 46791 44661
rect 46719 44604 46738 44638
rect 46772 44604 46791 44638
rect 45829 44533 45848 44567
rect 45882 44533 45901 44567
rect 45829 44477 45901 44533
rect 45829 44443 45848 44477
rect 45882 44443 45901 44477
rect 45829 44387 45901 44443
rect 45829 44353 45848 44387
rect 45882 44353 45901 44387
rect 45829 44297 45901 44353
rect 45829 44263 45848 44297
rect 45882 44263 45901 44297
rect 45829 44207 45901 44263
rect 45829 44173 45848 44207
rect 45882 44173 45901 44207
rect 45829 44117 45901 44173
rect 45829 44083 45848 44117
rect 45882 44083 45901 44117
rect 45829 44027 45901 44083
rect 45829 43993 45848 44027
rect 45882 43993 45901 44027
rect 45829 43937 45901 43993
rect 45829 43903 45848 43937
rect 45882 43903 45901 43937
rect 45963 44540 46657 44599
rect 45963 44506 46024 44540
rect 46058 44512 46114 44540
rect 46148 44512 46204 44540
rect 46238 44512 46294 44540
rect 46070 44506 46114 44512
rect 46170 44506 46204 44512
rect 46270 44506 46294 44512
rect 46328 44512 46384 44540
rect 46328 44506 46336 44512
rect 45963 44478 46036 44506
rect 46070 44478 46136 44506
rect 46170 44478 46236 44506
rect 46270 44478 46336 44506
rect 46370 44506 46384 44512
rect 46418 44512 46474 44540
rect 46418 44506 46436 44512
rect 46370 44478 46436 44506
rect 46470 44506 46474 44512
rect 46508 44512 46564 44540
rect 46508 44506 46536 44512
rect 46598 44506 46657 44540
rect 46470 44478 46536 44506
rect 46570 44478 46657 44506
rect 45963 44450 46657 44478
rect 45963 44416 46024 44450
rect 46058 44416 46114 44450
rect 46148 44416 46204 44450
rect 46238 44416 46294 44450
rect 46328 44416 46384 44450
rect 46418 44416 46474 44450
rect 46508 44416 46564 44450
rect 46598 44416 46657 44450
rect 45963 44412 46657 44416
rect 45963 44378 46036 44412
rect 46070 44378 46136 44412
rect 46170 44378 46236 44412
rect 46270 44378 46336 44412
rect 46370 44378 46436 44412
rect 46470 44378 46536 44412
rect 46570 44378 46657 44412
rect 45963 44360 46657 44378
rect 45963 44326 46024 44360
rect 46058 44326 46114 44360
rect 46148 44326 46204 44360
rect 46238 44326 46294 44360
rect 46328 44326 46384 44360
rect 46418 44326 46474 44360
rect 46508 44326 46564 44360
rect 46598 44326 46657 44360
rect 45963 44312 46657 44326
rect 45963 44278 46036 44312
rect 46070 44278 46136 44312
rect 46170 44278 46236 44312
rect 46270 44278 46336 44312
rect 46370 44278 46436 44312
rect 46470 44278 46536 44312
rect 46570 44278 46657 44312
rect 45963 44270 46657 44278
rect 45963 44236 46024 44270
rect 46058 44236 46114 44270
rect 46148 44236 46204 44270
rect 46238 44236 46294 44270
rect 46328 44236 46384 44270
rect 46418 44236 46474 44270
rect 46508 44236 46564 44270
rect 46598 44236 46657 44270
rect 45963 44212 46657 44236
rect 45963 44180 46036 44212
rect 46070 44180 46136 44212
rect 46170 44180 46236 44212
rect 46270 44180 46336 44212
rect 45963 44146 46024 44180
rect 46070 44178 46114 44180
rect 46170 44178 46204 44180
rect 46270 44178 46294 44180
rect 46058 44146 46114 44178
rect 46148 44146 46204 44178
rect 46238 44146 46294 44178
rect 46328 44178 46336 44180
rect 46370 44180 46436 44212
rect 46370 44178 46384 44180
rect 46328 44146 46384 44178
rect 46418 44178 46436 44180
rect 46470 44180 46536 44212
rect 46570 44180 46657 44212
rect 46470 44178 46474 44180
rect 46418 44146 46474 44178
rect 46508 44178 46536 44180
rect 46508 44146 46564 44178
rect 46598 44146 46657 44180
rect 45963 44112 46657 44146
rect 45963 44090 46036 44112
rect 46070 44090 46136 44112
rect 46170 44090 46236 44112
rect 46270 44090 46336 44112
rect 45963 44056 46024 44090
rect 46070 44078 46114 44090
rect 46170 44078 46204 44090
rect 46270 44078 46294 44090
rect 46058 44056 46114 44078
rect 46148 44056 46204 44078
rect 46238 44056 46294 44078
rect 46328 44078 46336 44090
rect 46370 44090 46436 44112
rect 46370 44078 46384 44090
rect 46328 44056 46384 44078
rect 46418 44078 46436 44090
rect 46470 44090 46536 44112
rect 46570 44090 46657 44112
rect 46470 44078 46474 44090
rect 46418 44056 46474 44078
rect 46508 44078 46536 44090
rect 46508 44056 46564 44078
rect 46598 44056 46657 44090
rect 45963 44012 46657 44056
rect 45963 44000 46036 44012
rect 46070 44000 46136 44012
rect 46170 44000 46236 44012
rect 46270 44000 46336 44012
rect 45963 43966 46024 44000
rect 46070 43978 46114 44000
rect 46170 43978 46204 44000
rect 46270 43978 46294 44000
rect 46058 43966 46114 43978
rect 46148 43966 46204 43978
rect 46238 43966 46294 43978
rect 46328 43978 46336 44000
rect 46370 44000 46436 44012
rect 46370 43978 46384 44000
rect 46328 43966 46384 43978
rect 46418 43978 46436 44000
rect 46470 44000 46536 44012
rect 46570 44000 46657 44012
rect 46470 43978 46474 44000
rect 46418 43966 46474 43978
rect 46508 43978 46536 44000
rect 46508 43966 46564 43978
rect 46598 43966 46657 44000
rect 45963 43905 46657 43966
rect 46719 44548 46791 44604
rect 46719 44514 46738 44548
rect 46772 44514 46791 44548
rect 46719 44458 46791 44514
rect 46719 44424 46738 44458
rect 46772 44424 46791 44458
rect 46719 44368 46791 44424
rect 46719 44334 46738 44368
rect 46772 44334 46791 44368
rect 46719 44278 46791 44334
rect 46719 44244 46738 44278
rect 46772 44244 46791 44278
rect 46719 44188 46791 44244
rect 46719 44154 46738 44188
rect 46772 44154 46791 44188
rect 46719 44098 46791 44154
rect 46719 44064 46738 44098
rect 46772 44064 46791 44098
rect 46719 44008 46791 44064
rect 46719 43974 46738 44008
rect 46772 43974 46791 44008
rect 46719 43918 46791 43974
rect 45829 43843 45901 43903
rect 46719 43884 46738 43918
rect 46772 43884 46791 43918
rect 46719 43843 46791 43884
rect 45829 43824 46791 43843
rect 45829 43790 45926 43824
rect 45960 43790 46016 43824
rect 46050 43790 46106 43824
rect 46140 43790 46196 43824
rect 46230 43790 46286 43824
rect 46320 43790 46376 43824
rect 46410 43790 46466 43824
rect 46500 43790 46556 43824
rect 46590 43790 46646 43824
rect 46680 43790 46791 43824
rect 45829 43771 46791 43790
rect 46855 44714 46887 44748
rect 46921 44714 47040 44748
rect 47074 44714 47105 44748
rect 48195 44748 48445 44797
rect 46855 44658 47105 44714
rect 46855 44624 46887 44658
rect 46921 44624 47040 44658
rect 47074 44624 47105 44658
rect 46855 44568 47105 44624
rect 46855 44534 46887 44568
rect 46921 44534 47040 44568
rect 47074 44534 47105 44568
rect 46855 44478 47105 44534
rect 46855 44444 46887 44478
rect 46921 44444 47040 44478
rect 47074 44444 47105 44478
rect 46855 44388 47105 44444
rect 46855 44354 46887 44388
rect 46921 44354 47040 44388
rect 47074 44354 47105 44388
rect 46855 44298 47105 44354
rect 46855 44264 46887 44298
rect 46921 44264 47040 44298
rect 47074 44264 47105 44298
rect 46855 44208 47105 44264
rect 46855 44174 46887 44208
rect 46921 44174 47040 44208
rect 47074 44174 47105 44208
rect 46855 44118 47105 44174
rect 46855 44084 46887 44118
rect 46921 44084 47040 44118
rect 47074 44084 47105 44118
rect 46855 44028 47105 44084
rect 46855 43994 46887 44028
rect 46921 43994 47040 44028
rect 47074 43994 47105 44028
rect 46855 43938 47105 43994
rect 46855 43904 46887 43938
rect 46921 43904 47040 43938
rect 47074 43904 47105 43938
rect 46855 43848 47105 43904
rect 46855 43814 46887 43848
rect 46921 43814 47040 43848
rect 47074 43814 47105 43848
rect 45515 43724 45547 43758
rect 45581 43724 45700 43758
rect 45734 43724 45765 43758
rect 45515 43707 45765 43724
rect 46855 43758 47105 43814
rect 47169 44716 48131 44733
rect 47169 44682 47190 44716
rect 47224 44682 47280 44716
rect 47314 44714 47370 44716
rect 47404 44714 47460 44716
rect 47494 44714 47550 44716
rect 47584 44714 47640 44716
rect 47674 44714 47730 44716
rect 47764 44714 47820 44716
rect 47854 44714 47910 44716
rect 47944 44714 48000 44716
rect 48034 44714 48090 44716
rect 47334 44682 47370 44714
rect 47424 44682 47460 44714
rect 47514 44682 47550 44714
rect 47604 44682 47640 44714
rect 47694 44682 47730 44714
rect 47784 44682 47820 44714
rect 47874 44682 47910 44714
rect 47964 44682 48000 44714
rect 48054 44682 48090 44714
rect 48124 44682 48131 44716
rect 47169 44680 47300 44682
rect 47334 44680 47390 44682
rect 47424 44680 47480 44682
rect 47514 44680 47570 44682
rect 47604 44680 47660 44682
rect 47694 44680 47750 44682
rect 47784 44680 47840 44682
rect 47874 44680 47930 44682
rect 47964 44680 48020 44682
rect 48054 44680 48131 44682
rect 47169 44661 48131 44680
rect 47169 44657 47241 44661
rect 47169 44623 47188 44657
rect 47222 44623 47241 44657
rect 47169 44567 47241 44623
rect 48059 44638 48131 44661
rect 48059 44604 48078 44638
rect 48112 44604 48131 44638
rect 47169 44533 47188 44567
rect 47222 44533 47241 44567
rect 47169 44477 47241 44533
rect 47169 44443 47188 44477
rect 47222 44443 47241 44477
rect 47169 44387 47241 44443
rect 47169 44353 47188 44387
rect 47222 44353 47241 44387
rect 47169 44297 47241 44353
rect 47169 44263 47188 44297
rect 47222 44263 47241 44297
rect 47169 44207 47241 44263
rect 47169 44173 47188 44207
rect 47222 44173 47241 44207
rect 47169 44117 47241 44173
rect 47169 44083 47188 44117
rect 47222 44083 47241 44117
rect 47169 44027 47241 44083
rect 47169 43993 47188 44027
rect 47222 43993 47241 44027
rect 47169 43937 47241 43993
rect 47169 43903 47188 43937
rect 47222 43903 47241 43937
rect 47303 44540 47997 44599
rect 47303 44506 47364 44540
rect 47398 44512 47454 44540
rect 47488 44512 47544 44540
rect 47578 44512 47634 44540
rect 47410 44506 47454 44512
rect 47510 44506 47544 44512
rect 47610 44506 47634 44512
rect 47668 44512 47724 44540
rect 47668 44506 47676 44512
rect 47303 44478 47376 44506
rect 47410 44478 47476 44506
rect 47510 44478 47576 44506
rect 47610 44478 47676 44506
rect 47710 44506 47724 44512
rect 47758 44512 47814 44540
rect 47758 44506 47776 44512
rect 47710 44478 47776 44506
rect 47810 44506 47814 44512
rect 47848 44512 47904 44540
rect 47848 44506 47876 44512
rect 47938 44506 47997 44540
rect 47810 44478 47876 44506
rect 47910 44478 47997 44506
rect 47303 44450 47997 44478
rect 47303 44416 47364 44450
rect 47398 44416 47454 44450
rect 47488 44416 47544 44450
rect 47578 44416 47634 44450
rect 47668 44416 47724 44450
rect 47758 44416 47814 44450
rect 47848 44416 47904 44450
rect 47938 44416 47997 44450
rect 47303 44412 47997 44416
rect 47303 44378 47376 44412
rect 47410 44378 47476 44412
rect 47510 44378 47576 44412
rect 47610 44378 47676 44412
rect 47710 44378 47776 44412
rect 47810 44378 47876 44412
rect 47910 44378 47997 44412
rect 47303 44360 47997 44378
rect 47303 44326 47364 44360
rect 47398 44326 47454 44360
rect 47488 44326 47544 44360
rect 47578 44326 47634 44360
rect 47668 44326 47724 44360
rect 47758 44326 47814 44360
rect 47848 44326 47904 44360
rect 47938 44326 47997 44360
rect 47303 44312 47997 44326
rect 47303 44278 47376 44312
rect 47410 44278 47476 44312
rect 47510 44278 47576 44312
rect 47610 44278 47676 44312
rect 47710 44278 47776 44312
rect 47810 44278 47876 44312
rect 47910 44278 47997 44312
rect 47303 44270 47997 44278
rect 47303 44236 47364 44270
rect 47398 44236 47454 44270
rect 47488 44236 47544 44270
rect 47578 44236 47634 44270
rect 47668 44236 47724 44270
rect 47758 44236 47814 44270
rect 47848 44236 47904 44270
rect 47938 44236 47997 44270
rect 47303 44212 47997 44236
rect 47303 44180 47376 44212
rect 47410 44180 47476 44212
rect 47510 44180 47576 44212
rect 47610 44180 47676 44212
rect 47303 44146 47364 44180
rect 47410 44178 47454 44180
rect 47510 44178 47544 44180
rect 47610 44178 47634 44180
rect 47398 44146 47454 44178
rect 47488 44146 47544 44178
rect 47578 44146 47634 44178
rect 47668 44178 47676 44180
rect 47710 44180 47776 44212
rect 47710 44178 47724 44180
rect 47668 44146 47724 44178
rect 47758 44178 47776 44180
rect 47810 44180 47876 44212
rect 47910 44180 47997 44212
rect 47810 44178 47814 44180
rect 47758 44146 47814 44178
rect 47848 44178 47876 44180
rect 47848 44146 47904 44178
rect 47938 44146 47997 44180
rect 47303 44112 47997 44146
rect 47303 44090 47376 44112
rect 47410 44090 47476 44112
rect 47510 44090 47576 44112
rect 47610 44090 47676 44112
rect 47303 44056 47364 44090
rect 47410 44078 47454 44090
rect 47510 44078 47544 44090
rect 47610 44078 47634 44090
rect 47398 44056 47454 44078
rect 47488 44056 47544 44078
rect 47578 44056 47634 44078
rect 47668 44078 47676 44090
rect 47710 44090 47776 44112
rect 47710 44078 47724 44090
rect 47668 44056 47724 44078
rect 47758 44078 47776 44090
rect 47810 44090 47876 44112
rect 47910 44090 47997 44112
rect 47810 44078 47814 44090
rect 47758 44056 47814 44078
rect 47848 44078 47876 44090
rect 47848 44056 47904 44078
rect 47938 44056 47997 44090
rect 47303 44012 47997 44056
rect 47303 44000 47376 44012
rect 47410 44000 47476 44012
rect 47510 44000 47576 44012
rect 47610 44000 47676 44012
rect 47303 43966 47364 44000
rect 47410 43978 47454 44000
rect 47510 43978 47544 44000
rect 47610 43978 47634 44000
rect 47398 43966 47454 43978
rect 47488 43966 47544 43978
rect 47578 43966 47634 43978
rect 47668 43978 47676 44000
rect 47710 44000 47776 44012
rect 47710 43978 47724 44000
rect 47668 43966 47724 43978
rect 47758 43978 47776 44000
rect 47810 44000 47876 44012
rect 47910 44000 47997 44012
rect 47810 43978 47814 44000
rect 47758 43966 47814 43978
rect 47848 43978 47876 44000
rect 47848 43966 47904 43978
rect 47938 43966 47997 44000
rect 47303 43905 47997 43966
rect 48059 44548 48131 44604
rect 48059 44514 48078 44548
rect 48112 44514 48131 44548
rect 48059 44458 48131 44514
rect 48059 44424 48078 44458
rect 48112 44424 48131 44458
rect 48059 44368 48131 44424
rect 48059 44334 48078 44368
rect 48112 44334 48131 44368
rect 48059 44278 48131 44334
rect 48059 44244 48078 44278
rect 48112 44244 48131 44278
rect 48059 44188 48131 44244
rect 48059 44154 48078 44188
rect 48112 44154 48131 44188
rect 48059 44098 48131 44154
rect 48059 44064 48078 44098
rect 48112 44064 48131 44098
rect 48059 44008 48131 44064
rect 48059 43974 48078 44008
rect 48112 43974 48131 44008
rect 48059 43918 48131 43974
rect 47169 43843 47241 43903
rect 48059 43884 48078 43918
rect 48112 43884 48131 43918
rect 48059 43843 48131 43884
rect 47169 43824 48131 43843
rect 47169 43790 47266 43824
rect 47300 43790 47356 43824
rect 47390 43790 47446 43824
rect 47480 43790 47536 43824
rect 47570 43790 47626 43824
rect 47660 43790 47716 43824
rect 47750 43790 47806 43824
rect 47840 43790 47896 43824
rect 47930 43790 47986 43824
rect 48020 43790 48131 43824
rect 47169 43771 48131 43790
rect 48195 44714 48227 44748
rect 48261 44714 48380 44748
rect 48414 44714 48445 44748
rect 49535 44748 49785 44797
rect 48195 44658 48445 44714
rect 48195 44624 48227 44658
rect 48261 44624 48380 44658
rect 48414 44624 48445 44658
rect 48195 44568 48445 44624
rect 48195 44534 48227 44568
rect 48261 44534 48380 44568
rect 48414 44534 48445 44568
rect 48195 44478 48445 44534
rect 48195 44444 48227 44478
rect 48261 44444 48380 44478
rect 48414 44444 48445 44478
rect 48195 44388 48445 44444
rect 48195 44354 48227 44388
rect 48261 44354 48380 44388
rect 48414 44354 48445 44388
rect 48195 44298 48445 44354
rect 48195 44264 48227 44298
rect 48261 44264 48380 44298
rect 48414 44264 48445 44298
rect 48195 44208 48445 44264
rect 48195 44174 48227 44208
rect 48261 44174 48380 44208
rect 48414 44174 48445 44208
rect 48195 44118 48445 44174
rect 48195 44084 48227 44118
rect 48261 44084 48380 44118
rect 48414 44084 48445 44118
rect 48195 44028 48445 44084
rect 48195 43994 48227 44028
rect 48261 43994 48380 44028
rect 48414 43994 48445 44028
rect 48195 43938 48445 43994
rect 48195 43904 48227 43938
rect 48261 43904 48380 43938
rect 48414 43904 48445 43938
rect 48195 43848 48445 43904
rect 48195 43814 48227 43848
rect 48261 43814 48380 43848
rect 48414 43814 48445 43848
rect 46855 43724 46887 43758
rect 46921 43724 47040 43758
rect 47074 43724 47105 43758
rect 46855 43707 47105 43724
rect 48195 43758 48445 43814
rect 48509 44716 49471 44733
rect 48509 44682 48530 44716
rect 48564 44682 48620 44716
rect 48654 44714 48710 44716
rect 48744 44714 48800 44716
rect 48834 44714 48890 44716
rect 48924 44714 48980 44716
rect 49014 44714 49070 44716
rect 49104 44714 49160 44716
rect 49194 44714 49250 44716
rect 49284 44714 49340 44716
rect 49374 44714 49430 44716
rect 48674 44682 48710 44714
rect 48764 44682 48800 44714
rect 48854 44682 48890 44714
rect 48944 44682 48980 44714
rect 49034 44682 49070 44714
rect 49124 44682 49160 44714
rect 49214 44682 49250 44714
rect 49304 44682 49340 44714
rect 49394 44682 49430 44714
rect 49464 44682 49471 44716
rect 48509 44680 48640 44682
rect 48674 44680 48730 44682
rect 48764 44680 48820 44682
rect 48854 44680 48910 44682
rect 48944 44680 49000 44682
rect 49034 44680 49090 44682
rect 49124 44680 49180 44682
rect 49214 44680 49270 44682
rect 49304 44680 49360 44682
rect 49394 44680 49471 44682
rect 48509 44661 49471 44680
rect 48509 44657 48581 44661
rect 48509 44623 48528 44657
rect 48562 44623 48581 44657
rect 48509 44567 48581 44623
rect 49399 44638 49471 44661
rect 49399 44604 49418 44638
rect 49452 44604 49471 44638
rect 48509 44533 48528 44567
rect 48562 44533 48581 44567
rect 48509 44477 48581 44533
rect 48509 44443 48528 44477
rect 48562 44443 48581 44477
rect 48509 44387 48581 44443
rect 48509 44353 48528 44387
rect 48562 44353 48581 44387
rect 48509 44297 48581 44353
rect 48509 44263 48528 44297
rect 48562 44263 48581 44297
rect 48509 44207 48581 44263
rect 48509 44173 48528 44207
rect 48562 44173 48581 44207
rect 48509 44117 48581 44173
rect 48509 44083 48528 44117
rect 48562 44083 48581 44117
rect 48509 44027 48581 44083
rect 48509 43993 48528 44027
rect 48562 43993 48581 44027
rect 48509 43937 48581 43993
rect 48509 43903 48528 43937
rect 48562 43903 48581 43937
rect 48643 44540 49337 44599
rect 48643 44506 48704 44540
rect 48738 44512 48794 44540
rect 48828 44512 48884 44540
rect 48918 44512 48974 44540
rect 48750 44506 48794 44512
rect 48850 44506 48884 44512
rect 48950 44506 48974 44512
rect 49008 44512 49064 44540
rect 49008 44506 49016 44512
rect 48643 44478 48716 44506
rect 48750 44478 48816 44506
rect 48850 44478 48916 44506
rect 48950 44478 49016 44506
rect 49050 44506 49064 44512
rect 49098 44512 49154 44540
rect 49098 44506 49116 44512
rect 49050 44478 49116 44506
rect 49150 44506 49154 44512
rect 49188 44512 49244 44540
rect 49188 44506 49216 44512
rect 49278 44506 49337 44540
rect 49150 44478 49216 44506
rect 49250 44478 49337 44506
rect 48643 44450 49337 44478
rect 48643 44416 48704 44450
rect 48738 44416 48794 44450
rect 48828 44416 48884 44450
rect 48918 44416 48974 44450
rect 49008 44416 49064 44450
rect 49098 44416 49154 44450
rect 49188 44416 49244 44450
rect 49278 44416 49337 44450
rect 48643 44412 49337 44416
rect 48643 44378 48716 44412
rect 48750 44378 48816 44412
rect 48850 44378 48916 44412
rect 48950 44378 49016 44412
rect 49050 44378 49116 44412
rect 49150 44378 49216 44412
rect 49250 44378 49337 44412
rect 48643 44360 49337 44378
rect 48643 44326 48704 44360
rect 48738 44326 48794 44360
rect 48828 44326 48884 44360
rect 48918 44326 48974 44360
rect 49008 44326 49064 44360
rect 49098 44326 49154 44360
rect 49188 44326 49244 44360
rect 49278 44326 49337 44360
rect 48643 44312 49337 44326
rect 48643 44278 48716 44312
rect 48750 44278 48816 44312
rect 48850 44278 48916 44312
rect 48950 44278 49016 44312
rect 49050 44278 49116 44312
rect 49150 44278 49216 44312
rect 49250 44278 49337 44312
rect 48643 44270 49337 44278
rect 48643 44236 48704 44270
rect 48738 44236 48794 44270
rect 48828 44236 48884 44270
rect 48918 44236 48974 44270
rect 49008 44236 49064 44270
rect 49098 44236 49154 44270
rect 49188 44236 49244 44270
rect 49278 44236 49337 44270
rect 48643 44212 49337 44236
rect 48643 44180 48716 44212
rect 48750 44180 48816 44212
rect 48850 44180 48916 44212
rect 48950 44180 49016 44212
rect 48643 44146 48704 44180
rect 48750 44178 48794 44180
rect 48850 44178 48884 44180
rect 48950 44178 48974 44180
rect 48738 44146 48794 44178
rect 48828 44146 48884 44178
rect 48918 44146 48974 44178
rect 49008 44178 49016 44180
rect 49050 44180 49116 44212
rect 49050 44178 49064 44180
rect 49008 44146 49064 44178
rect 49098 44178 49116 44180
rect 49150 44180 49216 44212
rect 49250 44180 49337 44212
rect 49150 44178 49154 44180
rect 49098 44146 49154 44178
rect 49188 44178 49216 44180
rect 49188 44146 49244 44178
rect 49278 44146 49337 44180
rect 48643 44112 49337 44146
rect 48643 44090 48716 44112
rect 48750 44090 48816 44112
rect 48850 44090 48916 44112
rect 48950 44090 49016 44112
rect 48643 44056 48704 44090
rect 48750 44078 48794 44090
rect 48850 44078 48884 44090
rect 48950 44078 48974 44090
rect 48738 44056 48794 44078
rect 48828 44056 48884 44078
rect 48918 44056 48974 44078
rect 49008 44078 49016 44090
rect 49050 44090 49116 44112
rect 49050 44078 49064 44090
rect 49008 44056 49064 44078
rect 49098 44078 49116 44090
rect 49150 44090 49216 44112
rect 49250 44090 49337 44112
rect 49150 44078 49154 44090
rect 49098 44056 49154 44078
rect 49188 44078 49216 44090
rect 49188 44056 49244 44078
rect 49278 44056 49337 44090
rect 48643 44012 49337 44056
rect 48643 44000 48716 44012
rect 48750 44000 48816 44012
rect 48850 44000 48916 44012
rect 48950 44000 49016 44012
rect 48643 43966 48704 44000
rect 48750 43978 48794 44000
rect 48850 43978 48884 44000
rect 48950 43978 48974 44000
rect 48738 43966 48794 43978
rect 48828 43966 48884 43978
rect 48918 43966 48974 43978
rect 49008 43978 49016 44000
rect 49050 44000 49116 44012
rect 49050 43978 49064 44000
rect 49008 43966 49064 43978
rect 49098 43978 49116 44000
rect 49150 44000 49216 44012
rect 49250 44000 49337 44012
rect 49150 43978 49154 44000
rect 49098 43966 49154 43978
rect 49188 43978 49216 44000
rect 49188 43966 49244 43978
rect 49278 43966 49337 44000
rect 48643 43905 49337 43966
rect 49399 44548 49471 44604
rect 49399 44514 49418 44548
rect 49452 44514 49471 44548
rect 49399 44458 49471 44514
rect 49399 44424 49418 44458
rect 49452 44424 49471 44458
rect 49399 44368 49471 44424
rect 49399 44334 49418 44368
rect 49452 44334 49471 44368
rect 49399 44278 49471 44334
rect 49399 44244 49418 44278
rect 49452 44244 49471 44278
rect 49399 44188 49471 44244
rect 49399 44154 49418 44188
rect 49452 44154 49471 44188
rect 49399 44098 49471 44154
rect 49399 44064 49418 44098
rect 49452 44064 49471 44098
rect 49399 44008 49471 44064
rect 49399 43974 49418 44008
rect 49452 43974 49471 44008
rect 49399 43918 49471 43974
rect 48509 43843 48581 43903
rect 49399 43884 49418 43918
rect 49452 43884 49471 43918
rect 49399 43843 49471 43884
rect 48509 43824 49471 43843
rect 48509 43790 48606 43824
rect 48640 43790 48696 43824
rect 48730 43790 48786 43824
rect 48820 43790 48876 43824
rect 48910 43790 48966 43824
rect 49000 43790 49056 43824
rect 49090 43790 49146 43824
rect 49180 43790 49236 43824
rect 49270 43790 49326 43824
rect 49360 43790 49471 43824
rect 48509 43771 49471 43790
rect 49535 44714 49567 44748
rect 49601 44714 49720 44748
rect 49754 44714 49785 44748
rect 50875 44748 51125 44797
rect 49535 44658 49785 44714
rect 49535 44624 49567 44658
rect 49601 44624 49720 44658
rect 49754 44624 49785 44658
rect 49535 44568 49785 44624
rect 49535 44534 49567 44568
rect 49601 44534 49720 44568
rect 49754 44534 49785 44568
rect 49535 44478 49785 44534
rect 49535 44444 49567 44478
rect 49601 44444 49720 44478
rect 49754 44444 49785 44478
rect 49535 44388 49785 44444
rect 49535 44354 49567 44388
rect 49601 44354 49720 44388
rect 49754 44354 49785 44388
rect 49535 44298 49785 44354
rect 49535 44264 49567 44298
rect 49601 44264 49720 44298
rect 49754 44264 49785 44298
rect 49535 44208 49785 44264
rect 49535 44174 49567 44208
rect 49601 44174 49720 44208
rect 49754 44174 49785 44208
rect 49535 44118 49785 44174
rect 49535 44084 49567 44118
rect 49601 44084 49720 44118
rect 49754 44084 49785 44118
rect 49535 44028 49785 44084
rect 49535 43994 49567 44028
rect 49601 43994 49720 44028
rect 49754 43994 49785 44028
rect 49535 43938 49785 43994
rect 49535 43904 49567 43938
rect 49601 43904 49720 43938
rect 49754 43904 49785 43938
rect 49535 43848 49785 43904
rect 49535 43814 49567 43848
rect 49601 43814 49720 43848
rect 49754 43814 49785 43848
rect 48195 43724 48227 43758
rect 48261 43724 48380 43758
rect 48414 43724 48445 43758
rect 48195 43707 48445 43724
rect 49535 43758 49785 43814
rect 49849 44716 50811 44733
rect 49849 44682 49870 44716
rect 49904 44682 49960 44716
rect 49994 44714 50050 44716
rect 50084 44714 50140 44716
rect 50174 44714 50230 44716
rect 50264 44714 50320 44716
rect 50354 44714 50410 44716
rect 50444 44714 50500 44716
rect 50534 44714 50590 44716
rect 50624 44714 50680 44716
rect 50714 44714 50770 44716
rect 50014 44682 50050 44714
rect 50104 44682 50140 44714
rect 50194 44682 50230 44714
rect 50284 44682 50320 44714
rect 50374 44682 50410 44714
rect 50464 44682 50500 44714
rect 50554 44682 50590 44714
rect 50644 44682 50680 44714
rect 50734 44682 50770 44714
rect 50804 44682 50811 44716
rect 49849 44680 49980 44682
rect 50014 44680 50070 44682
rect 50104 44680 50160 44682
rect 50194 44680 50250 44682
rect 50284 44680 50340 44682
rect 50374 44680 50430 44682
rect 50464 44680 50520 44682
rect 50554 44680 50610 44682
rect 50644 44680 50700 44682
rect 50734 44680 50811 44682
rect 49849 44661 50811 44680
rect 49849 44657 49921 44661
rect 49849 44623 49868 44657
rect 49902 44623 49921 44657
rect 49849 44567 49921 44623
rect 50739 44638 50811 44661
rect 50739 44604 50758 44638
rect 50792 44604 50811 44638
rect 49849 44533 49868 44567
rect 49902 44533 49921 44567
rect 49849 44477 49921 44533
rect 49849 44443 49868 44477
rect 49902 44443 49921 44477
rect 49849 44387 49921 44443
rect 49849 44353 49868 44387
rect 49902 44353 49921 44387
rect 49849 44297 49921 44353
rect 49849 44263 49868 44297
rect 49902 44263 49921 44297
rect 49849 44207 49921 44263
rect 49849 44173 49868 44207
rect 49902 44173 49921 44207
rect 49849 44117 49921 44173
rect 49849 44083 49868 44117
rect 49902 44083 49921 44117
rect 49849 44027 49921 44083
rect 49849 43993 49868 44027
rect 49902 43993 49921 44027
rect 49849 43937 49921 43993
rect 49849 43903 49868 43937
rect 49902 43903 49921 43937
rect 49983 44540 50677 44599
rect 49983 44506 50044 44540
rect 50078 44512 50134 44540
rect 50168 44512 50224 44540
rect 50258 44512 50314 44540
rect 50090 44506 50134 44512
rect 50190 44506 50224 44512
rect 50290 44506 50314 44512
rect 50348 44512 50404 44540
rect 50348 44506 50356 44512
rect 49983 44478 50056 44506
rect 50090 44478 50156 44506
rect 50190 44478 50256 44506
rect 50290 44478 50356 44506
rect 50390 44506 50404 44512
rect 50438 44512 50494 44540
rect 50438 44506 50456 44512
rect 50390 44478 50456 44506
rect 50490 44506 50494 44512
rect 50528 44512 50584 44540
rect 50528 44506 50556 44512
rect 50618 44506 50677 44540
rect 50490 44478 50556 44506
rect 50590 44478 50677 44506
rect 49983 44450 50677 44478
rect 49983 44416 50044 44450
rect 50078 44416 50134 44450
rect 50168 44416 50224 44450
rect 50258 44416 50314 44450
rect 50348 44416 50404 44450
rect 50438 44416 50494 44450
rect 50528 44416 50584 44450
rect 50618 44416 50677 44450
rect 49983 44412 50677 44416
rect 49983 44378 50056 44412
rect 50090 44378 50156 44412
rect 50190 44378 50256 44412
rect 50290 44378 50356 44412
rect 50390 44378 50456 44412
rect 50490 44378 50556 44412
rect 50590 44378 50677 44412
rect 49983 44360 50677 44378
rect 49983 44326 50044 44360
rect 50078 44326 50134 44360
rect 50168 44326 50224 44360
rect 50258 44326 50314 44360
rect 50348 44326 50404 44360
rect 50438 44326 50494 44360
rect 50528 44326 50584 44360
rect 50618 44326 50677 44360
rect 49983 44312 50677 44326
rect 49983 44278 50056 44312
rect 50090 44278 50156 44312
rect 50190 44278 50256 44312
rect 50290 44278 50356 44312
rect 50390 44278 50456 44312
rect 50490 44278 50556 44312
rect 50590 44278 50677 44312
rect 49983 44270 50677 44278
rect 49983 44236 50044 44270
rect 50078 44236 50134 44270
rect 50168 44236 50224 44270
rect 50258 44236 50314 44270
rect 50348 44236 50404 44270
rect 50438 44236 50494 44270
rect 50528 44236 50584 44270
rect 50618 44236 50677 44270
rect 49983 44212 50677 44236
rect 49983 44180 50056 44212
rect 50090 44180 50156 44212
rect 50190 44180 50256 44212
rect 50290 44180 50356 44212
rect 49983 44146 50044 44180
rect 50090 44178 50134 44180
rect 50190 44178 50224 44180
rect 50290 44178 50314 44180
rect 50078 44146 50134 44178
rect 50168 44146 50224 44178
rect 50258 44146 50314 44178
rect 50348 44178 50356 44180
rect 50390 44180 50456 44212
rect 50390 44178 50404 44180
rect 50348 44146 50404 44178
rect 50438 44178 50456 44180
rect 50490 44180 50556 44212
rect 50590 44180 50677 44212
rect 50490 44178 50494 44180
rect 50438 44146 50494 44178
rect 50528 44178 50556 44180
rect 50528 44146 50584 44178
rect 50618 44146 50677 44180
rect 49983 44112 50677 44146
rect 49983 44090 50056 44112
rect 50090 44090 50156 44112
rect 50190 44090 50256 44112
rect 50290 44090 50356 44112
rect 49983 44056 50044 44090
rect 50090 44078 50134 44090
rect 50190 44078 50224 44090
rect 50290 44078 50314 44090
rect 50078 44056 50134 44078
rect 50168 44056 50224 44078
rect 50258 44056 50314 44078
rect 50348 44078 50356 44090
rect 50390 44090 50456 44112
rect 50390 44078 50404 44090
rect 50348 44056 50404 44078
rect 50438 44078 50456 44090
rect 50490 44090 50556 44112
rect 50590 44090 50677 44112
rect 50490 44078 50494 44090
rect 50438 44056 50494 44078
rect 50528 44078 50556 44090
rect 50528 44056 50584 44078
rect 50618 44056 50677 44090
rect 49983 44012 50677 44056
rect 49983 44000 50056 44012
rect 50090 44000 50156 44012
rect 50190 44000 50256 44012
rect 50290 44000 50356 44012
rect 49983 43966 50044 44000
rect 50090 43978 50134 44000
rect 50190 43978 50224 44000
rect 50290 43978 50314 44000
rect 50078 43966 50134 43978
rect 50168 43966 50224 43978
rect 50258 43966 50314 43978
rect 50348 43978 50356 44000
rect 50390 44000 50456 44012
rect 50390 43978 50404 44000
rect 50348 43966 50404 43978
rect 50438 43978 50456 44000
rect 50490 44000 50556 44012
rect 50590 44000 50677 44012
rect 50490 43978 50494 44000
rect 50438 43966 50494 43978
rect 50528 43978 50556 44000
rect 50528 43966 50584 43978
rect 50618 43966 50677 44000
rect 49983 43905 50677 43966
rect 50739 44548 50811 44604
rect 50739 44514 50758 44548
rect 50792 44514 50811 44548
rect 50739 44458 50811 44514
rect 50739 44424 50758 44458
rect 50792 44424 50811 44458
rect 50739 44368 50811 44424
rect 50739 44334 50758 44368
rect 50792 44334 50811 44368
rect 50739 44278 50811 44334
rect 50739 44244 50758 44278
rect 50792 44244 50811 44278
rect 50739 44188 50811 44244
rect 50739 44154 50758 44188
rect 50792 44154 50811 44188
rect 50739 44098 50811 44154
rect 50739 44064 50758 44098
rect 50792 44064 50811 44098
rect 50739 44008 50811 44064
rect 50739 43974 50758 44008
rect 50792 43974 50811 44008
rect 50739 43918 50811 43974
rect 49849 43843 49921 43903
rect 50739 43884 50758 43918
rect 50792 43884 50811 43918
rect 50739 43843 50811 43884
rect 49849 43824 50811 43843
rect 49849 43790 49946 43824
rect 49980 43790 50036 43824
rect 50070 43790 50126 43824
rect 50160 43790 50216 43824
rect 50250 43790 50306 43824
rect 50340 43790 50396 43824
rect 50430 43790 50486 43824
rect 50520 43790 50576 43824
rect 50610 43790 50666 43824
rect 50700 43790 50811 43824
rect 49849 43771 50811 43790
rect 50875 44714 50907 44748
rect 50941 44714 51060 44748
rect 51094 44714 51125 44748
rect 52215 44748 52314 44797
rect 50875 44658 51125 44714
rect 50875 44624 50907 44658
rect 50941 44624 51060 44658
rect 51094 44624 51125 44658
rect 50875 44568 51125 44624
rect 50875 44534 50907 44568
rect 50941 44534 51060 44568
rect 51094 44534 51125 44568
rect 50875 44478 51125 44534
rect 50875 44444 50907 44478
rect 50941 44444 51060 44478
rect 51094 44444 51125 44478
rect 50875 44388 51125 44444
rect 50875 44354 50907 44388
rect 50941 44354 51060 44388
rect 51094 44354 51125 44388
rect 50875 44298 51125 44354
rect 50875 44264 50907 44298
rect 50941 44264 51060 44298
rect 51094 44264 51125 44298
rect 50875 44208 51125 44264
rect 50875 44174 50907 44208
rect 50941 44174 51060 44208
rect 51094 44174 51125 44208
rect 50875 44118 51125 44174
rect 50875 44084 50907 44118
rect 50941 44084 51060 44118
rect 51094 44084 51125 44118
rect 50875 44028 51125 44084
rect 50875 43994 50907 44028
rect 50941 43994 51060 44028
rect 51094 43994 51125 44028
rect 50875 43938 51125 43994
rect 50875 43904 50907 43938
rect 50941 43904 51060 43938
rect 51094 43904 51125 43938
rect 50875 43848 51125 43904
rect 50875 43814 50907 43848
rect 50941 43814 51060 43848
rect 51094 43814 51125 43848
rect 49535 43724 49567 43758
rect 49601 43724 49720 43758
rect 49754 43724 49785 43758
rect 49535 43707 49785 43724
rect 50875 43758 51125 43814
rect 51189 44716 52151 44733
rect 51189 44682 51210 44716
rect 51244 44682 51300 44716
rect 51334 44714 51390 44716
rect 51424 44714 51480 44716
rect 51514 44714 51570 44716
rect 51604 44714 51660 44716
rect 51694 44714 51750 44716
rect 51784 44714 51840 44716
rect 51874 44714 51930 44716
rect 51964 44714 52020 44716
rect 52054 44714 52110 44716
rect 51354 44682 51390 44714
rect 51444 44682 51480 44714
rect 51534 44682 51570 44714
rect 51624 44682 51660 44714
rect 51714 44682 51750 44714
rect 51804 44682 51840 44714
rect 51894 44682 51930 44714
rect 51984 44682 52020 44714
rect 52074 44682 52110 44714
rect 52144 44682 52151 44716
rect 51189 44680 51320 44682
rect 51354 44680 51410 44682
rect 51444 44680 51500 44682
rect 51534 44680 51590 44682
rect 51624 44680 51680 44682
rect 51714 44680 51770 44682
rect 51804 44680 51860 44682
rect 51894 44680 51950 44682
rect 51984 44680 52040 44682
rect 52074 44680 52151 44682
rect 51189 44661 52151 44680
rect 51189 44657 51261 44661
rect 51189 44623 51208 44657
rect 51242 44623 51261 44657
rect 51189 44567 51261 44623
rect 52079 44638 52151 44661
rect 52079 44604 52098 44638
rect 52132 44604 52151 44638
rect 51189 44533 51208 44567
rect 51242 44533 51261 44567
rect 51189 44477 51261 44533
rect 51189 44443 51208 44477
rect 51242 44443 51261 44477
rect 51189 44387 51261 44443
rect 51189 44353 51208 44387
rect 51242 44353 51261 44387
rect 51189 44297 51261 44353
rect 51189 44263 51208 44297
rect 51242 44263 51261 44297
rect 51189 44207 51261 44263
rect 51189 44173 51208 44207
rect 51242 44173 51261 44207
rect 51189 44117 51261 44173
rect 51189 44083 51208 44117
rect 51242 44083 51261 44117
rect 51189 44027 51261 44083
rect 51189 43993 51208 44027
rect 51242 43993 51261 44027
rect 51189 43937 51261 43993
rect 51189 43903 51208 43937
rect 51242 43903 51261 43937
rect 51323 44540 52017 44599
rect 51323 44506 51384 44540
rect 51418 44512 51474 44540
rect 51508 44512 51564 44540
rect 51598 44512 51654 44540
rect 51430 44506 51474 44512
rect 51530 44506 51564 44512
rect 51630 44506 51654 44512
rect 51688 44512 51744 44540
rect 51688 44506 51696 44512
rect 51323 44478 51396 44506
rect 51430 44478 51496 44506
rect 51530 44478 51596 44506
rect 51630 44478 51696 44506
rect 51730 44506 51744 44512
rect 51778 44512 51834 44540
rect 51778 44506 51796 44512
rect 51730 44478 51796 44506
rect 51830 44506 51834 44512
rect 51868 44512 51924 44540
rect 51868 44506 51896 44512
rect 51958 44506 52017 44540
rect 51830 44478 51896 44506
rect 51930 44478 52017 44506
rect 51323 44450 52017 44478
rect 51323 44416 51384 44450
rect 51418 44416 51474 44450
rect 51508 44416 51564 44450
rect 51598 44416 51654 44450
rect 51688 44416 51744 44450
rect 51778 44416 51834 44450
rect 51868 44416 51924 44450
rect 51958 44416 52017 44450
rect 51323 44412 52017 44416
rect 51323 44378 51396 44412
rect 51430 44378 51496 44412
rect 51530 44378 51596 44412
rect 51630 44378 51696 44412
rect 51730 44378 51796 44412
rect 51830 44378 51896 44412
rect 51930 44378 52017 44412
rect 51323 44360 52017 44378
rect 51323 44326 51384 44360
rect 51418 44326 51474 44360
rect 51508 44326 51564 44360
rect 51598 44326 51654 44360
rect 51688 44326 51744 44360
rect 51778 44326 51834 44360
rect 51868 44326 51924 44360
rect 51958 44326 52017 44360
rect 51323 44312 52017 44326
rect 51323 44278 51396 44312
rect 51430 44278 51496 44312
rect 51530 44278 51596 44312
rect 51630 44278 51696 44312
rect 51730 44278 51796 44312
rect 51830 44278 51896 44312
rect 51930 44278 52017 44312
rect 51323 44270 52017 44278
rect 51323 44236 51384 44270
rect 51418 44236 51474 44270
rect 51508 44236 51564 44270
rect 51598 44236 51654 44270
rect 51688 44236 51744 44270
rect 51778 44236 51834 44270
rect 51868 44236 51924 44270
rect 51958 44236 52017 44270
rect 51323 44212 52017 44236
rect 51323 44180 51396 44212
rect 51430 44180 51496 44212
rect 51530 44180 51596 44212
rect 51630 44180 51696 44212
rect 51323 44146 51384 44180
rect 51430 44178 51474 44180
rect 51530 44178 51564 44180
rect 51630 44178 51654 44180
rect 51418 44146 51474 44178
rect 51508 44146 51564 44178
rect 51598 44146 51654 44178
rect 51688 44178 51696 44180
rect 51730 44180 51796 44212
rect 51730 44178 51744 44180
rect 51688 44146 51744 44178
rect 51778 44178 51796 44180
rect 51830 44180 51896 44212
rect 51930 44180 52017 44212
rect 51830 44178 51834 44180
rect 51778 44146 51834 44178
rect 51868 44178 51896 44180
rect 51868 44146 51924 44178
rect 51958 44146 52017 44180
rect 51323 44112 52017 44146
rect 51323 44090 51396 44112
rect 51430 44090 51496 44112
rect 51530 44090 51596 44112
rect 51630 44090 51696 44112
rect 51323 44056 51384 44090
rect 51430 44078 51474 44090
rect 51530 44078 51564 44090
rect 51630 44078 51654 44090
rect 51418 44056 51474 44078
rect 51508 44056 51564 44078
rect 51598 44056 51654 44078
rect 51688 44078 51696 44090
rect 51730 44090 51796 44112
rect 51730 44078 51744 44090
rect 51688 44056 51744 44078
rect 51778 44078 51796 44090
rect 51830 44090 51896 44112
rect 51930 44090 52017 44112
rect 51830 44078 51834 44090
rect 51778 44056 51834 44078
rect 51868 44078 51896 44090
rect 51868 44056 51924 44078
rect 51958 44056 52017 44090
rect 51323 44012 52017 44056
rect 51323 44000 51396 44012
rect 51430 44000 51496 44012
rect 51530 44000 51596 44012
rect 51630 44000 51696 44012
rect 51323 43966 51384 44000
rect 51430 43978 51474 44000
rect 51530 43978 51564 44000
rect 51630 43978 51654 44000
rect 51418 43966 51474 43978
rect 51508 43966 51564 43978
rect 51598 43966 51654 43978
rect 51688 43978 51696 44000
rect 51730 44000 51796 44012
rect 51730 43978 51744 44000
rect 51688 43966 51744 43978
rect 51778 43978 51796 44000
rect 51830 44000 51896 44012
rect 51930 44000 52017 44012
rect 51830 43978 51834 44000
rect 51778 43966 51834 43978
rect 51868 43978 51896 44000
rect 51868 43966 51924 43978
rect 51958 43966 52017 44000
rect 51323 43905 52017 43966
rect 52079 44548 52151 44604
rect 52079 44514 52098 44548
rect 52132 44514 52151 44548
rect 52079 44458 52151 44514
rect 52079 44424 52098 44458
rect 52132 44424 52151 44458
rect 52079 44368 52151 44424
rect 52079 44334 52098 44368
rect 52132 44334 52151 44368
rect 52079 44278 52151 44334
rect 52079 44244 52098 44278
rect 52132 44244 52151 44278
rect 52079 44188 52151 44244
rect 52079 44154 52098 44188
rect 52132 44154 52151 44188
rect 52079 44098 52151 44154
rect 52079 44064 52098 44098
rect 52132 44064 52151 44098
rect 52079 44008 52151 44064
rect 52079 43974 52098 44008
rect 52132 43974 52151 44008
rect 52079 43918 52151 43974
rect 51189 43843 51261 43903
rect 52079 43884 52098 43918
rect 52132 43884 52151 43918
rect 52079 43843 52151 43884
rect 51189 43824 52151 43843
rect 51189 43790 51286 43824
rect 51320 43790 51376 43824
rect 51410 43790 51466 43824
rect 51500 43790 51556 43824
rect 51590 43790 51646 43824
rect 51680 43790 51736 43824
rect 51770 43790 51826 43824
rect 51860 43790 51916 43824
rect 51950 43790 52006 43824
rect 52040 43790 52151 43824
rect 51189 43771 52151 43790
rect 52215 44714 52247 44748
rect 52281 44714 52314 44748
rect 52215 44658 52314 44714
rect 52215 44624 52247 44658
rect 52281 44624 52314 44658
rect 52215 44568 52314 44624
rect 52215 44534 52247 44568
rect 52281 44534 52314 44568
rect 52215 44478 52314 44534
rect 52215 44444 52247 44478
rect 52281 44444 52314 44478
rect 52215 44388 52314 44444
rect 52215 44354 52247 44388
rect 52281 44354 52314 44388
rect 52215 44298 52314 44354
rect 52215 44264 52247 44298
rect 52281 44264 52314 44298
rect 52215 44208 52314 44264
rect 52215 44174 52247 44208
rect 52281 44174 52314 44208
rect 52215 44118 52314 44174
rect 52215 44084 52247 44118
rect 52281 44084 52314 44118
rect 52215 44028 52314 44084
rect 52215 43994 52247 44028
rect 52281 43994 52314 44028
rect 52215 43938 52314 43994
rect 52215 43904 52247 43938
rect 52281 43904 52314 43938
rect 52215 43848 52314 43904
rect 52215 43814 52247 43848
rect 52281 43814 52314 43848
rect 50875 43724 50907 43758
rect 50941 43724 51060 43758
rect 51094 43724 51125 43758
rect 50875 43707 51125 43724
rect 52215 43758 52314 43814
rect 52215 43724 52247 43758
rect 52281 43724 52314 43758
rect 52215 43707 52314 43724
rect 42986 43674 52314 43707
rect 42986 43640 43116 43674
rect 43150 43640 43206 43674
rect 43240 43640 43296 43674
rect 43330 43640 43386 43674
rect 43420 43640 43476 43674
rect 43510 43640 43566 43674
rect 43600 43640 43656 43674
rect 43690 43640 43746 43674
rect 43780 43640 43836 43674
rect 43870 43640 43926 43674
rect 43960 43640 44016 43674
rect 44050 43640 44106 43674
rect 44140 43640 44456 43674
rect 44490 43640 44546 43674
rect 44580 43640 44636 43674
rect 44670 43640 44726 43674
rect 44760 43640 44816 43674
rect 44850 43640 44906 43674
rect 44940 43640 44996 43674
rect 45030 43640 45086 43674
rect 45120 43640 45176 43674
rect 45210 43640 45266 43674
rect 45300 43640 45356 43674
rect 45390 43640 45446 43674
rect 45480 43640 45796 43674
rect 45830 43640 45886 43674
rect 45920 43640 45976 43674
rect 46010 43640 46066 43674
rect 46100 43640 46156 43674
rect 46190 43640 46246 43674
rect 46280 43640 46336 43674
rect 46370 43640 46426 43674
rect 46460 43640 46516 43674
rect 46550 43640 46606 43674
rect 46640 43640 46696 43674
rect 46730 43640 46786 43674
rect 46820 43640 47136 43674
rect 47170 43640 47226 43674
rect 47260 43640 47316 43674
rect 47350 43640 47406 43674
rect 47440 43640 47496 43674
rect 47530 43640 47586 43674
rect 47620 43640 47676 43674
rect 47710 43640 47766 43674
rect 47800 43640 47856 43674
rect 47890 43640 47946 43674
rect 47980 43640 48036 43674
rect 48070 43640 48126 43674
rect 48160 43640 48476 43674
rect 48510 43640 48566 43674
rect 48600 43640 48656 43674
rect 48690 43640 48746 43674
rect 48780 43640 48836 43674
rect 48870 43640 48926 43674
rect 48960 43640 49016 43674
rect 49050 43640 49106 43674
rect 49140 43640 49196 43674
rect 49230 43640 49286 43674
rect 49320 43640 49376 43674
rect 49410 43640 49466 43674
rect 49500 43640 49816 43674
rect 49850 43640 49906 43674
rect 49940 43640 49996 43674
rect 50030 43640 50086 43674
rect 50120 43640 50176 43674
rect 50210 43640 50266 43674
rect 50300 43640 50356 43674
rect 50390 43640 50446 43674
rect 50480 43640 50536 43674
rect 50570 43640 50626 43674
rect 50660 43640 50716 43674
rect 50750 43640 50806 43674
rect 50840 43640 51156 43674
rect 51190 43640 51246 43674
rect 51280 43640 51336 43674
rect 51370 43640 51426 43674
rect 51460 43640 51516 43674
rect 51550 43640 51606 43674
rect 51640 43640 51696 43674
rect 51730 43640 51786 43674
rect 51820 43640 51876 43674
rect 51910 43640 51966 43674
rect 52000 43640 52056 43674
rect 52090 43640 52146 43674
rect 52180 43640 52314 43674
rect 42986 43608 52314 43640
rect 15030 43571 42638 43582
rect 14048 43469 14108 43552
rect 15059 43537 42638 43571
rect 15030 43522 42638 43537
rect 14048 43435 14061 43469
rect 14095 43435 14108 43469
rect 14198 43503 14634 43516
rect 14198 43469 14301 43503
rect 14335 43469 14565 43503
rect 14599 43469 14634 43503
rect 14198 43456 14634 43469
rect 15030 43469 42638 43476
rect 15030 43463 29469 43469
rect 14048 43342 14108 43435
rect 15030 43429 15213 43463
rect 15247 43429 15613 43463
rect 15647 43429 16013 43463
rect 16047 43429 16413 43463
rect 16447 43429 16813 43463
rect 16847 43429 17213 43463
rect 17247 43429 17613 43463
rect 17647 43429 18013 43463
rect 18047 43429 18413 43463
rect 18447 43429 18813 43463
rect 18847 43429 19213 43463
rect 19247 43429 19613 43463
rect 19647 43429 20013 43463
rect 20047 43429 20413 43463
rect 20447 43429 20813 43463
rect 20847 43429 21213 43463
rect 21247 43429 21613 43463
rect 21647 43429 22013 43463
rect 22047 43429 22413 43463
rect 22447 43429 22813 43463
rect 22847 43429 23213 43463
rect 23247 43429 23613 43463
rect 23647 43429 24013 43463
rect 24047 43429 24413 43463
rect 24447 43429 24813 43463
rect 24847 43429 25213 43463
rect 25247 43429 25613 43463
rect 25647 43429 26013 43463
rect 26047 43429 26413 43463
rect 26447 43429 26813 43463
rect 26847 43429 27213 43463
rect 27247 43429 27613 43463
rect 27647 43429 28013 43463
rect 28047 43429 28413 43463
rect 28447 43429 28813 43463
rect 28847 43429 29213 43463
rect 29247 43435 29469 43463
rect 29503 43463 42638 43469
rect 29503 43435 29613 43463
rect 29247 43429 29613 43435
rect 29647 43429 30013 43463
rect 30047 43429 30413 43463
rect 30447 43429 30813 43463
rect 30847 43429 31213 43463
rect 31247 43429 31613 43463
rect 31647 43429 32013 43463
rect 32047 43429 32413 43463
rect 32447 43429 32813 43463
rect 32847 43429 33213 43463
rect 33247 43429 33613 43463
rect 33647 43429 34013 43463
rect 34047 43429 34413 43463
rect 34447 43429 34813 43463
rect 34847 43429 35213 43463
rect 35247 43429 35613 43463
rect 35647 43429 36013 43463
rect 36047 43429 36413 43463
rect 36447 43429 36813 43463
rect 36847 43429 37213 43463
rect 37247 43429 37613 43463
rect 37647 43429 38013 43463
rect 38047 43429 38413 43463
rect 38447 43429 38813 43463
rect 38847 43429 39213 43463
rect 39247 43429 39613 43463
rect 39647 43429 40013 43463
rect 40047 43429 40413 43463
rect 40447 43429 40813 43463
rect 40847 43429 41213 43463
rect 41247 43429 41613 43463
rect 41647 43429 42013 43463
rect 42047 43429 42413 43463
rect 42447 43429 42638 43463
rect 15030 43416 42638 43429
rect 5918 43329 13086 43342
rect 5918 43295 6101 43329
rect 6135 43295 6501 43329
rect 6535 43295 6901 43329
rect 6935 43295 7301 43329
rect 7335 43295 7701 43329
rect 7735 43295 8101 43329
rect 8135 43295 8501 43329
rect 8535 43295 8901 43329
rect 8935 43295 9301 43329
rect 9335 43295 9701 43329
rect 9735 43295 10101 43329
rect 10135 43295 10501 43329
rect 10535 43295 10901 43329
rect 10935 43295 11301 43329
rect 11335 43295 11701 43329
rect 11735 43295 12101 43329
rect 12135 43295 12501 43329
rect 12535 43295 12901 43329
rect 12935 43295 13086 43329
rect 5918 43282 13086 43295
rect 14020 43329 14634 43342
rect 14020 43295 14301 43329
rect 14335 43295 14634 43329
rect 14020 43282 14634 43295
rect 14932 43329 42638 43342
rect 14932 43295 15213 43329
rect 15247 43295 15613 43329
rect 15647 43295 16013 43329
rect 16047 43295 16413 43329
rect 16447 43295 16813 43329
rect 16847 43295 17213 43329
rect 17247 43295 17613 43329
rect 17647 43295 18013 43329
rect 18047 43295 18413 43329
rect 18447 43295 18813 43329
rect 18847 43295 19213 43329
rect 19247 43295 19613 43329
rect 19647 43295 20013 43329
rect 20047 43295 20413 43329
rect 20447 43295 20813 43329
rect 20847 43295 21213 43329
rect 21247 43295 21613 43329
rect 21647 43295 22013 43329
rect 22047 43295 22413 43329
rect 22447 43295 22813 43329
rect 22847 43295 23213 43329
rect 23247 43295 23613 43329
rect 23647 43295 24013 43329
rect 24047 43295 24413 43329
rect 24447 43295 24813 43329
rect 24847 43295 25213 43329
rect 25247 43295 25613 43329
rect 25647 43295 26013 43329
rect 26047 43295 26413 43329
rect 26447 43295 26813 43329
rect 26847 43295 27213 43329
rect 27247 43295 27613 43329
rect 27647 43295 28013 43329
rect 28047 43295 28413 43329
rect 28447 43295 28813 43329
rect 28847 43295 29213 43329
rect 29247 43295 29613 43329
rect 29647 43295 30013 43329
rect 30047 43295 30413 43329
rect 30447 43295 30813 43329
rect 30847 43295 31213 43329
rect 31247 43295 31613 43329
rect 31647 43295 32013 43329
rect 32047 43295 32413 43329
rect 32447 43295 32813 43329
rect 32847 43295 33213 43329
rect 33247 43295 33613 43329
rect 33647 43295 34013 43329
rect 34047 43295 34413 43329
rect 34447 43295 34813 43329
rect 34847 43295 35213 43329
rect 35247 43295 35613 43329
rect 35647 43295 36013 43329
rect 36047 43295 36413 43329
rect 36447 43295 36813 43329
rect 36847 43295 37213 43329
rect 37247 43295 37613 43329
rect 37647 43295 38013 43329
rect 38047 43295 38413 43329
rect 38447 43295 38813 43329
rect 38847 43295 39213 43329
rect 39247 43295 39613 43329
rect 39647 43295 40013 43329
rect 40047 43295 40413 43329
rect 40447 43295 40813 43329
rect 40847 43295 41213 43329
rect 41247 43295 41613 43329
rect 41647 43295 42013 43329
rect 42047 43295 42413 43329
rect 42447 43295 42638 43329
rect 14932 43282 42638 43295
rect 42960 43329 52340 43342
rect 42960 43295 43143 43329
rect 43177 43295 43343 43329
rect 43377 43295 43543 43329
rect 43577 43295 43743 43329
rect 43777 43295 43943 43329
rect 43977 43295 44143 43329
rect 44177 43295 44343 43329
rect 44377 43295 44543 43329
rect 44577 43295 44743 43329
rect 44777 43295 44943 43329
rect 44977 43295 45143 43329
rect 45177 43295 45343 43329
rect 45377 43295 45543 43329
rect 45577 43295 45743 43329
rect 45777 43295 45943 43329
rect 45977 43295 46143 43329
rect 46177 43295 46343 43329
rect 46377 43295 46543 43329
rect 46577 43295 46743 43329
rect 46777 43295 46943 43329
rect 46977 43295 47143 43329
rect 47177 43295 47343 43329
rect 47377 43295 47543 43329
rect 47577 43295 47743 43329
rect 47777 43295 47943 43329
rect 47977 43295 48143 43329
rect 48177 43295 48343 43329
rect 48377 43295 48543 43329
rect 48577 43295 48743 43329
rect 48777 43295 48943 43329
rect 48977 43295 49143 43329
rect 49177 43295 49343 43329
rect 49377 43295 49543 43329
rect 49577 43295 49743 43329
rect 49777 43295 49943 43329
rect 49977 43295 50143 43329
rect 50177 43295 50343 43329
rect 50377 43295 50543 43329
rect 50577 43295 50743 43329
rect 50777 43295 50943 43329
rect 50977 43295 51143 43329
rect 51177 43295 51343 43329
rect 51377 43295 51543 43329
rect 51577 43295 51743 43329
rect 51777 43295 51943 43329
rect 51977 43295 52143 43329
rect 52177 43295 52340 43329
rect 42960 43282 52340 43295
rect 6310 41449 13478 41462
rect 6310 41415 6493 41449
rect 6527 41415 6893 41449
rect 6927 41415 7293 41449
rect 7327 41415 7693 41449
rect 7727 41415 8093 41449
rect 8127 41415 8493 41449
rect 8527 41415 8893 41449
rect 8927 41415 9293 41449
rect 9327 41415 9693 41449
rect 9727 41415 10093 41449
rect 10127 41415 10493 41449
rect 10527 41415 10893 41449
rect 10927 41415 11293 41449
rect 11327 41415 11693 41449
rect 11727 41415 12093 41449
rect 12127 41415 12493 41449
rect 12527 41415 12893 41449
rect 12927 41415 13293 41449
rect 13327 41415 13478 41449
rect 6310 41402 13478 41415
rect 15130 41449 22298 41462
rect 15130 41415 15313 41449
rect 15347 41415 15713 41449
rect 15747 41415 16113 41449
rect 16147 41415 16513 41449
rect 16547 41415 16913 41449
rect 16947 41415 17313 41449
rect 17347 41415 17713 41449
rect 17747 41415 18113 41449
rect 18147 41415 18513 41449
rect 18547 41415 18913 41449
rect 18947 41415 19313 41449
rect 19347 41415 19713 41449
rect 19747 41415 20113 41449
rect 20147 41415 20513 41449
rect 20547 41415 20913 41449
rect 20947 41415 21313 41449
rect 21347 41415 21713 41449
rect 21747 41415 22113 41449
rect 22147 41415 22298 41449
rect 15130 41402 22298 41415
rect 22576 41449 28298 41462
rect 22576 41415 22857 41449
rect 22891 41415 23257 41449
rect 23291 41415 23657 41449
rect 23691 41415 24057 41449
rect 24091 41415 24457 41449
rect 24491 41415 24857 41449
rect 24891 41415 25257 41449
rect 25291 41415 25657 41449
rect 25691 41415 26057 41449
rect 26091 41415 26457 41449
rect 26491 41415 26857 41449
rect 26891 41415 27257 41449
rect 27291 41415 27657 41449
rect 27691 41415 28057 41449
rect 28091 41415 28298 41449
rect 22576 41402 28298 41415
rect 29240 41449 34962 41462
rect 29240 41415 29521 41449
rect 29555 41415 29921 41449
rect 29955 41415 30321 41449
rect 30355 41415 30721 41449
rect 30755 41415 31121 41449
rect 31155 41415 31521 41449
rect 31555 41415 31921 41449
rect 31955 41415 32321 41449
rect 32355 41415 32721 41449
rect 32755 41415 33121 41449
rect 33155 41415 33521 41449
rect 33555 41415 33921 41449
rect 33955 41415 34321 41449
rect 34355 41415 34721 41449
rect 34755 41415 34962 41449
rect 29240 41402 34962 41415
rect 37178 41449 41456 41462
rect 37178 41415 37459 41449
rect 37493 41415 37859 41449
rect 37893 41415 38259 41449
rect 38293 41415 38659 41449
rect 38693 41415 39059 41449
rect 39093 41415 39459 41449
rect 39493 41415 39859 41449
rect 39893 41415 40259 41449
rect 40293 41415 40659 41449
rect 40693 41415 41059 41449
rect 41093 41415 41456 41449
rect 37178 41402 41456 41415
rect 41784 41449 52504 41462
rect 41784 41415 41967 41449
rect 42001 41415 42167 41449
rect 42201 41415 42367 41449
rect 42401 41415 42567 41449
rect 42601 41415 42767 41449
rect 42801 41415 42967 41449
rect 43001 41415 43167 41449
rect 43201 41415 43367 41449
rect 43401 41415 43567 41449
rect 43601 41415 43767 41449
rect 43801 41415 43967 41449
rect 44001 41415 44167 41449
rect 44201 41415 44367 41449
rect 44401 41415 44567 41449
rect 44601 41415 44767 41449
rect 44801 41415 44967 41449
rect 45001 41415 45167 41449
rect 45201 41415 45367 41449
rect 45401 41415 45567 41449
rect 45601 41415 45767 41449
rect 45801 41415 45967 41449
rect 46001 41415 46167 41449
rect 46201 41415 46367 41449
rect 46401 41415 46567 41449
rect 46601 41415 46767 41449
rect 46801 41415 46967 41449
rect 47001 41415 47167 41449
rect 47201 41415 47367 41449
rect 47401 41415 47567 41449
rect 47601 41415 47767 41449
rect 47801 41415 47967 41449
rect 48001 41415 48167 41449
rect 48201 41415 48367 41449
rect 48401 41415 48567 41449
rect 48601 41415 48767 41449
rect 48801 41415 48967 41449
rect 49001 41415 49167 41449
rect 49201 41415 49367 41449
rect 49401 41415 49567 41449
rect 49601 41415 49767 41449
rect 49801 41415 49967 41449
rect 50001 41415 50167 41449
rect 50201 41415 50367 41449
rect 50401 41415 50567 41449
rect 50601 41415 50767 41449
rect 50801 41415 50967 41449
rect 51001 41415 51167 41449
rect 51201 41415 51367 41449
rect 51401 41415 51567 41449
rect 51601 41415 51767 41449
rect 51801 41415 51967 41449
rect 52001 41415 52167 41449
rect 52201 41415 52367 41449
rect 52401 41415 52504 41449
rect 41784 41402 52504 41415
rect 22604 41309 22664 41402
rect 23652 41359 23812 41402
rect 23652 41325 23717 41359
rect 23751 41325 23812 41359
rect 23652 41322 23812 41325
rect 24952 41359 25112 41402
rect 24952 41325 25017 41359
rect 25051 41325 25112 41359
rect 24952 41322 25112 41325
rect 26252 41359 26412 41402
rect 26252 41325 26317 41359
rect 26351 41325 26412 41359
rect 26252 41322 26412 41325
rect 22604 41275 22617 41309
rect 22651 41275 22664 41309
rect 29268 41309 29328 41402
rect 30316 41359 30476 41402
rect 30316 41325 30381 41359
rect 30415 41325 30476 41359
rect 30316 41322 30476 41325
rect 31616 41359 31776 41402
rect 31616 41325 31681 41359
rect 31715 41325 31776 41359
rect 31616 41322 31776 41325
rect 32916 41359 33076 41402
rect 32916 41325 32981 41359
rect 33015 41325 33076 41359
rect 32916 41322 33076 41325
rect 22604 41192 22664 41275
rect 22734 41259 28298 41282
rect 22734 41242 24869 41259
rect 22721 41181 22755 41201
rect 22721 41113 22755 41147
rect 22721 41045 22755 41075
rect 22721 40977 22755 41003
rect 22721 40909 22755 40931
rect 22721 40841 22755 40859
rect 22721 40773 22755 40787
rect 22721 40705 22755 40715
rect 22721 40637 22755 40643
rect 22721 40569 22755 40571
rect 22721 40533 22755 40535
rect 22721 40461 22755 40467
rect 22721 40389 22755 40399
rect 22721 40317 22755 40331
rect 22721 40245 22755 40263
rect 22721 40173 22755 40195
rect 22721 40101 22755 40127
rect 22721 40029 22755 40059
rect 22721 39957 22755 39991
rect 22721 39831 22755 39923
rect 23179 41181 23213 41242
rect 23179 41113 23213 41147
rect 23179 41045 23213 41075
rect 23179 40977 23213 41003
rect 23179 40909 23213 40931
rect 23179 40841 23213 40859
rect 23179 40773 23213 40787
rect 23179 40705 23213 40715
rect 23179 40637 23213 40643
rect 23179 40569 23213 40571
rect 23179 40533 23213 40535
rect 23179 40461 23213 40467
rect 23179 40389 23213 40399
rect 23179 40317 23213 40331
rect 23179 40245 23213 40263
rect 23179 40173 23213 40195
rect 23179 40101 23213 40127
rect 23179 40029 23213 40059
rect 23179 39957 23213 39991
rect 23179 39903 23213 39923
rect 23637 41181 23671 41201
rect 23637 41113 23671 41147
rect 23637 41045 23671 41075
rect 23637 40977 23671 41003
rect 23637 40909 23671 40931
rect 23637 40841 23671 40859
rect 23637 40773 23671 40787
rect 23637 40705 23671 40715
rect 23637 40637 23671 40643
rect 23637 40569 23671 40571
rect 23637 40533 23671 40535
rect 23637 40461 23671 40467
rect 23637 40389 23671 40399
rect 23637 40317 23671 40331
rect 23637 40245 23671 40263
rect 23637 40173 23671 40195
rect 23637 40101 23671 40127
rect 23637 40029 23671 40059
rect 23637 39957 23671 39991
rect 22721 39822 22753 39831
rect 22674 39797 22753 39822
rect 23637 39822 23671 39923
rect 24095 41181 24129 41242
rect 24903 41242 28298 41259
rect 29268 41275 29281 41309
rect 29315 41275 29328 41309
rect 24095 41113 24129 41147
rect 24095 41045 24129 41075
rect 24095 40977 24129 41003
rect 24095 40909 24129 40931
rect 24095 40841 24129 40859
rect 24095 40773 24129 40787
rect 24095 40705 24129 40715
rect 24095 40637 24129 40643
rect 24095 40569 24129 40571
rect 24095 40533 24129 40535
rect 24095 40461 24129 40467
rect 24095 40389 24129 40399
rect 24095 40317 24129 40331
rect 24095 40245 24129 40263
rect 24095 40173 24129 40195
rect 24095 40101 24129 40127
rect 24095 40029 24129 40059
rect 24095 39957 24129 39991
rect 24095 39903 24129 39923
rect 24553 41181 24587 41201
rect 24553 41113 24587 41147
rect 24553 41045 24587 41075
rect 24553 40977 24587 41003
rect 24553 40909 24587 40931
rect 24553 40841 24587 40859
rect 24553 40773 24587 40787
rect 24553 40705 24587 40715
rect 24553 40637 24587 40643
rect 24553 40569 24587 40571
rect 24553 40533 24587 40535
rect 24553 40461 24587 40467
rect 24553 40389 24587 40399
rect 24553 40317 24587 40331
rect 24553 40245 24587 40263
rect 24553 40173 24587 40195
rect 24553 40101 24587 40127
rect 24553 40029 24587 40059
rect 24553 39957 24587 39991
rect 24553 39822 24587 39923
rect 25011 41181 25045 41242
rect 25011 41113 25045 41147
rect 25011 41045 25045 41075
rect 25011 40977 25045 41003
rect 25011 40909 25045 40931
rect 25011 40841 25045 40859
rect 25011 40773 25045 40787
rect 25011 40705 25045 40715
rect 25011 40637 25045 40643
rect 25011 40569 25045 40571
rect 25011 40533 25045 40535
rect 25011 40461 25045 40467
rect 25011 40389 25045 40399
rect 25011 40317 25045 40331
rect 25011 40245 25045 40263
rect 25011 40173 25045 40195
rect 25011 40101 25045 40127
rect 25011 40029 25045 40059
rect 25011 39957 25045 39991
rect 25011 39903 25045 39923
rect 25469 41181 25503 41201
rect 25469 41113 25503 41147
rect 25469 41045 25503 41075
rect 25469 40977 25503 41003
rect 25469 40909 25503 40931
rect 25469 40841 25503 40859
rect 25469 40773 25503 40787
rect 25469 40705 25503 40715
rect 25469 40637 25503 40643
rect 25469 40569 25503 40571
rect 25469 40533 25503 40535
rect 25469 40461 25503 40467
rect 25469 40389 25503 40399
rect 25469 40317 25503 40331
rect 25469 40245 25503 40263
rect 25469 40173 25503 40195
rect 25469 40101 25503 40127
rect 25469 40029 25503 40059
rect 25469 39957 25503 39991
rect 25469 39822 25503 39923
rect 25927 41181 25961 41242
rect 25927 41113 25961 41147
rect 25927 41045 25961 41075
rect 25927 40977 25961 41003
rect 25927 40909 25961 40931
rect 25927 40841 25961 40859
rect 25927 40773 25961 40787
rect 25927 40705 25961 40715
rect 25927 40637 25961 40643
rect 25927 40569 25961 40571
rect 25927 40533 25961 40535
rect 25927 40461 25961 40467
rect 25927 40389 25961 40399
rect 25927 40317 25961 40331
rect 25927 40245 25961 40263
rect 25927 40173 25961 40195
rect 25927 40101 25961 40127
rect 25927 40029 25961 40059
rect 25927 39957 25961 39991
rect 25927 39903 25961 39923
rect 26385 41181 26419 41201
rect 26385 41113 26419 41147
rect 26385 41045 26419 41075
rect 26385 40977 26419 41003
rect 26385 40909 26419 40931
rect 26385 40841 26419 40859
rect 26385 40773 26419 40787
rect 26385 40705 26419 40715
rect 26385 40637 26419 40643
rect 26385 40569 26419 40571
rect 26385 40533 26419 40535
rect 26385 40461 26419 40467
rect 26385 40389 26419 40399
rect 26385 40317 26419 40331
rect 26385 40245 26419 40263
rect 26385 40173 26419 40195
rect 26385 40101 26419 40127
rect 26385 40029 26419 40059
rect 26385 39957 26419 39991
rect 26385 39822 26419 39923
rect 26843 41181 26877 41242
rect 26843 41113 26877 41147
rect 26843 41045 26877 41075
rect 26843 40977 26877 41003
rect 26843 40909 26877 40931
rect 26843 40841 26877 40859
rect 26843 40773 26877 40787
rect 26843 40705 26877 40715
rect 26843 40637 26877 40643
rect 26843 40569 26877 40571
rect 26843 40533 26877 40535
rect 26843 40461 26877 40467
rect 26843 40389 26877 40399
rect 26843 40317 26877 40331
rect 26843 40245 26877 40263
rect 26843 40173 26877 40195
rect 26843 40101 26877 40127
rect 26843 40029 26877 40059
rect 26843 39957 26877 39991
rect 26843 39903 26877 39923
rect 27301 41181 27335 41201
rect 27301 41113 27335 41147
rect 27301 41045 27335 41075
rect 27301 40977 27335 41003
rect 27301 40909 27335 40931
rect 27301 40841 27335 40859
rect 27301 40773 27335 40787
rect 27301 40705 27335 40715
rect 27301 40637 27335 40643
rect 27301 40569 27335 40571
rect 27301 40533 27335 40535
rect 27301 40461 27335 40467
rect 27301 40389 27335 40399
rect 27301 40317 27335 40331
rect 27301 40245 27335 40263
rect 27301 40173 27335 40195
rect 27301 40101 27335 40127
rect 27301 40029 27335 40059
rect 27301 39957 27335 39991
rect 27301 39822 27335 39923
rect 27759 41181 27793 41242
rect 27759 41113 27793 41147
rect 27759 41045 27793 41075
rect 27759 40977 27793 41003
rect 27759 40909 27793 40931
rect 27759 40841 27793 40859
rect 27759 40773 27793 40787
rect 27759 40705 27793 40715
rect 27759 40637 27793 40643
rect 27759 40569 27793 40571
rect 27759 40533 27793 40535
rect 27759 40461 27793 40467
rect 27759 40389 27793 40399
rect 27759 40317 27793 40331
rect 27759 40245 27793 40263
rect 27759 40173 27793 40195
rect 27759 40101 27793 40127
rect 27759 40029 27793 40059
rect 27759 39957 27793 39991
rect 27759 39903 27793 39923
rect 28217 41181 28251 41201
rect 29268 41192 29328 41275
rect 29398 41242 34962 41282
rect 37276 41242 41456 41302
rect 28217 41113 28251 41147
rect 28217 41045 28251 41075
rect 28217 40977 28251 41003
rect 28217 40909 28251 40931
rect 28217 40841 28251 40859
rect 28217 40773 28251 40787
rect 28217 40705 28251 40715
rect 28217 40637 28251 40643
rect 28217 40569 28251 40571
rect 28217 40533 28251 40535
rect 28217 40461 28251 40467
rect 28217 40389 28251 40399
rect 28217 40317 28251 40331
rect 28217 40245 28251 40263
rect 28217 40173 28251 40195
rect 28217 40101 28251 40127
rect 28217 40029 28251 40059
rect 28217 39957 28251 39991
rect 22787 39797 28089 39822
rect 28217 39822 28251 39923
rect 29385 41181 29419 41201
rect 29385 41113 29419 41147
rect 29385 41045 29419 41075
rect 29385 40977 29419 41003
rect 29385 40909 29419 40931
rect 29385 40841 29419 40859
rect 29385 40773 29419 40787
rect 29385 40705 29419 40715
rect 29385 40637 29419 40643
rect 29385 40569 29419 40571
rect 29385 40533 29419 40535
rect 29385 40461 29419 40467
rect 29385 40389 29419 40399
rect 29385 40317 29419 40331
rect 29385 40245 29419 40263
rect 29385 40173 29419 40195
rect 29385 40101 29419 40127
rect 29385 40029 29419 40059
rect 29385 39957 29419 39991
rect 29385 39822 29419 39923
rect 29843 41181 29877 41242
rect 29843 41113 29877 41147
rect 29843 41045 29877 41075
rect 29843 40977 29877 41003
rect 29843 40909 29877 40931
rect 29843 40841 29877 40859
rect 29843 40773 29877 40787
rect 29843 40705 29877 40715
rect 29843 40637 29877 40643
rect 29843 40569 29877 40571
rect 29843 40533 29877 40535
rect 29843 40461 29877 40467
rect 29843 40389 29877 40399
rect 29843 40317 29877 40331
rect 29843 40245 29877 40263
rect 29843 40173 29877 40195
rect 29843 40101 29877 40127
rect 29843 40029 29877 40059
rect 29843 39957 29877 39991
rect 29843 39903 29877 39923
rect 30301 41181 30335 41201
rect 30301 41113 30335 41147
rect 30301 41045 30335 41075
rect 30301 40977 30335 41003
rect 30301 40909 30335 40931
rect 30301 40841 30335 40859
rect 30301 40773 30335 40787
rect 30301 40705 30335 40715
rect 30301 40637 30335 40643
rect 30301 40569 30335 40571
rect 30301 40533 30335 40535
rect 30301 40461 30335 40467
rect 30301 40389 30335 40399
rect 30301 40317 30335 40331
rect 30301 40245 30335 40263
rect 30301 40173 30335 40195
rect 30301 40101 30335 40127
rect 30301 40029 30335 40059
rect 30301 39957 30335 39991
rect 30301 39822 30335 39923
rect 30759 41181 30793 41242
rect 30759 41113 30793 41147
rect 30759 41045 30793 41075
rect 30759 40977 30793 41003
rect 30759 40909 30793 40931
rect 30759 40841 30793 40859
rect 30759 40773 30793 40787
rect 30759 40705 30793 40715
rect 30759 40637 30793 40643
rect 30759 40569 30793 40571
rect 30759 40533 30793 40535
rect 30759 40461 30793 40467
rect 30759 40389 30793 40399
rect 30759 40317 30793 40331
rect 30759 40245 30793 40263
rect 30759 40173 30793 40195
rect 30759 40101 30793 40127
rect 30759 40029 30793 40059
rect 30759 39957 30793 39991
rect 30759 39903 30793 39923
rect 31217 41181 31251 41201
rect 31217 41113 31251 41147
rect 31217 41045 31251 41075
rect 31217 40977 31251 41003
rect 31217 40909 31251 40931
rect 31217 40841 31251 40859
rect 31217 40773 31251 40787
rect 31217 40705 31251 40715
rect 31217 40637 31251 40643
rect 31217 40569 31251 40571
rect 31217 40533 31251 40535
rect 31217 40461 31251 40467
rect 31217 40389 31251 40399
rect 31217 40317 31251 40331
rect 31217 40245 31251 40263
rect 31217 40173 31251 40195
rect 31217 40101 31251 40127
rect 31217 40029 31251 40059
rect 31217 39957 31251 39991
rect 31217 39822 31251 39923
rect 31675 41181 31709 41242
rect 31675 41113 31709 41147
rect 31675 41045 31709 41075
rect 31675 40977 31709 41003
rect 31675 40909 31709 40931
rect 31675 40841 31709 40859
rect 31675 40773 31709 40787
rect 31675 40705 31709 40715
rect 31675 40637 31709 40643
rect 31675 40569 31709 40571
rect 31675 40533 31709 40535
rect 31675 40461 31709 40467
rect 31675 40389 31709 40399
rect 31675 40317 31709 40331
rect 31675 40245 31709 40263
rect 31675 40173 31709 40195
rect 31675 40101 31709 40127
rect 31675 40029 31709 40059
rect 31675 39957 31709 39991
rect 31675 39903 31709 39923
rect 32133 41181 32167 41201
rect 32133 41113 32167 41147
rect 32133 41045 32167 41075
rect 32133 40977 32167 41003
rect 32133 40909 32167 40931
rect 32133 40841 32167 40859
rect 32133 40773 32167 40787
rect 32133 40705 32167 40715
rect 32133 40637 32167 40643
rect 32133 40569 32167 40571
rect 32133 40533 32167 40535
rect 32133 40461 32167 40467
rect 32133 40389 32167 40399
rect 32133 40317 32167 40331
rect 32133 40245 32167 40263
rect 32133 40173 32167 40195
rect 32133 40101 32167 40127
rect 32133 40029 32167 40059
rect 32133 39957 32167 39991
rect 32133 39822 32167 39923
rect 32591 41181 32625 41242
rect 32591 41113 32625 41147
rect 32591 41045 32625 41075
rect 32591 40977 32625 41003
rect 32591 40909 32625 40931
rect 32591 40841 32625 40859
rect 32591 40773 32625 40787
rect 32591 40705 32625 40715
rect 32591 40637 32625 40643
rect 32591 40569 32625 40571
rect 32591 40533 32625 40535
rect 32591 40461 32625 40467
rect 32591 40389 32625 40399
rect 32591 40317 32625 40331
rect 32591 40245 32625 40263
rect 32591 40173 32625 40195
rect 32591 40101 32625 40127
rect 32591 40029 32625 40059
rect 32591 39957 32625 39991
rect 32591 39903 32625 39923
rect 33049 41181 33083 41201
rect 33049 41113 33083 41147
rect 33049 41045 33083 41075
rect 33049 40977 33083 41003
rect 33049 40909 33083 40931
rect 33049 40841 33083 40859
rect 33049 40773 33083 40787
rect 33049 40705 33083 40715
rect 33049 40637 33083 40643
rect 33049 40569 33083 40571
rect 33049 40533 33083 40535
rect 33049 40461 33083 40467
rect 33049 40389 33083 40399
rect 33049 40317 33083 40331
rect 33049 40245 33083 40263
rect 33049 40173 33083 40195
rect 33049 40101 33083 40127
rect 33049 40029 33083 40059
rect 33049 39957 33083 39991
rect 33049 39822 33083 39923
rect 33507 41181 33541 41242
rect 33507 41113 33541 41147
rect 33507 41045 33541 41075
rect 33507 40977 33541 41003
rect 33507 40909 33541 40931
rect 33507 40841 33541 40859
rect 33507 40773 33541 40787
rect 33507 40705 33541 40715
rect 33507 40637 33541 40643
rect 33507 40569 33541 40571
rect 33507 40533 33541 40535
rect 33507 40461 33541 40467
rect 33507 40389 33541 40399
rect 33507 40317 33541 40331
rect 33507 40245 33541 40263
rect 33507 40173 33541 40195
rect 33507 40101 33541 40127
rect 33507 40029 33541 40059
rect 33507 39957 33541 39991
rect 33507 39903 33541 39923
rect 33965 41181 33999 41201
rect 33965 41113 33999 41147
rect 33965 41045 33999 41075
rect 33965 40977 33999 41003
rect 33965 40909 33999 40931
rect 33965 40841 33999 40859
rect 33965 40773 33999 40787
rect 33965 40705 33999 40715
rect 33965 40637 33999 40643
rect 33965 40569 33999 40571
rect 33965 40533 33999 40535
rect 33965 40461 33999 40467
rect 33965 40389 33999 40399
rect 33965 40317 33999 40331
rect 33965 40245 33999 40263
rect 33965 40173 33999 40195
rect 33965 40101 33999 40127
rect 33965 40029 33999 40059
rect 33965 39957 33999 39991
rect 33965 39822 33999 39923
rect 34423 41181 34457 41242
rect 34423 41113 34457 41147
rect 34423 41045 34457 41075
rect 34423 40977 34457 41003
rect 34423 40909 34457 40931
rect 34423 40841 34457 40859
rect 34423 40773 34457 40787
rect 34423 40705 34457 40715
rect 34423 40637 34457 40643
rect 34423 40569 34457 40571
rect 34423 40533 34457 40535
rect 34423 40461 34457 40467
rect 34423 40389 34457 40399
rect 34423 40317 34457 40331
rect 34423 40245 34457 40263
rect 34423 40173 34457 40195
rect 34423 40101 34457 40127
rect 34423 40029 34457 40059
rect 34423 39957 34457 39991
rect 34423 39903 34457 39923
rect 34881 41181 34915 41201
rect 34881 41113 34915 41147
rect 34881 41045 34915 41075
rect 34881 40977 34915 41003
rect 37745 40956 37779 41242
rect 38661 40956 38695 41242
rect 39577 40956 39611 41242
rect 40493 40956 40527 41242
rect 41409 40956 41443 41242
rect 41810 41116 52478 41136
rect 41810 41082 41830 41116
rect 41864 41082 41920 41116
rect 41954 41101 42010 41116
rect 42044 41101 42100 41116
rect 42134 41101 42190 41116
rect 42224 41101 42280 41116
rect 42314 41101 42370 41116
rect 42404 41101 42460 41116
rect 42494 41101 42550 41116
rect 42584 41101 42640 41116
rect 42674 41101 42730 41116
rect 42764 41101 42820 41116
rect 42854 41101 42910 41116
rect 42944 41101 43000 41116
rect 41974 41082 42010 41101
rect 42064 41082 42100 41101
rect 42154 41082 42190 41101
rect 42244 41082 42280 41101
rect 42334 41082 42370 41101
rect 42424 41082 42460 41101
rect 42514 41082 42550 41101
rect 42604 41082 42640 41101
rect 42694 41082 42730 41101
rect 42784 41082 42820 41101
rect 42874 41082 42910 41101
rect 42964 41082 43000 41101
rect 43034 41082 43170 41116
rect 43204 41082 43260 41116
rect 43294 41101 43350 41116
rect 43384 41101 43440 41116
rect 43474 41101 43530 41116
rect 43564 41101 43620 41116
rect 43654 41101 43710 41116
rect 43744 41101 43800 41116
rect 43834 41101 43890 41116
rect 43924 41101 43980 41116
rect 44014 41101 44070 41116
rect 44104 41101 44160 41116
rect 44194 41101 44250 41116
rect 44284 41101 44340 41116
rect 43314 41082 43350 41101
rect 43404 41082 43440 41101
rect 43494 41082 43530 41101
rect 43584 41082 43620 41101
rect 43674 41082 43710 41101
rect 43764 41082 43800 41101
rect 43854 41082 43890 41101
rect 43944 41082 43980 41101
rect 44034 41082 44070 41101
rect 44124 41082 44160 41101
rect 44214 41082 44250 41101
rect 44304 41082 44340 41101
rect 44374 41082 44510 41116
rect 44544 41082 44600 41116
rect 44634 41101 44690 41116
rect 44724 41101 44780 41116
rect 44814 41101 44870 41116
rect 44904 41101 44960 41116
rect 44994 41101 45050 41116
rect 45084 41101 45140 41116
rect 45174 41101 45230 41116
rect 45264 41101 45320 41116
rect 45354 41101 45410 41116
rect 45444 41101 45500 41116
rect 45534 41101 45590 41116
rect 45624 41101 45680 41116
rect 44654 41082 44690 41101
rect 44744 41082 44780 41101
rect 44834 41082 44870 41101
rect 44924 41082 44960 41101
rect 45014 41082 45050 41101
rect 45104 41082 45140 41101
rect 45194 41082 45230 41101
rect 45284 41082 45320 41101
rect 45374 41082 45410 41101
rect 45464 41082 45500 41101
rect 45554 41082 45590 41101
rect 45644 41082 45680 41101
rect 45714 41082 45850 41116
rect 45884 41082 45940 41116
rect 45974 41101 46030 41116
rect 46064 41101 46120 41116
rect 46154 41101 46210 41116
rect 46244 41101 46300 41116
rect 46334 41101 46390 41116
rect 46424 41101 46480 41116
rect 46514 41101 46570 41116
rect 46604 41101 46660 41116
rect 46694 41101 46750 41116
rect 46784 41101 46840 41116
rect 46874 41101 46930 41116
rect 46964 41101 47020 41116
rect 45994 41082 46030 41101
rect 46084 41082 46120 41101
rect 46174 41082 46210 41101
rect 46264 41082 46300 41101
rect 46354 41082 46390 41101
rect 46444 41082 46480 41101
rect 46534 41082 46570 41101
rect 46624 41082 46660 41101
rect 46714 41082 46750 41101
rect 46804 41082 46840 41101
rect 46894 41082 46930 41101
rect 46984 41082 47020 41101
rect 47054 41082 47190 41116
rect 47224 41082 47280 41116
rect 47314 41101 47370 41116
rect 47404 41101 47460 41116
rect 47494 41101 47550 41116
rect 47584 41101 47640 41116
rect 47674 41101 47730 41116
rect 47764 41101 47820 41116
rect 47854 41101 47910 41116
rect 47944 41101 48000 41116
rect 48034 41101 48090 41116
rect 48124 41101 48180 41116
rect 48214 41101 48270 41116
rect 48304 41101 48360 41116
rect 47334 41082 47370 41101
rect 47424 41082 47460 41101
rect 47514 41082 47550 41101
rect 47604 41082 47640 41101
rect 47694 41082 47730 41101
rect 47784 41082 47820 41101
rect 47874 41082 47910 41101
rect 47964 41082 48000 41101
rect 48054 41082 48090 41101
rect 48144 41082 48180 41101
rect 48234 41082 48270 41101
rect 48324 41082 48360 41101
rect 48394 41082 48530 41116
rect 48564 41082 48620 41116
rect 48654 41101 48710 41116
rect 48744 41101 48800 41116
rect 48834 41101 48890 41116
rect 48924 41101 48980 41116
rect 49014 41101 49070 41116
rect 49104 41101 49160 41116
rect 49194 41101 49250 41116
rect 49284 41101 49340 41116
rect 49374 41101 49430 41116
rect 49464 41101 49520 41116
rect 49554 41101 49610 41116
rect 49644 41101 49700 41116
rect 48674 41082 48710 41101
rect 48764 41082 48800 41101
rect 48854 41082 48890 41101
rect 48944 41082 48980 41101
rect 49034 41082 49070 41101
rect 49124 41082 49160 41101
rect 49214 41082 49250 41101
rect 49304 41082 49340 41101
rect 49394 41082 49430 41101
rect 49484 41082 49520 41101
rect 49574 41082 49610 41101
rect 49664 41082 49700 41101
rect 49734 41082 49870 41116
rect 49904 41082 49960 41116
rect 49994 41101 50050 41116
rect 50084 41101 50140 41116
rect 50174 41101 50230 41116
rect 50264 41101 50320 41116
rect 50354 41101 50410 41116
rect 50444 41101 50500 41116
rect 50534 41101 50590 41116
rect 50624 41101 50680 41116
rect 50714 41101 50770 41116
rect 50804 41101 50860 41116
rect 50894 41101 50950 41116
rect 50984 41101 51040 41116
rect 50014 41082 50050 41101
rect 50104 41082 50140 41101
rect 50194 41082 50230 41101
rect 50284 41082 50320 41101
rect 50374 41082 50410 41101
rect 50464 41082 50500 41101
rect 50554 41082 50590 41101
rect 50644 41082 50680 41101
rect 50734 41082 50770 41101
rect 50824 41082 50860 41101
rect 50914 41082 50950 41101
rect 51004 41082 51040 41101
rect 51074 41082 51210 41116
rect 51244 41082 51300 41116
rect 51334 41101 51390 41116
rect 51424 41101 51480 41116
rect 51514 41101 51570 41116
rect 51604 41101 51660 41116
rect 51694 41101 51750 41116
rect 51784 41101 51840 41116
rect 51874 41101 51930 41116
rect 51964 41101 52020 41116
rect 52054 41101 52110 41116
rect 52144 41101 52200 41116
rect 52234 41101 52290 41116
rect 52324 41101 52380 41116
rect 51354 41082 51390 41101
rect 51444 41082 51480 41101
rect 51534 41082 51570 41101
rect 51624 41082 51660 41101
rect 51714 41082 51750 41101
rect 51804 41082 51840 41101
rect 51894 41082 51930 41101
rect 51984 41082 52020 41101
rect 52074 41082 52110 41101
rect 52164 41082 52200 41101
rect 52254 41082 52290 41101
rect 52344 41082 52380 41101
rect 52414 41082 52478 41116
rect 41810 41078 41940 41082
rect 41810 41044 41844 41078
rect 41878 41067 41940 41078
rect 41974 41067 42030 41082
rect 42064 41067 42120 41082
rect 42154 41067 42210 41082
rect 42244 41067 42300 41082
rect 42334 41067 42390 41082
rect 42424 41067 42480 41082
rect 42514 41067 42570 41082
rect 42604 41067 42660 41082
rect 42694 41067 42750 41082
rect 42784 41067 42840 41082
rect 42874 41067 42930 41082
rect 42964 41078 43280 41082
rect 42964 41067 43031 41078
rect 41878 41044 43031 41067
rect 43065 41044 43184 41078
rect 43218 41067 43280 41078
rect 43314 41067 43370 41082
rect 43404 41067 43460 41082
rect 43494 41067 43550 41082
rect 43584 41067 43640 41082
rect 43674 41067 43730 41082
rect 43764 41067 43820 41082
rect 43854 41067 43910 41082
rect 43944 41067 44000 41082
rect 44034 41067 44090 41082
rect 44124 41067 44180 41082
rect 44214 41067 44270 41082
rect 44304 41078 44620 41082
rect 44304 41067 44371 41078
rect 43218 41044 44371 41067
rect 44405 41044 44524 41078
rect 44558 41067 44620 41078
rect 44654 41067 44710 41082
rect 44744 41067 44800 41082
rect 44834 41067 44890 41082
rect 44924 41067 44980 41082
rect 45014 41067 45070 41082
rect 45104 41067 45160 41082
rect 45194 41067 45250 41082
rect 45284 41067 45340 41082
rect 45374 41067 45430 41082
rect 45464 41067 45520 41082
rect 45554 41067 45610 41082
rect 45644 41078 45960 41082
rect 45644 41067 45711 41078
rect 44558 41044 45711 41067
rect 45745 41044 45864 41078
rect 45898 41067 45960 41078
rect 45994 41067 46050 41082
rect 46084 41067 46140 41082
rect 46174 41067 46230 41082
rect 46264 41067 46320 41082
rect 46354 41067 46410 41082
rect 46444 41067 46500 41082
rect 46534 41067 46590 41082
rect 46624 41067 46680 41082
rect 46714 41067 46770 41082
rect 46804 41067 46860 41082
rect 46894 41067 46950 41082
rect 46984 41078 47300 41082
rect 46984 41067 47051 41078
rect 45898 41044 47051 41067
rect 47085 41044 47204 41078
rect 47238 41067 47300 41078
rect 47334 41067 47390 41082
rect 47424 41067 47480 41082
rect 47514 41067 47570 41082
rect 47604 41067 47660 41082
rect 47694 41067 47750 41082
rect 47784 41067 47840 41082
rect 47874 41067 47930 41082
rect 47964 41067 48020 41082
rect 48054 41067 48110 41082
rect 48144 41067 48200 41082
rect 48234 41067 48290 41082
rect 48324 41078 48640 41082
rect 48324 41067 48391 41078
rect 47238 41044 48391 41067
rect 48425 41044 48544 41078
rect 48578 41067 48640 41078
rect 48674 41067 48730 41082
rect 48764 41067 48820 41082
rect 48854 41067 48910 41082
rect 48944 41067 49000 41082
rect 49034 41067 49090 41082
rect 49124 41067 49180 41082
rect 49214 41067 49270 41082
rect 49304 41067 49360 41082
rect 49394 41067 49450 41082
rect 49484 41067 49540 41082
rect 49574 41067 49630 41082
rect 49664 41078 49980 41082
rect 49664 41067 49731 41078
rect 48578 41044 49731 41067
rect 49765 41044 49884 41078
rect 49918 41067 49980 41078
rect 50014 41067 50070 41082
rect 50104 41067 50160 41082
rect 50194 41067 50250 41082
rect 50284 41067 50340 41082
rect 50374 41067 50430 41082
rect 50464 41067 50520 41082
rect 50554 41067 50610 41082
rect 50644 41067 50700 41082
rect 50734 41067 50790 41082
rect 50824 41067 50880 41082
rect 50914 41067 50970 41082
rect 51004 41078 51320 41082
rect 51004 41067 51071 41078
rect 49918 41044 51071 41067
rect 51105 41044 51224 41078
rect 51258 41067 51320 41078
rect 51354 41067 51410 41082
rect 51444 41067 51500 41082
rect 51534 41067 51590 41082
rect 51624 41067 51680 41082
rect 51714 41067 51770 41082
rect 51804 41067 51860 41082
rect 51894 41067 51950 41082
rect 51984 41067 52040 41082
rect 52074 41067 52130 41082
rect 52164 41067 52220 41082
rect 52254 41067 52310 41082
rect 52344 41078 52478 41082
rect 52344 41067 52411 41078
rect 51258 41044 52411 41067
rect 52445 41044 52478 41078
rect 41810 41037 52478 41044
rect 41810 40988 41909 41037
rect 34881 40909 34915 40931
rect 34881 40841 34915 40859
rect 34881 40773 34915 40787
rect 34881 40705 34915 40715
rect 34881 40637 34915 40643
rect 34881 40569 34915 40571
rect 34881 40533 34915 40535
rect 34881 40461 34915 40467
rect 34881 40389 34915 40399
rect 34881 40317 34915 40331
rect 34881 40245 34915 40263
rect 37288 40929 37322 40956
rect 37745 40938 37780 40956
rect 37288 40857 37322 40875
rect 37288 40785 37322 40807
rect 37288 40713 37322 40739
rect 37288 40641 37322 40671
rect 37288 40569 37322 40603
rect 37288 40501 37322 40535
rect 37288 40433 37322 40463
rect 37288 40365 37322 40391
rect 37288 40297 37322 40319
rect 37288 40229 37322 40247
rect 34881 40173 34915 40195
rect 34881 40101 34915 40127
rect 37287 40175 37288 40206
rect 37287 40148 37322 40175
rect 37746 40929 37780 40938
rect 37746 40857 37780 40875
rect 37746 40785 37780 40807
rect 37746 40713 37780 40739
rect 37746 40641 37780 40671
rect 37746 40569 37780 40603
rect 37746 40501 37780 40535
rect 37746 40433 37780 40463
rect 37746 40365 37780 40391
rect 37746 40297 37780 40319
rect 37746 40229 37780 40247
rect 38204 40929 38238 40956
rect 38661 40938 38696 40956
rect 38204 40857 38238 40875
rect 38204 40785 38238 40807
rect 38204 40713 38238 40739
rect 38204 40641 38238 40671
rect 38204 40569 38238 40603
rect 38204 40501 38238 40535
rect 38204 40433 38238 40463
rect 38204 40365 38238 40391
rect 38204 40297 38238 40319
rect 38204 40229 38238 40247
rect 37746 40148 37780 40175
rect 38203 40175 38204 40206
rect 38203 40148 38238 40175
rect 38662 40929 38696 40938
rect 38662 40857 38696 40875
rect 38662 40785 38696 40807
rect 38662 40713 38696 40739
rect 38662 40641 38696 40671
rect 38662 40569 38696 40603
rect 38662 40501 38696 40535
rect 38662 40433 38696 40463
rect 38662 40365 38696 40391
rect 38662 40297 38696 40319
rect 38662 40229 38696 40247
rect 39120 40929 39154 40956
rect 39577 40938 39612 40956
rect 39120 40857 39154 40875
rect 39120 40785 39154 40807
rect 39120 40713 39154 40739
rect 39120 40641 39154 40671
rect 39120 40569 39154 40603
rect 39120 40501 39154 40535
rect 39120 40433 39154 40463
rect 39120 40365 39154 40391
rect 39120 40297 39154 40319
rect 39120 40229 39154 40247
rect 38662 40148 38696 40175
rect 39119 40175 39120 40206
rect 39119 40148 39154 40175
rect 39578 40929 39612 40938
rect 39578 40857 39612 40875
rect 39578 40785 39612 40807
rect 39578 40713 39612 40739
rect 39578 40641 39612 40671
rect 39578 40569 39612 40603
rect 39578 40501 39612 40535
rect 39578 40433 39612 40463
rect 39578 40365 39612 40391
rect 39578 40297 39612 40319
rect 39578 40229 39612 40247
rect 40036 40929 40070 40956
rect 40493 40938 40528 40956
rect 40036 40857 40070 40875
rect 40036 40785 40070 40807
rect 40036 40713 40070 40739
rect 40036 40641 40070 40671
rect 40036 40569 40070 40603
rect 40036 40501 40070 40535
rect 40036 40433 40070 40463
rect 40036 40365 40070 40391
rect 40036 40297 40070 40319
rect 40036 40229 40070 40247
rect 39578 40148 39612 40175
rect 40035 40175 40036 40206
rect 40035 40148 40070 40175
rect 40494 40929 40528 40938
rect 40494 40857 40528 40875
rect 40494 40785 40528 40807
rect 40494 40713 40528 40739
rect 40494 40641 40528 40671
rect 40494 40569 40528 40603
rect 40494 40501 40528 40535
rect 40494 40433 40528 40463
rect 40494 40365 40528 40391
rect 40494 40297 40528 40319
rect 40494 40229 40528 40247
rect 40952 40929 40986 40956
rect 41409 40938 41444 40956
rect 40952 40857 40986 40875
rect 40952 40785 40986 40807
rect 40952 40713 40986 40739
rect 40952 40641 40986 40671
rect 40952 40569 40986 40603
rect 40952 40501 40986 40535
rect 40952 40433 40986 40463
rect 40952 40365 40986 40391
rect 40952 40297 40986 40319
rect 40952 40229 40986 40247
rect 40494 40148 40528 40175
rect 40951 40175 40952 40206
rect 40951 40148 40986 40175
rect 41410 40929 41444 40938
rect 41410 40857 41444 40875
rect 41410 40785 41444 40807
rect 41410 40713 41444 40739
rect 41410 40641 41444 40671
rect 41410 40569 41444 40603
rect 41410 40501 41444 40535
rect 41410 40433 41444 40463
rect 41410 40365 41444 40391
rect 41410 40297 41444 40319
rect 41410 40229 41444 40247
rect 41410 40148 41444 40175
rect 41810 40954 41844 40988
rect 41878 40954 41909 40988
rect 42999 40988 43249 41037
rect 41810 40898 41909 40954
rect 41810 40864 41844 40898
rect 41878 40864 41909 40898
rect 41810 40808 41909 40864
rect 41810 40774 41844 40808
rect 41878 40774 41909 40808
rect 41810 40718 41909 40774
rect 41810 40684 41844 40718
rect 41878 40684 41909 40718
rect 41810 40628 41909 40684
rect 41810 40594 41844 40628
rect 41878 40594 41909 40628
rect 41810 40538 41909 40594
rect 41810 40504 41844 40538
rect 41878 40504 41909 40538
rect 41810 40448 41909 40504
rect 41810 40414 41844 40448
rect 41878 40414 41909 40448
rect 41810 40358 41909 40414
rect 41810 40324 41844 40358
rect 41878 40324 41909 40358
rect 41810 40268 41909 40324
rect 41810 40234 41844 40268
rect 41878 40234 41909 40268
rect 41810 40178 41909 40234
rect 37287 40082 37321 40148
rect 38203 40082 38237 40148
rect 39119 40082 39153 40148
rect 40035 40082 40069 40148
rect 40951 40082 40985 40148
rect 41810 40144 41844 40178
rect 41878 40144 41909 40178
rect 41810 40088 41909 40144
rect 34881 40029 34915 40059
rect 37276 40022 41456 40082
rect 41810 40054 41844 40088
rect 41878 40054 41909 40088
rect 34881 39957 34915 39991
rect 34881 39822 34915 39923
rect 41810 39998 41909 40054
rect 41973 40956 42935 40973
rect 41973 40922 41994 40956
rect 42028 40922 42084 40956
rect 42118 40954 42174 40956
rect 42208 40954 42264 40956
rect 42298 40954 42354 40956
rect 42388 40954 42444 40956
rect 42478 40954 42534 40956
rect 42568 40954 42624 40956
rect 42658 40954 42714 40956
rect 42748 40954 42804 40956
rect 42838 40954 42894 40956
rect 42138 40922 42174 40954
rect 42228 40922 42264 40954
rect 42318 40922 42354 40954
rect 42408 40922 42444 40954
rect 42498 40922 42534 40954
rect 42588 40922 42624 40954
rect 42678 40922 42714 40954
rect 42768 40922 42804 40954
rect 42858 40922 42894 40954
rect 42928 40922 42935 40956
rect 41973 40920 42104 40922
rect 42138 40920 42194 40922
rect 42228 40920 42284 40922
rect 42318 40920 42374 40922
rect 42408 40920 42464 40922
rect 42498 40920 42554 40922
rect 42588 40920 42644 40922
rect 42678 40920 42734 40922
rect 42768 40920 42824 40922
rect 42858 40920 42935 40922
rect 41973 40901 42935 40920
rect 41973 40897 42045 40901
rect 41973 40863 41992 40897
rect 42026 40863 42045 40897
rect 41973 40807 42045 40863
rect 42863 40878 42935 40901
rect 42863 40844 42882 40878
rect 42916 40844 42935 40878
rect 41973 40773 41992 40807
rect 42026 40773 42045 40807
rect 41973 40717 42045 40773
rect 41973 40683 41992 40717
rect 42026 40683 42045 40717
rect 41973 40627 42045 40683
rect 41973 40593 41992 40627
rect 42026 40593 42045 40627
rect 41973 40537 42045 40593
rect 41973 40503 41992 40537
rect 42026 40503 42045 40537
rect 41973 40447 42045 40503
rect 41973 40413 41992 40447
rect 42026 40413 42045 40447
rect 41973 40357 42045 40413
rect 41973 40323 41992 40357
rect 42026 40323 42045 40357
rect 41973 40267 42045 40323
rect 41973 40233 41992 40267
rect 42026 40233 42045 40267
rect 41973 40177 42045 40233
rect 41973 40143 41992 40177
rect 42026 40143 42045 40177
rect 42107 40780 42801 40839
rect 42107 40746 42168 40780
rect 42202 40752 42258 40780
rect 42292 40752 42348 40780
rect 42382 40752 42438 40780
rect 42214 40746 42258 40752
rect 42314 40746 42348 40752
rect 42414 40746 42438 40752
rect 42472 40752 42528 40780
rect 42472 40746 42480 40752
rect 42107 40718 42180 40746
rect 42214 40718 42280 40746
rect 42314 40718 42380 40746
rect 42414 40718 42480 40746
rect 42514 40746 42528 40752
rect 42562 40752 42618 40780
rect 42562 40746 42580 40752
rect 42514 40718 42580 40746
rect 42614 40746 42618 40752
rect 42652 40752 42708 40780
rect 42652 40746 42680 40752
rect 42742 40746 42801 40780
rect 42614 40718 42680 40746
rect 42714 40718 42801 40746
rect 42107 40690 42801 40718
rect 42107 40656 42168 40690
rect 42202 40656 42258 40690
rect 42292 40656 42348 40690
rect 42382 40656 42438 40690
rect 42472 40656 42528 40690
rect 42562 40656 42618 40690
rect 42652 40656 42708 40690
rect 42742 40656 42801 40690
rect 42107 40652 42801 40656
rect 42107 40618 42180 40652
rect 42214 40618 42280 40652
rect 42314 40618 42380 40652
rect 42414 40618 42480 40652
rect 42514 40618 42580 40652
rect 42614 40618 42680 40652
rect 42714 40618 42801 40652
rect 42107 40600 42801 40618
rect 42107 40566 42168 40600
rect 42202 40566 42258 40600
rect 42292 40566 42348 40600
rect 42382 40566 42438 40600
rect 42472 40566 42528 40600
rect 42562 40566 42618 40600
rect 42652 40566 42708 40600
rect 42742 40566 42801 40600
rect 42107 40552 42801 40566
rect 42107 40518 42180 40552
rect 42214 40518 42280 40552
rect 42314 40518 42380 40552
rect 42414 40518 42480 40552
rect 42514 40518 42580 40552
rect 42614 40518 42680 40552
rect 42714 40518 42801 40552
rect 42107 40510 42801 40518
rect 42107 40476 42168 40510
rect 42202 40476 42258 40510
rect 42292 40476 42348 40510
rect 42382 40476 42438 40510
rect 42472 40476 42528 40510
rect 42562 40476 42618 40510
rect 42652 40476 42708 40510
rect 42742 40476 42801 40510
rect 42107 40452 42801 40476
rect 42107 40420 42180 40452
rect 42214 40420 42280 40452
rect 42314 40420 42380 40452
rect 42414 40420 42480 40452
rect 42107 40386 42168 40420
rect 42214 40418 42258 40420
rect 42314 40418 42348 40420
rect 42414 40418 42438 40420
rect 42202 40386 42258 40418
rect 42292 40386 42348 40418
rect 42382 40386 42438 40418
rect 42472 40418 42480 40420
rect 42514 40420 42580 40452
rect 42514 40418 42528 40420
rect 42472 40386 42528 40418
rect 42562 40418 42580 40420
rect 42614 40420 42680 40452
rect 42714 40420 42801 40452
rect 42614 40418 42618 40420
rect 42562 40386 42618 40418
rect 42652 40418 42680 40420
rect 42652 40386 42708 40418
rect 42742 40386 42801 40420
rect 42107 40352 42801 40386
rect 42107 40330 42180 40352
rect 42214 40330 42280 40352
rect 42314 40330 42380 40352
rect 42414 40330 42480 40352
rect 42107 40296 42168 40330
rect 42214 40318 42258 40330
rect 42314 40318 42348 40330
rect 42414 40318 42438 40330
rect 42202 40296 42258 40318
rect 42292 40296 42348 40318
rect 42382 40296 42438 40318
rect 42472 40318 42480 40330
rect 42514 40330 42580 40352
rect 42514 40318 42528 40330
rect 42472 40296 42528 40318
rect 42562 40318 42580 40330
rect 42614 40330 42680 40352
rect 42714 40330 42801 40352
rect 42614 40318 42618 40330
rect 42562 40296 42618 40318
rect 42652 40318 42680 40330
rect 42652 40296 42708 40318
rect 42742 40296 42801 40330
rect 42107 40252 42801 40296
rect 42107 40240 42180 40252
rect 42214 40240 42280 40252
rect 42314 40240 42380 40252
rect 42414 40240 42480 40252
rect 42107 40206 42168 40240
rect 42214 40218 42258 40240
rect 42314 40218 42348 40240
rect 42414 40218 42438 40240
rect 42202 40206 42258 40218
rect 42292 40206 42348 40218
rect 42382 40206 42438 40218
rect 42472 40218 42480 40240
rect 42514 40240 42580 40252
rect 42514 40218 42528 40240
rect 42472 40206 42528 40218
rect 42562 40218 42580 40240
rect 42614 40240 42680 40252
rect 42714 40240 42801 40252
rect 42614 40218 42618 40240
rect 42562 40206 42618 40218
rect 42652 40218 42680 40240
rect 42652 40206 42708 40218
rect 42742 40206 42801 40240
rect 42107 40145 42801 40206
rect 42863 40788 42935 40844
rect 42863 40754 42882 40788
rect 42916 40754 42935 40788
rect 42863 40698 42935 40754
rect 42863 40664 42882 40698
rect 42916 40664 42935 40698
rect 42863 40608 42935 40664
rect 42863 40574 42882 40608
rect 42916 40574 42935 40608
rect 42863 40518 42935 40574
rect 42863 40484 42882 40518
rect 42916 40484 42935 40518
rect 42863 40428 42935 40484
rect 42863 40394 42882 40428
rect 42916 40394 42935 40428
rect 42863 40338 42935 40394
rect 42863 40304 42882 40338
rect 42916 40304 42935 40338
rect 42863 40248 42935 40304
rect 42863 40214 42882 40248
rect 42916 40214 42935 40248
rect 42863 40158 42935 40214
rect 41973 40083 42045 40143
rect 42863 40124 42882 40158
rect 42916 40124 42935 40158
rect 42863 40083 42935 40124
rect 41973 40064 42935 40083
rect 41973 40030 42070 40064
rect 42104 40030 42160 40064
rect 42194 40030 42250 40064
rect 42284 40030 42340 40064
rect 42374 40030 42430 40064
rect 42464 40030 42520 40064
rect 42554 40030 42610 40064
rect 42644 40030 42700 40064
rect 42734 40030 42790 40064
rect 42824 40030 42935 40064
rect 41973 40011 42935 40030
rect 42999 40954 43031 40988
rect 43065 40954 43184 40988
rect 43218 40954 43249 40988
rect 44339 40988 44589 41037
rect 42999 40898 43249 40954
rect 42999 40864 43031 40898
rect 43065 40864 43184 40898
rect 43218 40864 43249 40898
rect 42999 40808 43249 40864
rect 42999 40774 43031 40808
rect 43065 40774 43184 40808
rect 43218 40774 43249 40808
rect 42999 40718 43249 40774
rect 42999 40684 43031 40718
rect 43065 40684 43184 40718
rect 43218 40684 43249 40718
rect 42999 40628 43249 40684
rect 42999 40594 43031 40628
rect 43065 40594 43184 40628
rect 43218 40594 43249 40628
rect 42999 40538 43249 40594
rect 42999 40504 43031 40538
rect 43065 40504 43184 40538
rect 43218 40504 43249 40538
rect 42999 40448 43249 40504
rect 42999 40414 43031 40448
rect 43065 40414 43184 40448
rect 43218 40414 43249 40448
rect 42999 40358 43249 40414
rect 42999 40324 43031 40358
rect 43065 40324 43184 40358
rect 43218 40324 43249 40358
rect 42999 40268 43249 40324
rect 42999 40234 43031 40268
rect 43065 40234 43184 40268
rect 43218 40234 43249 40268
rect 42999 40178 43249 40234
rect 42999 40144 43031 40178
rect 43065 40144 43184 40178
rect 43218 40144 43249 40178
rect 42999 40088 43249 40144
rect 42999 40054 43031 40088
rect 43065 40054 43184 40088
rect 43218 40054 43249 40088
rect 41810 39964 41844 39998
rect 41878 39964 41909 39998
rect 41810 39947 41909 39964
rect 42999 39998 43249 40054
rect 43313 40956 44275 40973
rect 43313 40922 43334 40956
rect 43368 40922 43424 40956
rect 43458 40954 43514 40956
rect 43548 40954 43604 40956
rect 43638 40954 43694 40956
rect 43728 40954 43784 40956
rect 43818 40954 43874 40956
rect 43908 40954 43964 40956
rect 43998 40954 44054 40956
rect 44088 40954 44144 40956
rect 44178 40954 44234 40956
rect 43478 40922 43514 40954
rect 43568 40922 43604 40954
rect 43658 40922 43694 40954
rect 43748 40922 43784 40954
rect 43838 40922 43874 40954
rect 43928 40922 43964 40954
rect 44018 40922 44054 40954
rect 44108 40922 44144 40954
rect 44198 40922 44234 40954
rect 44268 40922 44275 40956
rect 43313 40920 43444 40922
rect 43478 40920 43534 40922
rect 43568 40920 43624 40922
rect 43658 40920 43714 40922
rect 43748 40920 43804 40922
rect 43838 40920 43894 40922
rect 43928 40920 43984 40922
rect 44018 40920 44074 40922
rect 44108 40920 44164 40922
rect 44198 40920 44275 40922
rect 43313 40901 44275 40920
rect 43313 40897 43385 40901
rect 43313 40863 43332 40897
rect 43366 40863 43385 40897
rect 43313 40807 43385 40863
rect 44203 40878 44275 40901
rect 44203 40844 44222 40878
rect 44256 40844 44275 40878
rect 43313 40773 43332 40807
rect 43366 40773 43385 40807
rect 43313 40717 43385 40773
rect 43313 40683 43332 40717
rect 43366 40683 43385 40717
rect 43313 40627 43385 40683
rect 43313 40593 43332 40627
rect 43366 40593 43385 40627
rect 43313 40537 43385 40593
rect 43313 40503 43332 40537
rect 43366 40503 43385 40537
rect 43313 40447 43385 40503
rect 43313 40413 43332 40447
rect 43366 40413 43385 40447
rect 43313 40357 43385 40413
rect 43313 40323 43332 40357
rect 43366 40323 43385 40357
rect 43313 40267 43385 40323
rect 43313 40233 43332 40267
rect 43366 40233 43385 40267
rect 43313 40177 43385 40233
rect 43313 40143 43332 40177
rect 43366 40143 43385 40177
rect 43447 40780 44141 40839
rect 43447 40746 43508 40780
rect 43542 40752 43598 40780
rect 43632 40752 43688 40780
rect 43722 40752 43778 40780
rect 43554 40746 43598 40752
rect 43654 40746 43688 40752
rect 43754 40746 43778 40752
rect 43812 40752 43868 40780
rect 43812 40746 43820 40752
rect 43447 40718 43520 40746
rect 43554 40718 43620 40746
rect 43654 40718 43720 40746
rect 43754 40718 43820 40746
rect 43854 40746 43868 40752
rect 43902 40752 43958 40780
rect 43902 40746 43920 40752
rect 43854 40718 43920 40746
rect 43954 40746 43958 40752
rect 43992 40752 44048 40780
rect 43992 40746 44020 40752
rect 44082 40746 44141 40780
rect 43954 40718 44020 40746
rect 44054 40718 44141 40746
rect 43447 40690 44141 40718
rect 43447 40656 43508 40690
rect 43542 40656 43598 40690
rect 43632 40656 43688 40690
rect 43722 40656 43778 40690
rect 43812 40656 43868 40690
rect 43902 40656 43958 40690
rect 43992 40656 44048 40690
rect 44082 40656 44141 40690
rect 43447 40652 44141 40656
rect 43447 40618 43520 40652
rect 43554 40618 43620 40652
rect 43654 40618 43720 40652
rect 43754 40618 43820 40652
rect 43854 40618 43920 40652
rect 43954 40618 44020 40652
rect 44054 40618 44141 40652
rect 43447 40600 44141 40618
rect 43447 40566 43508 40600
rect 43542 40566 43598 40600
rect 43632 40566 43688 40600
rect 43722 40566 43778 40600
rect 43812 40566 43868 40600
rect 43902 40566 43958 40600
rect 43992 40566 44048 40600
rect 44082 40566 44141 40600
rect 43447 40552 44141 40566
rect 43447 40518 43520 40552
rect 43554 40518 43620 40552
rect 43654 40518 43720 40552
rect 43754 40518 43820 40552
rect 43854 40518 43920 40552
rect 43954 40518 44020 40552
rect 44054 40518 44141 40552
rect 43447 40510 44141 40518
rect 43447 40476 43508 40510
rect 43542 40476 43598 40510
rect 43632 40476 43688 40510
rect 43722 40476 43778 40510
rect 43812 40476 43868 40510
rect 43902 40476 43958 40510
rect 43992 40476 44048 40510
rect 44082 40476 44141 40510
rect 43447 40452 44141 40476
rect 43447 40420 43520 40452
rect 43554 40420 43620 40452
rect 43654 40420 43720 40452
rect 43754 40420 43820 40452
rect 43447 40386 43508 40420
rect 43554 40418 43598 40420
rect 43654 40418 43688 40420
rect 43754 40418 43778 40420
rect 43542 40386 43598 40418
rect 43632 40386 43688 40418
rect 43722 40386 43778 40418
rect 43812 40418 43820 40420
rect 43854 40420 43920 40452
rect 43854 40418 43868 40420
rect 43812 40386 43868 40418
rect 43902 40418 43920 40420
rect 43954 40420 44020 40452
rect 44054 40420 44141 40452
rect 43954 40418 43958 40420
rect 43902 40386 43958 40418
rect 43992 40418 44020 40420
rect 43992 40386 44048 40418
rect 44082 40386 44141 40420
rect 43447 40352 44141 40386
rect 43447 40330 43520 40352
rect 43554 40330 43620 40352
rect 43654 40330 43720 40352
rect 43754 40330 43820 40352
rect 43447 40296 43508 40330
rect 43554 40318 43598 40330
rect 43654 40318 43688 40330
rect 43754 40318 43778 40330
rect 43542 40296 43598 40318
rect 43632 40296 43688 40318
rect 43722 40296 43778 40318
rect 43812 40318 43820 40330
rect 43854 40330 43920 40352
rect 43854 40318 43868 40330
rect 43812 40296 43868 40318
rect 43902 40318 43920 40330
rect 43954 40330 44020 40352
rect 44054 40330 44141 40352
rect 43954 40318 43958 40330
rect 43902 40296 43958 40318
rect 43992 40318 44020 40330
rect 43992 40296 44048 40318
rect 44082 40296 44141 40330
rect 43447 40252 44141 40296
rect 43447 40240 43520 40252
rect 43554 40240 43620 40252
rect 43654 40240 43720 40252
rect 43754 40240 43820 40252
rect 43447 40206 43508 40240
rect 43554 40218 43598 40240
rect 43654 40218 43688 40240
rect 43754 40218 43778 40240
rect 43542 40206 43598 40218
rect 43632 40206 43688 40218
rect 43722 40206 43778 40218
rect 43812 40218 43820 40240
rect 43854 40240 43920 40252
rect 43854 40218 43868 40240
rect 43812 40206 43868 40218
rect 43902 40218 43920 40240
rect 43954 40240 44020 40252
rect 44054 40240 44141 40252
rect 43954 40218 43958 40240
rect 43902 40206 43958 40218
rect 43992 40218 44020 40240
rect 43992 40206 44048 40218
rect 44082 40206 44141 40240
rect 43447 40145 44141 40206
rect 44203 40788 44275 40844
rect 44203 40754 44222 40788
rect 44256 40754 44275 40788
rect 44203 40698 44275 40754
rect 44203 40664 44222 40698
rect 44256 40664 44275 40698
rect 44203 40608 44275 40664
rect 44203 40574 44222 40608
rect 44256 40574 44275 40608
rect 44203 40518 44275 40574
rect 44203 40484 44222 40518
rect 44256 40484 44275 40518
rect 44203 40428 44275 40484
rect 44203 40394 44222 40428
rect 44256 40394 44275 40428
rect 44203 40338 44275 40394
rect 44203 40304 44222 40338
rect 44256 40304 44275 40338
rect 44203 40248 44275 40304
rect 44203 40214 44222 40248
rect 44256 40214 44275 40248
rect 44203 40158 44275 40214
rect 43313 40083 43385 40143
rect 44203 40124 44222 40158
rect 44256 40124 44275 40158
rect 44203 40083 44275 40124
rect 43313 40064 44275 40083
rect 43313 40030 43410 40064
rect 43444 40030 43500 40064
rect 43534 40030 43590 40064
rect 43624 40030 43680 40064
rect 43714 40030 43770 40064
rect 43804 40030 43860 40064
rect 43894 40030 43950 40064
rect 43984 40030 44040 40064
rect 44074 40030 44130 40064
rect 44164 40030 44275 40064
rect 43313 40011 44275 40030
rect 44339 40954 44371 40988
rect 44405 40954 44524 40988
rect 44558 40954 44589 40988
rect 45679 40988 45929 41037
rect 44339 40898 44589 40954
rect 44339 40864 44371 40898
rect 44405 40864 44524 40898
rect 44558 40864 44589 40898
rect 44339 40808 44589 40864
rect 44339 40774 44371 40808
rect 44405 40774 44524 40808
rect 44558 40774 44589 40808
rect 44339 40718 44589 40774
rect 44339 40684 44371 40718
rect 44405 40684 44524 40718
rect 44558 40684 44589 40718
rect 44339 40628 44589 40684
rect 44339 40594 44371 40628
rect 44405 40594 44524 40628
rect 44558 40594 44589 40628
rect 44339 40538 44589 40594
rect 44339 40504 44371 40538
rect 44405 40504 44524 40538
rect 44558 40504 44589 40538
rect 44339 40448 44589 40504
rect 44339 40414 44371 40448
rect 44405 40414 44524 40448
rect 44558 40414 44589 40448
rect 44339 40358 44589 40414
rect 44339 40324 44371 40358
rect 44405 40324 44524 40358
rect 44558 40324 44589 40358
rect 44339 40268 44589 40324
rect 44339 40234 44371 40268
rect 44405 40234 44524 40268
rect 44558 40234 44589 40268
rect 44339 40178 44589 40234
rect 44339 40144 44371 40178
rect 44405 40144 44524 40178
rect 44558 40144 44589 40178
rect 44339 40088 44589 40144
rect 44339 40054 44371 40088
rect 44405 40054 44524 40088
rect 44558 40054 44589 40088
rect 42999 39964 43031 39998
rect 43065 39964 43184 39998
rect 43218 39964 43249 39998
rect 42999 39947 43249 39964
rect 44339 39998 44589 40054
rect 44653 40956 45615 40973
rect 44653 40922 44674 40956
rect 44708 40922 44764 40956
rect 44798 40954 44854 40956
rect 44888 40954 44944 40956
rect 44978 40954 45034 40956
rect 45068 40954 45124 40956
rect 45158 40954 45214 40956
rect 45248 40954 45304 40956
rect 45338 40954 45394 40956
rect 45428 40954 45484 40956
rect 45518 40954 45574 40956
rect 44818 40922 44854 40954
rect 44908 40922 44944 40954
rect 44998 40922 45034 40954
rect 45088 40922 45124 40954
rect 45178 40922 45214 40954
rect 45268 40922 45304 40954
rect 45358 40922 45394 40954
rect 45448 40922 45484 40954
rect 45538 40922 45574 40954
rect 45608 40922 45615 40956
rect 44653 40920 44784 40922
rect 44818 40920 44874 40922
rect 44908 40920 44964 40922
rect 44998 40920 45054 40922
rect 45088 40920 45144 40922
rect 45178 40920 45234 40922
rect 45268 40920 45324 40922
rect 45358 40920 45414 40922
rect 45448 40920 45504 40922
rect 45538 40920 45615 40922
rect 44653 40901 45615 40920
rect 44653 40897 44725 40901
rect 44653 40863 44672 40897
rect 44706 40863 44725 40897
rect 44653 40807 44725 40863
rect 45543 40878 45615 40901
rect 45543 40844 45562 40878
rect 45596 40844 45615 40878
rect 44653 40773 44672 40807
rect 44706 40773 44725 40807
rect 44653 40717 44725 40773
rect 44653 40683 44672 40717
rect 44706 40683 44725 40717
rect 44653 40627 44725 40683
rect 44653 40593 44672 40627
rect 44706 40593 44725 40627
rect 44653 40537 44725 40593
rect 44653 40503 44672 40537
rect 44706 40503 44725 40537
rect 44653 40447 44725 40503
rect 44653 40413 44672 40447
rect 44706 40413 44725 40447
rect 44653 40357 44725 40413
rect 44653 40323 44672 40357
rect 44706 40323 44725 40357
rect 44653 40267 44725 40323
rect 44653 40233 44672 40267
rect 44706 40233 44725 40267
rect 44653 40177 44725 40233
rect 44653 40143 44672 40177
rect 44706 40143 44725 40177
rect 44787 40780 45481 40839
rect 44787 40746 44848 40780
rect 44882 40752 44938 40780
rect 44972 40752 45028 40780
rect 45062 40752 45118 40780
rect 44894 40746 44938 40752
rect 44994 40746 45028 40752
rect 45094 40746 45118 40752
rect 45152 40752 45208 40780
rect 45152 40746 45160 40752
rect 44787 40718 44860 40746
rect 44894 40718 44960 40746
rect 44994 40718 45060 40746
rect 45094 40718 45160 40746
rect 45194 40746 45208 40752
rect 45242 40752 45298 40780
rect 45242 40746 45260 40752
rect 45194 40718 45260 40746
rect 45294 40746 45298 40752
rect 45332 40752 45388 40780
rect 45332 40746 45360 40752
rect 45422 40746 45481 40780
rect 45294 40718 45360 40746
rect 45394 40718 45481 40746
rect 44787 40690 45481 40718
rect 44787 40656 44848 40690
rect 44882 40656 44938 40690
rect 44972 40656 45028 40690
rect 45062 40656 45118 40690
rect 45152 40656 45208 40690
rect 45242 40656 45298 40690
rect 45332 40656 45388 40690
rect 45422 40656 45481 40690
rect 44787 40652 45481 40656
rect 44787 40618 44860 40652
rect 44894 40618 44960 40652
rect 44994 40618 45060 40652
rect 45094 40618 45160 40652
rect 45194 40618 45260 40652
rect 45294 40618 45360 40652
rect 45394 40618 45481 40652
rect 44787 40600 45481 40618
rect 44787 40566 44848 40600
rect 44882 40566 44938 40600
rect 44972 40566 45028 40600
rect 45062 40566 45118 40600
rect 45152 40566 45208 40600
rect 45242 40566 45298 40600
rect 45332 40566 45388 40600
rect 45422 40566 45481 40600
rect 44787 40552 45481 40566
rect 44787 40518 44860 40552
rect 44894 40518 44960 40552
rect 44994 40518 45060 40552
rect 45094 40518 45160 40552
rect 45194 40518 45260 40552
rect 45294 40518 45360 40552
rect 45394 40518 45481 40552
rect 44787 40510 45481 40518
rect 44787 40476 44848 40510
rect 44882 40476 44938 40510
rect 44972 40476 45028 40510
rect 45062 40476 45118 40510
rect 45152 40476 45208 40510
rect 45242 40476 45298 40510
rect 45332 40476 45388 40510
rect 45422 40476 45481 40510
rect 44787 40452 45481 40476
rect 44787 40420 44860 40452
rect 44894 40420 44960 40452
rect 44994 40420 45060 40452
rect 45094 40420 45160 40452
rect 44787 40386 44848 40420
rect 44894 40418 44938 40420
rect 44994 40418 45028 40420
rect 45094 40418 45118 40420
rect 44882 40386 44938 40418
rect 44972 40386 45028 40418
rect 45062 40386 45118 40418
rect 45152 40418 45160 40420
rect 45194 40420 45260 40452
rect 45194 40418 45208 40420
rect 45152 40386 45208 40418
rect 45242 40418 45260 40420
rect 45294 40420 45360 40452
rect 45394 40420 45481 40452
rect 45294 40418 45298 40420
rect 45242 40386 45298 40418
rect 45332 40418 45360 40420
rect 45332 40386 45388 40418
rect 45422 40386 45481 40420
rect 44787 40352 45481 40386
rect 44787 40330 44860 40352
rect 44894 40330 44960 40352
rect 44994 40330 45060 40352
rect 45094 40330 45160 40352
rect 44787 40296 44848 40330
rect 44894 40318 44938 40330
rect 44994 40318 45028 40330
rect 45094 40318 45118 40330
rect 44882 40296 44938 40318
rect 44972 40296 45028 40318
rect 45062 40296 45118 40318
rect 45152 40318 45160 40330
rect 45194 40330 45260 40352
rect 45194 40318 45208 40330
rect 45152 40296 45208 40318
rect 45242 40318 45260 40330
rect 45294 40330 45360 40352
rect 45394 40330 45481 40352
rect 45294 40318 45298 40330
rect 45242 40296 45298 40318
rect 45332 40318 45360 40330
rect 45332 40296 45388 40318
rect 45422 40296 45481 40330
rect 44787 40252 45481 40296
rect 44787 40240 44860 40252
rect 44894 40240 44960 40252
rect 44994 40240 45060 40252
rect 45094 40240 45160 40252
rect 44787 40206 44848 40240
rect 44894 40218 44938 40240
rect 44994 40218 45028 40240
rect 45094 40218 45118 40240
rect 44882 40206 44938 40218
rect 44972 40206 45028 40218
rect 45062 40206 45118 40218
rect 45152 40218 45160 40240
rect 45194 40240 45260 40252
rect 45194 40218 45208 40240
rect 45152 40206 45208 40218
rect 45242 40218 45260 40240
rect 45294 40240 45360 40252
rect 45394 40240 45481 40252
rect 45294 40218 45298 40240
rect 45242 40206 45298 40218
rect 45332 40218 45360 40240
rect 45332 40206 45388 40218
rect 45422 40206 45481 40240
rect 44787 40145 45481 40206
rect 45543 40788 45615 40844
rect 45543 40754 45562 40788
rect 45596 40754 45615 40788
rect 45543 40698 45615 40754
rect 45543 40664 45562 40698
rect 45596 40664 45615 40698
rect 45543 40608 45615 40664
rect 45543 40574 45562 40608
rect 45596 40574 45615 40608
rect 45543 40518 45615 40574
rect 45543 40484 45562 40518
rect 45596 40484 45615 40518
rect 45543 40428 45615 40484
rect 45543 40394 45562 40428
rect 45596 40394 45615 40428
rect 45543 40338 45615 40394
rect 45543 40304 45562 40338
rect 45596 40304 45615 40338
rect 45543 40248 45615 40304
rect 45543 40214 45562 40248
rect 45596 40214 45615 40248
rect 45543 40158 45615 40214
rect 44653 40083 44725 40143
rect 45543 40124 45562 40158
rect 45596 40124 45615 40158
rect 45543 40083 45615 40124
rect 44653 40064 45615 40083
rect 44653 40030 44750 40064
rect 44784 40030 44840 40064
rect 44874 40030 44930 40064
rect 44964 40030 45020 40064
rect 45054 40030 45110 40064
rect 45144 40030 45200 40064
rect 45234 40030 45290 40064
rect 45324 40030 45380 40064
rect 45414 40030 45470 40064
rect 45504 40030 45615 40064
rect 44653 40011 45615 40030
rect 45679 40954 45711 40988
rect 45745 40954 45864 40988
rect 45898 40954 45929 40988
rect 47019 40988 47269 41037
rect 45679 40898 45929 40954
rect 45679 40864 45711 40898
rect 45745 40864 45864 40898
rect 45898 40864 45929 40898
rect 45679 40808 45929 40864
rect 45679 40774 45711 40808
rect 45745 40774 45864 40808
rect 45898 40774 45929 40808
rect 45679 40718 45929 40774
rect 45679 40684 45711 40718
rect 45745 40684 45864 40718
rect 45898 40684 45929 40718
rect 45679 40628 45929 40684
rect 45679 40594 45711 40628
rect 45745 40594 45864 40628
rect 45898 40594 45929 40628
rect 45679 40538 45929 40594
rect 45679 40504 45711 40538
rect 45745 40504 45864 40538
rect 45898 40504 45929 40538
rect 45679 40448 45929 40504
rect 45679 40414 45711 40448
rect 45745 40414 45864 40448
rect 45898 40414 45929 40448
rect 45679 40358 45929 40414
rect 45679 40324 45711 40358
rect 45745 40324 45864 40358
rect 45898 40324 45929 40358
rect 45679 40268 45929 40324
rect 45679 40234 45711 40268
rect 45745 40234 45864 40268
rect 45898 40234 45929 40268
rect 45679 40178 45929 40234
rect 45679 40144 45711 40178
rect 45745 40144 45864 40178
rect 45898 40144 45929 40178
rect 45679 40088 45929 40144
rect 45679 40054 45711 40088
rect 45745 40054 45864 40088
rect 45898 40054 45929 40088
rect 44339 39964 44371 39998
rect 44405 39964 44524 39998
rect 44558 39964 44589 39998
rect 44339 39947 44589 39964
rect 45679 39998 45929 40054
rect 45993 40956 46955 40973
rect 45993 40922 46014 40956
rect 46048 40922 46104 40956
rect 46138 40954 46194 40956
rect 46228 40954 46284 40956
rect 46318 40954 46374 40956
rect 46408 40954 46464 40956
rect 46498 40954 46554 40956
rect 46588 40954 46644 40956
rect 46678 40954 46734 40956
rect 46768 40954 46824 40956
rect 46858 40954 46914 40956
rect 46158 40922 46194 40954
rect 46248 40922 46284 40954
rect 46338 40922 46374 40954
rect 46428 40922 46464 40954
rect 46518 40922 46554 40954
rect 46608 40922 46644 40954
rect 46698 40922 46734 40954
rect 46788 40922 46824 40954
rect 46878 40922 46914 40954
rect 46948 40922 46955 40956
rect 45993 40920 46124 40922
rect 46158 40920 46214 40922
rect 46248 40920 46304 40922
rect 46338 40920 46394 40922
rect 46428 40920 46484 40922
rect 46518 40920 46574 40922
rect 46608 40920 46664 40922
rect 46698 40920 46754 40922
rect 46788 40920 46844 40922
rect 46878 40920 46955 40922
rect 45993 40901 46955 40920
rect 45993 40897 46065 40901
rect 45993 40863 46012 40897
rect 46046 40863 46065 40897
rect 45993 40807 46065 40863
rect 46883 40878 46955 40901
rect 46883 40844 46902 40878
rect 46936 40844 46955 40878
rect 45993 40773 46012 40807
rect 46046 40773 46065 40807
rect 45993 40717 46065 40773
rect 45993 40683 46012 40717
rect 46046 40683 46065 40717
rect 45993 40627 46065 40683
rect 45993 40593 46012 40627
rect 46046 40593 46065 40627
rect 45993 40537 46065 40593
rect 45993 40503 46012 40537
rect 46046 40503 46065 40537
rect 45993 40447 46065 40503
rect 45993 40413 46012 40447
rect 46046 40413 46065 40447
rect 45993 40357 46065 40413
rect 45993 40323 46012 40357
rect 46046 40323 46065 40357
rect 45993 40267 46065 40323
rect 45993 40233 46012 40267
rect 46046 40233 46065 40267
rect 45993 40177 46065 40233
rect 45993 40143 46012 40177
rect 46046 40143 46065 40177
rect 46127 40780 46821 40839
rect 46127 40746 46188 40780
rect 46222 40752 46278 40780
rect 46312 40752 46368 40780
rect 46402 40752 46458 40780
rect 46234 40746 46278 40752
rect 46334 40746 46368 40752
rect 46434 40746 46458 40752
rect 46492 40752 46548 40780
rect 46492 40746 46500 40752
rect 46127 40718 46200 40746
rect 46234 40718 46300 40746
rect 46334 40718 46400 40746
rect 46434 40718 46500 40746
rect 46534 40746 46548 40752
rect 46582 40752 46638 40780
rect 46582 40746 46600 40752
rect 46534 40718 46600 40746
rect 46634 40746 46638 40752
rect 46672 40752 46728 40780
rect 46672 40746 46700 40752
rect 46762 40746 46821 40780
rect 46634 40718 46700 40746
rect 46734 40718 46821 40746
rect 46127 40690 46821 40718
rect 46127 40656 46188 40690
rect 46222 40656 46278 40690
rect 46312 40656 46368 40690
rect 46402 40656 46458 40690
rect 46492 40656 46548 40690
rect 46582 40656 46638 40690
rect 46672 40656 46728 40690
rect 46762 40656 46821 40690
rect 46127 40652 46821 40656
rect 46127 40618 46200 40652
rect 46234 40618 46300 40652
rect 46334 40618 46400 40652
rect 46434 40618 46500 40652
rect 46534 40618 46600 40652
rect 46634 40618 46700 40652
rect 46734 40618 46821 40652
rect 46127 40600 46821 40618
rect 46127 40566 46188 40600
rect 46222 40566 46278 40600
rect 46312 40566 46368 40600
rect 46402 40566 46458 40600
rect 46492 40566 46548 40600
rect 46582 40566 46638 40600
rect 46672 40566 46728 40600
rect 46762 40566 46821 40600
rect 46127 40552 46821 40566
rect 46127 40518 46200 40552
rect 46234 40518 46300 40552
rect 46334 40518 46400 40552
rect 46434 40518 46500 40552
rect 46534 40518 46600 40552
rect 46634 40518 46700 40552
rect 46734 40518 46821 40552
rect 46127 40510 46821 40518
rect 46127 40476 46188 40510
rect 46222 40476 46278 40510
rect 46312 40476 46368 40510
rect 46402 40476 46458 40510
rect 46492 40476 46548 40510
rect 46582 40476 46638 40510
rect 46672 40476 46728 40510
rect 46762 40476 46821 40510
rect 46127 40452 46821 40476
rect 46127 40420 46200 40452
rect 46234 40420 46300 40452
rect 46334 40420 46400 40452
rect 46434 40420 46500 40452
rect 46127 40386 46188 40420
rect 46234 40418 46278 40420
rect 46334 40418 46368 40420
rect 46434 40418 46458 40420
rect 46222 40386 46278 40418
rect 46312 40386 46368 40418
rect 46402 40386 46458 40418
rect 46492 40418 46500 40420
rect 46534 40420 46600 40452
rect 46534 40418 46548 40420
rect 46492 40386 46548 40418
rect 46582 40418 46600 40420
rect 46634 40420 46700 40452
rect 46734 40420 46821 40452
rect 46634 40418 46638 40420
rect 46582 40386 46638 40418
rect 46672 40418 46700 40420
rect 46672 40386 46728 40418
rect 46762 40386 46821 40420
rect 46127 40352 46821 40386
rect 46127 40330 46200 40352
rect 46234 40330 46300 40352
rect 46334 40330 46400 40352
rect 46434 40330 46500 40352
rect 46127 40296 46188 40330
rect 46234 40318 46278 40330
rect 46334 40318 46368 40330
rect 46434 40318 46458 40330
rect 46222 40296 46278 40318
rect 46312 40296 46368 40318
rect 46402 40296 46458 40318
rect 46492 40318 46500 40330
rect 46534 40330 46600 40352
rect 46534 40318 46548 40330
rect 46492 40296 46548 40318
rect 46582 40318 46600 40330
rect 46634 40330 46700 40352
rect 46734 40330 46821 40352
rect 46634 40318 46638 40330
rect 46582 40296 46638 40318
rect 46672 40318 46700 40330
rect 46672 40296 46728 40318
rect 46762 40296 46821 40330
rect 46127 40252 46821 40296
rect 46127 40240 46200 40252
rect 46234 40240 46300 40252
rect 46334 40240 46400 40252
rect 46434 40240 46500 40252
rect 46127 40206 46188 40240
rect 46234 40218 46278 40240
rect 46334 40218 46368 40240
rect 46434 40218 46458 40240
rect 46222 40206 46278 40218
rect 46312 40206 46368 40218
rect 46402 40206 46458 40218
rect 46492 40218 46500 40240
rect 46534 40240 46600 40252
rect 46534 40218 46548 40240
rect 46492 40206 46548 40218
rect 46582 40218 46600 40240
rect 46634 40240 46700 40252
rect 46734 40240 46821 40252
rect 46634 40218 46638 40240
rect 46582 40206 46638 40218
rect 46672 40218 46700 40240
rect 46672 40206 46728 40218
rect 46762 40206 46821 40240
rect 46127 40145 46821 40206
rect 46883 40788 46955 40844
rect 46883 40754 46902 40788
rect 46936 40754 46955 40788
rect 46883 40698 46955 40754
rect 46883 40664 46902 40698
rect 46936 40664 46955 40698
rect 46883 40608 46955 40664
rect 46883 40574 46902 40608
rect 46936 40574 46955 40608
rect 46883 40518 46955 40574
rect 46883 40484 46902 40518
rect 46936 40484 46955 40518
rect 46883 40428 46955 40484
rect 46883 40394 46902 40428
rect 46936 40394 46955 40428
rect 46883 40338 46955 40394
rect 46883 40304 46902 40338
rect 46936 40304 46955 40338
rect 46883 40248 46955 40304
rect 46883 40214 46902 40248
rect 46936 40214 46955 40248
rect 46883 40158 46955 40214
rect 45993 40083 46065 40143
rect 46883 40124 46902 40158
rect 46936 40124 46955 40158
rect 46883 40083 46955 40124
rect 45993 40064 46955 40083
rect 45993 40030 46090 40064
rect 46124 40030 46180 40064
rect 46214 40030 46270 40064
rect 46304 40030 46360 40064
rect 46394 40030 46450 40064
rect 46484 40030 46540 40064
rect 46574 40030 46630 40064
rect 46664 40030 46720 40064
rect 46754 40030 46810 40064
rect 46844 40030 46955 40064
rect 45993 40011 46955 40030
rect 47019 40954 47051 40988
rect 47085 40954 47204 40988
rect 47238 40954 47269 40988
rect 48359 40988 48609 41037
rect 47019 40898 47269 40954
rect 47019 40864 47051 40898
rect 47085 40864 47204 40898
rect 47238 40864 47269 40898
rect 47019 40808 47269 40864
rect 47019 40774 47051 40808
rect 47085 40774 47204 40808
rect 47238 40774 47269 40808
rect 47019 40718 47269 40774
rect 47019 40684 47051 40718
rect 47085 40684 47204 40718
rect 47238 40684 47269 40718
rect 47019 40628 47269 40684
rect 47019 40594 47051 40628
rect 47085 40594 47204 40628
rect 47238 40594 47269 40628
rect 47019 40538 47269 40594
rect 47019 40504 47051 40538
rect 47085 40504 47204 40538
rect 47238 40504 47269 40538
rect 47019 40448 47269 40504
rect 47019 40414 47051 40448
rect 47085 40414 47204 40448
rect 47238 40414 47269 40448
rect 47019 40358 47269 40414
rect 47019 40324 47051 40358
rect 47085 40324 47204 40358
rect 47238 40324 47269 40358
rect 47019 40268 47269 40324
rect 47019 40234 47051 40268
rect 47085 40234 47204 40268
rect 47238 40234 47269 40268
rect 47019 40178 47269 40234
rect 47019 40144 47051 40178
rect 47085 40144 47204 40178
rect 47238 40144 47269 40178
rect 47019 40088 47269 40144
rect 47019 40054 47051 40088
rect 47085 40054 47204 40088
rect 47238 40054 47269 40088
rect 45679 39964 45711 39998
rect 45745 39964 45864 39998
rect 45898 39964 45929 39998
rect 45679 39947 45929 39964
rect 47019 39998 47269 40054
rect 47333 40956 48295 40973
rect 47333 40922 47354 40956
rect 47388 40922 47444 40956
rect 47478 40954 47534 40956
rect 47568 40954 47624 40956
rect 47658 40954 47714 40956
rect 47748 40954 47804 40956
rect 47838 40954 47894 40956
rect 47928 40954 47984 40956
rect 48018 40954 48074 40956
rect 48108 40954 48164 40956
rect 48198 40954 48254 40956
rect 47498 40922 47534 40954
rect 47588 40922 47624 40954
rect 47678 40922 47714 40954
rect 47768 40922 47804 40954
rect 47858 40922 47894 40954
rect 47948 40922 47984 40954
rect 48038 40922 48074 40954
rect 48128 40922 48164 40954
rect 48218 40922 48254 40954
rect 48288 40922 48295 40956
rect 47333 40920 47464 40922
rect 47498 40920 47554 40922
rect 47588 40920 47644 40922
rect 47678 40920 47734 40922
rect 47768 40920 47824 40922
rect 47858 40920 47914 40922
rect 47948 40920 48004 40922
rect 48038 40920 48094 40922
rect 48128 40920 48184 40922
rect 48218 40920 48295 40922
rect 47333 40901 48295 40920
rect 47333 40897 47405 40901
rect 47333 40863 47352 40897
rect 47386 40863 47405 40897
rect 47333 40807 47405 40863
rect 48223 40878 48295 40901
rect 48223 40844 48242 40878
rect 48276 40844 48295 40878
rect 47333 40773 47352 40807
rect 47386 40773 47405 40807
rect 47333 40717 47405 40773
rect 47333 40683 47352 40717
rect 47386 40683 47405 40717
rect 47333 40627 47405 40683
rect 47333 40593 47352 40627
rect 47386 40593 47405 40627
rect 47333 40537 47405 40593
rect 47333 40503 47352 40537
rect 47386 40503 47405 40537
rect 47333 40447 47405 40503
rect 47333 40413 47352 40447
rect 47386 40413 47405 40447
rect 47333 40357 47405 40413
rect 47333 40323 47352 40357
rect 47386 40323 47405 40357
rect 47333 40267 47405 40323
rect 47333 40233 47352 40267
rect 47386 40233 47405 40267
rect 47333 40177 47405 40233
rect 47333 40143 47352 40177
rect 47386 40143 47405 40177
rect 47467 40780 48161 40839
rect 47467 40746 47528 40780
rect 47562 40752 47618 40780
rect 47652 40752 47708 40780
rect 47742 40752 47798 40780
rect 47574 40746 47618 40752
rect 47674 40746 47708 40752
rect 47774 40746 47798 40752
rect 47832 40752 47888 40780
rect 47832 40746 47840 40752
rect 47467 40718 47540 40746
rect 47574 40718 47640 40746
rect 47674 40718 47740 40746
rect 47774 40718 47840 40746
rect 47874 40746 47888 40752
rect 47922 40752 47978 40780
rect 47922 40746 47940 40752
rect 47874 40718 47940 40746
rect 47974 40746 47978 40752
rect 48012 40752 48068 40780
rect 48012 40746 48040 40752
rect 48102 40746 48161 40780
rect 47974 40718 48040 40746
rect 48074 40718 48161 40746
rect 47467 40690 48161 40718
rect 47467 40656 47528 40690
rect 47562 40656 47618 40690
rect 47652 40656 47708 40690
rect 47742 40656 47798 40690
rect 47832 40656 47888 40690
rect 47922 40656 47978 40690
rect 48012 40656 48068 40690
rect 48102 40656 48161 40690
rect 47467 40652 48161 40656
rect 47467 40618 47540 40652
rect 47574 40618 47640 40652
rect 47674 40618 47740 40652
rect 47774 40618 47840 40652
rect 47874 40618 47940 40652
rect 47974 40618 48040 40652
rect 48074 40618 48161 40652
rect 47467 40600 48161 40618
rect 47467 40566 47528 40600
rect 47562 40566 47618 40600
rect 47652 40566 47708 40600
rect 47742 40566 47798 40600
rect 47832 40566 47888 40600
rect 47922 40566 47978 40600
rect 48012 40566 48068 40600
rect 48102 40566 48161 40600
rect 47467 40552 48161 40566
rect 47467 40518 47540 40552
rect 47574 40518 47640 40552
rect 47674 40518 47740 40552
rect 47774 40518 47840 40552
rect 47874 40518 47940 40552
rect 47974 40518 48040 40552
rect 48074 40518 48161 40552
rect 47467 40510 48161 40518
rect 47467 40476 47528 40510
rect 47562 40476 47618 40510
rect 47652 40476 47708 40510
rect 47742 40476 47798 40510
rect 47832 40476 47888 40510
rect 47922 40476 47978 40510
rect 48012 40476 48068 40510
rect 48102 40476 48161 40510
rect 47467 40452 48161 40476
rect 47467 40420 47540 40452
rect 47574 40420 47640 40452
rect 47674 40420 47740 40452
rect 47774 40420 47840 40452
rect 47467 40386 47528 40420
rect 47574 40418 47618 40420
rect 47674 40418 47708 40420
rect 47774 40418 47798 40420
rect 47562 40386 47618 40418
rect 47652 40386 47708 40418
rect 47742 40386 47798 40418
rect 47832 40418 47840 40420
rect 47874 40420 47940 40452
rect 47874 40418 47888 40420
rect 47832 40386 47888 40418
rect 47922 40418 47940 40420
rect 47974 40420 48040 40452
rect 48074 40420 48161 40452
rect 47974 40418 47978 40420
rect 47922 40386 47978 40418
rect 48012 40418 48040 40420
rect 48012 40386 48068 40418
rect 48102 40386 48161 40420
rect 47467 40352 48161 40386
rect 47467 40330 47540 40352
rect 47574 40330 47640 40352
rect 47674 40330 47740 40352
rect 47774 40330 47840 40352
rect 47467 40296 47528 40330
rect 47574 40318 47618 40330
rect 47674 40318 47708 40330
rect 47774 40318 47798 40330
rect 47562 40296 47618 40318
rect 47652 40296 47708 40318
rect 47742 40296 47798 40318
rect 47832 40318 47840 40330
rect 47874 40330 47940 40352
rect 47874 40318 47888 40330
rect 47832 40296 47888 40318
rect 47922 40318 47940 40330
rect 47974 40330 48040 40352
rect 48074 40330 48161 40352
rect 47974 40318 47978 40330
rect 47922 40296 47978 40318
rect 48012 40318 48040 40330
rect 48012 40296 48068 40318
rect 48102 40296 48161 40330
rect 47467 40252 48161 40296
rect 47467 40240 47540 40252
rect 47574 40240 47640 40252
rect 47674 40240 47740 40252
rect 47774 40240 47840 40252
rect 47467 40206 47528 40240
rect 47574 40218 47618 40240
rect 47674 40218 47708 40240
rect 47774 40218 47798 40240
rect 47562 40206 47618 40218
rect 47652 40206 47708 40218
rect 47742 40206 47798 40218
rect 47832 40218 47840 40240
rect 47874 40240 47940 40252
rect 47874 40218 47888 40240
rect 47832 40206 47888 40218
rect 47922 40218 47940 40240
rect 47974 40240 48040 40252
rect 48074 40240 48161 40252
rect 47974 40218 47978 40240
rect 47922 40206 47978 40218
rect 48012 40218 48040 40240
rect 48012 40206 48068 40218
rect 48102 40206 48161 40240
rect 47467 40145 48161 40206
rect 48223 40788 48295 40844
rect 48223 40754 48242 40788
rect 48276 40754 48295 40788
rect 48223 40698 48295 40754
rect 48223 40664 48242 40698
rect 48276 40664 48295 40698
rect 48223 40608 48295 40664
rect 48223 40574 48242 40608
rect 48276 40574 48295 40608
rect 48223 40518 48295 40574
rect 48223 40484 48242 40518
rect 48276 40484 48295 40518
rect 48223 40428 48295 40484
rect 48223 40394 48242 40428
rect 48276 40394 48295 40428
rect 48223 40338 48295 40394
rect 48223 40304 48242 40338
rect 48276 40304 48295 40338
rect 48223 40248 48295 40304
rect 48223 40214 48242 40248
rect 48276 40214 48295 40248
rect 48223 40158 48295 40214
rect 47333 40083 47405 40143
rect 48223 40124 48242 40158
rect 48276 40124 48295 40158
rect 48223 40083 48295 40124
rect 47333 40064 48295 40083
rect 47333 40030 47430 40064
rect 47464 40030 47520 40064
rect 47554 40030 47610 40064
rect 47644 40030 47700 40064
rect 47734 40030 47790 40064
rect 47824 40030 47880 40064
rect 47914 40030 47970 40064
rect 48004 40030 48060 40064
rect 48094 40030 48150 40064
rect 48184 40030 48295 40064
rect 47333 40011 48295 40030
rect 48359 40954 48391 40988
rect 48425 40954 48544 40988
rect 48578 40954 48609 40988
rect 49699 40988 49949 41037
rect 48359 40898 48609 40954
rect 48359 40864 48391 40898
rect 48425 40864 48544 40898
rect 48578 40864 48609 40898
rect 48359 40808 48609 40864
rect 48359 40774 48391 40808
rect 48425 40774 48544 40808
rect 48578 40774 48609 40808
rect 48359 40718 48609 40774
rect 48359 40684 48391 40718
rect 48425 40684 48544 40718
rect 48578 40684 48609 40718
rect 48359 40628 48609 40684
rect 48359 40594 48391 40628
rect 48425 40594 48544 40628
rect 48578 40594 48609 40628
rect 48359 40538 48609 40594
rect 48359 40504 48391 40538
rect 48425 40504 48544 40538
rect 48578 40504 48609 40538
rect 48359 40448 48609 40504
rect 48359 40414 48391 40448
rect 48425 40414 48544 40448
rect 48578 40414 48609 40448
rect 48359 40358 48609 40414
rect 48359 40324 48391 40358
rect 48425 40324 48544 40358
rect 48578 40324 48609 40358
rect 48359 40268 48609 40324
rect 48359 40234 48391 40268
rect 48425 40234 48544 40268
rect 48578 40234 48609 40268
rect 48359 40178 48609 40234
rect 48359 40144 48391 40178
rect 48425 40144 48544 40178
rect 48578 40144 48609 40178
rect 48359 40088 48609 40144
rect 48359 40054 48391 40088
rect 48425 40054 48544 40088
rect 48578 40054 48609 40088
rect 47019 39964 47051 39998
rect 47085 39964 47204 39998
rect 47238 39964 47269 39998
rect 47019 39947 47269 39964
rect 48359 39998 48609 40054
rect 48673 40956 49635 40973
rect 48673 40922 48694 40956
rect 48728 40922 48784 40956
rect 48818 40954 48874 40956
rect 48908 40954 48964 40956
rect 48998 40954 49054 40956
rect 49088 40954 49144 40956
rect 49178 40954 49234 40956
rect 49268 40954 49324 40956
rect 49358 40954 49414 40956
rect 49448 40954 49504 40956
rect 49538 40954 49594 40956
rect 48838 40922 48874 40954
rect 48928 40922 48964 40954
rect 49018 40922 49054 40954
rect 49108 40922 49144 40954
rect 49198 40922 49234 40954
rect 49288 40922 49324 40954
rect 49378 40922 49414 40954
rect 49468 40922 49504 40954
rect 49558 40922 49594 40954
rect 49628 40922 49635 40956
rect 48673 40920 48804 40922
rect 48838 40920 48894 40922
rect 48928 40920 48984 40922
rect 49018 40920 49074 40922
rect 49108 40920 49164 40922
rect 49198 40920 49254 40922
rect 49288 40920 49344 40922
rect 49378 40920 49434 40922
rect 49468 40920 49524 40922
rect 49558 40920 49635 40922
rect 48673 40901 49635 40920
rect 48673 40897 48745 40901
rect 48673 40863 48692 40897
rect 48726 40863 48745 40897
rect 48673 40807 48745 40863
rect 49563 40878 49635 40901
rect 49563 40844 49582 40878
rect 49616 40844 49635 40878
rect 48673 40773 48692 40807
rect 48726 40773 48745 40807
rect 48673 40717 48745 40773
rect 48673 40683 48692 40717
rect 48726 40683 48745 40717
rect 48673 40627 48745 40683
rect 48673 40593 48692 40627
rect 48726 40593 48745 40627
rect 48673 40537 48745 40593
rect 48673 40503 48692 40537
rect 48726 40503 48745 40537
rect 48673 40447 48745 40503
rect 48673 40413 48692 40447
rect 48726 40413 48745 40447
rect 48673 40357 48745 40413
rect 48673 40323 48692 40357
rect 48726 40323 48745 40357
rect 48673 40267 48745 40323
rect 48673 40233 48692 40267
rect 48726 40233 48745 40267
rect 48673 40177 48745 40233
rect 48673 40143 48692 40177
rect 48726 40143 48745 40177
rect 48807 40780 49501 40839
rect 48807 40746 48868 40780
rect 48902 40752 48958 40780
rect 48992 40752 49048 40780
rect 49082 40752 49138 40780
rect 48914 40746 48958 40752
rect 49014 40746 49048 40752
rect 49114 40746 49138 40752
rect 49172 40752 49228 40780
rect 49172 40746 49180 40752
rect 48807 40718 48880 40746
rect 48914 40718 48980 40746
rect 49014 40718 49080 40746
rect 49114 40718 49180 40746
rect 49214 40746 49228 40752
rect 49262 40752 49318 40780
rect 49262 40746 49280 40752
rect 49214 40718 49280 40746
rect 49314 40746 49318 40752
rect 49352 40752 49408 40780
rect 49352 40746 49380 40752
rect 49442 40746 49501 40780
rect 49314 40718 49380 40746
rect 49414 40718 49501 40746
rect 48807 40690 49501 40718
rect 48807 40656 48868 40690
rect 48902 40656 48958 40690
rect 48992 40656 49048 40690
rect 49082 40656 49138 40690
rect 49172 40656 49228 40690
rect 49262 40656 49318 40690
rect 49352 40656 49408 40690
rect 49442 40656 49501 40690
rect 48807 40652 49501 40656
rect 48807 40618 48880 40652
rect 48914 40618 48980 40652
rect 49014 40618 49080 40652
rect 49114 40618 49180 40652
rect 49214 40618 49280 40652
rect 49314 40618 49380 40652
rect 49414 40618 49501 40652
rect 48807 40600 49501 40618
rect 48807 40566 48868 40600
rect 48902 40566 48958 40600
rect 48992 40566 49048 40600
rect 49082 40566 49138 40600
rect 49172 40566 49228 40600
rect 49262 40566 49318 40600
rect 49352 40566 49408 40600
rect 49442 40566 49501 40600
rect 48807 40552 49501 40566
rect 48807 40518 48880 40552
rect 48914 40518 48980 40552
rect 49014 40518 49080 40552
rect 49114 40518 49180 40552
rect 49214 40518 49280 40552
rect 49314 40518 49380 40552
rect 49414 40518 49501 40552
rect 48807 40510 49501 40518
rect 48807 40476 48868 40510
rect 48902 40476 48958 40510
rect 48992 40476 49048 40510
rect 49082 40476 49138 40510
rect 49172 40476 49228 40510
rect 49262 40476 49318 40510
rect 49352 40476 49408 40510
rect 49442 40476 49501 40510
rect 48807 40452 49501 40476
rect 48807 40420 48880 40452
rect 48914 40420 48980 40452
rect 49014 40420 49080 40452
rect 49114 40420 49180 40452
rect 48807 40386 48868 40420
rect 48914 40418 48958 40420
rect 49014 40418 49048 40420
rect 49114 40418 49138 40420
rect 48902 40386 48958 40418
rect 48992 40386 49048 40418
rect 49082 40386 49138 40418
rect 49172 40418 49180 40420
rect 49214 40420 49280 40452
rect 49214 40418 49228 40420
rect 49172 40386 49228 40418
rect 49262 40418 49280 40420
rect 49314 40420 49380 40452
rect 49414 40420 49501 40452
rect 49314 40418 49318 40420
rect 49262 40386 49318 40418
rect 49352 40418 49380 40420
rect 49352 40386 49408 40418
rect 49442 40386 49501 40420
rect 48807 40352 49501 40386
rect 48807 40330 48880 40352
rect 48914 40330 48980 40352
rect 49014 40330 49080 40352
rect 49114 40330 49180 40352
rect 48807 40296 48868 40330
rect 48914 40318 48958 40330
rect 49014 40318 49048 40330
rect 49114 40318 49138 40330
rect 48902 40296 48958 40318
rect 48992 40296 49048 40318
rect 49082 40296 49138 40318
rect 49172 40318 49180 40330
rect 49214 40330 49280 40352
rect 49214 40318 49228 40330
rect 49172 40296 49228 40318
rect 49262 40318 49280 40330
rect 49314 40330 49380 40352
rect 49414 40330 49501 40352
rect 49314 40318 49318 40330
rect 49262 40296 49318 40318
rect 49352 40318 49380 40330
rect 49352 40296 49408 40318
rect 49442 40296 49501 40330
rect 48807 40252 49501 40296
rect 48807 40240 48880 40252
rect 48914 40240 48980 40252
rect 49014 40240 49080 40252
rect 49114 40240 49180 40252
rect 48807 40206 48868 40240
rect 48914 40218 48958 40240
rect 49014 40218 49048 40240
rect 49114 40218 49138 40240
rect 48902 40206 48958 40218
rect 48992 40206 49048 40218
rect 49082 40206 49138 40218
rect 49172 40218 49180 40240
rect 49214 40240 49280 40252
rect 49214 40218 49228 40240
rect 49172 40206 49228 40218
rect 49262 40218 49280 40240
rect 49314 40240 49380 40252
rect 49414 40240 49501 40252
rect 49314 40218 49318 40240
rect 49262 40206 49318 40218
rect 49352 40218 49380 40240
rect 49352 40206 49408 40218
rect 49442 40206 49501 40240
rect 48807 40145 49501 40206
rect 49563 40788 49635 40844
rect 49563 40754 49582 40788
rect 49616 40754 49635 40788
rect 49563 40698 49635 40754
rect 49563 40664 49582 40698
rect 49616 40664 49635 40698
rect 49563 40608 49635 40664
rect 49563 40574 49582 40608
rect 49616 40574 49635 40608
rect 49563 40518 49635 40574
rect 49563 40484 49582 40518
rect 49616 40484 49635 40518
rect 49563 40428 49635 40484
rect 49563 40394 49582 40428
rect 49616 40394 49635 40428
rect 49563 40338 49635 40394
rect 49563 40304 49582 40338
rect 49616 40304 49635 40338
rect 49563 40248 49635 40304
rect 49563 40214 49582 40248
rect 49616 40214 49635 40248
rect 49563 40158 49635 40214
rect 48673 40083 48745 40143
rect 49563 40124 49582 40158
rect 49616 40124 49635 40158
rect 49563 40083 49635 40124
rect 48673 40064 49635 40083
rect 48673 40030 48770 40064
rect 48804 40030 48860 40064
rect 48894 40030 48950 40064
rect 48984 40030 49040 40064
rect 49074 40030 49130 40064
rect 49164 40030 49220 40064
rect 49254 40030 49310 40064
rect 49344 40030 49400 40064
rect 49434 40030 49490 40064
rect 49524 40030 49635 40064
rect 48673 40011 49635 40030
rect 49699 40954 49731 40988
rect 49765 40954 49884 40988
rect 49918 40954 49949 40988
rect 51039 40988 51289 41037
rect 49699 40898 49949 40954
rect 49699 40864 49731 40898
rect 49765 40864 49884 40898
rect 49918 40864 49949 40898
rect 49699 40808 49949 40864
rect 49699 40774 49731 40808
rect 49765 40774 49884 40808
rect 49918 40774 49949 40808
rect 49699 40718 49949 40774
rect 49699 40684 49731 40718
rect 49765 40684 49884 40718
rect 49918 40684 49949 40718
rect 49699 40628 49949 40684
rect 49699 40594 49731 40628
rect 49765 40594 49884 40628
rect 49918 40594 49949 40628
rect 49699 40538 49949 40594
rect 49699 40504 49731 40538
rect 49765 40504 49884 40538
rect 49918 40504 49949 40538
rect 49699 40448 49949 40504
rect 49699 40414 49731 40448
rect 49765 40414 49884 40448
rect 49918 40414 49949 40448
rect 49699 40358 49949 40414
rect 49699 40324 49731 40358
rect 49765 40324 49884 40358
rect 49918 40324 49949 40358
rect 49699 40268 49949 40324
rect 49699 40234 49731 40268
rect 49765 40234 49884 40268
rect 49918 40234 49949 40268
rect 49699 40178 49949 40234
rect 49699 40144 49731 40178
rect 49765 40144 49884 40178
rect 49918 40144 49949 40178
rect 49699 40088 49949 40144
rect 49699 40054 49731 40088
rect 49765 40054 49884 40088
rect 49918 40054 49949 40088
rect 48359 39964 48391 39998
rect 48425 39964 48544 39998
rect 48578 39964 48609 39998
rect 48359 39947 48609 39964
rect 49699 39998 49949 40054
rect 50013 40956 50975 40973
rect 50013 40922 50034 40956
rect 50068 40922 50124 40956
rect 50158 40954 50214 40956
rect 50248 40954 50304 40956
rect 50338 40954 50394 40956
rect 50428 40954 50484 40956
rect 50518 40954 50574 40956
rect 50608 40954 50664 40956
rect 50698 40954 50754 40956
rect 50788 40954 50844 40956
rect 50878 40954 50934 40956
rect 50178 40922 50214 40954
rect 50268 40922 50304 40954
rect 50358 40922 50394 40954
rect 50448 40922 50484 40954
rect 50538 40922 50574 40954
rect 50628 40922 50664 40954
rect 50718 40922 50754 40954
rect 50808 40922 50844 40954
rect 50898 40922 50934 40954
rect 50968 40922 50975 40956
rect 50013 40920 50144 40922
rect 50178 40920 50234 40922
rect 50268 40920 50324 40922
rect 50358 40920 50414 40922
rect 50448 40920 50504 40922
rect 50538 40920 50594 40922
rect 50628 40920 50684 40922
rect 50718 40920 50774 40922
rect 50808 40920 50864 40922
rect 50898 40920 50975 40922
rect 50013 40901 50975 40920
rect 50013 40897 50085 40901
rect 50013 40863 50032 40897
rect 50066 40863 50085 40897
rect 50013 40807 50085 40863
rect 50903 40878 50975 40901
rect 50903 40844 50922 40878
rect 50956 40844 50975 40878
rect 50013 40773 50032 40807
rect 50066 40773 50085 40807
rect 50013 40717 50085 40773
rect 50013 40683 50032 40717
rect 50066 40683 50085 40717
rect 50013 40627 50085 40683
rect 50013 40593 50032 40627
rect 50066 40593 50085 40627
rect 50013 40537 50085 40593
rect 50013 40503 50032 40537
rect 50066 40503 50085 40537
rect 50013 40447 50085 40503
rect 50013 40413 50032 40447
rect 50066 40413 50085 40447
rect 50013 40357 50085 40413
rect 50013 40323 50032 40357
rect 50066 40323 50085 40357
rect 50013 40267 50085 40323
rect 50013 40233 50032 40267
rect 50066 40233 50085 40267
rect 50013 40177 50085 40233
rect 50013 40143 50032 40177
rect 50066 40143 50085 40177
rect 50147 40780 50841 40839
rect 50147 40746 50208 40780
rect 50242 40752 50298 40780
rect 50332 40752 50388 40780
rect 50422 40752 50478 40780
rect 50254 40746 50298 40752
rect 50354 40746 50388 40752
rect 50454 40746 50478 40752
rect 50512 40752 50568 40780
rect 50512 40746 50520 40752
rect 50147 40718 50220 40746
rect 50254 40718 50320 40746
rect 50354 40718 50420 40746
rect 50454 40718 50520 40746
rect 50554 40746 50568 40752
rect 50602 40752 50658 40780
rect 50602 40746 50620 40752
rect 50554 40718 50620 40746
rect 50654 40746 50658 40752
rect 50692 40752 50748 40780
rect 50692 40746 50720 40752
rect 50782 40746 50841 40780
rect 50654 40718 50720 40746
rect 50754 40718 50841 40746
rect 50147 40690 50841 40718
rect 50147 40656 50208 40690
rect 50242 40656 50298 40690
rect 50332 40656 50388 40690
rect 50422 40656 50478 40690
rect 50512 40656 50568 40690
rect 50602 40656 50658 40690
rect 50692 40656 50748 40690
rect 50782 40656 50841 40690
rect 50147 40652 50841 40656
rect 50147 40618 50220 40652
rect 50254 40618 50320 40652
rect 50354 40618 50420 40652
rect 50454 40618 50520 40652
rect 50554 40618 50620 40652
rect 50654 40618 50720 40652
rect 50754 40618 50841 40652
rect 50147 40600 50841 40618
rect 50147 40566 50208 40600
rect 50242 40566 50298 40600
rect 50332 40566 50388 40600
rect 50422 40566 50478 40600
rect 50512 40566 50568 40600
rect 50602 40566 50658 40600
rect 50692 40566 50748 40600
rect 50782 40566 50841 40600
rect 50147 40552 50841 40566
rect 50147 40518 50220 40552
rect 50254 40518 50320 40552
rect 50354 40518 50420 40552
rect 50454 40518 50520 40552
rect 50554 40518 50620 40552
rect 50654 40518 50720 40552
rect 50754 40518 50841 40552
rect 50147 40510 50841 40518
rect 50147 40476 50208 40510
rect 50242 40476 50298 40510
rect 50332 40476 50388 40510
rect 50422 40476 50478 40510
rect 50512 40476 50568 40510
rect 50602 40476 50658 40510
rect 50692 40476 50748 40510
rect 50782 40476 50841 40510
rect 50147 40452 50841 40476
rect 50147 40420 50220 40452
rect 50254 40420 50320 40452
rect 50354 40420 50420 40452
rect 50454 40420 50520 40452
rect 50147 40386 50208 40420
rect 50254 40418 50298 40420
rect 50354 40418 50388 40420
rect 50454 40418 50478 40420
rect 50242 40386 50298 40418
rect 50332 40386 50388 40418
rect 50422 40386 50478 40418
rect 50512 40418 50520 40420
rect 50554 40420 50620 40452
rect 50554 40418 50568 40420
rect 50512 40386 50568 40418
rect 50602 40418 50620 40420
rect 50654 40420 50720 40452
rect 50754 40420 50841 40452
rect 50654 40418 50658 40420
rect 50602 40386 50658 40418
rect 50692 40418 50720 40420
rect 50692 40386 50748 40418
rect 50782 40386 50841 40420
rect 50147 40352 50841 40386
rect 50147 40330 50220 40352
rect 50254 40330 50320 40352
rect 50354 40330 50420 40352
rect 50454 40330 50520 40352
rect 50147 40296 50208 40330
rect 50254 40318 50298 40330
rect 50354 40318 50388 40330
rect 50454 40318 50478 40330
rect 50242 40296 50298 40318
rect 50332 40296 50388 40318
rect 50422 40296 50478 40318
rect 50512 40318 50520 40330
rect 50554 40330 50620 40352
rect 50554 40318 50568 40330
rect 50512 40296 50568 40318
rect 50602 40318 50620 40330
rect 50654 40330 50720 40352
rect 50754 40330 50841 40352
rect 50654 40318 50658 40330
rect 50602 40296 50658 40318
rect 50692 40318 50720 40330
rect 50692 40296 50748 40318
rect 50782 40296 50841 40330
rect 50147 40252 50841 40296
rect 50147 40240 50220 40252
rect 50254 40240 50320 40252
rect 50354 40240 50420 40252
rect 50454 40240 50520 40252
rect 50147 40206 50208 40240
rect 50254 40218 50298 40240
rect 50354 40218 50388 40240
rect 50454 40218 50478 40240
rect 50242 40206 50298 40218
rect 50332 40206 50388 40218
rect 50422 40206 50478 40218
rect 50512 40218 50520 40240
rect 50554 40240 50620 40252
rect 50554 40218 50568 40240
rect 50512 40206 50568 40218
rect 50602 40218 50620 40240
rect 50654 40240 50720 40252
rect 50754 40240 50841 40252
rect 50654 40218 50658 40240
rect 50602 40206 50658 40218
rect 50692 40218 50720 40240
rect 50692 40206 50748 40218
rect 50782 40206 50841 40240
rect 50147 40145 50841 40206
rect 50903 40788 50975 40844
rect 50903 40754 50922 40788
rect 50956 40754 50975 40788
rect 50903 40698 50975 40754
rect 50903 40664 50922 40698
rect 50956 40664 50975 40698
rect 50903 40608 50975 40664
rect 50903 40574 50922 40608
rect 50956 40574 50975 40608
rect 50903 40518 50975 40574
rect 50903 40484 50922 40518
rect 50956 40484 50975 40518
rect 50903 40428 50975 40484
rect 50903 40394 50922 40428
rect 50956 40394 50975 40428
rect 50903 40338 50975 40394
rect 50903 40304 50922 40338
rect 50956 40304 50975 40338
rect 50903 40248 50975 40304
rect 50903 40214 50922 40248
rect 50956 40214 50975 40248
rect 50903 40158 50975 40214
rect 50013 40083 50085 40143
rect 50903 40124 50922 40158
rect 50956 40124 50975 40158
rect 50903 40083 50975 40124
rect 50013 40064 50975 40083
rect 50013 40030 50110 40064
rect 50144 40030 50200 40064
rect 50234 40030 50290 40064
rect 50324 40030 50380 40064
rect 50414 40030 50470 40064
rect 50504 40030 50560 40064
rect 50594 40030 50650 40064
rect 50684 40030 50740 40064
rect 50774 40030 50830 40064
rect 50864 40030 50975 40064
rect 50013 40011 50975 40030
rect 51039 40954 51071 40988
rect 51105 40954 51224 40988
rect 51258 40954 51289 40988
rect 52379 40988 52478 41037
rect 51039 40898 51289 40954
rect 51039 40864 51071 40898
rect 51105 40864 51224 40898
rect 51258 40864 51289 40898
rect 51039 40808 51289 40864
rect 51039 40774 51071 40808
rect 51105 40774 51224 40808
rect 51258 40774 51289 40808
rect 51039 40718 51289 40774
rect 51039 40684 51071 40718
rect 51105 40684 51224 40718
rect 51258 40684 51289 40718
rect 51039 40628 51289 40684
rect 51039 40594 51071 40628
rect 51105 40594 51224 40628
rect 51258 40594 51289 40628
rect 51039 40538 51289 40594
rect 51039 40504 51071 40538
rect 51105 40504 51224 40538
rect 51258 40504 51289 40538
rect 51039 40448 51289 40504
rect 51039 40414 51071 40448
rect 51105 40414 51224 40448
rect 51258 40414 51289 40448
rect 51039 40358 51289 40414
rect 51039 40324 51071 40358
rect 51105 40324 51224 40358
rect 51258 40324 51289 40358
rect 51039 40268 51289 40324
rect 51039 40234 51071 40268
rect 51105 40234 51224 40268
rect 51258 40234 51289 40268
rect 51039 40178 51289 40234
rect 51039 40144 51071 40178
rect 51105 40144 51224 40178
rect 51258 40144 51289 40178
rect 51039 40088 51289 40144
rect 51039 40054 51071 40088
rect 51105 40054 51224 40088
rect 51258 40054 51289 40088
rect 49699 39964 49731 39998
rect 49765 39964 49884 39998
rect 49918 39964 49949 39998
rect 49699 39947 49949 39964
rect 51039 39998 51289 40054
rect 51353 40956 52315 40973
rect 51353 40922 51374 40956
rect 51408 40922 51464 40956
rect 51498 40954 51554 40956
rect 51588 40954 51644 40956
rect 51678 40954 51734 40956
rect 51768 40954 51824 40956
rect 51858 40954 51914 40956
rect 51948 40954 52004 40956
rect 52038 40954 52094 40956
rect 52128 40954 52184 40956
rect 52218 40954 52274 40956
rect 51518 40922 51554 40954
rect 51608 40922 51644 40954
rect 51698 40922 51734 40954
rect 51788 40922 51824 40954
rect 51878 40922 51914 40954
rect 51968 40922 52004 40954
rect 52058 40922 52094 40954
rect 52148 40922 52184 40954
rect 52238 40922 52274 40954
rect 52308 40922 52315 40956
rect 51353 40920 51484 40922
rect 51518 40920 51574 40922
rect 51608 40920 51664 40922
rect 51698 40920 51754 40922
rect 51788 40920 51844 40922
rect 51878 40920 51934 40922
rect 51968 40920 52024 40922
rect 52058 40920 52114 40922
rect 52148 40920 52204 40922
rect 52238 40920 52315 40922
rect 51353 40901 52315 40920
rect 51353 40897 51425 40901
rect 51353 40863 51372 40897
rect 51406 40863 51425 40897
rect 51353 40807 51425 40863
rect 52243 40878 52315 40901
rect 52243 40844 52262 40878
rect 52296 40844 52315 40878
rect 51353 40773 51372 40807
rect 51406 40773 51425 40807
rect 51353 40717 51425 40773
rect 51353 40683 51372 40717
rect 51406 40683 51425 40717
rect 51353 40627 51425 40683
rect 51353 40593 51372 40627
rect 51406 40593 51425 40627
rect 51353 40537 51425 40593
rect 51353 40503 51372 40537
rect 51406 40503 51425 40537
rect 51353 40447 51425 40503
rect 51353 40413 51372 40447
rect 51406 40413 51425 40447
rect 51353 40357 51425 40413
rect 51353 40323 51372 40357
rect 51406 40323 51425 40357
rect 51353 40267 51425 40323
rect 51353 40233 51372 40267
rect 51406 40233 51425 40267
rect 51353 40177 51425 40233
rect 51353 40143 51372 40177
rect 51406 40143 51425 40177
rect 51487 40780 52181 40839
rect 51487 40746 51548 40780
rect 51582 40752 51638 40780
rect 51672 40752 51728 40780
rect 51762 40752 51818 40780
rect 51594 40746 51638 40752
rect 51694 40746 51728 40752
rect 51794 40746 51818 40752
rect 51852 40752 51908 40780
rect 51852 40746 51860 40752
rect 51487 40718 51560 40746
rect 51594 40718 51660 40746
rect 51694 40718 51760 40746
rect 51794 40718 51860 40746
rect 51894 40746 51908 40752
rect 51942 40752 51998 40780
rect 51942 40746 51960 40752
rect 51894 40718 51960 40746
rect 51994 40746 51998 40752
rect 52032 40752 52088 40780
rect 52032 40746 52060 40752
rect 52122 40746 52181 40780
rect 51994 40718 52060 40746
rect 52094 40718 52181 40746
rect 51487 40690 52181 40718
rect 51487 40656 51548 40690
rect 51582 40656 51638 40690
rect 51672 40656 51728 40690
rect 51762 40656 51818 40690
rect 51852 40656 51908 40690
rect 51942 40656 51998 40690
rect 52032 40656 52088 40690
rect 52122 40656 52181 40690
rect 51487 40652 52181 40656
rect 51487 40618 51560 40652
rect 51594 40618 51660 40652
rect 51694 40618 51760 40652
rect 51794 40618 51860 40652
rect 51894 40618 51960 40652
rect 51994 40618 52060 40652
rect 52094 40618 52181 40652
rect 51487 40600 52181 40618
rect 51487 40566 51548 40600
rect 51582 40566 51638 40600
rect 51672 40566 51728 40600
rect 51762 40566 51818 40600
rect 51852 40566 51908 40600
rect 51942 40566 51998 40600
rect 52032 40566 52088 40600
rect 52122 40566 52181 40600
rect 51487 40552 52181 40566
rect 51487 40518 51560 40552
rect 51594 40518 51660 40552
rect 51694 40518 51760 40552
rect 51794 40518 51860 40552
rect 51894 40518 51960 40552
rect 51994 40518 52060 40552
rect 52094 40518 52181 40552
rect 51487 40510 52181 40518
rect 51487 40476 51548 40510
rect 51582 40476 51638 40510
rect 51672 40476 51728 40510
rect 51762 40476 51818 40510
rect 51852 40476 51908 40510
rect 51942 40476 51998 40510
rect 52032 40476 52088 40510
rect 52122 40476 52181 40510
rect 51487 40452 52181 40476
rect 51487 40420 51560 40452
rect 51594 40420 51660 40452
rect 51694 40420 51760 40452
rect 51794 40420 51860 40452
rect 51487 40386 51548 40420
rect 51594 40418 51638 40420
rect 51694 40418 51728 40420
rect 51794 40418 51818 40420
rect 51582 40386 51638 40418
rect 51672 40386 51728 40418
rect 51762 40386 51818 40418
rect 51852 40418 51860 40420
rect 51894 40420 51960 40452
rect 51894 40418 51908 40420
rect 51852 40386 51908 40418
rect 51942 40418 51960 40420
rect 51994 40420 52060 40452
rect 52094 40420 52181 40452
rect 51994 40418 51998 40420
rect 51942 40386 51998 40418
rect 52032 40418 52060 40420
rect 52032 40386 52088 40418
rect 52122 40386 52181 40420
rect 51487 40352 52181 40386
rect 51487 40330 51560 40352
rect 51594 40330 51660 40352
rect 51694 40330 51760 40352
rect 51794 40330 51860 40352
rect 51487 40296 51548 40330
rect 51594 40318 51638 40330
rect 51694 40318 51728 40330
rect 51794 40318 51818 40330
rect 51582 40296 51638 40318
rect 51672 40296 51728 40318
rect 51762 40296 51818 40318
rect 51852 40318 51860 40330
rect 51894 40330 51960 40352
rect 51894 40318 51908 40330
rect 51852 40296 51908 40318
rect 51942 40318 51960 40330
rect 51994 40330 52060 40352
rect 52094 40330 52181 40352
rect 51994 40318 51998 40330
rect 51942 40296 51998 40318
rect 52032 40318 52060 40330
rect 52032 40296 52088 40318
rect 52122 40296 52181 40330
rect 51487 40252 52181 40296
rect 51487 40240 51560 40252
rect 51594 40240 51660 40252
rect 51694 40240 51760 40252
rect 51794 40240 51860 40252
rect 51487 40206 51548 40240
rect 51594 40218 51638 40240
rect 51694 40218 51728 40240
rect 51794 40218 51818 40240
rect 51582 40206 51638 40218
rect 51672 40206 51728 40218
rect 51762 40206 51818 40218
rect 51852 40218 51860 40240
rect 51894 40240 51960 40252
rect 51894 40218 51908 40240
rect 51852 40206 51908 40218
rect 51942 40218 51960 40240
rect 51994 40240 52060 40252
rect 52094 40240 52181 40252
rect 51994 40218 51998 40240
rect 51942 40206 51998 40218
rect 52032 40218 52060 40240
rect 52032 40206 52088 40218
rect 52122 40206 52181 40240
rect 51487 40145 52181 40206
rect 52243 40788 52315 40844
rect 52243 40754 52262 40788
rect 52296 40754 52315 40788
rect 52243 40698 52315 40754
rect 52243 40664 52262 40698
rect 52296 40664 52315 40698
rect 52243 40608 52315 40664
rect 52243 40574 52262 40608
rect 52296 40574 52315 40608
rect 52243 40518 52315 40574
rect 52243 40484 52262 40518
rect 52296 40484 52315 40518
rect 52243 40428 52315 40484
rect 52243 40394 52262 40428
rect 52296 40394 52315 40428
rect 52243 40338 52315 40394
rect 52243 40304 52262 40338
rect 52296 40304 52315 40338
rect 52243 40248 52315 40304
rect 52243 40214 52262 40248
rect 52296 40214 52315 40248
rect 52243 40158 52315 40214
rect 51353 40083 51425 40143
rect 52243 40124 52262 40158
rect 52296 40124 52315 40158
rect 52243 40083 52315 40124
rect 51353 40064 52315 40083
rect 51353 40030 51450 40064
rect 51484 40030 51540 40064
rect 51574 40030 51630 40064
rect 51664 40030 51720 40064
rect 51754 40030 51810 40064
rect 51844 40030 51900 40064
rect 51934 40030 51990 40064
rect 52024 40030 52080 40064
rect 52114 40030 52170 40064
rect 52204 40030 52315 40064
rect 51353 40011 52315 40030
rect 52379 40954 52411 40988
rect 52445 40954 52478 40988
rect 52379 40898 52478 40954
rect 52379 40864 52411 40898
rect 52445 40864 52478 40898
rect 52379 40808 52478 40864
rect 52379 40774 52411 40808
rect 52445 40774 52478 40808
rect 52379 40718 52478 40774
rect 52379 40684 52411 40718
rect 52445 40684 52478 40718
rect 52379 40628 52478 40684
rect 52379 40594 52411 40628
rect 52445 40594 52478 40628
rect 52379 40538 52478 40594
rect 52379 40504 52411 40538
rect 52445 40504 52478 40538
rect 52379 40448 52478 40504
rect 52379 40414 52411 40448
rect 52445 40414 52478 40448
rect 52379 40358 52478 40414
rect 52379 40324 52411 40358
rect 52445 40324 52478 40358
rect 52379 40268 52478 40324
rect 52379 40234 52411 40268
rect 52445 40234 52478 40268
rect 52379 40178 52478 40234
rect 52379 40144 52411 40178
rect 52445 40144 52478 40178
rect 52379 40088 52478 40144
rect 52379 40054 52411 40088
rect 52445 40054 52478 40088
rect 51039 39964 51071 39998
rect 51105 39964 51224 39998
rect 51258 39964 51289 39998
rect 51039 39947 51289 39964
rect 52379 39998 52478 40054
rect 52379 39964 52411 39998
rect 52445 39964 52478 39998
rect 52379 39947 52478 39964
rect 37356 39903 41456 39916
rect 37356 39869 37459 39903
rect 37493 39869 37859 39903
rect 37893 39869 38259 39903
rect 38293 39869 38659 39903
rect 38693 39869 39059 39903
rect 39093 39869 39459 39903
rect 39493 39869 39859 39903
rect 39893 39869 40259 39903
rect 40293 39869 40659 39903
rect 40693 39869 41059 39903
rect 41093 39899 41456 39903
rect 41810 39914 52478 39947
rect 41093 39869 41429 39899
rect 37356 39865 41429 39869
rect 41810 39880 41940 39914
rect 41974 39880 42030 39914
rect 42064 39880 42120 39914
rect 42154 39880 42210 39914
rect 42244 39880 42300 39914
rect 42334 39880 42390 39914
rect 42424 39880 42480 39914
rect 42514 39880 42570 39914
rect 42604 39880 42660 39914
rect 42694 39880 42750 39914
rect 42784 39880 42840 39914
rect 42874 39880 42930 39914
rect 42964 39880 43280 39914
rect 43314 39880 43370 39914
rect 43404 39880 43460 39914
rect 43494 39880 43550 39914
rect 43584 39880 43640 39914
rect 43674 39880 43730 39914
rect 43764 39880 43820 39914
rect 43854 39880 43910 39914
rect 43944 39880 44000 39914
rect 44034 39880 44090 39914
rect 44124 39880 44180 39914
rect 44214 39880 44270 39914
rect 44304 39880 44620 39914
rect 44654 39880 44710 39914
rect 44744 39880 44800 39914
rect 44834 39880 44890 39914
rect 44924 39880 44980 39914
rect 45014 39880 45070 39914
rect 45104 39880 45160 39914
rect 45194 39880 45250 39914
rect 45284 39880 45340 39914
rect 45374 39880 45430 39914
rect 45464 39880 45520 39914
rect 45554 39880 45610 39914
rect 45644 39880 45960 39914
rect 45994 39880 46050 39914
rect 46084 39880 46140 39914
rect 46174 39880 46230 39914
rect 46264 39880 46320 39914
rect 46354 39880 46410 39914
rect 46444 39880 46500 39914
rect 46534 39880 46590 39914
rect 46624 39880 46680 39914
rect 46714 39880 46770 39914
rect 46804 39880 46860 39914
rect 46894 39880 46950 39914
rect 46984 39880 47300 39914
rect 47334 39880 47390 39914
rect 47424 39880 47480 39914
rect 47514 39880 47570 39914
rect 47604 39880 47660 39914
rect 47694 39880 47750 39914
rect 47784 39880 47840 39914
rect 47874 39880 47930 39914
rect 47964 39880 48020 39914
rect 48054 39880 48110 39914
rect 48144 39880 48200 39914
rect 48234 39880 48290 39914
rect 48324 39880 48640 39914
rect 48674 39880 48730 39914
rect 48764 39880 48820 39914
rect 48854 39880 48910 39914
rect 48944 39880 49000 39914
rect 49034 39880 49090 39914
rect 49124 39880 49180 39914
rect 49214 39880 49270 39914
rect 49304 39880 49360 39914
rect 49394 39880 49450 39914
rect 49484 39880 49540 39914
rect 49574 39880 49630 39914
rect 49664 39880 49980 39914
rect 50014 39880 50070 39914
rect 50104 39880 50160 39914
rect 50194 39880 50250 39914
rect 50284 39880 50340 39914
rect 50374 39880 50430 39914
rect 50464 39880 50520 39914
rect 50554 39880 50610 39914
rect 50644 39880 50700 39914
rect 50734 39880 50790 39914
rect 50824 39880 50880 39914
rect 50914 39880 50970 39914
rect 51004 39880 51320 39914
rect 51354 39880 51410 39914
rect 51444 39880 51500 39914
rect 51534 39880 51590 39914
rect 51624 39880 51680 39914
rect 51714 39880 51770 39914
rect 51804 39880 51860 39914
rect 51894 39880 51950 39914
rect 51984 39880 52040 39914
rect 52074 39880 52130 39914
rect 52164 39880 52220 39914
rect 52254 39880 52310 39914
rect 52344 39880 52478 39914
rect 37356 39856 41456 39865
rect 41810 39848 52478 39880
rect 28123 39797 28298 39822
rect 22674 39762 28298 39797
rect 29338 39762 34962 39822
rect 22674 39703 28298 39716
rect 22674 39669 22857 39703
rect 22891 39669 23257 39703
rect 23291 39669 23657 39703
rect 23691 39669 24057 39703
rect 24091 39669 24457 39703
rect 24491 39669 24857 39703
rect 24891 39669 25257 39703
rect 25291 39669 25657 39703
rect 25691 39669 26057 39703
rect 26091 39669 26457 39703
rect 26491 39669 26857 39703
rect 26891 39669 27257 39703
rect 27291 39669 27657 39703
rect 27691 39669 28057 39703
rect 28091 39695 28298 39703
rect 29338 39703 34962 39716
rect 29338 39695 29521 39703
rect 28091 39669 28273 39695
rect 22674 39661 28273 39669
rect 29338 39661 29469 39695
rect 29503 39669 29521 39695
rect 29555 39669 29921 39703
rect 29955 39669 30321 39703
rect 30355 39669 30721 39703
rect 30755 39669 31121 39703
rect 31155 39669 31521 39703
rect 31555 39669 31921 39703
rect 31955 39669 32321 39703
rect 32355 39669 32721 39703
rect 32755 39669 33121 39703
rect 33155 39669 33521 39703
rect 33555 39669 33921 39703
rect 33955 39669 34321 39703
rect 34355 39669 34721 39703
rect 34755 39669 34962 39703
rect 29503 39661 34962 39669
rect 22674 39656 28298 39661
rect 29338 39656 34962 39661
rect 37206 39709 37266 39792
rect 37206 39675 37219 39709
rect 37253 39675 37266 39709
rect 37206 39582 37266 39675
rect 38256 39679 38416 39702
rect 38256 39645 38321 39679
rect 38355 39645 38416 39679
rect 38256 39582 38416 39645
rect 39556 39679 39716 39702
rect 39556 39645 39621 39679
rect 39655 39645 39716 39679
rect 39556 39582 39716 39645
rect 6310 39569 13478 39582
rect 6310 39535 6493 39569
rect 6527 39535 6893 39569
rect 6927 39535 7293 39569
rect 7327 39535 7693 39569
rect 7727 39535 8093 39569
rect 8127 39535 8493 39569
rect 8527 39535 8893 39569
rect 8927 39535 9293 39569
rect 9327 39535 9693 39569
rect 9727 39535 10093 39569
rect 10127 39535 10493 39569
rect 10527 39535 10893 39569
rect 10927 39535 11293 39569
rect 11327 39535 11693 39569
rect 11727 39535 12093 39569
rect 12127 39535 12493 39569
rect 12527 39535 12893 39569
rect 12927 39535 13293 39569
rect 13327 39535 13478 39569
rect 6310 39522 13478 39535
rect 15130 39569 22298 39582
rect 15130 39535 15313 39569
rect 15347 39535 15713 39569
rect 15747 39535 16113 39569
rect 16147 39535 16513 39569
rect 16547 39535 16913 39569
rect 16947 39535 17313 39569
rect 17347 39535 17713 39569
rect 17747 39535 18113 39569
rect 18147 39535 18513 39569
rect 18547 39535 18913 39569
rect 18947 39535 19313 39569
rect 19347 39535 19713 39569
rect 19747 39535 20113 39569
rect 20147 39535 20513 39569
rect 20547 39535 20913 39569
rect 20947 39535 21313 39569
rect 21347 39535 21713 39569
rect 21747 39535 22113 39569
rect 22147 39535 22298 39569
rect 15130 39522 22298 39535
rect 22576 39569 28298 39582
rect 22576 39535 22857 39569
rect 22891 39535 23257 39569
rect 23291 39535 23657 39569
rect 23691 39535 24057 39569
rect 24091 39535 24457 39569
rect 24491 39535 24857 39569
rect 24891 39535 25257 39569
rect 25291 39535 25657 39569
rect 25691 39535 26057 39569
rect 26091 39535 26457 39569
rect 26491 39535 26857 39569
rect 26891 39535 27257 39569
rect 27291 39535 27657 39569
rect 27691 39535 28057 39569
rect 28091 39535 28298 39569
rect 22576 39522 28298 39535
rect 29240 39569 34962 39582
rect 29240 39535 29521 39569
rect 29555 39535 29921 39569
rect 29955 39535 30321 39569
rect 30355 39535 30721 39569
rect 30755 39535 31121 39569
rect 31155 39535 31521 39569
rect 31555 39535 31921 39569
rect 31955 39535 32321 39569
rect 32355 39535 32721 39569
rect 32755 39535 33121 39569
rect 33155 39535 33521 39569
rect 33555 39535 33921 39569
rect 33955 39535 34321 39569
rect 34355 39535 34721 39569
rect 34755 39535 34962 39569
rect 29240 39522 34962 39535
rect 37178 39569 41456 39582
rect 37178 39535 37459 39569
rect 37493 39535 37859 39569
rect 37893 39535 38259 39569
rect 38293 39535 38659 39569
rect 38693 39535 39059 39569
rect 39093 39535 39459 39569
rect 39493 39535 39859 39569
rect 39893 39535 40259 39569
rect 40293 39535 40659 39569
rect 40693 39535 41059 39569
rect 41093 39535 41456 39569
rect 37178 39522 41456 39535
rect 41784 39569 52504 39582
rect 41784 39535 41967 39569
rect 42001 39535 42167 39569
rect 42201 39535 42367 39569
rect 42401 39535 42567 39569
rect 42601 39535 42767 39569
rect 42801 39535 42967 39569
rect 43001 39535 43167 39569
rect 43201 39535 43367 39569
rect 43401 39535 43567 39569
rect 43601 39535 43767 39569
rect 43801 39535 43967 39569
rect 44001 39535 44167 39569
rect 44201 39535 44367 39569
rect 44401 39535 44567 39569
rect 44601 39535 44767 39569
rect 44801 39535 44967 39569
rect 45001 39535 45167 39569
rect 45201 39535 45367 39569
rect 45401 39535 45567 39569
rect 45601 39535 45767 39569
rect 45801 39535 45967 39569
rect 46001 39535 46167 39569
rect 46201 39535 46367 39569
rect 46401 39535 46567 39569
rect 46601 39535 46767 39569
rect 46801 39535 46967 39569
rect 47001 39535 47167 39569
rect 47201 39535 47367 39569
rect 47401 39535 47567 39569
rect 47601 39535 47767 39569
rect 47801 39535 47967 39569
rect 48001 39535 48167 39569
rect 48201 39535 48367 39569
rect 48401 39535 48567 39569
rect 48601 39535 48767 39569
rect 48801 39535 48967 39569
rect 49001 39535 49167 39569
rect 49201 39535 49367 39569
rect 49401 39535 49567 39569
rect 49601 39535 49767 39569
rect 49801 39535 49967 39569
rect 50001 39535 50167 39569
rect 50201 39535 50367 39569
rect 50401 39535 50567 39569
rect 50601 39535 50767 39569
rect 50801 39535 50967 39569
rect 51001 39535 51167 39569
rect 51201 39535 51367 39569
rect 51401 39535 51567 39569
rect 51601 39535 51767 39569
rect 51801 39535 51967 39569
rect 52001 39535 52167 39569
rect 52201 39535 52367 39569
rect 52401 39535 52504 39569
rect 41784 39522 52504 39535
rect 11992 37689 13332 37702
rect 11992 37655 12175 37689
rect 12209 37655 12375 37689
rect 12409 37655 12575 37689
rect 12609 37655 12775 37689
rect 12809 37655 12975 37689
rect 13009 37655 13175 37689
rect 13209 37655 13332 37689
rect 11992 37642 13332 37655
rect 13678 37689 16118 37702
rect 13678 37655 13861 37689
rect 13895 37655 14061 37689
rect 14095 37655 14261 37689
rect 14295 37655 14461 37689
rect 14495 37655 14661 37689
rect 14695 37655 14861 37689
rect 14895 37655 15061 37689
rect 15095 37655 15261 37689
rect 15295 37655 15461 37689
rect 15495 37655 15661 37689
rect 15695 37655 15861 37689
rect 15895 37655 16118 37689
rect 13678 37642 16118 37655
rect 16422 37689 18862 37702
rect 16422 37655 16605 37689
rect 16639 37655 16805 37689
rect 16839 37655 17005 37689
rect 17039 37655 17205 37689
rect 17239 37655 17405 37689
rect 17439 37655 17605 37689
rect 17639 37655 17805 37689
rect 17839 37655 18005 37689
rect 18039 37655 18205 37689
rect 18239 37655 18405 37689
rect 18439 37655 18605 37689
rect 18639 37655 18862 37689
rect 16422 37642 18862 37655
rect 19168 37689 22180 37702
rect 19168 37655 19351 37689
rect 19385 37655 19551 37689
rect 19585 37655 19751 37689
rect 19785 37655 19951 37689
rect 19985 37655 20151 37689
rect 20185 37655 20351 37689
rect 20385 37655 20551 37689
rect 20585 37655 20751 37689
rect 20785 37655 20951 37689
rect 20985 37655 21151 37689
rect 21185 37655 21351 37689
rect 21385 37655 21551 37689
rect 21585 37655 21751 37689
rect 21785 37655 21951 37689
rect 21985 37655 22180 37689
rect 19168 37642 22180 37655
rect 22498 37689 24938 37702
rect 22498 37655 22681 37689
rect 22715 37655 22881 37689
rect 22915 37655 23081 37689
rect 23115 37655 23281 37689
rect 23315 37655 23481 37689
rect 23515 37655 23681 37689
rect 23715 37655 23881 37689
rect 23915 37655 24081 37689
rect 24115 37655 24281 37689
rect 24315 37655 24481 37689
rect 24515 37655 24681 37689
rect 24715 37655 24938 37689
rect 22498 37642 24938 37655
rect 25320 37689 29598 37702
rect 25320 37655 25601 37689
rect 25635 37655 26001 37689
rect 26035 37655 26401 37689
rect 26435 37655 26801 37689
rect 26835 37655 27201 37689
rect 27235 37655 27601 37689
rect 27635 37655 28001 37689
rect 28035 37655 28401 37689
rect 28435 37655 28801 37689
rect 28835 37655 29201 37689
rect 29235 37655 29598 37689
rect 25320 37642 29598 37655
rect 29928 37689 37096 37702
rect 29928 37655 30111 37689
rect 30145 37655 30511 37689
rect 30545 37655 30911 37689
rect 30945 37655 31311 37689
rect 31345 37655 31711 37689
rect 31745 37655 32111 37689
rect 32145 37655 32511 37689
rect 32545 37655 32911 37689
rect 32945 37655 33311 37689
rect 33345 37655 33711 37689
rect 33745 37655 34111 37689
rect 34145 37655 34511 37689
rect 34545 37655 34911 37689
rect 34945 37655 35311 37689
rect 35345 37655 35711 37689
rect 35745 37655 36111 37689
rect 36145 37655 36511 37689
rect 36545 37655 36911 37689
rect 36945 37655 37096 37689
rect 29928 37642 37096 37655
rect 37374 37689 40348 37702
rect 37374 37655 37655 37689
rect 37689 37655 38055 37689
rect 38089 37655 38455 37689
rect 38489 37655 38855 37689
rect 38889 37655 39255 37689
rect 39289 37655 39655 37689
rect 39689 37655 40055 37689
rect 40089 37655 40348 37689
rect 37374 37642 40348 37655
rect 41784 37689 52504 37702
rect 41784 37655 41967 37689
rect 42001 37655 42167 37689
rect 42201 37655 42367 37689
rect 42401 37655 42567 37689
rect 42601 37655 42767 37689
rect 42801 37655 42967 37689
rect 43001 37655 43167 37689
rect 43201 37655 43367 37689
rect 43401 37655 43567 37689
rect 43601 37655 43767 37689
rect 43801 37655 43967 37689
rect 44001 37655 44167 37689
rect 44201 37655 44367 37689
rect 44401 37655 44567 37689
rect 44601 37655 44767 37689
rect 44801 37655 44967 37689
rect 45001 37655 45167 37689
rect 45201 37655 45367 37689
rect 45401 37655 45567 37689
rect 45601 37655 45767 37689
rect 45801 37655 45967 37689
rect 46001 37655 46167 37689
rect 46201 37655 46367 37689
rect 46401 37655 46567 37689
rect 46601 37655 46767 37689
rect 46801 37655 46967 37689
rect 47001 37655 47167 37689
rect 47201 37655 47367 37689
rect 47401 37655 47567 37689
rect 47601 37655 47767 37689
rect 47801 37655 47967 37689
rect 48001 37655 48167 37689
rect 48201 37655 48367 37689
rect 48401 37655 48567 37689
rect 48601 37655 48767 37689
rect 48801 37655 48967 37689
rect 49001 37655 49167 37689
rect 49201 37655 49367 37689
rect 49401 37655 49567 37689
rect 49601 37655 49767 37689
rect 49801 37655 49967 37689
rect 50001 37655 50167 37689
rect 50201 37655 50367 37689
rect 50401 37655 50567 37689
rect 50601 37655 50767 37689
rect 50801 37655 50967 37689
rect 51001 37655 51167 37689
rect 51201 37655 51367 37689
rect 51401 37655 51567 37689
rect 51601 37655 51767 37689
rect 51801 37655 51967 37689
rect 52001 37655 52167 37689
rect 52201 37655 52367 37689
rect 52401 37655 52504 37689
rect 41784 37642 52504 37655
rect 37402 37549 37462 37642
rect 38450 37599 38610 37642
rect 38450 37565 38515 37599
rect 38549 37565 38610 37599
rect 38450 37562 38610 37565
rect 25418 37482 29598 37542
rect 37402 37515 37415 37549
rect 37449 37515 37462 37549
rect 12018 37341 13306 37376
rect 12018 37318 12148 37341
rect 12018 37284 12052 37318
rect 12086 37307 12148 37318
rect 12182 37307 12238 37341
rect 12272 37307 12328 37341
rect 12362 37307 12418 37341
rect 12452 37307 12508 37341
rect 12542 37307 12598 37341
rect 12632 37307 12688 37341
rect 12722 37307 12778 37341
rect 12812 37307 12868 37341
rect 12902 37307 12958 37341
rect 12992 37307 13048 37341
rect 13082 37307 13138 37341
rect 13172 37318 13306 37341
rect 13172 37307 13239 37318
rect 12086 37284 13239 37307
rect 13273 37284 13306 37318
rect 12018 37277 13306 37284
rect 12018 37228 12117 37277
rect 12018 37194 12052 37228
rect 12086 37194 12117 37228
rect 13207 37228 13306 37277
rect 12018 37138 12117 37194
rect 12018 37104 12052 37138
rect 12086 37104 12117 37138
rect 12018 37048 12117 37104
rect 12018 37014 12052 37048
rect 12086 37014 12117 37048
rect 12018 36958 12117 37014
rect 12018 36924 12052 36958
rect 12086 36924 12117 36958
rect 12018 36868 12117 36924
rect 12018 36834 12052 36868
rect 12086 36834 12117 36868
rect 12018 36778 12117 36834
rect 12018 36744 12052 36778
rect 12086 36744 12117 36778
rect 12018 36688 12117 36744
rect 12018 36654 12052 36688
rect 12086 36654 12117 36688
rect 12018 36598 12117 36654
rect 12018 36564 12052 36598
rect 12086 36564 12117 36598
rect 12018 36508 12117 36564
rect 12018 36474 12052 36508
rect 12086 36474 12117 36508
rect 12018 36418 12117 36474
rect 12018 36384 12052 36418
rect 12086 36384 12117 36418
rect 12018 36328 12117 36384
rect 12018 36294 12052 36328
rect 12086 36294 12117 36328
rect 12018 36238 12117 36294
rect 12181 37194 13143 37213
rect 12181 37160 12312 37194
rect 12346 37160 12402 37194
rect 12436 37160 12492 37194
rect 12526 37160 12582 37194
rect 12616 37160 12672 37194
rect 12706 37160 12762 37194
rect 12796 37160 12852 37194
rect 12886 37160 12942 37194
rect 12976 37160 13032 37194
rect 13066 37160 13143 37194
rect 12181 37141 13143 37160
rect 12181 37137 12253 37141
rect 12181 37103 12200 37137
rect 12234 37103 12253 37137
rect 12181 37047 12253 37103
rect 13071 37118 13143 37141
rect 13071 37084 13090 37118
rect 13124 37084 13143 37118
rect 12181 37013 12200 37047
rect 12234 37013 12253 37047
rect 12181 36957 12253 37013
rect 12181 36923 12200 36957
rect 12234 36923 12253 36957
rect 12181 36867 12253 36923
rect 12181 36833 12200 36867
rect 12234 36833 12253 36867
rect 12181 36777 12253 36833
rect 12181 36743 12200 36777
rect 12234 36743 12253 36777
rect 12181 36687 12253 36743
rect 12181 36653 12200 36687
rect 12234 36653 12253 36687
rect 12181 36597 12253 36653
rect 12181 36563 12200 36597
rect 12234 36563 12253 36597
rect 12181 36507 12253 36563
rect 12181 36473 12200 36507
rect 12234 36473 12253 36507
rect 12181 36417 12253 36473
rect 12181 36383 12200 36417
rect 12234 36383 12253 36417
rect 12315 37020 13009 37079
rect 12315 36986 12376 37020
rect 12410 36992 12466 37020
rect 12500 36992 12556 37020
rect 12590 36992 12646 37020
rect 12422 36986 12466 36992
rect 12522 36986 12556 36992
rect 12622 36986 12646 36992
rect 12680 36992 12736 37020
rect 12680 36986 12688 36992
rect 12315 36958 12388 36986
rect 12422 36958 12488 36986
rect 12522 36958 12588 36986
rect 12622 36958 12688 36986
rect 12722 36986 12736 36992
rect 12770 36992 12826 37020
rect 12770 36986 12788 36992
rect 12722 36958 12788 36986
rect 12822 36986 12826 36992
rect 12860 36992 12916 37020
rect 12860 36986 12888 36992
rect 12950 36986 13009 37020
rect 12822 36958 12888 36986
rect 12922 36958 13009 36986
rect 12315 36930 13009 36958
rect 12315 36896 12376 36930
rect 12410 36896 12466 36930
rect 12500 36896 12556 36930
rect 12590 36896 12646 36930
rect 12680 36896 12736 36930
rect 12770 36896 12826 36930
rect 12860 36896 12916 36930
rect 12950 36896 13009 36930
rect 12315 36892 13009 36896
rect 12315 36858 12388 36892
rect 12422 36858 12488 36892
rect 12522 36858 12588 36892
rect 12622 36858 12688 36892
rect 12722 36858 12788 36892
rect 12822 36858 12888 36892
rect 12922 36858 13009 36892
rect 12315 36840 13009 36858
rect 12315 36806 12376 36840
rect 12410 36806 12466 36840
rect 12500 36806 12556 36840
rect 12590 36806 12646 36840
rect 12680 36806 12736 36840
rect 12770 36806 12826 36840
rect 12860 36806 12916 36840
rect 12950 36806 13009 36840
rect 12315 36792 13009 36806
rect 12315 36758 12388 36792
rect 12422 36758 12488 36792
rect 12522 36758 12588 36792
rect 12622 36758 12688 36792
rect 12722 36758 12788 36792
rect 12822 36758 12888 36792
rect 12922 36758 13009 36792
rect 12315 36750 13009 36758
rect 12315 36716 12376 36750
rect 12410 36716 12466 36750
rect 12500 36716 12556 36750
rect 12590 36716 12646 36750
rect 12680 36716 12736 36750
rect 12770 36716 12826 36750
rect 12860 36716 12916 36750
rect 12950 36716 13009 36750
rect 12315 36692 13009 36716
rect 12315 36660 12388 36692
rect 12422 36660 12488 36692
rect 12522 36660 12588 36692
rect 12622 36660 12688 36692
rect 12315 36626 12376 36660
rect 12422 36658 12466 36660
rect 12522 36658 12556 36660
rect 12622 36658 12646 36660
rect 12410 36626 12466 36658
rect 12500 36626 12556 36658
rect 12590 36626 12646 36658
rect 12680 36658 12688 36660
rect 12722 36660 12788 36692
rect 12722 36658 12736 36660
rect 12680 36626 12736 36658
rect 12770 36658 12788 36660
rect 12822 36660 12888 36692
rect 12922 36660 13009 36692
rect 12822 36658 12826 36660
rect 12770 36626 12826 36658
rect 12860 36658 12888 36660
rect 12860 36626 12916 36658
rect 12950 36626 13009 36660
rect 12315 36592 13009 36626
rect 12315 36570 12388 36592
rect 12422 36570 12488 36592
rect 12522 36570 12588 36592
rect 12622 36570 12688 36592
rect 12315 36536 12376 36570
rect 12422 36558 12466 36570
rect 12522 36558 12556 36570
rect 12622 36558 12646 36570
rect 12410 36536 12466 36558
rect 12500 36536 12556 36558
rect 12590 36536 12646 36558
rect 12680 36558 12688 36570
rect 12722 36570 12788 36592
rect 12722 36558 12736 36570
rect 12680 36536 12736 36558
rect 12770 36558 12788 36570
rect 12822 36570 12888 36592
rect 12922 36570 13009 36592
rect 12822 36558 12826 36570
rect 12770 36536 12826 36558
rect 12860 36558 12888 36570
rect 12860 36536 12916 36558
rect 12950 36536 13009 36570
rect 12315 36492 13009 36536
rect 12315 36480 12388 36492
rect 12422 36480 12488 36492
rect 12522 36480 12588 36492
rect 12622 36480 12688 36492
rect 12315 36446 12376 36480
rect 12422 36458 12466 36480
rect 12522 36458 12556 36480
rect 12622 36458 12646 36480
rect 12410 36446 12466 36458
rect 12500 36446 12556 36458
rect 12590 36446 12646 36458
rect 12680 36458 12688 36480
rect 12722 36480 12788 36492
rect 12722 36458 12736 36480
rect 12680 36446 12736 36458
rect 12770 36458 12788 36480
rect 12822 36480 12888 36492
rect 12922 36480 13009 36492
rect 12822 36458 12826 36480
rect 12770 36446 12826 36458
rect 12860 36458 12888 36480
rect 12860 36446 12916 36458
rect 12950 36446 13009 36480
rect 12315 36385 13009 36446
rect 13071 37028 13143 37084
rect 13071 36994 13090 37028
rect 13124 36994 13143 37028
rect 13071 36938 13143 36994
rect 13071 36904 13090 36938
rect 13124 36904 13143 36938
rect 13071 36848 13143 36904
rect 13071 36814 13090 36848
rect 13124 36814 13143 36848
rect 13071 36758 13143 36814
rect 13071 36724 13090 36758
rect 13124 36724 13143 36758
rect 13071 36668 13143 36724
rect 13071 36634 13090 36668
rect 13124 36634 13143 36668
rect 13071 36578 13143 36634
rect 13071 36544 13090 36578
rect 13124 36544 13143 36578
rect 13071 36488 13143 36544
rect 13071 36454 13090 36488
rect 13124 36454 13143 36488
rect 13071 36398 13143 36454
rect 12181 36323 12253 36383
rect 13071 36364 13090 36398
rect 13124 36364 13143 36398
rect 13071 36323 13143 36364
rect 12181 36304 13143 36323
rect 12181 36270 12278 36304
rect 12312 36270 12368 36304
rect 12402 36270 12458 36304
rect 12492 36270 12548 36304
rect 12582 36270 12638 36304
rect 12672 36270 12728 36304
rect 12762 36270 12818 36304
rect 12852 36270 12908 36304
rect 12942 36270 12998 36304
rect 13032 36295 13143 36304
rect 13032 36270 13093 36295
rect 12181 36261 13093 36270
rect 13127 36261 13143 36295
rect 12181 36251 13143 36261
rect 13207 37194 13239 37228
rect 13273 37194 13306 37228
rect 13207 37138 13306 37194
rect 13207 37104 13239 37138
rect 13273 37104 13306 37138
rect 13207 37048 13306 37104
rect 13207 37014 13239 37048
rect 13273 37014 13306 37048
rect 13207 36958 13306 37014
rect 13207 36924 13239 36958
rect 13273 36924 13306 36958
rect 13207 36868 13306 36924
rect 13207 36834 13239 36868
rect 13273 36834 13306 36868
rect 25887 37196 25921 37482
rect 26803 37196 26837 37482
rect 27719 37196 27753 37482
rect 28635 37196 28669 37482
rect 29551 37196 29585 37482
rect 37402 37432 37462 37515
rect 37532 37519 40348 37522
rect 37532 37485 37565 37519
rect 37599 37485 40348 37519
rect 37532 37482 40348 37485
rect 37519 37421 37553 37441
rect 37519 37353 37553 37387
rect 37519 37285 37553 37315
rect 37519 37217 37553 37243
rect 13207 36778 13306 36834
rect 13207 36744 13239 36778
rect 13273 36744 13306 36778
rect 13207 36688 13306 36744
rect 13207 36654 13239 36688
rect 13273 36654 13306 36688
rect 13207 36598 13306 36654
rect 13207 36564 13239 36598
rect 13273 36564 13306 36598
rect 13207 36508 13306 36564
rect 13207 36474 13239 36508
rect 13273 36474 13306 36508
rect 14590 36723 15206 36762
rect 14590 36621 14677 36723
rect 15119 36621 15206 36723
rect 13207 36418 13306 36474
rect 13207 36384 13239 36418
rect 13273 36384 13306 36418
rect 13207 36328 13306 36384
rect 13207 36294 13239 36328
rect 13273 36294 13306 36328
rect 12018 36204 12052 36238
rect 12086 36204 12117 36238
rect 12018 36187 12117 36204
rect 13207 36238 13306 36294
rect 13207 36204 13239 36238
rect 13273 36204 13306 36238
rect 13207 36187 13306 36204
rect 12018 36159 13306 36187
rect 12018 36154 13277 36159
rect 12018 36120 12148 36154
rect 12182 36120 12238 36154
rect 12272 36120 12328 36154
rect 12362 36120 12418 36154
rect 12452 36120 12508 36154
rect 12542 36120 12598 36154
rect 12632 36120 12688 36154
rect 12722 36120 12778 36154
rect 12812 36120 12868 36154
rect 12902 36120 12958 36154
rect 12992 36120 13048 36154
rect 13082 36120 13138 36154
rect 13172 36125 13277 36154
rect 13172 36120 13306 36125
rect 12018 36088 13306 36120
rect 14590 35822 15206 36621
rect 15686 36477 16118 36867
rect 17334 36723 17950 36762
rect 17334 36621 17421 36723
rect 17863 36621 17950 36723
rect 17334 35822 17950 36621
rect 18430 36477 18862 36867
rect 20366 36723 20982 36762
rect 20366 36621 20453 36723
rect 20895 36621 20982 36723
rect 20366 35822 20982 36621
rect 21749 36477 22181 36867
rect 23410 36723 24026 36762
rect 23410 36621 23497 36723
rect 23939 36621 24026 36723
rect 23410 35822 24026 36621
rect 24506 36477 24938 36867
rect 25430 37169 25464 37196
rect 25887 37178 25922 37196
rect 25430 37097 25464 37115
rect 25430 37025 25464 37047
rect 25430 36953 25464 36979
rect 25430 36881 25464 36911
rect 25430 36809 25464 36843
rect 25430 36741 25464 36775
rect 25430 36673 25464 36703
rect 25430 36605 25464 36631
rect 25430 36537 25464 36559
rect 25430 36469 25464 36487
rect 25429 36415 25430 36446
rect 25429 36388 25464 36415
rect 25888 37169 25922 37178
rect 25888 37097 25922 37115
rect 25888 37025 25922 37047
rect 25888 36953 25922 36979
rect 25888 36881 25922 36911
rect 25888 36809 25922 36843
rect 25888 36741 25922 36775
rect 25888 36673 25922 36703
rect 25888 36605 25922 36631
rect 25888 36537 25922 36559
rect 25888 36469 25922 36487
rect 26346 37169 26380 37196
rect 26803 37178 26838 37196
rect 26346 37097 26380 37115
rect 26346 37025 26380 37047
rect 26346 36953 26380 36979
rect 26346 36881 26380 36911
rect 26346 36809 26380 36843
rect 26346 36741 26380 36775
rect 26346 36673 26380 36703
rect 26346 36605 26380 36631
rect 26346 36537 26380 36559
rect 26346 36469 26380 36487
rect 25888 36388 25922 36415
rect 26345 36415 26346 36446
rect 26345 36388 26380 36415
rect 26804 37169 26838 37178
rect 26804 37097 26838 37115
rect 26804 37025 26838 37047
rect 26804 36953 26838 36979
rect 26804 36881 26838 36911
rect 26804 36809 26838 36843
rect 26804 36741 26838 36775
rect 26804 36673 26838 36703
rect 26804 36605 26838 36631
rect 26804 36537 26838 36559
rect 26804 36469 26838 36487
rect 27262 37169 27296 37196
rect 27719 37178 27754 37196
rect 27262 37097 27296 37115
rect 27262 37025 27296 37047
rect 27262 36953 27296 36979
rect 27262 36881 27296 36911
rect 27262 36809 27296 36843
rect 27262 36741 27296 36775
rect 27262 36673 27296 36703
rect 27262 36605 27296 36631
rect 27262 36537 27296 36559
rect 27262 36469 27296 36487
rect 26804 36388 26838 36415
rect 27261 36415 27262 36446
rect 27261 36388 27296 36415
rect 27720 37169 27754 37178
rect 27720 37097 27754 37115
rect 27720 37025 27754 37047
rect 27720 36953 27754 36979
rect 27720 36881 27754 36911
rect 27720 36809 27754 36843
rect 27720 36741 27754 36775
rect 27720 36673 27754 36703
rect 27720 36605 27754 36631
rect 27720 36537 27754 36559
rect 27720 36469 27754 36487
rect 28178 37169 28212 37196
rect 28635 37178 28670 37196
rect 28178 37097 28212 37115
rect 28178 37025 28212 37047
rect 28178 36953 28212 36979
rect 28178 36881 28212 36911
rect 28178 36809 28212 36843
rect 28178 36741 28212 36775
rect 28178 36673 28212 36703
rect 28178 36605 28212 36631
rect 28178 36537 28212 36559
rect 28178 36469 28212 36487
rect 27720 36388 27754 36415
rect 28177 36415 28178 36446
rect 28177 36388 28212 36415
rect 28636 37169 28670 37178
rect 28636 37097 28670 37115
rect 28636 37025 28670 37047
rect 28636 36953 28670 36979
rect 28636 36881 28670 36911
rect 28636 36809 28670 36843
rect 28636 36741 28670 36775
rect 28636 36673 28670 36703
rect 28636 36605 28670 36631
rect 28636 36537 28670 36559
rect 28636 36469 28670 36487
rect 29094 37169 29128 37196
rect 29551 37178 29586 37196
rect 29094 37097 29128 37115
rect 29094 37025 29128 37047
rect 29094 36953 29128 36979
rect 29094 36881 29128 36911
rect 29094 36809 29128 36843
rect 29094 36741 29128 36775
rect 29094 36673 29128 36703
rect 29094 36605 29128 36631
rect 29094 36537 29128 36559
rect 29094 36469 29128 36487
rect 28636 36388 28670 36415
rect 29093 36415 29094 36446
rect 29093 36388 29128 36415
rect 29552 37169 29586 37178
rect 29552 37097 29586 37115
rect 29552 37025 29586 37047
rect 29552 36953 29586 36979
rect 29552 36881 29586 36911
rect 29552 36809 29586 36843
rect 29552 36741 29586 36775
rect 29552 36673 29586 36703
rect 29552 36605 29586 36631
rect 29552 36537 29586 36559
rect 29552 36469 29586 36487
rect 29552 36388 29586 36415
rect 37519 37149 37553 37171
rect 37519 37081 37553 37099
rect 37519 37013 37553 37027
rect 37519 36945 37553 36955
rect 37519 36877 37553 36883
rect 37519 36809 37553 36811
rect 37519 36773 37553 36775
rect 37519 36701 37553 36707
rect 37519 36629 37553 36639
rect 37519 36557 37553 36571
rect 37519 36485 37553 36503
rect 37519 36413 37553 36435
rect 25429 36322 25463 36388
rect 26345 36322 26379 36388
rect 27261 36322 27295 36388
rect 28177 36322 28211 36388
rect 29093 36322 29127 36388
rect 37519 36341 37553 36367
rect 25418 36262 29598 36322
rect 37519 36269 37553 36299
rect 37519 36197 37553 36231
rect 25498 36143 28089 36156
rect 25498 36109 25601 36143
rect 25635 36109 26001 36143
rect 26035 36109 26401 36143
rect 26435 36109 26801 36143
rect 26835 36109 27201 36143
rect 27235 36109 27601 36143
rect 27635 36109 28001 36143
rect 28035 36125 28089 36143
rect 28123 36143 29598 36156
rect 28123 36125 28401 36143
rect 28035 36109 28401 36125
rect 28435 36109 28801 36143
rect 28835 36109 29201 36143
rect 29235 36109 29598 36143
rect 25498 36096 29598 36109
rect 37519 36062 37553 36163
rect 37977 37421 38011 37482
rect 37977 37353 38011 37387
rect 37977 37285 38011 37315
rect 37977 37217 38011 37243
rect 37977 37149 38011 37171
rect 37977 37081 38011 37099
rect 37977 37013 38011 37027
rect 37977 36945 38011 36955
rect 37977 36877 38011 36883
rect 37977 36809 38011 36811
rect 37977 36773 38011 36775
rect 37977 36701 38011 36707
rect 37977 36629 38011 36639
rect 37977 36557 38011 36571
rect 37977 36485 38011 36503
rect 37977 36413 38011 36435
rect 37977 36341 38011 36367
rect 37977 36269 38011 36299
rect 37977 36197 38011 36231
rect 37977 36143 38011 36163
rect 38435 37421 38469 37441
rect 38435 37353 38469 37387
rect 38435 37285 38469 37315
rect 38435 37217 38469 37243
rect 38435 37149 38469 37171
rect 38435 37081 38469 37099
rect 38435 37013 38469 37027
rect 38435 36945 38469 36955
rect 38435 36877 38469 36883
rect 38435 36809 38469 36811
rect 38435 36773 38469 36775
rect 38435 36701 38469 36707
rect 38435 36629 38469 36639
rect 38435 36557 38469 36571
rect 38435 36485 38469 36503
rect 38435 36413 38469 36435
rect 38435 36341 38469 36367
rect 38435 36269 38469 36299
rect 38435 36197 38469 36231
rect 38435 36062 38469 36163
rect 38893 37421 38927 37482
rect 38893 37353 38927 37387
rect 38893 37285 38927 37315
rect 38893 37217 38927 37243
rect 38893 37149 38927 37171
rect 38893 37081 38927 37099
rect 38893 37013 38927 37027
rect 38893 36945 38927 36955
rect 38893 36877 38927 36883
rect 38893 36809 38927 36811
rect 38893 36773 38927 36775
rect 38893 36701 38927 36707
rect 38893 36629 38927 36639
rect 38893 36557 38927 36571
rect 38893 36485 38927 36503
rect 38893 36413 38927 36435
rect 38893 36341 38927 36367
rect 38893 36269 38927 36299
rect 38893 36197 38927 36231
rect 38893 36143 38927 36163
rect 39351 37421 39385 37441
rect 39351 37353 39385 37387
rect 39351 37285 39385 37315
rect 39351 37217 39385 37243
rect 39351 37149 39385 37171
rect 39351 37081 39385 37099
rect 39351 37013 39385 37027
rect 39351 36945 39385 36955
rect 39351 36877 39385 36883
rect 39351 36809 39385 36811
rect 39351 36773 39385 36775
rect 39351 36701 39385 36707
rect 39351 36629 39385 36639
rect 39351 36557 39385 36571
rect 39351 36485 39385 36503
rect 39351 36413 39385 36435
rect 39351 36341 39385 36367
rect 39351 36269 39385 36299
rect 39351 36197 39385 36231
rect 39351 36062 39385 36163
rect 39809 37421 39843 37482
rect 39809 37353 39843 37387
rect 39809 37285 39843 37315
rect 39809 37217 39843 37243
rect 39809 37149 39843 37171
rect 39809 37081 39843 37099
rect 39809 37013 39843 37027
rect 39809 36945 39843 36955
rect 39809 36877 39843 36883
rect 39809 36809 39843 36811
rect 39809 36773 39843 36775
rect 39809 36701 39843 36707
rect 39809 36629 39843 36639
rect 39809 36557 39843 36571
rect 39809 36485 39843 36503
rect 39809 36413 39843 36435
rect 39809 36341 39843 36367
rect 39809 36269 39843 36299
rect 39809 36197 39843 36231
rect 39809 36143 39843 36163
rect 40267 37421 40301 37441
rect 40267 37353 40301 37387
rect 40267 37285 40301 37315
rect 40267 37217 40301 37243
rect 40267 37149 40301 37171
rect 40267 37081 40301 37099
rect 40267 37013 40301 37027
rect 40267 36945 40301 36955
rect 40267 36877 40301 36883
rect 40267 36809 40301 36811
rect 40267 36773 40301 36775
rect 40267 36701 40301 36707
rect 40267 36629 40301 36639
rect 40267 36557 40301 36571
rect 40267 36485 40301 36503
rect 40267 36413 40301 36435
rect 40267 36341 40301 36367
rect 40267 36269 40301 36299
rect 40267 36197 40301 36231
rect 40267 36062 40301 36163
rect 41810 37356 52478 37376
rect 41810 37322 41830 37356
rect 41864 37322 41920 37356
rect 41954 37341 42010 37356
rect 42044 37341 42100 37356
rect 42134 37341 42190 37356
rect 42224 37341 42280 37356
rect 42314 37341 42370 37356
rect 42404 37341 42460 37356
rect 42494 37341 42550 37356
rect 42584 37341 42640 37356
rect 42674 37341 42730 37356
rect 42764 37341 42820 37356
rect 42854 37341 42910 37356
rect 42944 37341 43000 37356
rect 41974 37322 42010 37341
rect 42064 37322 42100 37341
rect 42154 37322 42190 37341
rect 42244 37322 42280 37341
rect 42334 37322 42370 37341
rect 42424 37322 42460 37341
rect 42514 37322 42550 37341
rect 42604 37322 42640 37341
rect 42694 37322 42730 37341
rect 42784 37322 42820 37341
rect 42874 37322 42910 37341
rect 42964 37322 43000 37341
rect 43034 37322 43170 37356
rect 43204 37322 43260 37356
rect 43294 37341 43350 37356
rect 43384 37341 43440 37356
rect 43474 37341 43530 37356
rect 43564 37341 43620 37356
rect 43654 37341 43710 37356
rect 43744 37341 43800 37356
rect 43834 37341 43890 37356
rect 43924 37341 43980 37356
rect 44014 37341 44070 37356
rect 44104 37341 44160 37356
rect 44194 37341 44250 37356
rect 44284 37341 44340 37356
rect 43314 37322 43350 37341
rect 43404 37322 43440 37341
rect 43494 37322 43530 37341
rect 43584 37322 43620 37341
rect 43674 37322 43710 37341
rect 43764 37322 43800 37341
rect 43854 37322 43890 37341
rect 43944 37322 43980 37341
rect 44034 37322 44070 37341
rect 44124 37322 44160 37341
rect 44214 37322 44250 37341
rect 44304 37322 44340 37341
rect 44374 37322 44510 37356
rect 44544 37322 44600 37356
rect 44634 37341 44690 37356
rect 44724 37341 44780 37356
rect 44814 37341 44870 37356
rect 44904 37341 44960 37356
rect 44994 37341 45050 37356
rect 45084 37341 45140 37356
rect 45174 37341 45230 37356
rect 45264 37341 45320 37356
rect 45354 37341 45410 37356
rect 45444 37341 45500 37356
rect 45534 37341 45590 37356
rect 45624 37341 45680 37356
rect 44654 37322 44690 37341
rect 44744 37322 44780 37341
rect 44834 37322 44870 37341
rect 44924 37322 44960 37341
rect 45014 37322 45050 37341
rect 45104 37322 45140 37341
rect 45194 37322 45230 37341
rect 45284 37322 45320 37341
rect 45374 37322 45410 37341
rect 45464 37322 45500 37341
rect 45554 37322 45590 37341
rect 45644 37322 45680 37341
rect 45714 37322 45850 37356
rect 45884 37322 45940 37356
rect 45974 37341 46030 37356
rect 46064 37341 46120 37356
rect 46154 37341 46210 37356
rect 46244 37341 46300 37356
rect 46334 37341 46390 37356
rect 46424 37341 46480 37356
rect 46514 37341 46570 37356
rect 46604 37341 46660 37356
rect 46694 37341 46750 37356
rect 46784 37341 46840 37356
rect 46874 37341 46930 37356
rect 46964 37341 47020 37356
rect 45994 37322 46030 37341
rect 46084 37322 46120 37341
rect 46174 37322 46210 37341
rect 46264 37322 46300 37341
rect 46354 37322 46390 37341
rect 46444 37322 46480 37341
rect 46534 37322 46570 37341
rect 46624 37322 46660 37341
rect 46714 37322 46750 37341
rect 46804 37322 46840 37341
rect 46894 37322 46930 37341
rect 46984 37322 47020 37341
rect 47054 37322 47190 37356
rect 47224 37322 47280 37356
rect 47314 37341 47370 37356
rect 47404 37341 47460 37356
rect 47494 37341 47550 37356
rect 47584 37341 47640 37356
rect 47674 37341 47730 37356
rect 47764 37341 47820 37356
rect 47854 37341 47910 37356
rect 47944 37341 48000 37356
rect 48034 37341 48090 37356
rect 48124 37341 48180 37356
rect 48214 37341 48270 37356
rect 48304 37341 48360 37356
rect 47334 37322 47370 37341
rect 47424 37322 47460 37341
rect 47514 37322 47550 37341
rect 47604 37322 47640 37341
rect 47694 37322 47730 37341
rect 47784 37322 47820 37341
rect 47874 37322 47910 37341
rect 47964 37322 48000 37341
rect 48054 37322 48090 37341
rect 48144 37322 48180 37341
rect 48234 37322 48270 37341
rect 48324 37322 48360 37341
rect 48394 37322 48530 37356
rect 48564 37322 48620 37356
rect 48654 37341 48710 37356
rect 48744 37341 48800 37356
rect 48834 37341 48890 37356
rect 48924 37341 48980 37356
rect 49014 37341 49070 37356
rect 49104 37341 49160 37356
rect 49194 37341 49250 37356
rect 49284 37341 49340 37356
rect 49374 37341 49430 37356
rect 49464 37341 49520 37356
rect 49554 37341 49610 37356
rect 49644 37341 49700 37356
rect 48674 37322 48710 37341
rect 48764 37322 48800 37341
rect 48854 37322 48890 37341
rect 48944 37322 48980 37341
rect 49034 37322 49070 37341
rect 49124 37322 49160 37341
rect 49214 37322 49250 37341
rect 49304 37322 49340 37341
rect 49394 37322 49430 37341
rect 49484 37322 49520 37341
rect 49574 37322 49610 37341
rect 49664 37322 49700 37341
rect 49734 37322 49870 37356
rect 49904 37322 49960 37356
rect 49994 37341 50050 37356
rect 50084 37341 50140 37356
rect 50174 37341 50230 37356
rect 50264 37341 50320 37356
rect 50354 37341 50410 37356
rect 50444 37341 50500 37356
rect 50534 37341 50590 37356
rect 50624 37341 50680 37356
rect 50714 37341 50770 37356
rect 50804 37341 50860 37356
rect 50894 37341 50950 37356
rect 50984 37341 51040 37356
rect 50014 37322 50050 37341
rect 50104 37322 50140 37341
rect 50194 37322 50230 37341
rect 50284 37322 50320 37341
rect 50374 37322 50410 37341
rect 50464 37322 50500 37341
rect 50554 37322 50590 37341
rect 50644 37322 50680 37341
rect 50734 37322 50770 37341
rect 50824 37322 50860 37341
rect 50914 37322 50950 37341
rect 51004 37322 51040 37341
rect 51074 37322 51210 37356
rect 51244 37322 51300 37356
rect 51334 37341 51390 37356
rect 51424 37341 51480 37356
rect 51514 37341 51570 37356
rect 51604 37341 51660 37356
rect 51694 37341 51750 37356
rect 51784 37341 51840 37356
rect 51874 37341 51930 37356
rect 51964 37341 52020 37356
rect 52054 37341 52110 37356
rect 52144 37341 52200 37356
rect 52234 37341 52290 37356
rect 52324 37341 52380 37356
rect 51354 37322 51390 37341
rect 51444 37322 51480 37341
rect 51534 37322 51570 37341
rect 51624 37322 51660 37341
rect 51714 37322 51750 37341
rect 51804 37322 51840 37341
rect 51894 37322 51930 37341
rect 51984 37322 52020 37341
rect 52074 37322 52110 37341
rect 52164 37322 52200 37341
rect 52254 37322 52290 37341
rect 52344 37322 52380 37341
rect 52414 37322 52478 37356
rect 41810 37318 41940 37322
rect 41810 37284 41844 37318
rect 41878 37307 41940 37318
rect 41974 37307 42030 37322
rect 42064 37307 42120 37322
rect 42154 37307 42210 37322
rect 42244 37307 42300 37322
rect 42334 37307 42390 37322
rect 42424 37307 42480 37322
rect 42514 37307 42570 37322
rect 42604 37307 42660 37322
rect 42694 37307 42750 37322
rect 42784 37307 42840 37322
rect 42874 37307 42930 37322
rect 42964 37318 43280 37322
rect 42964 37307 43031 37318
rect 41878 37284 43031 37307
rect 43065 37284 43184 37318
rect 43218 37307 43280 37318
rect 43314 37307 43370 37322
rect 43404 37307 43460 37322
rect 43494 37307 43550 37322
rect 43584 37307 43640 37322
rect 43674 37307 43730 37322
rect 43764 37307 43820 37322
rect 43854 37307 43910 37322
rect 43944 37307 44000 37322
rect 44034 37307 44090 37322
rect 44124 37307 44180 37322
rect 44214 37307 44270 37322
rect 44304 37318 44620 37322
rect 44304 37307 44371 37318
rect 43218 37284 44371 37307
rect 44405 37284 44524 37318
rect 44558 37307 44620 37318
rect 44654 37307 44710 37322
rect 44744 37307 44800 37322
rect 44834 37307 44890 37322
rect 44924 37307 44980 37322
rect 45014 37307 45070 37322
rect 45104 37307 45160 37322
rect 45194 37307 45250 37322
rect 45284 37307 45340 37322
rect 45374 37307 45430 37322
rect 45464 37307 45520 37322
rect 45554 37307 45610 37322
rect 45644 37318 45960 37322
rect 45644 37307 45711 37318
rect 44558 37284 45711 37307
rect 45745 37284 45864 37318
rect 45898 37307 45960 37318
rect 45994 37307 46050 37322
rect 46084 37307 46140 37322
rect 46174 37307 46230 37322
rect 46264 37307 46320 37322
rect 46354 37307 46410 37322
rect 46444 37307 46500 37322
rect 46534 37307 46590 37322
rect 46624 37307 46680 37322
rect 46714 37307 46770 37322
rect 46804 37307 46860 37322
rect 46894 37307 46950 37322
rect 46984 37318 47300 37322
rect 46984 37307 47051 37318
rect 45898 37284 47051 37307
rect 47085 37284 47204 37318
rect 47238 37307 47300 37318
rect 47334 37307 47390 37322
rect 47424 37307 47480 37322
rect 47514 37307 47570 37322
rect 47604 37307 47660 37322
rect 47694 37307 47750 37322
rect 47784 37307 47840 37322
rect 47874 37307 47930 37322
rect 47964 37307 48020 37322
rect 48054 37307 48110 37322
rect 48144 37307 48200 37322
rect 48234 37307 48290 37322
rect 48324 37318 48640 37322
rect 48324 37307 48391 37318
rect 47238 37284 48391 37307
rect 48425 37284 48544 37318
rect 48578 37307 48640 37318
rect 48674 37307 48730 37322
rect 48764 37307 48820 37322
rect 48854 37307 48910 37322
rect 48944 37307 49000 37322
rect 49034 37307 49090 37322
rect 49124 37307 49180 37322
rect 49214 37307 49270 37322
rect 49304 37307 49360 37322
rect 49394 37307 49450 37322
rect 49484 37307 49540 37322
rect 49574 37307 49630 37322
rect 49664 37318 49980 37322
rect 49664 37307 49731 37318
rect 48578 37284 49731 37307
rect 49765 37284 49884 37318
rect 49918 37307 49980 37318
rect 50014 37307 50070 37322
rect 50104 37307 50160 37322
rect 50194 37307 50250 37322
rect 50284 37307 50340 37322
rect 50374 37307 50430 37322
rect 50464 37307 50520 37322
rect 50554 37307 50610 37322
rect 50644 37307 50700 37322
rect 50734 37307 50790 37322
rect 50824 37307 50880 37322
rect 50914 37307 50970 37322
rect 51004 37318 51320 37322
rect 51004 37307 51071 37318
rect 49918 37284 51071 37307
rect 51105 37284 51224 37318
rect 51258 37307 51320 37318
rect 51354 37307 51410 37322
rect 51444 37307 51500 37322
rect 51534 37307 51590 37322
rect 51624 37307 51680 37322
rect 51714 37307 51770 37322
rect 51804 37307 51860 37322
rect 51894 37307 51950 37322
rect 51984 37307 52040 37322
rect 52074 37307 52130 37322
rect 52164 37307 52220 37322
rect 52254 37307 52310 37322
rect 52344 37318 52478 37322
rect 52344 37307 52411 37318
rect 51258 37284 52411 37307
rect 52445 37284 52478 37318
rect 41810 37277 52478 37284
rect 41810 37228 41909 37277
rect 41810 37194 41844 37228
rect 41878 37194 41909 37228
rect 42999 37228 43249 37277
rect 41810 37138 41909 37194
rect 41810 37104 41844 37138
rect 41878 37104 41909 37138
rect 41810 37048 41909 37104
rect 41810 37014 41844 37048
rect 41878 37014 41909 37048
rect 41810 36958 41909 37014
rect 41810 36924 41844 36958
rect 41878 36924 41909 36958
rect 41810 36868 41909 36924
rect 41810 36834 41844 36868
rect 41878 36834 41909 36868
rect 41810 36778 41909 36834
rect 41810 36744 41844 36778
rect 41878 36744 41909 36778
rect 41810 36688 41909 36744
rect 41810 36654 41844 36688
rect 41878 36654 41909 36688
rect 41810 36598 41909 36654
rect 41810 36564 41844 36598
rect 41878 36564 41909 36598
rect 41810 36508 41909 36564
rect 41810 36474 41844 36508
rect 41878 36474 41909 36508
rect 41810 36418 41909 36474
rect 41810 36384 41844 36418
rect 41878 36384 41909 36418
rect 41810 36328 41909 36384
rect 41810 36294 41844 36328
rect 41878 36294 41909 36328
rect 41810 36238 41909 36294
rect 41973 37196 42935 37213
rect 41973 37162 41994 37196
rect 42028 37162 42084 37196
rect 42118 37194 42174 37196
rect 42208 37194 42264 37196
rect 42298 37194 42354 37196
rect 42388 37194 42444 37196
rect 42478 37194 42534 37196
rect 42568 37194 42624 37196
rect 42658 37194 42714 37196
rect 42748 37194 42804 37196
rect 42838 37194 42894 37196
rect 42138 37162 42174 37194
rect 42228 37162 42264 37194
rect 42318 37162 42354 37194
rect 42408 37162 42444 37194
rect 42498 37162 42534 37194
rect 42588 37162 42624 37194
rect 42678 37162 42714 37194
rect 42768 37162 42804 37194
rect 42858 37162 42894 37194
rect 42928 37162 42935 37196
rect 41973 37160 42104 37162
rect 42138 37160 42194 37162
rect 42228 37160 42284 37162
rect 42318 37160 42374 37162
rect 42408 37160 42464 37162
rect 42498 37160 42554 37162
rect 42588 37160 42644 37162
rect 42678 37160 42734 37162
rect 42768 37160 42824 37162
rect 42858 37160 42935 37162
rect 41973 37141 42935 37160
rect 41973 37137 42045 37141
rect 41973 37103 41992 37137
rect 42026 37103 42045 37137
rect 41973 37047 42045 37103
rect 42863 37118 42935 37141
rect 42863 37084 42882 37118
rect 42916 37084 42935 37118
rect 41973 37013 41992 37047
rect 42026 37013 42045 37047
rect 41973 36957 42045 37013
rect 41973 36923 41992 36957
rect 42026 36923 42045 36957
rect 41973 36867 42045 36923
rect 41973 36833 41992 36867
rect 42026 36833 42045 36867
rect 41973 36777 42045 36833
rect 41973 36743 41992 36777
rect 42026 36743 42045 36777
rect 41973 36687 42045 36743
rect 41973 36653 41992 36687
rect 42026 36653 42045 36687
rect 41973 36597 42045 36653
rect 41973 36563 41992 36597
rect 42026 36563 42045 36597
rect 41973 36507 42045 36563
rect 41973 36473 41992 36507
rect 42026 36473 42045 36507
rect 41973 36417 42045 36473
rect 41973 36383 41992 36417
rect 42026 36383 42045 36417
rect 42107 37020 42801 37079
rect 42107 36986 42168 37020
rect 42202 36992 42258 37020
rect 42292 36992 42348 37020
rect 42382 36992 42438 37020
rect 42214 36986 42258 36992
rect 42314 36986 42348 36992
rect 42414 36986 42438 36992
rect 42472 36992 42528 37020
rect 42472 36986 42480 36992
rect 42107 36958 42180 36986
rect 42214 36958 42280 36986
rect 42314 36958 42380 36986
rect 42414 36958 42480 36986
rect 42514 36986 42528 36992
rect 42562 36992 42618 37020
rect 42562 36986 42580 36992
rect 42514 36958 42580 36986
rect 42614 36986 42618 36992
rect 42652 36992 42708 37020
rect 42652 36986 42680 36992
rect 42742 36986 42801 37020
rect 42614 36958 42680 36986
rect 42714 36958 42801 36986
rect 42107 36930 42801 36958
rect 42107 36896 42168 36930
rect 42202 36896 42258 36930
rect 42292 36896 42348 36930
rect 42382 36896 42438 36930
rect 42472 36896 42528 36930
rect 42562 36896 42618 36930
rect 42652 36896 42708 36930
rect 42742 36896 42801 36930
rect 42107 36892 42801 36896
rect 42107 36858 42180 36892
rect 42214 36858 42280 36892
rect 42314 36858 42380 36892
rect 42414 36858 42480 36892
rect 42514 36858 42580 36892
rect 42614 36858 42680 36892
rect 42714 36858 42801 36892
rect 42107 36840 42801 36858
rect 42107 36806 42168 36840
rect 42202 36806 42258 36840
rect 42292 36806 42348 36840
rect 42382 36806 42438 36840
rect 42472 36806 42528 36840
rect 42562 36806 42618 36840
rect 42652 36806 42708 36840
rect 42742 36806 42801 36840
rect 42107 36792 42801 36806
rect 42107 36758 42180 36792
rect 42214 36758 42280 36792
rect 42314 36758 42380 36792
rect 42414 36758 42480 36792
rect 42514 36758 42580 36792
rect 42614 36758 42680 36792
rect 42714 36758 42801 36792
rect 42107 36750 42801 36758
rect 42107 36716 42168 36750
rect 42202 36716 42258 36750
rect 42292 36716 42348 36750
rect 42382 36716 42438 36750
rect 42472 36716 42528 36750
rect 42562 36716 42618 36750
rect 42652 36716 42708 36750
rect 42742 36716 42801 36750
rect 42107 36692 42801 36716
rect 42107 36660 42180 36692
rect 42214 36660 42280 36692
rect 42314 36660 42380 36692
rect 42414 36660 42480 36692
rect 42107 36626 42168 36660
rect 42214 36658 42258 36660
rect 42314 36658 42348 36660
rect 42414 36658 42438 36660
rect 42202 36626 42258 36658
rect 42292 36626 42348 36658
rect 42382 36626 42438 36658
rect 42472 36658 42480 36660
rect 42514 36660 42580 36692
rect 42514 36658 42528 36660
rect 42472 36626 42528 36658
rect 42562 36658 42580 36660
rect 42614 36660 42680 36692
rect 42714 36660 42801 36692
rect 42614 36658 42618 36660
rect 42562 36626 42618 36658
rect 42652 36658 42680 36660
rect 42652 36626 42708 36658
rect 42742 36626 42801 36660
rect 42107 36592 42801 36626
rect 42107 36570 42180 36592
rect 42214 36570 42280 36592
rect 42314 36570 42380 36592
rect 42414 36570 42480 36592
rect 42107 36536 42168 36570
rect 42214 36558 42258 36570
rect 42314 36558 42348 36570
rect 42414 36558 42438 36570
rect 42202 36536 42258 36558
rect 42292 36536 42348 36558
rect 42382 36536 42438 36558
rect 42472 36558 42480 36570
rect 42514 36570 42580 36592
rect 42514 36558 42528 36570
rect 42472 36536 42528 36558
rect 42562 36558 42580 36570
rect 42614 36570 42680 36592
rect 42714 36570 42801 36592
rect 42614 36558 42618 36570
rect 42562 36536 42618 36558
rect 42652 36558 42680 36570
rect 42652 36536 42708 36558
rect 42742 36536 42801 36570
rect 42107 36492 42801 36536
rect 42107 36480 42180 36492
rect 42214 36480 42280 36492
rect 42314 36480 42380 36492
rect 42414 36480 42480 36492
rect 42107 36446 42168 36480
rect 42214 36458 42258 36480
rect 42314 36458 42348 36480
rect 42414 36458 42438 36480
rect 42202 36446 42258 36458
rect 42292 36446 42348 36458
rect 42382 36446 42438 36458
rect 42472 36458 42480 36480
rect 42514 36480 42580 36492
rect 42514 36458 42528 36480
rect 42472 36446 42528 36458
rect 42562 36458 42580 36480
rect 42614 36480 42680 36492
rect 42714 36480 42801 36492
rect 42614 36458 42618 36480
rect 42562 36446 42618 36458
rect 42652 36458 42680 36480
rect 42652 36446 42708 36458
rect 42742 36446 42801 36480
rect 42107 36385 42801 36446
rect 42863 37028 42935 37084
rect 42863 36994 42882 37028
rect 42916 36994 42935 37028
rect 42863 36938 42935 36994
rect 42863 36904 42882 36938
rect 42916 36904 42935 36938
rect 42863 36848 42935 36904
rect 42863 36814 42882 36848
rect 42916 36814 42935 36848
rect 42863 36758 42935 36814
rect 42863 36724 42882 36758
rect 42916 36724 42935 36758
rect 42863 36668 42935 36724
rect 42863 36634 42882 36668
rect 42916 36634 42935 36668
rect 42863 36578 42935 36634
rect 42863 36544 42882 36578
rect 42916 36544 42935 36578
rect 42863 36488 42935 36544
rect 42863 36454 42882 36488
rect 42916 36454 42935 36488
rect 42863 36398 42935 36454
rect 41973 36323 42045 36383
rect 42863 36364 42882 36398
rect 42916 36364 42935 36398
rect 42863 36323 42935 36364
rect 41973 36304 42935 36323
rect 41973 36270 42070 36304
rect 42104 36270 42160 36304
rect 42194 36270 42250 36304
rect 42284 36270 42340 36304
rect 42374 36270 42430 36304
rect 42464 36270 42520 36304
rect 42554 36270 42610 36304
rect 42644 36270 42700 36304
rect 42734 36270 42790 36304
rect 42824 36270 42935 36304
rect 41973 36251 42935 36270
rect 42999 37194 43031 37228
rect 43065 37194 43184 37228
rect 43218 37194 43249 37228
rect 44339 37228 44589 37277
rect 42999 37138 43249 37194
rect 42999 37104 43031 37138
rect 43065 37104 43184 37138
rect 43218 37104 43249 37138
rect 42999 37048 43249 37104
rect 42999 37014 43031 37048
rect 43065 37014 43184 37048
rect 43218 37014 43249 37048
rect 42999 36958 43249 37014
rect 42999 36924 43031 36958
rect 43065 36924 43184 36958
rect 43218 36924 43249 36958
rect 42999 36868 43249 36924
rect 42999 36834 43031 36868
rect 43065 36834 43184 36868
rect 43218 36834 43249 36868
rect 42999 36778 43249 36834
rect 42999 36744 43031 36778
rect 43065 36744 43184 36778
rect 43218 36744 43249 36778
rect 42999 36688 43249 36744
rect 42999 36654 43031 36688
rect 43065 36654 43184 36688
rect 43218 36654 43249 36688
rect 42999 36598 43249 36654
rect 42999 36564 43031 36598
rect 43065 36564 43184 36598
rect 43218 36564 43249 36598
rect 42999 36508 43249 36564
rect 42999 36474 43031 36508
rect 43065 36474 43184 36508
rect 43218 36474 43249 36508
rect 42999 36418 43249 36474
rect 42999 36384 43031 36418
rect 43065 36384 43184 36418
rect 43218 36384 43249 36418
rect 42999 36328 43249 36384
rect 42999 36294 43031 36328
rect 43065 36294 43184 36328
rect 43218 36294 43249 36328
rect 41810 36204 41844 36238
rect 41878 36204 41909 36238
rect 41810 36187 41909 36204
rect 42999 36238 43249 36294
rect 43313 37196 44275 37213
rect 43313 37162 43334 37196
rect 43368 37162 43424 37196
rect 43458 37194 43514 37196
rect 43548 37194 43604 37196
rect 43638 37194 43694 37196
rect 43728 37194 43784 37196
rect 43818 37194 43874 37196
rect 43908 37194 43964 37196
rect 43998 37194 44054 37196
rect 44088 37194 44144 37196
rect 44178 37194 44234 37196
rect 43478 37162 43514 37194
rect 43568 37162 43604 37194
rect 43658 37162 43694 37194
rect 43748 37162 43784 37194
rect 43838 37162 43874 37194
rect 43928 37162 43964 37194
rect 44018 37162 44054 37194
rect 44108 37162 44144 37194
rect 44198 37162 44234 37194
rect 44268 37162 44275 37196
rect 43313 37160 43444 37162
rect 43478 37160 43534 37162
rect 43568 37160 43624 37162
rect 43658 37160 43714 37162
rect 43748 37160 43804 37162
rect 43838 37160 43894 37162
rect 43928 37160 43984 37162
rect 44018 37160 44074 37162
rect 44108 37160 44164 37162
rect 44198 37160 44275 37162
rect 43313 37141 44275 37160
rect 43313 37137 43385 37141
rect 43313 37103 43332 37137
rect 43366 37103 43385 37137
rect 43313 37047 43385 37103
rect 44203 37118 44275 37141
rect 44203 37084 44222 37118
rect 44256 37084 44275 37118
rect 43313 37013 43332 37047
rect 43366 37013 43385 37047
rect 43313 36957 43385 37013
rect 43313 36923 43332 36957
rect 43366 36923 43385 36957
rect 43313 36867 43385 36923
rect 43313 36833 43332 36867
rect 43366 36833 43385 36867
rect 43313 36777 43385 36833
rect 43313 36743 43332 36777
rect 43366 36743 43385 36777
rect 43313 36687 43385 36743
rect 43313 36653 43332 36687
rect 43366 36653 43385 36687
rect 43313 36597 43385 36653
rect 43313 36563 43332 36597
rect 43366 36563 43385 36597
rect 43313 36507 43385 36563
rect 43313 36473 43332 36507
rect 43366 36473 43385 36507
rect 43313 36417 43385 36473
rect 43313 36383 43332 36417
rect 43366 36383 43385 36417
rect 43447 37020 44141 37079
rect 43447 36986 43508 37020
rect 43542 36992 43598 37020
rect 43632 36992 43688 37020
rect 43722 36992 43778 37020
rect 43554 36986 43598 36992
rect 43654 36986 43688 36992
rect 43754 36986 43778 36992
rect 43812 36992 43868 37020
rect 43812 36986 43820 36992
rect 43447 36958 43520 36986
rect 43554 36958 43620 36986
rect 43654 36958 43720 36986
rect 43754 36958 43820 36986
rect 43854 36986 43868 36992
rect 43902 36992 43958 37020
rect 43902 36986 43920 36992
rect 43854 36958 43920 36986
rect 43954 36986 43958 36992
rect 43992 36992 44048 37020
rect 43992 36986 44020 36992
rect 44082 36986 44141 37020
rect 43954 36958 44020 36986
rect 44054 36958 44141 36986
rect 43447 36930 44141 36958
rect 43447 36896 43508 36930
rect 43542 36896 43598 36930
rect 43632 36896 43688 36930
rect 43722 36896 43778 36930
rect 43812 36896 43868 36930
rect 43902 36896 43958 36930
rect 43992 36896 44048 36930
rect 44082 36896 44141 36930
rect 43447 36892 44141 36896
rect 43447 36858 43520 36892
rect 43554 36858 43620 36892
rect 43654 36858 43720 36892
rect 43754 36858 43820 36892
rect 43854 36858 43920 36892
rect 43954 36858 44020 36892
rect 44054 36858 44141 36892
rect 43447 36840 44141 36858
rect 43447 36806 43508 36840
rect 43542 36806 43598 36840
rect 43632 36806 43688 36840
rect 43722 36806 43778 36840
rect 43812 36806 43868 36840
rect 43902 36806 43958 36840
rect 43992 36806 44048 36840
rect 44082 36806 44141 36840
rect 43447 36792 44141 36806
rect 43447 36758 43520 36792
rect 43554 36758 43620 36792
rect 43654 36758 43720 36792
rect 43754 36758 43820 36792
rect 43854 36758 43920 36792
rect 43954 36758 44020 36792
rect 44054 36758 44141 36792
rect 43447 36750 44141 36758
rect 43447 36716 43508 36750
rect 43542 36716 43598 36750
rect 43632 36716 43688 36750
rect 43722 36716 43778 36750
rect 43812 36716 43868 36750
rect 43902 36716 43958 36750
rect 43992 36716 44048 36750
rect 44082 36716 44141 36750
rect 43447 36692 44141 36716
rect 43447 36660 43520 36692
rect 43554 36660 43620 36692
rect 43654 36660 43720 36692
rect 43754 36660 43820 36692
rect 43447 36626 43508 36660
rect 43554 36658 43598 36660
rect 43654 36658 43688 36660
rect 43754 36658 43778 36660
rect 43542 36626 43598 36658
rect 43632 36626 43688 36658
rect 43722 36626 43778 36658
rect 43812 36658 43820 36660
rect 43854 36660 43920 36692
rect 43854 36658 43868 36660
rect 43812 36626 43868 36658
rect 43902 36658 43920 36660
rect 43954 36660 44020 36692
rect 44054 36660 44141 36692
rect 43954 36658 43958 36660
rect 43902 36626 43958 36658
rect 43992 36658 44020 36660
rect 43992 36626 44048 36658
rect 44082 36626 44141 36660
rect 43447 36592 44141 36626
rect 43447 36570 43520 36592
rect 43554 36570 43620 36592
rect 43654 36570 43720 36592
rect 43754 36570 43820 36592
rect 43447 36536 43508 36570
rect 43554 36558 43598 36570
rect 43654 36558 43688 36570
rect 43754 36558 43778 36570
rect 43542 36536 43598 36558
rect 43632 36536 43688 36558
rect 43722 36536 43778 36558
rect 43812 36558 43820 36570
rect 43854 36570 43920 36592
rect 43854 36558 43868 36570
rect 43812 36536 43868 36558
rect 43902 36558 43920 36570
rect 43954 36570 44020 36592
rect 44054 36570 44141 36592
rect 43954 36558 43958 36570
rect 43902 36536 43958 36558
rect 43992 36558 44020 36570
rect 43992 36536 44048 36558
rect 44082 36536 44141 36570
rect 43447 36492 44141 36536
rect 43447 36480 43520 36492
rect 43554 36480 43620 36492
rect 43654 36480 43720 36492
rect 43754 36480 43820 36492
rect 43447 36446 43508 36480
rect 43554 36458 43598 36480
rect 43654 36458 43688 36480
rect 43754 36458 43778 36480
rect 43542 36446 43598 36458
rect 43632 36446 43688 36458
rect 43722 36446 43778 36458
rect 43812 36458 43820 36480
rect 43854 36480 43920 36492
rect 43854 36458 43868 36480
rect 43812 36446 43868 36458
rect 43902 36458 43920 36480
rect 43954 36480 44020 36492
rect 44054 36480 44141 36492
rect 43954 36458 43958 36480
rect 43902 36446 43958 36458
rect 43992 36458 44020 36480
rect 43992 36446 44048 36458
rect 44082 36446 44141 36480
rect 43447 36385 44141 36446
rect 44203 37028 44275 37084
rect 44203 36994 44222 37028
rect 44256 36994 44275 37028
rect 44203 36938 44275 36994
rect 44203 36904 44222 36938
rect 44256 36904 44275 36938
rect 44203 36848 44275 36904
rect 44203 36814 44222 36848
rect 44256 36814 44275 36848
rect 44203 36758 44275 36814
rect 44203 36724 44222 36758
rect 44256 36724 44275 36758
rect 44203 36668 44275 36724
rect 44203 36634 44222 36668
rect 44256 36634 44275 36668
rect 44203 36578 44275 36634
rect 44203 36544 44222 36578
rect 44256 36544 44275 36578
rect 44203 36488 44275 36544
rect 44203 36454 44222 36488
rect 44256 36454 44275 36488
rect 44203 36398 44275 36454
rect 43313 36323 43385 36383
rect 44203 36364 44222 36398
rect 44256 36364 44275 36398
rect 44203 36323 44275 36364
rect 43313 36304 44275 36323
rect 43313 36270 43410 36304
rect 43444 36270 43500 36304
rect 43534 36270 43590 36304
rect 43624 36270 43680 36304
rect 43714 36270 43770 36304
rect 43804 36270 43860 36304
rect 43894 36270 43950 36304
rect 43984 36270 44040 36304
rect 44074 36270 44130 36304
rect 44164 36270 44275 36304
rect 43313 36251 44275 36270
rect 44339 37194 44371 37228
rect 44405 37194 44524 37228
rect 44558 37194 44589 37228
rect 45679 37228 45929 37277
rect 44339 37138 44589 37194
rect 44339 37104 44371 37138
rect 44405 37104 44524 37138
rect 44558 37104 44589 37138
rect 44339 37048 44589 37104
rect 44339 37014 44371 37048
rect 44405 37014 44524 37048
rect 44558 37014 44589 37048
rect 44339 36958 44589 37014
rect 44339 36924 44371 36958
rect 44405 36924 44524 36958
rect 44558 36924 44589 36958
rect 44339 36868 44589 36924
rect 44339 36834 44371 36868
rect 44405 36834 44524 36868
rect 44558 36834 44589 36868
rect 44339 36778 44589 36834
rect 44339 36744 44371 36778
rect 44405 36744 44524 36778
rect 44558 36744 44589 36778
rect 44339 36688 44589 36744
rect 44339 36654 44371 36688
rect 44405 36654 44524 36688
rect 44558 36654 44589 36688
rect 44339 36598 44589 36654
rect 44339 36564 44371 36598
rect 44405 36564 44524 36598
rect 44558 36564 44589 36598
rect 44339 36508 44589 36564
rect 44339 36474 44371 36508
rect 44405 36474 44524 36508
rect 44558 36474 44589 36508
rect 44339 36418 44589 36474
rect 44339 36384 44371 36418
rect 44405 36384 44524 36418
rect 44558 36384 44589 36418
rect 44339 36328 44589 36384
rect 44339 36294 44371 36328
rect 44405 36294 44524 36328
rect 44558 36294 44589 36328
rect 42999 36204 43031 36238
rect 43065 36204 43184 36238
rect 43218 36204 43249 36238
rect 42999 36187 43249 36204
rect 44339 36238 44589 36294
rect 44653 37196 45615 37213
rect 44653 37162 44674 37196
rect 44708 37162 44764 37196
rect 44798 37194 44854 37196
rect 44888 37194 44944 37196
rect 44978 37194 45034 37196
rect 45068 37194 45124 37196
rect 45158 37194 45214 37196
rect 45248 37194 45304 37196
rect 45338 37194 45394 37196
rect 45428 37194 45484 37196
rect 45518 37194 45574 37196
rect 44818 37162 44854 37194
rect 44908 37162 44944 37194
rect 44998 37162 45034 37194
rect 45088 37162 45124 37194
rect 45178 37162 45214 37194
rect 45268 37162 45304 37194
rect 45358 37162 45394 37194
rect 45448 37162 45484 37194
rect 45538 37162 45574 37194
rect 45608 37162 45615 37196
rect 44653 37160 44784 37162
rect 44818 37160 44874 37162
rect 44908 37160 44964 37162
rect 44998 37160 45054 37162
rect 45088 37160 45144 37162
rect 45178 37160 45234 37162
rect 45268 37160 45324 37162
rect 45358 37160 45414 37162
rect 45448 37160 45504 37162
rect 45538 37160 45615 37162
rect 44653 37141 45615 37160
rect 44653 37137 44725 37141
rect 44653 37103 44672 37137
rect 44706 37103 44725 37137
rect 44653 37047 44725 37103
rect 45543 37118 45615 37141
rect 45543 37084 45562 37118
rect 45596 37084 45615 37118
rect 44653 37013 44672 37047
rect 44706 37013 44725 37047
rect 44653 36957 44725 37013
rect 44653 36923 44672 36957
rect 44706 36923 44725 36957
rect 44653 36867 44725 36923
rect 44653 36833 44672 36867
rect 44706 36833 44725 36867
rect 44653 36777 44725 36833
rect 44653 36743 44672 36777
rect 44706 36743 44725 36777
rect 44653 36687 44725 36743
rect 44653 36653 44672 36687
rect 44706 36653 44725 36687
rect 44653 36597 44725 36653
rect 44653 36563 44672 36597
rect 44706 36563 44725 36597
rect 44653 36507 44725 36563
rect 44653 36473 44672 36507
rect 44706 36473 44725 36507
rect 44653 36417 44725 36473
rect 44653 36383 44672 36417
rect 44706 36383 44725 36417
rect 44787 37020 45481 37079
rect 44787 36986 44848 37020
rect 44882 36992 44938 37020
rect 44972 36992 45028 37020
rect 45062 36992 45118 37020
rect 44894 36986 44938 36992
rect 44994 36986 45028 36992
rect 45094 36986 45118 36992
rect 45152 36992 45208 37020
rect 45152 36986 45160 36992
rect 44787 36958 44860 36986
rect 44894 36958 44960 36986
rect 44994 36958 45060 36986
rect 45094 36958 45160 36986
rect 45194 36986 45208 36992
rect 45242 36992 45298 37020
rect 45242 36986 45260 36992
rect 45194 36958 45260 36986
rect 45294 36986 45298 36992
rect 45332 36992 45388 37020
rect 45332 36986 45360 36992
rect 45422 36986 45481 37020
rect 45294 36958 45360 36986
rect 45394 36958 45481 36986
rect 44787 36930 45481 36958
rect 44787 36896 44848 36930
rect 44882 36896 44938 36930
rect 44972 36896 45028 36930
rect 45062 36896 45118 36930
rect 45152 36896 45208 36930
rect 45242 36896 45298 36930
rect 45332 36896 45388 36930
rect 45422 36896 45481 36930
rect 44787 36892 45481 36896
rect 44787 36858 44860 36892
rect 44894 36858 44960 36892
rect 44994 36858 45060 36892
rect 45094 36858 45160 36892
rect 45194 36858 45260 36892
rect 45294 36858 45360 36892
rect 45394 36858 45481 36892
rect 44787 36840 45481 36858
rect 44787 36806 44848 36840
rect 44882 36806 44938 36840
rect 44972 36806 45028 36840
rect 45062 36806 45118 36840
rect 45152 36806 45208 36840
rect 45242 36806 45298 36840
rect 45332 36806 45388 36840
rect 45422 36806 45481 36840
rect 44787 36792 45481 36806
rect 44787 36758 44860 36792
rect 44894 36758 44960 36792
rect 44994 36758 45060 36792
rect 45094 36758 45160 36792
rect 45194 36758 45260 36792
rect 45294 36758 45360 36792
rect 45394 36758 45481 36792
rect 44787 36750 45481 36758
rect 44787 36716 44848 36750
rect 44882 36716 44938 36750
rect 44972 36716 45028 36750
rect 45062 36716 45118 36750
rect 45152 36716 45208 36750
rect 45242 36716 45298 36750
rect 45332 36716 45388 36750
rect 45422 36716 45481 36750
rect 44787 36692 45481 36716
rect 44787 36660 44860 36692
rect 44894 36660 44960 36692
rect 44994 36660 45060 36692
rect 45094 36660 45160 36692
rect 44787 36626 44848 36660
rect 44894 36658 44938 36660
rect 44994 36658 45028 36660
rect 45094 36658 45118 36660
rect 44882 36626 44938 36658
rect 44972 36626 45028 36658
rect 45062 36626 45118 36658
rect 45152 36658 45160 36660
rect 45194 36660 45260 36692
rect 45194 36658 45208 36660
rect 45152 36626 45208 36658
rect 45242 36658 45260 36660
rect 45294 36660 45360 36692
rect 45394 36660 45481 36692
rect 45294 36658 45298 36660
rect 45242 36626 45298 36658
rect 45332 36658 45360 36660
rect 45332 36626 45388 36658
rect 45422 36626 45481 36660
rect 44787 36592 45481 36626
rect 44787 36570 44860 36592
rect 44894 36570 44960 36592
rect 44994 36570 45060 36592
rect 45094 36570 45160 36592
rect 44787 36536 44848 36570
rect 44894 36558 44938 36570
rect 44994 36558 45028 36570
rect 45094 36558 45118 36570
rect 44882 36536 44938 36558
rect 44972 36536 45028 36558
rect 45062 36536 45118 36558
rect 45152 36558 45160 36570
rect 45194 36570 45260 36592
rect 45194 36558 45208 36570
rect 45152 36536 45208 36558
rect 45242 36558 45260 36570
rect 45294 36570 45360 36592
rect 45394 36570 45481 36592
rect 45294 36558 45298 36570
rect 45242 36536 45298 36558
rect 45332 36558 45360 36570
rect 45332 36536 45388 36558
rect 45422 36536 45481 36570
rect 44787 36492 45481 36536
rect 44787 36480 44860 36492
rect 44894 36480 44960 36492
rect 44994 36480 45060 36492
rect 45094 36480 45160 36492
rect 44787 36446 44848 36480
rect 44894 36458 44938 36480
rect 44994 36458 45028 36480
rect 45094 36458 45118 36480
rect 44882 36446 44938 36458
rect 44972 36446 45028 36458
rect 45062 36446 45118 36458
rect 45152 36458 45160 36480
rect 45194 36480 45260 36492
rect 45194 36458 45208 36480
rect 45152 36446 45208 36458
rect 45242 36458 45260 36480
rect 45294 36480 45360 36492
rect 45394 36480 45481 36492
rect 45294 36458 45298 36480
rect 45242 36446 45298 36458
rect 45332 36458 45360 36480
rect 45332 36446 45388 36458
rect 45422 36446 45481 36480
rect 44787 36385 45481 36446
rect 45543 37028 45615 37084
rect 45543 36994 45562 37028
rect 45596 36994 45615 37028
rect 45543 36938 45615 36994
rect 45543 36904 45562 36938
rect 45596 36904 45615 36938
rect 45543 36848 45615 36904
rect 45543 36814 45562 36848
rect 45596 36814 45615 36848
rect 45543 36758 45615 36814
rect 45543 36724 45562 36758
rect 45596 36724 45615 36758
rect 45543 36668 45615 36724
rect 45543 36634 45562 36668
rect 45596 36634 45615 36668
rect 45543 36578 45615 36634
rect 45543 36544 45562 36578
rect 45596 36544 45615 36578
rect 45543 36488 45615 36544
rect 45543 36454 45562 36488
rect 45596 36454 45615 36488
rect 45543 36398 45615 36454
rect 44653 36323 44725 36383
rect 45543 36364 45562 36398
rect 45596 36364 45615 36398
rect 45543 36323 45615 36364
rect 44653 36304 45615 36323
rect 44653 36270 44750 36304
rect 44784 36270 44840 36304
rect 44874 36270 44930 36304
rect 44964 36270 45020 36304
rect 45054 36270 45110 36304
rect 45144 36270 45200 36304
rect 45234 36270 45290 36304
rect 45324 36270 45380 36304
rect 45414 36270 45470 36304
rect 45504 36270 45615 36304
rect 44653 36251 45615 36270
rect 45679 37194 45711 37228
rect 45745 37194 45864 37228
rect 45898 37194 45929 37228
rect 47019 37228 47269 37277
rect 45679 37138 45929 37194
rect 45679 37104 45711 37138
rect 45745 37104 45864 37138
rect 45898 37104 45929 37138
rect 45679 37048 45929 37104
rect 45679 37014 45711 37048
rect 45745 37014 45864 37048
rect 45898 37014 45929 37048
rect 45679 36958 45929 37014
rect 45679 36924 45711 36958
rect 45745 36924 45864 36958
rect 45898 36924 45929 36958
rect 45679 36868 45929 36924
rect 45679 36834 45711 36868
rect 45745 36834 45864 36868
rect 45898 36834 45929 36868
rect 45679 36778 45929 36834
rect 45679 36744 45711 36778
rect 45745 36744 45864 36778
rect 45898 36744 45929 36778
rect 45679 36688 45929 36744
rect 45679 36654 45711 36688
rect 45745 36654 45864 36688
rect 45898 36654 45929 36688
rect 45679 36598 45929 36654
rect 45679 36564 45711 36598
rect 45745 36564 45864 36598
rect 45898 36564 45929 36598
rect 45679 36508 45929 36564
rect 45679 36474 45711 36508
rect 45745 36474 45864 36508
rect 45898 36474 45929 36508
rect 45679 36418 45929 36474
rect 45679 36384 45711 36418
rect 45745 36384 45864 36418
rect 45898 36384 45929 36418
rect 45679 36328 45929 36384
rect 45679 36294 45711 36328
rect 45745 36294 45864 36328
rect 45898 36294 45929 36328
rect 44339 36204 44371 36238
rect 44405 36204 44524 36238
rect 44558 36204 44589 36238
rect 44339 36187 44589 36204
rect 45679 36238 45929 36294
rect 45993 37196 46955 37213
rect 45993 37162 46014 37196
rect 46048 37162 46104 37196
rect 46138 37194 46194 37196
rect 46228 37194 46284 37196
rect 46318 37194 46374 37196
rect 46408 37194 46464 37196
rect 46498 37194 46554 37196
rect 46588 37194 46644 37196
rect 46678 37194 46734 37196
rect 46768 37194 46824 37196
rect 46858 37194 46914 37196
rect 46158 37162 46194 37194
rect 46248 37162 46284 37194
rect 46338 37162 46374 37194
rect 46428 37162 46464 37194
rect 46518 37162 46554 37194
rect 46608 37162 46644 37194
rect 46698 37162 46734 37194
rect 46788 37162 46824 37194
rect 46878 37162 46914 37194
rect 46948 37162 46955 37196
rect 45993 37160 46124 37162
rect 46158 37160 46214 37162
rect 46248 37160 46304 37162
rect 46338 37160 46394 37162
rect 46428 37160 46484 37162
rect 46518 37160 46574 37162
rect 46608 37160 46664 37162
rect 46698 37160 46754 37162
rect 46788 37160 46844 37162
rect 46878 37160 46955 37162
rect 45993 37141 46955 37160
rect 45993 37137 46065 37141
rect 45993 37103 46012 37137
rect 46046 37103 46065 37137
rect 45993 37047 46065 37103
rect 46883 37118 46955 37141
rect 46883 37084 46902 37118
rect 46936 37084 46955 37118
rect 45993 37013 46012 37047
rect 46046 37013 46065 37047
rect 45993 36957 46065 37013
rect 45993 36923 46012 36957
rect 46046 36923 46065 36957
rect 45993 36867 46065 36923
rect 45993 36833 46012 36867
rect 46046 36833 46065 36867
rect 45993 36777 46065 36833
rect 45993 36743 46012 36777
rect 46046 36743 46065 36777
rect 45993 36687 46065 36743
rect 45993 36653 46012 36687
rect 46046 36653 46065 36687
rect 45993 36597 46065 36653
rect 45993 36563 46012 36597
rect 46046 36563 46065 36597
rect 45993 36507 46065 36563
rect 45993 36473 46012 36507
rect 46046 36473 46065 36507
rect 45993 36417 46065 36473
rect 45993 36383 46012 36417
rect 46046 36383 46065 36417
rect 46127 37020 46821 37079
rect 46127 36986 46188 37020
rect 46222 36992 46278 37020
rect 46312 36992 46368 37020
rect 46402 36992 46458 37020
rect 46234 36986 46278 36992
rect 46334 36986 46368 36992
rect 46434 36986 46458 36992
rect 46492 36992 46548 37020
rect 46492 36986 46500 36992
rect 46127 36958 46200 36986
rect 46234 36958 46300 36986
rect 46334 36958 46400 36986
rect 46434 36958 46500 36986
rect 46534 36986 46548 36992
rect 46582 36992 46638 37020
rect 46582 36986 46600 36992
rect 46534 36958 46600 36986
rect 46634 36986 46638 36992
rect 46672 36992 46728 37020
rect 46672 36986 46700 36992
rect 46762 36986 46821 37020
rect 46634 36958 46700 36986
rect 46734 36958 46821 36986
rect 46127 36930 46821 36958
rect 46127 36896 46188 36930
rect 46222 36896 46278 36930
rect 46312 36896 46368 36930
rect 46402 36896 46458 36930
rect 46492 36896 46548 36930
rect 46582 36896 46638 36930
rect 46672 36896 46728 36930
rect 46762 36896 46821 36930
rect 46127 36892 46821 36896
rect 46127 36858 46200 36892
rect 46234 36858 46300 36892
rect 46334 36858 46400 36892
rect 46434 36858 46500 36892
rect 46534 36858 46600 36892
rect 46634 36858 46700 36892
rect 46734 36858 46821 36892
rect 46127 36840 46821 36858
rect 46127 36806 46188 36840
rect 46222 36806 46278 36840
rect 46312 36806 46368 36840
rect 46402 36806 46458 36840
rect 46492 36806 46548 36840
rect 46582 36806 46638 36840
rect 46672 36806 46728 36840
rect 46762 36806 46821 36840
rect 46127 36792 46821 36806
rect 46127 36758 46200 36792
rect 46234 36758 46300 36792
rect 46334 36758 46400 36792
rect 46434 36758 46500 36792
rect 46534 36758 46600 36792
rect 46634 36758 46700 36792
rect 46734 36758 46821 36792
rect 46127 36750 46821 36758
rect 46127 36716 46188 36750
rect 46222 36716 46278 36750
rect 46312 36716 46368 36750
rect 46402 36716 46458 36750
rect 46492 36716 46548 36750
rect 46582 36716 46638 36750
rect 46672 36716 46728 36750
rect 46762 36716 46821 36750
rect 46127 36692 46821 36716
rect 46127 36660 46200 36692
rect 46234 36660 46300 36692
rect 46334 36660 46400 36692
rect 46434 36660 46500 36692
rect 46127 36626 46188 36660
rect 46234 36658 46278 36660
rect 46334 36658 46368 36660
rect 46434 36658 46458 36660
rect 46222 36626 46278 36658
rect 46312 36626 46368 36658
rect 46402 36626 46458 36658
rect 46492 36658 46500 36660
rect 46534 36660 46600 36692
rect 46534 36658 46548 36660
rect 46492 36626 46548 36658
rect 46582 36658 46600 36660
rect 46634 36660 46700 36692
rect 46734 36660 46821 36692
rect 46634 36658 46638 36660
rect 46582 36626 46638 36658
rect 46672 36658 46700 36660
rect 46672 36626 46728 36658
rect 46762 36626 46821 36660
rect 46127 36592 46821 36626
rect 46127 36570 46200 36592
rect 46234 36570 46300 36592
rect 46334 36570 46400 36592
rect 46434 36570 46500 36592
rect 46127 36536 46188 36570
rect 46234 36558 46278 36570
rect 46334 36558 46368 36570
rect 46434 36558 46458 36570
rect 46222 36536 46278 36558
rect 46312 36536 46368 36558
rect 46402 36536 46458 36558
rect 46492 36558 46500 36570
rect 46534 36570 46600 36592
rect 46534 36558 46548 36570
rect 46492 36536 46548 36558
rect 46582 36558 46600 36570
rect 46634 36570 46700 36592
rect 46734 36570 46821 36592
rect 46634 36558 46638 36570
rect 46582 36536 46638 36558
rect 46672 36558 46700 36570
rect 46672 36536 46728 36558
rect 46762 36536 46821 36570
rect 46127 36492 46821 36536
rect 46127 36480 46200 36492
rect 46234 36480 46300 36492
rect 46334 36480 46400 36492
rect 46434 36480 46500 36492
rect 46127 36446 46188 36480
rect 46234 36458 46278 36480
rect 46334 36458 46368 36480
rect 46434 36458 46458 36480
rect 46222 36446 46278 36458
rect 46312 36446 46368 36458
rect 46402 36446 46458 36458
rect 46492 36458 46500 36480
rect 46534 36480 46600 36492
rect 46534 36458 46548 36480
rect 46492 36446 46548 36458
rect 46582 36458 46600 36480
rect 46634 36480 46700 36492
rect 46734 36480 46821 36492
rect 46634 36458 46638 36480
rect 46582 36446 46638 36458
rect 46672 36458 46700 36480
rect 46672 36446 46728 36458
rect 46762 36446 46821 36480
rect 46127 36385 46821 36446
rect 46883 37028 46955 37084
rect 46883 36994 46902 37028
rect 46936 36994 46955 37028
rect 46883 36938 46955 36994
rect 46883 36904 46902 36938
rect 46936 36904 46955 36938
rect 46883 36848 46955 36904
rect 46883 36814 46902 36848
rect 46936 36814 46955 36848
rect 46883 36758 46955 36814
rect 46883 36724 46902 36758
rect 46936 36724 46955 36758
rect 46883 36668 46955 36724
rect 46883 36634 46902 36668
rect 46936 36634 46955 36668
rect 46883 36578 46955 36634
rect 46883 36544 46902 36578
rect 46936 36544 46955 36578
rect 46883 36488 46955 36544
rect 46883 36454 46902 36488
rect 46936 36454 46955 36488
rect 46883 36398 46955 36454
rect 45993 36323 46065 36383
rect 46883 36364 46902 36398
rect 46936 36364 46955 36398
rect 46883 36323 46955 36364
rect 45993 36304 46955 36323
rect 45993 36270 46090 36304
rect 46124 36270 46180 36304
rect 46214 36270 46270 36304
rect 46304 36270 46360 36304
rect 46394 36270 46450 36304
rect 46484 36270 46540 36304
rect 46574 36270 46630 36304
rect 46664 36270 46720 36304
rect 46754 36270 46810 36304
rect 46844 36270 46955 36304
rect 45993 36251 46955 36270
rect 47019 37194 47051 37228
rect 47085 37194 47204 37228
rect 47238 37194 47269 37228
rect 48359 37228 48609 37277
rect 47019 37138 47269 37194
rect 47019 37104 47051 37138
rect 47085 37104 47204 37138
rect 47238 37104 47269 37138
rect 47019 37048 47269 37104
rect 47019 37014 47051 37048
rect 47085 37014 47204 37048
rect 47238 37014 47269 37048
rect 47019 36958 47269 37014
rect 47019 36924 47051 36958
rect 47085 36924 47204 36958
rect 47238 36924 47269 36958
rect 47019 36868 47269 36924
rect 47019 36834 47051 36868
rect 47085 36834 47204 36868
rect 47238 36834 47269 36868
rect 47019 36778 47269 36834
rect 47019 36744 47051 36778
rect 47085 36744 47204 36778
rect 47238 36744 47269 36778
rect 47019 36688 47269 36744
rect 47019 36654 47051 36688
rect 47085 36654 47204 36688
rect 47238 36654 47269 36688
rect 47019 36598 47269 36654
rect 47019 36564 47051 36598
rect 47085 36564 47204 36598
rect 47238 36564 47269 36598
rect 47019 36508 47269 36564
rect 47019 36474 47051 36508
rect 47085 36474 47204 36508
rect 47238 36474 47269 36508
rect 47019 36418 47269 36474
rect 47019 36384 47051 36418
rect 47085 36384 47204 36418
rect 47238 36384 47269 36418
rect 47019 36328 47269 36384
rect 47019 36294 47051 36328
rect 47085 36294 47204 36328
rect 47238 36294 47269 36328
rect 45679 36204 45711 36238
rect 45745 36204 45864 36238
rect 45898 36204 45929 36238
rect 45679 36187 45929 36204
rect 47019 36238 47269 36294
rect 47333 37196 48295 37213
rect 47333 37162 47354 37196
rect 47388 37162 47444 37196
rect 47478 37194 47534 37196
rect 47568 37194 47624 37196
rect 47658 37194 47714 37196
rect 47748 37194 47804 37196
rect 47838 37194 47894 37196
rect 47928 37194 47984 37196
rect 48018 37194 48074 37196
rect 48108 37194 48164 37196
rect 48198 37194 48254 37196
rect 47498 37162 47534 37194
rect 47588 37162 47624 37194
rect 47678 37162 47714 37194
rect 47768 37162 47804 37194
rect 47858 37162 47894 37194
rect 47948 37162 47984 37194
rect 48038 37162 48074 37194
rect 48128 37162 48164 37194
rect 48218 37162 48254 37194
rect 48288 37162 48295 37196
rect 47333 37160 47464 37162
rect 47498 37160 47554 37162
rect 47588 37160 47644 37162
rect 47678 37160 47734 37162
rect 47768 37160 47824 37162
rect 47858 37160 47914 37162
rect 47948 37160 48004 37162
rect 48038 37160 48094 37162
rect 48128 37160 48184 37162
rect 48218 37160 48295 37162
rect 47333 37141 48295 37160
rect 47333 37137 47405 37141
rect 47333 37103 47352 37137
rect 47386 37103 47405 37137
rect 47333 37047 47405 37103
rect 48223 37118 48295 37141
rect 48223 37084 48242 37118
rect 48276 37084 48295 37118
rect 47333 37013 47352 37047
rect 47386 37013 47405 37047
rect 47333 36957 47405 37013
rect 47333 36923 47352 36957
rect 47386 36923 47405 36957
rect 47333 36867 47405 36923
rect 47333 36833 47352 36867
rect 47386 36833 47405 36867
rect 47333 36777 47405 36833
rect 47333 36743 47352 36777
rect 47386 36743 47405 36777
rect 47333 36687 47405 36743
rect 47333 36653 47352 36687
rect 47386 36653 47405 36687
rect 47333 36597 47405 36653
rect 47333 36563 47352 36597
rect 47386 36563 47405 36597
rect 47333 36507 47405 36563
rect 47333 36473 47352 36507
rect 47386 36473 47405 36507
rect 47333 36417 47405 36473
rect 47333 36383 47352 36417
rect 47386 36383 47405 36417
rect 47467 37020 48161 37079
rect 47467 36986 47528 37020
rect 47562 36992 47618 37020
rect 47652 36992 47708 37020
rect 47742 36992 47798 37020
rect 47574 36986 47618 36992
rect 47674 36986 47708 36992
rect 47774 36986 47798 36992
rect 47832 36992 47888 37020
rect 47832 36986 47840 36992
rect 47467 36958 47540 36986
rect 47574 36958 47640 36986
rect 47674 36958 47740 36986
rect 47774 36958 47840 36986
rect 47874 36986 47888 36992
rect 47922 36992 47978 37020
rect 47922 36986 47940 36992
rect 47874 36958 47940 36986
rect 47974 36986 47978 36992
rect 48012 36992 48068 37020
rect 48012 36986 48040 36992
rect 48102 36986 48161 37020
rect 47974 36958 48040 36986
rect 48074 36958 48161 36986
rect 47467 36930 48161 36958
rect 47467 36896 47528 36930
rect 47562 36896 47618 36930
rect 47652 36896 47708 36930
rect 47742 36896 47798 36930
rect 47832 36896 47888 36930
rect 47922 36896 47978 36930
rect 48012 36896 48068 36930
rect 48102 36896 48161 36930
rect 47467 36892 48161 36896
rect 47467 36858 47540 36892
rect 47574 36858 47640 36892
rect 47674 36858 47740 36892
rect 47774 36858 47840 36892
rect 47874 36858 47940 36892
rect 47974 36858 48040 36892
rect 48074 36858 48161 36892
rect 47467 36840 48161 36858
rect 47467 36806 47528 36840
rect 47562 36806 47618 36840
rect 47652 36806 47708 36840
rect 47742 36806 47798 36840
rect 47832 36806 47888 36840
rect 47922 36806 47978 36840
rect 48012 36806 48068 36840
rect 48102 36806 48161 36840
rect 47467 36792 48161 36806
rect 47467 36758 47540 36792
rect 47574 36758 47640 36792
rect 47674 36758 47740 36792
rect 47774 36758 47840 36792
rect 47874 36758 47940 36792
rect 47974 36758 48040 36792
rect 48074 36758 48161 36792
rect 47467 36750 48161 36758
rect 47467 36716 47528 36750
rect 47562 36716 47618 36750
rect 47652 36716 47708 36750
rect 47742 36716 47798 36750
rect 47832 36716 47888 36750
rect 47922 36716 47978 36750
rect 48012 36716 48068 36750
rect 48102 36716 48161 36750
rect 47467 36692 48161 36716
rect 47467 36660 47540 36692
rect 47574 36660 47640 36692
rect 47674 36660 47740 36692
rect 47774 36660 47840 36692
rect 47467 36626 47528 36660
rect 47574 36658 47618 36660
rect 47674 36658 47708 36660
rect 47774 36658 47798 36660
rect 47562 36626 47618 36658
rect 47652 36626 47708 36658
rect 47742 36626 47798 36658
rect 47832 36658 47840 36660
rect 47874 36660 47940 36692
rect 47874 36658 47888 36660
rect 47832 36626 47888 36658
rect 47922 36658 47940 36660
rect 47974 36660 48040 36692
rect 48074 36660 48161 36692
rect 47974 36658 47978 36660
rect 47922 36626 47978 36658
rect 48012 36658 48040 36660
rect 48012 36626 48068 36658
rect 48102 36626 48161 36660
rect 47467 36592 48161 36626
rect 47467 36570 47540 36592
rect 47574 36570 47640 36592
rect 47674 36570 47740 36592
rect 47774 36570 47840 36592
rect 47467 36536 47528 36570
rect 47574 36558 47618 36570
rect 47674 36558 47708 36570
rect 47774 36558 47798 36570
rect 47562 36536 47618 36558
rect 47652 36536 47708 36558
rect 47742 36536 47798 36558
rect 47832 36558 47840 36570
rect 47874 36570 47940 36592
rect 47874 36558 47888 36570
rect 47832 36536 47888 36558
rect 47922 36558 47940 36570
rect 47974 36570 48040 36592
rect 48074 36570 48161 36592
rect 47974 36558 47978 36570
rect 47922 36536 47978 36558
rect 48012 36558 48040 36570
rect 48012 36536 48068 36558
rect 48102 36536 48161 36570
rect 47467 36492 48161 36536
rect 47467 36480 47540 36492
rect 47574 36480 47640 36492
rect 47674 36480 47740 36492
rect 47774 36480 47840 36492
rect 47467 36446 47528 36480
rect 47574 36458 47618 36480
rect 47674 36458 47708 36480
rect 47774 36458 47798 36480
rect 47562 36446 47618 36458
rect 47652 36446 47708 36458
rect 47742 36446 47798 36458
rect 47832 36458 47840 36480
rect 47874 36480 47940 36492
rect 47874 36458 47888 36480
rect 47832 36446 47888 36458
rect 47922 36458 47940 36480
rect 47974 36480 48040 36492
rect 48074 36480 48161 36492
rect 47974 36458 47978 36480
rect 47922 36446 47978 36458
rect 48012 36458 48040 36480
rect 48012 36446 48068 36458
rect 48102 36446 48161 36480
rect 47467 36385 48161 36446
rect 48223 37028 48295 37084
rect 48223 36994 48242 37028
rect 48276 36994 48295 37028
rect 48223 36938 48295 36994
rect 48223 36904 48242 36938
rect 48276 36904 48295 36938
rect 48223 36848 48295 36904
rect 48223 36814 48242 36848
rect 48276 36814 48295 36848
rect 48223 36758 48295 36814
rect 48223 36724 48242 36758
rect 48276 36724 48295 36758
rect 48223 36668 48295 36724
rect 48223 36634 48242 36668
rect 48276 36634 48295 36668
rect 48223 36578 48295 36634
rect 48223 36544 48242 36578
rect 48276 36544 48295 36578
rect 48223 36488 48295 36544
rect 48223 36454 48242 36488
rect 48276 36454 48295 36488
rect 48223 36398 48295 36454
rect 47333 36323 47405 36383
rect 48223 36364 48242 36398
rect 48276 36364 48295 36398
rect 48223 36323 48295 36364
rect 47333 36304 48295 36323
rect 47333 36270 47430 36304
rect 47464 36270 47520 36304
rect 47554 36270 47610 36304
rect 47644 36270 47700 36304
rect 47734 36270 47790 36304
rect 47824 36270 47880 36304
rect 47914 36270 47970 36304
rect 48004 36270 48060 36304
rect 48094 36270 48150 36304
rect 48184 36270 48295 36304
rect 47333 36251 48295 36270
rect 48359 37194 48391 37228
rect 48425 37194 48544 37228
rect 48578 37194 48609 37228
rect 49699 37228 49949 37277
rect 48359 37138 48609 37194
rect 48359 37104 48391 37138
rect 48425 37104 48544 37138
rect 48578 37104 48609 37138
rect 48359 37048 48609 37104
rect 48359 37014 48391 37048
rect 48425 37014 48544 37048
rect 48578 37014 48609 37048
rect 48359 36958 48609 37014
rect 48359 36924 48391 36958
rect 48425 36924 48544 36958
rect 48578 36924 48609 36958
rect 48359 36868 48609 36924
rect 48359 36834 48391 36868
rect 48425 36834 48544 36868
rect 48578 36834 48609 36868
rect 48359 36778 48609 36834
rect 48359 36744 48391 36778
rect 48425 36744 48544 36778
rect 48578 36744 48609 36778
rect 48359 36688 48609 36744
rect 48359 36654 48391 36688
rect 48425 36654 48544 36688
rect 48578 36654 48609 36688
rect 48359 36598 48609 36654
rect 48359 36564 48391 36598
rect 48425 36564 48544 36598
rect 48578 36564 48609 36598
rect 48359 36508 48609 36564
rect 48359 36474 48391 36508
rect 48425 36474 48544 36508
rect 48578 36474 48609 36508
rect 48359 36418 48609 36474
rect 48359 36384 48391 36418
rect 48425 36384 48544 36418
rect 48578 36384 48609 36418
rect 48359 36328 48609 36384
rect 48359 36294 48391 36328
rect 48425 36294 48544 36328
rect 48578 36294 48609 36328
rect 47019 36204 47051 36238
rect 47085 36204 47204 36238
rect 47238 36204 47269 36238
rect 47019 36187 47269 36204
rect 48359 36238 48609 36294
rect 48673 37196 49635 37213
rect 48673 37162 48694 37196
rect 48728 37162 48784 37196
rect 48818 37194 48874 37196
rect 48908 37194 48964 37196
rect 48998 37194 49054 37196
rect 49088 37194 49144 37196
rect 49178 37194 49234 37196
rect 49268 37194 49324 37196
rect 49358 37194 49414 37196
rect 49448 37194 49504 37196
rect 49538 37194 49594 37196
rect 48838 37162 48874 37194
rect 48928 37162 48964 37194
rect 49018 37162 49054 37194
rect 49108 37162 49144 37194
rect 49198 37162 49234 37194
rect 49288 37162 49324 37194
rect 49378 37162 49414 37194
rect 49468 37162 49504 37194
rect 49558 37162 49594 37194
rect 49628 37162 49635 37196
rect 48673 37160 48804 37162
rect 48838 37160 48894 37162
rect 48928 37160 48984 37162
rect 49018 37160 49074 37162
rect 49108 37160 49164 37162
rect 49198 37160 49254 37162
rect 49288 37160 49344 37162
rect 49378 37160 49434 37162
rect 49468 37160 49524 37162
rect 49558 37160 49635 37162
rect 48673 37141 49635 37160
rect 48673 37137 48745 37141
rect 48673 37103 48692 37137
rect 48726 37103 48745 37137
rect 48673 37047 48745 37103
rect 49563 37118 49635 37141
rect 49563 37084 49582 37118
rect 49616 37084 49635 37118
rect 48673 37013 48692 37047
rect 48726 37013 48745 37047
rect 48673 36957 48745 37013
rect 48673 36923 48692 36957
rect 48726 36923 48745 36957
rect 48673 36867 48745 36923
rect 48673 36833 48692 36867
rect 48726 36833 48745 36867
rect 48673 36777 48745 36833
rect 48673 36743 48692 36777
rect 48726 36743 48745 36777
rect 48673 36687 48745 36743
rect 48673 36653 48692 36687
rect 48726 36653 48745 36687
rect 48673 36597 48745 36653
rect 48673 36563 48692 36597
rect 48726 36563 48745 36597
rect 48673 36507 48745 36563
rect 48673 36473 48692 36507
rect 48726 36473 48745 36507
rect 48673 36417 48745 36473
rect 48673 36383 48692 36417
rect 48726 36383 48745 36417
rect 48807 37020 49501 37079
rect 48807 36986 48868 37020
rect 48902 36992 48958 37020
rect 48992 36992 49048 37020
rect 49082 36992 49138 37020
rect 48914 36986 48958 36992
rect 49014 36986 49048 36992
rect 49114 36986 49138 36992
rect 49172 36992 49228 37020
rect 49172 36986 49180 36992
rect 48807 36958 48880 36986
rect 48914 36958 48980 36986
rect 49014 36958 49080 36986
rect 49114 36958 49180 36986
rect 49214 36986 49228 36992
rect 49262 36992 49318 37020
rect 49262 36986 49280 36992
rect 49214 36958 49280 36986
rect 49314 36986 49318 36992
rect 49352 36992 49408 37020
rect 49352 36986 49380 36992
rect 49442 36986 49501 37020
rect 49314 36958 49380 36986
rect 49414 36958 49501 36986
rect 48807 36930 49501 36958
rect 48807 36896 48868 36930
rect 48902 36896 48958 36930
rect 48992 36896 49048 36930
rect 49082 36896 49138 36930
rect 49172 36896 49228 36930
rect 49262 36896 49318 36930
rect 49352 36896 49408 36930
rect 49442 36896 49501 36930
rect 48807 36892 49501 36896
rect 48807 36858 48880 36892
rect 48914 36858 48980 36892
rect 49014 36858 49080 36892
rect 49114 36858 49180 36892
rect 49214 36858 49280 36892
rect 49314 36858 49380 36892
rect 49414 36858 49501 36892
rect 48807 36840 49501 36858
rect 48807 36806 48868 36840
rect 48902 36806 48958 36840
rect 48992 36806 49048 36840
rect 49082 36806 49138 36840
rect 49172 36806 49228 36840
rect 49262 36806 49318 36840
rect 49352 36806 49408 36840
rect 49442 36806 49501 36840
rect 48807 36792 49501 36806
rect 48807 36758 48880 36792
rect 48914 36758 48980 36792
rect 49014 36758 49080 36792
rect 49114 36758 49180 36792
rect 49214 36758 49280 36792
rect 49314 36758 49380 36792
rect 49414 36758 49501 36792
rect 48807 36750 49501 36758
rect 48807 36716 48868 36750
rect 48902 36716 48958 36750
rect 48992 36716 49048 36750
rect 49082 36716 49138 36750
rect 49172 36716 49228 36750
rect 49262 36716 49318 36750
rect 49352 36716 49408 36750
rect 49442 36716 49501 36750
rect 48807 36692 49501 36716
rect 48807 36660 48880 36692
rect 48914 36660 48980 36692
rect 49014 36660 49080 36692
rect 49114 36660 49180 36692
rect 48807 36626 48868 36660
rect 48914 36658 48958 36660
rect 49014 36658 49048 36660
rect 49114 36658 49138 36660
rect 48902 36626 48958 36658
rect 48992 36626 49048 36658
rect 49082 36626 49138 36658
rect 49172 36658 49180 36660
rect 49214 36660 49280 36692
rect 49214 36658 49228 36660
rect 49172 36626 49228 36658
rect 49262 36658 49280 36660
rect 49314 36660 49380 36692
rect 49414 36660 49501 36692
rect 49314 36658 49318 36660
rect 49262 36626 49318 36658
rect 49352 36658 49380 36660
rect 49352 36626 49408 36658
rect 49442 36626 49501 36660
rect 48807 36592 49501 36626
rect 48807 36570 48880 36592
rect 48914 36570 48980 36592
rect 49014 36570 49080 36592
rect 49114 36570 49180 36592
rect 48807 36536 48868 36570
rect 48914 36558 48958 36570
rect 49014 36558 49048 36570
rect 49114 36558 49138 36570
rect 48902 36536 48958 36558
rect 48992 36536 49048 36558
rect 49082 36536 49138 36558
rect 49172 36558 49180 36570
rect 49214 36570 49280 36592
rect 49214 36558 49228 36570
rect 49172 36536 49228 36558
rect 49262 36558 49280 36570
rect 49314 36570 49380 36592
rect 49414 36570 49501 36592
rect 49314 36558 49318 36570
rect 49262 36536 49318 36558
rect 49352 36558 49380 36570
rect 49352 36536 49408 36558
rect 49442 36536 49501 36570
rect 48807 36492 49501 36536
rect 48807 36480 48880 36492
rect 48914 36480 48980 36492
rect 49014 36480 49080 36492
rect 49114 36480 49180 36492
rect 48807 36446 48868 36480
rect 48914 36458 48958 36480
rect 49014 36458 49048 36480
rect 49114 36458 49138 36480
rect 48902 36446 48958 36458
rect 48992 36446 49048 36458
rect 49082 36446 49138 36458
rect 49172 36458 49180 36480
rect 49214 36480 49280 36492
rect 49214 36458 49228 36480
rect 49172 36446 49228 36458
rect 49262 36458 49280 36480
rect 49314 36480 49380 36492
rect 49414 36480 49501 36492
rect 49314 36458 49318 36480
rect 49262 36446 49318 36458
rect 49352 36458 49380 36480
rect 49352 36446 49408 36458
rect 49442 36446 49501 36480
rect 48807 36385 49501 36446
rect 49563 37028 49635 37084
rect 49563 36994 49582 37028
rect 49616 36994 49635 37028
rect 49563 36938 49635 36994
rect 49563 36904 49582 36938
rect 49616 36904 49635 36938
rect 49563 36848 49635 36904
rect 49563 36814 49582 36848
rect 49616 36814 49635 36848
rect 49563 36758 49635 36814
rect 49563 36724 49582 36758
rect 49616 36724 49635 36758
rect 49563 36668 49635 36724
rect 49563 36634 49582 36668
rect 49616 36634 49635 36668
rect 49563 36578 49635 36634
rect 49563 36544 49582 36578
rect 49616 36544 49635 36578
rect 49563 36488 49635 36544
rect 49563 36454 49582 36488
rect 49616 36454 49635 36488
rect 49563 36398 49635 36454
rect 48673 36323 48745 36383
rect 49563 36364 49582 36398
rect 49616 36364 49635 36398
rect 49563 36323 49635 36364
rect 48673 36304 49635 36323
rect 48673 36270 48770 36304
rect 48804 36270 48860 36304
rect 48894 36270 48950 36304
rect 48984 36270 49040 36304
rect 49074 36270 49130 36304
rect 49164 36270 49220 36304
rect 49254 36270 49310 36304
rect 49344 36270 49400 36304
rect 49434 36270 49490 36304
rect 49524 36270 49635 36304
rect 48673 36251 49635 36270
rect 49699 37194 49731 37228
rect 49765 37194 49884 37228
rect 49918 37194 49949 37228
rect 51039 37228 51289 37277
rect 49699 37138 49949 37194
rect 49699 37104 49731 37138
rect 49765 37104 49884 37138
rect 49918 37104 49949 37138
rect 49699 37048 49949 37104
rect 49699 37014 49731 37048
rect 49765 37014 49884 37048
rect 49918 37014 49949 37048
rect 49699 36958 49949 37014
rect 49699 36924 49731 36958
rect 49765 36924 49884 36958
rect 49918 36924 49949 36958
rect 49699 36868 49949 36924
rect 49699 36834 49731 36868
rect 49765 36834 49884 36868
rect 49918 36834 49949 36868
rect 49699 36778 49949 36834
rect 49699 36744 49731 36778
rect 49765 36744 49884 36778
rect 49918 36744 49949 36778
rect 49699 36688 49949 36744
rect 49699 36654 49731 36688
rect 49765 36654 49884 36688
rect 49918 36654 49949 36688
rect 49699 36598 49949 36654
rect 49699 36564 49731 36598
rect 49765 36564 49884 36598
rect 49918 36564 49949 36598
rect 49699 36508 49949 36564
rect 49699 36474 49731 36508
rect 49765 36474 49884 36508
rect 49918 36474 49949 36508
rect 49699 36418 49949 36474
rect 49699 36384 49731 36418
rect 49765 36384 49884 36418
rect 49918 36384 49949 36418
rect 49699 36328 49949 36384
rect 49699 36294 49731 36328
rect 49765 36294 49884 36328
rect 49918 36294 49949 36328
rect 48359 36204 48391 36238
rect 48425 36204 48544 36238
rect 48578 36204 48609 36238
rect 48359 36187 48609 36204
rect 49699 36238 49949 36294
rect 50013 37196 50975 37213
rect 50013 37162 50034 37196
rect 50068 37162 50124 37196
rect 50158 37194 50214 37196
rect 50248 37194 50304 37196
rect 50338 37194 50394 37196
rect 50428 37194 50484 37196
rect 50518 37194 50574 37196
rect 50608 37194 50664 37196
rect 50698 37194 50754 37196
rect 50788 37194 50844 37196
rect 50878 37194 50934 37196
rect 50178 37162 50214 37194
rect 50268 37162 50304 37194
rect 50358 37162 50394 37194
rect 50448 37162 50484 37194
rect 50538 37162 50574 37194
rect 50628 37162 50664 37194
rect 50718 37162 50754 37194
rect 50808 37162 50844 37194
rect 50898 37162 50934 37194
rect 50968 37162 50975 37196
rect 50013 37160 50144 37162
rect 50178 37160 50234 37162
rect 50268 37160 50324 37162
rect 50358 37160 50414 37162
rect 50448 37160 50504 37162
rect 50538 37160 50594 37162
rect 50628 37160 50684 37162
rect 50718 37160 50774 37162
rect 50808 37160 50864 37162
rect 50898 37160 50975 37162
rect 50013 37141 50975 37160
rect 50013 37137 50085 37141
rect 50013 37103 50032 37137
rect 50066 37103 50085 37137
rect 50013 37047 50085 37103
rect 50903 37118 50975 37141
rect 50903 37084 50922 37118
rect 50956 37084 50975 37118
rect 50013 37013 50032 37047
rect 50066 37013 50085 37047
rect 50013 36957 50085 37013
rect 50013 36923 50032 36957
rect 50066 36923 50085 36957
rect 50013 36867 50085 36923
rect 50013 36833 50032 36867
rect 50066 36833 50085 36867
rect 50013 36777 50085 36833
rect 50013 36743 50032 36777
rect 50066 36743 50085 36777
rect 50013 36687 50085 36743
rect 50013 36653 50032 36687
rect 50066 36653 50085 36687
rect 50013 36597 50085 36653
rect 50013 36563 50032 36597
rect 50066 36563 50085 36597
rect 50013 36507 50085 36563
rect 50013 36473 50032 36507
rect 50066 36473 50085 36507
rect 50013 36417 50085 36473
rect 50013 36383 50032 36417
rect 50066 36383 50085 36417
rect 50147 37020 50841 37079
rect 50147 36986 50208 37020
rect 50242 36992 50298 37020
rect 50332 36992 50388 37020
rect 50422 36992 50478 37020
rect 50254 36986 50298 36992
rect 50354 36986 50388 36992
rect 50454 36986 50478 36992
rect 50512 36992 50568 37020
rect 50512 36986 50520 36992
rect 50147 36958 50220 36986
rect 50254 36958 50320 36986
rect 50354 36958 50420 36986
rect 50454 36958 50520 36986
rect 50554 36986 50568 36992
rect 50602 36992 50658 37020
rect 50602 36986 50620 36992
rect 50554 36958 50620 36986
rect 50654 36986 50658 36992
rect 50692 36992 50748 37020
rect 50692 36986 50720 36992
rect 50782 36986 50841 37020
rect 50654 36958 50720 36986
rect 50754 36958 50841 36986
rect 50147 36930 50841 36958
rect 50147 36896 50208 36930
rect 50242 36896 50298 36930
rect 50332 36896 50388 36930
rect 50422 36896 50478 36930
rect 50512 36896 50568 36930
rect 50602 36896 50658 36930
rect 50692 36896 50748 36930
rect 50782 36896 50841 36930
rect 50147 36892 50841 36896
rect 50147 36858 50220 36892
rect 50254 36858 50320 36892
rect 50354 36858 50420 36892
rect 50454 36858 50520 36892
rect 50554 36858 50620 36892
rect 50654 36858 50720 36892
rect 50754 36858 50841 36892
rect 50147 36840 50841 36858
rect 50147 36806 50208 36840
rect 50242 36806 50298 36840
rect 50332 36806 50388 36840
rect 50422 36806 50478 36840
rect 50512 36806 50568 36840
rect 50602 36806 50658 36840
rect 50692 36806 50748 36840
rect 50782 36806 50841 36840
rect 50147 36792 50841 36806
rect 50147 36758 50220 36792
rect 50254 36758 50320 36792
rect 50354 36758 50420 36792
rect 50454 36758 50520 36792
rect 50554 36758 50620 36792
rect 50654 36758 50720 36792
rect 50754 36758 50841 36792
rect 50147 36750 50841 36758
rect 50147 36716 50208 36750
rect 50242 36716 50298 36750
rect 50332 36716 50388 36750
rect 50422 36716 50478 36750
rect 50512 36716 50568 36750
rect 50602 36716 50658 36750
rect 50692 36716 50748 36750
rect 50782 36716 50841 36750
rect 50147 36692 50841 36716
rect 50147 36660 50220 36692
rect 50254 36660 50320 36692
rect 50354 36660 50420 36692
rect 50454 36660 50520 36692
rect 50147 36626 50208 36660
rect 50254 36658 50298 36660
rect 50354 36658 50388 36660
rect 50454 36658 50478 36660
rect 50242 36626 50298 36658
rect 50332 36626 50388 36658
rect 50422 36626 50478 36658
rect 50512 36658 50520 36660
rect 50554 36660 50620 36692
rect 50554 36658 50568 36660
rect 50512 36626 50568 36658
rect 50602 36658 50620 36660
rect 50654 36660 50720 36692
rect 50754 36660 50841 36692
rect 50654 36658 50658 36660
rect 50602 36626 50658 36658
rect 50692 36658 50720 36660
rect 50692 36626 50748 36658
rect 50782 36626 50841 36660
rect 50147 36592 50841 36626
rect 50147 36570 50220 36592
rect 50254 36570 50320 36592
rect 50354 36570 50420 36592
rect 50454 36570 50520 36592
rect 50147 36536 50208 36570
rect 50254 36558 50298 36570
rect 50354 36558 50388 36570
rect 50454 36558 50478 36570
rect 50242 36536 50298 36558
rect 50332 36536 50388 36558
rect 50422 36536 50478 36558
rect 50512 36558 50520 36570
rect 50554 36570 50620 36592
rect 50554 36558 50568 36570
rect 50512 36536 50568 36558
rect 50602 36558 50620 36570
rect 50654 36570 50720 36592
rect 50754 36570 50841 36592
rect 50654 36558 50658 36570
rect 50602 36536 50658 36558
rect 50692 36558 50720 36570
rect 50692 36536 50748 36558
rect 50782 36536 50841 36570
rect 50147 36492 50841 36536
rect 50147 36480 50220 36492
rect 50254 36480 50320 36492
rect 50354 36480 50420 36492
rect 50454 36480 50520 36492
rect 50147 36446 50208 36480
rect 50254 36458 50298 36480
rect 50354 36458 50388 36480
rect 50454 36458 50478 36480
rect 50242 36446 50298 36458
rect 50332 36446 50388 36458
rect 50422 36446 50478 36458
rect 50512 36458 50520 36480
rect 50554 36480 50620 36492
rect 50554 36458 50568 36480
rect 50512 36446 50568 36458
rect 50602 36458 50620 36480
rect 50654 36480 50720 36492
rect 50754 36480 50841 36492
rect 50654 36458 50658 36480
rect 50602 36446 50658 36458
rect 50692 36458 50720 36480
rect 50692 36446 50748 36458
rect 50782 36446 50841 36480
rect 50147 36385 50841 36446
rect 50903 37028 50975 37084
rect 50903 36994 50922 37028
rect 50956 36994 50975 37028
rect 50903 36938 50975 36994
rect 50903 36904 50922 36938
rect 50956 36904 50975 36938
rect 50903 36848 50975 36904
rect 50903 36814 50922 36848
rect 50956 36814 50975 36848
rect 50903 36758 50975 36814
rect 50903 36724 50922 36758
rect 50956 36724 50975 36758
rect 50903 36668 50975 36724
rect 50903 36634 50922 36668
rect 50956 36634 50975 36668
rect 50903 36578 50975 36634
rect 50903 36544 50922 36578
rect 50956 36544 50975 36578
rect 50903 36488 50975 36544
rect 50903 36454 50922 36488
rect 50956 36454 50975 36488
rect 50903 36398 50975 36454
rect 50013 36323 50085 36383
rect 50903 36364 50922 36398
rect 50956 36364 50975 36398
rect 50903 36323 50975 36364
rect 50013 36304 50975 36323
rect 50013 36270 50110 36304
rect 50144 36270 50200 36304
rect 50234 36270 50290 36304
rect 50324 36270 50380 36304
rect 50414 36270 50470 36304
rect 50504 36270 50560 36304
rect 50594 36270 50650 36304
rect 50684 36270 50740 36304
rect 50774 36270 50830 36304
rect 50864 36270 50975 36304
rect 50013 36251 50975 36270
rect 51039 37194 51071 37228
rect 51105 37194 51224 37228
rect 51258 37194 51289 37228
rect 52379 37228 52478 37277
rect 51039 37138 51289 37194
rect 51039 37104 51071 37138
rect 51105 37104 51224 37138
rect 51258 37104 51289 37138
rect 51039 37048 51289 37104
rect 51039 37014 51071 37048
rect 51105 37014 51224 37048
rect 51258 37014 51289 37048
rect 51039 36958 51289 37014
rect 51039 36924 51071 36958
rect 51105 36924 51224 36958
rect 51258 36924 51289 36958
rect 51039 36868 51289 36924
rect 51039 36834 51071 36868
rect 51105 36834 51224 36868
rect 51258 36834 51289 36868
rect 51039 36778 51289 36834
rect 51039 36744 51071 36778
rect 51105 36744 51224 36778
rect 51258 36744 51289 36778
rect 51039 36688 51289 36744
rect 51039 36654 51071 36688
rect 51105 36654 51224 36688
rect 51258 36654 51289 36688
rect 51039 36598 51289 36654
rect 51039 36564 51071 36598
rect 51105 36564 51224 36598
rect 51258 36564 51289 36598
rect 51039 36508 51289 36564
rect 51039 36474 51071 36508
rect 51105 36474 51224 36508
rect 51258 36474 51289 36508
rect 51039 36418 51289 36474
rect 51039 36384 51071 36418
rect 51105 36384 51224 36418
rect 51258 36384 51289 36418
rect 51039 36328 51289 36384
rect 51039 36294 51071 36328
rect 51105 36294 51224 36328
rect 51258 36294 51289 36328
rect 49699 36204 49731 36238
rect 49765 36204 49884 36238
rect 49918 36204 49949 36238
rect 49699 36187 49949 36204
rect 51039 36238 51289 36294
rect 51353 37196 52315 37213
rect 51353 37162 51374 37196
rect 51408 37162 51464 37196
rect 51498 37194 51554 37196
rect 51588 37194 51644 37196
rect 51678 37194 51734 37196
rect 51768 37194 51824 37196
rect 51858 37194 51914 37196
rect 51948 37194 52004 37196
rect 52038 37194 52094 37196
rect 52128 37194 52184 37196
rect 52218 37194 52274 37196
rect 51518 37162 51554 37194
rect 51608 37162 51644 37194
rect 51698 37162 51734 37194
rect 51788 37162 51824 37194
rect 51878 37162 51914 37194
rect 51968 37162 52004 37194
rect 52058 37162 52094 37194
rect 52148 37162 52184 37194
rect 52238 37162 52274 37194
rect 52308 37162 52315 37196
rect 51353 37160 51484 37162
rect 51518 37160 51574 37162
rect 51608 37160 51664 37162
rect 51698 37160 51754 37162
rect 51788 37160 51844 37162
rect 51878 37160 51934 37162
rect 51968 37160 52024 37162
rect 52058 37160 52114 37162
rect 52148 37160 52204 37162
rect 52238 37160 52315 37162
rect 51353 37141 52315 37160
rect 51353 37137 51425 37141
rect 51353 37103 51372 37137
rect 51406 37103 51425 37137
rect 51353 37047 51425 37103
rect 52243 37118 52315 37141
rect 52243 37084 52262 37118
rect 52296 37084 52315 37118
rect 51353 37013 51372 37047
rect 51406 37013 51425 37047
rect 51353 36957 51425 37013
rect 51353 36923 51372 36957
rect 51406 36923 51425 36957
rect 51353 36867 51425 36923
rect 51353 36833 51372 36867
rect 51406 36833 51425 36867
rect 51353 36777 51425 36833
rect 51353 36743 51372 36777
rect 51406 36743 51425 36777
rect 51353 36687 51425 36743
rect 51353 36653 51372 36687
rect 51406 36653 51425 36687
rect 51353 36597 51425 36653
rect 51353 36563 51372 36597
rect 51406 36563 51425 36597
rect 51353 36507 51425 36563
rect 51353 36473 51372 36507
rect 51406 36473 51425 36507
rect 51353 36417 51425 36473
rect 51353 36383 51372 36417
rect 51406 36383 51425 36417
rect 51487 37020 52181 37079
rect 51487 36986 51548 37020
rect 51582 36992 51638 37020
rect 51672 36992 51728 37020
rect 51762 36992 51818 37020
rect 51594 36986 51638 36992
rect 51694 36986 51728 36992
rect 51794 36986 51818 36992
rect 51852 36992 51908 37020
rect 51852 36986 51860 36992
rect 51487 36958 51560 36986
rect 51594 36958 51660 36986
rect 51694 36958 51760 36986
rect 51794 36958 51860 36986
rect 51894 36986 51908 36992
rect 51942 36992 51998 37020
rect 51942 36986 51960 36992
rect 51894 36958 51960 36986
rect 51994 36986 51998 36992
rect 52032 36992 52088 37020
rect 52032 36986 52060 36992
rect 52122 36986 52181 37020
rect 51994 36958 52060 36986
rect 52094 36958 52181 36986
rect 51487 36930 52181 36958
rect 51487 36896 51548 36930
rect 51582 36896 51638 36930
rect 51672 36896 51728 36930
rect 51762 36896 51818 36930
rect 51852 36896 51908 36930
rect 51942 36896 51998 36930
rect 52032 36896 52088 36930
rect 52122 36896 52181 36930
rect 51487 36892 52181 36896
rect 51487 36858 51560 36892
rect 51594 36858 51660 36892
rect 51694 36858 51760 36892
rect 51794 36858 51860 36892
rect 51894 36858 51960 36892
rect 51994 36858 52060 36892
rect 52094 36858 52181 36892
rect 51487 36840 52181 36858
rect 51487 36806 51548 36840
rect 51582 36806 51638 36840
rect 51672 36806 51728 36840
rect 51762 36806 51818 36840
rect 51852 36806 51908 36840
rect 51942 36806 51998 36840
rect 52032 36806 52088 36840
rect 52122 36806 52181 36840
rect 51487 36792 52181 36806
rect 51487 36758 51560 36792
rect 51594 36758 51660 36792
rect 51694 36758 51760 36792
rect 51794 36758 51860 36792
rect 51894 36758 51960 36792
rect 51994 36758 52060 36792
rect 52094 36758 52181 36792
rect 51487 36750 52181 36758
rect 51487 36716 51548 36750
rect 51582 36716 51638 36750
rect 51672 36716 51728 36750
rect 51762 36716 51818 36750
rect 51852 36716 51908 36750
rect 51942 36716 51998 36750
rect 52032 36716 52088 36750
rect 52122 36716 52181 36750
rect 51487 36692 52181 36716
rect 51487 36660 51560 36692
rect 51594 36660 51660 36692
rect 51694 36660 51760 36692
rect 51794 36660 51860 36692
rect 51487 36626 51548 36660
rect 51594 36658 51638 36660
rect 51694 36658 51728 36660
rect 51794 36658 51818 36660
rect 51582 36626 51638 36658
rect 51672 36626 51728 36658
rect 51762 36626 51818 36658
rect 51852 36658 51860 36660
rect 51894 36660 51960 36692
rect 51894 36658 51908 36660
rect 51852 36626 51908 36658
rect 51942 36658 51960 36660
rect 51994 36660 52060 36692
rect 52094 36660 52181 36692
rect 51994 36658 51998 36660
rect 51942 36626 51998 36658
rect 52032 36658 52060 36660
rect 52032 36626 52088 36658
rect 52122 36626 52181 36660
rect 51487 36592 52181 36626
rect 51487 36570 51560 36592
rect 51594 36570 51660 36592
rect 51694 36570 51760 36592
rect 51794 36570 51860 36592
rect 51487 36536 51548 36570
rect 51594 36558 51638 36570
rect 51694 36558 51728 36570
rect 51794 36558 51818 36570
rect 51582 36536 51638 36558
rect 51672 36536 51728 36558
rect 51762 36536 51818 36558
rect 51852 36558 51860 36570
rect 51894 36570 51960 36592
rect 51894 36558 51908 36570
rect 51852 36536 51908 36558
rect 51942 36558 51960 36570
rect 51994 36570 52060 36592
rect 52094 36570 52181 36592
rect 51994 36558 51998 36570
rect 51942 36536 51998 36558
rect 52032 36558 52060 36570
rect 52032 36536 52088 36558
rect 52122 36536 52181 36570
rect 51487 36492 52181 36536
rect 51487 36480 51560 36492
rect 51594 36480 51660 36492
rect 51694 36480 51760 36492
rect 51794 36480 51860 36492
rect 51487 36446 51548 36480
rect 51594 36458 51638 36480
rect 51694 36458 51728 36480
rect 51794 36458 51818 36480
rect 51582 36446 51638 36458
rect 51672 36446 51728 36458
rect 51762 36446 51818 36458
rect 51852 36458 51860 36480
rect 51894 36480 51960 36492
rect 51894 36458 51908 36480
rect 51852 36446 51908 36458
rect 51942 36458 51960 36480
rect 51994 36480 52060 36492
rect 52094 36480 52181 36492
rect 51994 36458 51998 36480
rect 51942 36446 51998 36458
rect 52032 36458 52060 36480
rect 52032 36446 52088 36458
rect 52122 36446 52181 36480
rect 51487 36385 52181 36446
rect 52243 37028 52315 37084
rect 52243 36994 52262 37028
rect 52296 36994 52315 37028
rect 52243 36938 52315 36994
rect 52243 36904 52262 36938
rect 52296 36904 52315 36938
rect 52243 36848 52315 36904
rect 52243 36814 52262 36848
rect 52296 36814 52315 36848
rect 52243 36758 52315 36814
rect 52243 36724 52262 36758
rect 52296 36724 52315 36758
rect 52243 36668 52315 36724
rect 52243 36634 52262 36668
rect 52296 36634 52315 36668
rect 52243 36578 52315 36634
rect 52243 36544 52262 36578
rect 52296 36544 52315 36578
rect 52243 36488 52315 36544
rect 52243 36454 52262 36488
rect 52296 36454 52315 36488
rect 52243 36398 52315 36454
rect 51353 36323 51425 36383
rect 52243 36364 52262 36398
rect 52296 36364 52315 36398
rect 52243 36323 52315 36364
rect 51353 36304 52315 36323
rect 51353 36270 51450 36304
rect 51484 36270 51540 36304
rect 51574 36270 51630 36304
rect 51664 36270 51720 36304
rect 51754 36270 51810 36304
rect 51844 36270 51900 36304
rect 51934 36270 51990 36304
rect 52024 36270 52080 36304
rect 52114 36270 52170 36304
rect 52204 36270 52315 36304
rect 51353 36251 52315 36270
rect 52379 37194 52411 37228
rect 52445 37194 52478 37228
rect 52379 37138 52478 37194
rect 52379 37104 52411 37138
rect 52445 37104 52478 37138
rect 52379 37048 52478 37104
rect 52379 37014 52411 37048
rect 52445 37014 52478 37048
rect 52379 36958 52478 37014
rect 52379 36924 52411 36958
rect 52445 36924 52478 36958
rect 52379 36868 52478 36924
rect 52379 36834 52411 36868
rect 52445 36834 52478 36868
rect 52379 36778 52478 36834
rect 52379 36744 52411 36778
rect 52445 36744 52478 36778
rect 52379 36688 52478 36744
rect 52379 36654 52411 36688
rect 52445 36654 52478 36688
rect 52379 36598 52478 36654
rect 52379 36564 52411 36598
rect 52445 36564 52478 36598
rect 52379 36508 52478 36564
rect 52379 36474 52411 36508
rect 52445 36474 52478 36508
rect 52379 36418 52478 36474
rect 52379 36384 52411 36418
rect 52445 36384 52478 36418
rect 52379 36328 52478 36384
rect 52379 36294 52411 36328
rect 52445 36294 52478 36328
rect 51039 36204 51071 36238
rect 51105 36204 51224 36238
rect 51258 36204 51289 36238
rect 51039 36187 51289 36204
rect 52379 36238 52478 36294
rect 52379 36204 52411 36238
rect 52445 36204 52478 36238
rect 52379 36187 52478 36204
rect 41810 36154 52478 36187
rect 41810 36120 41940 36154
rect 41974 36120 42030 36154
rect 42064 36120 42120 36154
rect 42154 36120 42210 36154
rect 42244 36120 42300 36154
rect 42334 36120 42390 36154
rect 42424 36120 42480 36154
rect 42514 36120 42570 36154
rect 42604 36120 42660 36154
rect 42694 36120 42750 36154
rect 42784 36120 42840 36154
rect 42874 36120 42930 36154
rect 42964 36120 43280 36154
rect 43314 36120 43370 36154
rect 43404 36120 43460 36154
rect 43494 36120 43550 36154
rect 43584 36120 43640 36154
rect 43674 36120 43730 36154
rect 43764 36120 43820 36154
rect 43854 36120 43910 36154
rect 43944 36120 44000 36154
rect 44034 36120 44090 36154
rect 44124 36120 44180 36154
rect 44214 36120 44270 36154
rect 44304 36120 44620 36154
rect 44654 36120 44710 36154
rect 44744 36120 44800 36154
rect 44834 36120 44890 36154
rect 44924 36120 44980 36154
rect 45014 36120 45070 36154
rect 45104 36120 45160 36154
rect 45194 36120 45250 36154
rect 45284 36120 45340 36154
rect 45374 36120 45430 36154
rect 45464 36120 45520 36154
rect 45554 36120 45610 36154
rect 45644 36120 45960 36154
rect 45994 36120 46050 36154
rect 46084 36120 46140 36154
rect 46174 36120 46230 36154
rect 46264 36120 46320 36154
rect 46354 36120 46410 36154
rect 46444 36120 46500 36154
rect 46534 36120 46590 36154
rect 46624 36120 46680 36154
rect 46714 36120 46770 36154
rect 46804 36120 46860 36154
rect 46894 36120 46950 36154
rect 46984 36120 47300 36154
rect 47334 36120 47390 36154
rect 47424 36120 47480 36154
rect 47514 36120 47570 36154
rect 47604 36120 47660 36154
rect 47694 36120 47750 36154
rect 47784 36120 47840 36154
rect 47874 36120 47930 36154
rect 47964 36120 48020 36154
rect 48054 36120 48110 36154
rect 48144 36120 48200 36154
rect 48234 36120 48290 36154
rect 48324 36120 48640 36154
rect 48674 36120 48730 36154
rect 48764 36120 48820 36154
rect 48854 36120 48910 36154
rect 48944 36120 49000 36154
rect 49034 36120 49090 36154
rect 49124 36120 49180 36154
rect 49214 36120 49270 36154
rect 49304 36120 49360 36154
rect 49394 36120 49450 36154
rect 49484 36120 49540 36154
rect 49574 36120 49630 36154
rect 49664 36120 49980 36154
rect 50014 36120 50070 36154
rect 50104 36120 50160 36154
rect 50194 36120 50250 36154
rect 50284 36120 50340 36154
rect 50374 36120 50430 36154
rect 50464 36120 50520 36154
rect 50554 36120 50610 36154
rect 50644 36120 50700 36154
rect 50734 36120 50790 36154
rect 50824 36120 50880 36154
rect 50914 36120 50970 36154
rect 51004 36120 51320 36154
rect 51354 36120 51410 36154
rect 51444 36120 51500 36154
rect 51534 36120 51590 36154
rect 51624 36120 51680 36154
rect 51714 36120 51770 36154
rect 51804 36120 51860 36154
rect 51894 36120 51950 36154
rect 51984 36120 52040 36154
rect 52074 36120 52130 36154
rect 52164 36120 52220 36154
rect 52254 36120 52310 36154
rect 52344 36120 52478 36154
rect 41810 36088 52478 36120
rect 37472 36057 40348 36062
rect 25348 35949 25408 36032
rect 37472 36023 37565 36057
rect 37599 36023 40348 36057
rect 37472 36002 40348 36023
rect 25348 35915 25361 35949
rect 25395 35915 25408 35949
rect 37472 35955 40348 35956
rect 37472 35943 38577 35955
rect 25348 35822 25408 35915
rect 26398 35919 26558 35942
rect 26398 35885 26463 35919
rect 26497 35885 26558 35919
rect 26398 35822 26558 35885
rect 27698 35919 27858 35942
rect 27698 35885 27763 35919
rect 27797 35885 27858 35919
rect 37472 35909 37655 35943
rect 37689 35909 38055 35943
rect 38089 35909 38455 35943
rect 38489 35921 38577 35943
rect 38611 35943 40348 35955
rect 38611 35921 38855 35943
rect 38489 35909 38855 35921
rect 38889 35909 39255 35943
rect 39289 35909 39655 35943
rect 39689 35909 40055 35943
rect 40089 35909 40348 35943
rect 37472 35896 40348 35909
rect 27698 35822 27858 35885
rect 11992 35809 13332 35822
rect 11992 35775 12175 35809
rect 12209 35775 12375 35809
rect 12409 35775 12575 35809
rect 12609 35775 12775 35809
rect 12809 35775 12975 35809
rect 13009 35775 13175 35809
rect 13209 35775 13332 35809
rect 11992 35762 13332 35775
rect 13678 35809 16118 35822
rect 13678 35775 13861 35809
rect 13895 35775 14061 35809
rect 14095 35775 14261 35809
rect 14295 35775 14461 35809
rect 14495 35775 14661 35809
rect 14695 35775 14861 35809
rect 14895 35775 15061 35809
rect 15095 35775 15261 35809
rect 15295 35775 15461 35809
rect 15495 35775 15661 35809
rect 15695 35775 15861 35809
rect 15895 35775 16118 35809
rect 13678 35762 16118 35775
rect 16422 35809 18862 35822
rect 16422 35775 16605 35809
rect 16639 35775 16805 35809
rect 16839 35775 17005 35809
rect 17039 35775 17205 35809
rect 17239 35775 17405 35809
rect 17439 35775 17605 35809
rect 17639 35775 17805 35809
rect 17839 35775 18005 35809
rect 18039 35775 18205 35809
rect 18239 35775 18405 35809
rect 18439 35775 18605 35809
rect 18639 35775 18862 35809
rect 16422 35762 18862 35775
rect 19168 35809 22180 35822
rect 19168 35775 19351 35809
rect 19385 35775 19551 35809
rect 19585 35775 19751 35809
rect 19785 35775 19951 35809
rect 19985 35775 20151 35809
rect 20185 35775 20351 35809
rect 20385 35775 20551 35809
rect 20585 35775 20751 35809
rect 20785 35775 20951 35809
rect 20985 35775 21151 35809
rect 21185 35775 21351 35809
rect 21385 35775 21551 35809
rect 21585 35775 21751 35809
rect 21785 35775 21951 35809
rect 21985 35775 22180 35809
rect 19168 35762 22180 35775
rect 22498 35809 24938 35822
rect 22498 35775 22681 35809
rect 22715 35775 22881 35809
rect 22915 35775 23081 35809
rect 23115 35775 23281 35809
rect 23315 35775 23481 35809
rect 23515 35775 23681 35809
rect 23715 35775 23881 35809
rect 23915 35775 24081 35809
rect 24115 35775 24281 35809
rect 24315 35775 24481 35809
rect 24515 35775 24681 35809
rect 24715 35775 24938 35809
rect 22498 35762 24938 35775
rect 25320 35809 29598 35822
rect 25320 35775 25601 35809
rect 25635 35775 26001 35809
rect 26035 35775 26401 35809
rect 26435 35775 26801 35809
rect 26835 35775 27201 35809
rect 27235 35775 27601 35809
rect 27635 35775 28001 35809
rect 28035 35775 28401 35809
rect 28435 35775 28801 35809
rect 28835 35775 29201 35809
rect 29235 35775 29598 35809
rect 25320 35762 29598 35775
rect 29928 35809 37096 35822
rect 29928 35775 30111 35809
rect 30145 35775 30511 35809
rect 30545 35775 30911 35809
rect 30945 35775 31311 35809
rect 31345 35775 31711 35809
rect 31745 35775 32111 35809
rect 32145 35775 32511 35809
rect 32545 35775 32911 35809
rect 32945 35775 33311 35809
rect 33345 35775 33711 35809
rect 33745 35775 34111 35809
rect 34145 35775 34511 35809
rect 34545 35775 34911 35809
rect 34945 35775 35311 35809
rect 35345 35775 35711 35809
rect 35745 35775 36111 35809
rect 36145 35775 36511 35809
rect 36545 35775 36911 35809
rect 36945 35775 37096 35809
rect 29928 35762 37096 35775
rect 37374 35809 40348 35822
rect 37374 35775 37655 35809
rect 37689 35775 38055 35809
rect 38089 35775 38455 35809
rect 38489 35775 38855 35809
rect 38889 35775 39255 35809
rect 39289 35775 39655 35809
rect 39689 35775 40055 35809
rect 40089 35775 40348 35809
rect 37374 35762 40348 35775
rect 41784 35809 52504 35822
rect 41784 35775 41967 35809
rect 42001 35775 42167 35809
rect 42201 35775 42367 35809
rect 42401 35775 42567 35809
rect 42601 35775 42767 35809
rect 42801 35775 42967 35809
rect 43001 35775 43167 35809
rect 43201 35775 43367 35809
rect 43401 35775 43567 35809
rect 43601 35775 43767 35809
rect 43801 35775 43967 35809
rect 44001 35775 44167 35809
rect 44201 35775 44367 35809
rect 44401 35775 44567 35809
rect 44601 35775 44767 35809
rect 44801 35775 44967 35809
rect 45001 35775 45167 35809
rect 45201 35775 45367 35809
rect 45401 35775 45567 35809
rect 45601 35775 45767 35809
rect 45801 35775 45967 35809
rect 46001 35775 46167 35809
rect 46201 35775 46367 35809
rect 46401 35775 46567 35809
rect 46601 35775 46767 35809
rect 46801 35775 46967 35809
rect 47001 35775 47167 35809
rect 47201 35775 47367 35809
rect 47401 35775 47567 35809
rect 47601 35775 47767 35809
rect 47801 35775 47967 35809
rect 48001 35775 48167 35809
rect 48201 35775 48367 35809
rect 48401 35775 48567 35809
rect 48601 35775 48767 35809
rect 48801 35775 48967 35809
rect 49001 35775 49167 35809
rect 49201 35775 49367 35809
rect 49401 35775 49567 35809
rect 49601 35775 49767 35809
rect 49801 35775 49967 35809
rect 50001 35775 50167 35809
rect 50201 35775 50367 35809
rect 50401 35775 50567 35809
rect 50601 35775 50767 35809
rect 50801 35775 50967 35809
rect 51001 35775 51167 35809
rect 51201 35775 51367 35809
rect 51401 35775 51567 35809
rect 51601 35775 51767 35809
rect 51801 35775 51967 35809
rect 52001 35775 52167 35809
rect 52201 35775 52367 35809
rect 52401 35775 52504 35809
rect 41784 35762 52504 35775
rect 19264 33929 21704 33942
rect 19264 33895 19447 33929
rect 19481 33895 19647 33929
rect 19681 33895 19847 33929
rect 19881 33895 20047 33929
rect 20081 33895 20247 33929
rect 20281 33895 20447 33929
rect 20481 33895 20647 33929
rect 20681 33895 20847 33929
rect 20881 33895 21047 33929
rect 21081 33895 21247 33929
rect 21281 33895 21447 33929
rect 21481 33895 21704 33929
rect 19264 33882 21704 33895
rect 22010 33929 25022 33942
rect 22010 33895 22193 33929
rect 22227 33895 22393 33929
rect 22427 33895 22593 33929
rect 22627 33895 22793 33929
rect 22827 33895 22993 33929
rect 23027 33895 23193 33929
rect 23227 33895 23393 33929
rect 23427 33895 23593 33929
rect 23627 33895 23793 33929
rect 23827 33895 23993 33929
rect 24027 33895 24193 33929
rect 24227 33895 24393 33929
rect 24427 33895 24593 33929
rect 24627 33895 24793 33929
rect 24827 33895 25022 33929
rect 22010 33882 25022 33895
rect 26204 33929 33372 33942
rect 26204 33895 26387 33929
rect 26421 33895 26787 33929
rect 26821 33895 27187 33929
rect 27221 33895 27587 33929
rect 27621 33895 27987 33929
rect 28021 33895 28387 33929
rect 28421 33895 28787 33929
rect 28821 33895 29187 33929
rect 29221 33895 29587 33929
rect 29621 33895 29987 33929
rect 30021 33895 30387 33929
rect 30421 33895 30787 33929
rect 30821 33895 31187 33929
rect 31221 33895 31587 33929
rect 31621 33895 31987 33929
rect 32021 33895 32387 33929
rect 32421 33895 32787 33929
rect 32821 33895 33187 33929
rect 33221 33895 33372 33929
rect 26204 33882 33372 33895
rect 33652 33929 40820 33942
rect 33652 33895 33835 33929
rect 33869 33895 34235 33929
rect 34269 33895 34635 33929
rect 34669 33895 35035 33929
rect 35069 33895 35435 33929
rect 35469 33895 35835 33929
rect 35869 33895 36235 33929
rect 36269 33895 36635 33929
rect 36669 33895 37035 33929
rect 37069 33895 37435 33929
rect 37469 33895 37835 33929
rect 37869 33895 38235 33929
rect 38269 33895 38635 33929
rect 38669 33895 39035 33929
rect 39069 33895 39435 33929
rect 39469 33895 39835 33929
rect 39869 33895 40235 33929
rect 40269 33895 40635 33929
rect 40669 33895 40820 33929
rect 33652 33882 40820 33895
rect 41784 33929 52504 33942
rect 41784 33895 41967 33929
rect 42001 33895 42167 33929
rect 42201 33895 42367 33929
rect 42401 33895 42567 33929
rect 42601 33895 42767 33929
rect 42801 33895 42967 33929
rect 43001 33895 43167 33929
rect 43201 33895 43367 33929
rect 43401 33895 43567 33929
rect 43601 33895 43767 33929
rect 43801 33895 43967 33929
rect 44001 33895 44167 33929
rect 44201 33895 44367 33929
rect 44401 33895 44567 33929
rect 44601 33895 44767 33929
rect 44801 33895 44967 33929
rect 45001 33895 45167 33929
rect 45201 33895 45367 33929
rect 45401 33895 45567 33929
rect 45601 33895 45767 33929
rect 45801 33895 45967 33929
rect 46001 33895 46167 33929
rect 46201 33895 46367 33929
rect 46401 33895 46567 33929
rect 46601 33895 46767 33929
rect 46801 33895 46967 33929
rect 47001 33895 47167 33929
rect 47201 33895 47367 33929
rect 47401 33895 47567 33929
rect 47601 33895 47767 33929
rect 47801 33895 47967 33929
rect 48001 33895 48167 33929
rect 48201 33895 48367 33929
rect 48401 33895 48567 33929
rect 48601 33895 48767 33929
rect 48801 33895 48967 33929
rect 49001 33895 49167 33929
rect 49201 33895 49367 33929
rect 49401 33895 49567 33929
rect 49601 33895 49767 33929
rect 49801 33895 49967 33929
rect 50001 33895 50167 33929
rect 50201 33895 50367 33929
rect 50401 33895 50567 33929
rect 50601 33895 50767 33929
rect 50801 33895 50967 33929
rect 51001 33895 51167 33929
rect 51201 33895 51367 33929
rect 51401 33895 51567 33929
rect 51601 33895 51767 33929
rect 51801 33895 51967 33929
rect 52001 33895 52167 33929
rect 52201 33895 52367 33929
rect 52401 33895 52504 33929
rect 41784 33882 52504 33895
rect 20176 32963 20792 33002
rect 20176 32861 20263 32963
rect 20705 32861 20792 32963
rect 20176 32062 20792 32861
rect 21272 32717 21704 33107
rect 23208 32963 23824 33002
rect 23208 32861 23295 32963
rect 23737 32861 23824 32963
rect 23208 32062 23824 32861
rect 24591 32717 25023 33107
rect 41810 33596 52478 33616
rect 41810 33562 41830 33596
rect 41864 33562 41920 33596
rect 41954 33581 42010 33596
rect 42044 33581 42100 33596
rect 42134 33581 42190 33596
rect 42224 33581 42280 33596
rect 42314 33581 42370 33596
rect 42404 33581 42460 33596
rect 42494 33581 42550 33596
rect 42584 33581 42640 33596
rect 42674 33581 42730 33596
rect 42764 33581 42820 33596
rect 42854 33581 42910 33596
rect 42944 33581 43000 33596
rect 41974 33562 42010 33581
rect 42064 33562 42100 33581
rect 42154 33562 42190 33581
rect 42244 33562 42280 33581
rect 42334 33562 42370 33581
rect 42424 33562 42460 33581
rect 42514 33562 42550 33581
rect 42604 33562 42640 33581
rect 42694 33562 42730 33581
rect 42784 33562 42820 33581
rect 42874 33562 42910 33581
rect 42964 33562 43000 33581
rect 43034 33562 43170 33596
rect 43204 33562 43260 33596
rect 43294 33581 43350 33596
rect 43384 33581 43440 33596
rect 43474 33581 43530 33596
rect 43564 33581 43620 33596
rect 43654 33581 43710 33596
rect 43744 33581 43800 33596
rect 43834 33581 43890 33596
rect 43924 33581 43980 33596
rect 44014 33581 44070 33596
rect 44104 33581 44160 33596
rect 44194 33581 44250 33596
rect 44284 33581 44340 33596
rect 43314 33562 43350 33581
rect 43404 33562 43440 33581
rect 43494 33562 43530 33581
rect 43584 33562 43620 33581
rect 43674 33562 43710 33581
rect 43764 33562 43800 33581
rect 43854 33562 43890 33581
rect 43944 33562 43980 33581
rect 44034 33562 44070 33581
rect 44124 33562 44160 33581
rect 44214 33562 44250 33581
rect 44304 33562 44340 33581
rect 44374 33562 44510 33596
rect 44544 33562 44600 33596
rect 44634 33581 44690 33596
rect 44724 33581 44780 33596
rect 44814 33581 44870 33596
rect 44904 33581 44960 33596
rect 44994 33581 45050 33596
rect 45084 33581 45140 33596
rect 45174 33581 45230 33596
rect 45264 33581 45320 33596
rect 45354 33581 45410 33596
rect 45444 33581 45500 33596
rect 45534 33581 45590 33596
rect 45624 33581 45680 33596
rect 44654 33562 44690 33581
rect 44744 33562 44780 33581
rect 44834 33562 44870 33581
rect 44924 33562 44960 33581
rect 45014 33562 45050 33581
rect 45104 33562 45140 33581
rect 45194 33562 45230 33581
rect 45284 33562 45320 33581
rect 45374 33562 45410 33581
rect 45464 33562 45500 33581
rect 45554 33562 45590 33581
rect 45644 33562 45680 33581
rect 45714 33562 45850 33596
rect 45884 33562 45940 33596
rect 45974 33581 46030 33596
rect 46064 33581 46120 33596
rect 46154 33581 46210 33596
rect 46244 33581 46300 33596
rect 46334 33581 46390 33596
rect 46424 33581 46480 33596
rect 46514 33581 46570 33596
rect 46604 33581 46660 33596
rect 46694 33581 46750 33596
rect 46784 33581 46840 33596
rect 46874 33581 46930 33596
rect 46964 33581 47020 33596
rect 45994 33562 46030 33581
rect 46084 33562 46120 33581
rect 46174 33562 46210 33581
rect 46264 33562 46300 33581
rect 46354 33562 46390 33581
rect 46444 33562 46480 33581
rect 46534 33562 46570 33581
rect 46624 33562 46660 33581
rect 46714 33562 46750 33581
rect 46804 33562 46840 33581
rect 46894 33562 46930 33581
rect 46984 33562 47020 33581
rect 47054 33562 47190 33596
rect 47224 33562 47280 33596
rect 47314 33581 47370 33596
rect 47404 33581 47460 33596
rect 47494 33581 47550 33596
rect 47584 33581 47640 33596
rect 47674 33581 47730 33596
rect 47764 33581 47820 33596
rect 47854 33581 47910 33596
rect 47944 33581 48000 33596
rect 48034 33581 48090 33596
rect 48124 33581 48180 33596
rect 48214 33581 48270 33596
rect 48304 33581 48360 33596
rect 47334 33562 47370 33581
rect 47424 33562 47460 33581
rect 47514 33562 47550 33581
rect 47604 33562 47640 33581
rect 47694 33562 47730 33581
rect 47784 33562 47820 33581
rect 47874 33562 47910 33581
rect 47964 33562 48000 33581
rect 48054 33562 48090 33581
rect 48144 33562 48180 33581
rect 48234 33562 48270 33581
rect 48324 33562 48360 33581
rect 48394 33562 48530 33596
rect 48564 33562 48620 33596
rect 48654 33581 48710 33596
rect 48744 33581 48800 33596
rect 48834 33581 48890 33596
rect 48924 33581 48980 33596
rect 49014 33581 49070 33596
rect 49104 33581 49160 33596
rect 49194 33581 49250 33596
rect 49284 33581 49340 33596
rect 49374 33581 49430 33596
rect 49464 33581 49520 33596
rect 49554 33581 49610 33596
rect 49644 33581 49700 33596
rect 48674 33562 48710 33581
rect 48764 33562 48800 33581
rect 48854 33562 48890 33581
rect 48944 33562 48980 33581
rect 49034 33562 49070 33581
rect 49124 33562 49160 33581
rect 49214 33562 49250 33581
rect 49304 33562 49340 33581
rect 49394 33562 49430 33581
rect 49484 33562 49520 33581
rect 49574 33562 49610 33581
rect 49664 33562 49700 33581
rect 49734 33562 49870 33596
rect 49904 33562 49960 33596
rect 49994 33581 50050 33596
rect 50084 33581 50140 33596
rect 50174 33581 50230 33596
rect 50264 33581 50320 33596
rect 50354 33581 50410 33596
rect 50444 33581 50500 33596
rect 50534 33581 50590 33596
rect 50624 33581 50680 33596
rect 50714 33581 50770 33596
rect 50804 33581 50860 33596
rect 50894 33581 50950 33596
rect 50984 33581 51040 33596
rect 50014 33562 50050 33581
rect 50104 33562 50140 33581
rect 50194 33562 50230 33581
rect 50284 33562 50320 33581
rect 50374 33562 50410 33581
rect 50464 33562 50500 33581
rect 50554 33562 50590 33581
rect 50644 33562 50680 33581
rect 50734 33562 50770 33581
rect 50824 33562 50860 33581
rect 50914 33562 50950 33581
rect 51004 33562 51040 33581
rect 51074 33562 51210 33596
rect 51244 33562 51300 33596
rect 51334 33581 51390 33596
rect 51424 33581 51480 33596
rect 51514 33581 51570 33596
rect 51604 33581 51660 33596
rect 51694 33581 51750 33596
rect 51784 33581 51840 33596
rect 51874 33581 51930 33596
rect 51964 33581 52020 33596
rect 52054 33581 52110 33596
rect 52144 33581 52200 33596
rect 52234 33581 52290 33596
rect 52324 33581 52380 33596
rect 51354 33562 51390 33581
rect 51444 33562 51480 33581
rect 51534 33562 51570 33581
rect 51624 33562 51660 33581
rect 51714 33562 51750 33581
rect 51804 33562 51840 33581
rect 51894 33562 51930 33581
rect 51984 33562 52020 33581
rect 52074 33562 52110 33581
rect 52164 33562 52200 33581
rect 52254 33562 52290 33581
rect 52344 33562 52380 33581
rect 52414 33562 52478 33596
rect 41810 33558 41940 33562
rect 41810 33524 41844 33558
rect 41878 33547 41940 33558
rect 41974 33547 42030 33562
rect 42064 33547 42120 33562
rect 42154 33547 42210 33562
rect 42244 33547 42300 33562
rect 42334 33547 42390 33562
rect 42424 33547 42480 33562
rect 42514 33547 42570 33562
rect 42604 33547 42660 33562
rect 42694 33547 42750 33562
rect 42784 33547 42840 33562
rect 42874 33547 42930 33562
rect 42964 33558 43280 33562
rect 42964 33547 43031 33558
rect 41878 33524 43031 33547
rect 43065 33524 43184 33558
rect 43218 33547 43280 33558
rect 43314 33547 43370 33562
rect 43404 33547 43460 33562
rect 43494 33547 43550 33562
rect 43584 33547 43640 33562
rect 43674 33547 43730 33562
rect 43764 33547 43820 33562
rect 43854 33547 43910 33562
rect 43944 33547 44000 33562
rect 44034 33547 44090 33562
rect 44124 33547 44180 33562
rect 44214 33547 44270 33562
rect 44304 33558 44620 33562
rect 44304 33547 44371 33558
rect 43218 33524 44371 33547
rect 44405 33524 44524 33558
rect 44558 33547 44620 33558
rect 44654 33547 44710 33562
rect 44744 33547 44800 33562
rect 44834 33547 44890 33562
rect 44924 33547 44980 33562
rect 45014 33547 45070 33562
rect 45104 33547 45160 33562
rect 45194 33547 45250 33562
rect 45284 33547 45340 33562
rect 45374 33547 45430 33562
rect 45464 33547 45520 33562
rect 45554 33547 45610 33562
rect 45644 33558 45960 33562
rect 45644 33547 45711 33558
rect 44558 33524 45711 33547
rect 45745 33524 45864 33558
rect 45898 33547 45960 33558
rect 45994 33547 46050 33562
rect 46084 33547 46140 33562
rect 46174 33547 46230 33562
rect 46264 33547 46320 33562
rect 46354 33547 46410 33562
rect 46444 33547 46500 33562
rect 46534 33547 46590 33562
rect 46624 33547 46680 33562
rect 46714 33547 46770 33562
rect 46804 33547 46860 33562
rect 46894 33547 46950 33562
rect 46984 33558 47300 33562
rect 46984 33547 47051 33558
rect 45898 33524 47051 33547
rect 47085 33524 47204 33558
rect 47238 33547 47300 33558
rect 47334 33547 47390 33562
rect 47424 33547 47480 33562
rect 47514 33547 47570 33562
rect 47604 33547 47660 33562
rect 47694 33547 47750 33562
rect 47784 33547 47840 33562
rect 47874 33547 47930 33562
rect 47964 33547 48020 33562
rect 48054 33547 48110 33562
rect 48144 33547 48200 33562
rect 48234 33547 48290 33562
rect 48324 33558 48640 33562
rect 48324 33547 48391 33558
rect 47238 33524 48391 33547
rect 48425 33524 48544 33558
rect 48578 33547 48640 33558
rect 48674 33547 48730 33562
rect 48764 33547 48820 33562
rect 48854 33547 48910 33562
rect 48944 33547 49000 33562
rect 49034 33547 49090 33562
rect 49124 33547 49180 33562
rect 49214 33547 49270 33562
rect 49304 33547 49360 33562
rect 49394 33547 49450 33562
rect 49484 33547 49540 33562
rect 49574 33547 49630 33562
rect 49664 33558 49980 33562
rect 49664 33547 49731 33558
rect 48578 33524 49731 33547
rect 49765 33524 49884 33558
rect 49918 33547 49980 33558
rect 50014 33547 50070 33562
rect 50104 33547 50160 33562
rect 50194 33547 50250 33562
rect 50284 33547 50340 33562
rect 50374 33547 50430 33562
rect 50464 33547 50520 33562
rect 50554 33547 50610 33562
rect 50644 33547 50700 33562
rect 50734 33547 50790 33562
rect 50824 33547 50880 33562
rect 50914 33547 50970 33562
rect 51004 33558 51320 33562
rect 51004 33547 51071 33558
rect 49918 33524 51071 33547
rect 51105 33524 51224 33558
rect 51258 33547 51320 33558
rect 51354 33547 51410 33562
rect 51444 33547 51500 33562
rect 51534 33547 51590 33562
rect 51624 33547 51680 33562
rect 51714 33547 51770 33562
rect 51804 33547 51860 33562
rect 51894 33547 51950 33562
rect 51984 33547 52040 33562
rect 52074 33547 52130 33562
rect 52164 33547 52220 33562
rect 52254 33547 52310 33562
rect 52344 33558 52478 33562
rect 52344 33547 52411 33558
rect 51258 33524 52411 33547
rect 52445 33524 52478 33558
rect 41810 33517 52478 33524
rect 41810 33468 41909 33517
rect 41810 33434 41844 33468
rect 41878 33434 41909 33468
rect 42999 33468 43249 33517
rect 41810 33378 41909 33434
rect 41810 33344 41844 33378
rect 41878 33344 41909 33378
rect 41810 33288 41909 33344
rect 41810 33254 41844 33288
rect 41878 33254 41909 33288
rect 41810 33198 41909 33254
rect 41810 33164 41844 33198
rect 41878 33164 41909 33198
rect 41810 33108 41909 33164
rect 41810 33074 41844 33108
rect 41878 33074 41909 33108
rect 41810 33018 41909 33074
rect 41810 32984 41844 33018
rect 41878 32984 41909 33018
rect 41810 32928 41909 32984
rect 41810 32894 41844 32928
rect 41878 32894 41909 32928
rect 41810 32838 41909 32894
rect 41810 32804 41844 32838
rect 41878 32804 41909 32838
rect 41810 32748 41909 32804
rect 41810 32714 41844 32748
rect 41878 32714 41909 32748
rect 41810 32658 41909 32714
rect 41810 32624 41844 32658
rect 41878 32624 41909 32658
rect 41810 32568 41909 32624
rect 41810 32534 41844 32568
rect 41878 32534 41909 32568
rect 41810 32478 41909 32534
rect 41973 33436 42935 33453
rect 41973 33402 41994 33436
rect 42028 33402 42084 33436
rect 42118 33434 42174 33436
rect 42208 33434 42264 33436
rect 42298 33434 42354 33436
rect 42388 33434 42444 33436
rect 42478 33434 42534 33436
rect 42568 33434 42624 33436
rect 42658 33434 42714 33436
rect 42748 33434 42804 33436
rect 42838 33434 42894 33436
rect 42138 33402 42174 33434
rect 42228 33402 42264 33434
rect 42318 33402 42354 33434
rect 42408 33402 42444 33434
rect 42498 33402 42534 33434
rect 42588 33402 42624 33434
rect 42678 33402 42714 33434
rect 42768 33402 42804 33434
rect 42858 33402 42894 33434
rect 42928 33402 42935 33436
rect 41973 33400 42104 33402
rect 42138 33400 42194 33402
rect 42228 33400 42284 33402
rect 42318 33400 42374 33402
rect 42408 33400 42464 33402
rect 42498 33400 42554 33402
rect 42588 33400 42644 33402
rect 42678 33400 42734 33402
rect 42768 33400 42824 33402
rect 42858 33400 42935 33402
rect 41973 33381 42935 33400
rect 41973 33377 42045 33381
rect 41973 33343 41992 33377
rect 42026 33343 42045 33377
rect 41973 33287 42045 33343
rect 42863 33358 42935 33381
rect 42863 33324 42882 33358
rect 42916 33324 42935 33358
rect 41973 33253 41992 33287
rect 42026 33253 42045 33287
rect 41973 33197 42045 33253
rect 41973 33163 41992 33197
rect 42026 33163 42045 33197
rect 41973 33107 42045 33163
rect 41973 33073 41992 33107
rect 42026 33073 42045 33107
rect 41973 33017 42045 33073
rect 41973 32983 41992 33017
rect 42026 32983 42045 33017
rect 41973 32927 42045 32983
rect 41973 32893 41992 32927
rect 42026 32893 42045 32927
rect 41973 32837 42045 32893
rect 41973 32803 41992 32837
rect 42026 32803 42045 32837
rect 41973 32747 42045 32803
rect 41973 32713 41992 32747
rect 42026 32713 42045 32747
rect 41973 32657 42045 32713
rect 41973 32623 41992 32657
rect 42026 32623 42045 32657
rect 42107 33260 42801 33319
rect 42107 33226 42168 33260
rect 42202 33232 42258 33260
rect 42292 33232 42348 33260
rect 42382 33232 42438 33260
rect 42214 33226 42258 33232
rect 42314 33226 42348 33232
rect 42414 33226 42438 33232
rect 42472 33232 42528 33260
rect 42472 33226 42480 33232
rect 42107 33198 42180 33226
rect 42214 33198 42280 33226
rect 42314 33198 42380 33226
rect 42414 33198 42480 33226
rect 42514 33226 42528 33232
rect 42562 33232 42618 33260
rect 42562 33226 42580 33232
rect 42514 33198 42580 33226
rect 42614 33226 42618 33232
rect 42652 33232 42708 33260
rect 42652 33226 42680 33232
rect 42742 33226 42801 33260
rect 42614 33198 42680 33226
rect 42714 33198 42801 33226
rect 42107 33170 42801 33198
rect 42107 33136 42168 33170
rect 42202 33136 42258 33170
rect 42292 33136 42348 33170
rect 42382 33136 42438 33170
rect 42472 33136 42528 33170
rect 42562 33136 42618 33170
rect 42652 33136 42708 33170
rect 42742 33136 42801 33170
rect 42107 33132 42801 33136
rect 42107 33098 42180 33132
rect 42214 33098 42280 33132
rect 42314 33098 42380 33132
rect 42414 33098 42480 33132
rect 42514 33098 42580 33132
rect 42614 33098 42680 33132
rect 42714 33098 42801 33132
rect 42107 33080 42801 33098
rect 42107 33046 42168 33080
rect 42202 33046 42258 33080
rect 42292 33046 42348 33080
rect 42382 33046 42438 33080
rect 42472 33046 42528 33080
rect 42562 33046 42618 33080
rect 42652 33046 42708 33080
rect 42742 33046 42801 33080
rect 42107 33032 42801 33046
rect 42107 32998 42180 33032
rect 42214 32998 42280 33032
rect 42314 32998 42380 33032
rect 42414 32998 42480 33032
rect 42514 32998 42580 33032
rect 42614 32998 42680 33032
rect 42714 32998 42801 33032
rect 42107 32990 42801 32998
rect 42107 32956 42168 32990
rect 42202 32956 42258 32990
rect 42292 32956 42348 32990
rect 42382 32956 42438 32990
rect 42472 32956 42528 32990
rect 42562 32956 42618 32990
rect 42652 32956 42708 32990
rect 42742 32956 42801 32990
rect 42107 32932 42801 32956
rect 42107 32900 42180 32932
rect 42214 32900 42280 32932
rect 42314 32900 42380 32932
rect 42414 32900 42480 32932
rect 42107 32866 42168 32900
rect 42214 32898 42258 32900
rect 42314 32898 42348 32900
rect 42414 32898 42438 32900
rect 42202 32866 42258 32898
rect 42292 32866 42348 32898
rect 42382 32866 42438 32898
rect 42472 32898 42480 32900
rect 42514 32900 42580 32932
rect 42514 32898 42528 32900
rect 42472 32866 42528 32898
rect 42562 32898 42580 32900
rect 42614 32900 42680 32932
rect 42714 32900 42801 32932
rect 42614 32898 42618 32900
rect 42562 32866 42618 32898
rect 42652 32898 42680 32900
rect 42652 32866 42708 32898
rect 42742 32866 42801 32900
rect 42107 32832 42801 32866
rect 42107 32810 42180 32832
rect 42214 32810 42280 32832
rect 42314 32810 42380 32832
rect 42414 32810 42480 32832
rect 42107 32776 42168 32810
rect 42214 32798 42258 32810
rect 42314 32798 42348 32810
rect 42414 32798 42438 32810
rect 42202 32776 42258 32798
rect 42292 32776 42348 32798
rect 42382 32776 42438 32798
rect 42472 32798 42480 32810
rect 42514 32810 42580 32832
rect 42514 32798 42528 32810
rect 42472 32776 42528 32798
rect 42562 32798 42580 32810
rect 42614 32810 42680 32832
rect 42714 32810 42801 32832
rect 42614 32798 42618 32810
rect 42562 32776 42618 32798
rect 42652 32798 42680 32810
rect 42652 32776 42708 32798
rect 42742 32776 42801 32810
rect 42107 32732 42801 32776
rect 42107 32720 42180 32732
rect 42214 32720 42280 32732
rect 42314 32720 42380 32732
rect 42414 32720 42480 32732
rect 42107 32686 42168 32720
rect 42214 32698 42258 32720
rect 42314 32698 42348 32720
rect 42414 32698 42438 32720
rect 42202 32686 42258 32698
rect 42292 32686 42348 32698
rect 42382 32686 42438 32698
rect 42472 32698 42480 32720
rect 42514 32720 42580 32732
rect 42514 32698 42528 32720
rect 42472 32686 42528 32698
rect 42562 32698 42580 32720
rect 42614 32720 42680 32732
rect 42714 32720 42801 32732
rect 42614 32698 42618 32720
rect 42562 32686 42618 32698
rect 42652 32698 42680 32720
rect 42652 32686 42708 32698
rect 42742 32686 42801 32720
rect 42107 32625 42801 32686
rect 42863 33268 42935 33324
rect 42863 33234 42882 33268
rect 42916 33234 42935 33268
rect 42863 33178 42935 33234
rect 42863 33144 42882 33178
rect 42916 33144 42935 33178
rect 42863 33088 42935 33144
rect 42863 33054 42882 33088
rect 42916 33054 42935 33088
rect 42863 32998 42935 33054
rect 42863 32964 42882 32998
rect 42916 32964 42935 32998
rect 42863 32908 42935 32964
rect 42863 32874 42882 32908
rect 42916 32874 42935 32908
rect 42863 32818 42935 32874
rect 42863 32784 42882 32818
rect 42916 32784 42935 32818
rect 42863 32728 42935 32784
rect 42863 32694 42882 32728
rect 42916 32694 42935 32728
rect 42863 32638 42935 32694
rect 41973 32563 42045 32623
rect 42863 32604 42882 32638
rect 42916 32604 42935 32638
rect 42863 32563 42935 32604
rect 41973 32544 42935 32563
rect 41973 32510 42070 32544
rect 42104 32510 42160 32544
rect 42194 32510 42250 32544
rect 42284 32510 42340 32544
rect 42374 32510 42430 32544
rect 42464 32510 42520 32544
rect 42554 32510 42610 32544
rect 42644 32510 42700 32544
rect 42734 32510 42790 32544
rect 42824 32510 42935 32544
rect 41973 32491 42935 32510
rect 42999 33434 43031 33468
rect 43065 33434 43184 33468
rect 43218 33434 43249 33468
rect 44339 33468 44589 33517
rect 42999 33378 43249 33434
rect 42999 33344 43031 33378
rect 43065 33344 43184 33378
rect 43218 33344 43249 33378
rect 42999 33288 43249 33344
rect 42999 33254 43031 33288
rect 43065 33254 43184 33288
rect 43218 33254 43249 33288
rect 42999 33198 43249 33254
rect 42999 33164 43031 33198
rect 43065 33164 43184 33198
rect 43218 33164 43249 33198
rect 42999 33108 43249 33164
rect 42999 33074 43031 33108
rect 43065 33074 43184 33108
rect 43218 33074 43249 33108
rect 42999 33018 43249 33074
rect 42999 32984 43031 33018
rect 43065 32984 43184 33018
rect 43218 32984 43249 33018
rect 42999 32928 43249 32984
rect 42999 32894 43031 32928
rect 43065 32894 43184 32928
rect 43218 32894 43249 32928
rect 42999 32838 43249 32894
rect 42999 32804 43031 32838
rect 43065 32804 43184 32838
rect 43218 32804 43249 32838
rect 42999 32748 43249 32804
rect 42999 32714 43031 32748
rect 43065 32714 43184 32748
rect 43218 32714 43249 32748
rect 42999 32658 43249 32714
rect 42999 32624 43031 32658
rect 43065 32624 43184 32658
rect 43218 32624 43249 32658
rect 42999 32568 43249 32624
rect 42999 32534 43031 32568
rect 43065 32534 43184 32568
rect 43218 32534 43249 32568
rect 41810 32444 41844 32478
rect 41878 32444 41909 32478
rect 41810 32427 41909 32444
rect 42999 32478 43249 32534
rect 43313 33436 44275 33453
rect 43313 33402 43334 33436
rect 43368 33402 43424 33436
rect 43458 33434 43514 33436
rect 43548 33434 43604 33436
rect 43638 33434 43694 33436
rect 43728 33434 43784 33436
rect 43818 33434 43874 33436
rect 43908 33434 43964 33436
rect 43998 33434 44054 33436
rect 44088 33434 44144 33436
rect 44178 33434 44234 33436
rect 43478 33402 43514 33434
rect 43568 33402 43604 33434
rect 43658 33402 43694 33434
rect 43748 33402 43784 33434
rect 43838 33402 43874 33434
rect 43928 33402 43964 33434
rect 44018 33402 44054 33434
rect 44108 33402 44144 33434
rect 44198 33402 44234 33434
rect 44268 33402 44275 33436
rect 43313 33400 43444 33402
rect 43478 33400 43534 33402
rect 43568 33400 43624 33402
rect 43658 33400 43714 33402
rect 43748 33400 43804 33402
rect 43838 33400 43894 33402
rect 43928 33400 43984 33402
rect 44018 33400 44074 33402
rect 44108 33400 44164 33402
rect 44198 33400 44275 33402
rect 43313 33381 44275 33400
rect 43313 33377 43385 33381
rect 43313 33343 43332 33377
rect 43366 33343 43385 33377
rect 43313 33287 43385 33343
rect 44203 33358 44275 33381
rect 44203 33324 44222 33358
rect 44256 33324 44275 33358
rect 43313 33253 43332 33287
rect 43366 33253 43385 33287
rect 43313 33197 43385 33253
rect 43313 33163 43332 33197
rect 43366 33163 43385 33197
rect 43313 33107 43385 33163
rect 43313 33073 43332 33107
rect 43366 33073 43385 33107
rect 43313 33017 43385 33073
rect 43313 32983 43332 33017
rect 43366 32983 43385 33017
rect 43313 32927 43385 32983
rect 43313 32893 43332 32927
rect 43366 32893 43385 32927
rect 43313 32837 43385 32893
rect 43313 32803 43332 32837
rect 43366 32803 43385 32837
rect 43313 32747 43385 32803
rect 43313 32713 43332 32747
rect 43366 32713 43385 32747
rect 43313 32657 43385 32713
rect 43313 32623 43332 32657
rect 43366 32623 43385 32657
rect 43447 33260 44141 33319
rect 43447 33226 43508 33260
rect 43542 33232 43598 33260
rect 43632 33232 43688 33260
rect 43722 33232 43778 33260
rect 43554 33226 43598 33232
rect 43654 33226 43688 33232
rect 43754 33226 43778 33232
rect 43812 33232 43868 33260
rect 43812 33226 43820 33232
rect 43447 33198 43520 33226
rect 43554 33198 43620 33226
rect 43654 33198 43720 33226
rect 43754 33198 43820 33226
rect 43854 33226 43868 33232
rect 43902 33232 43958 33260
rect 43902 33226 43920 33232
rect 43854 33198 43920 33226
rect 43954 33226 43958 33232
rect 43992 33232 44048 33260
rect 43992 33226 44020 33232
rect 44082 33226 44141 33260
rect 43954 33198 44020 33226
rect 44054 33198 44141 33226
rect 43447 33170 44141 33198
rect 43447 33136 43508 33170
rect 43542 33136 43598 33170
rect 43632 33136 43688 33170
rect 43722 33136 43778 33170
rect 43812 33136 43868 33170
rect 43902 33136 43958 33170
rect 43992 33136 44048 33170
rect 44082 33136 44141 33170
rect 43447 33132 44141 33136
rect 43447 33098 43520 33132
rect 43554 33098 43620 33132
rect 43654 33098 43720 33132
rect 43754 33098 43820 33132
rect 43854 33098 43920 33132
rect 43954 33098 44020 33132
rect 44054 33098 44141 33132
rect 43447 33080 44141 33098
rect 43447 33046 43508 33080
rect 43542 33046 43598 33080
rect 43632 33046 43688 33080
rect 43722 33046 43778 33080
rect 43812 33046 43868 33080
rect 43902 33046 43958 33080
rect 43992 33046 44048 33080
rect 44082 33046 44141 33080
rect 43447 33032 44141 33046
rect 43447 32998 43520 33032
rect 43554 32998 43620 33032
rect 43654 32998 43720 33032
rect 43754 32998 43820 33032
rect 43854 32998 43920 33032
rect 43954 32998 44020 33032
rect 44054 32998 44141 33032
rect 43447 32990 44141 32998
rect 43447 32956 43508 32990
rect 43542 32956 43598 32990
rect 43632 32956 43688 32990
rect 43722 32956 43778 32990
rect 43812 32956 43868 32990
rect 43902 32956 43958 32990
rect 43992 32956 44048 32990
rect 44082 32956 44141 32990
rect 43447 32932 44141 32956
rect 43447 32900 43520 32932
rect 43554 32900 43620 32932
rect 43654 32900 43720 32932
rect 43754 32900 43820 32932
rect 43447 32866 43508 32900
rect 43554 32898 43598 32900
rect 43654 32898 43688 32900
rect 43754 32898 43778 32900
rect 43542 32866 43598 32898
rect 43632 32866 43688 32898
rect 43722 32866 43778 32898
rect 43812 32898 43820 32900
rect 43854 32900 43920 32932
rect 43854 32898 43868 32900
rect 43812 32866 43868 32898
rect 43902 32898 43920 32900
rect 43954 32900 44020 32932
rect 44054 32900 44141 32932
rect 43954 32898 43958 32900
rect 43902 32866 43958 32898
rect 43992 32898 44020 32900
rect 43992 32866 44048 32898
rect 44082 32866 44141 32900
rect 43447 32832 44141 32866
rect 43447 32810 43520 32832
rect 43554 32810 43620 32832
rect 43654 32810 43720 32832
rect 43754 32810 43820 32832
rect 43447 32776 43508 32810
rect 43554 32798 43598 32810
rect 43654 32798 43688 32810
rect 43754 32798 43778 32810
rect 43542 32776 43598 32798
rect 43632 32776 43688 32798
rect 43722 32776 43778 32798
rect 43812 32798 43820 32810
rect 43854 32810 43920 32832
rect 43854 32798 43868 32810
rect 43812 32776 43868 32798
rect 43902 32798 43920 32810
rect 43954 32810 44020 32832
rect 44054 32810 44141 32832
rect 43954 32798 43958 32810
rect 43902 32776 43958 32798
rect 43992 32798 44020 32810
rect 43992 32776 44048 32798
rect 44082 32776 44141 32810
rect 43447 32732 44141 32776
rect 43447 32720 43520 32732
rect 43554 32720 43620 32732
rect 43654 32720 43720 32732
rect 43754 32720 43820 32732
rect 43447 32686 43508 32720
rect 43554 32698 43598 32720
rect 43654 32698 43688 32720
rect 43754 32698 43778 32720
rect 43542 32686 43598 32698
rect 43632 32686 43688 32698
rect 43722 32686 43778 32698
rect 43812 32698 43820 32720
rect 43854 32720 43920 32732
rect 43854 32698 43868 32720
rect 43812 32686 43868 32698
rect 43902 32698 43920 32720
rect 43954 32720 44020 32732
rect 44054 32720 44141 32732
rect 43954 32698 43958 32720
rect 43902 32686 43958 32698
rect 43992 32698 44020 32720
rect 43992 32686 44048 32698
rect 44082 32686 44141 32720
rect 43447 32625 44141 32686
rect 44203 33268 44275 33324
rect 44203 33234 44222 33268
rect 44256 33234 44275 33268
rect 44203 33178 44275 33234
rect 44203 33144 44222 33178
rect 44256 33144 44275 33178
rect 44203 33088 44275 33144
rect 44203 33054 44222 33088
rect 44256 33054 44275 33088
rect 44203 32998 44275 33054
rect 44203 32964 44222 32998
rect 44256 32964 44275 32998
rect 44203 32908 44275 32964
rect 44203 32874 44222 32908
rect 44256 32874 44275 32908
rect 44203 32818 44275 32874
rect 44203 32784 44222 32818
rect 44256 32784 44275 32818
rect 44203 32728 44275 32784
rect 44203 32694 44222 32728
rect 44256 32694 44275 32728
rect 44203 32638 44275 32694
rect 43313 32563 43385 32623
rect 44203 32604 44222 32638
rect 44256 32604 44275 32638
rect 44203 32563 44275 32604
rect 43313 32544 44275 32563
rect 43313 32510 43410 32544
rect 43444 32510 43500 32544
rect 43534 32510 43590 32544
rect 43624 32510 43680 32544
rect 43714 32510 43770 32544
rect 43804 32510 43860 32544
rect 43894 32510 43950 32544
rect 43984 32510 44040 32544
rect 44074 32510 44130 32544
rect 44164 32510 44275 32544
rect 43313 32491 44275 32510
rect 44339 33434 44371 33468
rect 44405 33434 44524 33468
rect 44558 33434 44589 33468
rect 45679 33468 45929 33517
rect 44339 33378 44589 33434
rect 44339 33344 44371 33378
rect 44405 33344 44524 33378
rect 44558 33344 44589 33378
rect 44339 33288 44589 33344
rect 44339 33254 44371 33288
rect 44405 33254 44524 33288
rect 44558 33254 44589 33288
rect 44339 33198 44589 33254
rect 44339 33164 44371 33198
rect 44405 33164 44524 33198
rect 44558 33164 44589 33198
rect 44339 33108 44589 33164
rect 44339 33074 44371 33108
rect 44405 33074 44524 33108
rect 44558 33074 44589 33108
rect 44339 33018 44589 33074
rect 44339 32984 44371 33018
rect 44405 32984 44524 33018
rect 44558 32984 44589 33018
rect 44339 32928 44589 32984
rect 44339 32894 44371 32928
rect 44405 32894 44524 32928
rect 44558 32894 44589 32928
rect 44339 32838 44589 32894
rect 44339 32804 44371 32838
rect 44405 32804 44524 32838
rect 44558 32804 44589 32838
rect 44339 32748 44589 32804
rect 44339 32714 44371 32748
rect 44405 32714 44524 32748
rect 44558 32714 44589 32748
rect 44339 32658 44589 32714
rect 44339 32624 44371 32658
rect 44405 32624 44524 32658
rect 44558 32624 44589 32658
rect 44339 32568 44589 32624
rect 44339 32534 44371 32568
rect 44405 32534 44524 32568
rect 44558 32534 44589 32568
rect 42999 32444 43031 32478
rect 43065 32444 43184 32478
rect 43218 32444 43249 32478
rect 42999 32427 43249 32444
rect 44339 32478 44589 32534
rect 44653 33436 45615 33453
rect 44653 33402 44674 33436
rect 44708 33402 44764 33436
rect 44798 33434 44854 33436
rect 44888 33434 44944 33436
rect 44978 33434 45034 33436
rect 45068 33434 45124 33436
rect 45158 33434 45214 33436
rect 45248 33434 45304 33436
rect 45338 33434 45394 33436
rect 45428 33434 45484 33436
rect 45518 33434 45574 33436
rect 44818 33402 44854 33434
rect 44908 33402 44944 33434
rect 44998 33402 45034 33434
rect 45088 33402 45124 33434
rect 45178 33402 45214 33434
rect 45268 33402 45304 33434
rect 45358 33402 45394 33434
rect 45448 33402 45484 33434
rect 45538 33402 45574 33434
rect 45608 33402 45615 33436
rect 44653 33400 44784 33402
rect 44818 33400 44874 33402
rect 44908 33400 44964 33402
rect 44998 33400 45054 33402
rect 45088 33400 45144 33402
rect 45178 33400 45234 33402
rect 45268 33400 45324 33402
rect 45358 33400 45414 33402
rect 45448 33400 45504 33402
rect 45538 33400 45615 33402
rect 44653 33381 45615 33400
rect 44653 33377 44725 33381
rect 44653 33343 44672 33377
rect 44706 33343 44725 33377
rect 44653 33287 44725 33343
rect 45543 33358 45615 33381
rect 45543 33324 45562 33358
rect 45596 33324 45615 33358
rect 44653 33253 44672 33287
rect 44706 33253 44725 33287
rect 44653 33197 44725 33253
rect 44653 33163 44672 33197
rect 44706 33163 44725 33197
rect 44653 33107 44725 33163
rect 44653 33073 44672 33107
rect 44706 33073 44725 33107
rect 44653 33017 44725 33073
rect 44653 32983 44672 33017
rect 44706 32983 44725 33017
rect 44653 32927 44725 32983
rect 44653 32893 44672 32927
rect 44706 32893 44725 32927
rect 44653 32837 44725 32893
rect 44653 32803 44672 32837
rect 44706 32803 44725 32837
rect 44653 32747 44725 32803
rect 44653 32713 44672 32747
rect 44706 32713 44725 32747
rect 44653 32657 44725 32713
rect 44653 32623 44672 32657
rect 44706 32623 44725 32657
rect 44787 33260 45481 33319
rect 44787 33226 44848 33260
rect 44882 33232 44938 33260
rect 44972 33232 45028 33260
rect 45062 33232 45118 33260
rect 44894 33226 44938 33232
rect 44994 33226 45028 33232
rect 45094 33226 45118 33232
rect 45152 33232 45208 33260
rect 45152 33226 45160 33232
rect 44787 33198 44860 33226
rect 44894 33198 44960 33226
rect 44994 33198 45060 33226
rect 45094 33198 45160 33226
rect 45194 33226 45208 33232
rect 45242 33232 45298 33260
rect 45242 33226 45260 33232
rect 45194 33198 45260 33226
rect 45294 33226 45298 33232
rect 45332 33232 45388 33260
rect 45332 33226 45360 33232
rect 45422 33226 45481 33260
rect 45294 33198 45360 33226
rect 45394 33198 45481 33226
rect 44787 33170 45481 33198
rect 44787 33136 44848 33170
rect 44882 33136 44938 33170
rect 44972 33136 45028 33170
rect 45062 33136 45118 33170
rect 45152 33136 45208 33170
rect 45242 33136 45298 33170
rect 45332 33136 45388 33170
rect 45422 33136 45481 33170
rect 44787 33132 45481 33136
rect 44787 33098 44860 33132
rect 44894 33098 44960 33132
rect 44994 33098 45060 33132
rect 45094 33098 45160 33132
rect 45194 33098 45260 33132
rect 45294 33098 45360 33132
rect 45394 33098 45481 33132
rect 44787 33080 45481 33098
rect 44787 33046 44848 33080
rect 44882 33046 44938 33080
rect 44972 33046 45028 33080
rect 45062 33046 45118 33080
rect 45152 33046 45208 33080
rect 45242 33046 45298 33080
rect 45332 33046 45388 33080
rect 45422 33046 45481 33080
rect 44787 33032 45481 33046
rect 44787 32998 44860 33032
rect 44894 32998 44960 33032
rect 44994 32998 45060 33032
rect 45094 32998 45160 33032
rect 45194 32998 45260 33032
rect 45294 32998 45360 33032
rect 45394 32998 45481 33032
rect 44787 32990 45481 32998
rect 44787 32956 44848 32990
rect 44882 32956 44938 32990
rect 44972 32956 45028 32990
rect 45062 32956 45118 32990
rect 45152 32956 45208 32990
rect 45242 32956 45298 32990
rect 45332 32956 45388 32990
rect 45422 32956 45481 32990
rect 44787 32932 45481 32956
rect 44787 32900 44860 32932
rect 44894 32900 44960 32932
rect 44994 32900 45060 32932
rect 45094 32900 45160 32932
rect 44787 32866 44848 32900
rect 44894 32898 44938 32900
rect 44994 32898 45028 32900
rect 45094 32898 45118 32900
rect 44882 32866 44938 32898
rect 44972 32866 45028 32898
rect 45062 32866 45118 32898
rect 45152 32898 45160 32900
rect 45194 32900 45260 32932
rect 45194 32898 45208 32900
rect 45152 32866 45208 32898
rect 45242 32898 45260 32900
rect 45294 32900 45360 32932
rect 45394 32900 45481 32932
rect 45294 32898 45298 32900
rect 45242 32866 45298 32898
rect 45332 32898 45360 32900
rect 45332 32866 45388 32898
rect 45422 32866 45481 32900
rect 44787 32832 45481 32866
rect 44787 32810 44860 32832
rect 44894 32810 44960 32832
rect 44994 32810 45060 32832
rect 45094 32810 45160 32832
rect 44787 32776 44848 32810
rect 44894 32798 44938 32810
rect 44994 32798 45028 32810
rect 45094 32798 45118 32810
rect 44882 32776 44938 32798
rect 44972 32776 45028 32798
rect 45062 32776 45118 32798
rect 45152 32798 45160 32810
rect 45194 32810 45260 32832
rect 45194 32798 45208 32810
rect 45152 32776 45208 32798
rect 45242 32798 45260 32810
rect 45294 32810 45360 32832
rect 45394 32810 45481 32832
rect 45294 32798 45298 32810
rect 45242 32776 45298 32798
rect 45332 32798 45360 32810
rect 45332 32776 45388 32798
rect 45422 32776 45481 32810
rect 44787 32732 45481 32776
rect 44787 32720 44860 32732
rect 44894 32720 44960 32732
rect 44994 32720 45060 32732
rect 45094 32720 45160 32732
rect 44787 32686 44848 32720
rect 44894 32698 44938 32720
rect 44994 32698 45028 32720
rect 45094 32698 45118 32720
rect 44882 32686 44938 32698
rect 44972 32686 45028 32698
rect 45062 32686 45118 32698
rect 45152 32698 45160 32720
rect 45194 32720 45260 32732
rect 45194 32698 45208 32720
rect 45152 32686 45208 32698
rect 45242 32698 45260 32720
rect 45294 32720 45360 32732
rect 45394 32720 45481 32732
rect 45294 32698 45298 32720
rect 45242 32686 45298 32698
rect 45332 32698 45360 32720
rect 45332 32686 45388 32698
rect 45422 32686 45481 32720
rect 44787 32625 45481 32686
rect 45543 33268 45615 33324
rect 45543 33234 45562 33268
rect 45596 33234 45615 33268
rect 45543 33178 45615 33234
rect 45543 33144 45562 33178
rect 45596 33144 45615 33178
rect 45543 33088 45615 33144
rect 45543 33054 45562 33088
rect 45596 33054 45615 33088
rect 45543 32998 45615 33054
rect 45543 32964 45562 32998
rect 45596 32964 45615 32998
rect 45543 32908 45615 32964
rect 45543 32874 45562 32908
rect 45596 32874 45615 32908
rect 45543 32818 45615 32874
rect 45543 32784 45562 32818
rect 45596 32784 45615 32818
rect 45543 32728 45615 32784
rect 45543 32694 45562 32728
rect 45596 32694 45615 32728
rect 45543 32638 45615 32694
rect 44653 32563 44725 32623
rect 45543 32604 45562 32638
rect 45596 32604 45615 32638
rect 45543 32563 45615 32604
rect 44653 32544 45615 32563
rect 44653 32510 44750 32544
rect 44784 32510 44840 32544
rect 44874 32510 44930 32544
rect 44964 32510 45020 32544
rect 45054 32510 45110 32544
rect 45144 32510 45200 32544
rect 45234 32510 45290 32544
rect 45324 32510 45380 32544
rect 45414 32510 45470 32544
rect 45504 32510 45615 32544
rect 44653 32491 45615 32510
rect 45679 33434 45711 33468
rect 45745 33434 45864 33468
rect 45898 33434 45929 33468
rect 47019 33468 47269 33517
rect 45679 33378 45929 33434
rect 45679 33344 45711 33378
rect 45745 33344 45864 33378
rect 45898 33344 45929 33378
rect 45679 33288 45929 33344
rect 45679 33254 45711 33288
rect 45745 33254 45864 33288
rect 45898 33254 45929 33288
rect 45679 33198 45929 33254
rect 45679 33164 45711 33198
rect 45745 33164 45864 33198
rect 45898 33164 45929 33198
rect 45679 33108 45929 33164
rect 45679 33074 45711 33108
rect 45745 33074 45864 33108
rect 45898 33074 45929 33108
rect 45679 33018 45929 33074
rect 45679 32984 45711 33018
rect 45745 32984 45864 33018
rect 45898 32984 45929 33018
rect 45679 32928 45929 32984
rect 45679 32894 45711 32928
rect 45745 32894 45864 32928
rect 45898 32894 45929 32928
rect 45679 32838 45929 32894
rect 45679 32804 45711 32838
rect 45745 32804 45864 32838
rect 45898 32804 45929 32838
rect 45679 32748 45929 32804
rect 45679 32714 45711 32748
rect 45745 32714 45864 32748
rect 45898 32714 45929 32748
rect 45679 32658 45929 32714
rect 45679 32624 45711 32658
rect 45745 32624 45864 32658
rect 45898 32624 45929 32658
rect 45679 32568 45929 32624
rect 45679 32534 45711 32568
rect 45745 32534 45864 32568
rect 45898 32534 45929 32568
rect 44339 32444 44371 32478
rect 44405 32444 44524 32478
rect 44558 32444 44589 32478
rect 44339 32427 44589 32444
rect 45679 32478 45929 32534
rect 45993 33436 46955 33453
rect 45993 33402 46014 33436
rect 46048 33402 46104 33436
rect 46138 33434 46194 33436
rect 46228 33434 46284 33436
rect 46318 33434 46374 33436
rect 46408 33434 46464 33436
rect 46498 33434 46554 33436
rect 46588 33434 46644 33436
rect 46678 33434 46734 33436
rect 46768 33434 46824 33436
rect 46858 33434 46914 33436
rect 46158 33402 46194 33434
rect 46248 33402 46284 33434
rect 46338 33402 46374 33434
rect 46428 33402 46464 33434
rect 46518 33402 46554 33434
rect 46608 33402 46644 33434
rect 46698 33402 46734 33434
rect 46788 33402 46824 33434
rect 46878 33402 46914 33434
rect 46948 33402 46955 33436
rect 45993 33400 46124 33402
rect 46158 33400 46214 33402
rect 46248 33400 46304 33402
rect 46338 33400 46394 33402
rect 46428 33400 46484 33402
rect 46518 33400 46574 33402
rect 46608 33400 46664 33402
rect 46698 33400 46754 33402
rect 46788 33400 46844 33402
rect 46878 33400 46955 33402
rect 45993 33381 46955 33400
rect 45993 33377 46065 33381
rect 45993 33343 46012 33377
rect 46046 33343 46065 33377
rect 45993 33287 46065 33343
rect 46883 33358 46955 33381
rect 46883 33324 46902 33358
rect 46936 33324 46955 33358
rect 45993 33253 46012 33287
rect 46046 33253 46065 33287
rect 45993 33197 46065 33253
rect 45993 33163 46012 33197
rect 46046 33163 46065 33197
rect 45993 33107 46065 33163
rect 45993 33073 46012 33107
rect 46046 33073 46065 33107
rect 45993 33017 46065 33073
rect 45993 32983 46012 33017
rect 46046 32983 46065 33017
rect 45993 32927 46065 32983
rect 45993 32893 46012 32927
rect 46046 32893 46065 32927
rect 45993 32837 46065 32893
rect 45993 32803 46012 32837
rect 46046 32803 46065 32837
rect 45993 32747 46065 32803
rect 45993 32713 46012 32747
rect 46046 32713 46065 32747
rect 45993 32657 46065 32713
rect 45993 32623 46012 32657
rect 46046 32623 46065 32657
rect 46127 33260 46821 33319
rect 46127 33226 46188 33260
rect 46222 33232 46278 33260
rect 46312 33232 46368 33260
rect 46402 33232 46458 33260
rect 46234 33226 46278 33232
rect 46334 33226 46368 33232
rect 46434 33226 46458 33232
rect 46492 33232 46548 33260
rect 46492 33226 46500 33232
rect 46127 33198 46200 33226
rect 46234 33198 46300 33226
rect 46334 33198 46400 33226
rect 46434 33198 46500 33226
rect 46534 33226 46548 33232
rect 46582 33232 46638 33260
rect 46582 33226 46600 33232
rect 46534 33198 46600 33226
rect 46634 33226 46638 33232
rect 46672 33232 46728 33260
rect 46672 33226 46700 33232
rect 46762 33226 46821 33260
rect 46634 33198 46700 33226
rect 46734 33198 46821 33226
rect 46127 33170 46821 33198
rect 46127 33136 46188 33170
rect 46222 33136 46278 33170
rect 46312 33136 46368 33170
rect 46402 33136 46458 33170
rect 46492 33136 46548 33170
rect 46582 33136 46638 33170
rect 46672 33136 46728 33170
rect 46762 33136 46821 33170
rect 46127 33132 46821 33136
rect 46127 33098 46200 33132
rect 46234 33098 46300 33132
rect 46334 33098 46400 33132
rect 46434 33098 46500 33132
rect 46534 33098 46600 33132
rect 46634 33098 46700 33132
rect 46734 33098 46821 33132
rect 46127 33080 46821 33098
rect 46127 33046 46188 33080
rect 46222 33046 46278 33080
rect 46312 33046 46368 33080
rect 46402 33046 46458 33080
rect 46492 33046 46548 33080
rect 46582 33046 46638 33080
rect 46672 33046 46728 33080
rect 46762 33046 46821 33080
rect 46127 33032 46821 33046
rect 46127 32998 46200 33032
rect 46234 32998 46300 33032
rect 46334 32998 46400 33032
rect 46434 32998 46500 33032
rect 46534 32998 46600 33032
rect 46634 32998 46700 33032
rect 46734 32998 46821 33032
rect 46127 32990 46821 32998
rect 46127 32956 46188 32990
rect 46222 32956 46278 32990
rect 46312 32956 46368 32990
rect 46402 32956 46458 32990
rect 46492 32956 46548 32990
rect 46582 32956 46638 32990
rect 46672 32956 46728 32990
rect 46762 32956 46821 32990
rect 46127 32932 46821 32956
rect 46127 32900 46200 32932
rect 46234 32900 46300 32932
rect 46334 32900 46400 32932
rect 46434 32900 46500 32932
rect 46127 32866 46188 32900
rect 46234 32898 46278 32900
rect 46334 32898 46368 32900
rect 46434 32898 46458 32900
rect 46222 32866 46278 32898
rect 46312 32866 46368 32898
rect 46402 32866 46458 32898
rect 46492 32898 46500 32900
rect 46534 32900 46600 32932
rect 46534 32898 46548 32900
rect 46492 32866 46548 32898
rect 46582 32898 46600 32900
rect 46634 32900 46700 32932
rect 46734 32900 46821 32932
rect 46634 32898 46638 32900
rect 46582 32866 46638 32898
rect 46672 32898 46700 32900
rect 46672 32866 46728 32898
rect 46762 32866 46821 32900
rect 46127 32832 46821 32866
rect 46127 32810 46200 32832
rect 46234 32810 46300 32832
rect 46334 32810 46400 32832
rect 46434 32810 46500 32832
rect 46127 32776 46188 32810
rect 46234 32798 46278 32810
rect 46334 32798 46368 32810
rect 46434 32798 46458 32810
rect 46222 32776 46278 32798
rect 46312 32776 46368 32798
rect 46402 32776 46458 32798
rect 46492 32798 46500 32810
rect 46534 32810 46600 32832
rect 46534 32798 46548 32810
rect 46492 32776 46548 32798
rect 46582 32798 46600 32810
rect 46634 32810 46700 32832
rect 46734 32810 46821 32832
rect 46634 32798 46638 32810
rect 46582 32776 46638 32798
rect 46672 32798 46700 32810
rect 46672 32776 46728 32798
rect 46762 32776 46821 32810
rect 46127 32732 46821 32776
rect 46127 32720 46200 32732
rect 46234 32720 46300 32732
rect 46334 32720 46400 32732
rect 46434 32720 46500 32732
rect 46127 32686 46188 32720
rect 46234 32698 46278 32720
rect 46334 32698 46368 32720
rect 46434 32698 46458 32720
rect 46222 32686 46278 32698
rect 46312 32686 46368 32698
rect 46402 32686 46458 32698
rect 46492 32698 46500 32720
rect 46534 32720 46600 32732
rect 46534 32698 46548 32720
rect 46492 32686 46548 32698
rect 46582 32698 46600 32720
rect 46634 32720 46700 32732
rect 46734 32720 46821 32732
rect 46634 32698 46638 32720
rect 46582 32686 46638 32698
rect 46672 32698 46700 32720
rect 46672 32686 46728 32698
rect 46762 32686 46821 32720
rect 46127 32625 46821 32686
rect 46883 33268 46955 33324
rect 46883 33234 46902 33268
rect 46936 33234 46955 33268
rect 46883 33178 46955 33234
rect 46883 33144 46902 33178
rect 46936 33144 46955 33178
rect 46883 33088 46955 33144
rect 46883 33054 46902 33088
rect 46936 33054 46955 33088
rect 46883 32998 46955 33054
rect 46883 32964 46902 32998
rect 46936 32964 46955 32998
rect 46883 32908 46955 32964
rect 46883 32874 46902 32908
rect 46936 32874 46955 32908
rect 46883 32818 46955 32874
rect 46883 32784 46902 32818
rect 46936 32784 46955 32818
rect 46883 32728 46955 32784
rect 46883 32694 46902 32728
rect 46936 32694 46955 32728
rect 46883 32638 46955 32694
rect 45993 32563 46065 32623
rect 46883 32604 46902 32638
rect 46936 32604 46955 32638
rect 46883 32563 46955 32604
rect 45993 32544 46955 32563
rect 45993 32510 46090 32544
rect 46124 32510 46180 32544
rect 46214 32510 46270 32544
rect 46304 32510 46360 32544
rect 46394 32510 46450 32544
rect 46484 32510 46540 32544
rect 46574 32510 46630 32544
rect 46664 32510 46720 32544
rect 46754 32510 46810 32544
rect 46844 32510 46955 32544
rect 45993 32491 46955 32510
rect 47019 33434 47051 33468
rect 47085 33434 47204 33468
rect 47238 33434 47269 33468
rect 48359 33468 48609 33517
rect 47019 33378 47269 33434
rect 47019 33344 47051 33378
rect 47085 33344 47204 33378
rect 47238 33344 47269 33378
rect 47019 33288 47269 33344
rect 47019 33254 47051 33288
rect 47085 33254 47204 33288
rect 47238 33254 47269 33288
rect 47019 33198 47269 33254
rect 47019 33164 47051 33198
rect 47085 33164 47204 33198
rect 47238 33164 47269 33198
rect 47019 33108 47269 33164
rect 47019 33074 47051 33108
rect 47085 33074 47204 33108
rect 47238 33074 47269 33108
rect 47019 33018 47269 33074
rect 47019 32984 47051 33018
rect 47085 32984 47204 33018
rect 47238 32984 47269 33018
rect 47019 32928 47269 32984
rect 47019 32894 47051 32928
rect 47085 32894 47204 32928
rect 47238 32894 47269 32928
rect 47019 32838 47269 32894
rect 47019 32804 47051 32838
rect 47085 32804 47204 32838
rect 47238 32804 47269 32838
rect 47019 32748 47269 32804
rect 47019 32714 47051 32748
rect 47085 32714 47204 32748
rect 47238 32714 47269 32748
rect 47019 32658 47269 32714
rect 47019 32624 47051 32658
rect 47085 32624 47204 32658
rect 47238 32624 47269 32658
rect 47019 32568 47269 32624
rect 47019 32534 47051 32568
rect 47085 32534 47204 32568
rect 47238 32534 47269 32568
rect 45679 32444 45711 32478
rect 45745 32444 45864 32478
rect 45898 32444 45929 32478
rect 45679 32427 45929 32444
rect 47019 32478 47269 32534
rect 47333 33436 48295 33453
rect 47333 33402 47354 33436
rect 47388 33402 47444 33436
rect 47478 33434 47534 33436
rect 47568 33434 47624 33436
rect 47658 33434 47714 33436
rect 47748 33434 47804 33436
rect 47838 33434 47894 33436
rect 47928 33434 47984 33436
rect 48018 33434 48074 33436
rect 48108 33434 48164 33436
rect 48198 33434 48254 33436
rect 47498 33402 47534 33434
rect 47588 33402 47624 33434
rect 47678 33402 47714 33434
rect 47768 33402 47804 33434
rect 47858 33402 47894 33434
rect 47948 33402 47984 33434
rect 48038 33402 48074 33434
rect 48128 33402 48164 33434
rect 48218 33402 48254 33434
rect 48288 33402 48295 33436
rect 47333 33400 47464 33402
rect 47498 33400 47554 33402
rect 47588 33400 47644 33402
rect 47678 33400 47734 33402
rect 47768 33400 47824 33402
rect 47858 33400 47914 33402
rect 47948 33400 48004 33402
rect 48038 33400 48094 33402
rect 48128 33400 48184 33402
rect 48218 33400 48295 33402
rect 47333 33381 48295 33400
rect 47333 33377 47405 33381
rect 47333 33343 47352 33377
rect 47386 33343 47405 33377
rect 47333 33287 47405 33343
rect 48223 33358 48295 33381
rect 48223 33324 48242 33358
rect 48276 33324 48295 33358
rect 47333 33253 47352 33287
rect 47386 33253 47405 33287
rect 47333 33197 47405 33253
rect 47333 33163 47352 33197
rect 47386 33163 47405 33197
rect 47333 33107 47405 33163
rect 47333 33073 47352 33107
rect 47386 33073 47405 33107
rect 47333 33017 47405 33073
rect 47333 32983 47352 33017
rect 47386 32983 47405 33017
rect 47333 32927 47405 32983
rect 47333 32893 47352 32927
rect 47386 32893 47405 32927
rect 47333 32837 47405 32893
rect 47333 32803 47352 32837
rect 47386 32803 47405 32837
rect 47333 32747 47405 32803
rect 47333 32713 47352 32747
rect 47386 32713 47405 32747
rect 47333 32657 47405 32713
rect 47333 32623 47352 32657
rect 47386 32623 47405 32657
rect 47467 33260 48161 33319
rect 47467 33226 47528 33260
rect 47562 33232 47618 33260
rect 47652 33232 47708 33260
rect 47742 33232 47798 33260
rect 47574 33226 47618 33232
rect 47674 33226 47708 33232
rect 47774 33226 47798 33232
rect 47832 33232 47888 33260
rect 47832 33226 47840 33232
rect 47467 33198 47540 33226
rect 47574 33198 47640 33226
rect 47674 33198 47740 33226
rect 47774 33198 47840 33226
rect 47874 33226 47888 33232
rect 47922 33232 47978 33260
rect 47922 33226 47940 33232
rect 47874 33198 47940 33226
rect 47974 33226 47978 33232
rect 48012 33232 48068 33260
rect 48012 33226 48040 33232
rect 48102 33226 48161 33260
rect 47974 33198 48040 33226
rect 48074 33198 48161 33226
rect 47467 33170 48161 33198
rect 47467 33136 47528 33170
rect 47562 33136 47618 33170
rect 47652 33136 47708 33170
rect 47742 33136 47798 33170
rect 47832 33136 47888 33170
rect 47922 33136 47978 33170
rect 48012 33136 48068 33170
rect 48102 33136 48161 33170
rect 47467 33132 48161 33136
rect 47467 33098 47540 33132
rect 47574 33098 47640 33132
rect 47674 33098 47740 33132
rect 47774 33098 47840 33132
rect 47874 33098 47940 33132
rect 47974 33098 48040 33132
rect 48074 33098 48161 33132
rect 47467 33080 48161 33098
rect 47467 33046 47528 33080
rect 47562 33046 47618 33080
rect 47652 33046 47708 33080
rect 47742 33046 47798 33080
rect 47832 33046 47888 33080
rect 47922 33046 47978 33080
rect 48012 33046 48068 33080
rect 48102 33046 48161 33080
rect 47467 33032 48161 33046
rect 47467 32998 47540 33032
rect 47574 32998 47640 33032
rect 47674 32998 47740 33032
rect 47774 32998 47840 33032
rect 47874 32998 47940 33032
rect 47974 32998 48040 33032
rect 48074 32998 48161 33032
rect 47467 32990 48161 32998
rect 47467 32956 47528 32990
rect 47562 32956 47618 32990
rect 47652 32956 47708 32990
rect 47742 32956 47798 32990
rect 47832 32956 47888 32990
rect 47922 32956 47978 32990
rect 48012 32956 48068 32990
rect 48102 32956 48161 32990
rect 47467 32932 48161 32956
rect 47467 32900 47540 32932
rect 47574 32900 47640 32932
rect 47674 32900 47740 32932
rect 47774 32900 47840 32932
rect 47467 32866 47528 32900
rect 47574 32898 47618 32900
rect 47674 32898 47708 32900
rect 47774 32898 47798 32900
rect 47562 32866 47618 32898
rect 47652 32866 47708 32898
rect 47742 32866 47798 32898
rect 47832 32898 47840 32900
rect 47874 32900 47940 32932
rect 47874 32898 47888 32900
rect 47832 32866 47888 32898
rect 47922 32898 47940 32900
rect 47974 32900 48040 32932
rect 48074 32900 48161 32932
rect 47974 32898 47978 32900
rect 47922 32866 47978 32898
rect 48012 32898 48040 32900
rect 48012 32866 48068 32898
rect 48102 32866 48161 32900
rect 47467 32832 48161 32866
rect 47467 32810 47540 32832
rect 47574 32810 47640 32832
rect 47674 32810 47740 32832
rect 47774 32810 47840 32832
rect 47467 32776 47528 32810
rect 47574 32798 47618 32810
rect 47674 32798 47708 32810
rect 47774 32798 47798 32810
rect 47562 32776 47618 32798
rect 47652 32776 47708 32798
rect 47742 32776 47798 32798
rect 47832 32798 47840 32810
rect 47874 32810 47940 32832
rect 47874 32798 47888 32810
rect 47832 32776 47888 32798
rect 47922 32798 47940 32810
rect 47974 32810 48040 32832
rect 48074 32810 48161 32832
rect 47974 32798 47978 32810
rect 47922 32776 47978 32798
rect 48012 32798 48040 32810
rect 48012 32776 48068 32798
rect 48102 32776 48161 32810
rect 47467 32732 48161 32776
rect 47467 32720 47540 32732
rect 47574 32720 47640 32732
rect 47674 32720 47740 32732
rect 47774 32720 47840 32732
rect 47467 32686 47528 32720
rect 47574 32698 47618 32720
rect 47674 32698 47708 32720
rect 47774 32698 47798 32720
rect 47562 32686 47618 32698
rect 47652 32686 47708 32698
rect 47742 32686 47798 32698
rect 47832 32698 47840 32720
rect 47874 32720 47940 32732
rect 47874 32698 47888 32720
rect 47832 32686 47888 32698
rect 47922 32698 47940 32720
rect 47974 32720 48040 32732
rect 48074 32720 48161 32732
rect 47974 32698 47978 32720
rect 47922 32686 47978 32698
rect 48012 32698 48040 32720
rect 48012 32686 48068 32698
rect 48102 32686 48161 32720
rect 47467 32625 48161 32686
rect 48223 33268 48295 33324
rect 48223 33234 48242 33268
rect 48276 33234 48295 33268
rect 48223 33178 48295 33234
rect 48223 33144 48242 33178
rect 48276 33144 48295 33178
rect 48223 33088 48295 33144
rect 48223 33054 48242 33088
rect 48276 33054 48295 33088
rect 48223 32998 48295 33054
rect 48223 32964 48242 32998
rect 48276 32964 48295 32998
rect 48223 32908 48295 32964
rect 48223 32874 48242 32908
rect 48276 32874 48295 32908
rect 48223 32818 48295 32874
rect 48223 32784 48242 32818
rect 48276 32784 48295 32818
rect 48223 32728 48295 32784
rect 48223 32694 48242 32728
rect 48276 32694 48295 32728
rect 48223 32638 48295 32694
rect 47333 32563 47405 32623
rect 48223 32604 48242 32638
rect 48276 32604 48295 32638
rect 48223 32563 48295 32604
rect 47333 32544 48295 32563
rect 47333 32510 47430 32544
rect 47464 32510 47520 32544
rect 47554 32510 47610 32544
rect 47644 32510 47700 32544
rect 47734 32510 47790 32544
rect 47824 32510 47880 32544
rect 47914 32510 47970 32544
rect 48004 32510 48060 32544
rect 48094 32510 48150 32544
rect 48184 32510 48295 32544
rect 47333 32491 48295 32510
rect 48359 33434 48391 33468
rect 48425 33434 48544 33468
rect 48578 33434 48609 33468
rect 49699 33468 49949 33517
rect 48359 33378 48609 33434
rect 48359 33344 48391 33378
rect 48425 33344 48544 33378
rect 48578 33344 48609 33378
rect 48359 33288 48609 33344
rect 48359 33254 48391 33288
rect 48425 33254 48544 33288
rect 48578 33254 48609 33288
rect 48359 33198 48609 33254
rect 48359 33164 48391 33198
rect 48425 33164 48544 33198
rect 48578 33164 48609 33198
rect 48359 33108 48609 33164
rect 48359 33074 48391 33108
rect 48425 33074 48544 33108
rect 48578 33074 48609 33108
rect 48359 33018 48609 33074
rect 48359 32984 48391 33018
rect 48425 32984 48544 33018
rect 48578 32984 48609 33018
rect 48359 32928 48609 32984
rect 48359 32894 48391 32928
rect 48425 32894 48544 32928
rect 48578 32894 48609 32928
rect 48359 32838 48609 32894
rect 48359 32804 48391 32838
rect 48425 32804 48544 32838
rect 48578 32804 48609 32838
rect 48359 32748 48609 32804
rect 48359 32714 48391 32748
rect 48425 32714 48544 32748
rect 48578 32714 48609 32748
rect 48359 32658 48609 32714
rect 48359 32624 48391 32658
rect 48425 32624 48544 32658
rect 48578 32624 48609 32658
rect 48359 32568 48609 32624
rect 48359 32534 48391 32568
rect 48425 32534 48544 32568
rect 48578 32534 48609 32568
rect 47019 32444 47051 32478
rect 47085 32444 47204 32478
rect 47238 32444 47269 32478
rect 47019 32427 47269 32444
rect 48359 32478 48609 32534
rect 48673 33436 49635 33453
rect 48673 33402 48694 33436
rect 48728 33402 48784 33436
rect 48818 33434 48874 33436
rect 48908 33434 48964 33436
rect 48998 33434 49054 33436
rect 49088 33434 49144 33436
rect 49178 33434 49234 33436
rect 49268 33434 49324 33436
rect 49358 33434 49414 33436
rect 49448 33434 49504 33436
rect 49538 33434 49594 33436
rect 48838 33402 48874 33434
rect 48928 33402 48964 33434
rect 49018 33402 49054 33434
rect 49108 33402 49144 33434
rect 49198 33402 49234 33434
rect 49288 33402 49324 33434
rect 49378 33402 49414 33434
rect 49468 33402 49504 33434
rect 49558 33402 49594 33434
rect 49628 33402 49635 33436
rect 48673 33400 48804 33402
rect 48838 33400 48894 33402
rect 48928 33400 48984 33402
rect 49018 33400 49074 33402
rect 49108 33400 49164 33402
rect 49198 33400 49254 33402
rect 49288 33400 49344 33402
rect 49378 33400 49434 33402
rect 49468 33400 49524 33402
rect 49558 33400 49635 33402
rect 48673 33381 49635 33400
rect 48673 33377 48745 33381
rect 48673 33343 48692 33377
rect 48726 33343 48745 33377
rect 48673 33287 48745 33343
rect 49563 33358 49635 33381
rect 49563 33324 49582 33358
rect 49616 33324 49635 33358
rect 48673 33253 48692 33287
rect 48726 33253 48745 33287
rect 48673 33197 48745 33253
rect 48673 33163 48692 33197
rect 48726 33163 48745 33197
rect 48673 33107 48745 33163
rect 48673 33073 48692 33107
rect 48726 33073 48745 33107
rect 48673 33017 48745 33073
rect 48673 32983 48692 33017
rect 48726 32983 48745 33017
rect 48673 32927 48745 32983
rect 48673 32893 48692 32927
rect 48726 32893 48745 32927
rect 48673 32837 48745 32893
rect 48673 32803 48692 32837
rect 48726 32803 48745 32837
rect 48673 32747 48745 32803
rect 48673 32713 48692 32747
rect 48726 32713 48745 32747
rect 48673 32657 48745 32713
rect 48673 32623 48692 32657
rect 48726 32623 48745 32657
rect 48807 33260 49501 33319
rect 48807 33226 48868 33260
rect 48902 33232 48958 33260
rect 48992 33232 49048 33260
rect 49082 33232 49138 33260
rect 48914 33226 48958 33232
rect 49014 33226 49048 33232
rect 49114 33226 49138 33232
rect 49172 33232 49228 33260
rect 49172 33226 49180 33232
rect 48807 33198 48880 33226
rect 48914 33198 48980 33226
rect 49014 33198 49080 33226
rect 49114 33198 49180 33226
rect 49214 33226 49228 33232
rect 49262 33232 49318 33260
rect 49262 33226 49280 33232
rect 49214 33198 49280 33226
rect 49314 33226 49318 33232
rect 49352 33232 49408 33260
rect 49352 33226 49380 33232
rect 49442 33226 49501 33260
rect 49314 33198 49380 33226
rect 49414 33198 49501 33226
rect 48807 33170 49501 33198
rect 48807 33136 48868 33170
rect 48902 33136 48958 33170
rect 48992 33136 49048 33170
rect 49082 33136 49138 33170
rect 49172 33136 49228 33170
rect 49262 33136 49318 33170
rect 49352 33136 49408 33170
rect 49442 33136 49501 33170
rect 48807 33132 49501 33136
rect 48807 33098 48880 33132
rect 48914 33098 48980 33132
rect 49014 33098 49080 33132
rect 49114 33098 49180 33132
rect 49214 33098 49280 33132
rect 49314 33098 49380 33132
rect 49414 33098 49501 33132
rect 48807 33080 49501 33098
rect 48807 33046 48868 33080
rect 48902 33046 48958 33080
rect 48992 33046 49048 33080
rect 49082 33046 49138 33080
rect 49172 33046 49228 33080
rect 49262 33046 49318 33080
rect 49352 33046 49408 33080
rect 49442 33046 49501 33080
rect 48807 33032 49501 33046
rect 48807 32998 48880 33032
rect 48914 32998 48980 33032
rect 49014 32998 49080 33032
rect 49114 32998 49180 33032
rect 49214 32998 49280 33032
rect 49314 32998 49380 33032
rect 49414 32998 49501 33032
rect 48807 32990 49501 32998
rect 48807 32956 48868 32990
rect 48902 32956 48958 32990
rect 48992 32956 49048 32990
rect 49082 32956 49138 32990
rect 49172 32956 49228 32990
rect 49262 32956 49318 32990
rect 49352 32956 49408 32990
rect 49442 32956 49501 32990
rect 48807 32932 49501 32956
rect 48807 32900 48880 32932
rect 48914 32900 48980 32932
rect 49014 32900 49080 32932
rect 49114 32900 49180 32932
rect 48807 32866 48868 32900
rect 48914 32898 48958 32900
rect 49014 32898 49048 32900
rect 49114 32898 49138 32900
rect 48902 32866 48958 32898
rect 48992 32866 49048 32898
rect 49082 32866 49138 32898
rect 49172 32898 49180 32900
rect 49214 32900 49280 32932
rect 49214 32898 49228 32900
rect 49172 32866 49228 32898
rect 49262 32898 49280 32900
rect 49314 32900 49380 32932
rect 49414 32900 49501 32932
rect 49314 32898 49318 32900
rect 49262 32866 49318 32898
rect 49352 32898 49380 32900
rect 49352 32866 49408 32898
rect 49442 32866 49501 32900
rect 48807 32832 49501 32866
rect 48807 32810 48880 32832
rect 48914 32810 48980 32832
rect 49014 32810 49080 32832
rect 49114 32810 49180 32832
rect 48807 32776 48868 32810
rect 48914 32798 48958 32810
rect 49014 32798 49048 32810
rect 49114 32798 49138 32810
rect 48902 32776 48958 32798
rect 48992 32776 49048 32798
rect 49082 32776 49138 32798
rect 49172 32798 49180 32810
rect 49214 32810 49280 32832
rect 49214 32798 49228 32810
rect 49172 32776 49228 32798
rect 49262 32798 49280 32810
rect 49314 32810 49380 32832
rect 49414 32810 49501 32832
rect 49314 32798 49318 32810
rect 49262 32776 49318 32798
rect 49352 32798 49380 32810
rect 49352 32776 49408 32798
rect 49442 32776 49501 32810
rect 48807 32732 49501 32776
rect 48807 32720 48880 32732
rect 48914 32720 48980 32732
rect 49014 32720 49080 32732
rect 49114 32720 49180 32732
rect 48807 32686 48868 32720
rect 48914 32698 48958 32720
rect 49014 32698 49048 32720
rect 49114 32698 49138 32720
rect 48902 32686 48958 32698
rect 48992 32686 49048 32698
rect 49082 32686 49138 32698
rect 49172 32698 49180 32720
rect 49214 32720 49280 32732
rect 49214 32698 49228 32720
rect 49172 32686 49228 32698
rect 49262 32698 49280 32720
rect 49314 32720 49380 32732
rect 49414 32720 49501 32732
rect 49314 32698 49318 32720
rect 49262 32686 49318 32698
rect 49352 32698 49380 32720
rect 49352 32686 49408 32698
rect 49442 32686 49501 32720
rect 48807 32625 49501 32686
rect 49563 33268 49635 33324
rect 49563 33234 49582 33268
rect 49616 33234 49635 33268
rect 49563 33178 49635 33234
rect 49563 33144 49582 33178
rect 49616 33144 49635 33178
rect 49563 33088 49635 33144
rect 49563 33054 49582 33088
rect 49616 33054 49635 33088
rect 49563 32998 49635 33054
rect 49563 32964 49582 32998
rect 49616 32964 49635 32998
rect 49563 32908 49635 32964
rect 49563 32874 49582 32908
rect 49616 32874 49635 32908
rect 49563 32818 49635 32874
rect 49563 32784 49582 32818
rect 49616 32784 49635 32818
rect 49563 32728 49635 32784
rect 49563 32694 49582 32728
rect 49616 32694 49635 32728
rect 49563 32638 49635 32694
rect 48673 32563 48745 32623
rect 49563 32604 49582 32638
rect 49616 32604 49635 32638
rect 49563 32563 49635 32604
rect 48673 32544 49635 32563
rect 48673 32510 48770 32544
rect 48804 32510 48860 32544
rect 48894 32510 48950 32544
rect 48984 32510 49040 32544
rect 49074 32510 49130 32544
rect 49164 32510 49220 32544
rect 49254 32510 49310 32544
rect 49344 32510 49400 32544
rect 49434 32510 49490 32544
rect 49524 32510 49635 32544
rect 48673 32491 49635 32510
rect 49699 33434 49731 33468
rect 49765 33434 49884 33468
rect 49918 33434 49949 33468
rect 51039 33468 51289 33517
rect 49699 33378 49949 33434
rect 49699 33344 49731 33378
rect 49765 33344 49884 33378
rect 49918 33344 49949 33378
rect 49699 33288 49949 33344
rect 49699 33254 49731 33288
rect 49765 33254 49884 33288
rect 49918 33254 49949 33288
rect 49699 33198 49949 33254
rect 49699 33164 49731 33198
rect 49765 33164 49884 33198
rect 49918 33164 49949 33198
rect 49699 33108 49949 33164
rect 49699 33074 49731 33108
rect 49765 33074 49884 33108
rect 49918 33074 49949 33108
rect 49699 33018 49949 33074
rect 49699 32984 49731 33018
rect 49765 32984 49884 33018
rect 49918 32984 49949 33018
rect 49699 32928 49949 32984
rect 49699 32894 49731 32928
rect 49765 32894 49884 32928
rect 49918 32894 49949 32928
rect 49699 32838 49949 32894
rect 49699 32804 49731 32838
rect 49765 32804 49884 32838
rect 49918 32804 49949 32838
rect 49699 32748 49949 32804
rect 49699 32714 49731 32748
rect 49765 32714 49884 32748
rect 49918 32714 49949 32748
rect 49699 32658 49949 32714
rect 49699 32624 49731 32658
rect 49765 32624 49884 32658
rect 49918 32624 49949 32658
rect 49699 32568 49949 32624
rect 49699 32534 49731 32568
rect 49765 32534 49884 32568
rect 49918 32534 49949 32568
rect 48359 32444 48391 32478
rect 48425 32444 48544 32478
rect 48578 32444 48609 32478
rect 48359 32427 48609 32444
rect 49699 32478 49949 32534
rect 50013 33436 50975 33453
rect 50013 33402 50034 33436
rect 50068 33402 50124 33436
rect 50158 33434 50214 33436
rect 50248 33434 50304 33436
rect 50338 33434 50394 33436
rect 50428 33434 50484 33436
rect 50518 33434 50574 33436
rect 50608 33434 50664 33436
rect 50698 33434 50754 33436
rect 50788 33434 50844 33436
rect 50878 33434 50934 33436
rect 50178 33402 50214 33434
rect 50268 33402 50304 33434
rect 50358 33402 50394 33434
rect 50448 33402 50484 33434
rect 50538 33402 50574 33434
rect 50628 33402 50664 33434
rect 50718 33402 50754 33434
rect 50808 33402 50844 33434
rect 50898 33402 50934 33434
rect 50968 33402 50975 33436
rect 50013 33400 50144 33402
rect 50178 33400 50234 33402
rect 50268 33400 50324 33402
rect 50358 33400 50414 33402
rect 50448 33400 50504 33402
rect 50538 33400 50594 33402
rect 50628 33400 50684 33402
rect 50718 33400 50774 33402
rect 50808 33400 50864 33402
rect 50898 33400 50975 33402
rect 50013 33381 50975 33400
rect 50013 33377 50085 33381
rect 50013 33343 50032 33377
rect 50066 33343 50085 33377
rect 50013 33287 50085 33343
rect 50903 33358 50975 33381
rect 50903 33324 50922 33358
rect 50956 33324 50975 33358
rect 50013 33253 50032 33287
rect 50066 33253 50085 33287
rect 50013 33197 50085 33253
rect 50013 33163 50032 33197
rect 50066 33163 50085 33197
rect 50013 33107 50085 33163
rect 50013 33073 50032 33107
rect 50066 33073 50085 33107
rect 50013 33017 50085 33073
rect 50013 32983 50032 33017
rect 50066 32983 50085 33017
rect 50013 32927 50085 32983
rect 50013 32893 50032 32927
rect 50066 32893 50085 32927
rect 50013 32837 50085 32893
rect 50013 32803 50032 32837
rect 50066 32803 50085 32837
rect 50013 32747 50085 32803
rect 50013 32713 50032 32747
rect 50066 32713 50085 32747
rect 50013 32657 50085 32713
rect 50013 32623 50032 32657
rect 50066 32623 50085 32657
rect 50147 33260 50841 33319
rect 50147 33226 50208 33260
rect 50242 33232 50298 33260
rect 50332 33232 50388 33260
rect 50422 33232 50478 33260
rect 50254 33226 50298 33232
rect 50354 33226 50388 33232
rect 50454 33226 50478 33232
rect 50512 33232 50568 33260
rect 50512 33226 50520 33232
rect 50147 33198 50220 33226
rect 50254 33198 50320 33226
rect 50354 33198 50420 33226
rect 50454 33198 50520 33226
rect 50554 33226 50568 33232
rect 50602 33232 50658 33260
rect 50602 33226 50620 33232
rect 50554 33198 50620 33226
rect 50654 33226 50658 33232
rect 50692 33232 50748 33260
rect 50692 33226 50720 33232
rect 50782 33226 50841 33260
rect 50654 33198 50720 33226
rect 50754 33198 50841 33226
rect 50147 33170 50841 33198
rect 50147 33136 50208 33170
rect 50242 33136 50298 33170
rect 50332 33136 50388 33170
rect 50422 33136 50478 33170
rect 50512 33136 50568 33170
rect 50602 33136 50658 33170
rect 50692 33136 50748 33170
rect 50782 33136 50841 33170
rect 50147 33132 50841 33136
rect 50147 33098 50220 33132
rect 50254 33098 50320 33132
rect 50354 33098 50420 33132
rect 50454 33098 50520 33132
rect 50554 33098 50620 33132
rect 50654 33098 50720 33132
rect 50754 33098 50841 33132
rect 50147 33080 50841 33098
rect 50147 33046 50208 33080
rect 50242 33046 50298 33080
rect 50332 33046 50388 33080
rect 50422 33046 50478 33080
rect 50512 33046 50568 33080
rect 50602 33046 50658 33080
rect 50692 33046 50748 33080
rect 50782 33046 50841 33080
rect 50147 33032 50841 33046
rect 50147 32998 50220 33032
rect 50254 32998 50320 33032
rect 50354 32998 50420 33032
rect 50454 32998 50520 33032
rect 50554 32998 50620 33032
rect 50654 32998 50720 33032
rect 50754 32998 50841 33032
rect 50147 32990 50841 32998
rect 50147 32956 50208 32990
rect 50242 32956 50298 32990
rect 50332 32956 50388 32990
rect 50422 32956 50478 32990
rect 50512 32956 50568 32990
rect 50602 32956 50658 32990
rect 50692 32956 50748 32990
rect 50782 32956 50841 32990
rect 50147 32932 50841 32956
rect 50147 32900 50220 32932
rect 50254 32900 50320 32932
rect 50354 32900 50420 32932
rect 50454 32900 50520 32932
rect 50147 32866 50208 32900
rect 50254 32898 50298 32900
rect 50354 32898 50388 32900
rect 50454 32898 50478 32900
rect 50242 32866 50298 32898
rect 50332 32866 50388 32898
rect 50422 32866 50478 32898
rect 50512 32898 50520 32900
rect 50554 32900 50620 32932
rect 50554 32898 50568 32900
rect 50512 32866 50568 32898
rect 50602 32898 50620 32900
rect 50654 32900 50720 32932
rect 50754 32900 50841 32932
rect 50654 32898 50658 32900
rect 50602 32866 50658 32898
rect 50692 32898 50720 32900
rect 50692 32866 50748 32898
rect 50782 32866 50841 32900
rect 50147 32832 50841 32866
rect 50147 32810 50220 32832
rect 50254 32810 50320 32832
rect 50354 32810 50420 32832
rect 50454 32810 50520 32832
rect 50147 32776 50208 32810
rect 50254 32798 50298 32810
rect 50354 32798 50388 32810
rect 50454 32798 50478 32810
rect 50242 32776 50298 32798
rect 50332 32776 50388 32798
rect 50422 32776 50478 32798
rect 50512 32798 50520 32810
rect 50554 32810 50620 32832
rect 50554 32798 50568 32810
rect 50512 32776 50568 32798
rect 50602 32798 50620 32810
rect 50654 32810 50720 32832
rect 50754 32810 50841 32832
rect 50654 32798 50658 32810
rect 50602 32776 50658 32798
rect 50692 32798 50720 32810
rect 50692 32776 50748 32798
rect 50782 32776 50841 32810
rect 50147 32732 50841 32776
rect 50147 32720 50220 32732
rect 50254 32720 50320 32732
rect 50354 32720 50420 32732
rect 50454 32720 50520 32732
rect 50147 32686 50208 32720
rect 50254 32698 50298 32720
rect 50354 32698 50388 32720
rect 50454 32698 50478 32720
rect 50242 32686 50298 32698
rect 50332 32686 50388 32698
rect 50422 32686 50478 32698
rect 50512 32698 50520 32720
rect 50554 32720 50620 32732
rect 50554 32698 50568 32720
rect 50512 32686 50568 32698
rect 50602 32698 50620 32720
rect 50654 32720 50720 32732
rect 50754 32720 50841 32732
rect 50654 32698 50658 32720
rect 50602 32686 50658 32698
rect 50692 32698 50720 32720
rect 50692 32686 50748 32698
rect 50782 32686 50841 32720
rect 50147 32625 50841 32686
rect 50903 33268 50975 33324
rect 50903 33234 50922 33268
rect 50956 33234 50975 33268
rect 50903 33178 50975 33234
rect 50903 33144 50922 33178
rect 50956 33144 50975 33178
rect 50903 33088 50975 33144
rect 50903 33054 50922 33088
rect 50956 33054 50975 33088
rect 50903 32998 50975 33054
rect 50903 32964 50922 32998
rect 50956 32964 50975 32998
rect 50903 32908 50975 32964
rect 50903 32874 50922 32908
rect 50956 32874 50975 32908
rect 50903 32818 50975 32874
rect 50903 32784 50922 32818
rect 50956 32784 50975 32818
rect 50903 32728 50975 32784
rect 50903 32694 50922 32728
rect 50956 32694 50975 32728
rect 50903 32638 50975 32694
rect 50013 32563 50085 32623
rect 50903 32604 50922 32638
rect 50956 32604 50975 32638
rect 50903 32563 50975 32604
rect 50013 32544 50975 32563
rect 50013 32510 50110 32544
rect 50144 32510 50200 32544
rect 50234 32510 50290 32544
rect 50324 32510 50380 32544
rect 50414 32510 50470 32544
rect 50504 32510 50560 32544
rect 50594 32510 50650 32544
rect 50684 32510 50740 32544
rect 50774 32510 50830 32544
rect 50864 32510 50975 32544
rect 50013 32491 50975 32510
rect 51039 33434 51071 33468
rect 51105 33434 51224 33468
rect 51258 33434 51289 33468
rect 52379 33468 52478 33517
rect 51039 33378 51289 33434
rect 51039 33344 51071 33378
rect 51105 33344 51224 33378
rect 51258 33344 51289 33378
rect 51039 33288 51289 33344
rect 51039 33254 51071 33288
rect 51105 33254 51224 33288
rect 51258 33254 51289 33288
rect 51039 33198 51289 33254
rect 51039 33164 51071 33198
rect 51105 33164 51224 33198
rect 51258 33164 51289 33198
rect 51039 33108 51289 33164
rect 51039 33074 51071 33108
rect 51105 33074 51224 33108
rect 51258 33074 51289 33108
rect 51039 33018 51289 33074
rect 51039 32984 51071 33018
rect 51105 32984 51224 33018
rect 51258 32984 51289 33018
rect 51039 32928 51289 32984
rect 51039 32894 51071 32928
rect 51105 32894 51224 32928
rect 51258 32894 51289 32928
rect 51039 32838 51289 32894
rect 51039 32804 51071 32838
rect 51105 32804 51224 32838
rect 51258 32804 51289 32838
rect 51039 32748 51289 32804
rect 51039 32714 51071 32748
rect 51105 32714 51224 32748
rect 51258 32714 51289 32748
rect 51039 32658 51289 32714
rect 51039 32624 51071 32658
rect 51105 32624 51224 32658
rect 51258 32624 51289 32658
rect 51039 32568 51289 32624
rect 51039 32534 51071 32568
rect 51105 32534 51224 32568
rect 51258 32534 51289 32568
rect 49699 32444 49731 32478
rect 49765 32444 49884 32478
rect 49918 32444 49949 32478
rect 49699 32427 49949 32444
rect 51039 32478 51289 32534
rect 51353 33436 52315 33453
rect 51353 33402 51374 33436
rect 51408 33402 51464 33436
rect 51498 33434 51554 33436
rect 51588 33434 51644 33436
rect 51678 33434 51734 33436
rect 51768 33434 51824 33436
rect 51858 33434 51914 33436
rect 51948 33434 52004 33436
rect 52038 33434 52094 33436
rect 52128 33434 52184 33436
rect 52218 33434 52274 33436
rect 51518 33402 51554 33434
rect 51608 33402 51644 33434
rect 51698 33402 51734 33434
rect 51788 33402 51824 33434
rect 51878 33402 51914 33434
rect 51968 33402 52004 33434
rect 52058 33402 52094 33434
rect 52148 33402 52184 33434
rect 52238 33402 52274 33434
rect 52308 33402 52315 33436
rect 51353 33400 51484 33402
rect 51518 33400 51574 33402
rect 51608 33400 51664 33402
rect 51698 33400 51754 33402
rect 51788 33400 51844 33402
rect 51878 33400 51934 33402
rect 51968 33400 52024 33402
rect 52058 33400 52114 33402
rect 52148 33400 52204 33402
rect 52238 33400 52315 33402
rect 51353 33381 52315 33400
rect 51353 33377 51425 33381
rect 51353 33343 51372 33377
rect 51406 33343 51425 33377
rect 51353 33287 51425 33343
rect 52243 33358 52315 33381
rect 52243 33324 52262 33358
rect 52296 33324 52315 33358
rect 51353 33253 51372 33287
rect 51406 33253 51425 33287
rect 51353 33197 51425 33253
rect 51353 33163 51372 33197
rect 51406 33163 51425 33197
rect 51353 33107 51425 33163
rect 51353 33073 51372 33107
rect 51406 33073 51425 33107
rect 51353 33017 51425 33073
rect 51353 32983 51372 33017
rect 51406 32983 51425 33017
rect 51353 32927 51425 32983
rect 51353 32893 51372 32927
rect 51406 32893 51425 32927
rect 51353 32837 51425 32893
rect 51353 32803 51372 32837
rect 51406 32803 51425 32837
rect 51353 32747 51425 32803
rect 51353 32713 51372 32747
rect 51406 32713 51425 32747
rect 51353 32657 51425 32713
rect 51353 32623 51372 32657
rect 51406 32623 51425 32657
rect 51487 33260 52181 33319
rect 51487 33226 51548 33260
rect 51582 33232 51638 33260
rect 51672 33232 51728 33260
rect 51762 33232 51818 33260
rect 51594 33226 51638 33232
rect 51694 33226 51728 33232
rect 51794 33226 51818 33232
rect 51852 33232 51908 33260
rect 51852 33226 51860 33232
rect 51487 33198 51560 33226
rect 51594 33198 51660 33226
rect 51694 33198 51760 33226
rect 51794 33198 51860 33226
rect 51894 33226 51908 33232
rect 51942 33232 51998 33260
rect 51942 33226 51960 33232
rect 51894 33198 51960 33226
rect 51994 33226 51998 33232
rect 52032 33232 52088 33260
rect 52032 33226 52060 33232
rect 52122 33226 52181 33260
rect 51994 33198 52060 33226
rect 52094 33198 52181 33226
rect 51487 33170 52181 33198
rect 51487 33136 51548 33170
rect 51582 33136 51638 33170
rect 51672 33136 51728 33170
rect 51762 33136 51818 33170
rect 51852 33136 51908 33170
rect 51942 33136 51998 33170
rect 52032 33136 52088 33170
rect 52122 33136 52181 33170
rect 51487 33132 52181 33136
rect 51487 33098 51560 33132
rect 51594 33098 51660 33132
rect 51694 33098 51760 33132
rect 51794 33098 51860 33132
rect 51894 33098 51960 33132
rect 51994 33098 52060 33132
rect 52094 33098 52181 33132
rect 51487 33080 52181 33098
rect 51487 33046 51548 33080
rect 51582 33046 51638 33080
rect 51672 33046 51728 33080
rect 51762 33046 51818 33080
rect 51852 33046 51908 33080
rect 51942 33046 51998 33080
rect 52032 33046 52088 33080
rect 52122 33046 52181 33080
rect 51487 33032 52181 33046
rect 51487 32998 51560 33032
rect 51594 32998 51660 33032
rect 51694 32998 51760 33032
rect 51794 32998 51860 33032
rect 51894 32998 51960 33032
rect 51994 32998 52060 33032
rect 52094 32998 52181 33032
rect 51487 32990 52181 32998
rect 51487 32956 51548 32990
rect 51582 32956 51638 32990
rect 51672 32956 51728 32990
rect 51762 32956 51818 32990
rect 51852 32956 51908 32990
rect 51942 32956 51998 32990
rect 52032 32956 52088 32990
rect 52122 32956 52181 32990
rect 51487 32932 52181 32956
rect 51487 32900 51560 32932
rect 51594 32900 51660 32932
rect 51694 32900 51760 32932
rect 51794 32900 51860 32932
rect 51487 32866 51548 32900
rect 51594 32898 51638 32900
rect 51694 32898 51728 32900
rect 51794 32898 51818 32900
rect 51582 32866 51638 32898
rect 51672 32866 51728 32898
rect 51762 32866 51818 32898
rect 51852 32898 51860 32900
rect 51894 32900 51960 32932
rect 51894 32898 51908 32900
rect 51852 32866 51908 32898
rect 51942 32898 51960 32900
rect 51994 32900 52060 32932
rect 52094 32900 52181 32932
rect 51994 32898 51998 32900
rect 51942 32866 51998 32898
rect 52032 32898 52060 32900
rect 52032 32866 52088 32898
rect 52122 32866 52181 32900
rect 51487 32832 52181 32866
rect 51487 32810 51560 32832
rect 51594 32810 51660 32832
rect 51694 32810 51760 32832
rect 51794 32810 51860 32832
rect 51487 32776 51548 32810
rect 51594 32798 51638 32810
rect 51694 32798 51728 32810
rect 51794 32798 51818 32810
rect 51582 32776 51638 32798
rect 51672 32776 51728 32798
rect 51762 32776 51818 32798
rect 51852 32798 51860 32810
rect 51894 32810 51960 32832
rect 51894 32798 51908 32810
rect 51852 32776 51908 32798
rect 51942 32798 51960 32810
rect 51994 32810 52060 32832
rect 52094 32810 52181 32832
rect 51994 32798 51998 32810
rect 51942 32776 51998 32798
rect 52032 32798 52060 32810
rect 52032 32776 52088 32798
rect 52122 32776 52181 32810
rect 51487 32732 52181 32776
rect 51487 32720 51560 32732
rect 51594 32720 51660 32732
rect 51694 32720 51760 32732
rect 51794 32720 51860 32732
rect 51487 32686 51548 32720
rect 51594 32698 51638 32720
rect 51694 32698 51728 32720
rect 51794 32698 51818 32720
rect 51582 32686 51638 32698
rect 51672 32686 51728 32698
rect 51762 32686 51818 32698
rect 51852 32698 51860 32720
rect 51894 32720 51960 32732
rect 51894 32698 51908 32720
rect 51852 32686 51908 32698
rect 51942 32698 51960 32720
rect 51994 32720 52060 32732
rect 52094 32720 52181 32732
rect 51994 32698 51998 32720
rect 51942 32686 51998 32698
rect 52032 32698 52060 32720
rect 52032 32686 52088 32698
rect 52122 32686 52181 32720
rect 51487 32625 52181 32686
rect 52243 33268 52315 33324
rect 52243 33234 52262 33268
rect 52296 33234 52315 33268
rect 52243 33178 52315 33234
rect 52243 33144 52262 33178
rect 52296 33144 52315 33178
rect 52243 33088 52315 33144
rect 52243 33054 52262 33088
rect 52296 33054 52315 33088
rect 52243 32998 52315 33054
rect 52243 32964 52262 32998
rect 52296 32964 52315 32998
rect 52243 32908 52315 32964
rect 52243 32874 52262 32908
rect 52296 32874 52315 32908
rect 52243 32818 52315 32874
rect 52243 32784 52262 32818
rect 52296 32784 52315 32818
rect 52243 32728 52315 32784
rect 52243 32694 52262 32728
rect 52296 32694 52315 32728
rect 52243 32638 52315 32694
rect 51353 32563 51425 32623
rect 52243 32604 52262 32638
rect 52296 32604 52315 32638
rect 52243 32563 52315 32604
rect 51353 32544 52315 32563
rect 51353 32510 51450 32544
rect 51484 32510 51540 32544
rect 51574 32510 51630 32544
rect 51664 32510 51720 32544
rect 51754 32510 51810 32544
rect 51844 32510 51900 32544
rect 51934 32510 51990 32544
rect 52024 32510 52080 32544
rect 52114 32510 52170 32544
rect 52204 32510 52315 32544
rect 51353 32491 52315 32510
rect 52379 33434 52411 33468
rect 52445 33434 52478 33468
rect 52379 33378 52478 33434
rect 52379 33344 52411 33378
rect 52445 33344 52478 33378
rect 52379 33288 52478 33344
rect 52379 33254 52411 33288
rect 52445 33254 52478 33288
rect 52379 33198 52478 33254
rect 52379 33164 52411 33198
rect 52445 33164 52478 33198
rect 52379 33108 52478 33164
rect 52379 33074 52411 33108
rect 52445 33074 52478 33108
rect 52379 33018 52478 33074
rect 52379 32984 52411 33018
rect 52445 32984 52478 33018
rect 52379 32928 52478 32984
rect 52379 32894 52411 32928
rect 52445 32894 52478 32928
rect 52379 32838 52478 32894
rect 52379 32804 52411 32838
rect 52445 32804 52478 32838
rect 52379 32748 52478 32804
rect 52379 32714 52411 32748
rect 52445 32714 52478 32748
rect 52379 32658 52478 32714
rect 52379 32624 52411 32658
rect 52445 32624 52478 32658
rect 52379 32568 52478 32624
rect 52379 32534 52411 32568
rect 52445 32534 52478 32568
rect 51039 32444 51071 32478
rect 51105 32444 51224 32478
rect 51258 32444 51289 32478
rect 51039 32427 51289 32444
rect 52379 32478 52478 32534
rect 52379 32444 52411 32478
rect 52445 32444 52478 32478
rect 52379 32427 52478 32444
rect 41810 32394 52478 32427
rect 41810 32360 41940 32394
rect 41974 32360 42030 32394
rect 42064 32360 42120 32394
rect 42154 32360 42210 32394
rect 42244 32360 42300 32394
rect 42334 32360 42390 32394
rect 42424 32360 42480 32394
rect 42514 32360 42570 32394
rect 42604 32360 42660 32394
rect 42694 32360 42750 32394
rect 42784 32360 42840 32394
rect 42874 32360 42930 32394
rect 42964 32360 43280 32394
rect 43314 32360 43370 32394
rect 43404 32360 43460 32394
rect 43494 32360 43550 32394
rect 43584 32360 43640 32394
rect 43674 32360 43730 32394
rect 43764 32360 43820 32394
rect 43854 32360 43910 32394
rect 43944 32360 44000 32394
rect 44034 32360 44090 32394
rect 44124 32360 44180 32394
rect 44214 32360 44270 32394
rect 44304 32360 44620 32394
rect 44654 32360 44710 32394
rect 44744 32360 44800 32394
rect 44834 32360 44890 32394
rect 44924 32360 44980 32394
rect 45014 32360 45070 32394
rect 45104 32360 45160 32394
rect 45194 32360 45250 32394
rect 45284 32360 45340 32394
rect 45374 32360 45430 32394
rect 45464 32360 45520 32394
rect 45554 32360 45610 32394
rect 45644 32360 45960 32394
rect 45994 32360 46050 32394
rect 46084 32360 46140 32394
rect 46174 32360 46230 32394
rect 46264 32360 46320 32394
rect 46354 32360 46410 32394
rect 46444 32360 46500 32394
rect 46534 32360 46590 32394
rect 46624 32360 46680 32394
rect 46714 32360 46770 32394
rect 46804 32360 46860 32394
rect 46894 32360 46950 32394
rect 46984 32360 47300 32394
rect 47334 32360 47390 32394
rect 47424 32360 47480 32394
rect 47514 32360 47570 32394
rect 47604 32360 47660 32394
rect 47694 32360 47750 32394
rect 47784 32360 47840 32394
rect 47874 32360 47930 32394
rect 47964 32360 48020 32394
rect 48054 32360 48110 32394
rect 48144 32360 48200 32394
rect 48234 32360 48290 32394
rect 48324 32360 48640 32394
rect 48674 32360 48730 32394
rect 48764 32360 48820 32394
rect 48854 32360 48910 32394
rect 48944 32360 49000 32394
rect 49034 32360 49090 32394
rect 49124 32360 49180 32394
rect 49214 32360 49270 32394
rect 49304 32360 49360 32394
rect 49394 32360 49450 32394
rect 49484 32360 49540 32394
rect 49574 32360 49630 32394
rect 49664 32360 49980 32394
rect 50014 32360 50070 32394
rect 50104 32360 50160 32394
rect 50194 32360 50250 32394
rect 50284 32360 50340 32394
rect 50374 32360 50430 32394
rect 50464 32360 50520 32394
rect 50554 32360 50610 32394
rect 50644 32360 50700 32394
rect 50734 32360 50790 32394
rect 50824 32360 50880 32394
rect 50914 32360 50970 32394
rect 51004 32360 51320 32394
rect 51354 32360 51410 32394
rect 51444 32360 51500 32394
rect 51534 32360 51590 32394
rect 51624 32360 51680 32394
rect 51714 32360 51770 32394
rect 51804 32360 51860 32394
rect 51894 32360 51950 32394
rect 51984 32360 52040 32394
rect 52074 32360 52130 32394
rect 52164 32360 52220 32394
rect 52254 32360 52310 32394
rect 52344 32360 52478 32394
rect 41810 32328 52478 32360
rect 19264 32049 21704 32062
rect 19264 32015 19447 32049
rect 19481 32015 19647 32049
rect 19681 32015 19847 32049
rect 19881 32015 20047 32049
rect 20081 32015 20247 32049
rect 20281 32015 20447 32049
rect 20481 32015 20647 32049
rect 20681 32015 20847 32049
rect 20881 32015 21047 32049
rect 21081 32015 21247 32049
rect 21281 32015 21447 32049
rect 21481 32015 21704 32049
rect 19264 32002 21704 32015
rect 22010 32049 25022 32062
rect 22010 32015 22193 32049
rect 22227 32015 22393 32049
rect 22427 32015 22593 32049
rect 22627 32015 22793 32049
rect 22827 32015 22993 32049
rect 23027 32015 23193 32049
rect 23227 32015 23393 32049
rect 23427 32015 23593 32049
rect 23627 32015 23793 32049
rect 23827 32015 23993 32049
rect 24027 32015 24193 32049
rect 24227 32015 24393 32049
rect 24427 32015 24593 32049
rect 24627 32015 24793 32049
rect 24827 32015 25022 32049
rect 22010 32002 25022 32015
rect 26204 32049 33372 32062
rect 26204 32015 26387 32049
rect 26421 32015 26787 32049
rect 26821 32015 27187 32049
rect 27221 32015 27587 32049
rect 27621 32015 27987 32049
rect 28021 32015 28387 32049
rect 28421 32015 28787 32049
rect 28821 32015 29187 32049
rect 29221 32015 29587 32049
rect 29621 32015 29987 32049
rect 30021 32015 30387 32049
rect 30421 32015 30787 32049
rect 30821 32015 31187 32049
rect 31221 32015 31587 32049
rect 31621 32015 31987 32049
rect 32021 32015 32387 32049
rect 32421 32015 32787 32049
rect 32821 32015 33187 32049
rect 33221 32015 33372 32049
rect 26204 32002 33372 32015
rect 33652 32049 40820 32062
rect 33652 32015 33835 32049
rect 33869 32015 34235 32049
rect 34269 32015 34635 32049
rect 34669 32015 35035 32049
rect 35069 32015 35435 32049
rect 35469 32015 35835 32049
rect 35869 32015 36235 32049
rect 36269 32015 36635 32049
rect 36669 32015 37035 32049
rect 37069 32015 37435 32049
rect 37469 32015 37835 32049
rect 37869 32015 38235 32049
rect 38269 32015 38635 32049
rect 38669 32015 39035 32049
rect 39069 32015 39435 32049
rect 39469 32015 39835 32049
rect 39869 32015 40235 32049
rect 40269 32015 40635 32049
rect 40669 32015 40820 32049
rect 33652 32002 40820 32015
rect 41784 32049 52504 32062
rect 41784 32015 41967 32049
rect 42001 32015 42167 32049
rect 42201 32015 42367 32049
rect 42401 32015 42567 32049
rect 42601 32015 42767 32049
rect 42801 32015 42967 32049
rect 43001 32015 43167 32049
rect 43201 32015 43367 32049
rect 43401 32015 43567 32049
rect 43601 32015 43767 32049
rect 43801 32015 43967 32049
rect 44001 32015 44167 32049
rect 44201 32015 44367 32049
rect 44401 32015 44567 32049
rect 44601 32015 44767 32049
rect 44801 32015 44967 32049
rect 45001 32015 45167 32049
rect 45201 32015 45367 32049
rect 45401 32015 45567 32049
rect 45601 32015 45767 32049
rect 45801 32015 45967 32049
rect 46001 32015 46167 32049
rect 46201 32015 46367 32049
rect 46401 32015 46567 32049
rect 46601 32015 46767 32049
rect 46801 32015 46967 32049
rect 47001 32015 47167 32049
rect 47201 32015 47367 32049
rect 47401 32015 47567 32049
rect 47601 32015 47767 32049
rect 47801 32015 47967 32049
rect 48001 32015 48167 32049
rect 48201 32015 48367 32049
rect 48401 32015 48567 32049
rect 48601 32015 48767 32049
rect 48801 32015 48967 32049
rect 49001 32015 49167 32049
rect 49201 32015 49367 32049
rect 49401 32015 49567 32049
rect 49601 32015 49767 32049
rect 49801 32015 49967 32049
rect 50001 32015 50167 32049
rect 50201 32015 50367 32049
rect 50401 32015 50567 32049
rect 50601 32015 50767 32049
rect 50801 32015 50967 32049
rect 51001 32015 51167 32049
rect 51201 32015 51367 32049
rect 51401 32015 51567 32049
rect 51601 32015 51767 32049
rect 51801 32015 51967 32049
rect 52001 32015 52167 32049
rect 52201 32015 52367 32049
rect 52401 32015 52504 32049
rect 41784 32002 52504 32015
rect 16520 30169 18960 30182
rect 16520 30135 16703 30169
rect 16737 30135 16903 30169
rect 16937 30135 17103 30169
rect 17137 30135 17303 30169
rect 17337 30135 17503 30169
rect 17537 30135 17703 30169
rect 17737 30135 17903 30169
rect 17937 30135 18103 30169
rect 18137 30135 18303 30169
rect 18337 30135 18503 30169
rect 18537 30135 18703 30169
rect 18737 30135 18960 30169
rect 16520 30122 18960 30135
rect 19264 30169 21704 30182
rect 19264 30135 19447 30169
rect 19481 30135 19647 30169
rect 19681 30135 19847 30169
rect 19881 30135 20047 30169
rect 20081 30135 20247 30169
rect 20281 30135 20447 30169
rect 20481 30135 20647 30169
rect 20681 30135 20847 30169
rect 20881 30135 21047 30169
rect 21081 30135 21247 30169
rect 21281 30135 21447 30169
rect 21481 30135 21704 30169
rect 19264 30122 21704 30135
rect 22008 30169 24448 30182
rect 22008 30135 22191 30169
rect 22225 30135 22391 30169
rect 22425 30135 22591 30169
rect 22625 30135 22791 30169
rect 22825 30135 22991 30169
rect 23025 30135 23191 30169
rect 23225 30135 23391 30169
rect 23425 30135 23591 30169
rect 23625 30135 23791 30169
rect 23825 30135 23991 30169
rect 24025 30135 24191 30169
rect 24225 30135 24448 30169
rect 22008 30122 24448 30135
rect 27202 30169 29642 30182
rect 27202 30135 27385 30169
rect 27419 30135 27585 30169
rect 27619 30135 27785 30169
rect 27819 30135 27985 30169
rect 28019 30135 28185 30169
rect 28219 30135 28385 30169
rect 28419 30135 28585 30169
rect 28619 30135 28785 30169
rect 28819 30135 28985 30169
rect 29019 30135 29185 30169
rect 29219 30135 29385 30169
rect 29419 30135 29642 30169
rect 27202 30122 29642 30135
rect 29928 30169 37096 30182
rect 29928 30135 30111 30169
rect 30145 30135 30511 30169
rect 30545 30135 30911 30169
rect 30945 30135 31311 30169
rect 31345 30135 31711 30169
rect 31745 30135 32111 30169
rect 32145 30135 32511 30169
rect 32545 30135 32911 30169
rect 32945 30135 33311 30169
rect 33345 30135 33711 30169
rect 33745 30135 34111 30169
rect 34145 30135 34511 30169
rect 34545 30135 34911 30169
rect 34945 30135 35311 30169
rect 35345 30135 35711 30169
rect 35745 30135 36111 30169
rect 36145 30135 36511 30169
rect 36545 30135 36911 30169
rect 36945 30135 37096 30169
rect 29928 30122 37096 30135
rect 37374 30169 40348 30182
rect 37374 30135 37655 30169
rect 37689 30135 38055 30169
rect 38089 30135 38455 30169
rect 38489 30135 38855 30169
rect 38889 30135 39255 30169
rect 39289 30135 39655 30169
rect 39689 30135 40055 30169
rect 40089 30135 40348 30169
rect 37374 30122 40348 30135
rect 41784 30169 52504 30182
rect 41784 30135 41967 30169
rect 42001 30135 42167 30169
rect 42201 30135 42367 30169
rect 42401 30135 42567 30169
rect 42601 30135 42767 30169
rect 42801 30135 42967 30169
rect 43001 30135 43167 30169
rect 43201 30135 43367 30169
rect 43401 30135 43567 30169
rect 43601 30135 43767 30169
rect 43801 30135 43967 30169
rect 44001 30135 44167 30169
rect 44201 30135 44367 30169
rect 44401 30135 44567 30169
rect 44601 30135 44767 30169
rect 44801 30135 44967 30169
rect 45001 30135 45167 30169
rect 45201 30135 45367 30169
rect 45401 30135 45567 30169
rect 45601 30135 45767 30169
rect 45801 30135 45967 30169
rect 46001 30135 46167 30169
rect 46201 30135 46367 30169
rect 46401 30135 46567 30169
rect 46601 30135 46767 30169
rect 46801 30135 46967 30169
rect 47001 30135 47167 30169
rect 47201 30135 47367 30169
rect 47401 30135 47567 30169
rect 47601 30135 47767 30169
rect 47801 30135 47967 30169
rect 48001 30135 48167 30169
rect 48201 30135 48367 30169
rect 48401 30135 48567 30169
rect 48601 30135 48767 30169
rect 48801 30135 48967 30169
rect 49001 30135 49167 30169
rect 49201 30135 49367 30169
rect 49401 30135 49567 30169
rect 49601 30135 49767 30169
rect 49801 30135 49967 30169
rect 50001 30135 50167 30169
rect 50201 30135 50367 30169
rect 50401 30135 50567 30169
rect 50601 30135 50767 30169
rect 50801 30135 50967 30169
rect 51001 30135 51167 30169
rect 51201 30135 51367 30169
rect 51401 30135 51567 30169
rect 51601 30135 51767 30169
rect 51801 30135 51967 30169
rect 52001 30135 52167 30169
rect 52201 30135 52367 30169
rect 52401 30135 52504 30169
rect 41784 30122 52504 30135
rect 37402 30029 37462 30122
rect 38450 30079 38610 30122
rect 38450 30045 38515 30079
rect 38549 30045 38610 30079
rect 38450 30042 38610 30045
rect 37402 29995 37415 30029
rect 37449 29995 37462 30029
rect 37402 29912 37462 29995
rect 37532 29999 40348 30002
rect 37532 29965 40325 29999
rect 37532 29962 40348 29965
rect 17432 29203 18048 29242
rect 17432 29101 17519 29203
rect 17961 29101 18048 29203
rect 17432 28302 18048 29101
rect 18528 28957 18960 29347
rect 20176 29203 20792 29242
rect 20176 29101 20263 29203
rect 20705 29101 20792 29203
rect 20176 28302 20792 29101
rect 21272 28957 21704 29347
rect 22920 29203 23536 29242
rect 22920 29101 23007 29203
rect 23449 29101 23536 29203
rect 22920 28302 23536 29101
rect 24016 28957 24448 29347
rect 28114 29203 28730 29242
rect 28114 29101 28201 29203
rect 28643 29101 28730 29203
rect 28114 28302 28730 29101
rect 29210 28957 29642 29347
rect 37519 29901 37553 29921
rect 37519 29833 37553 29867
rect 37519 29765 37553 29795
rect 37519 29697 37553 29723
rect 37519 29629 37553 29651
rect 37519 29561 37553 29579
rect 37519 29493 37553 29507
rect 37519 29425 37553 29435
rect 37519 29357 37553 29363
rect 37519 29289 37553 29291
rect 37519 29253 37553 29255
rect 37519 29181 37553 29187
rect 37519 29109 37553 29119
rect 37519 29037 37553 29051
rect 37519 28965 37553 28983
rect 37519 28893 37553 28915
rect 37519 28821 37553 28847
rect 37519 28749 37553 28779
rect 37519 28677 37553 28711
rect 37519 28542 37553 28643
rect 37977 29901 38011 29962
rect 37977 29833 38011 29867
rect 37977 29765 38011 29795
rect 37977 29697 38011 29723
rect 37977 29629 38011 29651
rect 37977 29561 38011 29579
rect 37977 29493 38011 29507
rect 37977 29425 38011 29435
rect 37977 29357 38011 29363
rect 37977 29289 38011 29291
rect 37977 29253 38011 29255
rect 37977 29181 38011 29187
rect 37977 29109 38011 29119
rect 37977 29037 38011 29051
rect 37977 28965 38011 28983
rect 37977 28893 38011 28915
rect 37977 28821 38011 28847
rect 37977 28749 38011 28779
rect 37977 28677 38011 28711
rect 37977 28623 38011 28643
rect 38435 29901 38469 29921
rect 38435 29833 38469 29867
rect 38435 29765 38469 29795
rect 38435 29697 38469 29723
rect 38435 29629 38469 29651
rect 38435 29561 38469 29579
rect 38435 29493 38469 29507
rect 38435 29425 38469 29435
rect 38435 29357 38469 29363
rect 38435 29289 38469 29291
rect 38435 29253 38469 29255
rect 38435 29181 38469 29187
rect 38435 29109 38469 29119
rect 38435 29037 38469 29051
rect 38435 28965 38469 28983
rect 38435 28893 38469 28915
rect 38435 28821 38469 28847
rect 38435 28749 38469 28779
rect 38435 28677 38469 28711
rect 38435 28542 38469 28643
rect 38893 29901 38927 29962
rect 38893 29833 38927 29867
rect 38893 29765 38927 29795
rect 38893 29697 38927 29723
rect 38893 29629 38927 29651
rect 38893 29561 38927 29579
rect 38893 29493 38927 29507
rect 38893 29425 38927 29435
rect 38893 29357 38927 29363
rect 38893 29289 38927 29291
rect 38893 29253 38927 29255
rect 38893 29181 38927 29187
rect 38893 29109 38927 29119
rect 38893 29037 38927 29051
rect 38893 28965 38927 28983
rect 38893 28893 38927 28915
rect 38893 28821 38927 28847
rect 38893 28749 38927 28779
rect 38893 28677 38927 28711
rect 38893 28623 38927 28643
rect 39351 29901 39385 29921
rect 39351 29833 39385 29867
rect 39351 29765 39385 29795
rect 39351 29697 39385 29723
rect 39351 29629 39385 29651
rect 39351 29561 39385 29579
rect 39351 29493 39385 29507
rect 39351 29425 39385 29435
rect 39351 29357 39385 29363
rect 39351 29289 39385 29291
rect 39351 29253 39385 29255
rect 39351 29181 39385 29187
rect 39351 29109 39385 29119
rect 39351 29037 39385 29051
rect 39351 28965 39385 28983
rect 39351 28893 39385 28915
rect 39351 28821 39385 28847
rect 39351 28749 39385 28779
rect 39351 28677 39385 28711
rect 37472 28509 38577 28542
rect 39351 28542 39385 28643
rect 39809 29901 39843 29962
rect 39809 29833 39843 29867
rect 39809 29765 39843 29795
rect 39809 29697 39843 29723
rect 39809 29629 39843 29651
rect 39809 29561 39843 29579
rect 39809 29493 39843 29507
rect 39809 29425 39843 29435
rect 39809 29357 39843 29363
rect 39809 29289 39843 29291
rect 39809 29253 39843 29255
rect 39809 29181 39843 29187
rect 39809 29109 39843 29119
rect 39809 29037 39843 29051
rect 39809 28965 39843 28983
rect 39809 28893 39843 28915
rect 39809 28821 39843 28847
rect 39809 28749 39843 28779
rect 39809 28677 39843 28711
rect 39809 28623 39843 28643
rect 40267 29901 40301 29921
rect 40267 29833 40301 29867
rect 40267 29765 40301 29795
rect 40267 29697 40301 29723
rect 40267 29629 40301 29651
rect 40267 29561 40301 29579
rect 40267 29493 40301 29507
rect 40267 29425 40301 29435
rect 40267 29357 40301 29363
rect 40267 29289 40301 29291
rect 40267 29253 40301 29255
rect 40267 29181 40301 29187
rect 40267 29109 40301 29119
rect 40267 29037 40301 29051
rect 40267 28965 40301 28983
rect 40267 28893 40301 28915
rect 40267 28821 40301 28847
rect 40267 28749 40301 28779
rect 40267 28677 40301 28711
rect 40267 28542 40301 28643
rect 41810 29836 52478 29856
rect 41810 29802 41830 29836
rect 41864 29802 41920 29836
rect 41954 29821 42010 29836
rect 42044 29821 42100 29836
rect 42134 29821 42190 29836
rect 42224 29821 42280 29836
rect 42314 29821 42370 29836
rect 42404 29821 42460 29836
rect 42494 29821 42550 29836
rect 42584 29821 42640 29836
rect 42674 29821 42730 29836
rect 42764 29821 42820 29836
rect 42854 29821 42910 29836
rect 42944 29821 43000 29836
rect 41974 29802 42010 29821
rect 42064 29802 42100 29821
rect 42154 29802 42190 29821
rect 42244 29802 42280 29821
rect 42334 29802 42370 29821
rect 42424 29802 42460 29821
rect 42514 29802 42550 29821
rect 42604 29802 42640 29821
rect 42694 29802 42730 29821
rect 42784 29802 42820 29821
rect 42874 29802 42910 29821
rect 42964 29802 43000 29821
rect 43034 29802 43170 29836
rect 43204 29802 43260 29836
rect 43294 29821 43350 29836
rect 43384 29821 43440 29836
rect 43474 29821 43530 29836
rect 43564 29821 43620 29836
rect 43654 29821 43710 29836
rect 43744 29821 43800 29836
rect 43834 29821 43890 29836
rect 43924 29821 43980 29836
rect 44014 29821 44070 29836
rect 44104 29821 44160 29836
rect 44194 29821 44250 29836
rect 44284 29821 44340 29836
rect 43314 29802 43350 29821
rect 43404 29802 43440 29821
rect 43494 29802 43530 29821
rect 43584 29802 43620 29821
rect 43674 29802 43710 29821
rect 43764 29802 43800 29821
rect 43854 29802 43890 29821
rect 43944 29802 43980 29821
rect 44034 29802 44070 29821
rect 44124 29802 44160 29821
rect 44214 29802 44250 29821
rect 44304 29802 44340 29821
rect 44374 29802 44510 29836
rect 44544 29802 44600 29836
rect 44634 29821 44690 29836
rect 44724 29821 44780 29836
rect 44814 29821 44870 29836
rect 44904 29821 44960 29836
rect 44994 29821 45050 29836
rect 45084 29821 45140 29836
rect 45174 29821 45230 29836
rect 45264 29821 45320 29836
rect 45354 29821 45410 29836
rect 45444 29821 45500 29836
rect 45534 29821 45590 29836
rect 45624 29821 45680 29836
rect 44654 29802 44690 29821
rect 44744 29802 44780 29821
rect 44834 29802 44870 29821
rect 44924 29802 44960 29821
rect 45014 29802 45050 29821
rect 45104 29802 45140 29821
rect 45194 29802 45230 29821
rect 45284 29802 45320 29821
rect 45374 29802 45410 29821
rect 45464 29802 45500 29821
rect 45554 29802 45590 29821
rect 45644 29802 45680 29821
rect 45714 29802 45850 29836
rect 45884 29802 45940 29836
rect 45974 29821 46030 29836
rect 46064 29821 46120 29836
rect 46154 29821 46210 29836
rect 46244 29821 46300 29836
rect 46334 29821 46390 29836
rect 46424 29821 46480 29836
rect 46514 29821 46570 29836
rect 46604 29821 46660 29836
rect 46694 29821 46750 29836
rect 46784 29821 46840 29836
rect 46874 29821 46930 29836
rect 46964 29821 47020 29836
rect 45994 29802 46030 29821
rect 46084 29802 46120 29821
rect 46174 29802 46210 29821
rect 46264 29802 46300 29821
rect 46354 29802 46390 29821
rect 46444 29802 46480 29821
rect 46534 29802 46570 29821
rect 46624 29802 46660 29821
rect 46714 29802 46750 29821
rect 46804 29802 46840 29821
rect 46894 29802 46930 29821
rect 46984 29802 47020 29821
rect 47054 29802 47190 29836
rect 47224 29802 47280 29836
rect 47314 29821 47370 29836
rect 47404 29821 47460 29836
rect 47494 29821 47550 29836
rect 47584 29821 47640 29836
rect 47674 29821 47730 29836
rect 47764 29821 47820 29836
rect 47854 29821 47910 29836
rect 47944 29821 48000 29836
rect 48034 29821 48090 29836
rect 48124 29821 48180 29836
rect 48214 29821 48270 29836
rect 48304 29821 48360 29836
rect 47334 29802 47370 29821
rect 47424 29802 47460 29821
rect 47514 29802 47550 29821
rect 47604 29802 47640 29821
rect 47694 29802 47730 29821
rect 47784 29802 47820 29821
rect 47874 29802 47910 29821
rect 47964 29802 48000 29821
rect 48054 29802 48090 29821
rect 48144 29802 48180 29821
rect 48234 29802 48270 29821
rect 48324 29802 48360 29821
rect 48394 29802 48530 29836
rect 48564 29802 48620 29836
rect 48654 29821 48710 29836
rect 48744 29821 48800 29836
rect 48834 29821 48890 29836
rect 48924 29821 48980 29836
rect 49014 29821 49070 29836
rect 49104 29821 49160 29836
rect 49194 29821 49250 29836
rect 49284 29821 49340 29836
rect 49374 29821 49430 29836
rect 49464 29821 49520 29836
rect 49554 29821 49610 29836
rect 49644 29821 49700 29836
rect 48674 29802 48710 29821
rect 48764 29802 48800 29821
rect 48854 29802 48890 29821
rect 48944 29802 48980 29821
rect 49034 29802 49070 29821
rect 49124 29802 49160 29821
rect 49214 29802 49250 29821
rect 49304 29802 49340 29821
rect 49394 29802 49430 29821
rect 49484 29802 49520 29821
rect 49574 29802 49610 29821
rect 49664 29802 49700 29821
rect 49734 29802 49870 29836
rect 49904 29802 49960 29836
rect 49994 29821 50050 29836
rect 50084 29821 50140 29836
rect 50174 29821 50230 29836
rect 50264 29821 50320 29836
rect 50354 29821 50410 29836
rect 50444 29821 50500 29836
rect 50534 29821 50590 29836
rect 50624 29821 50680 29836
rect 50714 29821 50770 29836
rect 50804 29821 50860 29836
rect 50894 29821 50950 29836
rect 50984 29821 51040 29836
rect 50014 29802 50050 29821
rect 50104 29802 50140 29821
rect 50194 29802 50230 29821
rect 50284 29802 50320 29821
rect 50374 29802 50410 29821
rect 50464 29802 50500 29821
rect 50554 29802 50590 29821
rect 50644 29802 50680 29821
rect 50734 29802 50770 29821
rect 50824 29802 50860 29821
rect 50914 29802 50950 29821
rect 51004 29802 51040 29821
rect 51074 29802 51210 29836
rect 51244 29802 51300 29836
rect 51334 29821 51390 29836
rect 51424 29821 51480 29836
rect 51514 29821 51570 29836
rect 51604 29821 51660 29836
rect 51694 29821 51750 29836
rect 51784 29821 51840 29836
rect 51874 29821 51930 29836
rect 51964 29821 52020 29836
rect 52054 29821 52110 29836
rect 52144 29821 52200 29836
rect 52234 29821 52290 29836
rect 52324 29821 52380 29836
rect 51354 29802 51390 29821
rect 51444 29802 51480 29821
rect 51534 29802 51570 29821
rect 51624 29802 51660 29821
rect 51714 29802 51750 29821
rect 51804 29802 51840 29821
rect 51894 29802 51930 29821
rect 51984 29802 52020 29821
rect 52074 29802 52110 29821
rect 52164 29802 52200 29821
rect 52254 29802 52290 29821
rect 52344 29802 52380 29821
rect 52414 29802 52478 29836
rect 41810 29798 41940 29802
rect 41810 29764 41844 29798
rect 41878 29787 41940 29798
rect 41974 29787 42030 29802
rect 42064 29787 42120 29802
rect 42154 29787 42210 29802
rect 42244 29787 42300 29802
rect 42334 29787 42390 29802
rect 42424 29787 42480 29802
rect 42514 29787 42570 29802
rect 42604 29787 42660 29802
rect 42694 29787 42750 29802
rect 42784 29787 42840 29802
rect 42874 29787 42930 29802
rect 42964 29798 43280 29802
rect 42964 29787 43031 29798
rect 41878 29764 43031 29787
rect 43065 29764 43184 29798
rect 43218 29787 43280 29798
rect 43314 29787 43370 29802
rect 43404 29787 43460 29802
rect 43494 29787 43550 29802
rect 43584 29787 43640 29802
rect 43674 29787 43730 29802
rect 43764 29787 43820 29802
rect 43854 29787 43910 29802
rect 43944 29787 44000 29802
rect 44034 29787 44090 29802
rect 44124 29787 44180 29802
rect 44214 29787 44270 29802
rect 44304 29798 44620 29802
rect 44304 29787 44371 29798
rect 43218 29764 44371 29787
rect 44405 29764 44524 29798
rect 44558 29787 44620 29798
rect 44654 29787 44710 29802
rect 44744 29787 44800 29802
rect 44834 29787 44890 29802
rect 44924 29787 44980 29802
rect 45014 29787 45070 29802
rect 45104 29787 45160 29802
rect 45194 29787 45250 29802
rect 45284 29787 45340 29802
rect 45374 29787 45430 29802
rect 45464 29787 45520 29802
rect 45554 29787 45610 29802
rect 45644 29798 45960 29802
rect 45644 29787 45711 29798
rect 44558 29764 45711 29787
rect 45745 29764 45864 29798
rect 45898 29787 45960 29798
rect 45994 29787 46050 29802
rect 46084 29787 46140 29802
rect 46174 29787 46230 29802
rect 46264 29787 46320 29802
rect 46354 29787 46410 29802
rect 46444 29787 46500 29802
rect 46534 29787 46590 29802
rect 46624 29787 46680 29802
rect 46714 29787 46770 29802
rect 46804 29787 46860 29802
rect 46894 29787 46950 29802
rect 46984 29798 47300 29802
rect 46984 29787 47051 29798
rect 45898 29764 47051 29787
rect 47085 29764 47204 29798
rect 47238 29787 47300 29798
rect 47334 29787 47390 29802
rect 47424 29787 47480 29802
rect 47514 29787 47570 29802
rect 47604 29787 47660 29802
rect 47694 29787 47750 29802
rect 47784 29787 47840 29802
rect 47874 29787 47930 29802
rect 47964 29787 48020 29802
rect 48054 29787 48110 29802
rect 48144 29787 48200 29802
rect 48234 29787 48290 29802
rect 48324 29798 48640 29802
rect 48324 29787 48391 29798
rect 47238 29764 48391 29787
rect 48425 29764 48544 29798
rect 48578 29787 48640 29798
rect 48674 29787 48730 29802
rect 48764 29787 48820 29802
rect 48854 29787 48910 29802
rect 48944 29787 49000 29802
rect 49034 29787 49090 29802
rect 49124 29787 49180 29802
rect 49214 29787 49270 29802
rect 49304 29787 49360 29802
rect 49394 29787 49450 29802
rect 49484 29787 49540 29802
rect 49574 29787 49630 29802
rect 49664 29798 49980 29802
rect 49664 29787 49731 29798
rect 48578 29764 49731 29787
rect 49765 29764 49884 29798
rect 49918 29787 49980 29798
rect 50014 29787 50070 29802
rect 50104 29787 50160 29802
rect 50194 29787 50250 29802
rect 50284 29787 50340 29802
rect 50374 29787 50430 29802
rect 50464 29787 50520 29802
rect 50554 29787 50610 29802
rect 50644 29787 50700 29802
rect 50734 29787 50790 29802
rect 50824 29787 50880 29802
rect 50914 29787 50970 29802
rect 51004 29798 51320 29802
rect 51004 29787 51071 29798
rect 49918 29764 51071 29787
rect 51105 29764 51224 29798
rect 51258 29787 51320 29798
rect 51354 29787 51410 29802
rect 51444 29787 51500 29802
rect 51534 29787 51590 29802
rect 51624 29787 51680 29802
rect 51714 29787 51770 29802
rect 51804 29787 51860 29802
rect 51894 29787 51950 29802
rect 51984 29787 52040 29802
rect 52074 29787 52130 29802
rect 52164 29787 52220 29802
rect 52254 29787 52310 29802
rect 52344 29798 52478 29802
rect 52344 29787 52411 29798
rect 51258 29764 52411 29787
rect 52445 29764 52478 29798
rect 41810 29757 52478 29764
rect 41810 29708 41909 29757
rect 41810 29674 41844 29708
rect 41878 29674 41909 29708
rect 42999 29708 43249 29757
rect 41810 29618 41909 29674
rect 41810 29584 41844 29618
rect 41878 29584 41909 29618
rect 41810 29528 41909 29584
rect 41810 29494 41844 29528
rect 41878 29494 41909 29528
rect 41810 29438 41909 29494
rect 41810 29404 41844 29438
rect 41878 29404 41909 29438
rect 41810 29348 41909 29404
rect 41810 29314 41844 29348
rect 41878 29314 41909 29348
rect 41810 29258 41909 29314
rect 41810 29224 41844 29258
rect 41878 29224 41909 29258
rect 41810 29168 41909 29224
rect 41810 29134 41844 29168
rect 41878 29134 41909 29168
rect 41810 29078 41909 29134
rect 41810 29044 41844 29078
rect 41878 29044 41909 29078
rect 41810 28988 41909 29044
rect 41810 28954 41844 28988
rect 41878 28954 41909 28988
rect 41810 28898 41909 28954
rect 41810 28864 41844 28898
rect 41878 28864 41909 28898
rect 41810 28808 41909 28864
rect 41810 28774 41844 28808
rect 41878 28774 41909 28808
rect 41810 28718 41909 28774
rect 41973 29676 42935 29693
rect 41973 29642 41994 29676
rect 42028 29642 42084 29676
rect 42118 29674 42174 29676
rect 42208 29674 42264 29676
rect 42298 29674 42354 29676
rect 42388 29674 42444 29676
rect 42478 29674 42534 29676
rect 42568 29674 42624 29676
rect 42658 29674 42714 29676
rect 42748 29674 42804 29676
rect 42838 29674 42894 29676
rect 42138 29642 42174 29674
rect 42228 29642 42264 29674
rect 42318 29642 42354 29674
rect 42408 29642 42444 29674
rect 42498 29642 42534 29674
rect 42588 29642 42624 29674
rect 42678 29642 42714 29674
rect 42768 29642 42804 29674
rect 42858 29642 42894 29674
rect 42928 29642 42935 29676
rect 41973 29640 42104 29642
rect 42138 29640 42194 29642
rect 42228 29640 42284 29642
rect 42318 29640 42374 29642
rect 42408 29640 42464 29642
rect 42498 29640 42554 29642
rect 42588 29640 42644 29642
rect 42678 29640 42734 29642
rect 42768 29640 42824 29642
rect 42858 29640 42935 29642
rect 41973 29621 42935 29640
rect 41973 29617 42045 29621
rect 41973 29583 41992 29617
rect 42026 29583 42045 29617
rect 41973 29527 42045 29583
rect 42863 29598 42935 29621
rect 42863 29564 42882 29598
rect 42916 29564 42935 29598
rect 41973 29493 41992 29527
rect 42026 29493 42045 29527
rect 41973 29437 42045 29493
rect 41973 29403 41992 29437
rect 42026 29403 42045 29437
rect 41973 29347 42045 29403
rect 41973 29313 41992 29347
rect 42026 29313 42045 29347
rect 41973 29257 42045 29313
rect 41973 29223 41992 29257
rect 42026 29223 42045 29257
rect 41973 29167 42045 29223
rect 41973 29133 41992 29167
rect 42026 29133 42045 29167
rect 41973 29077 42045 29133
rect 41973 29043 41992 29077
rect 42026 29043 42045 29077
rect 41973 28987 42045 29043
rect 41973 28953 41992 28987
rect 42026 28953 42045 28987
rect 41973 28897 42045 28953
rect 41973 28863 41992 28897
rect 42026 28863 42045 28897
rect 42107 29500 42801 29559
rect 42107 29466 42168 29500
rect 42202 29472 42258 29500
rect 42292 29472 42348 29500
rect 42382 29472 42438 29500
rect 42214 29466 42258 29472
rect 42314 29466 42348 29472
rect 42414 29466 42438 29472
rect 42472 29472 42528 29500
rect 42472 29466 42480 29472
rect 42107 29438 42180 29466
rect 42214 29438 42280 29466
rect 42314 29438 42380 29466
rect 42414 29438 42480 29466
rect 42514 29466 42528 29472
rect 42562 29472 42618 29500
rect 42562 29466 42580 29472
rect 42514 29438 42580 29466
rect 42614 29466 42618 29472
rect 42652 29472 42708 29500
rect 42652 29466 42680 29472
rect 42742 29466 42801 29500
rect 42614 29438 42680 29466
rect 42714 29438 42801 29466
rect 42107 29410 42801 29438
rect 42107 29376 42168 29410
rect 42202 29376 42258 29410
rect 42292 29376 42348 29410
rect 42382 29376 42438 29410
rect 42472 29376 42528 29410
rect 42562 29376 42618 29410
rect 42652 29376 42708 29410
rect 42742 29376 42801 29410
rect 42107 29372 42801 29376
rect 42107 29338 42180 29372
rect 42214 29338 42280 29372
rect 42314 29338 42380 29372
rect 42414 29338 42480 29372
rect 42514 29338 42580 29372
rect 42614 29338 42680 29372
rect 42714 29338 42801 29372
rect 42107 29320 42801 29338
rect 42107 29286 42168 29320
rect 42202 29286 42258 29320
rect 42292 29286 42348 29320
rect 42382 29286 42438 29320
rect 42472 29286 42528 29320
rect 42562 29286 42618 29320
rect 42652 29286 42708 29320
rect 42742 29286 42801 29320
rect 42107 29272 42801 29286
rect 42107 29238 42180 29272
rect 42214 29238 42280 29272
rect 42314 29238 42380 29272
rect 42414 29238 42480 29272
rect 42514 29238 42580 29272
rect 42614 29238 42680 29272
rect 42714 29238 42801 29272
rect 42107 29230 42801 29238
rect 42107 29196 42168 29230
rect 42202 29196 42258 29230
rect 42292 29196 42348 29230
rect 42382 29196 42438 29230
rect 42472 29196 42528 29230
rect 42562 29196 42618 29230
rect 42652 29196 42708 29230
rect 42742 29196 42801 29230
rect 42107 29172 42801 29196
rect 42107 29140 42180 29172
rect 42214 29140 42280 29172
rect 42314 29140 42380 29172
rect 42414 29140 42480 29172
rect 42107 29106 42168 29140
rect 42214 29138 42258 29140
rect 42314 29138 42348 29140
rect 42414 29138 42438 29140
rect 42202 29106 42258 29138
rect 42292 29106 42348 29138
rect 42382 29106 42438 29138
rect 42472 29138 42480 29140
rect 42514 29140 42580 29172
rect 42514 29138 42528 29140
rect 42472 29106 42528 29138
rect 42562 29138 42580 29140
rect 42614 29140 42680 29172
rect 42714 29140 42801 29172
rect 42614 29138 42618 29140
rect 42562 29106 42618 29138
rect 42652 29138 42680 29140
rect 42652 29106 42708 29138
rect 42742 29106 42801 29140
rect 42107 29072 42801 29106
rect 42107 29050 42180 29072
rect 42214 29050 42280 29072
rect 42314 29050 42380 29072
rect 42414 29050 42480 29072
rect 42107 29016 42168 29050
rect 42214 29038 42258 29050
rect 42314 29038 42348 29050
rect 42414 29038 42438 29050
rect 42202 29016 42258 29038
rect 42292 29016 42348 29038
rect 42382 29016 42438 29038
rect 42472 29038 42480 29050
rect 42514 29050 42580 29072
rect 42514 29038 42528 29050
rect 42472 29016 42528 29038
rect 42562 29038 42580 29050
rect 42614 29050 42680 29072
rect 42714 29050 42801 29072
rect 42614 29038 42618 29050
rect 42562 29016 42618 29038
rect 42652 29038 42680 29050
rect 42652 29016 42708 29038
rect 42742 29016 42801 29050
rect 42107 28972 42801 29016
rect 42107 28960 42180 28972
rect 42214 28960 42280 28972
rect 42314 28960 42380 28972
rect 42414 28960 42480 28972
rect 42107 28926 42168 28960
rect 42214 28938 42258 28960
rect 42314 28938 42348 28960
rect 42414 28938 42438 28960
rect 42202 28926 42258 28938
rect 42292 28926 42348 28938
rect 42382 28926 42438 28938
rect 42472 28938 42480 28960
rect 42514 28960 42580 28972
rect 42514 28938 42528 28960
rect 42472 28926 42528 28938
rect 42562 28938 42580 28960
rect 42614 28960 42680 28972
rect 42714 28960 42801 28972
rect 42614 28938 42618 28960
rect 42562 28926 42618 28938
rect 42652 28938 42680 28960
rect 42652 28926 42708 28938
rect 42742 28926 42801 28960
rect 42107 28865 42801 28926
rect 42863 29508 42935 29564
rect 42863 29474 42882 29508
rect 42916 29474 42935 29508
rect 42863 29418 42935 29474
rect 42863 29384 42882 29418
rect 42916 29384 42935 29418
rect 42863 29328 42935 29384
rect 42863 29294 42882 29328
rect 42916 29294 42935 29328
rect 42863 29238 42935 29294
rect 42863 29204 42882 29238
rect 42916 29204 42935 29238
rect 42863 29148 42935 29204
rect 42863 29114 42882 29148
rect 42916 29114 42935 29148
rect 42863 29058 42935 29114
rect 42863 29024 42882 29058
rect 42916 29024 42935 29058
rect 42863 28968 42935 29024
rect 42863 28934 42882 28968
rect 42916 28934 42935 28968
rect 42863 28878 42935 28934
rect 41973 28803 42045 28863
rect 42863 28844 42882 28878
rect 42916 28844 42935 28878
rect 42863 28803 42935 28844
rect 41973 28784 42935 28803
rect 41973 28750 42070 28784
rect 42104 28750 42160 28784
rect 42194 28750 42250 28784
rect 42284 28750 42340 28784
rect 42374 28750 42430 28784
rect 42464 28750 42520 28784
rect 42554 28750 42610 28784
rect 42644 28750 42700 28784
rect 42734 28750 42790 28784
rect 42824 28750 42935 28784
rect 41973 28731 42935 28750
rect 42999 29674 43031 29708
rect 43065 29674 43184 29708
rect 43218 29674 43249 29708
rect 44339 29708 44589 29757
rect 42999 29618 43249 29674
rect 42999 29584 43031 29618
rect 43065 29584 43184 29618
rect 43218 29584 43249 29618
rect 42999 29528 43249 29584
rect 42999 29494 43031 29528
rect 43065 29494 43184 29528
rect 43218 29494 43249 29528
rect 42999 29438 43249 29494
rect 42999 29404 43031 29438
rect 43065 29404 43184 29438
rect 43218 29404 43249 29438
rect 42999 29348 43249 29404
rect 42999 29314 43031 29348
rect 43065 29314 43184 29348
rect 43218 29314 43249 29348
rect 42999 29258 43249 29314
rect 42999 29224 43031 29258
rect 43065 29224 43184 29258
rect 43218 29224 43249 29258
rect 42999 29168 43249 29224
rect 42999 29134 43031 29168
rect 43065 29134 43184 29168
rect 43218 29134 43249 29168
rect 42999 29078 43249 29134
rect 42999 29044 43031 29078
rect 43065 29044 43184 29078
rect 43218 29044 43249 29078
rect 42999 28988 43249 29044
rect 42999 28954 43031 28988
rect 43065 28954 43184 28988
rect 43218 28954 43249 28988
rect 42999 28898 43249 28954
rect 42999 28864 43031 28898
rect 43065 28864 43184 28898
rect 43218 28864 43249 28898
rect 42999 28808 43249 28864
rect 42999 28774 43031 28808
rect 43065 28774 43184 28808
rect 43218 28774 43249 28808
rect 41810 28684 41844 28718
rect 41878 28684 41909 28718
rect 41810 28667 41909 28684
rect 42999 28718 43249 28774
rect 43313 29676 44275 29693
rect 43313 29642 43334 29676
rect 43368 29642 43424 29676
rect 43458 29674 43514 29676
rect 43548 29674 43604 29676
rect 43638 29674 43694 29676
rect 43728 29674 43784 29676
rect 43818 29674 43874 29676
rect 43908 29674 43964 29676
rect 43998 29674 44054 29676
rect 44088 29674 44144 29676
rect 44178 29674 44234 29676
rect 43478 29642 43514 29674
rect 43568 29642 43604 29674
rect 43658 29642 43694 29674
rect 43748 29642 43784 29674
rect 43838 29642 43874 29674
rect 43928 29642 43964 29674
rect 44018 29642 44054 29674
rect 44108 29642 44144 29674
rect 44198 29642 44234 29674
rect 44268 29642 44275 29676
rect 43313 29640 43444 29642
rect 43478 29640 43534 29642
rect 43568 29640 43624 29642
rect 43658 29640 43714 29642
rect 43748 29640 43804 29642
rect 43838 29640 43894 29642
rect 43928 29640 43984 29642
rect 44018 29640 44074 29642
rect 44108 29640 44164 29642
rect 44198 29640 44275 29642
rect 43313 29621 44275 29640
rect 43313 29617 43385 29621
rect 43313 29583 43332 29617
rect 43366 29583 43385 29617
rect 43313 29527 43385 29583
rect 44203 29598 44275 29621
rect 44203 29564 44222 29598
rect 44256 29564 44275 29598
rect 43313 29493 43332 29527
rect 43366 29493 43385 29527
rect 43313 29437 43385 29493
rect 43313 29403 43332 29437
rect 43366 29403 43385 29437
rect 43313 29347 43385 29403
rect 43313 29313 43332 29347
rect 43366 29313 43385 29347
rect 43313 29257 43385 29313
rect 43313 29223 43332 29257
rect 43366 29223 43385 29257
rect 43313 29167 43385 29223
rect 43313 29133 43332 29167
rect 43366 29133 43385 29167
rect 43313 29077 43385 29133
rect 43313 29043 43332 29077
rect 43366 29043 43385 29077
rect 43313 28987 43385 29043
rect 43313 28953 43332 28987
rect 43366 28953 43385 28987
rect 43313 28897 43385 28953
rect 43313 28863 43332 28897
rect 43366 28863 43385 28897
rect 43447 29500 44141 29559
rect 43447 29466 43508 29500
rect 43542 29472 43598 29500
rect 43632 29472 43688 29500
rect 43722 29472 43778 29500
rect 43554 29466 43598 29472
rect 43654 29466 43688 29472
rect 43754 29466 43778 29472
rect 43812 29472 43868 29500
rect 43812 29466 43820 29472
rect 43447 29438 43520 29466
rect 43554 29438 43620 29466
rect 43654 29438 43720 29466
rect 43754 29438 43820 29466
rect 43854 29466 43868 29472
rect 43902 29472 43958 29500
rect 43902 29466 43920 29472
rect 43854 29438 43920 29466
rect 43954 29466 43958 29472
rect 43992 29472 44048 29500
rect 43992 29466 44020 29472
rect 44082 29466 44141 29500
rect 43954 29438 44020 29466
rect 44054 29438 44141 29466
rect 43447 29410 44141 29438
rect 43447 29376 43508 29410
rect 43542 29376 43598 29410
rect 43632 29376 43688 29410
rect 43722 29376 43778 29410
rect 43812 29376 43868 29410
rect 43902 29376 43958 29410
rect 43992 29376 44048 29410
rect 44082 29376 44141 29410
rect 43447 29372 44141 29376
rect 43447 29338 43520 29372
rect 43554 29338 43620 29372
rect 43654 29338 43720 29372
rect 43754 29338 43820 29372
rect 43854 29338 43920 29372
rect 43954 29338 44020 29372
rect 44054 29338 44141 29372
rect 43447 29320 44141 29338
rect 43447 29286 43508 29320
rect 43542 29286 43598 29320
rect 43632 29286 43688 29320
rect 43722 29286 43778 29320
rect 43812 29286 43868 29320
rect 43902 29286 43958 29320
rect 43992 29286 44048 29320
rect 44082 29286 44141 29320
rect 43447 29272 44141 29286
rect 43447 29238 43520 29272
rect 43554 29238 43620 29272
rect 43654 29238 43720 29272
rect 43754 29238 43820 29272
rect 43854 29238 43920 29272
rect 43954 29238 44020 29272
rect 44054 29238 44141 29272
rect 43447 29230 44141 29238
rect 43447 29196 43508 29230
rect 43542 29196 43598 29230
rect 43632 29196 43688 29230
rect 43722 29196 43778 29230
rect 43812 29196 43868 29230
rect 43902 29196 43958 29230
rect 43992 29196 44048 29230
rect 44082 29196 44141 29230
rect 43447 29172 44141 29196
rect 43447 29140 43520 29172
rect 43554 29140 43620 29172
rect 43654 29140 43720 29172
rect 43754 29140 43820 29172
rect 43447 29106 43508 29140
rect 43554 29138 43598 29140
rect 43654 29138 43688 29140
rect 43754 29138 43778 29140
rect 43542 29106 43598 29138
rect 43632 29106 43688 29138
rect 43722 29106 43778 29138
rect 43812 29138 43820 29140
rect 43854 29140 43920 29172
rect 43854 29138 43868 29140
rect 43812 29106 43868 29138
rect 43902 29138 43920 29140
rect 43954 29140 44020 29172
rect 44054 29140 44141 29172
rect 43954 29138 43958 29140
rect 43902 29106 43958 29138
rect 43992 29138 44020 29140
rect 43992 29106 44048 29138
rect 44082 29106 44141 29140
rect 43447 29072 44141 29106
rect 43447 29050 43520 29072
rect 43554 29050 43620 29072
rect 43654 29050 43720 29072
rect 43754 29050 43820 29072
rect 43447 29016 43508 29050
rect 43554 29038 43598 29050
rect 43654 29038 43688 29050
rect 43754 29038 43778 29050
rect 43542 29016 43598 29038
rect 43632 29016 43688 29038
rect 43722 29016 43778 29038
rect 43812 29038 43820 29050
rect 43854 29050 43920 29072
rect 43854 29038 43868 29050
rect 43812 29016 43868 29038
rect 43902 29038 43920 29050
rect 43954 29050 44020 29072
rect 44054 29050 44141 29072
rect 43954 29038 43958 29050
rect 43902 29016 43958 29038
rect 43992 29038 44020 29050
rect 43992 29016 44048 29038
rect 44082 29016 44141 29050
rect 43447 28972 44141 29016
rect 43447 28960 43520 28972
rect 43554 28960 43620 28972
rect 43654 28960 43720 28972
rect 43754 28960 43820 28972
rect 43447 28926 43508 28960
rect 43554 28938 43598 28960
rect 43654 28938 43688 28960
rect 43754 28938 43778 28960
rect 43542 28926 43598 28938
rect 43632 28926 43688 28938
rect 43722 28926 43778 28938
rect 43812 28938 43820 28960
rect 43854 28960 43920 28972
rect 43854 28938 43868 28960
rect 43812 28926 43868 28938
rect 43902 28938 43920 28960
rect 43954 28960 44020 28972
rect 44054 28960 44141 28972
rect 43954 28938 43958 28960
rect 43902 28926 43958 28938
rect 43992 28938 44020 28960
rect 43992 28926 44048 28938
rect 44082 28926 44141 28960
rect 43447 28865 44141 28926
rect 44203 29508 44275 29564
rect 44203 29474 44222 29508
rect 44256 29474 44275 29508
rect 44203 29418 44275 29474
rect 44203 29384 44222 29418
rect 44256 29384 44275 29418
rect 44203 29328 44275 29384
rect 44203 29294 44222 29328
rect 44256 29294 44275 29328
rect 44203 29238 44275 29294
rect 44203 29204 44222 29238
rect 44256 29204 44275 29238
rect 44203 29148 44275 29204
rect 44203 29114 44222 29148
rect 44256 29114 44275 29148
rect 44203 29058 44275 29114
rect 44203 29024 44222 29058
rect 44256 29024 44275 29058
rect 44203 28968 44275 29024
rect 44203 28934 44222 28968
rect 44256 28934 44275 28968
rect 44203 28878 44275 28934
rect 43313 28803 43385 28863
rect 44203 28844 44222 28878
rect 44256 28844 44275 28878
rect 44203 28803 44275 28844
rect 43313 28784 44275 28803
rect 43313 28750 43410 28784
rect 43444 28750 43500 28784
rect 43534 28750 43590 28784
rect 43624 28750 43680 28784
rect 43714 28750 43770 28784
rect 43804 28750 43860 28784
rect 43894 28750 43950 28784
rect 43984 28750 44040 28784
rect 44074 28750 44130 28784
rect 44164 28750 44275 28784
rect 43313 28731 44275 28750
rect 44339 29674 44371 29708
rect 44405 29674 44524 29708
rect 44558 29674 44589 29708
rect 45679 29708 45929 29757
rect 44339 29618 44589 29674
rect 44339 29584 44371 29618
rect 44405 29584 44524 29618
rect 44558 29584 44589 29618
rect 44339 29528 44589 29584
rect 44339 29494 44371 29528
rect 44405 29494 44524 29528
rect 44558 29494 44589 29528
rect 44339 29438 44589 29494
rect 44339 29404 44371 29438
rect 44405 29404 44524 29438
rect 44558 29404 44589 29438
rect 44339 29348 44589 29404
rect 44339 29314 44371 29348
rect 44405 29314 44524 29348
rect 44558 29314 44589 29348
rect 44339 29258 44589 29314
rect 44339 29224 44371 29258
rect 44405 29224 44524 29258
rect 44558 29224 44589 29258
rect 44339 29168 44589 29224
rect 44339 29134 44371 29168
rect 44405 29134 44524 29168
rect 44558 29134 44589 29168
rect 44339 29078 44589 29134
rect 44339 29044 44371 29078
rect 44405 29044 44524 29078
rect 44558 29044 44589 29078
rect 44339 28988 44589 29044
rect 44339 28954 44371 28988
rect 44405 28954 44524 28988
rect 44558 28954 44589 28988
rect 44339 28898 44589 28954
rect 44339 28864 44371 28898
rect 44405 28864 44524 28898
rect 44558 28864 44589 28898
rect 44339 28808 44589 28864
rect 44339 28774 44371 28808
rect 44405 28774 44524 28808
rect 44558 28774 44589 28808
rect 42999 28684 43031 28718
rect 43065 28684 43184 28718
rect 43218 28684 43249 28718
rect 42999 28667 43249 28684
rect 44339 28718 44589 28774
rect 44653 29676 45615 29693
rect 44653 29642 44674 29676
rect 44708 29642 44764 29676
rect 44798 29674 44854 29676
rect 44888 29674 44944 29676
rect 44978 29674 45034 29676
rect 45068 29674 45124 29676
rect 45158 29674 45214 29676
rect 45248 29674 45304 29676
rect 45338 29674 45394 29676
rect 45428 29674 45484 29676
rect 45518 29674 45574 29676
rect 44818 29642 44854 29674
rect 44908 29642 44944 29674
rect 44998 29642 45034 29674
rect 45088 29642 45124 29674
rect 45178 29642 45214 29674
rect 45268 29642 45304 29674
rect 45358 29642 45394 29674
rect 45448 29642 45484 29674
rect 45538 29642 45574 29674
rect 45608 29642 45615 29676
rect 44653 29640 44784 29642
rect 44818 29640 44874 29642
rect 44908 29640 44964 29642
rect 44998 29640 45054 29642
rect 45088 29640 45144 29642
rect 45178 29640 45234 29642
rect 45268 29640 45324 29642
rect 45358 29640 45414 29642
rect 45448 29640 45504 29642
rect 45538 29640 45615 29642
rect 44653 29621 45615 29640
rect 44653 29617 44725 29621
rect 44653 29583 44672 29617
rect 44706 29583 44725 29617
rect 44653 29527 44725 29583
rect 45543 29598 45615 29621
rect 45543 29564 45562 29598
rect 45596 29564 45615 29598
rect 44653 29493 44672 29527
rect 44706 29493 44725 29527
rect 44653 29437 44725 29493
rect 44653 29403 44672 29437
rect 44706 29403 44725 29437
rect 44653 29347 44725 29403
rect 44653 29313 44672 29347
rect 44706 29313 44725 29347
rect 44653 29257 44725 29313
rect 44653 29223 44672 29257
rect 44706 29223 44725 29257
rect 44653 29167 44725 29223
rect 44653 29133 44672 29167
rect 44706 29133 44725 29167
rect 44653 29077 44725 29133
rect 44653 29043 44672 29077
rect 44706 29043 44725 29077
rect 44653 28987 44725 29043
rect 44653 28953 44672 28987
rect 44706 28953 44725 28987
rect 44653 28897 44725 28953
rect 44653 28863 44672 28897
rect 44706 28863 44725 28897
rect 44787 29500 45481 29559
rect 44787 29466 44848 29500
rect 44882 29472 44938 29500
rect 44972 29472 45028 29500
rect 45062 29472 45118 29500
rect 44894 29466 44938 29472
rect 44994 29466 45028 29472
rect 45094 29466 45118 29472
rect 45152 29472 45208 29500
rect 45152 29466 45160 29472
rect 44787 29438 44860 29466
rect 44894 29438 44960 29466
rect 44994 29438 45060 29466
rect 45094 29438 45160 29466
rect 45194 29466 45208 29472
rect 45242 29472 45298 29500
rect 45242 29466 45260 29472
rect 45194 29438 45260 29466
rect 45294 29466 45298 29472
rect 45332 29472 45388 29500
rect 45332 29466 45360 29472
rect 45422 29466 45481 29500
rect 45294 29438 45360 29466
rect 45394 29438 45481 29466
rect 44787 29410 45481 29438
rect 44787 29376 44848 29410
rect 44882 29376 44938 29410
rect 44972 29376 45028 29410
rect 45062 29376 45118 29410
rect 45152 29376 45208 29410
rect 45242 29376 45298 29410
rect 45332 29376 45388 29410
rect 45422 29376 45481 29410
rect 44787 29372 45481 29376
rect 44787 29338 44860 29372
rect 44894 29338 44960 29372
rect 44994 29338 45060 29372
rect 45094 29338 45160 29372
rect 45194 29338 45260 29372
rect 45294 29338 45360 29372
rect 45394 29338 45481 29372
rect 44787 29320 45481 29338
rect 44787 29286 44848 29320
rect 44882 29286 44938 29320
rect 44972 29286 45028 29320
rect 45062 29286 45118 29320
rect 45152 29286 45208 29320
rect 45242 29286 45298 29320
rect 45332 29286 45388 29320
rect 45422 29286 45481 29320
rect 44787 29272 45481 29286
rect 44787 29238 44860 29272
rect 44894 29238 44960 29272
rect 44994 29238 45060 29272
rect 45094 29238 45160 29272
rect 45194 29238 45260 29272
rect 45294 29238 45360 29272
rect 45394 29238 45481 29272
rect 44787 29230 45481 29238
rect 44787 29196 44848 29230
rect 44882 29196 44938 29230
rect 44972 29196 45028 29230
rect 45062 29196 45118 29230
rect 45152 29196 45208 29230
rect 45242 29196 45298 29230
rect 45332 29196 45388 29230
rect 45422 29196 45481 29230
rect 44787 29172 45481 29196
rect 44787 29140 44860 29172
rect 44894 29140 44960 29172
rect 44994 29140 45060 29172
rect 45094 29140 45160 29172
rect 44787 29106 44848 29140
rect 44894 29138 44938 29140
rect 44994 29138 45028 29140
rect 45094 29138 45118 29140
rect 44882 29106 44938 29138
rect 44972 29106 45028 29138
rect 45062 29106 45118 29138
rect 45152 29138 45160 29140
rect 45194 29140 45260 29172
rect 45194 29138 45208 29140
rect 45152 29106 45208 29138
rect 45242 29138 45260 29140
rect 45294 29140 45360 29172
rect 45394 29140 45481 29172
rect 45294 29138 45298 29140
rect 45242 29106 45298 29138
rect 45332 29138 45360 29140
rect 45332 29106 45388 29138
rect 45422 29106 45481 29140
rect 44787 29072 45481 29106
rect 44787 29050 44860 29072
rect 44894 29050 44960 29072
rect 44994 29050 45060 29072
rect 45094 29050 45160 29072
rect 44787 29016 44848 29050
rect 44894 29038 44938 29050
rect 44994 29038 45028 29050
rect 45094 29038 45118 29050
rect 44882 29016 44938 29038
rect 44972 29016 45028 29038
rect 45062 29016 45118 29038
rect 45152 29038 45160 29050
rect 45194 29050 45260 29072
rect 45194 29038 45208 29050
rect 45152 29016 45208 29038
rect 45242 29038 45260 29050
rect 45294 29050 45360 29072
rect 45394 29050 45481 29072
rect 45294 29038 45298 29050
rect 45242 29016 45298 29038
rect 45332 29038 45360 29050
rect 45332 29016 45388 29038
rect 45422 29016 45481 29050
rect 44787 28972 45481 29016
rect 44787 28960 44860 28972
rect 44894 28960 44960 28972
rect 44994 28960 45060 28972
rect 45094 28960 45160 28972
rect 44787 28926 44848 28960
rect 44894 28938 44938 28960
rect 44994 28938 45028 28960
rect 45094 28938 45118 28960
rect 44882 28926 44938 28938
rect 44972 28926 45028 28938
rect 45062 28926 45118 28938
rect 45152 28938 45160 28960
rect 45194 28960 45260 28972
rect 45194 28938 45208 28960
rect 45152 28926 45208 28938
rect 45242 28938 45260 28960
rect 45294 28960 45360 28972
rect 45394 28960 45481 28972
rect 45294 28938 45298 28960
rect 45242 28926 45298 28938
rect 45332 28938 45360 28960
rect 45332 28926 45388 28938
rect 45422 28926 45481 28960
rect 44787 28865 45481 28926
rect 45543 29508 45615 29564
rect 45543 29474 45562 29508
rect 45596 29474 45615 29508
rect 45543 29418 45615 29474
rect 45543 29384 45562 29418
rect 45596 29384 45615 29418
rect 45543 29328 45615 29384
rect 45543 29294 45562 29328
rect 45596 29294 45615 29328
rect 45543 29238 45615 29294
rect 45543 29204 45562 29238
rect 45596 29204 45615 29238
rect 45543 29148 45615 29204
rect 45543 29114 45562 29148
rect 45596 29114 45615 29148
rect 45543 29058 45615 29114
rect 45543 29024 45562 29058
rect 45596 29024 45615 29058
rect 45543 28968 45615 29024
rect 45543 28934 45562 28968
rect 45596 28934 45615 28968
rect 45543 28878 45615 28934
rect 44653 28803 44725 28863
rect 45543 28844 45562 28878
rect 45596 28844 45615 28878
rect 45543 28803 45615 28844
rect 44653 28784 45615 28803
rect 44653 28750 44750 28784
rect 44784 28750 44840 28784
rect 44874 28750 44930 28784
rect 44964 28750 45020 28784
rect 45054 28750 45110 28784
rect 45144 28750 45200 28784
rect 45234 28750 45290 28784
rect 45324 28750 45380 28784
rect 45414 28750 45470 28784
rect 45504 28750 45615 28784
rect 44653 28731 45615 28750
rect 45679 29674 45711 29708
rect 45745 29674 45864 29708
rect 45898 29674 45929 29708
rect 47019 29708 47269 29757
rect 45679 29618 45929 29674
rect 45679 29584 45711 29618
rect 45745 29584 45864 29618
rect 45898 29584 45929 29618
rect 45679 29528 45929 29584
rect 45679 29494 45711 29528
rect 45745 29494 45864 29528
rect 45898 29494 45929 29528
rect 45679 29438 45929 29494
rect 45679 29404 45711 29438
rect 45745 29404 45864 29438
rect 45898 29404 45929 29438
rect 45679 29348 45929 29404
rect 45679 29314 45711 29348
rect 45745 29314 45864 29348
rect 45898 29314 45929 29348
rect 45679 29258 45929 29314
rect 45679 29224 45711 29258
rect 45745 29224 45864 29258
rect 45898 29224 45929 29258
rect 45679 29168 45929 29224
rect 45679 29134 45711 29168
rect 45745 29134 45864 29168
rect 45898 29134 45929 29168
rect 45679 29078 45929 29134
rect 45679 29044 45711 29078
rect 45745 29044 45864 29078
rect 45898 29044 45929 29078
rect 45679 28988 45929 29044
rect 45679 28954 45711 28988
rect 45745 28954 45864 28988
rect 45898 28954 45929 28988
rect 45679 28898 45929 28954
rect 45679 28864 45711 28898
rect 45745 28864 45864 28898
rect 45898 28864 45929 28898
rect 45679 28808 45929 28864
rect 45679 28774 45711 28808
rect 45745 28774 45864 28808
rect 45898 28774 45929 28808
rect 44339 28684 44371 28718
rect 44405 28684 44524 28718
rect 44558 28684 44589 28718
rect 44339 28667 44589 28684
rect 45679 28718 45929 28774
rect 45993 29676 46955 29693
rect 45993 29642 46014 29676
rect 46048 29642 46104 29676
rect 46138 29674 46194 29676
rect 46228 29674 46284 29676
rect 46318 29674 46374 29676
rect 46408 29674 46464 29676
rect 46498 29674 46554 29676
rect 46588 29674 46644 29676
rect 46678 29674 46734 29676
rect 46768 29674 46824 29676
rect 46858 29674 46914 29676
rect 46158 29642 46194 29674
rect 46248 29642 46284 29674
rect 46338 29642 46374 29674
rect 46428 29642 46464 29674
rect 46518 29642 46554 29674
rect 46608 29642 46644 29674
rect 46698 29642 46734 29674
rect 46788 29642 46824 29674
rect 46878 29642 46914 29674
rect 46948 29642 46955 29676
rect 45993 29640 46124 29642
rect 46158 29640 46214 29642
rect 46248 29640 46304 29642
rect 46338 29640 46394 29642
rect 46428 29640 46484 29642
rect 46518 29640 46574 29642
rect 46608 29640 46664 29642
rect 46698 29640 46754 29642
rect 46788 29640 46844 29642
rect 46878 29640 46955 29642
rect 45993 29621 46955 29640
rect 45993 29617 46065 29621
rect 45993 29583 46012 29617
rect 46046 29583 46065 29617
rect 45993 29527 46065 29583
rect 46883 29598 46955 29621
rect 46883 29564 46902 29598
rect 46936 29564 46955 29598
rect 45993 29493 46012 29527
rect 46046 29493 46065 29527
rect 45993 29437 46065 29493
rect 45993 29403 46012 29437
rect 46046 29403 46065 29437
rect 45993 29347 46065 29403
rect 45993 29313 46012 29347
rect 46046 29313 46065 29347
rect 45993 29257 46065 29313
rect 45993 29223 46012 29257
rect 46046 29223 46065 29257
rect 45993 29167 46065 29223
rect 45993 29133 46012 29167
rect 46046 29133 46065 29167
rect 45993 29077 46065 29133
rect 45993 29043 46012 29077
rect 46046 29043 46065 29077
rect 45993 28987 46065 29043
rect 45993 28953 46012 28987
rect 46046 28953 46065 28987
rect 45993 28897 46065 28953
rect 45993 28863 46012 28897
rect 46046 28863 46065 28897
rect 46127 29500 46821 29559
rect 46127 29466 46188 29500
rect 46222 29472 46278 29500
rect 46312 29472 46368 29500
rect 46402 29472 46458 29500
rect 46234 29466 46278 29472
rect 46334 29466 46368 29472
rect 46434 29466 46458 29472
rect 46492 29472 46548 29500
rect 46492 29466 46500 29472
rect 46127 29438 46200 29466
rect 46234 29438 46300 29466
rect 46334 29438 46400 29466
rect 46434 29438 46500 29466
rect 46534 29466 46548 29472
rect 46582 29472 46638 29500
rect 46582 29466 46600 29472
rect 46534 29438 46600 29466
rect 46634 29466 46638 29472
rect 46672 29472 46728 29500
rect 46672 29466 46700 29472
rect 46762 29466 46821 29500
rect 46634 29438 46700 29466
rect 46734 29438 46821 29466
rect 46127 29410 46821 29438
rect 46127 29376 46188 29410
rect 46222 29376 46278 29410
rect 46312 29376 46368 29410
rect 46402 29376 46458 29410
rect 46492 29376 46548 29410
rect 46582 29376 46638 29410
rect 46672 29376 46728 29410
rect 46762 29376 46821 29410
rect 46127 29372 46821 29376
rect 46127 29338 46200 29372
rect 46234 29338 46300 29372
rect 46334 29338 46400 29372
rect 46434 29338 46500 29372
rect 46534 29338 46600 29372
rect 46634 29338 46700 29372
rect 46734 29338 46821 29372
rect 46127 29320 46821 29338
rect 46127 29286 46188 29320
rect 46222 29286 46278 29320
rect 46312 29286 46368 29320
rect 46402 29286 46458 29320
rect 46492 29286 46548 29320
rect 46582 29286 46638 29320
rect 46672 29286 46728 29320
rect 46762 29286 46821 29320
rect 46127 29272 46821 29286
rect 46127 29238 46200 29272
rect 46234 29238 46300 29272
rect 46334 29238 46400 29272
rect 46434 29238 46500 29272
rect 46534 29238 46600 29272
rect 46634 29238 46700 29272
rect 46734 29238 46821 29272
rect 46127 29230 46821 29238
rect 46127 29196 46188 29230
rect 46222 29196 46278 29230
rect 46312 29196 46368 29230
rect 46402 29196 46458 29230
rect 46492 29196 46548 29230
rect 46582 29196 46638 29230
rect 46672 29196 46728 29230
rect 46762 29196 46821 29230
rect 46127 29172 46821 29196
rect 46127 29140 46200 29172
rect 46234 29140 46300 29172
rect 46334 29140 46400 29172
rect 46434 29140 46500 29172
rect 46127 29106 46188 29140
rect 46234 29138 46278 29140
rect 46334 29138 46368 29140
rect 46434 29138 46458 29140
rect 46222 29106 46278 29138
rect 46312 29106 46368 29138
rect 46402 29106 46458 29138
rect 46492 29138 46500 29140
rect 46534 29140 46600 29172
rect 46534 29138 46548 29140
rect 46492 29106 46548 29138
rect 46582 29138 46600 29140
rect 46634 29140 46700 29172
rect 46734 29140 46821 29172
rect 46634 29138 46638 29140
rect 46582 29106 46638 29138
rect 46672 29138 46700 29140
rect 46672 29106 46728 29138
rect 46762 29106 46821 29140
rect 46127 29072 46821 29106
rect 46127 29050 46200 29072
rect 46234 29050 46300 29072
rect 46334 29050 46400 29072
rect 46434 29050 46500 29072
rect 46127 29016 46188 29050
rect 46234 29038 46278 29050
rect 46334 29038 46368 29050
rect 46434 29038 46458 29050
rect 46222 29016 46278 29038
rect 46312 29016 46368 29038
rect 46402 29016 46458 29038
rect 46492 29038 46500 29050
rect 46534 29050 46600 29072
rect 46534 29038 46548 29050
rect 46492 29016 46548 29038
rect 46582 29038 46600 29050
rect 46634 29050 46700 29072
rect 46734 29050 46821 29072
rect 46634 29038 46638 29050
rect 46582 29016 46638 29038
rect 46672 29038 46700 29050
rect 46672 29016 46728 29038
rect 46762 29016 46821 29050
rect 46127 28972 46821 29016
rect 46127 28960 46200 28972
rect 46234 28960 46300 28972
rect 46334 28960 46400 28972
rect 46434 28960 46500 28972
rect 46127 28926 46188 28960
rect 46234 28938 46278 28960
rect 46334 28938 46368 28960
rect 46434 28938 46458 28960
rect 46222 28926 46278 28938
rect 46312 28926 46368 28938
rect 46402 28926 46458 28938
rect 46492 28938 46500 28960
rect 46534 28960 46600 28972
rect 46534 28938 46548 28960
rect 46492 28926 46548 28938
rect 46582 28938 46600 28960
rect 46634 28960 46700 28972
rect 46734 28960 46821 28972
rect 46634 28938 46638 28960
rect 46582 28926 46638 28938
rect 46672 28938 46700 28960
rect 46672 28926 46728 28938
rect 46762 28926 46821 28960
rect 46127 28865 46821 28926
rect 46883 29508 46955 29564
rect 46883 29474 46902 29508
rect 46936 29474 46955 29508
rect 46883 29418 46955 29474
rect 46883 29384 46902 29418
rect 46936 29384 46955 29418
rect 46883 29328 46955 29384
rect 46883 29294 46902 29328
rect 46936 29294 46955 29328
rect 46883 29238 46955 29294
rect 46883 29204 46902 29238
rect 46936 29204 46955 29238
rect 46883 29148 46955 29204
rect 46883 29114 46902 29148
rect 46936 29114 46955 29148
rect 46883 29058 46955 29114
rect 46883 29024 46902 29058
rect 46936 29024 46955 29058
rect 46883 28968 46955 29024
rect 46883 28934 46902 28968
rect 46936 28934 46955 28968
rect 46883 28878 46955 28934
rect 45993 28803 46065 28863
rect 46883 28844 46902 28878
rect 46936 28844 46955 28878
rect 46883 28803 46955 28844
rect 45993 28784 46955 28803
rect 45993 28750 46090 28784
rect 46124 28750 46180 28784
rect 46214 28750 46270 28784
rect 46304 28750 46360 28784
rect 46394 28750 46450 28784
rect 46484 28750 46540 28784
rect 46574 28750 46630 28784
rect 46664 28750 46720 28784
rect 46754 28750 46810 28784
rect 46844 28750 46955 28784
rect 45993 28731 46955 28750
rect 47019 29674 47051 29708
rect 47085 29674 47204 29708
rect 47238 29674 47269 29708
rect 48359 29708 48609 29757
rect 47019 29618 47269 29674
rect 47019 29584 47051 29618
rect 47085 29584 47204 29618
rect 47238 29584 47269 29618
rect 47019 29528 47269 29584
rect 47019 29494 47051 29528
rect 47085 29494 47204 29528
rect 47238 29494 47269 29528
rect 47019 29438 47269 29494
rect 47019 29404 47051 29438
rect 47085 29404 47204 29438
rect 47238 29404 47269 29438
rect 47019 29348 47269 29404
rect 47019 29314 47051 29348
rect 47085 29314 47204 29348
rect 47238 29314 47269 29348
rect 47019 29258 47269 29314
rect 47019 29224 47051 29258
rect 47085 29224 47204 29258
rect 47238 29224 47269 29258
rect 47019 29168 47269 29224
rect 47019 29134 47051 29168
rect 47085 29134 47204 29168
rect 47238 29134 47269 29168
rect 47019 29078 47269 29134
rect 47019 29044 47051 29078
rect 47085 29044 47204 29078
rect 47238 29044 47269 29078
rect 47019 28988 47269 29044
rect 47019 28954 47051 28988
rect 47085 28954 47204 28988
rect 47238 28954 47269 28988
rect 47019 28898 47269 28954
rect 47019 28864 47051 28898
rect 47085 28864 47204 28898
rect 47238 28864 47269 28898
rect 47019 28808 47269 28864
rect 47019 28774 47051 28808
rect 47085 28774 47204 28808
rect 47238 28774 47269 28808
rect 45679 28684 45711 28718
rect 45745 28684 45864 28718
rect 45898 28684 45929 28718
rect 45679 28667 45929 28684
rect 47019 28718 47269 28774
rect 47333 29676 48295 29693
rect 47333 29642 47354 29676
rect 47388 29642 47444 29676
rect 47478 29674 47534 29676
rect 47568 29674 47624 29676
rect 47658 29674 47714 29676
rect 47748 29674 47804 29676
rect 47838 29674 47894 29676
rect 47928 29674 47984 29676
rect 48018 29674 48074 29676
rect 48108 29674 48164 29676
rect 48198 29674 48254 29676
rect 47498 29642 47534 29674
rect 47588 29642 47624 29674
rect 47678 29642 47714 29674
rect 47768 29642 47804 29674
rect 47858 29642 47894 29674
rect 47948 29642 47984 29674
rect 48038 29642 48074 29674
rect 48128 29642 48164 29674
rect 48218 29642 48254 29674
rect 48288 29642 48295 29676
rect 47333 29640 47464 29642
rect 47498 29640 47554 29642
rect 47588 29640 47644 29642
rect 47678 29640 47734 29642
rect 47768 29640 47824 29642
rect 47858 29640 47914 29642
rect 47948 29640 48004 29642
rect 48038 29640 48094 29642
rect 48128 29640 48184 29642
rect 48218 29640 48295 29642
rect 47333 29621 48295 29640
rect 47333 29617 47405 29621
rect 47333 29583 47352 29617
rect 47386 29583 47405 29617
rect 47333 29527 47405 29583
rect 48223 29598 48295 29621
rect 48223 29564 48242 29598
rect 48276 29564 48295 29598
rect 47333 29493 47352 29527
rect 47386 29493 47405 29527
rect 47333 29437 47405 29493
rect 47333 29403 47352 29437
rect 47386 29403 47405 29437
rect 47333 29347 47405 29403
rect 47333 29313 47352 29347
rect 47386 29313 47405 29347
rect 47333 29257 47405 29313
rect 47333 29223 47352 29257
rect 47386 29223 47405 29257
rect 47333 29167 47405 29223
rect 47333 29133 47352 29167
rect 47386 29133 47405 29167
rect 47333 29077 47405 29133
rect 47333 29043 47352 29077
rect 47386 29043 47405 29077
rect 47333 28987 47405 29043
rect 47333 28953 47352 28987
rect 47386 28953 47405 28987
rect 47333 28897 47405 28953
rect 47333 28863 47352 28897
rect 47386 28863 47405 28897
rect 47467 29500 48161 29559
rect 47467 29466 47528 29500
rect 47562 29472 47618 29500
rect 47652 29472 47708 29500
rect 47742 29472 47798 29500
rect 47574 29466 47618 29472
rect 47674 29466 47708 29472
rect 47774 29466 47798 29472
rect 47832 29472 47888 29500
rect 47832 29466 47840 29472
rect 47467 29438 47540 29466
rect 47574 29438 47640 29466
rect 47674 29438 47740 29466
rect 47774 29438 47840 29466
rect 47874 29466 47888 29472
rect 47922 29472 47978 29500
rect 47922 29466 47940 29472
rect 47874 29438 47940 29466
rect 47974 29466 47978 29472
rect 48012 29472 48068 29500
rect 48012 29466 48040 29472
rect 48102 29466 48161 29500
rect 47974 29438 48040 29466
rect 48074 29438 48161 29466
rect 47467 29410 48161 29438
rect 47467 29376 47528 29410
rect 47562 29376 47618 29410
rect 47652 29376 47708 29410
rect 47742 29376 47798 29410
rect 47832 29376 47888 29410
rect 47922 29376 47978 29410
rect 48012 29376 48068 29410
rect 48102 29376 48161 29410
rect 47467 29372 48161 29376
rect 47467 29338 47540 29372
rect 47574 29338 47640 29372
rect 47674 29338 47740 29372
rect 47774 29338 47840 29372
rect 47874 29338 47940 29372
rect 47974 29338 48040 29372
rect 48074 29338 48161 29372
rect 47467 29320 48161 29338
rect 47467 29286 47528 29320
rect 47562 29286 47618 29320
rect 47652 29286 47708 29320
rect 47742 29286 47798 29320
rect 47832 29286 47888 29320
rect 47922 29286 47978 29320
rect 48012 29286 48068 29320
rect 48102 29286 48161 29320
rect 47467 29272 48161 29286
rect 47467 29238 47540 29272
rect 47574 29238 47640 29272
rect 47674 29238 47740 29272
rect 47774 29238 47840 29272
rect 47874 29238 47940 29272
rect 47974 29238 48040 29272
rect 48074 29238 48161 29272
rect 47467 29230 48161 29238
rect 47467 29196 47528 29230
rect 47562 29196 47618 29230
rect 47652 29196 47708 29230
rect 47742 29196 47798 29230
rect 47832 29196 47888 29230
rect 47922 29196 47978 29230
rect 48012 29196 48068 29230
rect 48102 29196 48161 29230
rect 47467 29172 48161 29196
rect 47467 29140 47540 29172
rect 47574 29140 47640 29172
rect 47674 29140 47740 29172
rect 47774 29140 47840 29172
rect 47467 29106 47528 29140
rect 47574 29138 47618 29140
rect 47674 29138 47708 29140
rect 47774 29138 47798 29140
rect 47562 29106 47618 29138
rect 47652 29106 47708 29138
rect 47742 29106 47798 29138
rect 47832 29138 47840 29140
rect 47874 29140 47940 29172
rect 47874 29138 47888 29140
rect 47832 29106 47888 29138
rect 47922 29138 47940 29140
rect 47974 29140 48040 29172
rect 48074 29140 48161 29172
rect 47974 29138 47978 29140
rect 47922 29106 47978 29138
rect 48012 29138 48040 29140
rect 48012 29106 48068 29138
rect 48102 29106 48161 29140
rect 47467 29072 48161 29106
rect 47467 29050 47540 29072
rect 47574 29050 47640 29072
rect 47674 29050 47740 29072
rect 47774 29050 47840 29072
rect 47467 29016 47528 29050
rect 47574 29038 47618 29050
rect 47674 29038 47708 29050
rect 47774 29038 47798 29050
rect 47562 29016 47618 29038
rect 47652 29016 47708 29038
rect 47742 29016 47798 29038
rect 47832 29038 47840 29050
rect 47874 29050 47940 29072
rect 47874 29038 47888 29050
rect 47832 29016 47888 29038
rect 47922 29038 47940 29050
rect 47974 29050 48040 29072
rect 48074 29050 48161 29072
rect 47974 29038 47978 29050
rect 47922 29016 47978 29038
rect 48012 29038 48040 29050
rect 48012 29016 48068 29038
rect 48102 29016 48161 29050
rect 47467 28972 48161 29016
rect 47467 28960 47540 28972
rect 47574 28960 47640 28972
rect 47674 28960 47740 28972
rect 47774 28960 47840 28972
rect 47467 28926 47528 28960
rect 47574 28938 47618 28960
rect 47674 28938 47708 28960
rect 47774 28938 47798 28960
rect 47562 28926 47618 28938
rect 47652 28926 47708 28938
rect 47742 28926 47798 28938
rect 47832 28938 47840 28960
rect 47874 28960 47940 28972
rect 47874 28938 47888 28960
rect 47832 28926 47888 28938
rect 47922 28938 47940 28960
rect 47974 28960 48040 28972
rect 48074 28960 48161 28972
rect 47974 28938 47978 28960
rect 47922 28926 47978 28938
rect 48012 28938 48040 28960
rect 48012 28926 48068 28938
rect 48102 28926 48161 28960
rect 47467 28865 48161 28926
rect 48223 29508 48295 29564
rect 48223 29474 48242 29508
rect 48276 29474 48295 29508
rect 48223 29418 48295 29474
rect 48223 29384 48242 29418
rect 48276 29384 48295 29418
rect 48223 29328 48295 29384
rect 48223 29294 48242 29328
rect 48276 29294 48295 29328
rect 48223 29238 48295 29294
rect 48223 29204 48242 29238
rect 48276 29204 48295 29238
rect 48223 29148 48295 29204
rect 48223 29114 48242 29148
rect 48276 29114 48295 29148
rect 48223 29058 48295 29114
rect 48223 29024 48242 29058
rect 48276 29024 48295 29058
rect 48223 28968 48295 29024
rect 48223 28934 48242 28968
rect 48276 28934 48295 28968
rect 48223 28878 48295 28934
rect 47333 28803 47405 28863
rect 48223 28844 48242 28878
rect 48276 28844 48295 28878
rect 48223 28803 48295 28844
rect 47333 28784 48295 28803
rect 47333 28750 47430 28784
rect 47464 28750 47520 28784
rect 47554 28750 47610 28784
rect 47644 28750 47700 28784
rect 47734 28750 47790 28784
rect 47824 28750 47880 28784
rect 47914 28750 47970 28784
rect 48004 28750 48060 28784
rect 48094 28750 48150 28784
rect 48184 28750 48295 28784
rect 47333 28731 48295 28750
rect 48359 29674 48391 29708
rect 48425 29674 48544 29708
rect 48578 29674 48609 29708
rect 49699 29708 49949 29757
rect 48359 29618 48609 29674
rect 48359 29584 48391 29618
rect 48425 29584 48544 29618
rect 48578 29584 48609 29618
rect 48359 29528 48609 29584
rect 48359 29494 48391 29528
rect 48425 29494 48544 29528
rect 48578 29494 48609 29528
rect 48359 29438 48609 29494
rect 48359 29404 48391 29438
rect 48425 29404 48544 29438
rect 48578 29404 48609 29438
rect 48359 29348 48609 29404
rect 48359 29314 48391 29348
rect 48425 29314 48544 29348
rect 48578 29314 48609 29348
rect 48359 29258 48609 29314
rect 48359 29224 48391 29258
rect 48425 29224 48544 29258
rect 48578 29224 48609 29258
rect 48359 29168 48609 29224
rect 48359 29134 48391 29168
rect 48425 29134 48544 29168
rect 48578 29134 48609 29168
rect 48359 29078 48609 29134
rect 48359 29044 48391 29078
rect 48425 29044 48544 29078
rect 48578 29044 48609 29078
rect 48359 28988 48609 29044
rect 48359 28954 48391 28988
rect 48425 28954 48544 28988
rect 48578 28954 48609 28988
rect 48359 28898 48609 28954
rect 48359 28864 48391 28898
rect 48425 28864 48544 28898
rect 48578 28864 48609 28898
rect 48359 28808 48609 28864
rect 48359 28774 48391 28808
rect 48425 28774 48544 28808
rect 48578 28774 48609 28808
rect 47019 28684 47051 28718
rect 47085 28684 47204 28718
rect 47238 28684 47269 28718
rect 47019 28667 47269 28684
rect 48359 28718 48609 28774
rect 48673 29676 49635 29693
rect 48673 29642 48694 29676
rect 48728 29642 48784 29676
rect 48818 29674 48874 29676
rect 48908 29674 48964 29676
rect 48998 29674 49054 29676
rect 49088 29674 49144 29676
rect 49178 29674 49234 29676
rect 49268 29674 49324 29676
rect 49358 29674 49414 29676
rect 49448 29674 49504 29676
rect 49538 29674 49594 29676
rect 48838 29642 48874 29674
rect 48928 29642 48964 29674
rect 49018 29642 49054 29674
rect 49108 29642 49144 29674
rect 49198 29642 49234 29674
rect 49288 29642 49324 29674
rect 49378 29642 49414 29674
rect 49468 29642 49504 29674
rect 49558 29642 49594 29674
rect 49628 29642 49635 29676
rect 48673 29640 48804 29642
rect 48838 29640 48894 29642
rect 48928 29640 48984 29642
rect 49018 29640 49074 29642
rect 49108 29640 49164 29642
rect 49198 29640 49254 29642
rect 49288 29640 49344 29642
rect 49378 29640 49434 29642
rect 49468 29640 49524 29642
rect 49558 29640 49635 29642
rect 48673 29621 49635 29640
rect 48673 29617 48745 29621
rect 48673 29583 48692 29617
rect 48726 29583 48745 29617
rect 48673 29527 48745 29583
rect 49563 29598 49635 29621
rect 49563 29564 49582 29598
rect 49616 29564 49635 29598
rect 48673 29493 48692 29527
rect 48726 29493 48745 29527
rect 48673 29437 48745 29493
rect 48673 29403 48692 29437
rect 48726 29403 48745 29437
rect 48673 29347 48745 29403
rect 48673 29313 48692 29347
rect 48726 29313 48745 29347
rect 48673 29257 48745 29313
rect 48673 29223 48692 29257
rect 48726 29223 48745 29257
rect 48673 29167 48745 29223
rect 48673 29133 48692 29167
rect 48726 29133 48745 29167
rect 48673 29077 48745 29133
rect 48673 29043 48692 29077
rect 48726 29043 48745 29077
rect 48673 28987 48745 29043
rect 48673 28953 48692 28987
rect 48726 28953 48745 28987
rect 48673 28897 48745 28953
rect 48673 28863 48692 28897
rect 48726 28863 48745 28897
rect 48807 29500 49501 29559
rect 48807 29466 48868 29500
rect 48902 29472 48958 29500
rect 48992 29472 49048 29500
rect 49082 29472 49138 29500
rect 48914 29466 48958 29472
rect 49014 29466 49048 29472
rect 49114 29466 49138 29472
rect 49172 29472 49228 29500
rect 49172 29466 49180 29472
rect 48807 29438 48880 29466
rect 48914 29438 48980 29466
rect 49014 29438 49080 29466
rect 49114 29438 49180 29466
rect 49214 29466 49228 29472
rect 49262 29472 49318 29500
rect 49262 29466 49280 29472
rect 49214 29438 49280 29466
rect 49314 29466 49318 29472
rect 49352 29472 49408 29500
rect 49352 29466 49380 29472
rect 49442 29466 49501 29500
rect 49314 29438 49380 29466
rect 49414 29438 49501 29466
rect 48807 29410 49501 29438
rect 48807 29376 48868 29410
rect 48902 29376 48958 29410
rect 48992 29376 49048 29410
rect 49082 29376 49138 29410
rect 49172 29376 49228 29410
rect 49262 29376 49318 29410
rect 49352 29376 49408 29410
rect 49442 29376 49501 29410
rect 48807 29372 49501 29376
rect 48807 29338 48880 29372
rect 48914 29338 48980 29372
rect 49014 29338 49080 29372
rect 49114 29338 49180 29372
rect 49214 29338 49280 29372
rect 49314 29338 49380 29372
rect 49414 29338 49501 29372
rect 48807 29320 49501 29338
rect 48807 29286 48868 29320
rect 48902 29286 48958 29320
rect 48992 29286 49048 29320
rect 49082 29286 49138 29320
rect 49172 29286 49228 29320
rect 49262 29286 49318 29320
rect 49352 29286 49408 29320
rect 49442 29286 49501 29320
rect 48807 29272 49501 29286
rect 48807 29238 48880 29272
rect 48914 29238 48980 29272
rect 49014 29238 49080 29272
rect 49114 29238 49180 29272
rect 49214 29238 49280 29272
rect 49314 29238 49380 29272
rect 49414 29238 49501 29272
rect 48807 29230 49501 29238
rect 48807 29196 48868 29230
rect 48902 29196 48958 29230
rect 48992 29196 49048 29230
rect 49082 29196 49138 29230
rect 49172 29196 49228 29230
rect 49262 29196 49318 29230
rect 49352 29196 49408 29230
rect 49442 29196 49501 29230
rect 48807 29172 49501 29196
rect 48807 29140 48880 29172
rect 48914 29140 48980 29172
rect 49014 29140 49080 29172
rect 49114 29140 49180 29172
rect 48807 29106 48868 29140
rect 48914 29138 48958 29140
rect 49014 29138 49048 29140
rect 49114 29138 49138 29140
rect 48902 29106 48958 29138
rect 48992 29106 49048 29138
rect 49082 29106 49138 29138
rect 49172 29138 49180 29140
rect 49214 29140 49280 29172
rect 49214 29138 49228 29140
rect 49172 29106 49228 29138
rect 49262 29138 49280 29140
rect 49314 29140 49380 29172
rect 49414 29140 49501 29172
rect 49314 29138 49318 29140
rect 49262 29106 49318 29138
rect 49352 29138 49380 29140
rect 49352 29106 49408 29138
rect 49442 29106 49501 29140
rect 48807 29072 49501 29106
rect 48807 29050 48880 29072
rect 48914 29050 48980 29072
rect 49014 29050 49080 29072
rect 49114 29050 49180 29072
rect 48807 29016 48868 29050
rect 48914 29038 48958 29050
rect 49014 29038 49048 29050
rect 49114 29038 49138 29050
rect 48902 29016 48958 29038
rect 48992 29016 49048 29038
rect 49082 29016 49138 29038
rect 49172 29038 49180 29050
rect 49214 29050 49280 29072
rect 49214 29038 49228 29050
rect 49172 29016 49228 29038
rect 49262 29038 49280 29050
rect 49314 29050 49380 29072
rect 49414 29050 49501 29072
rect 49314 29038 49318 29050
rect 49262 29016 49318 29038
rect 49352 29038 49380 29050
rect 49352 29016 49408 29038
rect 49442 29016 49501 29050
rect 48807 28972 49501 29016
rect 48807 28960 48880 28972
rect 48914 28960 48980 28972
rect 49014 28960 49080 28972
rect 49114 28960 49180 28972
rect 48807 28926 48868 28960
rect 48914 28938 48958 28960
rect 49014 28938 49048 28960
rect 49114 28938 49138 28960
rect 48902 28926 48958 28938
rect 48992 28926 49048 28938
rect 49082 28926 49138 28938
rect 49172 28938 49180 28960
rect 49214 28960 49280 28972
rect 49214 28938 49228 28960
rect 49172 28926 49228 28938
rect 49262 28938 49280 28960
rect 49314 28960 49380 28972
rect 49414 28960 49501 28972
rect 49314 28938 49318 28960
rect 49262 28926 49318 28938
rect 49352 28938 49380 28960
rect 49352 28926 49408 28938
rect 49442 28926 49501 28960
rect 48807 28865 49501 28926
rect 49563 29508 49635 29564
rect 49563 29474 49582 29508
rect 49616 29474 49635 29508
rect 49563 29418 49635 29474
rect 49563 29384 49582 29418
rect 49616 29384 49635 29418
rect 49563 29328 49635 29384
rect 49563 29294 49582 29328
rect 49616 29294 49635 29328
rect 49563 29238 49635 29294
rect 49563 29204 49582 29238
rect 49616 29204 49635 29238
rect 49563 29148 49635 29204
rect 49563 29114 49582 29148
rect 49616 29114 49635 29148
rect 49563 29058 49635 29114
rect 49563 29024 49582 29058
rect 49616 29024 49635 29058
rect 49563 28968 49635 29024
rect 49563 28934 49582 28968
rect 49616 28934 49635 28968
rect 49563 28878 49635 28934
rect 48673 28803 48745 28863
rect 49563 28844 49582 28878
rect 49616 28844 49635 28878
rect 49563 28803 49635 28844
rect 48673 28784 49635 28803
rect 48673 28750 48770 28784
rect 48804 28750 48860 28784
rect 48894 28750 48950 28784
rect 48984 28750 49040 28784
rect 49074 28750 49130 28784
rect 49164 28750 49220 28784
rect 49254 28750 49310 28784
rect 49344 28750 49400 28784
rect 49434 28750 49490 28784
rect 49524 28750 49635 28784
rect 48673 28731 49635 28750
rect 49699 29674 49731 29708
rect 49765 29674 49884 29708
rect 49918 29674 49949 29708
rect 51039 29708 51289 29757
rect 49699 29618 49949 29674
rect 49699 29584 49731 29618
rect 49765 29584 49884 29618
rect 49918 29584 49949 29618
rect 49699 29528 49949 29584
rect 49699 29494 49731 29528
rect 49765 29494 49884 29528
rect 49918 29494 49949 29528
rect 49699 29438 49949 29494
rect 49699 29404 49731 29438
rect 49765 29404 49884 29438
rect 49918 29404 49949 29438
rect 49699 29348 49949 29404
rect 49699 29314 49731 29348
rect 49765 29314 49884 29348
rect 49918 29314 49949 29348
rect 49699 29258 49949 29314
rect 49699 29224 49731 29258
rect 49765 29224 49884 29258
rect 49918 29224 49949 29258
rect 49699 29168 49949 29224
rect 49699 29134 49731 29168
rect 49765 29134 49884 29168
rect 49918 29134 49949 29168
rect 49699 29078 49949 29134
rect 49699 29044 49731 29078
rect 49765 29044 49884 29078
rect 49918 29044 49949 29078
rect 49699 28988 49949 29044
rect 49699 28954 49731 28988
rect 49765 28954 49884 28988
rect 49918 28954 49949 28988
rect 49699 28898 49949 28954
rect 49699 28864 49731 28898
rect 49765 28864 49884 28898
rect 49918 28864 49949 28898
rect 49699 28808 49949 28864
rect 49699 28774 49731 28808
rect 49765 28774 49884 28808
rect 49918 28774 49949 28808
rect 48359 28684 48391 28718
rect 48425 28684 48544 28718
rect 48578 28684 48609 28718
rect 48359 28667 48609 28684
rect 49699 28718 49949 28774
rect 50013 29676 50975 29693
rect 50013 29642 50034 29676
rect 50068 29642 50124 29676
rect 50158 29674 50214 29676
rect 50248 29674 50304 29676
rect 50338 29674 50394 29676
rect 50428 29674 50484 29676
rect 50518 29674 50574 29676
rect 50608 29674 50664 29676
rect 50698 29674 50754 29676
rect 50788 29674 50844 29676
rect 50878 29674 50934 29676
rect 50178 29642 50214 29674
rect 50268 29642 50304 29674
rect 50358 29642 50394 29674
rect 50448 29642 50484 29674
rect 50538 29642 50574 29674
rect 50628 29642 50664 29674
rect 50718 29642 50754 29674
rect 50808 29642 50844 29674
rect 50898 29642 50934 29674
rect 50968 29642 50975 29676
rect 50013 29640 50144 29642
rect 50178 29640 50234 29642
rect 50268 29640 50324 29642
rect 50358 29640 50414 29642
rect 50448 29640 50504 29642
rect 50538 29640 50594 29642
rect 50628 29640 50684 29642
rect 50718 29640 50774 29642
rect 50808 29640 50864 29642
rect 50898 29640 50975 29642
rect 50013 29621 50975 29640
rect 50013 29617 50085 29621
rect 50013 29583 50032 29617
rect 50066 29583 50085 29617
rect 50013 29527 50085 29583
rect 50903 29598 50975 29621
rect 50903 29564 50922 29598
rect 50956 29564 50975 29598
rect 50013 29493 50032 29527
rect 50066 29493 50085 29527
rect 50013 29437 50085 29493
rect 50013 29403 50032 29437
rect 50066 29403 50085 29437
rect 50013 29347 50085 29403
rect 50013 29313 50032 29347
rect 50066 29313 50085 29347
rect 50013 29257 50085 29313
rect 50013 29223 50032 29257
rect 50066 29223 50085 29257
rect 50013 29167 50085 29223
rect 50013 29133 50032 29167
rect 50066 29133 50085 29167
rect 50013 29077 50085 29133
rect 50013 29043 50032 29077
rect 50066 29043 50085 29077
rect 50013 28987 50085 29043
rect 50013 28953 50032 28987
rect 50066 28953 50085 28987
rect 50013 28897 50085 28953
rect 50013 28863 50032 28897
rect 50066 28863 50085 28897
rect 50147 29500 50841 29559
rect 50147 29466 50208 29500
rect 50242 29472 50298 29500
rect 50332 29472 50388 29500
rect 50422 29472 50478 29500
rect 50254 29466 50298 29472
rect 50354 29466 50388 29472
rect 50454 29466 50478 29472
rect 50512 29472 50568 29500
rect 50512 29466 50520 29472
rect 50147 29438 50220 29466
rect 50254 29438 50320 29466
rect 50354 29438 50420 29466
rect 50454 29438 50520 29466
rect 50554 29466 50568 29472
rect 50602 29472 50658 29500
rect 50602 29466 50620 29472
rect 50554 29438 50620 29466
rect 50654 29466 50658 29472
rect 50692 29472 50748 29500
rect 50692 29466 50720 29472
rect 50782 29466 50841 29500
rect 50654 29438 50720 29466
rect 50754 29438 50841 29466
rect 50147 29410 50841 29438
rect 50147 29376 50208 29410
rect 50242 29376 50298 29410
rect 50332 29376 50388 29410
rect 50422 29376 50478 29410
rect 50512 29376 50568 29410
rect 50602 29376 50658 29410
rect 50692 29376 50748 29410
rect 50782 29376 50841 29410
rect 50147 29372 50841 29376
rect 50147 29338 50220 29372
rect 50254 29338 50320 29372
rect 50354 29338 50420 29372
rect 50454 29338 50520 29372
rect 50554 29338 50620 29372
rect 50654 29338 50720 29372
rect 50754 29338 50841 29372
rect 50147 29320 50841 29338
rect 50147 29286 50208 29320
rect 50242 29286 50298 29320
rect 50332 29286 50388 29320
rect 50422 29286 50478 29320
rect 50512 29286 50568 29320
rect 50602 29286 50658 29320
rect 50692 29286 50748 29320
rect 50782 29286 50841 29320
rect 50147 29272 50841 29286
rect 50147 29238 50220 29272
rect 50254 29238 50320 29272
rect 50354 29238 50420 29272
rect 50454 29238 50520 29272
rect 50554 29238 50620 29272
rect 50654 29238 50720 29272
rect 50754 29238 50841 29272
rect 50147 29230 50841 29238
rect 50147 29196 50208 29230
rect 50242 29196 50298 29230
rect 50332 29196 50388 29230
rect 50422 29196 50478 29230
rect 50512 29196 50568 29230
rect 50602 29196 50658 29230
rect 50692 29196 50748 29230
rect 50782 29196 50841 29230
rect 50147 29172 50841 29196
rect 50147 29140 50220 29172
rect 50254 29140 50320 29172
rect 50354 29140 50420 29172
rect 50454 29140 50520 29172
rect 50147 29106 50208 29140
rect 50254 29138 50298 29140
rect 50354 29138 50388 29140
rect 50454 29138 50478 29140
rect 50242 29106 50298 29138
rect 50332 29106 50388 29138
rect 50422 29106 50478 29138
rect 50512 29138 50520 29140
rect 50554 29140 50620 29172
rect 50554 29138 50568 29140
rect 50512 29106 50568 29138
rect 50602 29138 50620 29140
rect 50654 29140 50720 29172
rect 50754 29140 50841 29172
rect 50654 29138 50658 29140
rect 50602 29106 50658 29138
rect 50692 29138 50720 29140
rect 50692 29106 50748 29138
rect 50782 29106 50841 29140
rect 50147 29072 50841 29106
rect 50147 29050 50220 29072
rect 50254 29050 50320 29072
rect 50354 29050 50420 29072
rect 50454 29050 50520 29072
rect 50147 29016 50208 29050
rect 50254 29038 50298 29050
rect 50354 29038 50388 29050
rect 50454 29038 50478 29050
rect 50242 29016 50298 29038
rect 50332 29016 50388 29038
rect 50422 29016 50478 29038
rect 50512 29038 50520 29050
rect 50554 29050 50620 29072
rect 50554 29038 50568 29050
rect 50512 29016 50568 29038
rect 50602 29038 50620 29050
rect 50654 29050 50720 29072
rect 50754 29050 50841 29072
rect 50654 29038 50658 29050
rect 50602 29016 50658 29038
rect 50692 29038 50720 29050
rect 50692 29016 50748 29038
rect 50782 29016 50841 29050
rect 50147 28972 50841 29016
rect 50147 28960 50220 28972
rect 50254 28960 50320 28972
rect 50354 28960 50420 28972
rect 50454 28960 50520 28972
rect 50147 28926 50208 28960
rect 50254 28938 50298 28960
rect 50354 28938 50388 28960
rect 50454 28938 50478 28960
rect 50242 28926 50298 28938
rect 50332 28926 50388 28938
rect 50422 28926 50478 28938
rect 50512 28938 50520 28960
rect 50554 28960 50620 28972
rect 50554 28938 50568 28960
rect 50512 28926 50568 28938
rect 50602 28938 50620 28960
rect 50654 28960 50720 28972
rect 50754 28960 50841 28972
rect 50654 28938 50658 28960
rect 50602 28926 50658 28938
rect 50692 28938 50720 28960
rect 50692 28926 50748 28938
rect 50782 28926 50841 28960
rect 50147 28865 50841 28926
rect 50903 29508 50975 29564
rect 50903 29474 50922 29508
rect 50956 29474 50975 29508
rect 50903 29418 50975 29474
rect 50903 29384 50922 29418
rect 50956 29384 50975 29418
rect 50903 29328 50975 29384
rect 50903 29294 50922 29328
rect 50956 29294 50975 29328
rect 50903 29238 50975 29294
rect 50903 29204 50922 29238
rect 50956 29204 50975 29238
rect 50903 29148 50975 29204
rect 50903 29114 50922 29148
rect 50956 29114 50975 29148
rect 50903 29058 50975 29114
rect 50903 29024 50922 29058
rect 50956 29024 50975 29058
rect 50903 28968 50975 29024
rect 50903 28934 50922 28968
rect 50956 28934 50975 28968
rect 50903 28878 50975 28934
rect 50013 28803 50085 28863
rect 50903 28844 50922 28878
rect 50956 28844 50975 28878
rect 50903 28803 50975 28844
rect 50013 28784 50975 28803
rect 50013 28750 50110 28784
rect 50144 28750 50200 28784
rect 50234 28750 50290 28784
rect 50324 28750 50380 28784
rect 50414 28750 50470 28784
rect 50504 28750 50560 28784
rect 50594 28750 50650 28784
rect 50684 28750 50740 28784
rect 50774 28750 50830 28784
rect 50864 28750 50975 28784
rect 50013 28731 50975 28750
rect 51039 29674 51071 29708
rect 51105 29674 51224 29708
rect 51258 29674 51289 29708
rect 52379 29708 52478 29757
rect 51039 29618 51289 29674
rect 51039 29584 51071 29618
rect 51105 29584 51224 29618
rect 51258 29584 51289 29618
rect 51039 29528 51289 29584
rect 51039 29494 51071 29528
rect 51105 29494 51224 29528
rect 51258 29494 51289 29528
rect 51039 29438 51289 29494
rect 51039 29404 51071 29438
rect 51105 29404 51224 29438
rect 51258 29404 51289 29438
rect 51039 29348 51289 29404
rect 51039 29314 51071 29348
rect 51105 29314 51224 29348
rect 51258 29314 51289 29348
rect 51039 29258 51289 29314
rect 51039 29224 51071 29258
rect 51105 29224 51224 29258
rect 51258 29224 51289 29258
rect 51039 29168 51289 29224
rect 51039 29134 51071 29168
rect 51105 29134 51224 29168
rect 51258 29134 51289 29168
rect 51039 29078 51289 29134
rect 51039 29044 51071 29078
rect 51105 29044 51224 29078
rect 51258 29044 51289 29078
rect 51039 28988 51289 29044
rect 51039 28954 51071 28988
rect 51105 28954 51224 28988
rect 51258 28954 51289 28988
rect 51039 28898 51289 28954
rect 51039 28864 51071 28898
rect 51105 28864 51224 28898
rect 51258 28864 51289 28898
rect 51039 28808 51289 28864
rect 51039 28774 51071 28808
rect 51105 28774 51224 28808
rect 51258 28774 51289 28808
rect 49699 28684 49731 28718
rect 49765 28684 49884 28718
rect 49918 28684 49949 28718
rect 49699 28667 49949 28684
rect 51039 28718 51289 28774
rect 51353 29676 52315 29693
rect 51353 29642 51374 29676
rect 51408 29642 51464 29676
rect 51498 29674 51554 29676
rect 51588 29674 51644 29676
rect 51678 29674 51734 29676
rect 51768 29674 51824 29676
rect 51858 29674 51914 29676
rect 51948 29674 52004 29676
rect 52038 29674 52094 29676
rect 52128 29674 52184 29676
rect 52218 29674 52274 29676
rect 51518 29642 51554 29674
rect 51608 29642 51644 29674
rect 51698 29642 51734 29674
rect 51788 29642 51824 29674
rect 51878 29642 51914 29674
rect 51968 29642 52004 29674
rect 52058 29642 52094 29674
rect 52148 29642 52184 29674
rect 52238 29642 52274 29674
rect 52308 29642 52315 29676
rect 51353 29640 51484 29642
rect 51518 29640 51574 29642
rect 51608 29640 51664 29642
rect 51698 29640 51754 29642
rect 51788 29640 51844 29642
rect 51878 29640 51934 29642
rect 51968 29640 52024 29642
rect 52058 29640 52114 29642
rect 52148 29640 52204 29642
rect 52238 29640 52315 29642
rect 51353 29621 52315 29640
rect 51353 29617 51425 29621
rect 51353 29583 51372 29617
rect 51406 29583 51425 29617
rect 51353 29527 51425 29583
rect 52243 29598 52315 29621
rect 52243 29564 52262 29598
rect 52296 29564 52315 29598
rect 51353 29493 51372 29527
rect 51406 29493 51425 29527
rect 51353 29437 51425 29493
rect 51353 29403 51372 29437
rect 51406 29403 51425 29437
rect 51353 29347 51425 29403
rect 51353 29313 51372 29347
rect 51406 29313 51425 29347
rect 51353 29257 51425 29313
rect 51353 29223 51372 29257
rect 51406 29223 51425 29257
rect 51353 29167 51425 29223
rect 51353 29133 51372 29167
rect 51406 29133 51425 29167
rect 51353 29077 51425 29133
rect 51353 29043 51372 29077
rect 51406 29043 51425 29077
rect 51353 28987 51425 29043
rect 51353 28953 51372 28987
rect 51406 28953 51425 28987
rect 51353 28897 51425 28953
rect 51353 28863 51372 28897
rect 51406 28863 51425 28897
rect 51487 29500 52181 29559
rect 51487 29466 51548 29500
rect 51582 29472 51638 29500
rect 51672 29472 51728 29500
rect 51762 29472 51818 29500
rect 51594 29466 51638 29472
rect 51694 29466 51728 29472
rect 51794 29466 51818 29472
rect 51852 29472 51908 29500
rect 51852 29466 51860 29472
rect 51487 29438 51560 29466
rect 51594 29438 51660 29466
rect 51694 29438 51760 29466
rect 51794 29438 51860 29466
rect 51894 29466 51908 29472
rect 51942 29472 51998 29500
rect 51942 29466 51960 29472
rect 51894 29438 51960 29466
rect 51994 29466 51998 29472
rect 52032 29472 52088 29500
rect 52032 29466 52060 29472
rect 52122 29466 52181 29500
rect 51994 29438 52060 29466
rect 52094 29438 52181 29466
rect 51487 29410 52181 29438
rect 51487 29376 51548 29410
rect 51582 29376 51638 29410
rect 51672 29376 51728 29410
rect 51762 29376 51818 29410
rect 51852 29376 51908 29410
rect 51942 29376 51998 29410
rect 52032 29376 52088 29410
rect 52122 29376 52181 29410
rect 51487 29372 52181 29376
rect 51487 29338 51560 29372
rect 51594 29338 51660 29372
rect 51694 29338 51760 29372
rect 51794 29338 51860 29372
rect 51894 29338 51960 29372
rect 51994 29338 52060 29372
rect 52094 29338 52181 29372
rect 51487 29320 52181 29338
rect 51487 29286 51548 29320
rect 51582 29286 51638 29320
rect 51672 29286 51728 29320
rect 51762 29286 51818 29320
rect 51852 29286 51908 29320
rect 51942 29286 51998 29320
rect 52032 29286 52088 29320
rect 52122 29286 52181 29320
rect 51487 29272 52181 29286
rect 51487 29238 51560 29272
rect 51594 29238 51660 29272
rect 51694 29238 51760 29272
rect 51794 29238 51860 29272
rect 51894 29238 51960 29272
rect 51994 29238 52060 29272
rect 52094 29238 52181 29272
rect 51487 29230 52181 29238
rect 51487 29196 51548 29230
rect 51582 29196 51638 29230
rect 51672 29196 51728 29230
rect 51762 29196 51818 29230
rect 51852 29196 51908 29230
rect 51942 29196 51998 29230
rect 52032 29196 52088 29230
rect 52122 29196 52181 29230
rect 51487 29172 52181 29196
rect 51487 29140 51560 29172
rect 51594 29140 51660 29172
rect 51694 29140 51760 29172
rect 51794 29140 51860 29172
rect 51487 29106 51548 29140
rect 51594 29138 51638 29140
rect 51694 29138 51728 29140
rect 51794 29138 51818 29140
rect 51582 29106 51638 29138
rect 51672 29106 51728 29138
rect 51762 29106 51818 29138
rect 51852 29138 51860 29140
rect 51894 29140 51960 29172
rect 51894 29138 51908 29140
rect 51852 29106 51908 29138
rect 51942 29138 51960 29140
rect 51994 29140 52060 29172
rect 52094 29140 52181 29172
rect 51994 29138 51998 29140
rect 51942 29106 51998 29138
rect 52032 29138 52060 29140
rect 52032 29106 52088 29138
rect 52122 29106 52181 29140
rect 51487 29072 52181 29106
rect 51487 29050 51560 29072
rect 51594 29050 51660 29072
rect 51694 29050 51760 29072
rect 51794 29050 51860 29072
rect 51487 29016 51548 29050
rect 51594 29038 51638 29050
rect 51694 29038 51728 29050
rect 51794 29038 51818 29050
rect 51582 29016 51638 29038
rect 51672 29016 51728 29038
rect 51762 29016 51818 29038
rect 51852 29038 51860 29050
rect 51894 29050 51960 29072
rect 51894 29038 51908 29050
rect 51852 29016 51908 29038
rect 51942 29038 51960 29050
rect 51994 29050 52060 29072
rect 52094 29050 52181 29072
rect 51994 29038 51998 29050
rect 51942 29016 51998 29038
rect 52032 29038 52060 29050
rect 52032 29016 52088 29038
rect 52122 29016 52181 29050
rect 51487 28972 52181 29016
rect 51487 28960 51560 28972
rect 51594 28960 51660 28972
rect 51694 28960 51760 28972
rect 51794 28960 51860 28972
rect 51487 28926 51548 28960
rect 51594 28938 51638 28960
rect 51694 28938 51728 28960
rect 51794 28938 51818 28960
rect 51582 28926 51638 28938
rect 51672 28926 51728 28938
rect 51762 28926 51818 28938
rect 51852 28938 51860 28960
rect 51894 28960 51960 28972
rect 51894 28938 51908 28960
rect 51852 28926 51908 28938
rect 51942 28938 51960 28960
rect 51994 28960 52060 28972
rect 52094 28960 52181 28972
rect 51994 28938 51998 28960
rect 51942 28926 51998 28938
rect 52032 28938 52060 28960
rect 52032 28926 52088 28938
rect 52122 28926 52181 28960
rect 51487 28865 52181 28926
rect 52243 29508 52315 29564
rect 52243 29474 52262 29508
rect 52296 29474 52315 29508
rect 52243 29418 52315 29474
rect 52243 29384 52262 29418
rect 52296 29384 52315 29418
rect 52243 29328 52315 29384
rect 52243 29294 52262 29328
rect 52296 29294 52315 29328
rect 52243 29238 52315 29294
rect 52243 29204 52262 29238
rect 52296 29204 52315 29238
rect 52243 29148 52315 29204
rect 52243 29114 52262 29148
rect 52296 29114 52315 29148
rect 52243 29058 52315 29114
rect 52243 29024 52262 29058
rect 52296 29024 52315 29058
rect 52243 28968 52315 29024
rect 52243 28934 52262 28968
rect 52296 28934 52315 28968
rect 52243 28878 52315 28934
rect 51353 28803 51425 28863
rect 52243 28844 52262 28878
rect 52296 28844 52315 28878
rect 52243 28803 52315 28844
rect 51353 28784 52315 28803
rect 51353 28750 51450 28784
rect 51484 28750 51540 28784
rect 51574 28750 51630 28784
rect 51664 28750 51720 28784
rect 51754 28750 51810 28784
rect 51844 28750 51900 28784
rect 51934 28750 51990 28784
rect 52024 28750 52080 28784
rect 52114 28750 52170 28784
rect 52204 28750 52315 28784
rect 51353 28731 52315 28750
rect 52379 29674 52411 29708
rect 52445 29674 52478 29708
rect 52379 29618 52478 29674
rect 52379 29584 52411 29618
rect 52445 29584 52478 29618
rect 52379 29528 52478 29584
rect 52379 29494 52411 29528
rect 52445 29494 52478 29528
rect 52379 29438 52478 29494
rect 52379 29404 52411 29438
rect 52445 29404 52478 29438
rect 52379 29348 52478 29404
rect 52379 29314 52411 29348
rect 52445 29314 52478 29348
rect 52379 29258 52478 29314
rect 52379 29224 52411 29258
rect 52445 29224 52478 29258
rect 52379 29168 52478 29224
rect 52379 29134 52411 29168
rect 52445 29134 52478 29168
rect 52379 29078 52478 29134
rect 52379 29044 52411 29078
rect 52445 29044 52478 29078
rect 52379 28988 52478 29044
rect 52379 28954 52411 28988
rect 52445 28954 52478 28988
rect 52379 28898 52478 28954
rect 52379 28864 52411 28898
rect 52445 28864 52478 28898
rect 52379 28808 52478 28864
rect 52379 28774 52411 28808
rect 52445 28774 52478 28808
rect 51039 28684 51071 28718
rect 51105 28684 51224 28718
rect 51258 28684 51289 28718
rect 51039 28667 51289 28684
rect 52379 28718 52478 28774
rect 52379 28684 52411 28718
rect 52445 28684 52478 28718
rect 52379 28667 52478 28684
rect 41810 28634 52478 28667
rect 41810 28600 41940 28634
rect 41974 28600 42030 28634
rect 42064 28600 42120 28634
rect 42154 28600 42210 28634
rect 42244 28600 42300 28634
rect 42334 28600 42390 28634
rect 42424 28600 42480 28634
rect 42514 28600 42570 28634
rect 42604 28600 42660 28634
rect 42694 28600 42750 28634
rect 42784 28600 42840 28634
rect 42874 28600 42930 28634
rect 42964 28600 43280 28634
rect 43314 28600 43370 28634
rect 43404 28600 43460 28634
rect 43494 28600 43550 28634
rect 43584 28600 43640 28634
rect 43674 28600 43730 28634
rect 43764 28600 43820 28634
rect 43854 28600 43910 28634
rect 43944 28600 44000 28634
rect 44034 28600 44090 28634
rect 44124 28600 44180 28634
rect 44214 28600 44270 28634
rect 44304 28600 44620 28634
rect 44654 28600 44710 28634
rect 44744 28600 44800 28634
rect 44834 28600 44890 28634
rect 44924 28600 44980 28634
rect 45014 28600 45070 28634
rect 45104 28600 45160 28634
rect 45194 28600 45250 28634
rect 45284 28600 45340 28634
rect 45374 28600 45430 28634
rect 45464 28600 45520 28634
rect 45554 28600 45610 28634
rect 45644 28600 45960 28634
rect 45994 28600 46050 28634
rect 46084 28600 46140 28634
rect 46174 28600 46230 28634
rect 46264 28600 46320 28634
rect 46354 28600 46410 28634
rect 46444 28600 46500 28634
rect 46534 28600 46590 28634
rect 46624 28600 46680 28634
rect 46714 28600 46770 28634
rect 46804 28600 46860 28634
rect 46894 28600 46950 28634
rect 46984 28600 47300 28634
rect 47334 28600 47390 28634
rect 47424 28600 47480 28634
rect 47514 28600 47570 28634
rect 47604 28600 47660 28634
rect 47694 28600 47750 28634
rect 47784 28600 47840 28634
rect 47874 28600 47930 28634
rect 47964 28600 48020 28634
rect 48054 28600 48110 28634
rect 48144 28600 48200 28634
rect 48234 28600 48290 28634
rect 48324 28600 48640 28634
rect 48674 28600 48730 28634
rect 48764 28600 48820 28634
rect 48854 28600 48910 28634
rect 48944 28600 49000 28634
rect 49034 28600 49090 28634
rect 49124 28600 49180 28634
rect 49214 28600 49270 28634
rect 49304 28600 49360 28634
rect 49394 28600 49450 28634
rect 49484 28600 49540 28634
rect 49574 28600 49630 28634
rect 49664 28600 49980 28634
rect 50014 28600 50070 28634
rect 50104 28600 50160 28634
rect 50194 28600 50250 28634
rect 50284 28600 50340 28634
rect 50374 28600 50430 28634
rect 50464 28600 50520 28634
rect 50554 28600 50610 28634
rect 50644 28600 50700 28634
rect 50734 28600 50790 28634
rect 50824 28600 50880 28634
rect 50914 28600 50970 28634
rect 51004 28600 51320 28634
rect 51354 28600 51410 28634
rect 51444 28600 51500 28634
rect 51534 28600 51590 28634
rect 51624 28600 51680 28634
rect 51714 28600 51770 28634
rect 51804 28600 51860 28634
rect 51894 28600 51950 28634
rect 51984 28600 52040 28634
rect 52074 28600 52130 28634
rect 52164 28600 52220 28634
rect 52254 28600 52310 28634
rect 52344 28600 52478 28634
rect 41810 28568 52478 28600
rect 38611 28509 40348 28542
rect 37472 28482 40348 28509
rect 37472 28423 40348 28436
rect 37472 28389 37655 28423
rect 37689 28389 38055 28423
rect 38089 28389 38455 28423
rect 38489 28407 38855 28423
rect 38489 28389 38577 28407
rect 37472 28376 38577 28389
rect 38611 28389 38855 28407
rect 38889 28389 39255 28423
rect 39289 28389 39655 28423
rect 39689 28389 40055 28423
rect 40089 28389 40348 28423
rect 38611 28376 40348 28389
rect 16520 28289 18960 28302
rect 16520 28255 16703 28289
rect 16737 28255 16903 28289
rect 16937 28255 17103 28289
rect 17137 28255 17303 28289
rect 17337 28255 17503 28289
rect 17537 28255 17703 28289
rect 17737 28255 17903 28289
rect 17937 28255 18103 28289
rect 18137 28255 18303 28289
rect 18337 28255 18503 28289
rect 18537 28255 18703 28289
rect 18737 28255 18960 28289
rect 16520 28242 18960 28255
rect 19264 28289 21704 28302
rect 19264 28255 19447 28289
rect 19481 28255 19647 28289
rect 19681 28255 19847 28289
rect 19881 28255 20047 28289
rect 20081 28255 20247 28289
rect 20281 28255 20447 28289
rect 20481 28255 20647 28289
rect 20681 28255 20847 28289
rect 20881 28255 21047 28289
rect 21081 28255 21247 28289
rect 21281 28255 21447 28289
rect 21481 28255 21704 28289
rect 19264 28242 21704 28255
rect 22008 28289 24448 28302
rect 22008 28255 22191 28289
rect 22225 28255 22391 28289
rect 22425 28255 22591 28289
rect 22625 28255 22791 28289
rect 22825 28255 22991 28289
rect 23025 28255 23191 28289
rect 23225 28255 23391 28289
rect 23425 28255 23591 28289
rect 23625 28255 23791 28289
rect 23825 28255 23991 28289
rect 24025 28255 24191 28289
rect 24225 28255 24448 28289
rect 22008 28242 24448 28255
rect 27202 28289 29642 28302
rect 27202 28255 27385 28289
rect 27419 28255 27585 28289
rect 27619 28255 27785 28289
rect 27819 28255 27985 28289
rect 28019 28255 28185 28289
rect 28219 28255 28385 28289
rect 28419 28255 28585 28289
rect 28619 28255 28785 28289
rect 28819 28255 28985 28289
rect 29019 28255 29185 28289
rect 29219 28255 29385 28289
rect 29419 28255 29642 28289
rect 27202 28242 29642 28255
rect 29928 28289 37096 28302
rect 29928 28255 30111 28289
rect 30145 28255 30511 28289
rect 30545 28255 30911 28289
rect 30945 28255 31311 28289
rect 31345 28255 31711 28289
rect 31745 28255 32111 28289
rect 32145 28255 32511 28289
rect 32545 28255 32911 28289
rect 32945 28255 33311 28289
rect 33345 28255 33711 28289
rect 33745 28255 34111 28289
rect 34145 28255 34511 28289
rect 34545 28255 34911 28289
rect 34945 28255 35311 28289
rect 35345 28255 35711 28289
rect 35745 28255 36111 28289
rect 36145 28255 36511 28289
rect 36545 28255 36911 28289
rect 36945 28255 37096 28289
rect 29928 28242 37096 28255
rect 37374 28289 40348 28302
rect 37374 28255 37655 28289
rect 37689 28255 38055 28289
rect 38089 28255 38455 28289
rect 38489 28255 38855 28289
rect 38889 28255 39255 28289
rect 39289 28255 39655 28289
rect 39689 28255 40055 28289
rect 40089 28255 40348 28289
rect 37374 28242 40348 28255
rect 41784 28289 52504 28302
rect 41784 28255 41967 28289
rect 42001 28255 42167 28289
rect 42201 28255 42367 28289
rect 42401 28255 42567 28289
rect 42601 28255 42767 28289
rect 42801 28255 42967 28289
rect 43001 28255 43167 28289
rect 43201 28255 43367 28289
rect 43401 28255 43567 28289
rect 43601 28255 43767 28289
rect 43801 28255 43967 28289
rect 44001 28255 44167 28289
rect 44201 28255 44367 28289
rect 44401 28255 44567 28289
rect 44601 28255 44767 28289
rect 44801 28255 44967 28289
rect 45001 28255 45167 28289
rect 45201 28255 45367 28289
rect 45401 28255 45567 28289
rect 45601 28255 45767 28289
rect 45801 28255 45967 28289
rect 46001 28255 46167 28289
rect 46201 28255 46367 28289
rect 46401 28255 46567 28289
rect 46601 28255 46767 28289
rect 46801 28255 46967 28289
rect 47001 28255 47167 28289
rect 47201 28255 47367 28289
rect 47401 28255 47567 28289
rect 47601 28255 47767 28289
rect 47801 28255 47967 28289
rect 48001 28255 48167 28289
rect 48201 28255 48367 28289
rect 48401 28255 48567 28289
rect 48601 28255 48767 28289
rect 48801 28255 48967 28289
rect 49001 28255 49167 28289
rect 49201 28255 49367 28289
rect 49401 28255 49567 28289
rect 49601 28255 49767 28289
rect 49801 28255 49967 28289
rect 50001 28255 50167 28289
rect 50201 28255 50367 28289
rect 50401 28255 50567 28289
rect 50601 28255 50767 28289
rect 50801 28255 50967 28289
rect 51001 28255 51167 28289
rect 51201 28255 51367 28289
rect 51401 28255 51567 28289
rect 51601 28255 51767 28289
rect 51801 28255 51967 28289
rect 52001 28255 52167 28289
rect 52201 28255 52367 28289
rect 52401 28255 52504 28289
rect 41784 28242 52504 28255
rect 22400 26409 24840 26422
rect 22400 26375 22583 26409
rect 22617 26375 22783 26409
rect 22817 26375 22983 26409
rect 23017 26375 23183 26409
rect 23217 26375 23383 26409
rect 23417 26375 23583 26409
rect 23617 26375 23783 26409
rect 23817 26375 23983 26409
rect 24017 26375 24183 26409
rect 24217 26375 24383 26409
rect 24417 26375 24583 26409
rect 24617 26375 24840 26409
rect 22400 26362 24840 26375
rect 25320 26409 29598 26422
rect 25320 26375 25601 26409
rect 25635 26375 26001 26409
rect 26035 26375 26401 26409
rect 26435 26375 26801 26409
rect 26835 26375 27201 26409
rect 27235 26375 27601 26409
rect 27635 26375 28001 26409
rect 28035 26375 28401 26409
rect 28435 26375 28801 26409
rect 28835 26375 29201 26409
rect 29235 26375 29598 26409
rect 25320 26362 29598 26375
rect 29928 26409 37096 26422
rect 29928 26375 30111 26409
rect 30145 26375 30511 26409
rect 30545 26375 30911 26409
rect 30945 26375 31311 26409
rect 31345 26375 31711 26409
rect 31745 26375 32111 26409
rect 32145 26375 32511 26409
rect 32545 26375 32911 26409
rect 32945 26375 33311 26409
rect 33345 26375 33711 26409
rect 33745 26375 34111 26409
rect 34145 26375 34511 26409
rect 34545 26375 34911 26409
rect 34945 26375 35311 26409
rect 35345 26375 35711 26409
rect 35745 26375 36111 26409
rect 36145 26375 36511 26409
rect 36545 26375 36911 26409
rect 36945 26375 37096 26409
rect 29928 26362 37096 26375
rect 37394 26409 39834 26422
rect 37394 26375 37577 26409
rect 37611 26375 37777 26409
rect 37811 26375 37977 26409
rect 38011 26375 38177 26409
rect 38211 26375 38377 26409
rect 38411 26375 38577 26409
rect 38611 26375 38777 26409
rect 38811 26375 38977 26409
rect 39011 26375 39177 26409
rect 39211 26375 39377 26409
rect 39411 26375 39577 26409
rect 39611 26375 39834 26409
rect 37394 26362 39834 26375
rect 40138 26409 42578 26422
rect 40138 26375 40321 26409
rect 40355 26375 40521 26409
rect 40555 26375 40721 26409
rect 40755 26375 40921 26409
rect 40955 26375 41121 26409
rect 41155 26375 41321 26409
rect 41355 26375 41521 26409
rect 41555 26375 41721 26409
rect 41755 26375 41921 26409
rect 41955 26375 42121 26409
rect 42155 26375 42321 26409
rect 42355 26375 42578 26409
rect 40138 26362 42578 26375
rect 42882 26409 45322 26422
rect 42882 26375 43065 26409
rect 43099 26375 43265 26409
rect 43299 26375 43465 26409
rect 43499 26375 43665 26409
rect 43699 26375 43865 26409
rect 43899 26375 44065 26409
rect 44099 26375 44265 26409
rect 44299 26375 44465 26409
rect 44499 26375 44665 26409
rect 44699 26375 44865 26409
rect 44899 26375 45065 26409
rect 45099 26375 45322 26409
rect 42882 26362 45322 26375
rect 45626 26409 48066 26422
rect 45626 26375 45809 26409
rect 45843 26375 46009 26409
rect 46043 26375 46209 26409
rect 46243 26375 46409 26409
rect 46443 26375 46609 26409
rect 46643 26375 46809 26409
rect 46843 26375 47009 26409
rect 47043 26375 47209 26409
rect 47243 26375 47409 26409
rect 47443 26375 47609 26409
rect 47643 26375 47809 26409
rect 47843 26375 48066 26409
rect 45626 26362 48066 26375
rect 48370 26409 50810 26422
rect 48370 26375 48553 26409
rect 48587 26375 48753 26409
rect 48787 26375 48953 26409
rect 48987 26375 49153 26409
rect 49187 26375 49353 26409
rect 49387 26375 49553 26409
rect 49587 26375 49753 26409
rect 49787 26375 49953 26409
rect 49987 26375 50153 26409
rect 50187 26375 50353 26409
rect 50387 26375 50553 26409
rect 50587 26375 50810 26409
rect 48370 26362 50810 26375
rect 25418 26202 29598 26262
rect 25887 25916 25921 26202
rect 26803 25916 26837 26202
rect 27719 25916 27753 26202
rect 28635 25916 28669 26202
rect 29551 25916 29585 26202
rect 23312 25443 23928 25482
rect 23312 25341 23399 25443
rect 23841 25341 23928 25443
rect 23312 24542 23928 25341
rect 24408 25197 24840 25587
rect 25430 25889 25464 25916
rect 25887 25898 25922 25916
rect 25430 25817 25464 25835
rect 25430 25745 25464 25767
rect 25430 25673 25464 25699
rect 25430 25601 25464 25631
rect 25430 25529 25464 25563
rect 25430 25461 25464 25495
rect 25430 25393 25464 25423
rect 25430 25325 25464 25351
rect 25430 25257 25464 25279
rect 25430 25189 25464 25207
rect 25429 25135 25430 25166
rect 25429 25108 25464 25135
rect 25888 25889 25922 25898
rect 25888 25817 25922 25835
rect 25888 25745 25922 25767
rect 25888 25673 25922 25699
rect 25888 25601 25922 25631
rect 25888 25529 25922 25563
rect 25888 25461 25922 25495
rect 25888 25393 25922 25423
rect 25888 25325 25922 25351
rect 25888 25257 25922 25279
rect 25888 25189 25922 25207
rect 26346 25889 26380 25916
rect 26803 25898 26838 25916
rect 26346 25817 26380 25835
rect 26346 25745 26380 25767
rect 26346 25673 26380 25699
rect 26346 25601 26380 25631
rect 26346 25529 26380 25563
rect 26346 25461 26380 25495
rect 26346 25393 26380 25423
rect 26346 25325 26380 25351
rect 26346 25257 26380 25279
rect 26346 25189 26380 25207
rect 25888 25108 25922 25135
rect 26345 25135 26346 25166
rect 26345 25108 26380 25135
rect 26804 25889 26838 25898
rect 26804 25817 26838 25835
rect 26804 25745 26838 25767
rect 26804 25673 26838 25699
rect 26804 25601 26838 25631
rect 26804 25529 26838 25563
rect 26804 25461 26838 25495
rect 26804 25393 26838 25423
rect 26804 25325 26838 25351
rect 26804 25257 26838 25279
rect 26804 25189 26838 25207
rect 27262 25889 27296 25916
rect 27719 25898 27754 25916
rect 27262 25817 27296 25835
rect 27262 25745 27296 25767
rect 27262 25673 27296 25699
rect 27262 25601 27296 25631
rect 27262 25529 27296 25563
rect 27262 25461 27296 25495
rect 27262 25393 27296 25423
rect 27262 25325 27296 25351
rect 27262 25257 27296 25279
rect 27262 25189 27296 25207
rect 26804 25108 26838 25135
rect 27261 25135 27262 25166
rect 27261 25108 27296 25135
rect 27720 25889 27754 25898
rect 27720 25817 27754 25835
rect 27720 25745 27754 25767
rect 27720 25673 27754 25699
rect 27720 25601 27754 25631
rect 27720 25529 27754 25563
rect 27720 25461 27754 25495
rect 27720 25393 27754 25423
rect 27720 25325 27754 25351
rect 27720 25257 27754 25279
rect 27720 25189 27754 25207
rect 28178 25889 28212 25916
rect 28635 25898 28670 25916
rect 28178 25817 28212 25835
rect 28178 25745 28212 25767
rect 28178 25673 28212 25699
rect 28178 25601 28212 25631
rect 28178 25529 28212 25563
rect 28178 25461 28212 25495
rect 28178 25393 28212 25423
rect 28178 25325 28212 25351
rect 28178 25257 28212 25279
rect 28178 25189 28212 25207
rect 27720 25108 27754 25135
rect 28177 25135 28178 25166
rect 28177 25108 28212 25135
rect 28636 25889 28670 25898
rect 28636 25817 28670 25835
rect 28636 25745 28670 25767
rect 28636 25673 28670 25699
rect 28636 25601 28670 25631
rect 28636 25529 28670 25563
rect 28636 25461 28670 25495
rect 28636 25393 28670 25423
rect 28636 25325 28670 25351
rect 28636 25257 28670 25279
rect 28636 25189 28670 25207
rect 29094 25889 29128 25916
rect 29551 25898 29586 25916
rect 29094 25817 29128 25835
rect 29094 25745 29128 25767
rect 29094 25673 29128 25699
rect 29094 25601 29128 25631
rect 29094 25529 29128 25563
rect 29094 25461 29128 25495
rect 29094 25393 29128 25423
rect 29094 25325 29128 25351
rect 29094 25257 29128 25279
rect 29094 25189 29128 25207
rect 28636 25108 28670 25135
rect 29093 25135 29094 25166
rect 29093 25108 29128 25135
rect 29552 25889 29586 25898
rect 29552 25817 29586 25835
rect 29552 25745 29586 25767
rect 29552 25673 29586 25699
rect 29552 25601 29586 25631
rect 29552 25529 29586 25563
rect 29552 25461 29586 25495
rect 29552 25393 29586 25423
rect 29552 25325 29586 25351
rect 29552 25257 29586 25279
rect 29552 25189 29586 25207
rect 38306 25443 38922 25482
rect 38306 25341 38393 25443
rect 38835 25341 38922 25443
rect 29552 25108 29586 25135
rect 25429 25042 25463 25108
rect 26345 25042 26379 25108
rect 27261 25042 27295 25108
rect 28177 25042 28211 25108
rect 29093 25042 29127 25108
rect 25418 24982 29598 25042
rect 25498 24871 29598 24876
rect 25498 24863 27537 24871
rect 25498 24829 25601 24863
rect 25635 24829 26001 24863
rect 26035 24829 26401 24863
rect 26435 24829 26801 24863
rect 26835 24829 27201 24863
rect 27235 24837 27537 24863
rect 27571 24863 29598 24871
rect 27571 24837 27601 24863
rect 27235 24829 27601 24837
rect 27635 24829 28001 24863
rect 28035 24829 28401 24863
rect 28435 24829 28801 24863
rect 28835 24829 29201 24863
rect 29235 24829 29598 24863
rect 25498 24816 29598 24829
rect 25348 24669 25408 24752
rect 25348 24635 25361 24669
rect 25395 24635 25408 24669
rect 25348 24542 25408 24635
rect 26398 24639 26558 24662
rect 26398 24605 26463 24639
rect 26497 24605 26558 24639
rect 26398 24542 26558 24605
rect 27698 24639 27858 24662
rect 27698 24605 27763 24639
rect 27797 24605 27858 24639
rect 27698 24542 27858 24605
rect 38306 24542 38922 25341
rect 39402 25197 39834 25587
rect 41050 25443 41666 25482
rect 41050 25341 41137 25443
rect 41579 25341 41666 25443
rect 41050 24542 41666 25341
rect 42146 25197 42578 25587
rect 43794 25443 44410 25482
rect 43794 25341 43881 25443
rect 44323 25341 44410 25443
rect 43794 24542 44410 25341
rect 44890 25197 45322 25587
rect 46538 25443 47154 25482
rect 46538 25341 46625 25443
rect 47067 25341 47154 25443
rect 46538 24542 47154 25341
rect 47634 25197 48066 25587
rect 49282 25443 49898 25482
rect 49282 25341 49369 25443
rect 49811 25341 49898 25443
rect 49282 24542 49898 25341
rect 50378 25197 50810 25587
rect 22400 24529 24840 24542
rect 22400 24495 22583 24529
rect 22617 24495 22783 24529
rect 22817 24495 22983 24529
rect 23017 24495 23183 24529
rect 23217 24495 23383 24529
rect 23417 24495 23583 24529
rect 23617 24495 23783 24529
rect 23817 24495 23983 24529
rect 24017 24495 24183 24529
rect 24217 24495 24383 24529
rect 24417 24495 24583 24529
rect 24617 24495 24840 24529
rect 22400 24482 24840 24495
rect 25320 24529 29598 24542
rect 25320 24495 25601 24529
rect 25635 24495 26001 24529
rect 26035 24495 26401 24529
rect 26435 24495 26801 24529
rect 26835 24495 27201 24529
rect 27235 24495 27601 24529
rect 27635 24495 28001 24529
rect 28035 24495 28401 24529
rect 28435 24495 28801 24529
rect 28835 24495 29201 24529
rect 29235 24495 29598 24529
rect 25320 24482 29598 24495
rect 29928 24529 37096 24542
rect 29928 24495 30111 24529
rect 30145 24495 30511 24529
rect 30545 24495 30911 24529
rect 30945 24495 31311 24529
rect 31345 24495 31711 24529
rect 31745 24495 32111 24529
rect 32145 24495 32511 24529
rect 32545 24495 32911 24529
rect 32945 24495 33311 24529
rect 33345 24495 33711 24529
rect 33745 24495 34111 24529
rect 34145 24495 34511 24529
rect 34545 24495 34911 24529
rect 34945 24495 35311 24529
rect 35345 24495 35711 24529
rect 35745 24495 36111 24529
rect 36145 24495 36511 24529
rect 36545 24495 36911 24529
rect 36945 24495 37096 24529
rect 29928 24482 37096 24495
rect 37394 24529 39834 24542
rect 37394 24495 37577 24529
rect 37611 24495 37777 24529
rect 37811 24495 37977 24529
rect 38011 24495 38177 24529
rect 38211 24495 38377 24529
rect 38411 24495 38577 24529
rect 38611 24495 38777 24529
rect 38811 24495 38977 24529
rect 39011 24495 39177 24529
rect 39211 24495 39377 24529
rect 39411 24495 39577 24529
rect 39611 24495 39834 24529
rect 37394 24482 39834 24495
rect 40138 24529 42578 24542
rect 40138 24495 40321 24529
rect 40355 24495 40521 24529
rect 40555 24495 40721 24529
rect 40755 24495 40921 24529
rect 40955 24495 41121 24529
rect 41155 24495 41321 24529
rect 41355 24495 41521 24529
rect 41555 24495 41721 24529
rect 41755 24495 41921 24529
rect 41955 24495 42121 24529
rect 42155 24495 42321 24529
rect 42355 24495 42578 24529
rect 40138 24482 42578 24495
rect 42882 24529 45322 24542
rect 42882 24495 43065 24529
rect 43099 24495 43265 24529
rect 43299 24495 43465 24529
rect 43499 24495 43665 24529
rect 43699 24495 43865 24529
rect 43899 24495 44065 24529
rect 44099 24495 44265 24529
rect 44299 24495 44465 24529
rect 44499 24495 44665 24529
rect 44699 24495 44865 24529
rect 44899 24495 45065 24529
rect 45099 24495 45322 24529
rect 42882 24482 45322 24495
rect 45626 24529 48066 24542
rect 45626 24495 45809 24529
rect 45843 24495 46009 24529
rect 46043 24495 46209 24529
rect 46243 24495 46409 24529
rect 46443 24495 46609 24529
rect 46643 24495 46809 24529
rect 46843 24495 47009 24529
rect 47043 24495 47209 24529
rect 47243 24495 47409 24529
rect 47443 24495 47609 24529
rect 47643 24495 47809 24529
rect 47843 24495 48066 24529
rect 45626 24482 48066 24495
rect 48370 24529 50810 24542
rect 48370 24495 48553 24529
rect 48587 24495 48753 24529
rect 48787 24495 48953 24529
rect 48987 24495 49153 24529
rect 49187 24495 49353 24529
rect 49387 24495 49553 24529
rect 49587 24495 49753 24529
rect 49787 24495 49953 24529
rect 49987 24495 50153 24529
rect 50187 24495 50353 24529
rect 50387 24495 50553 24529
rect 50587 24495 50810 24529
rect 48370 24482 50810 24495
rect 23870 22649 26310 22662
rect 23870 22615 24053 22649
rect 24087 22615 24253 22649
rect 24287 22615 24453 22649
rect 24487 22615 24653 22649
rect 24687 22615 24853 22649
rect 24887 22615 25053 22649
rect 25087 22615 25253 22649
rect 25287 22615 25453 22649
rect 25487 22615 25653 22649
rect 25687 22615 25853 22649
rect 25887 22615 26053 22649
rect 26087 22615 26310 22649
rect 23870 22602 26310 22615
rect 27202 22649 29642 22662
rect 27202 22615 27385 22649
rect 27419 22615 27585 22649
rect 27619 22615 27785 22649
rect 27819 22615 27985 22649
rect 28019 22615 28185 22649
rect 28219 22615 28385 22649
rect 28419 22615 28585 22649
rect 28619 22615 28785 22649
rect 28819 22615 28985 22649
rect 29019 22615 29185 22649
rect 29219 22615 29385 22649
rect 29419 22615 29642 22649
rect 27202 22602 29642 22615
rect 29946 22649 32386 22662
rect 29946 22615 30129 22649
rect 30163 22615 30329 22649
rect 30363 22615 30529 22649
rect 30563 22615 30729 22649
rect 30763 22615 30929 22649
rect 30963 22615 31129 22649
rect 31163 22615 31329 22649
rect 31363 22615 31529 22649
rect 31563 22615 31729 22649
rect 31763 22615 31929 22649
rect 31963 22615 32129 22649
rect 32163 22615 32386 22649
rect 29946 22602 32386 22615
rect 33180 22649 35620 22662
rect 33180 22615 33363 22649
rect 33397 22615 33563 22649
rect 33597 22615 33763 22649
rect 33797 22615 33963 22649
rect 33997 22615 34163 22649
rect 34197 22615 34363 22649
rect 34397 22615 34563 22649
rect 34597 22615 34763 22649
rect 34797 22615 34963 22649
rect 34997 22615 35163 22649
rect 35197 22615 35363 22649
rect 35397 22615 35620 22649
rect 33180 22602 35620 22615
rect 37394 22649 39834 22662
rect 37394 22615 37577 22649
rect 37611 22615 37777 22649
rect 37811 22615 37977 22649
rect 38011 22615 38177 22649
rect 38211 22615 38377 22649
rect 38411 22615 38577 22649
rect 38611 22615 38777 22649
rect 38811 22615 38977 22649
rect 39011 22615 39177 22649
rect 39211 22615 39377 22649
rect 39411 22615 39577 22649
rect 39611 22615 39834 22649
rect 37394 22602 39834 22615
rect 40138 22649 42578 22662
rect 40138 22615 40321 22649
rect 40355 22615 40521 22649
rect 40555 22615 40721 22649
rect 40755 22615 40921 22649
rect 40955 22615 41121 22649
rect 41155 22615 41321 22649
rect 41355 22615 41521 22649
rect 41555 22615 41721 22649
rect 41755 22615 41921 22649
rect 41955 22615 42121 22649
rect 42155 22615 42321 22649
rect 42355 22615 42578 22649
rect 40138 22602 42578 22615
rect 48370 22649 50810 22662
rect 48370 22615 48553 22649
rect 48587 22615 48753 22649
rect 48787 22615 48953 22649
rect 48987 22615 49153 22649
rect 49187 22615 49353 22649
rect 49387 22615 49553 22649
rect 49587 22615 49753 22649
rect 49787 22615 49953 22649
rect 49987 22615 50153 22649
rect 50187 22615 50353 22649
rect 50387 22615 50553 22649
rect 50587 22615 50810 22649
rect 48370 22602 50810 22615
rect 24782 21683 25398 21722
rect 24782 21581 24869 21683
rect 25311 21581 25398 21683
rect 24782 20782 25398 21581
rect 25878 21437 26310 21827
rect 28114 21683 28730 21722
rect 28114 21581 28201 21683
rect 28643 21581 28730 21683
rect 28114 20782 28730 21581
rect 29210 21437 29642 21827
rect 30858 21683 31474 21722
rect 30858 21581 30945 21683
rect 31387 21581 31474 21683
rect 30858 20782 31474 21581
rect 31954 21437 32386 21827
rect 34092 21683 34708 21722
rect 34092 21581 34179 21683
rect 34621 21581 34708 21683
rect 34092 20782 34708 21581
rect 35188 21437 35620 21827
rect 38306 21683 38922 21722
rect 38306 21581 38393 21683
rect 38835 21581 38922 21683
rect 38306 20782 38922 21581
rect 39402 21437 39834 21827
rect 41050 21683 41666 21722
rect 41050 21581 41137 21683
rect 41579 21581 41666 21683
rect 41050 20782 41666 21581
rect 42146 21437 42578 21827
rect 49282 21683 49898 21722
rect 49282 21581 49369 21683
rect 49811 21581 49898 21683
rect 49282 20782 49898 21581
rect 50378 21437 50810 21827
rect 23870 20769 26310 20782
rect 23870 20735 24053 20769
rect 24087 20735 24253 20769
rect 24287 20735 24453 20769
rect 24487 20735 24653 20769
rect 24687 20735 24853 20769
rect 24887 20735 25053 20769
rect 25087 20735 25253 20769
rect 25287 20735 25453 20769
rect 25487 20735 25653 20769
rect 25687 20735 25853 20769
rect 25887 20735 26053 20769
rect 26087 20735 26310 20769
rect 23870 20722 26310 20735
rect 27202 20769 29642 20782
rect 27202 20735 27385 20769
rect 27419 20735 27585 20769
rect 27619 20735 27785 20769
rect 27819 20735 27985 20769
rect 28019 20735 28185 20769
rect 28219 20735 28385 20769
rect 28419 20735 28585 20769
rect 28619 20735 28785 20769
rect 28819 20735 28985 20769
rect 29019 20735 29185 20769
rect 29219 20735 29385 20769
rect 29419 20735 29642 20769
rect 27202 20722 29642 20735
rect 29946 20769 32386 20782
rect 29946 20735 30129 20769
rect 30163 20735 30329 20769
rect 30363 20735 30529 20769
rect 30563 20735 30729 20769
rect 30763 20735 30929 20769
rect 30963 20735 31129 20769
rect 31163 20735 31329 20769
rect 31363 20735 31529 20769
rect 31563 20735 31729 20769
rect 31763 20735 31929 20769
rect 31963 20735 32129 20769
rect 32163 20735 32386 20769
rect 29946 20722 32386 20735
rect 33180 20769 35620 20782
rect 33180 20735 33363 20769
rect 33397 20735 33563 20769
rect 33597 20735 33763 20769
rect 33797 20735 33963 20769
rect 33997 20735 34163 20769
rect 34197 20735 34363 20769
rect 34397 20735 34563 20769
rect 34597 20735 34763 20769
rect 34797 20735 34963 20769
rect 34997 20735 35163 20769
rect 35197 20735 35363 20769
rect 35397 20735 35620 20769
rect 33180 20722 35620 20735
rect 37394 20769 39834 20782
rect 37394 20735 37577 20769
rect 37611 20735 37777 20769
rect 37811 20735 37977 20769
rect 38011 20735 38177 20769
rect 38211 20735 38377 20769
rect 38411 20735 38577 20769
rect 38611 20735 38777 20769
rect 38811 20735 38977 20769
rect 39011 20735 39177 20769
rect 39211 20735 39377 20769
rect 39411 20735 39577 20769
rect 39611 20735 39834 20769
rect 37394 20722 39834 20735
rect 40138 20769 42578 20782
rect 40138 20735 40321 20769
rect 40355 20735 40521 20769
rect 40555 20735 40721 20769
rect 40755 20735 40921 20769
rect 40955 20735 41121 20769
rect 41155 20735 41321 20769
rect 41355 20735 41521 20769
rect 41555 20735 41721 20769
rect 41755 20735 41921 20769
rect 41955 20735 42121 20769
rect 42155 20735 42321 20769
rect 42355 20735 42578 20769
rect 40138 20722 42578 20735
rect 48370 20769 50810 20782
rect 48370 20735 48553 20769
rect 48587 20735 48753 20769
rect 48787 20735 48953 20769
rect 48987 20735 49153 20769
rect 49187 20735 49353 20769
rect 49387 20735 49553 20769
rect 49587 20735 49753 20769
rect 49787 20735 49953 20769
rect 49987 20735 50153 20769
rect 50187 20735 50353 20769
rect 50387 20735 50553 20769
rect 50587 20735 50810 20769
rect 48370 20722 50810 20735
rect 24732 18889 52438 18902
rect 24732 18855 25013 18889
rect 25047 18855 25413 18889
rect 25447 18855 25813 18889
rect 25847 18855 26213 18889
rect 26247 18855 26613 18889
rect 26647 18855 27013 18889
rect 27047 18855 27413 18889
rect 27447 18855 27813 18889
rect 27847 18855 28213 18889
rect 28247 18855 28613 18889
rect 28647 18855 29013 18889
rect 29047 18855 29413 18889
rect 29447 18855 29813 18889
rect 29847 18855 30213 18889
rect 30247 18855 30613 18889
rect 30647 18855 31013 18889
rect 31047 18855 31413 18889
rect 31447 18855 31813 18889
rect 31847 18855 32213 18889
rect 32247 18855 32613 18889
rect 32647 18855 33013 18889
rect 33047 18855 33413 18889
rect 33447 18855 33813 18889
rect 33847 18855 34213 18889
rect 34247 18855 34613 18889
rect 34647 18855 35013 18889
rect 35047 18855 35413 18889
rect 35447 18855 35813 18889
rect 35847 18855 36213 18889
rect 36247 18855 36613 18889
rect 36647 18855 37013 18889
rect 37047 18855 37413 18889
rect 37447 18855 37813 18889
rect 37847 18855 38213 18889
rect 38247 18855 38613 18889
rect 38647 18855 39013 18889
rect 39047 18855 39413 18889
rect 39447 18855 39813 18889
rect 39847 18855 40213 18889
rect 40247 18855 40613 18889
rect 40647 18855 41013 18889
rect 41047 18855 41413 18889
rect 41447 18855 41813 18889
rect 41847 18855 42213 18889
rect 42247 18855 42613 18889
rect 42647 18855 43013 18889
rect 43047 18855 43413 18889
rect 43447 18855 43813 18889
rect 43847 18855 44213 18889
rect 44247 18855 44613 18889
rect 44647 18855 45013 18889
rect 45047 18855 45413 18889
rect 45447 18855 45813 18889
rect 45847 18855 46213 18889
rect 46247 18855 46613 18889
rect 46647 18855 47013 18889
rect 47047 18855 47413 18889
rect 47447 18855 47813 18889
rect 47847 18855 48213 18889
rect 48247 18855 48613 18889
rect 48647 18855 49013 18889
rect 49047 18855 49413 18889
rect 49447 18855 49813 18889
rect 49847 18855 50213 18889
rect 50247 18855 50613 18889
rect 50647 18855 51013 18889
rect 51047 18855 51413 18889
rect 51447 18855 51813 18889
rect 51847 18855 52213 18889
rect 52247 18855 52438 18889
rect 24732 18842 52438 18855
rect 24760 18749 24820 18842
rect 25808 18799 25968 18842
rect 25808 18765 25873 18799
rect 25907 18765 25968 18799
rect 25808 18762 25968 18765
rect 27108 18799 27268 18842
rect 27108 18765 27173 18799
rect 27207 18765 27268 18799
rect 27108 18762 27268 18765
rect 28408 18799 28568 18842
rect 28408 18765 28473 18799
rect 28507 18765 28568 18799
rect 28408 18762 28568 18765
rect 29708 18799 29868 18842
rect 29708 18765 29773 18799
rect 29807 18765 29868 18799
rect 29708 18762 29868 18765
rect 31008 18799 31168 18842
rect 31008 18765 31073 18799
rect 31107 18765 31168 18799
rect 31008 18762 31168 18765
rect 32308 18799 32468 18842
rect 32308 18765 32373 18799
rect 32407 18765 32468 18799
rect 32308 18762 32468 18765
rect 33608 18799 33768 18842
rect 33608 18765 33673 18799
rect 33707 18765 33768 18799
rect 33608 18762 33768 18765
rect 34908 18799 35068 18842
rect 34908 18765 34973 18799
rect 35007 18765 35068 18799
rect 34908 18762 35068 18765
rect 36208 18799 36368 18842
rect 36208 18765 36273 18799
rect 36307 18765 36368 18799
rect 36208 18762 36368 18765
rect 37508 18799 37668 18842
rect 37508 18765 37573 18799
rect 37607 18765 37668 18799
rect 37508 18762 37668 18765
rect 38808 18799 38968 18842
rect 38808 18765 38873 18799
rect 38907 18765 38968 18799
rect 38808 18762 38968 18765
rect 40108 18799 40268 18842
rect 40108 18765 40173 18799
rect 40207 18765 40268 18799
rect 40108 18762 40268 18765
rect 41408 18799 41568 18842
rect 41408 18765 41473 18799
rect 41507 18765 41568 18799
rect 41408 18762 41568 18765
rect 42708 18799 42868 18842
rect 42708 18765 42773 18799
rect 42807 18765 42868 18799
rect 42708 18762 42868 18765
rect 44008 18799 44168 18842
rect 44008 18765 44073 18799
rect 44107 18765 44168 18799
rect 44008 18762 44168 18765
rect 45308 18799 45468 18842
rect 45308 18765 45373 18799
rect 45407 18765 45468 18799
rect 45308 18762 45468 18765
rect 46608 18799 46768 18842
rect 46608 18765 46673 18799
rect 46707 18765 46768 18799
rect 46608 18762 46768 18765
rect 47908 18799 48068 18842
rect 47908 18765 47973 18799
rect 48007 18765 48068 18799
rect 47908 18762 48068 18765
rect 49208 18799 49368 18842
rect 49208 18765 49273 18799
rect 49307 18765 49368 18799
rect 49208 18762 49368 18765
rect 50508 18799 50668 18842
rect 50508 18765 50573 18799
rect 50607 18765 50668 18799
rect 50508 18762 50668 18765
rect 24760 18715 24773 18749
rect 24807 18715 24820 18749
rect 24760 18632 24820 18715
rect 24890 18682 52438 18722
rect 24877 18621 24911 18641
rect 24877 18553 24911 18587
rect 24877 18485 24911 18515
rect 24877 18417 24911 18443
rect 24877 18349 24911 18371
rect 24877 18281 24911 18299
rect 24877 18213 24911 18227
rect 24877 18145 24911 18155
rect 24877 18077 24911 18083
rect 24877 18009 24911 18011
rect 24877 17973 24911 17975
rect 24877 17901 24911 17907
rect 24877 17829 24911 17839
rect 24877 17757 24911 17771
rect 24877 17685 24911 17703
rect 24877 17613 24911 17635
rect 24877 17541 24911 17567
rect 24877 17469 24911 17499
rect 24877 17397 24911 17431
rect 24877 17262 24911 17363
rect 25335 18621 25369 18682
rect 25335 18553 25369 18587
rect 25335 18485 25369 18515
rect 25335 18417 25369 18443
rect 25335 18349 25369 18371
rect 25335 18281 25369 18299
rect 25335 18213 25369 18227
rect 25335 18145 25369 18155
rect 25335 18077 25369 18083
rect 25335 18009 25369 18011
rect 25335 17973 25369 17975
rect 25335 17901 25369 17907
rect 25335 17829 25369 17839
rect 25335 17757 25369 17771
rect 25335 17685 25369 17703
rect 25335 17613 25369 17635
rect 25335 17541 25369 17567
rect 25335 17469 25369 17499
rect 25335 17397 25369 17431
rect 25335 17343 25369 17363
rect 25793 18621 25827 18641
rect 25793 18553 25827 18587
rect 25793 18485 25827 18515
rect 25793 18417 25827 18443
rect 25793 18349 25827 18371
rect 25793 18281 25827 18299
rect 25793 18213 25827 18227
rect 25793 18145 25827 18155
rect 25793 18077 25827 18083
rect 25793 18009 25827 18011
rect 25793 17973 25827 17975
rect 25793 17901 25827 17907
rect 25793 17829 25827 17839
rect 25793 17757 25827 17771
rect 25793 17685 25827 17703
rect 25793 17613 25827 17635
rect 25793 17541 25827 17567
rect 25793 17469 25827 17499
rect 25793 17397 25827 17431
rect 25793 17262 25827 17363
rect 26251 18621 26285 18682
rect 26251 18553 26285 18587
rect 26251 18485 26285 18515
rect 26251 18417 26285 18443
rect 26251 18349 26285 18371
rect 26251 18281 26285 18299
rect 26251 18213 26285 18227
rect 26251 18145 26285 18155
rect 26251 18077 26285 18083
rect 26251 18009 26285 18011
rect 26251 17973 26285 17975
rect 26251 17901 26285 17907
rect 26251 17829 26285 17839
rect 26251 17757 26285 17771
rect 26251 17685 26285 17703
rect 26251 17613 26285 17635
rect 26251 17541 26285 17567
rect 26251 17469 26285 17499
rect 26251 17397 26285 17431
rect 26251 17343 26285 17363
rect 26709 18621 26743 18641
rect 26709 18553 26743 18587
rect 26709 18485 26743 18515
rect 26709 18417 26743 18443
rect 26709 18349 26743 18371
rect 26709 18281 26743 18299
rect 26709 18213 26743 18227
rect 26709 18145 26743 18155
rect 26709 18077 26743 18083
rect 26709 18009 26743 18011
rect 26709 17973 26743 17975
rect 26709 17901 26743 17907
rect 26709 17829 26743 17839
rect 26709 17757 26743 17771
rect 26709 17685 26743 17703
rect 26709 17613 26743 17635
rect 26709 17541 26743 17567
rect 26709 17469 26743 17499
rect 26709 17397 26743 17431
rect 26709 17262 26743 17363
rect 27167 18621 27201 18682
rect 27167 18553 27201 18587
rect 27167 18485 27201 18515
rect 27167 18417 27201 18443
rect 27167 18349 27201 18371
rect 27167 18281 27201 18299
rect 27167 18213 27201 18227
rect 27167 18145 27201 18155
rect 27167 18077 27201 18083
rect 27167 18009 27201 18011
rect 27167 17973 27201 17975
rect 27167 17901 27201 17907
rect 27167 17829 27201 17839
rect 27167 17757 27201 17771
rect 27167 17685 27201 17703
rect 27167 17613 27201 17635
rect 27167 17541 27201 17567
rect 27167 17469 27201 17499
rect 27167 17397 27201 17431
rect 27167 17343 27201 17363
rect 27625 18621 27659 18641
rect 27625 18553 27659 18587
rect 27625 18485 27659 18515
rect 27625 18417 27659 18443
rect 27625 18349 27659 18371
rect 27625 18281 27659 18299
rect 27625 18213 27659 18227
rect 27625 18145 27659 18155
rect 27625 18077 27659 18083
rect 27625 18009 27659 18011
rect 27625 17973 27659 17975
rect 27625 17901 27659 17907
rect 27625 17829 27659 17839
rect 27625 17757 27659 17771
rect 27625 17685 27659 17703
rect 27625 17613 27659 17635
rect 27625 17541 27659 17567
rect 27625 17469 27659 17499
rect 27625 17397 27659 17431
rect 27625 17262 27659 17363
rect 28083 18621 28117 18682
rect 28083 18553 28117 18587
rect 28083 18485 28117 18515
rect 28083 18417 28117 18443
rect 28083 18349 28117 18371
rect 28083 18281 28117 18299
rect 28083 18213 28117 18227
rect 28083 18145 28117 18155
rect 28083 18077 28117 18083
rect 28083 18009 28117 18011
rect 28083 17973 28117 17975
rect 28083 17901 28117 17907
rect 28083 17829 28117 17839
rect 28083 17757 28117 17771
rect 28083 17685 28117 17703
rect 28083 17613 28117 17635
rect 28083 17541 28117 17567
rect 28083 17469 28117 17499
rect 28083 17397 28117 17431
rect 28083 17343 28117 17363
rect 28541 18621 28575 18641
rect 28541 18553 28575 18587
rect 28541 18485 28575 18515
rect 28541 18417 28575 18443
rect 28541 18349 28575 18371
rect 28541 18281 28575 18299
rect 28541 18213 28575 18227
rect 28541 18145 28575 18155
rect 28541 18077 28575 18083
rect 28541 18009 28575 18011
rect 28541 17973 28575 17975
rect 28541 17901 28575 17907
rect 28541 17829 28575 17839
rect 28541 17757 28575 17771
rect 28541 17685 28575 17703
rect 28541 17613 28575 17635
rect 28541 17541 28575 17567
rect 28541 17469 28575 17499
rect 28541 17397 28575 17431
rect 28541 17262 28575 17363
rect 28999 18621 29033 18682
rect 28999 18553 29033 18587
rect 28999 18485 29033 18515
rect 28999 18417 29033 18443
rect 28999 18349 29033 18371
rect 28999 18281 29033 18299
rect 28999 18213 29033 18227
rect 28999 18145 29033 18155
rect 28999 18077 29033 18083
rect 28999 18009 29033 18011
rect 28999 17973 29033 17975
rect 28999 17901 29033 17907
rect 28999 17829 29033 17839
rect 28999 17757 29033 17771
rect 28999 17685 29033 17703
rect 28999 17613 29033 17635
rect 28999 17541 29033 17567
rect 28999 17469 29033 17499
rect 28999 17397 29033 17431
rect 28999 17343 29033 17363
rect 29457 18621 29491 18641
rect 29457 18553 29491 18587
rect 29457 18485 29491 18515
rect 29457 18417 29491 18443
rect 29457 18349 29491 18371
rect 29457 18281 29491 18299
rect 29457 18213 29491 18227
rect 29457 18145 29491 18155
rect 29457 18077 29491 18083
rect 29457 18009 29491 18011
rect 29457 17973 29491 17975
rect 29457 17901 29491 17907
rect 29457 17829 29491 17839
rect 29457 17757 29491 17771
rect 29457 17685 29491 17703
rect 29457 17613 29491 17635
rect 29457 17541 29491 17567
rect 29457 17469 29491 17499
rect 29457 17397 29491 17431
rect 29457 17262 29491 17363
rect 29915 18621 29949 18682
rect 29915 18553 29949 18587
rect 29915 18485 29949 18515
rect 29915 18417 29949 18443
rect 29915 18349 29949 18371
rect 29915 18281 29949 18299
rect 29915 18213 29949 18227
rect 29915 18145 29949 18155
rect 29915 18077 29949 18083
rect 29915 18009 29949 18011
rect 29915 17973 29949 17975
rect 29915 17901 29949 17907
rect 29915 17829 29949 17839
rect 29915 17757 29949 17771
rect 29915 17685 29949 17703
rect 29915 17613 29949 17635
rect 29915 17541 29949 17567
rect 29915 17469 29949 17499
rect 29915 17397 29949 17431
rect 29915 17343 29949 17363
rect 30373 18621 30407 18641
rect 30373 18553 30407 18587
rect 30373 18485 30407 18515
rect 30373 18417 30407 18443
rect 30373 18349 30407 18371
rect 30373 18281 30407 18299
rect 30373 18213 30407 18227
rect 30373 18145 30407 18155
rect 30373 18077 30407 18083
rect 30373 18009 30407 18011
rect 30373 17973 30407 17975
rect 30373 17901 30407 17907
rect 30373 17829 30407 17839
rect 30373 17757 30407 17771
rect 30373 17685 30407 17703
rect 30373 17613 30407 17635
rect 30373 17541 30407 17567
rect 30373 17469 30407 17499
rect 30373 17397 30407 17431
rect 30373 17262 30407 17363
rect 30831 18621 30865 18682
rect 30831 18553 30865 18587
rect 30831 18485 30865 18515
rect 30831 18417 30865 18443
rect 30831 18349 30865 18371
rect 30831 18281 30865 18299
rect 30831 18213 30865 18227
rect 30831 18145 30865 18155
rect 30831 18077 30865 18083
rect 30831 18009 30865 18011
rect 30831 17973 30865 17975
rect 30831 17901 30865 17907
rect 30831 17829 30865 17839
rect 30831 17757 30865 17771
rect 30831 17685 30865 17703
rect 30831 17613 30865 17635
rect 30831 17541 30865 17567
rect 30831 17469 30865 17499
rect 30831 17397 30865 17431
rect 30831 17343 30865 17363
rect 31289 18621 31323 18641
rect 31289 18553 31323 18587
rect 31289 18485 31323 18515
rect 31289 18417 31323 18443
rect 31289 18349 31323 18371
rect 31289 18281 31323 18299
rect 31289 18213 31323 18227
rect 31289 18145 31323 18155
rect 31289 18077 31323 18083
rect 31289 18009 31323 18011
rect 31289 17973 31323 17975
rect 31289 17901 31323 17907
rect 31289 17829 31323 17839
rect 31289 17757 31323 17771
rect 31289 17685 31323 17703
rect 31289 17613 31323 17635
rect 31289 17541 31323 17567
rect 31289 17469 31323 17499
rect 31289 17397 31323 17431
rect 31289 17262 31323 17363
rect 31747 18621 31781 18682
rect 31747 18553 31781 18587
rect 31747 18485 31781 18515
rect 31747 18417 31781 18443
rect 31747 18349 31781 18371
rect 31747 18281 31781 18299
rect 31747 18213 31781 18227
rect 31747 18145 31781 18155
rect 31747 18077 31781 18083
rect 31747 18009 31781 18011
rect 31747 17973 31781 17975
rect 31747 17901 31781 17907
rect 31747 17829 31781 17839
rect 31747 17757 31781 17771
rect 31747 17685 31781 17703
rect 31747 17613 31781 17635
rect 31747 17541 31781 17567
rect 31747 17469 31781 17499
rect 31747 17397 31781 17431
rect 31747 17343 31781 17363
rect 32205 18621 32239 18641
rect 32205 18553 32239 18587
rect 32205 18485 32239 18515
rect 32205 18417 32239 18443
rect 32205 18349 32239 18371
rect 32205 18281 32239 18299
rect 32205 18213 32239 18227
rect 32205 18145 32239 18155
rect 32205 18077 32239 18083
rect 32205 18009 32239 18011
rect 32205 17973 32239 17975
rect 32205 17901 32239 17907
rect 32205 17829 32239 17839
rect 32205 17757 32239 17771
rect 32205 17685 32239 17703
rect 32205 17613 32239 17635
rect 32205 17541 32239 17567
rect 32205 17469 32239 17499
rect 32205 17397 32239 17431
rect 32205 17262 32239 17363
rect 32663 18621 32697 18682
rect 32663 18553 32697 18587
rect 32663 18485 32697 18515
rect 32663 18417 32697 18443
rect 32663 18349 32697 18371
rect 32663 18281 32697 18299
rect 32663 18213 32697 18227
rect 32663 18145 32697 18155
rect 32663 18077 32697 18083
rect 32663 18009 32697 18011
rect 32663 17973 32697 17975
rect 32663 17901 32697 17907
rect 32663 17829 32697 17839
rect 32663 17757 32697 17771
rect 32663 17685 32697 17703
rect 32663 17613 32697 17635
rect 32663 17541 32697 17567
rect 32663 17469 32697 17499
rect 32663 17397 32697 17431
rect 32663 17343 32697 17363
rect 33121 18621 33155 18641
rect 33121 18553 33155 18587
rect 33121 18485 33155 18515
rect 33121 18417 33155 18443
rect 33121 18349 33155 18371
rect 33121 18281 33155 18299
rect 33121 18213 33155 18227
rect 33121 18145 33155 18155
rect 33121 18077 33155 18083
rect 33121 18009 33155 18011
rect 33121 17973 33155 17975
rect 33121 17901 33155 17907
rect 33121 17829 33155 17839
rect 33121 17757 33155 17771
rect 33121 17685 33155 17703
rect 33121 17613 33155 17635
rect 33121 17541 33155 17567
rect 33121 17469 33155 17499
rect 33121 17397 33155 17431
rect 33121 17262 33155 17363
rect 33579 18621 33613 18682
rect 33579 18553 33613 18587
rect 33579 18485 33613 18515
rect 33579 18417 33613 18443
rect 33579 18349 33613 18371
rect 33579 18281 33613 18299
rect 33579 18213 33613 18227
rect 33579 18145 33613 18155
rect 33579 18077 33613 18083
rect 33579 18009 33613 18011
rect 33579 17973 33613 17975
rect 33579 17901 33613 17907
rect 33579 17829 33613 17839
rect 33579 17757 33613 17771
rect 33579 17685 33613 17703
rect 33579 17613 33613 17635
rect 33579 17541 33613 17567
rect 33579 17469 33613 17499
rect 33579 17397 33613 17431
rect 33579 17343 33613 17363
rect 34037 18621 34071 18641
rect 34037 18553 34071 18587
rect 34037 18485 34071 18515
rect 34037 18417 34071 18443
rect 34037 18349 34071 18371
rect 34037 18281 34071 18299
rect 34037 18213 34071 18227
rect 34037 18145 34071 18155
rect 34037 18077 34071 18083
rect 34037 18009 34071 18011
rect 34037 17973 34071 17975
rect 34037 17901 34071 17907
rect 34037 17829 34071 17839
rect 34037 17757 34071 17771
rect 34037 17685 34071 17703
rect 34037 17613 34071 17635
rect 34037 17541 34071 17567
rect 34037 17469 34071 17499
rect 34037 17397 34071 17431
rect 34037 17262 34071 17363
rect 34495 18621 34529 18682
rect 34495 18553 34529 18587
rect 34495 18485 34529 18515
rect 34495 18417 34529 18443
rect 34495 18349 34529 18371
rect 34495 18281 34529 18299
rect 34495 18213 34529 18227
rect 34495 18145 34529 18155
rect 34495 18077 34529 18083
rect 34495 18009 34529 18011
rect 34495 17973 34529 17975
rect 34495 17901 34529 17907
rect 34495 17829 34529 17839
rect 34495 17757 34529 17771
rect 34495 17685 34529 17703
rect 34495 17613 34529 17635
rect 34495 17541 34529 17567
rect 34495 17469 34529 17499
rect 34495 17397 34529 17431
rect 34495 17343 34529 17363
rect 34953 18621 34987 18641
rect 34953 18553 34987 18587
rect 34953 18485 34987 18515
rect 34953 18417 34987 18443
rect 34953 18349 34987 18371
rect 34953 18281 34987 18299
rect 34953 18213 34987 18227
rect 34953 18145 34987 18155
rect 34953 18077 34987 18083
rect 34953 18009 34987 18011
rect 34953 17973 34987 17975
rect 34953 17901 34987 17907
rect 34953 17829 34987 17839
rect 34953 17757 34987 17771
rect 34953 17685 34987 17703
rect 34953 17613 34987 17635
rect 34953 17541 34987 17567
rect 34953 17469 34987 17499
rect 34953 17397 34987 17431
rect 34953 17262 34987 17363
rect 35411 18621 35445 18682
rect 35411 18553 35445 18587
rect 35411 18485 35445 18515
rect 35411 18417 35445 18443
rect 35411 18349 35445 18371
rect 35411 18281 35445 18299
rect 35411 18213 35445 18227
rect 35411 18145 35445 18155
rect 35411 18077 35445 18083
rect 35411 18009 35445 18011
rect 35411 17973 35445 17975
rect 35411 17901 35445 17907
rect 35411 17829 35445 17839
rect 35411 17757 35445 17771
rect 35411 17685 35445 17703
rect 35411 17613 35445 17635
rect 35411 17541 35445 17567
rect 35411 17469 35445 17499
rect 35411 17397 35445 17431
rect 35411 17343 35445 17363
rect 35869 18621 35903 18641
rect 35869 18553 35903 18587
rect 35869 18485 35903 18515
rect 35869 18417 35903 18443
rect 35869 18349 35903 18371
rect 35869 18281 35903 18299
rect 35869 18213 35903 18227
rect 35869 18145 35903 18155
rect 35869 18077 35903 18083
rect 35869 18009 35903 18011
rect 35869 17973 35903 17975
rect 35869 17901 35903 17907
rect 35869 17829 35903 17839
rect 35869 17757 35903 17771
rect 35869 17685 35903 17703
rect 35869 17613 35903 17635
rect 35869 17541 35903 17567
rect 35869 17469 35903 17499
rect 35869 17397 35903 17431
rect 35869 17262 35903 17363
rect 36327 18621 36361 18682
rect 36327 18553 36361 18587
rect 36327 18485 36361 18515
rect 36327 18417 36361 18443
rect 36327 18349 36361 18371
rect 36327 18281 36361 18299
rect 36327 18213 36361 18227
rect 36327 18145 36361 18155
rect 36327 18077 36361 18083
rect 36327 18009 36361 18011
rect 36327 17973 36361 17975
rect 36327 17901 36361 17907
rect 36327 17829 36361 17839
rect 36327 17757 36361 17771
rect 36327 17685 36361 17703
rect 36327 17613 36361 17635
rect 36327 17541 36361 17567
rect 36327 17469 36361 17499
rect 36327 17397 36361 17431
rect 36327 17343 36361 17363
rect 36785 18621 36819 18641
rect 36785 18553 36819 18587
rect 36785 18485 36819 18515
rect 36785 18417 36819 18443
rect 36785 18349 36819 18371
rect 36785 18281 36819 18299
rect 36785 18213 36819 18227
rect 36785 18145 36819 18155
rect 36785 18077 36819 18083
rect 36785 18009 36819 18011
rect 36785 17973 36819 17975
rect 36785 17901 36819 17907
rect 36785 17829 36819 17839
rect 36785 17757 36819 17771
rect 36785 17685 36819 17703
rect 36785 17613 36819 17635
rect 36785 17541 36819 17567
rect 36785 17469 36819 17499
rect 36785 17397 36819 17431
rect 36785 17262 36819 17363
rect 37243 18621 37277 18682
rect 37243 18553 37277 18587
rect 37243 18485 37277 18515
rect 37243 18417 37277 18443
rect 37243 18349 37277 18371
rect 37243 18281 37277 18299
rect 37243 18213 37277 18227
rect 37243 18145 37277 18155
rect 37243 18077 37277 18083
rect 37243 18009 37277 18011
rect 37243 17973 37277 17975
rect 37243 17901 37277 17907
rect 37243 17829 37277 17839
rect 37243 17757 37277 17771
rect 37243 17685 37277 17703
rect 37243 17613 37277 17635
rect 37243 17541 37277 17567
rect 37243 17469 37277 17499
rect 37243 17397 37277 17431
rect 37243 17343 37277 17363
rect 37701 18621 37735 18641
rect 37701 18553 37735 18587
rect 37701 18485 37735 18515
rect 37701 18417 37735 18443
rect 37701 18349 37735 18371
rect 37701 18281 37735 18299
rect 37701 18213 37735 18227
rect 37701 18145 37735 18155
rect 37701 18077 37735 18083
rect 37701 18009 37735 18011
rect 37701 17973 37735 17975
rect 37701 17901 37735 17907
rect 37701 17829 37735 17839
rect 37701 17757 37735 17771
rect 37701 17685 37735 17703
rect 37701 17613 37735 17635
rect 37701 17541 37735 17567
rect 37701 17469 37735 17499
rect 37701 17397 37735 17431
rect 37701 17262 37735 17363
rect 38159 18621 38193 18682
rect 38159 18553 38193 18587
rect 38159 18485 38193 18515
rect 38159 18417 38193 18443
rect 38159 18349 38193 18371
rect 38159 18281 38193 18299
rect 38159 18213 38193 18227
rect 38159 18145 38193 18155
rect 38159 18077 38193 18083
rect 38159 18009 38193 18011
rect 38159 17973 38193 17975
rect 38159 17901 38193 17907
rect 38159 17829 38193 17839
rect 38159 17757 38193 17771
rect 38159 17685 38193 17703
rect 38159 17613 38193 17635
rect 38159 17541 38193 17567
rect 38159 17469 38193 17499
rect 38159 17397 38193 17431
rect 38159 17343 38193 17363
rect 38617 18621 38651 18641
rect 38617 18553 38651 18587
rect 38617 18485 38651 18515
rect 38617 18417 38651 18443
rect 38617 18349 38651 18371
rect 38617 18281 38651 18299
rect 38617 18213 38651 18227
rect 38617 18145 38651 18155
rect 38617 18077 38651 18083
rect 38617 18009 38651 18011
rect 38617 17973 38651 17975
rect 38617 17901 38651 17907
rect 38617 17829 38651 17839
rect 38617 17757 38651 17771
rect 38617 17685 38651 17703
rect 38617 17613 38651 17635
rect 38617 17541 38651 17567
rect 38617 17469 38651 17499
rect 38617 17397 38651 17431
rect 38617 17262 38651 17363
rect 39075 18621 39109 18682
rect 39075 18553 39109 18587
rect 39075 18485 39109 18515
rect 39075 18417 39109 18443
rect 39075 18349 39109 18371
rect 39075 18281 39109 18299
rect 39075 18213 39109 18227
rect 39075 18145 39109 18155
rect 39075 18077 39109 18083
rect 39075 18009 39109 18011
rect 39075 17973 39109 17975
rect 39075 17901 39109 17907
rect 39075 17829 39109 17839
rect 39075 17757 39109 17771
rect 39075 17685 39109 17703
rect 39075 17613 39109 17635
rect 39075 17541 39109 17567
rect 39075 17469 39109 17499
rect 39075 17397 39109 17431
rect 39075 17343 39109 17363
rect 39533 18621 39567 18641
rect 39533 18553 39567 18587
rect 39533 18485 39567 18515
rect 39533 18417 39567 18443
rect 39533 18349 39567 18371
rect 39533 18281 39567 18299
rect 39533 18213 39567 18227
rect 39533 18145 39567 18155
rect 39533 18077 39567 18083
rect 39533 18009 39567 18011
rect 39533 17973 39567 17975
rect 39533 17901 39567 17907
rect 39533 17829 39567 17839
rect 39533 17757 39567 17771
rect 39533 17685 39567 17703
rect 39533 17613 39567 17635
rect 39533 17541 39567 17567
rect 39533 17469 39567 17499
rect 39533 17397 39567 17431
rect 39533 17262 39567 17363
rect 39991 18621 40025 18682
rect 39991 18553 40025 18587
rect 39991 18485 40025 18515
rect 39991 18417 40025 18443
rect 39991 18349 40025 18371
rect 39991 18281 40025 18299
rect 39991 18213 40025 18227
rect 39991 18145 40025 18155
rect 39991 18077 40025 18083
rect 39991 18009 40025 18011
rect 39991 17973 40025 17975
rect 39991 17901 40025 17907
rect 39991 17829 40025 17839
rect 39991 17757 40025 17771
rect 39991 17685 40025 17703
rect 39991 17613 40025 17635
rect 39991 17541 40025 17567
rect 39991 17469 40025 17499
rect 39991 17397 40025 17431
rect 39991 17343 40025 17363
rect 40449 18621 40483 18641
rect 40449 18553 40483 18587
rect 40449 18485 40483 18515
rect 40449 18417 40483 18443
rect 40449 18349 40483 18371
rect 40449 18281 40483 18299
rect 40449 18213 40483 18227
rect 40449 18145 40483 18155
rect 40449 18077 40483 18083
rect 40449 18009 40483 18011
rect 40449 17973 40483 17975
rect 40449 17901 40483 17907
rect 40449 17829 40483 17839
rect 40449 17757 40483 17771
rect 40449 17685 40483 17703
rect 40449 17613 40483 17635
rect 40449 17541 40483 17567
rect 40449 17469 40483 17499
rect 40449 17397 40483 17431
rect 40449 17262 40483 17363
rect 40907 18621 40941 18682
rect 40907 18553 40941 18587
rect 40907 18485 40941 18515
rect 40907 18417 40941 18443
rect 40907 18349 40941 18371
rect 40907 18281 40941 18299
rect 40907 18213 40941 18227
rect 40907 18145 40941 18155
rect 40907 18077 40941 18083
rect 40907 18009 40941 18011
rect 40907 17973 40941 17975
rect 40907 17901 40941 17907
rect 40907 17829 40941 17839
rect 40907 17757 40941 17771
rect 40907 17685 40941 17703
rect 40907 17613 40941 17635
rect 40907 17541 40941 17567
rect 40907 17469 40941 17499
rect 40907 17397 40941 17431
rect 40907 17343 40941 17363
rect 41365 18621 41399 18641
rect 41365 18553 41399 18587
rect 41365 18485 41399 18515
rect 41365 18417 41399 18443
rect 41365 18349 41399 18371
rect 41365 18281 41399 18299
rect 41365 18213 41399 18227
rect 41365 18145 41399 18155
rect 41365 18077 41399 18083
rect 41365 18009 41399 18011
rect 41365 17973 41399 17975
rect 41365 17901 41399 17907
rect 41365 17829 41399 17839
rect 41365 17757 41399 17771
rect 41365 17685 41399 17703
rect 41365 17613 41399 17635
rect 41365 17541 41399 17567
rect 41365 17469 41399 17499
rect 41365 17397 41399 17431
rect 41365 17262 41399 17363
rect 41823 18621 41857 18682
rect 41823 18553 41857 18587
rect 41823 18485 41857 18515
rect 41823 18417 41857 18443
rect 41823 18349 41857 18371
rect 41823 18281 41857 18299
rect 41823 18213 41857 18227
rect 41823 18145 41857 18155
rect 41823 18077 41857 18083
rect 41823 18009 41857 18011
rect 41823 17973 41857 17975
rect 41823 17901 41857 17907
rect 41823 17829 41857 17839
rect 41823 17757 41857 17771
rect 41823 17685 41857 17703
rect 41823 17613 41857 17635
rect 41823 17541 41857 17567
rect 41823 17469 41857 17499
rect 41823 17397 41857 17431
rect 41823 17343 41857 17363
rect 42281 18621 42315 18641
rect 42281 18553 42315 18587
rect 42281 18485 42315 18515
rect 42281 18417 42315 18443
rect 42281 18349 42315 18371
rect 42281 18281 42315 18299
rect 42281 18213 42315 18227
rect 42281 18145 42315 18155
rect 42281 18077 42315 18083
rect 42281 18009 42315 18011
rect 42281 17973 42315 17975
rect 42281 17901 42315 17907
rect 42281 17829 42315 17839
rect 42281 17757 42315 17771
rect 42281 17685 42315 17703
rect 42281 17613 42315 17635
rect 42281 17541 42315 17567
rect 42281 17469 42315 17499
rect 42281 17397 42315 17431
rect 42281 17262 42315 17363
rect 42739 18621 42773 18682
rect 42739 18553 42773 18587
rect 42739 18485 42773 18515
rect 42739 18417 42773 18443
rect 42739 18349 42773 18371
rect 42739 18281 42773 18299
rect 42739 18213 42773 18227
rect 42739 18145 42773 18155
rect 42739 18077 42773 18083
rect 42739 18009 42773 18011
rect 42739 17973 42773 17975
rect 42739 17901 42773 17907
rect 42739 17829 42773 17839
rect 42739 17757 42773 17771
rect 42739 17685 42773 17703
rect 42739 17613 42773 17635
rect 42739 17541 42773 17567
rect 42739 17469 42773 17499
rect 42739 17397 42773 17431
rect 42739 17343 42773 17363
rect 43197 18621 43231 18641
rect 43197 18553 43231 18587
rect 43197 18485 43231 18515
rect 43197 18417 43231 18443
rect 43197 18349 43231 18371
rect 43197 18281 43231 18299
rect 43197 18213 43231 18227
rect 43197 18145 43231 18155
rect 43197 18077 43231 18083
rect 43197 18009 43231 18011
rect 43197 17973 43231 17975
rect 43197 17901 43231 17907
rect 43197 17829 43231 17839
rect 43197 17757 43231 17771
rect 43197 17685 43231 17703
rect 43197 17613 43231 17635
rect 43197 17541 43231 17567
rect 43197 17469 43231 17499
rect 43197 17397 43231 17431
rect 43197 17262 43231 17363
rect 43655 18621 43689 18682
rect 43655 18553 43689 18587
rect 43655 18485 43689 18515
rect 43655 18417 43689 18443
rect 43655 18349 43689 18371
rect 43655 18281 43689 18299
rect 43655 18213 43689 18227
rect 43655 18145 43689 18155
rect 43655 18077 43689 18083
rect 43655 18009 43689 18011
rect 43655 17973 43689 17975
rect 43655 17901 43689 17907
rect 43655 17829 43689 17839
rect 43655 17757 43689 17771
rect 43655 17685 43689 17703
rect 43655 17613 43689 17635
rect 43655 17541 43689 17567
rect 43655 17469 43689 17499
rect 43655 17397 43689 17431
rect 43655 17343 43689 17363
rect 44113 18621 44147 18641
rect 44113 18553 44147 18587
rect 44113 18485 44147 18515
rect 44113 18417 44147 18443
rect 44113 18349 44147 18371
rect 44113 18281 44147 18299
rect 44113 18213 44147 18227
rect 44113 18145 44147 18155
rect 44113 18077 44147 18083
rect 44113 18009 44147 18011
rect 44113 17973 44147 17975
rect 44113 17901 44147 17907
rect 44113 17829 44147 17839
rect 44113 17757 44147 17771
rect 44113 17685 44147 17703
rect 44113 17613 44147 17635
rect 44113 17541 44147 17567
rect 44113 17469 44147 17499
rect 44113 17397 44147 17431
rect 44113 17262 44147 17363
rect 44571 18621 44605 18682
rect 44571 18553 44605 18587
rect 44571 18485 44605 18515
rect 44571 18417 44605 18443
rect 44571 18349 44605 18371
rect 44571 18281 44605 18299
rect 44571 18213 44605 18227
rect 44571 18145 44605 18155
rect 44571 18077 44605 18083
rect 44571 18009 44605 18011
rect 44571 17973 44605 17975
rect 44571 17901 44605 17907
rect 44571 17829 44605 17839
rect 44571 17757 44605 17771
rect 44571 17685 44605 17703
rect 44571 17613 44605 17635
rect 44571 17541 44605 17567
rect 44571 17469 44605 17499
rect 44571 17397 44605 17431
rect 44571 17343 44605 17363
rect 45029 18621 45063 18641
rect 45029 18553 45063 18587
rect 45029 18485 45063 18515
rect 45029 18417 45063 18443
rect 45029 18349 45063 18371
rect 45029 18281 45063 18299
rect 45029 18213 45063 18227
rect 45029 18145 45063 18155
rect 45029 18077 45063 18083
rect 45029 18009 45063 18011
rect 45029 17973 45063 17975
rect 45029 17901 45063 17907
rect 45029 17829 45063 17839
rect 45029 17757 45063 17771
rect 45029 17685 45063 17703
rect 45029 17613 45063 17635
rect 45029 17541 45063 17567
rect 45029 17469 45063 17499
rect 45029 17397 45063 17431
rect 45029 17262 45063 17363
rect 45487 18621 45521 18682
rect 45487 18553 45521 18587
rect 45487 18485 45521 18515
rect 45487 18417 45521 18443
rect 45487 18349 45521 18371
rect 45487 18281 45521 18299
rect 45487 18213 45521 18227
rect 45487 18145 45521 18155
rect 45487 18077 45521 18083
rect 45487 18009 45521 18011
rect 45487 17973 45521 17975
rect 45487 17901 45521 17907
rect 45487 17829 45521 17839
rect 45487 17757 45521 17771
rect 45487 17685 45521 17703
rect 45487 17613 45521 17635
rect 45487 17541 45521 17567
rect 45487 17469 45521 17499
rect 45487 17397 45521 17431
rect 45487 17343 45521 17363
rect 45945 18621 45979 18641
rect 45945 18553 45979 18587
rect 45945 18485 45979 18515
rect 45945 18417 45979 18443
rect 45945 18349 45979 18371
rect 45945 18281 45979 18299
rect 45945 18213 45979 18227
rect 45945 18145 45979 18155
rect 45945 18077 45979 18083
rect 45945 18009 45979 18011
rect 45945 17973 45979 17975
rect 45945 17901 45979 17907
rect 45945 17829 45979 17839
rect 45945 17757 45979 17771
rect 45945 17685 45979 17703
rect 45945 17613 45979 17635
rect 45945 17541 45979 17567
rect 45945 17469 45979 17499
rect 45945 17397 45979 17431
rect 45945 17262 45979 17363
rect 46403 18621 46437 18682
rect 46403 18553 46437 18587
rect 46403 18485 46437 18515
rect 46403 18417 46437 18443
rect 46403 18349 46437 18371
rect 46403 18281 46437 18299
rect 46403 18213 46437 18227
rect 46403 18145 46437 18155
rect 46403 18077 46437 18083
rect 46403 18009 46437 18011
rect 46403 17973 46437 17975
rect 46403 17901 46437 17907
rect 46403 17829 46437 17839
rect 46403 17757 46437 17771
rect 46403 17685 46437 17703
rect 46403 17613 46437 17635
rect 46403 17541 46437 17567
rect 46403 17469 46437 17499
rect 46403 17397 46437 17431
rect 46403 17343 46437 17363
rect 46861 18621 46895 18641
rect 46861 18553 46895 18587
rect 46861 18485 46895 18515
rect 46861 18417 46895 18443
rect 46861 18349 46895 18371
rect 46861 18281 46895 18299
rect 46861 18213 46895 18227
rect 46861 18145 46895 18155
rect 46861 18077 46895 18083
rect 46861 18009 46895 18011
rect 46861 17973 46895 17975
rect 46861 17901 46895 17907
rect 46861 17829 46895 17839
rect 46861 17757 46895 17771
rect 46861 17685 46895 17703
rect 46861 17613 46895 17635
rect 46861 17541 46895 17567
rect 46861 17469 46895 17499
rect 46861 17397 46895 17431
rect 46861 17262 46895 17363
rect 47319 18621 47353 18682
rect 47319 18553 47353 18587
rect 47319 18485 47353 18515
rect 47319 18417 47353 18443
rect 47319 18349 47353 18371
rect 47319 18281 47353 18299
rect 47319 18213 47353 18227
rect 47319 18145 47353 18155
rect 47319 18077 47353 18083
rect 47319 18009 47353 18011
rect 47319 17973 47353 17975
rect 47319 17901 47353 17907
rect 47319 17829 47353 17839
rect 47319 17757 47353 17771
rect 47319 17685 47353 17703
rect 47319 17613 47353 17635
rect 47319 17541 47353 17567
rect 47319 17469 47353 17499
rect 47319 17397 47353 17431
rect 47319 17343 47353 17363
rect 47777 18621 47811 18641
rect 47777 18553 47811 18587
rect 47777 18485 47811 18515
rect 47777 18417 47811 18443
rect 47777 18349 47811 18371
rect 47777 18281 47811 18299
rect 47777 18213 47811 18227
rect 47777 18145 47811 18155
rect 47777 18077 47811 18083
rect 47777 18009 47811 18011
rect 47777 17973 47811 17975
rect 47777 17901 47811 17907
rect 47777 17829 47811 17839
rect 47777 17757 47811 17771
rect 47777 17685 47811 17703
rect 47777 17613 47811 17635
rect 47777 17541 47811 17567
rect 47777 17469 47811 17499
rect 47777 17397 47811 17431
rect 47777 17262 47811 17363
rect 48235 18621 48269 18682
rect 48235 18553 48269 18587
rect 48235 18485 48269 18515
rect 48235 18417 48269 18443
rect 48235 18349 48269 18371
rect 48235 18281 48269 18299
rect 48235 18213 48269 18227
rect 48235 18145 48269 18155
rect 48235 18077 48269 18083
rect 48235 18009 48269 18011
rect 48235 17973 48269 17975
rect 48235 17901 48269 17907
rect 48235 17829 48269 17839
rect 48235 17757 48269 17771
rect 48235 17685 48269 17703
rect 48235 17613 48269 17635
rect 48235 17541 48269 17567
rect 48235 17469 48269 17499
rect 48235 17397 48269 17431
rect 48235 17343 48269 17363
rect 48693 18621 48727 18641
rect 48693 18553 48727 18587
rect 48693 18485 48727 18515
rect 48693 18417 48727 18443
rect 48693 18349 48727 18371
rect 48693 18281 48727 18299
rect 48693 18213 48727 18227
rect 48693 18145 48727 18155
rect 48693 18077 48727 18083
rect 48693 18009 48727 18011
rect 48693 17973 48727 17975
rect 48693 17901 48727 17907
rect 48693 17829 48727 17839
rect 48693 17757 48727 17771
rect 48693 17685 48727 17703
rect 48693 17613 48727 17635
rect 48693 17541 48727 17567
rect 48693 17469 48727 17499
rect 48693 17397 48727 17431
rect 48693 17262 48727 17363
rect 49151 18621 49185 18682
rect 49151 18553 49185 18587
rect 49151 18485 49185 18515
rect 49151 18417 49185 18443
rect 49151 18349 49185 18371
rect 49151 18281 49185 18299
rect 49151 18213 49185 18227
rect 49151 18145 49185 18155
rect 49151 18077 49185 18083
rect 49151 18009 49185 18011
rect 49151 17973 49185 17975
rect 49151 17901 49185 17907
rect 49151 17829 49185 17839
rect 49151 17757 49185 17771
rect 49151 17685 49185 17703
rect 49151 17613 49185 17635
rect 49151 17541 49185 17567
rect 49151 17469 49185 17499
rect 49151 17397 49185 17431
rect 49151 17343 49185 17363
rect 49609 18621 49643 18641
rect 49609 18553 49643 18587
rect 49609 18485 49643 18515
rect 49609 18417 49643 18443
rect 49609 18349 49643 18371
rect 49609 18281 49643 18299
rect 49609 18213 49643 18227
rect 49609 18145 49643 18155
rect 49609 18077 49643 18083
rect 49609 18009 49643 18011
rect 49609 17973 49643 17975
rect 49609 17901 49643 17907
rect 49609 17829 49643 17839
rect 49609 17757 49643 17771
rect 49609 17685 49643 17703
rect 49609 17613 49643 17635
rect 49609 17541 49643 17567
rect 49609 17469 49643 17499
rect 49609 17397 49643 17431
rect 49609 17262 49643 17363
rect 50067 18621 50101 18682
rect 50067 18553 50101 18587
rect 50067 18485 50101 18515
rect 50067 18417 50101 18443
rect 50067 18349 50101 18371
rect 50067 18281 50101 18299
rect 50067 18213 50101 18227
rect 50067 18145 50101 18155
rect 50067 18077 50101 18083
rect 50067 18009 50101 18011
rect 50067 17973 50101 17975
rect 50067 17901 50101 17907
rect 50067 17829 50101 17839
rect 50067 17757 50101 17771
rect 50067 17685 50101 17703
rect 50067 17613 50101 17635
rect 50067 17541 50101 17567
rect 50067 17469 50101 17499
rect 50067 17397 50101 17431
rect 50067 17343 50101 17363
rect 50525 18621 50559 18641
rect 50525 18553 50559 18587
rect 50525 18485 50559 18515
rect 50525 18417 50559 18443
rect 50525 18349 50559 18371
rect 50525 18281 50559 18299
rect 50525 18213 50559 18227
rect 50525 18145 50559 18155
rect 50525 18077 50559 18083
rect 50525 18009 50559 18011
rect 50525 17973 50559 17975
rect 50525 17901 50559 17907
rect 50525 17829 50559 17839
rect 50525 17757 50559 17771
rect 50525 17685 50559 17703
rect 50525 17613 50559 17635
rect 50525 17541 50559 17567
rect 50525 17469 50559 17499
rect 50525 17397 50559 17431
rect 50525 17262 50559 17363
rect 50983 18621 51017 18682
rect 50983 18553 51017 18587
rect 50983 18485 51017 18515
rect 50983 18417 51017 18443
rect 50983 18349 51017 18371
rect 50983 18281 51017 18299
rect 50983 18213 51017 18227
rect 50983 18145 51017 18155
rect 50983 18077 51017 18083
rect 50983 18009 51017 18011
rect 50983 17973 51017 17975
rect 50983 17901 51017 17907
rect 50983 17829 51017 17839
rect 50983 17757 51017 17771
rect 50983 17685 51017 17703
rect 50983 17613 51017 17635
rect 50983 17541 51017 17567
rect 50983 17469 51017 17499
rect 50983 17397 51017 17431
rect 50983 17343 51017 17363
rect 51441 18621 51475 18641
rect 51441 18553 51475 18587
rect 51441 18485 51475 18515
rect 51441 18417 51475 18443
rect 51441 18349 51475 18371
rect 51441 18281 51475 18299
rect 51441 18213 51475 18227
rect 51441 18145 51475 18155
rect 51441 18077 51475 18083
rect 51441 18009 51475 18011
rect 51441 17973 51475 17975
rect 51441 17901 51475 17907
rect 51441 17829 51475 17839
rect 51441 17757 51475 17771
rect 51441 17685 51475 17703
rect 51441 17613 51475 17635
rect 51441 17541 51475 17567
rect 51441 17469 51475 17499
rect 51441 17397 51475 17431
rect 51441 17262 51475 17363
rect 51899 18621 51933 18682
rect 51899 18553 51933 18587
rect 51899 18485 51933 18515
rect 51899 18417 51933 18443
rect 51899 18349 51933 18371
rect 51899 18281 51933 18299
rect 51899 18213 51933 18227
rect 51899 18145 51933 18155
rect 51899 18077 51933 18083
rect 51899 18009 51933 18011
rect 51899 17973 51933 17975
rect 51899 17901 51933 17907
rect 51899 17829 51933 17839
rect 51899 17757 51933 17771
rect 51899 17685 51933 17703
rect 51899 17613 51933 17635
rect 51899 17541 51933 17567
rect 51899 17469 51933 17499
rect 51899 17397 51933 17431
rect 51899 17343 51933 17363
rect 52357 18621 52391 18641
rect 52357 18553 52391 18587
rect 52357 18485 52391 18515
rect 52357 18417 52391 18443
rect 52357 18349 52391 18371
rect 52357 18281 52391 18299
rect 52357 18213 52391 18227
rect 52357 18145 52391 18155
rect 52357 18077 52391 18083
rect 52357 18009 52391 18011
rect 52357 17973 52391 17975
rect 52357 17901 52391 17907
rect 52357 17829 52391 17839
rect 52357 17757 52391 17771
rect 52357 17685 52391 17703
rect 52357 17613 52391 17635
rect 52357 17541 52391 17567
rect 52357 17469 52391 17499
rect 52357 17397 52391 17431
rect 52357 17262 52391 17363
rect 24830 17255 52438 17262
rect 24830 17221 34345 17255
rect 34379 17221 52438 17255
rect 24830 17202 52438 17221
rect 24830 17153 52438 17156
rect 24830 17143 25421 17153
rect 25455 17143 52438 17153
rect 24830 17109 25013 17143
rect 25047 17109 25413 17143
rect 25455 17119 25813 17143
rect 25447 17109 25813 17119
rect 25847 17109 26213 17143
rect 26247 17109 26613 17143
rect 26647 17109 27013 17143
rect 27047 17109 27413 17143
rect 27447 17109 27813 17143
rect 27847 17109 28213 17143
rect 28247 17109 28613 17143
rect 28647 17109 29013 17143
rect 29047 17109 29413 17143
rect 29447 17109 29813 17143
rect 29847 17109 30213 17143
rect 30247 17109 30613 17143
rect 30647 17109 31013 17143
rect 31047 17109 31413 17143
rect 31447 17109 31813 17143
rect 31847 17109 32213 17143
rect 32247 17109 32613 17143
rect 32647 17109 33013 17143
rect 33047 17109 33413 17143
rect 33447 17109 33813 17143
rect 33847 17109 34213 17143
rect 34247 17109 34613 17143
rect 34647 17109 35013 17143
rect 35047 17109 35413 17143
rect 35447 17109 35813 17143
rect 35847 17109 36213 17143
rect 36247 17109 36613 17143
rect 36647 17109 37013 17143
rect 37047 17109 37413 17143
rect 37447 17109 37813 17143
rect 37847 17109 38213 17143
rect 38247 17109 38613 17143
rect 38647 17109 39013 17143
rect 39047 17109 39413 17143
rect 39447 17109 39813 17143
rect 39847 17109 40213 17143
rect 40247 17109 40613 17143
rect 40647 17109 41013 17143
rect 41047 17109 41413 17143
rect 41447 17109 41813 17143
rect 41847 17109 42213 17143
rect 42247 17109 42613 17143
rect 42647 17109 43013 17143
rect 43047 17109 43413 17143
rect 43447 17109 43813 17143
rect 43847 17109 44213 17143
rect 44247 17109 44613 17143
rect 44647 17109 45013 17143
rect 45047 17109 45413 17143
rect 45447 17109 45813 17143
rect 45847 17109 46213 17143
rect 46247 17109 46613 17143
rect 46647 17109 47013 17143
rect 47047 17109 47413 17143
rect 47447 17109 47813 17143
rect 47847 17109 48213 17143
rect 48247 17109 48613 17143
rect 48647 17109 49013 17143
rect 49047 17109 49413 17143
rect 49447 17109 49813 17143
rect 49847 17109 50213 17143
rect 50247 17109 50613 17143
rect 50647 17109 51013 17143
rect 51047 17109 51413 17143
rect 51447 17109 51813 17143
rect 51847 17109 52213 17143
rect 52247 17109 52438 17143
rect 24830 17096 52438 17109
rect 24732 17009 52438 17022
rect 24732 16975 25013 17009
rect 25047 16975 25413 17009
rect 25447 16975 25813 17009
rect 25847 16975 26213 17009
rect 26247 16975 26613 17009
rect 26647 16975 27013 17009
rect 27047 16975 27413 17009
rect 27447 16975 27813 17009
rect 27847 16975 28213 17009
rect 28247 16975 28613 17009
rect 28647 16975 29013 17009
rect 29047 16975 29413 17009
rect 29447 16975 29813 17009
rect 29847 16975 30213 17009
rect 30247 16975 30613 17009
rect 30647 16975 31013 17009
rect 31047 16975 31413 17009
rect 31447 16975 31813 17009
rect 31847 16975 32213 17009
rect 32247 16975 32613 17009
rect 32647 16975 33013 17009
rect 33047 16975 33413 17009
rect 33447 16975 33813 17009
rect 33847 16975 34213 17009
rect 34247 16975 34613 17009
rect 34647 16975 35013 17009
rect 35047 16975 35413 17009
rect 35447 16975 35813 17009
rect 35847 16975 36213 17009
rect 36247 16975 36613 17009
rect 36647 16975 37013 17009
rect 37047 16975 37413 17009
rect 37447 16975 37813 17009
rect 37847 16975 38213 17009
rect 38247 16975 38613 17009
rect 38647 16975 39013 17009
rect 39047 16975 39413 17009
rect 39447 16975 39813 17009
rect 39847 16975 40213 17009
rect 40247 16975 40613 17009
rect 40647 16975 41013 17009
rect 41047 16975 41413 17009
rect 41447 16975 41813 17009
rect 41847 16975 42213 17009
rect 42247 16975 42613 17009
rect 42647 16975 43013 17009
rect 43047 16975 43413 17009
rect 43447 16975 43813 17009
rect 43847 16975 44213 17009
rect 44247 16975 44613 17009
rect 44647 16975 45013 17009
rect 45047 16975 45413 17009
rect 45447 16975 45813 17009
rect 45847 16975 46213 17009
rect 46247 16975 46613 17009
rect 46647 16975 47013 17009
rect 47047 16975 47413 17009
rect 47447 16975 47813 17009
rect 47847 16975 48213 17009
rect 48247 16975 48613 17009
rect 48647 16975 49013 17009
rect 49047 16975 49413 17009
rect 49447 16975 49813 17009
rect 49847 16975 50213 17009
rect 50247 16975 50613 17009
rect 50647 16975 51013 17009
rect 51047 16975 51413 17009
rect 51447 16975 51813 17009
rect 51847 16975 52213 17009
rect 52247 16975 52438 17009
rect 24732 16962 52438 16975
rect 43862 15129 46302 15142
rect 43862 15095 44045 15129
rect 44079 15095 44245 15129
rect 44279 15095 44445 15129
rect 44479 15095 44645 15129
rect 44679 15095 44845 15129
rect 44879 15095 45045 15129
rect 45079 15095 45245 15129
rect 45279 15095 45445 15129
rect 45479 15095 45645 15129
rect 45679 15095 45845 15129
rect 45879 15095 46045 15129
rect 46079 15095 46302 15129
rect 43862 15082 46302 15095
rect 46606 15129 49046 15142
rect 46606 15095 46789 15129
rect 46823 15095 46989 15129
rect 47023 15095 47189 15129
rect 47223 15095 47389 15129
rect 47423 15095 47589 15129
rect 47623 15095 47789 15129
rect 47823 15095 47989 15129
rect 48023 15095 48189 15129
rect 48223 15095 48389 15129
rect 48423 15095 48589 15129
rect 48623 15095 48789 15129
rect 48823 15095 49046 15129
rect 46606 15082 49046 15095
rect 49350 15129 51790 15142
rect 49350 15095 49533 15129
rect 49567 15095 49733 15129
rect 49767 15095 49933 15129
rect 49967 15095 50133 15129
rect 50167 15095 50333 15129
rect 50367 15095 50533 15129
rect 50567 15095 50733 15129
rect 50767 15095 50933 15129
rect 50967 15095 51133 15129
rect 51167 15095 51333 15129
rect 51367 15095 51533 15129
rect 51567 15095 51790 15129
rect 49350 15082 51790 15095
rect 44774 14163 45390 14202
rect 44774 14061 44861 14163
rect 45303 14061 45390 14163
rect 44774 13262 45390 14061
rect 45870 13917 46302 14307
rect 47518 14163 48134 14202
rect 47518 14061 47605 14163
rect 48047 14061 48134 14163
rect 47518 13262 48134 14061
rect 48614 13917 49046 14307
rect 50262 14163 50878 14202
rect 50262 14061 50349 14163
rect 50791 14061 50878 14163
rect 50262 13262 50878 14061
rect 51358 13917 51790 14307
rect 43862 13249 46302 13262
rect 43862 13215 44045 13249
rect 44079 13215 44245 13249
rect 44279 13215 44445 13249
rect 44479 13215 44645 13249
rect 44679 13215 44845 13249
rect 44879 13215 45045 13249
rect 45079 13215 45245 13249
rect 45279 13215 45445 13249
rect 45479 13215 45645 13249
rect 45679 13215 45845 13249
rect 45879 13215 46045 13249
rect 46079 13215 46302 13249
rect 43862 13202 46302 13215
rect 46606 13249 49046 13262
rect 46606 13215 46789 13249
rect 46823 13215 46989 13249
rect 47023 13215 47189 13249
rect 47223 13215 47389 13249
rect 47423 13215 47589 13249
rect 47623 13215 47789 13249
rect 47823 13215 47989 13249
rect 48023 13215 48189 13249
rect 48223 13215 48389 13249
rect 48423 13215 48589 13249
rect 48623 13215 48789 13249
rect 48823 13215 49046 13249
rect 46606 13202 49046 13215
rect 49350 13249 51790 13262
rect 49350 13215 49533 13249
rect 49567 13215 49733 13249
rect 49767 13215 49933 13249
rect 49967 13215 50133 13249
rect 50167 13215 50333 13249
rect 50367 13215 50533 13249
rect 50567 13215 50733 13249
rect 50767 13215 50933 13249
rect 50967 13215 51133 13249
rect 51167 13215 51333 13249
rect 51367 13215 51533 13249
rect 51567 13215 51790 13249
rect 49350 13202 51790 13215
rect 43764 11369 46204 11382
rect 43764 11335 43947 11369
rect 43981 11335 44147 11369
rect 44181 11335 44347 11369
rect 44381 11335 44547 11369
rect 44581 11335 44747 11369
rect 44781 11335 44947 11369
rect 44981 11335 45147 11369
rect 45181 11335 45347 11369
rect 45381 11335 45547 11369
rect 45581 11335 45747 11369
rect 45781 11335 45947 11369
rect 45981 11335 46204 11369
rect 43764 11322 46204 11335
rect 46508 11369 48948 11382
rect 46508 11335 46691 11369
rect 46725 11335 46891 11369
rect 46925 11335 47091 11369
rect 47125 11335 47291 11369
rect 47325 11335 47491 11369
rect 47525 11335 47691 11369
rect 47725 11335 47891 11369
rect 47925 11335 48091 11369
rect 48125 11335 48291 11369
rect 48325 11335 48491 11369
rect 48525 11335 48691 11369
rect 48725 11335 48948 11369
rect 46508 11322 48948 11335
rect 49252 11369 51692 11382
rect 49252 11335 49435 11369
rect 49469 11335 49635 11369
rect 49669 11335 49835 11369
rect 49869 11335 50035 11369
rect 50069 11335 50235 11369
rect 50269 11335 50435 11369
rect 50469 11335 50635 11369
rect 50669 11335 50835 11369
rect 50869 11335 51035 11369
rect 51069 11335 51235 11369
rect 51269 11335 51435 11369
rect 51469 11335 51692 11369
rect 49252 11322 51692 11335
rect 44676 10403 45292 10442
rect 44676 10301 44763 10403
rect 45205 10301 45292 10403
rect 44676 9502 45292 10301
rect 45772 10157 46204 10547
rect 47420 10403 48036 10442
rect 47420 10301 47507 10403
rect 47949 10301 48036 10403
rect 47420 9502 48036 10301
rect 48516 10157 48948 10547
rect 50164 10403 50780 10442
rect 50164 10301 50251 10403
rect 50693 10301 50780 10403
rect 50164 9502 50780 10301
rect 51260 10157 51692 10547
rect 43764 9489 46204 9502
rect 43764 9455 43947 9489
rect 43981 9455 44147 9489
rect 44181 9455 44347 9489
rect 44381 9455 44547 9489
rect 44581 9455 44747 9489
rect 44781 9455 44947 9489
rect 44981 9455 45147 9489
rect 45181 9455 45347 9489
rect 45381 9455 45547 9489
rect 45581 9455 45747 9489
rect 45781 9455 45947 9489
rect 45981 9455 46204 9489
rect 43764 9442 46204 9455
rect 46508 9489 48948 9502
rect 46508 9455 46691 9489
rect 46725 9455 46891 9489
rect 46925 9455 47091 9489
rect 47125 9455 47291 9489
rect 47325 9455 47491 9489
rect 47525 9455 47691 9489
rect 47725 9455 47891 9489
rect 47925 9455 48091 9489
rect 48125 9455 48291 9489
rect 48325 9455 48491 9489
rect 48525 9455 48691 9489
rect 48725 9455 48948 9489
rect 46508 9442 48948 9455
rect 49252 9489 51692 9502
rect 49252 9455 49435 9489
rect 49469 9455 49635 9489
rect 49669 9455 49835 9489
rect 49869 9455 50035 9489
rect 50069 9455 50235 9489
rect 50269 9455 50435 9489
rect 50469 9455 50635 9489
rect 50669 9455 50835 9489
rect 50869 9455 51035 9489
rect 51069 9455 51235 9489
rect 51269 9455 51435 9489
rect 51469 9455 51692 9489
rect 49252 9442 51692 9455
rect 44548 7609 46988 7622
rect 44548 7575 44731 7609
rect 44765 7575 44931 7609
rect 44965 7575 45131 7609
rect 45165 7575 45331 7609
rect 45365 7575 45531 7609
rect 45565 7575 45731 7609
rect 45765 7575 45931 7609
rect 45965 7575 46131 7609
rect 46165 7575 46331 7609
rect 46365 7575 46531 7609
rect 46565 7575 46731 7609
rect 46765 7575 46988 7609
rect 44548 7562 46988 7575
rect 47292 7609 49732 7622
rect 47292 7575 47475 7609
rect 47509 7575 47675 7609
rect 47709 7575 47875 7609
rect 47909 7575 48075 7609
rect 48109 7575 48275 7609
rect 48309 7575 48475 7609
rect 48509 7575 48675 7609
rect 48709 7575 48875 7609
rect 48909 7575 49075 7609
rect 49109 7575 49275 7609
rect 49309 7575 49475 7609
rect 49509 7575 49732 7609
rect 47292 7562 49732 7575
rect 50036 7609 52476 7622
rect 50036 7575 50219 7609
rect 50253 7575 50419 7609
rect 50453 7575 50619 7609
rect 50653 7575 50819 7609
rect 50853 7575 51019 7609
rect 51053 7575 51219 7609
rect 51253 7575 51419 7609
rect 51453 7575 51619 7609
rect 51653 7575 51819 7609
rect 51853 7575 52019 7609
rect 52053 7575 52219 7609
rect 52253 7575 52476 7609
rect 50036 7562 52476 7575
rect 45460 6643 46076 6682
rect 45460 6541 45547 6643
rect 45989 6541 46076 6643
rect 45460 5742 46076 6541
rect 46556 6397 46988 6787
rect 48204 6643 48820 6682
rect 48204 6541 48291 6643
rect 48733 6541 48820 6643
rect 48204 5742 48820 6541
rect 49300 6397 49732 6787
rect 50948 6643 51564 6682
rect 50948 6541 51035 6643
rect 51477 6541 51564 6643
rect 50948 5742 51564 6541
rect 52044 6397 52476 6787
rect 44548 5729 46988 5742
rect 44548 5695 44731 5729
rect 44765 5695 44931 5729
rect 44965 5695 45131 5729
rect 45165 5695 45331 5729
rect 45365 5695 45531 5729
rect 45565 5695 45731 5729
rect 45765 5695 45931 5729
rect 45965 5695 46131 5729
rect 46165 5695 46331 5729
rect 46365 5695 46531 5729
rect 46565 5695 46731 5729
rect 46765 5695 46988 5729
rect 44548 5682 46988 5695
rect 47292 5729 49732 5742
rect 47292 5695 47475 5729
rect 47509 5695 47675 5729
rect 47709 5695 47875 5729
rect 47909 5695 48075 5729
rect 48109 5695 48275 5729
rect 48309 5695 48475 5729
rect 48509 5695 48675 5729
rect 48709 5695 48875 5729
rect 48909 5695 49075 5729
rect 49109 5695 49275 5729
rect 49309 5695 49475 5729
rect 49509 5695 49732 5729
rect 47292 5682 49732 5695
rect 50036 5729 52476 5742
rect 50036 5695 50219 5729
rect 50253 5695 50419 5729
rect 50453 5695 50619 5729
rect 50653 5695 50819 5729
rect 50853 5695 51019 5729
rect 51053 5695 51219 5729
rect 51253 5695 51419 5729
rect 51453 5695 51619 5729
rect 51653 5695 51819 5729
rect 51853 5695 52019 5729
rect 52053 5695 52219 5729
rect 52253 5695 52476 5729
rect 50036 5682 52476 5695
<< viali >>
rect 6101 48935 6135 48969
rect 6501 48935 6535 48969
rect 6901 48935 6935 48969
rect 7301 48935 7335 48969
rect 7701 48935 7735 48969
rect 8101 48935 8135 48969
rect 8501 48935 8535 48969
rect 8901 48935 8935 48969
rect 9301 48935 9335 48969
rect 9701 48935 9735 48969
rect 10101 48935 10135 48969
rect 10501 48935 10535 48969
rect 10901 48935 10935 48969
rect 11301 48935 11335 48969
rect 11701 48935 11735 48969
rect 12101 48935 12135 48969
rect 12501 48935 12535 48969
rect 12901 48935 12935 48969
rect 13549 48935 13583 48969
rect 13949 48935 13983 48969
rect 14349 48935 14383 48969
rect 14749 48935 14783 48969
rect 15149 48935 15183 48969
rect 15549 48935 15583 48969
rect 15949 48935 15983 48969
rect 16349 48935 16383 48969
rect 16749 48935 16783 48969
rect 17149 48935 17183 48969
rect 17549 48935 17583 48969
rect 17949 48935 17983 48969
rect 18349 48935 18383 48969
rect 18749 48935 18783 48969
rect 19149 48935 19183 48969
rect 19549 48935 19583 48969
rect 19949 48935 19983 48969
rect 20349 48935 20383 48969
rect 21015 48935 21049 48969
rect 21215 48935 21249 48969
rect 21415 48935 21449 48969
rect 21615 48935 21649 48969
rect 21815 48935 21849 48969
rect 22015 48935 22049 48969
rect 22215 48935 22249 48969
rect 22415 48935 22449 48969
rect 22615 48935 22649 48969
rect 22815 48935 22849 48969
rect 23015 48935 23049 48969
rect 24101 48935 24135 48969
rect 25013 48935 25047 48969
rect 25413 48935 25447 48969
rect 25813 48935 25847 48969
rect 26213 48935 26247 48969
rect 26613 48935 26647 48969
rect 27013 48935 27047 48969
rect 27413 48935 27447 48969
rect 27813 48935 27847 48969
rect 28213 48935 28247 48969
rect 28613 48935 28647 48969
rect 29013 48935 29047 48969
rect 29413 48935 29447 48969
rect 29813 48935 29847 48969
rect 30213 48935 30247 48969
rect 30613 48935 30647 48969
rect 31013 48935 31047 48969
rect 31413 48935 31447 48969
rect 31813 48935 31847 48969
rect 32213 48935 32247 48969
rect 32613 48935 32647 48969
rect 33013 48935 33047 48969
rect 33413 48935 33447 48969
rect 33813 48935 33847 48969
rect 34213 48935 34247 48969
rect 34613 48935 34647 48969
rect 35013 48935 35047 48969
rect 35413 48935 35447 48969
rect 35813 48935 35847 48969
rect 36213 48935 36247 48969
rect 36613 48935 36647 48969
rect 37013 48935 37047 48969
rect 37413 48935 37447 48969
rect 37813 48935 37847 48969
rect 38213 48935 38247 48969
rect 38613 48935 38647 48969
rect 39013 48935 39047 48969
rect 39413 48935 39447 48969
rect 39813 48935 39847 48969
rect 40213 48935 40247 48969
rect 40613 48935 40647 48969
rect 41013 48935 41047 48969
rect 41413 48935 41447 48969
rect 41813 48935 41847 48969
rect 42213 48935 42247 48969
rect 42613 48935 42647 48969
rect 43013 48935 43047 48969
rect 43413 48935 43447 48969
rect 43813 48935 43847 48969
rect 44213 48935 44247 48969
rect 44613 48935 44647 48969
rect 45013 48935 45047 48969
rect 45413 48935 45447 48969
rect 45813 48935 45847 48969
rect 46213 48935 46247 48969
rect 46613 48935 46647 48969
rect 47013 48935 47047 48969
rect 47413 48935 47447 48969
rect 47813 48935 47847 48969
rect 48213 48935 48247 48969
rect 48613 48935 48647 48969
rect 49013 48935 49047 48969
rect 49413 48935 49447 48969
rect 49813 48935 49847 48969
rect 50213 48935 50247 48969
rect 50613 48935 50647 48969
rect 51013 48935 51047 48969
rect 51413 48935 51447 48969
rect 51813 48935 51847 48969
rect 52213 48935 52247 48969
rect 20851 48163 21245 48701
rect 22858 48163 23252 48701
rect 24877 48667 24911 48701
rect 24877 48599 24911 48629
rect 24877 48595 24911 48599
rect 24877 48531 24911 48557
rect 24877 48523 24911 48531
rect 20851 47203 21245 47741
rect 22858 47203 23252 47741
rect 23930 48429 23964 48449
rect 23930 48415 23964 48429
rect 23930 48361 23964 48377
rect 23930 48343 23964 48361
rect 23930 48293 23964 48305
rect 23930 48271 23964 48293
rect 23930 48225 23964 48233
rect 23930 48199 23964 48225
rect 23930 48157 23964 48161
rect 23930 48127 23964 48157
rect 23930 48055 23964 48089
rect 23930 47987 23964 48017
rect 23930 47983 23964 47987
rect 23930 47919 23964 47945
rect 23930 47911 23964 47919
rect 23930 47851 23964 47873
rect 23930 47839 23964 47851
rect 23930 47783 23964 47801
rect 23930 47767 23964 47783
rect 23930 47715 23964 47729
rect 23930 47695 23964 47715
rect 24388 48429 24422 48449
rect 24388 48415 24422 48429
rect 24388 48361 24422 48377
rect 24388 48343 24422 48361
rect 24388 48293 24422 48305
rect 24388 48271 24422 48293
rect 24388 48225 24422 48233
rect 24388 48199 24422 48225
rect 24388 48157 24422 48161
rect 24388 48127 24422 48157
rect 24388 48055 24422 48089
rect 24388 47987 24422 48017
rect 24388 47983 24422 47987
rect 24388 47919 24422 47945
rect 24388 47911 24422 47919
rect 24388 47851 24422 47873
rect 24388 47839 24422 47851
rect 24388 47783 24422 47801
rect 24388 47767 24422 47783
rect 24388 47715 24422 47729
rect 24388 47695 24422 47715
rect 24877 48463 24911 48485
rect 24877 48451 24911 48463
rect 24877 48395 24911 48413
rect 24877 48379 24911 48395
rect 24877 48327 24911 48341
rect 24877 48307 24911 48327
rect 24877 48259 24911 48269
rect 24877 48235 24911 48259
rect 24877 48191 24911 48197
rect 24877 48163 24911 48191
rect 24877 48123 24911 48125
rect 24877 48091 24911 48123
rect 24877 48021 24911 48053
rect 24877 48019 24911 48021
rect 24877 47953 24911 47981
rect 24877 47947 24911 47953
rect 24877 47885 24911 47909
rect 24877 47875 24911 47885
rect 24877 47817 24911 47837
rect 24877 47803 24911 47817
rect 24877 47749 24911 47765
rect 24877 47731 24911 47749
rect 24877 47681 24911 47693
rect 24877 47659 24911 47681
rect 24877 47613 24911 47621
rect 24877 47587 24911 47613
rect 24877 47545 24911 47549
rect 24877 47515 24911 47545
rect 24877 47443 24911 47477
rect 25335 48667 25369 48701
rect 25335 48599 25369 48629
rect 25335 48595 25369 48599
rect 25335 48531 25369 48557
rect 25335 48523 25369 48531
rect 25335 48463 25369 48485
rect 25335 48451 25369 48463
rect 25335 48395 25369 48413
rect 25335 48379 25369 48395
rect 25335 48327 25369 48341
rect 25335 48307 25369 48327
rect 25335 48259 25369 48269
rect 25335 48235 25369 48259
rect 25335 48191 25369 48197
rect 25335 48163 25369 48191
rect 25335 48123 25369 48125
rect 25335 48091 25369 48123
rect 25335 48021 25369 48053
rect 25335 48019 25369 48021
rect 25335 47953 25369 47981
rect 25335 47947 25369 47953
rect 25335 47885 25369 47909
rect 25335 47875 25369 47885
rect 25335 47817 25369 47837
rect 25335 47803 25369 47817
rect 25335 47749 25369 47765
rect 25335 47731 25369 47749
rect 25335 47681 25369 47693
rect 25335 47659 25369 47681
rect 25335 47613 25369 47621
rect 25335 47587 25369 47613
rect 25335 47545 25369 47549
rect 25335 47515 25369 47545
rect 25335 47443 25369 47477
rect 25793 48667 25827 48701
rect 25793 48599 25827 48629
rect 25793 48595 25827 48599
rect 25793 48531 25827 48557
rect 25793 48523 25827 48531
rect 25793 48463 25827 48485
rect 25793 48451 25827 48463
rect 25793 48395 25827 48413
rect 25793 48379 25827 48395
rect 25793 48327 25827 48341
rect 25793 48307 25827 48327
rect 25793 48259 25827 48269
rect 25793 48235 25827 48259
rect 25793 48191 25827 48197
rect 25793 48163 25827 48191
rect 25793 48123 25827 48125
rect 25793 48091 25827 48123
rect 25793 48021 25827 48053
rect 25793 48019 25827 48021
rect 25793 47953 25827 47981
rect 25793 47947 25827 47953
rect 25793 47885 25827 47909
rect 25793 47875 25827 47885
rect 25793 47817 25827 47837
rect 25793 47803 25827 47817
rect 25793 47749 25827 47765
rect 25793 47731 25827 47749
rect 25793 47681 25827 47693
rect 25793 47659 25827 47681
rect 25793 47613 25827 47621
rect 25793 47587 25827 47613
rect 25793 47545 25827 47549
rect 25793 47515 25827 47545
rect 25793 47443 25827 47477
rect 26251 48667 26285 48701
rect 26251 48599 26285 48629
rect 26251 48595 26285 48599
rect 26251 48531 26285 48557
rect 26251 48523 26285 48531
rect 26251 48463 26285 48485
rect 26251 48451 26285 48463
rect 26251 48395 26285 48413
rect 26251 48379 26285 48395
rect 26251 48327 26285 48341
rect 26251 48307 26285 48327
rect 26251 48259 26285 48269
rect 26251 48235 26285 48259
rect 26251 48191 26285 48197
rect 26251 48163 26285 48191
rect 26251 48123 26285 48125
rect 26251 48091 26285 48123
rect 26251 48021 26285 48053
rect 26251 48019 26285 48021
rect 26251 47953 26285 47981
rect 26251 47947 26285 47953
rect 26251 47885 26285 47909
rect 26251 47875 26285 47885
rect 26251 47817 26285 47837
rect 26251 47803 26285 47817
rect 26251 47749 26285 47765
rect 26251 47731 26285 47749
rect 26251 47681 26285 47693
rect 26251 47659 26285 47681
rect 26251 47613 26285 47621
rect 26251 47587 26285 47613
rect 26251 47545 26285 47549
rect 26251 47515 26285 47545
rect 26251 47443 26285 47477
rect 26709 48667 26743 48701
rect 26709 48599 26743 48629
rect 26709 48595 26743 48599
rect 26709 48531 26743 48557
rect 26709 48523 26743 48531
rect 26709 48463 26743 48485
rect 26709 48451 26743 48463
rect 26709 48395 26743 48413
rect 26709 48379 26743 48395
rect 26709 48327 26743 48341
rect 26709 48307 26743 48327
rect 26709 48259 26743 48269
rect 26709 48235 26743 48259
rect 26709 48191 26743 48197
rect 26709 48163 26743 48191
rect 26709 48123 26743 48125
rect 26709 48091 26743 48123
rect 26709 48021 26743 48053
rect 26709 48019 26743 48021
rect 26709 47953 26743 47981
rect 26709 47947 26743 47953
rect 26709 47885 26743 47909
rect 26709 47875 26743 47885
rect 26709 47817 26743 47837
rect 26709 47803 26743 47817
rect 26709 47749 26743 47765
rect 26709 47731 26743 47749
rect 26709 47681 26743 47693
rect 26709 47659 26743 47681
rect 26709 47613 26743 47621
rect 26709 47587 26743 47613
rect 26709 47545 26743 47549
rect 26709 47515 26743 47545
rect 26709 47443 26743 47477
rect 27167 48667 27201 48701
rect 27167 48599 27201 48629
rect 27167 48595 27201 48599
rect 27167 48531 27201 48557
rect 27167 48523 27201 48531
rect 27167 48463 27201 48485
rect 27167 48451 27201 48463
rect 27167 48395 27201 48413
rect 27167 48379 27201 48395
rect 27167 48327 27201 48341
rect 27167 48307 27201 48327
rect 27167 48259 27201 48269
rect 27167 48235 27201 48259
rect 27167 48191 27201 48197
rect 27167 48163 27201 48191
rect 27167 48123 27201 48125
rect 27167 48091 27201 48123
rect 27167 48021 27201 48053
rect 27167 48019 27201 48021
rect 27167 47953 27201 47981
rect 27167 47947 27201 47953
rect 27167 47885 27201 47909
rect 27167 47875 27201 47885
rect 27167 47817 27201 47837
rect 27167 47803 27201 47817
rect 27167 47749 27201 47765
rect 27167 47731 27201 47749
rect 27167 47681 27201 47693
rect 27167 47659 27201 47681
rect 27167 47613 27201 47621
rect 27167 47587 27201 47613
rect 27167 47545 27201 47549
rect 27167 47515 27201 47545
rect 27167 47443 27201 47477
rect 27625 48667 27659 48701
rect 27625 48599 27659 48629
rect 27625 48595 27659 48599
rect 27625 48531 27659 48557
rect 27625 48523 27659 48531
rect 27625 48463 27659 48485
rect 27625 48451 27659 48463
rect 27625 48395 27659 48413
rect 27625 48379 27659 48395
rect 27625 48327 27659 48341
rect 27625 48307 27659 48327
rect 27625 48259 27659 48269
rect 27625 48235 27659 48259
rect 27625 48191 27659 48197
rect 27625 48163 27659 48191
rect 27625 48123 27659 48125
rect 27625 48091 27659 48123
rect 27625 48021 27659 48053
rect 27625 48019 27659 48021
rect 27625 47953 27659 47981
rect 27625 47947 27659 47953
rect 27625 47885 27659 47909
rect 27625 47875 27659 47885
rect 27625 47817 27659 47837
rect 27625 47803 27659 47817
rect 27625 47749 27659 47765
rect 27625 47731 27659 47749
rect 27625 47681 27659 47693
rect 27625 47659 27659 47681
rect 27625 47613 27659 47621
rect 27625 47587 27659 47613
rect 27625 47545 27659 47549
rect 27625 47515 27659 47545
rect 27625 47443 27659 47477
rect 28083 48667 28117 48701
rect 28083 48599 28117 48629
rect 28083 48595 28117 48599
rect 28083 48531 28117 48557
rect 28083 48523 28117 48531
rect 28083 48463 28117 48485
rect 28083 48451 28117 48463
rect 28083 48395 28117 48413
rect 28083 48379 28117 48395
rect 28083 48327 28117 48341
rect 28083 48307 28117 48327
rect 28083 48259 28117 48269
rect 28083 48235 28117 48259
rect 28083 48191 28117 48197
rect 28083 48163 28117 48191
rect 28083 48123 28117 48125
rect 28083 48091 28117 48123
rect 28083 48021 28117 48053
rect 28083 48019 28117 48021
rect 28083 47953 28117 47981
rect 28083 47947 28117 47953
rect 28083 47885 28117 47909
rect 28083 47875 28117 47885
rect 28083 47817 28117 47837
rect 28083 47803 28117 47817
rect 28083 47749 28117 47765
rect 28083 47731 28117 47749
rect 28083 47681 28117 47693
rect 28083 47659 28117 47681
rect 28083 47613 28117 47621
rect 28083 47587 28117 47613
rect 28083 47545 28117 47549
rect 28083 47515 28117 47545
rect 28083 47443 28117 47477
rect 28541 48667 28575 48701
rect 28541 48599 28575 48629
rect 28541 48595 28575 48599
rect 28541 48531 28575 48557
rect 28541 48523 28575 48531
rect 28541 48463 28575 48485
rect 28541 48451 28575 48463
rect 28541 48395 28575 48413
rect 28541 48379 28575 48395
rect 28541 48327 28575 48341
rect 28541 48307 28575 48327
rect 28541 48259 28575 48269
rect 28541 48235 28575 48259
rect 28541 48191 28575 48197
rect 28541 48163 28575 48191
rect 28541 48123 28575 48125
rect 28541 48091 28575 48123
rect 28541 48021 28575 48053
rect 28541 48019 28575 48021
rect 28541 47953 28575 47981
rect 28541 47947 28575 47953
rect 28541 47885 28575 47909
rect 28541 47875 28575 47885
rect 28541 47817 28575 47837
rect 28541 47803 28575 47817
rect 28541 47749 28575 47765
rect 28541 47731 28575 47749
rect 28541 47681 28575 47693
rect 28541 47659 28575 47681
rect 28541 47613 28575 47621
rect 28541 47587 28575 47613
rect 28541 47545 28575 47549
rect 28541 47515 28575 47545
rect 28541 47443 28575 47477
rect 28999 48667 29033 48701
rect 28999 48599 29033 48629
rect 28999 48595 29033 48599
rect 28999 48531 29033 48557
rect 28999 48523 29033 48531
rect 28999 48463 29033 48485
rect 28999 48451 29033 48463
rect 28999 48395 29033 48413
rect 28999 48379 29033 48395
rect 28999 48327 29033 48341
rect 28999 48307 29033 48327
rect 28999 48259 29033 48269
rect 28999 48235 29033 48259
rect 28999 48191 29033 48197
rect 28999 48163 29033 48191
rect 28999 48123 29033 48125
rect 28999 48091 29033 48123
rect 28999 48021 29033 48053
rect 28999 48019 29033 48021
rect 28999 47953 29033 47981
rect 28999 47947 29033 47953
rect 28999 47885 29033 47909
rect 28999 47875 29033 47885
rect 28999 47817 29033 47837
rect 28999 47803 29033 47817
rect 28999 47749 29033 47765
rect 28999 47731 29033 47749
rect 28999 47681 29033 47693
rect 28999 47659 29033 47681
rect 28999 47613 29033 47621
rect 28999 47587 29033 47613
rect 28999 47545 29033 47549
rect 28999 47515 29033 47545
rect 28999 47443 29033 47477
rect 29457 48667 29491 48701
rect 29457 48599 29491 48629
rect 29457 48595 29491 48599
rect 29457 48531 29491 48557
rect 29457 48523 29491 48531
rect 29457 48463 29491 48485
rect 29457 48451 29491 48463
rect 29457 48395 29491 48413
rect 29457 48379 29491 48395
rect 29457 48327 29491 48341
rect 29457 48307 29491 48327
rect 29457 48259 29491 48269
rect 29457 48235 29491 48259
rect 29457 48191 29491 48197
rect 29457 48163 29491 48191
rect 29457 48123 29491 48125
rect 29457 48091 29491 48123
rect 29457 48021 29491 48053
rect 29457 48019 29491 48021
rect 29457 47953 29491 47981
rect 29457 47947 29491 47953
rect 29457 47885 29491 47909
rect 29457 47875 29491 47885
rect 29457 47817 29491 47837
rect 29457 47803 29491 47817
rect 29457 47749 29491 47765
rect 29457 47731 29491 47749
rect 29457 47681 29491 47693
rect 29457 47659 29491 47681
rect 29457 47613 29491 47621
rect 29457 47587 29491 47613
rect 29457 47545 29491 47549
rect 29457 47515 29491 47545
rect 29457 47443 29491 47477
rect 29915 48667 29949 48701
rect 29915 48599 29949 48629
rect 29915 48595 29949 48599
rect 29915 48531 29949 48557
rect 29915 48523 29949 48531
rect 29915 48463 29949 48485
rect 29915 48451 29949 48463
rect 29915 48395 29949 48413
rect 29915 48379 29949 48395
rect 29915 48327 29949 48341
rect 29915 48307 29949 48327
rect 29915 48259 29949 48269
rect 29915 48235 29949 48259
rect 29915 48191 29949 48197
rect 29915 48163 29949 48191
rect 29915 48123 29949 48125
rect 29915 48091 29949 48123
rect 29915 48021 29949 48053
rect 29915 48019 29949 48021
rect 29915 47953 29949 47981
rect 29915 47947 29949 47953
rect 29915 47885 29949 47909
rect 29915 47875 29949 47885
rect 29915 47817 29949 47837
rect 29915 47803 29949 47817
rect 29915 47749 29949 47765
rect 29915 47731 29949 47749
rect 29915 47681 29949 47693
rect 29915 47659 29949 47681
rect 29915 47613 29949 47621
rect 29915 47587 29949 47613
rect 29915 47545 29949 47549
rect 29915 47515 29949 47545
rect 29915 47443 29949 47477
rect 30373 48667 30407 48701
rect 30373 48599 30407 48629
rect 30373 48595 30407 48599
rect 30373 48531 30407 48557
rect 30373 48523 30407 48531
rect 30373 48463 30407 48485
rect 30373 48451 30407 48463
rect 30373 48395 30407 48413
rect 30373 48379 30407 48395
rect 30373 48327 30407 48341
rect 30373 48307 30407 48327
rect 30373 48259 30407 48269
rect 30373 48235 30407 48259
rect 30373 48191 30407 48197
rect 30373 48163 30407 48191
rect 30373 48123 30407 48125
rect 30373 48091 30407 48123
rect 30373 48021 30407 48053
rect 30373 48019 30407 48021
rect 30373 47953 30407 47981
rect 30373 47947 30407 47953
rect 30373 47885 30407 47909
rect 30373 47875 30407 47885
rect 30373 47817 30407 47837
rect 30373 47803 30407 47817
rect 30373 47749 30407 47765
rect 30373 47731 30407 47749
rect 30373 47681 30407 47693
rect 30373 47659 30407 47681
rect 30373 47613 30407 47621
rect 30373 47587 30407 47613
rect 30373 47545 30407 47549
rect 30373 47515 30407 47545
rect 30373 47443 30407 47477
rect 30831 48667 30865 48701
rect 30831 48599 30865 48629
rect 30831 48595 30865 48599
rect 30831 48531 30865 48557
rect 30831 48523 30865 48531
rect 30831 48463 30865 48485
rect 30831 48451 30865 48463
rect 30831 48395 30865 48413
rect 30831 48379 30865 48395
rect 30831 48327 30865 48341
rect 30831 48307 30865 48327
rect 30831 48259 30865 48269
rect 30831 48235 30865 48259
rect 30831 48191 30865 48197
rect 30831 48163 30865 48191
rect 30831 48123 30865 48125
rect 30831 48091 30865 48123
rect 30831 48021 30865 48053
rect 30831 48019 30865 48021
rect 30831 47953 30865 47981
rect 30831 47947 30865 47953
rect 30831 47885 30865 47909
rect 30831 47875 30865 47885
rect 30831 47817 30865 47837
rect 30831 47803 30865 47817
rect 30831 47749 30865 47765
rect 30831 47731 30865 47749
rect 30831 47681 30865 47693
rect 30831 47659 30865 47681
rect 30831 47613 30865 47621
rect 30831 47587 30865 47613
rect 30831 47545 30865 47549
rect 30831 47515 30865 47545
rect 30831 47443 30865 47477
rect 31289 48667 31323 48701
rect 31289 48599 31323 48629
rect 31289 48595 31323 48599
rect 31289 48531 31323 48557
rect 31289 48523 31323 48531
rect 31289 48463 31323 48485
rect 31289 48451 31323 48463
rect 31289 48395 31323 48413
rect 31289 48379 31323 48395
rect 31289 48327 31323 48341
rect 31289 48307 31323 48327
rect 31289 48259 31323 48269
rect 31289 48235 31323 48259
rect 31289 48191 31323 48197
rect 31289 48163 31323 48191
rect 31289 48123 31323 48125
rect 31289 48091 31323 48123
rect 31289 48021 31323 48053
rect 31289 48019 31323 48021
rect 31289 47953 31323 47981
rect 31289 47947 31323 47953
rect 31289 47885 31323 47909
rect 31289 47875 31323 47885
rect 31289 47817 31323 47837
rect 31289 47803 31323 47817
rect 31289 47749 31323 47765
rect 31289 47731 31323 47749
rect 31289 47681 31323 47693
rect 31289 47659 31323 47681
rect 31289 47613 31323 47621
rect 31289 47587 31323 47613
rect 31289 47545 31323 47549
rect 31289 47515 31323 47545
rect 31289 47443 31323 47477
rect 31747 48667 31781 48701
rect 31747 48599 31781 48629
rect 31747 48595 31781 48599
rect 31747 48531 31781 48557
rect 31747 48523 31781 48531
rect 31747 48463 31781 48485
rect 31747 48451 31781 48463
rect 31747 48395 31781 48413
rect 31747 48379 31781 48395
rect 31747 48327 31781 48341
rect 31747 48307 31781 48327
rect 31747 48259 31781 48269
rect 31747 48235 31781 48259
rect 31747 48191 31781 48197
rect 31747 48163 31781 48191
rect 31747 48123 31781 48125
rect 31747 48091 31781 48123
rect 31747 48021 31781 48053
rect 31747 48019 31781 48021
rect 31747 47953 31781 47981
rect 31747 47947 31781 47953
rect 31747 47885 31781 47909
rect 31747 47875 31781 47885
rect 31747 47817 31781 47837
rect 31747 47803 31781 47817
rect 31747 47749 31781 47765
rect 31747 47731 31781 47749
rect 31747 47681 31781 47693
rect 31747 47659 31781 47681
rect 31747 47613 31781 47621
rect 31747 47587 31781 47613
rect 31747 47545 31781 47549
rect 31747 47515 31781 47545
rect 31747 47443 31781 47477
rect 32205 48667 32239 48701
rect 32205 48599 32239 48629
rect 32205 48595 32239 48599
rect 32205 48531 32239 48557
rect 32205 48523 32239 48531
rect 32205 48463 32239 48485
rect 32205 48451 32239 48463
rect 32205 48395 32239 48413
rect 32205 48379 32239 48395
rect 32205 48327 32239 48341
rect 32205 48307 32239 48327
rect 32205 48259 32239 48269
rect 32205 48235 32239 48259
rect 32205 48191 32239 48197
rect 32205 48163 32239 48191
rect 32205 48123 32239 48125
rect 32205 48091 32239 48123
rect 32205 48021 32239 48053
rect 32205 48019 32239 48021
rect 32205 47953 32239 47981
rect 32205 47947 32239 47953
rect 32205 47885 32239 47909
rect 32205 47875 32239 47885
rect 32205 47817 32239 47837
rect 32205 47803 32239 47817
rect 32205 47749 32239 47765
rect 32205 47731 32239 47749
rect 32205 47681 32239 47693
rect 32205 47659 32239 47681
rect 32205 47613 32239 47621
rect 32205 47587 32239 47613
rect 32205 47545 32239 47549
rect 32205 47515 32239 47545
rect 32205 47443 32239 47477
rect 32663 48667 32697 48701
rect 32663 48599 32697 48629
rect 32663 48595 32697 48599
rect 32663 48531 32697 48557
rect 32663 48523 32697 48531
rect 32663 48463 32697 48485
rect 32663 48451 32697 48463
rect 32663 48395 32697 48413
rect 32663 48379 32697 48395
rect 32663 48327 32697 48341
rect 32663 48307 32697 48327
rect 32663 48259 32697 48269
rect 32663 48235 32697 48259
rect 32663 48191 32697 48197
rect 32663 48163 32697 48191
rect 32663 48123 32697 48125
rect 32663 48091 32697 48123
rect 32663 48021 32697 48053
rect 32663 48019 32697 48021
rect 32663 47953 32697 47981
rect 32663 47947 32697 47953
rect 32663 47885 32697 47909
rect 32663 47875 32697 47885
rect 32663 47817 32697 47837
rect 32663 47803 32697 47817
rect 32663 47749 32697 47765
rect 32663 47731 32697 47749
rect 32663 47681 32697 47693
rect 32663 47659 32697 47681
rect 32663 47613 32697 47621
rect 32663 47587 32697 47613
rect 32663 47545 32697 47549
rect 32663 47515 32697 47545
rect 32663 47443 32697 47477
rect 33121 48667 33155 48701
rect 33121 48599 33155 48629
rect 33121 48595 33155 48599
rect 33121 48531 33155 48557
rect 33121 48523 33155 48531
rect 33121 48463 33155 48485
rect 33121 48451 33155 48463
rect 33121 48395 33155 48413
rect 33121 48379 33155 48395
rect 33121 48327 33155 48341
rect 33121 48307 33155 48327
rect 33121 48259 33155 48269
rect 33121 48235 33155 48259
rect 33121 48191 33155 48197
rect 33121 48163 33155 48191
rect 33121 48123 33155 48125
rect 33121 48091 33155 48123
rect 33121 48021 33155 48053
rect 33121 48019 33155 48021
rect 33121 47953 33155 47981
rect 33121 47947 33155 47953
rect 33121 47885 33155 47909
rect 33121 47875 33155 47885
rect 33121 47817 33155 47837
rect 33121 47803 33155 47817
rect 33121 47749 33155 47765
rect 33121 47731 33155 47749
rect 33121 47681 33155 47693
rect 33121 47659 33155 47681
rect 33121 47613 33155 47621
rect 33121 47587 33155 47613
rect 33121 47545 33155 47549
rect 33121 47515 33155 47545
rect 33121 47443 33155 47477
rect 33579 48667 33613 48701
rect 33579 48599 33613 48629
rect 33579 48595 33613 48599
rect 33579 48531 33613 48557
rect 33579 48523 33613 48531
rect 33579 48463 33613 48485
rect 33579 48451 33613 48463
rect 33579 48395 33613 48413
rect 33579 48379 33613 48395
rect 33579 48327 33613 48341
rect 33579 48307 33613 48327
rect 33579 48259 33613 48269
rect 33579 48235 33613 48259
rect 33579 48191 33613 48197
rect 33579 48163 33613 48191
rect 33579 48123 33613 48125
rect 33579 48091 33613 48123
rect 33579 48021 33613 48053
rect 33579 48019 33613 48021
rect 33579 47953 33613 47981
rect 33579 47947 33613 47953
rect 33579 47885 33613 47909
rect 33579 47875 33613 47885
rect 33579 47817 33613 47837
rect 33579 47803 33613 47817
rect 33579 47749 33613 47765
rect 33579 47731 33613 47749
rect 33579 47681 33613 47693
rect 33579 47659 33613 47681
rect 33579 47613 33613 47621
rect 33579 47587 33613 47613
rect 33579 47545 33613 47549
rect 33579 47515 33613 47545
rect 33579 47443 33613 47477
rect 34037 48667 34071 48701
rect 34037 48599 34071 48629
rect 34037 48595 34071 48599
rect 34037 48531 34071 48557
rect 34037 48523 34071 48531
rect 34037 48463 34071 48485
rect 34037 48451 34071 48463
rect 34037 48395 34071 48413
rect 34037 48379 34071 48395
rect 34037 48327 34071 48341
rect 34037 48307 34071 48327
rect 34037 48259 34071 48269
rect 34037 48235 34071 48259
rect 34037 48191 34071 48197
rect 34037 48163 34071 48191
rect 34037 48123 34071 48125
rect 34037 48091 34071 48123
rect 34037 48021 34071 48053
rect 34037 48019 34071 48021
rect 34037 47953 34071 47981
rect 34037 47947 34071 47953
rect 34037 47885 34071 47909
rect 34037 47875 34071 47885
rect 34037 47817 34071 47837
rect 34037 47803 34071 47817
rect 34037 47749 34071 47765
rect 34037 47731 34071 47749
rect 34037 47681 34071 47693
rect 34037 47659 34071 47681
rect 34037 47613 34071 47621
rect 34037 47587 34071 47613
rect 34037 47545 34071 47549
rect 34037 47515 34071 47545
rect 34037 47443 34071 47477
rect 34495 48667 34529 48701
rect 34495 48599 34529 48629
rect 34495 48595 34529 48599
rect 34495 48531 34529 48557
rect 34495 48523 34529 48531
rect 34495 48463 34529 48485
rect 34495 48451 34529 48463
rect 34495 48395 34529 48413
rect 34495 48379 34529 48395
rect 34495 48327 34529 48341
rect 34495 48307 34529 48327
rect 34495 48259 34529 48269
rect 34495 48235 34529 48259
rect 34495 48191 34529 48197
rect 34495 48163 34529 48191
rect 34495 48123 34529 48125
rect 34495 48091 34529 48123
rect 34495 48021 34529 48053
rect 34495 48019 34529 48021
rect 34495 47953 34529 47981
rect 34495 47947 34529 47953
rect 34495 47885 34529 47909
rect 34495 47875 34529 47885
rect 34495 47817 34529 47837
rect 34495 47803 34529 47817
rect 34495 47749 34529 47765
rect 34495 47731 34529 47749
rect 34495 47681 34529 47693
rect 34495 47659 34529 47681
rect 34495 47613 34529 47621
rect 34495 47587 34529 47613
rect 34495 47545 34529 47549
rect 34495 47515 34529 47545
rect 34495 47443 34529 47477
rect 34953 48667 34987 48701
rect 34953 48599 34987 48629
rect 34953 48595 34987 48599
rect 34953 48531 34987 48557
rect 34953 48523 34987 48531
rect 34953 48463 34987 48485
rect 34953 48451 34987 48463
rect 34953 48395 34987 48413
rect 34953 48379 34987 48395
rect 34953 48327 34987 48341
rect 34953 48307 34987 48327
rect 34953 48259 34987 48269
rect 34953 48235 34987 48259
rect 34953 48191 34987 48197
rect 34953 48163 34987 48191
rect 34953 48123 34987 48125
rect 34953 48091 34987 48123
rect 34953 48021 34987 48053
rect 34953 48019 34987 48021
rect 34953 47953 34987 47981
rect 34953 47947 34987 47953
rect 34953 47885 34987 47909
rect 34953 47875 34987 47885
rect 34953 47817 34987 47837
rect 34953 47803 34987 47817
rect 34953 47749 34987 47765
rect 34953 47731 34987 47749
rect 34953 47681 34987 47693
rect 34953 47659 34987 47681
rect 34953 47613 34987 47621
rect 34953 47587 34987 47613
rect 34953 47545 34987 47549
rect 34953 47515 34987 47545
rect 34953 47443 34987 47477
rect 35411 48667 35445 48701
rect 35411 48599 35445 48629
rect 35411 48595 35445 48599
rect 35411 48531 35445 48557
rect 35411 48523 35445 48531
rect 35411 48463 35445 48485
rect 35411 48451 35445 48463
rect 35411 48395 35445 48413
rect 35411 48379 35445 48395
rect 35411 48327 35445 48341
rect 35411 48307 35445 48327
rect 35411 48259 35445 48269
rect 35411 48235 35445 48259
rect 35411 48191 35445 48197
rect 35411 48163 35445 48191
rect 35411 48123 35445 48125
rect 35411 48091 35445 48123
rect 35411 48021 35445 48053
rect 35411 48019 35445 48021
rect 35411 47953 35445 47981
rect 35411 47947 35445 47953
rect 35411 47885 35445 47909
rect 35411 47875 35445 47885
rect 35411 47817 35445 47837
rect 35411 47803 35445 47817
rect 35411 47749 35445 47765
rect 35411 47731 35445 47749
rect 35411 47681 35445 47693
rect 35411 47659 35445 47681
rect 35411 47613 35445 47621
rect 35411 47587 35445 47613
rect 35411 47545 35445 47549
rect 35411 47515 35445 47545
rect 35411 47443 35445 47477
rect 35869 48667 35903 48701
rect 35869 48599 35903 48629
rect 35869 48595 35903 48599
rect 35869 48531 35903 48557
rect 35869 48523 35903 48531
rect 35869 48463 35903 48485
rect 35869 48451 35903 48463
rect 35869 48395 35903 48413
rect 35869 48379 35903 48395
rect 35869 48327 35903 48341
rect 35869 48307 35903 48327
rect 35869 48259 35903 48269
rect 35869 48235 35903 48259
rect 35869 48191 35903 48197
rect 35869 48163 35903 48191
rect 35869 48123 35903 48125
rect 35869 48091 35903 48123
rect 35869 48021 35903 48053
rect 35869 48019 35903 48021
rect 35869 47953 35903 47981
rect 35869 47947 35903 47953
rect 35869 47885 35903 47909
rect 35869 47875 35903 47885
rect 35869 47817 35903 47837
rect 35869 47803 35903 47817
rect 35869 47749 35903 47765
rect 35869 47731 35903 47749
rect 35869 47681 35903 47693
rect 35869 47659 35903 47681
rect 35869 47613 35903 47621
rect 35869 47587 35903 47613
rect 35869 47545 35903 47549
rect 35869 47515 35903 47545
rect 35869 47443 35903 47477
rect 36327 48667 36361 48701
rect 36327 48599 36361 48629
rect 36327 48595 36361 48599
rect 36327 48531 36361 48557
rect 36327 48523 36361 48531
rect 36327 48463 36361 48485
rect 36327 48451 36361 48463
rect 36327 48395 36361 48413
rect 36327 48379 36361 48395
rect 36327 48327 36361 48341
rect 36327 48307 36361 48327
rect 36327 48259 36361 48269
rect 36327 48235 36361 48259
rect 36327 48191 36361 48197
rect 36327 48163 36361 48191
rect 36327 48123 36361 48125
rect 36327 48091 36361 48123
rect 36327 48021 36361 48053
rect 36327 48019 36361 48021
rect 36327 47953 36361 47981
rect 36327 47947 36361 47953
rect 36327 47885 36361 47909
rect 36327 47875 36361 47885
rect 36327 47817 36361 47837
rect 36327 47803 36361 47817
rect 36327 47749 36361 47765
rect 36327 47731 36361 47749
rect 36327 47681 36361 47693
rect 36327 47659 36361 47681
rect 36327 47613 36361 47621
rect 36327 47587 36361 47613
rect 36327 47545 36361 47549
rect 36327 47515 36361 47545
rect 36327 47443 36361 47477
rect 36785 48667 36819 48701
rect 36785 48599 36819 48629
rect 36785 48595 36819 48599
rect 36785 48531 36819 48557
rect 36785 48523 36819 48531
rect 36785 48463 36819 48485
rect 36785 48451 36819 48463
rect 36785 48395 36819 48413
rect 36785 48379 36819 48395
rect 36785 48327 36819 48341
rect 36785 48307 36819 48327
rect 36785 48259 36819 48269
rect 36785 48235 36819 48259
rect 36785 48191 36819 48197
rect 36785 48163 36819 48191
rect 36785 48123 36819 48125
rect 36785 48091 36819 48123
rect 36785 48021 36819 48053
rect 36785 48019 36819 48021
rect 36785 47953 36819 47981
rect 36785 47947 36819 47953
rect 36785 47885 36819 47909
rect 36785 47875 36819 47885
rect 36785 47817 36819 47837
rect 36785 47803 36819 47817
rect 36785 47749 36819 47765
rect 36785 47731 36819 47749
rect 36785 47681 36819 47693
rect 36785 47659 36819 47681
rect 36785 47613 36819 47621
rect 36785 47587 36819 47613
rect 36785 47545 36819 47549
rect 36785 47515 36819 47545
rect 36785 47443 36819 47477
rect 37243 48667 37277 48701
rect 37243 48599 37277 48629
rect 37243 48595 37277 48599
rect 37243 48531 37277 48557
rect 37243 48523 37277 48531
rect 37243 48463 37277 48485
rect 37243 48451 37277 48463
rect 37243 48395 37277 48413
rect 37243 48379 37277 48395
rect 37243 48327 37277 48341
rect 37243 48307 37277 48327
rect 37243 48259 37277 48269
rect 37243 48235 37277 48259
rect 37243 48191 37277 48197
rect 37243 48163 37277 48191
rect 37243 48123 37277 48125
rect 37243 48091 37277 48123
rect 37243 48021 37277 48053
rect 37243 48019 37277 48021
rect 37243 47953 37277 47981
rect 37243 47947 37277 47953
rect 37243 47885 37277 47909
rect 37243 47875 37277 47885
rect 37243 47817 37277 47837
rect 37243 47803 37277 47817
rect 37243 47749 37277 47765
rect 37243 47731 37277 47749
rect 37243 47681 37277 47693
rect 37243 47659 37277 47681
rect 37243 47613 37277 47621
rect 37243 47587 37277 47613
rect 37243 47545 37277 47549
rect 37243 47515 37277 47545
rect 37243 47443 37277 47477
rect 37701 48667 37735 48701
rect 37701 48599 37735 48629
rect 37701 48595 37735 48599
rect 37701 48531 37735 48557
rect 37701 48523 37735 48531
rect 37701 48463 37735 48485
rect 37701 48451 37735 48463
rect 37701 48395 37735 48413
rect 37701 48379 37735 48395
rect 37701 48327 37735 48341
rect 37701 48307 37735 48327
rect 37701 48259 37735 48269
rect 37701 48235 37735 48259
rect 37701 48191 37735 48197
rect 37701 48163 37735 48191
rect 37701 48123 37735 48125
rect 37701 48091 37735 48123
rect 37701 48021 37735 48053
rect 37701 48019 37735 48021
rect 37701 47953 37735 47981
rect 37701 47947 37735 47953
rect 37701 47885 37735 47909
rect 37701 47875 37735 47885
rect 37701 47817 37735 47837
rect 37701 47803 37735 47817
rect 37701 47749 37735 47765
rect 37701 47731 37735 47749
rect 37701 47681 37735 47693
rect 37701 47659 37735 47681
rect 37701 47613 37735 47621
rect 37701 47587 37735 47613
rect 37701 47545 37735 47549
rect 37701 47515 37735 47545
rect 37701 47443 37735 47477
rect 38159 48667 38193 48701
rect 38159 48599 38193 48629
rect 38159 48595 38193 48599
rect 38159 48531 38193 48557
rect 38159 48523 38193 48531
rect 38159 48463 38193 48485
rect 38159 48451 38193 48463
rect 38159 48395 38193 48413
rect 38159 48379 38193 48395
rect 38159 48327 38193 48341
rect 38159 48307 38193 48327
rect 38159 48259 38193 48269
rect 38159 48235 38193 48259
rect 38159 48191 38193 48197
rect 38159 48163 38193 48191
rect 38159 48123 38193 48125
rect 38159 48091 38193 48123
rect 38159 48021 38193 48053
rect 38159 48019 38193 48021
rect 38159 47953 38193 47981
rect 38159 47947 38193 47953
rect 38159 47885 38193 47909
rect 38159 47875 38193 47885
rect 38159 47817 38193 47837
rect 38159 47803 38193 47817
rect 38159 47749 38193 47765
rect 38159 47731 38193 47749
rect 38159 47681 38193 47693
rect 38159 47659 38193 47681
rect 38159 47613 38193 47621
rect 38159 47587 38193 47613
rect 38159 47545 38193 47549
rect 38159 47515 38193 47545
rect 38159 47443 38193 47477
rect 38617 48667 38651 48701
rect 38617 48599 38651 48629
rect 38617 48595 38651 48599
rect 38617 48531 38651 48557
rect 38617 48523 38651 48531
rect 38617 48463 38651 48485
rect 38617 48451 38651 48463
rect 38617 48395 38651 48413
rect 38617 48379 38651 48395
rect 38617 48327 38651 48341
rect 38617 48307 38651 48327
rect 38617 48259 38651 48269
rect 38617 48235 38651 48259
rect 38617 48191 38651 48197
rect 38617 48163 38651 48191
rect 38617 48123 38651 48125
rect 38617 48091 38651 48123
rect 38617 48021 38651 48053
rect 38617 48019 38651 48021
rect 38617 47953 38651 47981
rect 38617 47947 38651 47953
rect 38617 47885 38651 47909
rect 38617 47875 38651 47885
rect 38617 47817 38651 47837
rect 38617 47803 38651 47817
rect 38617 47749 38651 47765
rect 38617 47731 38651 47749
rect 38617 47681 38651 47693
rect 38617 47659 38651 47681
rect 38617 47613 38651 47621
rect 38617 47587 38651 47613
rect 38617 47545 38651 47549
rect 38617 47515 38651 47545
rect 38617 47443 38651 47477
rect 39075 48667 39109 48701
rect 39075 48599 39109 48629
rect 39075 48595 39109 48599
rect 39075 48531 39109 48557
rect 39075 48523 39109 48531
rect 39075 48463 39109 48485
rect 39075 48451 39109 48463
rect 39075 48395 39109 48413
rect 39075 48379 39109 48395
rect 39075 48327 39109 48341
rect 39075 48307 39109 48327
rect 39075 48259 39109 48269
rect 39075 48235 39109 48259
rect 39075 48191 39109 48197
rect 39075 48163 39109 48191
rect 39075 48123 39109 48125
rect 39075 48091 39109 48123
rect 39075 48021 39109 48053
rect 39075 48019 39109 48021
rect 39075 47953 39109 47981
rect 39075 47947 39109 47953
rect 39075 47885 39109 47909
rect 39075 47875 39109 47885
rect 39075 47817 39109 47837
rect 39075 47803 39109 47817
rect 39075 47749 39109 47765
rect 39075 47731 39109 47749
rect 39075 47681 39109 47693
rect 39075 47659 39109 47681
rect 39075 47613 39109 47621
rect 39075 47587 39109 47613
rect 39075 47545 39109 47549
rect 39075 47515 39109 47545
rect 39075 47443 39109 47477
rect 39533 48667 39567 48701
rect 39533 48599 39567 48629
rect 39533 48595 39567 48599
rect 39533 48531 39567 48557
rect 39533 48523 39567 48531
rect 39533 48463 39567 48485
rect 39533 48451 39567 48463
rect 39533 48395 39567 48413
rect 39533 48379 39567 48395
rect 39533 48327 39567 48341
rect 39533 48307 39567 48327
rect 39533 48259 39567 48269
rect 39533 48235 39567 48259
rect 39533 48191 39567 48197
rect 39533 48163 39567 48191
rect 39533 48123 39567 48125
rect 39533 48091 39567 48123
rect 39533 48021 39567 48053
rect 39533 48019 39567 48021
rect 39533 47953 39567 47981
rect 39533 47947 39567 47953
rect 39533 47885 39567 47909
rect 39533 47875 39567 47885
rect 39533 47817 39567 47837
rect 39533 47803 39567 47817
rect 39533 47749 39567 47765
rect 39533 47731 39567 47749
rect 39533 47681 39567 47693
rect 39533 47659 39567 47681
rect 39533 47613 39567 47621
rect 39533 47587 39567 47613
rect 39533 47545 39567 47549
rect 39533 47515 39567 47545
rect 39533 47443 39567 47477
rect 39991 48667 40025 48701
rect 39991 48599 40025 48629
rect 39991 48595 40025 48599
rect 39991 48531 40025 48557
rect 39991 48523 40025 48531
rect 39991 48463 40025 48485
rect 39991 48451 40025 48463
rect 39991 48395 40025 48413
rect 39991 48379 40025 48395
rect 39991 48327 40025 48341
rect 39991 48307 40025 48327
rect 39991 48259 40025 48269
rect 39991 48235 40025 48259
rect 39991 48191 40025 48197
rect 39991 48163 40025 48191
rect 39991 48123 40025 48125
rect 39991 48091 40025 48123
rect 39991 48021 40025 48053
rect 39991 48019 40025 48021
rect 39991 47953 40025 47981
rect 39991 47947 40025 47953
rect 39991 47885 40025 47909
rect 39991 47875 40025 47885
rect 39991 47817 40025 47837
rect 39991 47803 40025 47817
rect 39991 47749 40025 47765
rect 39991 47731 40025 47749
rect 39991 47681 40025 47693
rect 39991 47659 40025 47681
rect 39991 47613 40025 47621
rect 39991 47587 40025 47613
rect 39991 47545 40025 47549
rect 39991 47515 40025 47545
rect 39991 47443 40025 47477
rect 40449 48667 40483 48701
rect 40449 48599 40483 48629
rect 40449 48595 40483 48599
rect 40449 48531 40483 48557
rect 40449 48523 40483 48531
rect 40449 48463 40483 48485
rect 40449 48451 40483 48463
rect 40449 48395 40483 48413
rect 40449 48379 40483 48395
rect 40449 48327 40483 48341
rect 40449 48307 40483 48327
rect 40449 48259 40483 48269
rect 40449 48235 40483 48259
rect 40449 48191 40483 48197
rect 40449 48163 40483 48191
rect 40449 48123 40483 48125
rect 40449 48091 40483 48123
rect 40449 48021 40483 48053
rect 40449 48019 40483 48021
rect 40449 47953 40483 47981
rect 40449 47947 40483 47953
rect 40449 47885 40483 47909
rect 40449 47875 40483 47885
rect 40449 47817 40483 47837
rect 40449 47803 40483 47817
rect 40449 47749 40483 47765
rect 40449 47731 40483 47749
rect 40449 47681 40483 47693
rect 40449 47659 40483 47681
rect 40449 47613 40483 47621
rect 40449 47587 40483 47613
rect 40449 47545 40483 47549
rect 40449 47515 40483 47545
rect 40449 47443 40483 47477
rect 40907 48667 40941 48701
rect 40907 48599 40941 48629
rect 40907 48595 40941 48599
rect 40907 48531 40941 48557
rect 40907 48523 40941 48531
rect 40907 48463 40941 48485
rect 40907 48451 40941 48463
rect 40907 48395 40941 48413
rect 40907 48379 40941 48395
rect 40907 48327 40941 48341
rect 40907 48307 40941 48327
rect 40907 48259 40941 48269
rect 40907 48235 40941 48259
rect 40907 48191 40941 48197
rect 40907 48163 40941 48191
rect 40907 48123 40941 48125
rect 40907 48091 40941 48123
rect 40907 48021 40941 48053
rect 40907 48019 40941 48021
rect 40907 47953 40941 47981
rect 40907 47947 40941 47953
rect 40907 47885 40941 47909
rect 40907 47875 40941 47885
rect 40907 47817 40941 47837
rect 40907 47803 40941 47817
rect 40907 47749 40941 47765
rect 40907 47731 40941 47749
rect 40907 47681 40941 47693
rect 40907 47659 40941 47681
rect 40907 47613 40941 47621
rect 40907 47587 40941 47613
rect 40907 47545 40941 47549
rect 40907 47515 40941 47545
rect 40907 47443 40941 47477
rect 41365 48667 41399 48701
rect 41365 48599 41399 48629
rect 41365 48595 41399 48599
rect 41365 48531 41399 48557
rect 41365 48523 41399 48531
rect 41365 48463 41399 48485
rect 41365 48451 41399 48463
rect 41365 48395 41399 48413
rect 41365 48379 41399 48395
rect 41365 48327 41399 48341
rect 41365 48307 41399 48327
rect 41365 48259 41399 48269
rect 41365 48235 41399 48259
rect 41365 48191 41399 48197
rect 41365 48163 41399 48191
rect 41365 48123 41399 48125
rect 41365 48091 41399 48123
rect 41365 48021 41399 48053
rect 41365 48019 41399 48021
rect 41365 47953 41399 47981
rect 41365 47947 41399 47953
rect 41365 47885 41399 47909
rect 41365 47875 41399 47885
rect 41365 47817 41399 47837
rect 41365 47803 41399 47817
rect 41365 47749 41399 47765
rect 41365 47731 41399 47749
rect 41365 47681 41399 47693
rect 41365 47659 41399 47681
rect 41365 47613 41399 47621
rect 41365 47587 41399 47613
rect 41365 47545 41399 47549
rect 41365 47515 41399 47545
rect 41365 47443 41399 47477
rect 41823 48667 41857 48701
rect 41823 48599 41857 48629
rect 41823 48595 41857 48599
rect 41823 48531 41857 48557
rect 41823 48523 41857 48531
rect 41823 48463 41857 48485
rect 41823 48451 41857 48463
rect 41823 48395 41857 48413
rect 41823 48379 41857 48395
rect 41823 48327 41857 48341
rect 41823 48307 41857 48327
rect 41823 48259 41857 48269
rect 41823 48235 41857 48259
rect 41823 48191 41857 48197
rect 41823 48163 41857 48191
rect 41823 48123 41857 48125
rect 41823 48091 41857 48123
rect 41823 48021 41857 48053
rect 41823 48019 41857 48021
rect 41823 47953 41857 47981
rect 41823 47947 41857 47953
rect 41823 47885 41857 47909
rect 41823 47875 41857 47885
rect 41823 47817 41857 47837
rect 41823 47803 41857 47817
rect 41823 47749 41857 47765
rect 41823 47731 41857 47749
rect 41823 47681 41857 47693
rect 41823 47659 41857 47681
rect 41823 47613 41857 47621
rect 41823 47587 41857 47613
rect 41823 47545 41857 47549
rect 41823 47515 41857 47545
rect 41823 47443 41857 47477
rect 42281 48667 42315 48701
rect 42281 48599 42315 48629
rect 42281 48595 42315 48599
rect 42281 48531 42315 48557
rect 42281 48523 42315 48531
rect 42281 48463 42315 48485
rect 42281 48451 42315 48463
rect 42281 48395 42315 48413
rect 42281 48379 42315 48395
rect 42281 48327 42315 48341
rect 42281 48307 42315 48327
rect 42281 48259 42315 48269
rect 42281 48235 42315 48259
rect 42281 48191 42315 48197
rect 42281 48163 42315 48191
rect 42281 48123 42315 48125
rect 42281 48091 42315 48123
rect 42281 48021 42315 48053
rect 42281 48019 42315 48021
rect 42281 47953 42315 47981
rect 42281 47947 42315 47953
rect 42281 47885 42315 47909
rect 42281 47875 42315 47885
rect 42281 47817 42315 47837
rect 42281 47803 42315 47817
rect 42281 47749 42315 47765
rect 42281 47731 42315 47749
rect 42281 47681 42315 47693
rect 42281 47659 42315 47681
rect 42281 47613 42315 47621
rect 42281 47587 42315 47613
rect 42281 47545 42315 47549
rect 42281 47515 42315 47545
rect 42281 47443 42315 47477
rect 42739 48667 42773 48701
rect 42739 48599 42773 48629
rect 42739 48595 42773 48599
rect 42739 48531 42773 48557
rect 42739 48523 42773 48531
rect 42739 48463 42773 48485
rect 42739 48451 42773 48463
rect 42739 48395 42773 48413
rect 42739 48379 42773 48395
rect 42739 48327 42773 48341
rect 42739 48307 42773 48327
rect 42739 48259 42773 48269
rect 42739 48235 42773 48259
rect 42739 48191 42773 48197
rect 42739 48163 42773 48191
rect 42739 48123 42773 48125
rect 42739 48091 42773 48123
rect 42739 48021 42773 48053
rect 42739 48019 42773 48021
rect 42739 47953 42773 47981
rect 42739 47947 42773 47953
rect 42739 47885 42773 47909
rect 42739 47875 42773 47885
rect 42739 47817 42773 47837
rect 42739 47803 42773 47817
rect 42739 47749 42773 47765
rect 42739 47731 42773 47749
rect 42739 47681 42773 47693
rect 42739 47659 42773 47681
rect 42739 47613 42773 47621
rect 42739 47587 42773 47613
rect 42739 47545 42773 47549
rect 42739 47515 42773 47545
rect 42739 47443 42773 47477
rect 43197 48667 43231 48701
rect 43197 48599 43231 48629
rect 43197 48595 43231 48599
rect 43197 48531 43231 48557
rect 43197 48523 43231 48531
rect 43197 48463 43231 48485
rect 43197 48451 43231 48463
rect 43197 48395 43231 48413
rect 43197 48379 43231 48395
rect 43197 48327 43231 48341
rect 43197 48307 43231 48327
rect 43197 48259 43231 48269
rect 43197 48235 43231 48259
rect 43197 48191 43231 48197
rect 43197 48163 43231 48191
rect 43197 48123 43231 48125
rect 43197 48091 43231 48123
rect 43197 48021 43231 48053
rect 43197 48019 43231 48021
rect 43197 47953 43231 47981
rect 43197 47947 43231 47953
rect 43197 47885 43231 47909
rect 43197 47875 43231 47885
rect 43197 47817 43231 47837
rect 43197 47803 43231 47817
rect 43197 47749 43231 47765
rect 43197 47731 43231 47749
rect 43197 47681 43231 47693
rect 43197 47659 43231 47681
rect 43197 47613 43231 47621
rect 43197 47587 43231 47613
rect 43197 47545 43231 47549
rect 43197 47515 43231 47545
rect 43197 47443 43231 47477
rect 43655 48667 43689 48701
rect 43655 48599 43689 48629
rect 43655 48595 43689 48599
rect 43655 48531 43689 48557
rect 43655 48523 43689 48531
rect 43655 48463 43689 48485
rect 43655 48451 43689 48463
rect 43655 48395 43689 48413
rect 43655 48379 43689 48395
rect 43655 48327 43689 48341
rect 43655 48307 43689 48327
rect 43655 48259 43689 48269
rect 43655 48235 43689 48259
rect 43655 48191 43689 48197
rect 43655 48163 43689 48191
rect 43655 48123 43689 48125
rect 43655 48091 43689 48123
rect 43655 48021 43689 48053
rect 43655 48019 43689 48021
rect 43655 47953 43689 47981
rect 43655 47947 43689 47953
rect 43655 47885 43689 47909
rect 43655 47875 43689 47885
rect 43655 47817 43689 47837
rect 43655 47803 43689 47817
rect 43655 47749 43689 47765
rect 43655 47731 43689 47749
rect 43655 47681 43689 47693
rect 43655 47659 43689 47681
rect 43655 47613 43689 47621
rect 43655 47587 43689 47613
rect 43655 47545 43689 47549
rect 43655 47515 43689 47545
rect 43655 47443 43689 47477
rect 44113 48667 44147 48701
rect 44113 48599 44147 48629
rect 44113 48595 44147 48599
rect 44113 48531 44147 48557
rect 44113 48523 44147 48531
rect 44113 48463 44147 48485
rect 44113 48451 44147 48463
rect 44113 48395 44147 48413
rect 44113 48379 44147 48395
rect 44113 48327 44147 48341
rect 44113 48307 44147 48327
rect 44113 48259 44147 48269
rect 44113 48235 44147 48259
rect 44113 48191 44147 48197
rect 44113 48163 44147 48191
rect 44113 48123 44147 48125
rect 44113 48091 44147 48123
rect 44113 48021 44147 48053
rect 44113 48019 44147 48021
rect 44113 47953 44147 47981
rect 44113 47947 44147 47953
rect 44113 47885 44147 47909
rect 44113 47875 44147 47885
rect 44113 47817 44147 47837
rect 44113 47803 44147 47817
rect 44113 47749 44147 47765
rect 44113 47731 44147 47749
rect 44113 47681 44147 47693
rect 44113 47659 44147 47681
rect 44113 47613 44147 47621
rect 44113 47587 44147 47613
rect 44113 47545 44147 47549
rect 44113 47515 44147 47545
rect 44113 47443 44147 47477
rect 44571 48667 44605 48701
rect 44571 48599 44605 48629
rect 44571 48595 44605 48599
rect 44571 48531 44605 48557
rect 44571 48523 44605 48531
rect 44571 48463 44605 48485
rect 44571 48451 44605 48463
rect 44571 48395 44605 48413
rect 44571 48379 44605 48395
rect 44571 48327 44605 48341
rect 44571 48307 44605 48327
rect 44571 48259 44605 48269
rect 44571 48235 44605 48259
rect 44571 48191 44605 48197
rect 44571 48163 44605 48191
rect 44571 48123 44605 48125
rect 44571 48091 44605 48123
rect 44571 48021 44605 48053
rect 44571 48019 44605 48021
rect 44571 47953 44605 47981
rect 44571 47947 44605 47953
rect 44571 47885 44605 47909
rect 44571 47875 44605 47885
rect 44571 47817 44605 47837
rect 44571 47803 44605 47817
rect 44571 47749 44605 47765
rect 44571 47731 44605 47749
rect 44571 47681 44605 47693
rect 44571 47659 44605 47681
rect 44571 47613 44605 47621
rect 44571 47587 44605 47613
rect 44571 47545 44605 47549
rect 44571 47515 44605 47545
rect 44571 47443 44605 47477
rect 45029 48667 45063 48701
rect 45029 48599 45063 48629
rect 45029 48595 45063 48599
rect 45029 48531 45063 48557
rect 45029 48523 45063 48531
rect 45029 48463 45063 48485
rect 45029 48451 45063 48463
rect 45029 48395 45063 48413
rect 45029 48379 45063 48395
rect 45029 48327 45063 48341
rect 45029 48307 45063 48327
rect 45029 48259 45063 48269
rect 45029 48235 45063 48259
rect 45029 48191 45063 48197
rect 45029 48163 45063 48191
rect 45029 48123 45063 48125
rect 45029 48091 45063 48123
rect 45029 48021 45063 48053
rect 45029 48019 45063 48021
rect 45029 47953 45063 47981
rect 45029 47947 45063 47953
rect 45029 47885 45063 47909
rect 45029 47875 45063 47885
rect 45029 47817 45063 47837
rect 45029 47803 45063 47817
rect 45029 47749 45063 47765
rect 45029 47731 45063 47749
rect 45029 47681 45063 47693
rect 45029 47659 45063 47681
rect 45029 47613 45063 47621
rect 45029 47587 45063 47613
rect 45029 47545 45063 47549
rect 45029 47515 45063 47545
rect 45029 47443 45063 47477
rect 45487 48667 45521 48701
rect 45487 48599 45521 48629
rect 45487 48595 45521 48599
rect 45487 48531 45521 48557
rect 45487 48523 45521 48531
rect 45487 48463 45521 48485
rect 45487 48451 45521 48463
rect 45487 48395 45521 48413
rect 45487 48379 45521 48395
rect 45487 48327 45521 48341
rect 45487 48307 45521 48327
rect 45487 48259 45521 48269
rect 45487 48235 45521 48259
rect 45487 48191 45521 48197
rect 45487 48163 45521 48191
rect 45487 48123 45521 48125
rect 45487 48091 45521 48123
rect 45487 48021 45521 48053
rect 45487 48019 45521 48021
rect 45487 47953 45521 47981
rect 45487 47947 45521 47953
rect 45487 47885 45521 47909
rect 45487 47875 45521 47885
rect 45487 47817 45521 47837
rect 45487 47803 45521 47817
rect 45487 47749 45521 47765
rect 45487 47731 45521 47749
rect 45487 47681 45521 47693
rect 45487 47659 45521 47681
rect 45487 47613 45521 47621
rect 45487 47587 45521 47613
rect 45487 47545 45521 47549
rect 45487 47515 45521 47545
rect 45487 47443 45521 47477
rect 45945 48667 45979 48701
rect 45945 48599 45979 48629
rect 45945 48595 45979 48599
rect 45945 48531 45979 48557
rect 45945 48523 45979 48531
rect 45945 48463 45979 48485
rect 45945 48451 45979 48463
rect 45945 48395 45979 48413
rect 45945 48379 45979 48395
rect 45945 48327 45979 48341
rect 45945 48307 45979 48327
rect 45945 48259 45979 48269
rect 45945 48235 45979 48259
rect 45945 48191 45979 48197
rect 45945 48163 45979 48191
rect 45945 48123 45979 48125
rect 45945 48091 45979 48123
rect 45945 48021 45979 48053
rect 45945 48019 45979 48021
rect 45945 47953 45979 47981
rect 45945 47947 45979 47953
rect 45945 47885 45979 47909
rect 45945 47875 45979 47885
rect 45945 47817 45979 47837
rect 45945 47803 45979 47817
rect 45945 47749 45979 47765
rect 45945 47731 45979 47749
rect 45945 47681 45979 47693
rect 45945 47659 45979 47681
rect 45945 47613 45979 47621
rect 45945 47587 45979 47613
rect 45945 47545 45979 47549
rect 45945 47515 45979 47545
rect 45945 47443 45979 47477
rect 46403 48667 46437 48701
rect 46403 48599 46437 48629
rect 46403 48595 46437 48599
rect 46403 48531 46437 48557
rect 46403 48523 46437 48531
rect 46403 48463 46437 48485
rect 46403 48451 46437 48463
rect 46403 48395 46437 48413
rect 46403 48379 46437 48395
rect 46403 48327 46437 48341
rect 46403 48307 46437 48327
rect 46403 48259 46437 48269
rect 46403 48235 46437 48259
rect 46403 48191 46437 48197
rect 46403 48163 46437 48191
rect 46403 48123 46437 48125
rect 46403 48091 46437 48123
rect 46403 48021 46437 48053
rect 46403 48019 46437 48021
rect 46403 47953 46437 47981
rect 46403 47947 46437 47953
rect 46403 47885 46437 47909
rect 46403 47875 46437 47885
rect 46403 47817 46437 47837
rect 46403 47803 46437 47817
rect 46403 47749 46437 47765
rect 46403 47731 46437 47749
rect 46403 47681 46437 47693
rect 46403 47659 46437 47681
rect 46403 47613 46437 47621
rect 46403 47587 46437 47613
rect 46403 47545 46437 47549
rect 46403 47515 46437 47545
rect 46403 47443 46437 47477
rect 46861 48667 46895 48701
rect 46861 48599 46895 48629
rect 46861 48595 46895 48599
rect 46861 48531 46895 48557
rect 46861 48523 46895 48531
rect 46861 48463 46895 48485
rect 46861 48451 46895 48463
rect 46861 48395 46895 48413
rect 46861 48379 46895 48395
rect 46861 48327 46895 48341
rect 46861 48307 46895 48327
rect 46861 48259 46895 48269
rect 46861 48235 46895 48259
rect 46861 48191 46895 48197
rect 46861 48163 46895 48191
rect 46861 48123 46895 48125
rect 46861 48091 46895 48123
rect 46861 48021 46895 48053
rect 46861 48019 46895 48021
rect 46861 47953 46895 47981
rect 46861 47947 46895 47953
rect 46861 47885 46895 47909
rect 46861 47875 46895 47885
rect 46861 47817 46895 47837
rect 46861 47803 46895 47817
rect 46861 47749 46895 47765
rect 46861 47731 46895 47749
rect 46861 47681 46895 47693
rect 46861 47659 46895 47681
rect 46861 47613 46895 47621
rect 46861 47587 46895 47613
rect 46861 47545 46895 47549
rect 46861 47515 46895 47545
rect 46861 47443 46895 47477
rect 47319 48667 47353 48701
rect 47319 48599 47353 48629
rect 47319 48595 47353 48599
rect 47319 48531 47353 48557
rect 47319 48523 47353 48531
rect 47319 48463 47353 48485
rect 47319 48451 47353 48463
rect 47319 48395 47353 48413
rect 47319 48379 47353 48395
rect 47319 48327 47353 48341
rect 47319 48307 47353 48327
rect 47319 48259 47353 48269
rect 47319 48235 47353 48259
rect 47319 48191 47353 48197
rect 47319 48163 47353 48191
rect 47319 48123 47353 48125
rect 47319 48091 47353 48123
rect 47319 48021 47353 48053
rect 47319 48019 47353 48021
rect 47319 47953 47353 47981
rect 47319 47947 47353 47953
rect 47319 47885 47353 47909
rect 47319 47875 47353 47885
rect 47319 47817 47353 47837
rect 47319 47803 47353 47817
rect 47319 47749 47353 47765
rect 47319 47731 47353 47749
rect 47319 47681 47353 47693
rect 47319 47659 47353 47681
rect 47319 47613 47353 47621
rect 47319 47587 47353 47613
rect 47319 47545 47353 47549
rect 47319 47515 47353 47545
rect 47319 47443 47353 47477
rect 47777 48667 47811 48701
rect 47777 48599 47811 48629
rect 47777 48595 47811 48599
rect 47777 48531 47811 48557
rect 47777 48523 47811 48531
rect 47777 48463 47811 48485
rect 47777 48451 47811 48463
rect 47777 48395 47811 48413
rect 47777 48379 47811 48395
rect 47777 48327 47811 48341
rect 47777 48307 47811 48327
rect 47777 48259 47811 48269
rect 47777 48235 47811 48259
rect 47777 48191 47811 48197
rect 47777 48163 47811 48191
rect 47777 48123 47811 48125
rect 47777 48091 47811 48123
rect 47777 48021 47811 48053
rect 47777 48019 47811 48021
rect 47777 47953 47811 47981
rect 47777 47947 47811 47953
rect 47777 47885 47811 47909
rect 47777 47875 47811 47885
rect 47777 47817 47811 47837
rect 47777 47803 47811 47817
rect 47777 47749 47811 47765
rect 47777 47731 47811 47749
rect 47777 47681 47811 47693
rect 47777 47659 47811 47681
rect 47777 47613 47811 47621
rect 47777 47587 47811 47613
rect 47777 47545 47811 47549
rect 47777 47515 47811 47545
rect 47777 47443 47811 47477
rect 48235 48667 48269 48701
rect 48235 48599 48269 48629
rect 48235 48595 48269 48599
rect 48235 48531 48269 48557
rect 48235 48523 48269 48531
rect 48235 48463 48269 48485
rect 48235 48451 48269 48463
rect 48235 48395 48269 48413
rect 48235 48379 48269 48395
rect 48235 48327 48269 48341
rect 48235 48307 48269 48327
rect 48235 48259 48269 48269
rect 48235 48235 48269 48259
rect 48235 48191 48269 48197
rect 48235 48163 48269 48191
rect 48235 48123 48269 48125
rect 48235 48091 48269 48123
rect 48235 48021 48269 48053
rect 48235 48019 48269 48021
rect 48235 47953 48269 47981
rect 48235 47947 48269 47953
rect 48235 47885 48269 47909
rect 48235 47875 48269 47885
rect 48235 47817 48269 47837
rect 48235 47803 48269 47817
rect 48235 47749 48269 47765
rect 48235 47731 48269 47749
rect 48235 47681 48269 47693
rect 48235 47659 48269 47681
rect 48235 47613 48269 47621
rect 48235 47587 48269 47613
rect 48235 47545 48269 47549
rect 48235 47515 48269 47545
rect 48235 47443 48269 47477
rect 48693 48667 48727 48701
rect 48693 48599 48727 48629
rect 48693 48595 48727 48599
rect 48693 48531 48727 48557
rect 48693 48523 48727 48531
rect 48693 48463 48727 48485
rect 48693 48451 48727 48463
rect 48693 48395 48727 48413
rect 48693 48379 48727 48395
rect 48693 48327 48727 48341
rect 48693 48307 48727 48327
rect 48693 48259 48727 48269
rect 48693 48235 48727 48259
rect 48693 48191 48727 48197
rect 48693 48163 48727 48191
rect 48693 48123 48727 48125
rect 48693 48091 48727 48123
rect 48693 48021 48727 48053
rect 48693 48019 48727 48021
rect 48693 47953 48727 47981
rect 48693 47947 48727 47953
rect 48693 47885 48727 47909
rect 48693 47875 48727 47885
rect 48693 47817 48727 47837
rect 48693 47803 48727 47817
rect 48693 47749 48727 47765
rect 48693 47731 48727 47749
rect 48693 47681 48727 47693
rect 48693 47659 48727 47681
rect 48693 47613 48727 47621
rect 48693 47587 48727 47613
rect 48693 47545 48727 47549
rect 48693 47515 48727 47545
rect 48693 47443 48727 47477
rect 49151 48667 49185 48701
rect 49151 48599 49185 48629
rect 49151 48595 49185 48599
rect 49151 48531 49185 48557
rect 49151 48523 49185 48531
rect 49151 48463 49185 48485
rect 49151 48451 49185 48463
rect 49151 48395 49185 48413
rect 49151 48379 49185 48395
rect 49151 48327 49185 48341
rect 49151 48307 49185 48327
rect 49151 48259 49185 48269
rect 49151 48235 49185 48259
rect 49151 48191 49185 48197
rect 49151 48163 49185 48191
rect 49151 48123 49185 48125
rect 49151 48091 49185 48123
rect 49151 48021 49185 48053
rect 49151 48019 49185 48021
rect 49151 47953 49185 47981
rect 49151 47947 49185 47953
rect 49151 47885 49185 47909
rect 49151 47875 49185 47885
rect 49151 47817 49185 47837
rect 49151 47803 49185 47817
rect 49151 47749 49185 47765
rect 49151 47731 49185 47749
rect 49151 47681 49185 47693
rect 49151 47659 49185 47681
rect 49151 47613 49185 47621
rect 49151 47587 49185 47613
rect 49151 47545 49185 47549
rect 49151 47515 49185 47545
rect 49151 47443 49185 47477
rect 49609 48667 49643 48701
rect 49609 48599 49643 48629
rect 49609 48595 49643 48599
rect 49609 48531 49643 48557
rect 49609 48523 49643 48531
rect 49609 48463 49643 48485
rect 49609 48451 49643 48463
rect 49609 48395 49643 48413
rect 49609 48379 49643 48395
rect 49609 48327 49643 48341
rect 49609 48307 49643 48327
rect 49609 48259 49643 48269
rect 49609 48235 49643 48259
rect 49609 48191 49643 48197
rect 49609 48163 49643 48191
rect 49609 48123 49643 48125
rect 49609 48091 49643 48123
rect 49609 48021 49643 48053
rect 49609 48019 49643 48021
rect 49609 47953 49643 47981
rect 49609 47947 49643 47953
rect 49609 47885 49643 47909
rect 49609 47875 49643 47885
rect 49609 47817 49643 47837
rect 49609 47803 49643 47817
rect 49609 47749 49643 47765
rect 49609 47731 49643 47749
rect 49609 47681 49643 47693
rect 49609 47659 49643 47681
rect 49609 47613 49643 47621
rect 49609 47587 49643 47613
rect 49609 47545 49643 47549
rect 49609 47515 49643 47545
rect 49609 47443 49643 47477
rect 50067 48667 50101 48701
rect 50067 48599 50101 48629
rect 50067 48595 50101 48599
rect 50067 48531 50101 48557
rect 50067 48523 50101 48531
rect 50067 48463 50101 48485
rect 50067 48451 50101 48463
rect 50067 48395 50101 48413
rect 50067 48379 50101 48395
rect 50067 48327 50101 48341
rect 50067 48307 50101 48327
rect 50067 48259 50101 48269
rect 50067 48235 50101 48259
rect 50067 48191 50101 48197
rect 50067 48163 50101 48191
rect 50067 48123 50101 48125
rect 50067 48091 50101 48123
rect 50067 48021 50101 48053
rect 50067 48019 50101 48021
rect 50067 47953 50101 47981
rect 50067 47947 50101 47953
rect 50067 47885 50101 47909
rect 50067 47875 50101 47885
rect 50067 47817 50101 47837
rect 50067 47803 50101 47817
rect 50067 47749 50101 47765
rect 50067 47731 50101 47749
rect 50067 47681 50101 47693
rect 50067 47659 50101 47681
rect 50067 47613 50101 47621
rect 50067 47587 50101 47613
rect 50067 47545 50101 47549
rect 50067 47515 50101 47545
rect 50067 47443 50101 47477
rect 50525 48667 50559 48701
rect 50525 48599 50559 48629
rect 50525 48595 50559 48599
rect 50525 48531 50559 48557
rect 50525 48523 50559 48531
rect 50525 48463 50559 48485
rect 50525 48451 50559 48463
rect 50525 48395 50559 48413
rect 50525 48379 50559 48395
rect 50525 48327 50559 48341
rect 50525 48307 50559 48327
rect 50525 48259 50559 48269
rect 50525 48235 50559 48259
rect 50525 48191 50559 48197
rect 50525 48163 50559 48191
rect 50525 48123 50559 48125
rect 50525 48091 50559 48123
rect 50525 48021 50559 48053
rect 50525 48019 50559 48021
rect 50525 47953 50559 47981
rect 50525 47947 50559 47953
rect 50525 47885 50559 47909
rect 50525 47875 50559 47885
rect 50525 47817 50559 47837
rect 50525 47803 50559 47817
rect 50525 47749 50559 47765
rect 50525 47731 50559 47749
rect 50525 47681 50559 47693
rect 50525 47659 50559 47681
rect 50525 47613 50559 47621
rect 50525 47587 50559 47613
rect 50525 47545 50559 47549
rect 50525 47515 50559 47545
rect 50525 47443 50559 47477
rect 50983 48667 51017 48701
rect 50983 48599 51017 48629
rect 50983 48595 51017 48599
rect 50983 48531 51017 48557
rect 50983 48523 51017 48531
rect 50983 48463 51017 48485
rect 50983 48451 51017 48463
rect 50983 48395 51017 48413
rect 50983 48379 51017 48395
rect 50983 48327 51017 48341
rect 50983 48307 51017 48327
rect 50983 48259 51017 48269
rect 50983 48235 51017 48259
rect 50983 48191 51017 48197
rect 50983 48163 51017 48191
rect 50983 48123 51017 48125
rect 50983 48091 51017 48123
rect 50983 48021 51017 48053
rect 50983 48019 51017 48021
rect 50983 47953 51017 47981
rect 50983 47947 51017 47953
rect 50983 47885 51017 47909
rect 50983 47875 51017 47885
rect 50983 47817 51017 47837
rect 50983 47803 51017 47817
rect 50983 47749 51017 47765
rect 50983 47731 51017 47749
rect 50983 47681 51017 47693
rect 50983 47659 51017 47681
rect 50983 47613 51017 47621
rect 50983 47587 51017 47613
rect 50983 47545 51017 47549
rect 50983 47515 51017 47545
rect 50983 47443 51017 47477
rect 51441 48667 51475 48701
rect 51441 48599 51475 48629
rect 51441 48595 51475 48599
rect 51441 48531 51475 48557
rect 51441 48523 51475 48531
rect 51441 48463 51475 48485
rect 51441 48451 51475 48463
rect 51441 48395 51475 48413
rect 51441 48379 51475 48395
rect 51441 48327 51475 48341
rect 51441 48307 51475 48327
rect 51441 48259 51475 48269
rect 51441 48235 51475 48259
rect 51441 48191 51475 48197
rect 51441 48163 51475 48191
rect 51441 48123 51475 48125
rect 51441 48091 51475 48123
rect 51441 48021 51475 48053
rect 51441 48019 51475 48021
rect 51441 47953 51475 47981
rect 51441 47947 51475 47953
rect 51441 47885 51475 47909
rect 51441 47875 51475 47885
rect 51441 47817 51475 47837
rect 51441 47803 51475 47817
rect 51441 47749 51475 47765
rect 51441 47731 51475 47749
rect 51441 47681 51475 47693
rect 51441 47659 51475 47681
rect 51441 47613 51475 47621
rect 51441 47587 51475 47613
rect 51441 47545 51475 47549
rect 51441 47515 51475 47545
rect 51441 47443 51475 47477
rect 51899 48667 51933 48701
rect 51899 48599 51933 48629
rect 51899 48595 51933 48599
rect 51899 48531 51933 48557
rect 51899 48523 51933 48531
rect 51899 48463 51933 48485
rect 51899 48451 51933 48463
rect 51899 48395 51933 48413
rect 51899 48379 51933 48395
rect 51899 48327 51933 48341
rect 51899 48307 51933 48327
rect 51899 48259 51933 48269
rect 51899 48235 51933 48259
rect 51899 48191 51933 48197
rect 51899 48163 51933 48191
rect 51899 48123 51933 48125
rect 51899 48091 51933 48123
rect 51899 48021 51933 48053
rect 51899 48019 51933 48021
rect 51899 47953 51933 47981
rect 51899 47947 51933 47953
rect 51899 47885 51933 47909
rect 51899 47875 51933 47885
rect 51899 47817 51933 47837
rect 51899 47803 51933 47817
rect 51899 47749 51933 47765
rect 51899 47731 51933 47749
rect 51899 47681 51933 47693
rect 51899 47659 51933 47681
rect 51899 47613 51933 47621
rect 51899 47587 51933 47613
rect 51899 47545 51933 47549
rect 51899 47515 51933 47545
rect 51899 47443 51933 47477
rect 52357 48667 52391 48701
rect 52357 48599 52391 48629
rect 52357 48595 52391 48599
rect 52357 48531 52391 48557
rect 52357 48523 52391 48531
rect 52357 48463 52391 48485
rect 52357 48451 52391 48463
rect 52357 48395 52391 48413
rect 52357 48379 52391 48395
rect 52357 48327 52391 48341
rect 52357 48307 52391 48327
rect 52357 48259 52391 48269
rect 52357 48235 52391 48259
rect 52357 48191 52391 48197
rect 52357 48163 52391 48191
rect 52357 48123 52391 48125
rect 52357 48091 52391 48123
rect 52357 48021 52391 48053
rect 52357 48019 52391 48021
rect 52357 47953 52391 47981
rect 52357 47947 52391 47953
rect 52357 47885 52391 47909
rect 52357 47875 52391 47885
rect 52357 47817 52391 47837
rect 52357 47803 52391 47817
rect 52357 47749 52391 47765
rect 52357 47731 52391 47749
rect 52357 47681 52391 47693
rect 52357 47659 52391 47681
rect 52357 47613 52391 47621
rect 52357 47587 52391 47613
rect 52357 47545 52391 47549
rect 52357 47515 52391 47545
rect 52357 47443 52391 47477
rect 24041 47209 24075 47243
rect 29469 47209 29503 47243
rect 6101 47055 6135 47089
rect 6501 47055 6535 47089
rect 6901 47055 6935 47089
rect 7301 47055 7335 47089
rect 7701 47055 7735 47089
rect 8101 47055 8135 47089
rect 8501 47055 8535 47089
rect 8901 47055 8935 47089
rect 9301 47055 9335 47089
rect 9701 47055 9735 47089
rect 10101 47055 10135 47089
rect 10501 47055 10535 47089
rect 10901 47055 10935 47089
rect 11301 47055 11335 47089
rect 11701 47055 11735 47089
rect 12101 47055 12135 47089
rect 12501 47055 12535 47089
rect 12901 47055 12935 47089
rect 13549 47055 13583 47089
rect 13949 47055 13983 47089
rect 14349 47055 14383 47089
rect 14749 47055 14783 47089
rect 15149 47055 15183 47089
rect 15549 47055 15583 47089
rect 15949 47055 15983 47089
rect 16349 47055 16383 47089
rect 16749 47055 16783 47089
rect 17149 47055 17183 47089
rect 17549 47055 17583 47089
rect 17949 47055 17983 47089
rect 18349 47055 18383 47089
rect 18749 47055 18783 47089
rect 19149 47055 19183 47089
rect 19549 47055 19583 47089
rect 19949 47055 19983 47089
rect 20349 47055 20383 47089
rect 21015 47055 21049 47089
rect 21215 47055 21249 47089
rect 21415 47055 21449 47089
rect 21615 47055 21649 47089
rect 21815 47055 21849 47089
rect 22015 47055 22049 47089
rect 22215 47055 22249 47089
rect 22415 47055 22449 47089
rect 22615 47055 22649 47089
rect 22815 47055 22849 47089
rect 23015 47055 23049 47089
rect 24101 47055 24135 47089
rect 25013 47055 25047 47089
rect 25413 47055 25447 47089
rect 25813 47055 25847 47089
rect 26213 47055 26247 47089
rect 26613 47055 26647 47089
rect 27013 47055 27047 47089
rect 27413 47055 27447 47089
rect 27813 47055 27847 47089
rect 28213 47055 28247 47089
rect 28613 47055 28647 47089
rect 29013 47055 29047 47089
rect 29413 47055 29447 47089
rect 29813 47055 29847 47089
rect 30213 47055 30247 47089
rect 30613 47055 30647 47089
rect 31013 47055 31047 47089
rect 31413 47055 31447 47089
rect 31813 47055 31847 47089
rect 32213 47055 32247 47089
rect 32613 47055 32647 47089
rect 33013 47055 33047 47089
rect 33413 47055 33447 47089
rect 33813 47055 33847 47089
rect 34213 47055 34247 47089
rect 34613 47055 34647 47089
rect 35013 47055 35047 47089
rect 35413 47055 35447 47089
rect 35813 47055 35847 47089
rect 36213 47055 36247 47089
rect 36613 47055 36647 47089
rect 37013 47055 37047 47089
rect 37413 47055 37447 47089
rect 37813 47055 37847 47089
rect 38213 47055 38247 47089
rect 38613 47055 38647 47089
rect 39013 47055 39047 47089
rect 39413 47055 39447 47089
rect 39813 47055 39847 47089
rect 40213 47055 40247 47089
rect 40613 47055 40647 47089
rect 41013 47055 41047 47089
rect 41413 47055 41447 47089
rect 41813 47055 41847 47089
rect 42213 47055 42247 47089
rect 42613 47055 42647 47089
rect 43013 47055 43047 47089
rect 43413 47055 43447 47089
rect 43813 47055 43847 47089
rect 44213 47055 44247 47089
rect 44613 47055 44647 47089
rect 45013 47055 45047 47089
rect 45413 47055 45447 47089
rect 45813 47055 45847 47089
rect 46213 47055 46247 47089
rect 46613 47055 46647 47089
rect 47013 47055 47047 47089
rect 47413 47055 47447 47089
rect 47813 47055 47847 47089
rect 48213 47055 48247 47089
rect 48613 47055 48647 47089
rect 49013 47055 49047 47089
rect 49413 47055 49447 47089
rect 49813 47055 49847 47089
rect 50213 47055 50247 47089
rect 50613 47055 50647 47089
rect 51013 47055 51047 47089
rect 51413 47055 51447 47089
rect 51813 47055 51847 47089
rect 52213 47055 52247 47089
rect 6101 45175 6135 45209
rect 6501 45175 6535 45209
rect 6901 45175 6935 45209
rect 7301 45175 7335 45209
rect 7701 45175 7735 45209
rect 8101 45175 8135 45209
rect 8501 45175 8535 45209
rect 8901 45175 8935 45209
rect 9301 45175 9335 45209
rect 9701 45175 9735 45209
rect 10101 45175 10135 45209
rect 10501 45175 10535 45209
rect 10901 45175 10935 45209
rect 11301 45175 11335 45209
rect 11701 45175 11735 45209
rect 12101 45175 12135 45209
rect 12501 45175 12535 45209
rect 12901 45175 12935 45209
rect 14301 45175 14335 45209
rect 15213 45175 15247 45209
rect 15613 45175 15647 45209
rect 16013 45175 16047 45209
rect 16413 45175 16447 45209
rect 16813 45175 16847 45209
rect 17213 45175 17247 45209
rect 17613 45175 17647 45209
rect 18013 45175 18047 45209
rect 18413 45175 18447 45209
rect 18813 45175 18847 45209
rect 19213 45175 19247 45209
rect 19613 45175 19647 45209
rect 20013 45175 20047 45209
rect 20413 45175 20447 45209
rect 20813 45175 20847 45209
rect 21213 45175 21247 45209
rect 21613 45175 21647 45209
rect 22013 45175 22047 45209
rect 22413 45175 22447 45209
rect 22813 45175 22847 45209
rect 23213 45175 23247 45209
rect 23613 45175 23647 45209
rect 24013 45175 24047 45209
rect 24413 45175 24447 45209
rect 24813 45175 24847 45209
rect 25213 45175 25247 45209
rect 25613 45175 25647 45209
rect 26013 45175 26047 45209
rect 26413 45175 26447 45209
rect 26813 45175 26847 45209
rect 27213 45175 27247 45209
rect 27613 45175 27647 45209
rect 28013 45175 28047 45209
rect 28413 45175 28447 45209
rect 28813 45175 28847 45209
rect 29213 45175 29247 45209
rect 29613 45175 29647 45209
rect 30013 45175 30047 45209
rect 30413 45175 30447 45209
rect 30813 45175 30847 45209
rect 31213 45175 31247 45209
rect 31613 45175 31647 45209
rect 32013 45175 32047 45209
rect 32413 45175 32447 45209
rect 32813 45175 32847 45209
rect 33213 45175 33247 45209
rect 33613 45175 33647 45209
rect 34013 45175 34047 45209
rect 34413 45175 34447 45209
rect 34813 45175 34847 45209
rect 35213 45175 35247 45209
rect 35613 45175 35647 45209
rect 36013 45175 36047 45209
rect 36413 45175 36447 45209
rect 36813 45175 36847 45209
rect 37213 45175 37247 45209
rect 37613 45175 37647 45209
rect 38013 45175 38047 45209
rect 38413 45175 38447 45209
rect 38813 45175 38847 45209
rect 39213 45175 39247 45209
rect 39613 45175 39647 45209
rect 40013 45175 40047 45209
rect 40413 45175 40447 45209
rect 40813 45175 40847 45209
rect 41213 45175 41247 45209
rect 41613 45175 41647 45209
rect 42013 45175 42047 45209
rect 42413 45175 42447 45209
rect 43143 45175 43177 45209
rect 43343 45175 43377 45209
rect 43543 45175 43577 45209
rect 43743 45175 43777 45209
rect 43943 45175 43977 45209
rect 44143 45175 44177 45209
rect 44343 45175 44377 45209
rect 44543 45175 44577 45209
rect 44743 45175 44777 45209
rect 44943 45175 44977 45209
rect 45143 45175 45177 45209
rect 45343 45175 45377 45209
rect 45543 45175 45577 45209
rect 45743 45175 45777 45209
rect 45943 45175 45977 45209
rect 46143 45175 46177 45209
rect 46343 45175 46377 45209
rect 46543 45175 46577 45209
rect 46743 45175 46777 45209
rect 46943 45175 46977 45209
rect 47143 45175 47177 45209
rect 47343 45175 47377 45209
rect 47543 45175 47577 45209
rect 47743 45175 47777 45209
rect 47943 45175 47977 45209
rect 48143 45175 48177 45209
rect 48343 45175 48377 45209
rect 48543 45175 48577 45209
rect 48743 45175 48777 45209
rect 48943 45175 48977 45209
rect 49143 45175 49177 45209
rect 49343 45175 49377 45209
rect 49543 45175 49577 45209
rect 49743 45175 49777 45209
rect 49943 45175 49977 45209
rect 50143 45175 50177 45209
rect 50343 45175 50377 45209
rect 50543 45175 50577 45209
rect 50743 45175 50777 45209
rect 50943 45175 50977 45209
rect 51143 45175 51177 45209
rect 51343 45175 51377 45209
rect 51543 45175 51577 45209
rect 51743 45175 51777 45209
rect 51943 45175 51977 45209
rect 52143 45175 52177 45209
rect 15077 44907 15111 44941
rect 15077 44839 15111 44869
rect 15077 44835 15111 44839
rect 15077 44771 15111 44797
rect 15077 44763 15111 44771
rect 14130 44669 14164 44689
rect 14130 44655 14164 44669
rect 14130 44601 14164 44617
rect 14130 44583 14164 44601
rect 14130 44533 14164 44545
rect 14130 44511 14164 44533
rect 14130 44465 14164 44473
rect 14130 44439 14164 44465
rect 14130 44397 14164 44401
rect 14130 44367 14164 44397
rect 14130 44295 14164 44329
rect 14130 44227 14164 44257
rect 14130 44223 14164 44227
rect 14130 44159 14164 44185
rect 14130 44151 14164 44159
rect 14130 44091 14164 44113
rect 14130 44079 14164 44091
rect 14130 44023 14164 44041
rect 14130 44007 14164 44023
rect 14130 43955 14164 43969
rect 14130 43935 14164 43955
rect 14588 44669 14622 44689
rect 14588 44655 14622 44669
rect 14588 44601 14622 44617
rect 14588 44583 14622 44601
rect 14588 44533 14622 44545
rect 14588 44511 14622 44533
rect 14588 44465 14622 44473
rect 14588 44439 14622 44465
rect 14588 44397 14622 44401
rect 14588 44367 14622 44397
rect 14588 44295 14622 44329
rect 14588 44227 14622 44257
rect 14588 44223 14622 44227
rect 14588 44159 14622 44185
rect 14588 44151 14622 44159
rect 14588 44091 14622 44113
rect 14588 44079 14622 44091
rect 14588 44023 14622 44041
rect 14588 44007 14622 44023
rect 14588 43955 14622 43969
rect 14588 43935 14622 43955
rect 15077 44703 15111 44725
rect 15077 44691 15111 44703
rect 15077 44635 15111 44653
rect 15077 44619 15111 44635
rect 15077 44567 15111 44581
rect 15077 44547 15111 44567
rect 15077 44499 15111 44509
rect 15077 44475 15111 44499
rect 15077 44431 15111 44437
rect 15077 44403 15111 44431
rect 15077 44363 15111 44365
rect 15077 44331 15111 44363
rect 15077 44261 15111 44293
rect 15077 44259 15111 44261
rect 15077 44193 15111 44221
rect 15077 44187 15111 44193
rect 15077 44125 15111 44149
rect 15077 44115 15111 44125
rect 15077 44057 15111 44077
rect 15077 44043 15111 44057
rect 15077 43989 15111 44005
rect 15077 43971 15111 43989
rect 15077 43921 15111 43933
rect 15077 43899 15111 43921
rect 15077 43853 15111 43861
rect 15077 43827 15111 43853
rect 15077 43785 15111 43789
rect 15077 43755 15111 43785
rect 14381 43673 14415 43707
rect 15077 43683 15111 43717
rect 15535 44907 15569 44941
rect 15535 44839 15569 44869
rect 15535 44835 15569 44839
rect 15535 44771 15569 44797
rect 15535 44763 15569 44771
rect 15535 44703 15569 44725
rect 15535 44691 15569 44703
rect 15535 44635 15569 44653
rect 15535 44619 15569 44635
rect 15535 44567 15569 44581
rect 15535 44547 15569 44567
rect 15535 44499 15569 44509
rect 15535 44475 15569 44499
rect 15535 44431 15569 44437
rect 15535 44403 15569 44431
rect 15535 44363 15569 44365
rect 15535 44331 15569 44363
rect 15535 44261 15569 44293
rect 15535 44259 15569 44261
rect 15535 44193 15569 44221
rect 15535 44187 15569 44193
rect 15535 44125 15569 44149
rect 15535 44115 15569 44125
rect 15535 44057 15569 44077
rect 15535 44043 15569 44057
rect 15535 43989 15569 44005
rect 15535 43971 15569 43989
rect 15535 43921 15569 43933
rect 15535 43899 15569 43921
rect 15535 43853 15569 43861
rect 15535 43827 15569 43853
rect 15535 43785 15569 43789
rect 15535 43755 15569 43785
rect 15535 43683 15569 43717
rect 15993 44907 16027 44941
rect 15993 44839 16027 44869
rect 15993 44835 16027 44839
rect 15993 44771 16027 44797
rect 15993 44763 16027 44771
rect 15993 44703 16027 44725
rect 15993 44691 16027 44703
rect 15993 44635 16027 44653
rect 15993 44619 16027 44635
rect 15993 44567 16027 44581
rect 15993 44547 16027 44567
rect 15993 44499 16027 44509
rect 15993 44475 16027 44499
rect 15993 44431 16027 44437
rect 15993 44403 16027 44431
rect 15993 44363 16027 44365
rect 15993 44331 16027 44363
rect 15993 44261 16027 44293
rect 15993 44259 16027 44261
rect 15993 44193 16027 44221
rect 15993 44187 16027 44193
rect 15993 44125 16027 44149
rect 15993 44115 16027 44125
rect 15993 44057 16027 44077
rect 15993 44043 16027 44057
rect 15993 43989 16027 44005
rect 15993 43971 16027 43989
rect 15993 43921 16027 43933
rect 15993 43899 16027 43921
rect 15993 43853 16027 43861
rect 15993 43827 16027 43853
rect 15993 43785 16027 43789
rect 15993 43755 16027 43785
rect 15993 43683 16027 43717
rect 16451 44907 16485 44941
rect 16451 44839 16485 44869
rect 16451 44835 16485 44839
rect 16451 44771 16485 44797
rect 16451 44763 16485 44771
rect 16451 44703 16485 44725
rect 16451 44691 16485 44703
rect 16451 44635 16485 44653
rect 16451 44619 16485 44635
rect 16451 44567 16485 44581
rect 16451 44547 16485 44567
rect 16451 44499 16485 44509
rect 16451 44475 16485 44499
rect 16451 44431 16485 44437
rect 16451 44403 16485 44431
rect 16451 44363 16485 44365
rect 16451 44331 16485 44363
rect 16451 44261 16485 44293
rect 16451 44259 16485 44261
rect 16451 44193 16485 44221
rect 16451 44187 16485 44193
rect 16451 44125 16485 44149
rect 16451 44115 16485 44125
rect 16451 44057 16485 44077
rect 16451 44043 16485 44057
rect 16451 43989 16485 44005
rect 16451 43971 16485 43989
rect 16451 43921 16485 43933
rect 16451 43899 16485 43921
rect 16451 43853 16485 43861
rect 16451 43827 16485 43853
rect 16451 43785 16485 43789
rect 16451 43755 16485 43785
rect 16451 43683 16485 43717
rect 16909 44907 16943 44941
rect 16909 44839 16943 44869
rect 16909 44835 16943 44839
rect 16909 44771 16943 44797
rect 16909 44763 16943 44771
rect 16909 44703 16943 44725
rect 16909 44691 16943 44703
rect 16909 44635 16943 44653
rect 16909 44619 16943 44635
rect 16909 44567 16943 44581
rect 16909 44547 16943 44567
rect 16909 44499 16943 44509
rect 16909 44475 16943 44499
rect 16909 44431 16943 44437
rect 16909 44403 16943 44431
rect 16909 44363 16943 44365
rect 16909 44331 16943 44363
rect 16909 44261 16943 44293
rect 16909 44259 16943 44261
rect 16909 44193 16943 44221
rect 16909 44187 16943 44193
rect 16909 44125 16943 44149
rect 16909 44115 16943 44125
rect 16909 44057 16943 44077
rect 16909 44043 16943 44057
rect 16909 43989 16943 44005
rect 16909 43971 16943 43989
rect 16909 43921 16943 43933
rect 16909 43899 16943 43921
rect 16909 43853 16943 43861
rect 16909 43827 16943 43853
rect 16909 43785 16943 43789
rect 16909 43755 16943 43785
rect 16909 43683 16943 43717
rect 17367 44907 17401 44941
rect 17367 44839 17401 44869
rect 17367 44835 17401 44839
rect 17367 44771 17401 44797
rect 17367 44763 17401 44771
rect 17367 44703 17401 44725
rect 17367 44691 17401 44703
rect 17367 44635 17401 44653
rect 17367 44619 17401 44635
rect 17367 44567 17401 44581
rect 17367 44547 17401 44567
rect 17367 44499 17401 44509
rect 17367 44475 17401 44499
rect 17367 44431 17401 44437
rect 17367 44403 17401 44431
rect 17367 44363 17401 44365
rect 17367 44331 17401 44363
rect 17367 44261 17401 44293
rect 17367 44259 17401 44261
rect 17367 44193 17401 44221
rect 17367 44187 17401 44193
rect 17367 44125 17401 44149
rect 17367 44115 17401 44125
rect 17367 44057 17401 44077
rect 17367 44043 17401 44057
rect 17367 43989 17401 44005
rect 17367 43971 17401 43989
rect 17367 43921 17401 43933
rect 17367 43899 17401 43921
rect 17367 43853 17401 43861
rect 17367 43827 17401 43853
rect 17367 43785 17401 43789
rect 17367 43755 17401 43785
rect 17367 43683 17401 43717
rect 17825 44907 17859 44941
rect 17825 44839 17859 44869
rect 17825 44835 17859 44839
rect 17825 44771 17859 44797
rect 17825 44763 17859 44771
rect 17825 44703 17859 44725
rect 17825 44691 17859 44703
rect 17825 44635 17859 44653
rect 17825 44619 17859 44635
rect 17825 44567 17859 44581
rect 17825 44547 17859 44567
rect 17825 44499 17859 44509
rect 17825 44475 17859 44499
rect 17825 44431 17859 44437
rect 17825 44403 17859 44431
rect 17825 44363 17859 44365
rect 17825 44331 17859 44363
rect 17825 44261 17859 44293
rect 17825 44259 17859 44261
rect 17825 44193 17859 44221
rect 17825 44187 17859 44193
rect 17825 44125 17859 44149
rect 17825 44115 17859 44125
rect 17825 44057 17859 44077
rect 17825 44043 17859 44057
rect 17825 43989 17859 44005
rect 17825 43971 17859 43989
rect 17825 43921 17859 43933
rect 17825 43899 17859 43921
rect 17825 43853 17859 43861
rect 17825 43827 17859 43853
rect 17825 43785 17859 43789
rect 17825 43755 17859 43785
rect 17825 43683 17859 43717
rect 18283 44907 18317 44941
rect 18283 44839 18317 44869
rect 18283 44835 18317 44839
rect 18283 44771 18317 44797
rect 18283 44763 18317 44771
rect 18283 44703 18317 44725
rect 18283 44691 18317 44703
rect 18283 44635 18317 44653
rect 18283 44619 18317 44635
rect 18283 44567 18317 44581
rect 18283 44547 18317 44567
rect 18283 44499 18317 44509
rect 18283 44475 18317 44499
rect 18283 44431 18317 44437
rect 18283 44403 18317 44431
rect 18283 44363 18317 44365
rect 18283 44331 18317 44363
rect 18283 44261 18317 44293
rect 18283 44259 18317 44261
rect 18283 44193 18317 44221
rect 18283 44187 18317 44193
rect 18283 44125 18317 44149
rect 18283 44115 18317 44125
rect 18283 44057 18317 44077
rect 18283 44043 18317 44057
rect 18283 43989 18317 44005
rect 18283 43971 18317 43989
rect 18283 43921 18317 43933
rect 18283 43899 18317 43921
rect 18283 43853 18317 43861
rect 18283 43827 18317 43853
rect 18283 43785 18317 43789
rect 18283 43755 18317 43785
rect 18283 43683 18317 43717
rect 18741 44907 18775 44941
rect 18741 44839 18775 44869
rect 18741 44835 18775 44839
rect 18741 44771 18775 44797
rect 18741 44763 18775 44771
rect 18741 44703 18775 44725
rect 18741 44691 18775 44703
rect 18741 44635 18775 44653
rect 18741 44619 18775 44635
rect 18741 44567 18775 44581
rect 18741 44547 18775 44567
rect 18741 44499 18775 44509
rect 18741 44475 18775 44499
rect 18741 44431 18775 44437
rect 18741 44403 18775 44431
rect 18741 44363 18775 44365
rect 18741 44331 18775 44363
rect 18741 44261 18775 44293
rect 18741 44259 18775 44261
rect 18741 44193 18775 44221
rect 18741 44187 18775 44193
rect 18741 44125 18775 44149
rect 18741 44115 18775 44125
rect 18741 44057 18775 44077
rect 18741 44043 18775 44057
rect 18741 43989 18775 44005
rect 18741 43971 18775 43989
rect 18741 43921 18775 43933
rect 18741 43899 18775 43921
rect 18741 43853 18775 43861
rect 18741 43827 18775 43853
rect 18741 43785 18775 43789
rect 18741 43755 18775 43785
rect 18741 43683 18775 43717
rect 19199 44907 19233 44941
rect 19199 44839 19233 44869
rect 19199 44835 19233 44839
rect 19199 44771 19233 44797
rect 19199 44763 19233 44771
rect 19199 44703 19233 44725
rect 19199 44691 19233 44703
rect 19199 44635 19233 44653
rect 19199 44619 19233 44635
rect 19199 44567 19233 44581
rect 19199 44547 19233 44567
rect 19199 44499 19233 44509
rect 19199 44475 19233 44499
rect 19199 44431 19233 44437
rect 19199 44403 19233 44431
rect 19199 44363 19233 44365
rect 19199 44331 19233 44363
rect 19199 44261 19233 44293
rect 19199 44259 19233 44261
rect 19199 44193 19233 44221
rect 19199 44187 19233 44193
rect 19199 44125 19233 44149
rect 19199 44115 19233 44125
rect 19199 44057 19233 44077
rect 19199 44043 19233 44057
rect 19199 43989 19233 44005
rect 19199 43971 19233 43989
rect 19199 43921 19233 43933
rect 19199 43899 19233 43921
rect 19199 43853 19233 43861
rect 19199 43827 19233 43853
rect 19199 43785 19233 43789
rect 19199 43755 19233 43785
rect 19199 43683 19233 43717
rect 19657 44907 19691 44941
rect 19657 44839 19691 44869
rect 19657 44835 19691 44839
rect 19657 44771 19691 44797
rect 19657 44763 19691 44771
rect 19657 44703 19691 44725
rect 19657 44691 19691 44703
rect 19657 44635 19691 44653
rect 19657 44619 19691 44635
rect 19657 44567 19691 44581
rect 19657 44547 19691 44567
rect 19657 44499 19691 44509
rect 19657 44475 19691 44499
rect 19657 44431 19691 44437
rect 19657 44403 19691 44431
rect 19657 44363 19691 44365
rect 19657 44331 19691 44363
rect 19657 44261 19691 44293
rect 19657 44259 19691 44261
rect 19657 44193 19691 44221
rect 19657 44187 19691 44193
rect 19657 44125 19691 44149
rect 19657 44115 19691 44125
rect 19657 44057 19691 44077
rect 19657 44043 19691 44057
rect 19657 43989 19691 44005
rect 19657 43971 19691 43989
rect 19657 43921 19691 43933
rect 19657 43899 19691 43921
rect 19657 43853 19691 43861
rect 19657 43827 19691 43853
rect 19657 43785 19691 43789
rect 19657 43755 19691 43785
rect 19657 43683 19691 43717
rect 20115 44907 20149 44941
rect 20115 44839 20149 44869
rect 20115 44835 20149 44839
rect 20115 44771 20149 44797
rect 20115 44763 20149 44771
rect 20115 44703 20149 44725
rect 20115 44691 20149 44703
rect 20115 44635 20149 44653
rect 20115 44619 20149 44635
rect 20115 44567 20149 44581
rect 20115 44547 20149 44567
rect 20115 44499 20149 44509
rect 20115 44475 20149 44499
rect 20115 44431 20149 44437
rect 20115 44403 20149 44431
rect 20115 44363 20149 44365
rect 20115 44331 20149 44363
rect 20115 44261 20149 44293
rect 20115 44259 20149 44261
rect 20115 44193 20149 44221
rect 20115 44187 20149 44193
rect 20115 44125 20149 44149
rect 20115 44115 20149 44125
rect 20115 44057 20149 44077
rect 20115 44043 20149 44057
rect 20115 43989 20149 44005
rect 20115 43971 20149 43989
rect 20115 43921 20149 43933
rect 20115 43899 20149 43921
rect 20115 43853 20149 43861
rect 20115 43827 20149 43853
rect 20115 43785 20149 43789
rect 20115 43755 20149 43785
rect 20115 43683 20149 43717
rect 20573 44907 20607 44941
rect 20573 44839 20607 44869
rect 20573 44835 20607 44839
rect 20573 44771 20607 44797
rect 20573 44763 20607 44771
rect 20573 44703 20607 44725
rect 20573 44691 20607 44703
rect 20573 44635 20607 44653
rect 20573 44619 20607 44635
rect 20573 44567 20607 44581
rect 20573 44547 20607 44567
rect 20573 44499 20607 44509
rect 20573 44475 20607 44499
rect 20573 44431 20607 44437
rect 20573 44403 20607 44431
rect 20573 44363 20607 44365
rect 20573 44331 20607 44363
rect 20573 44261 20607 44293
rect 20573 44259 20607 44261
rect 20573 44193 20607 44221
rect 20573 44187 20607 44193
rect 20573 44125 20607 44149
rect 20573 44115 20607 44125
rect 20573 44057 20607 44077
rect 20573 44043 20607 44057
rect 20573 43989 20607 44005
rect 20573 43971 20607 43989
rect 20573 43921 20607 43933
rect 20573 43899 20607 43921
rect 20573 43853 20607 43861
rect 20573 43827 20607 43853
rect 20573 43785 20607 43789
rect 20573 43755 20607 43785
rect 20573 43683 20607 43717
rect 21031 44907 21065 44941
rect 21031 44839 21065 44869
rect 21031 44835 21065 44839
rect 21031 44771 21065 44797
rect 21031 44763 21065 44771
rect 21031 44703 21065 44725
rect 21031 44691 21065 44703
rect 21031 44635 21065 44653
rect 21031 44619 21065 44635
rect 21031 44567 21065 44581
rect 21031 44547 21065 44567
rect 21031 44499 21065 44509
rect 21031 44475 21065 44499
rect 21031 44431 21065 44437
rect 21031 44403 21065 44431
rect 21031 44363 21065 44365
rect 21031 44331 21065 44363
rect 21031 44261 21065 44293
rect 21031 44259 21065 44261
rect 21031 44193 21065 44221
rect 21031 44187 21065 44193
rect 21031 44125 21065 44149
rect 21031 44115 21065 44125
rect 21031 44057 21065 44077
rect 21031 44043 21065 44057
rect 21031 43989 21065 44005
rect 21031 43971 21065 43989
rect 21031 43921 21065 43933
rect 21031 43899 21065 43921
rect 21031 43853 21065 43861
rect 21031 43827 21065 43853
rect 21031 43785 21065 43789
rect 21031 43755 21065 43785
rect 21031 43683 21065 43717
rect 21489 44907 21523 44941
rect 21489 44839 21523 44869
rect 21489 44835 21523 44839
rect 21489 44771 21523 44797
rect 21489 44763 21523 44771
rect 21489 44703 21523 44725
rect 21489 44691 21523 44703
rect 21489 44635 21523 44653
rect 21489 44619 21523 44635
rect 21489 44567 21523 44581
rect 21489 44547 21523 44567
rect 21489 44499 21523 44509
rect 21489 44475 21523 44499
rect 21489 44431 21523 44437
rect 21489 44403 21523 44431
rect 21489 44363 21523 44365
rect 21489 44331 21523 44363
rect 21489 44261 21523 44293
rect 21489 44259 21523 44261
rect 21489 44193 21523 44221
rect 21489 44187 21523 44193
rect 21489 44125 21523 44149
rect 21489 44115 21523 44125
rect 21489 44057 21523 44077
rect 21489 44043 21523 44057
rect 21489 43989 21523 44005
rect 21489 43971 21523 43989
rect 21489 43921 21523 43933
rect 21489 43899 21523 43921
rect 21489 43853 21523 43861
rect 21489 43827 21523 43853
rect 21489 43785 21523 43789
rect 21489 43755 21523 43785
rect 21489 43683 21523 43717
rect 21947 44907 21981 44941
rect 21947 44839 21981 44869
rect 21947 44835 21981 44839
rect 21947 44771 21981 44797
rect 21947 44763 21981 44771
rect 21947 44703 21981 44725
rect 21947 44691 21981 44703
rect 21947 44635 21981 44653
rect 21947 44619 21981 44635
rect 21947 44567 21981 44581
rect 21947 44547 21981 44567
rect 21947 44499 21981 44509
rect 21947 44475 21981 44499
rect 21947 44431 21981 44437
rect 21947 44403 21981 44431
rect 21947 44363 21981 44365
rect 21947 44331 21981 44363
rect 21947 44261 21981 44293
rect 21947 44259 21981 44261
rect 21947 44193 21981 44221
rect 21947 44187 21981 44193
rect 21947 44125 21981 44149
rect 21947 44115 21981 44125
rect 21947 44057 21981 44077
rect 21947 44043 21981 44057
rect 21947 43989 21981 44005
rect 21947 43971 21981 43989
rect 21947 43921 21981 43933
rect 21947 43899 21981 43921
rect 21947 43853 21981 43861
rect 21947 43827 21981 43853
rect 21947 43785 21981 43789
rect 21947 43755 21981 43785
rect 21947 43683 21981 43717
rect 22405 44907 22439 44941
rect 22405 44839 22439 44869
rect 22405 44835 22439 44839
rect 22405 44771 22439 44797
rect 22405 44763 22439 44771
rect 22405 44703 22439 44725
rect 22405 44691 22439 44703
rect 22405 44635 22439 44653
rect 22405 44619 22439 44635
rect 22405 44567 22439 44581
rect 22405 44547 22439 44567
rect 22405 44499 22439 44509
rect 22405 44475 22439 44499
rect 22405 44431 22439 44437
rect 22405 44403 22439 44431
rect 22405 44363 22439 44365
rect 22405 44331 22439 44363
rect 22405 44261 22439 44293
rect 22405 44259 22439 44261
rect 22405 44193 22439 44221
rect 22405 44187 22439 44193
rect 22405 44125 22439 44149
rect 22405 44115 22439 44125
rect 22405 44057 22439 44077
rect 22405 44043 22439 44057
rect 22405 43989 22439 44005
rect 22405 43971 22439 43989
rect 22405 43921 22439 43933
rect 22405 43899 22439 43921
rect 22405 43853 22439 43861
rect 22405 43827 22439 43853
rect 22405 43785 22439 43789
rect 22405 43755 22439 43785
rect 22405 43683 22439 43717
rect 22863 44907 22897 44941
rect 22863 44839 22897 44869
rect 22863 44835 22897 44839
rect 22863 44771 22897 44797
rect 22863 44763 22897 44771
rect 22863 44703 22897 44725
rect 22863 44691 22897 44703
rect 22863 44635 22897 44653
rect 22863 44619 22897 44635
rect 22863 44567 22897 44581
rect 22863 44547 22897 44567
rect 22863 44499 22897 44509
rect 22863 44475 22897 44499
rect 22863 44431 22897 44437
rect 22863 44403 22897 44431
rect 22863 44363 22897 44365
rect 22863 44331 22897 44363
rect 22863 44261 22897 44293
rect 22863 44259 22897 44261
rect 22863 44193 22897 44221
rect 22863 44187 22897 44193
rect 22863 44125 22897 44149
rect 22863 44115 22897 44125
rect 22863 44057 22897 44077
rect 22863 44043 22897 44057
rect 22863 43989 22897 44005
rect 22863 43971 22897 43989
rect 22863 43921 22897 43933
rect 22863 43899 22897 43921
rect 22863 43853 22897 43861
rect 22863 43827 22897 43853
rect 22863 43785 22897 43789
rect 22863 43755 22897 43785
rect 22863 43683 22897 43717
rect 23321 44907 23355 44941
rect 23321 44839 23355 44869
rect 23321 44835 23355 44839
rect 23321 44771 23355 44797
rect 23321 44763 23355 44771
rect 23321 44703 23355 44725
rect 23321 44691 23355 44703
rect 23321 44635 23355 44653
rect 23321 44619 23355 44635
rect 23321 44567 23355 44581
rect 23321 44547 23355 44567
rect 23321 44499 23355 44509
rect 23321 44475 23355 44499
rect 23321 44431 23355 44437
rect 23321 44403 23355 44431
rect 23321 44363 23355 44365
rect 23321 44331 23355 44363
rect 23321 44261 23355 44293
rect 23321 44259 23355 44261
rect 23321 44193 23355 44221
rect 23321 44187 23355 44193
rect 23321 44125 23355 44149
rect 23321 44115 23355 44125
rect 23321 44057 23355 44077
rect 23321 44043 23355 44057
rect 23321 43989 23355 44005
rect 23321 43971 23355 43989
rect 23321 43921 23355 43933
rect 23321 43899 23355 43921
rect 23321 43853 23355 43861
rect 23321 43827 23355 43853
rect 23321 43785 23355 43789
rect 23321 43755 23355 43785
rect 23321 43683 23355 43717
rect 23779 44907 23813 44941
rect 23779 44839 23813 44869
rect 23779 44835 23813 44839
rect 23779 44771 23813 44797
rect 23779 44763 23813 44771
rect 23779 44703 23813 44725
rect 23779 44691 23813 44703
rect 23779 44635 23813 44653
rect 23779 44619 23813 44635
rect 23779 44567 23813 44581
rect 23779 44547 23813 44567
rect 23779 44499 23813 44509
rect 23779 44475 23813 44499
rect 23779 44431 23813 44437
rect 23779 44403 23813 44431
rect 23779 44363 23813 44365
rect 23779 44331 23813 44363
rect 23779 44261 23813 44293
rect 23779 44259 23813 44261
rect 23779 44193 23813 44221
rect 23779 44187 23813 44193
rect 23779 44125 23813 44149
rect 23779 44115 23813 44125
rect 23779 44057 23813 44077
rect 23779 44043 23813 44057
rect 23779 43989 23813 44005
rect 23779 43971 23813 43989
rect 23779 43921 23813 43933
rect 23779 43899 23813 43921
rect 23779 43853 23813 43861
rect 23779 43827 23813 43853
rect 23779 43785 23813 43789
rect 23779 43755 23813 43785
rect 23779 43683 23813 43717
rect 24237 44907 24271 44941
rect 24237 44839 24271 44869
rect 24237 44835 24271 44839
rect 24237 44771 24271 44797
rect 24237 44763 24271 44771
rect 24237 44703 24271 44725
rect 24237 44691 24271 44703
rect 24237 44635 24271 44653
rect 24237 44619 24271 44635
rect 24237 44567 24271 44581
rect 24237 44547 24271 44567
rect 24237 44499 24271 44509
rect 24237 44475 24271 44499
rect 24237 44431 24271 44437
rect 24237 44403 24271 44431
rect 24237 44363 24271 44365
rect 24237 44331 24271 44363
rect 24237 44261 24271 44293
rect 24237 44259 24271 44261
rect 24237 44193 24271 44221
rect 24237 44187 24271 44193
rect 24237 44125 24271 44149
rect 24237 44115 24271 44125
rect 24237 44057 24271 44077
rect 24237 44043 24271 44057
rect 24237 43989 24271 44005
rect 24237 43971 24271 43989
rect 24237 43921 24271 43933
rect 24237 43899 24271 43921
rect 24237 43853 24271 43861
rect 24237 43827 24271 43853
rect 24237 43785 24271 43789
rect 24237 43755 24271 43785
rect 24237 43683 24271 43717
rect 24695 44907 24729 44941
rect 24695 44839 24729 44869
rect 24695 44835 24729 44839
rect 24695 44771 24729 44797
rect 24695 44763 24729 44771
rect 24695 44703 24729 44725
rect 24695 44691 24729 44703
rect 24695 44635 24729 44653
rect 24695 44619 24729 44635
rect 24695 44567 24729 44581
rect 24695 44547 24729 44567
rect 24695 44499 24729 44509
rect 24695 44475 24729 44499
rect 24695 44431 24729 44437
rect 24695 44403 24729 44431
rect 24695 44363 24729 44365
rect 24695 44331 24729 44363
rect 24695 44261 24729 44293
rect 24695 44259 24729 44261
rect 24695 44193 24729 44221
rect 24695 44187 24729 44193
rect 24695 44125 24729 44149
rect 24695 44115 24729 44125
rect 24695 44057 24729 44077
rect 24695 44043 24729 44057
rect 24695 43989 24729 44005
rect 24695 43971 24729 43989
rect 24695 43921 24729 43933
rect 24695 43899 24729 43921
rect 24695 43853 24729 43861
rect 24695 43827 24729 43853
rect 24695 43785 24729 43789
rect 24695 43755 24729 43785
rect 24695 43683 24729 43717
rect 25153 44907 25187 44941
rect 25153 44839 25187 44869
rect 25153 44835 25187 44839
rect 25153 44771 25187 44797
rect 25153 44763 25187 44771
rect 25153 44703 25187 44725
rect 25153 44691 25187 44703
rect 25153 44635 25187 44653
rect 25153 44619 25187 44635
rect 25153 44567 25187 44581
rect 25153 44547 25187 44567
rect 25153 44499 25187 44509
rect 25153 44475 25187 44499
rect 25153 44431 25187 44437
rect 25153 44403 25187 44431
rect 25153 44363 25187 44365
rect 25153 44331 25187 44363
rect 25153 44261 25187 44293
rect 25153 44259 25187 44261
rect 25153 44193 25187 44221
rect 25153 44187 25187 44193
rect 25153 44125 25187 44149
rect 25153 44115 25187 44125
rect 25153 44057 25187 44077
rect 25153 44043 25187 44057
rect 25153 43989 25187 44005
rect 25153 43971 25187 43989
rect 25153 43921 25187 43933
rect 25153 43899 25187 43921
rect 25153 43853 25187 43861
rect 25153 43827 25187 43853
rect 25153 43785 25187 43789
rect 25153 43755 25187 43785
rect 25153 43683 25187 43717
rect 25611 44907 25645 44941
rect 25611 44839 25645 44869
rect 25611 44835 25645 44839
rect 25611 44771 25645 44797
rect 25611 44763 25645 44771
rect 25611 44703 25645 44725
rect 25611 44691 25645 44703
rect 25611 44635 25645 44653
rect 25611 44619 25645 44635
rect 25611 44567 25645 44581
rect 25611 44547 25645 44567
rect 25611 44499 25645 44509
rect 25611 44475 25645 44499
rect 25611 44431 25645 44437
rect 25611 44403 25645 44431
rect 25611 44363 25645 44365
rect 25611 44331 25645 44363
rect 25611 44261 25645 44293
rect 25611 44259 25645 44261
rect 25611 44193 25645 44221
rect 25611 44187 25645 44193
rect 25611 44125 25645 44149
rect 25611 44115 25645 44125
rect 25611 44057 25645 44077
rect 25611 44043 25645 44057
rect 25611 43989 25645 44005
rect 25611 43971 25645 43989
rect 25611 43921 25645 43933
rect 25611 43899 25645 43921
rect 25611 43853 25645 43861
rect 25611 43827 25645 43853
rect 25611 43785 25645 43789
rect 25611 43755 25645 43785
rect 25611 43683 25645 43717
rect 26069 44907 26103 44941
rect 26069 44839 26103 44869
rect 26069 44835 26103 44839
rect 26069 44771 26103 44797
rect 26069 44763 26103 44771
rect 26069 44703 26103 44725
rect 26069 44691 26103 44703
rect 26069 44635 26103 44653
rect 26069 44619 26103 44635
rect 26069 44567 26103 44581
rect 26069 44547 26103 44567
rect 26069 44499 26103 44509
rect 26069 44475 26103 44499
rect 26069 44431 26103 44437
rect 26069 44403 26103 44431
rect 26069 44363 26103 44365
rect 26069 44331 26103 44363
rect 26069 44261 26103 44293
rect 26069 44259 26103 44261
rect 26069 44193 26103 44221
rect 26069 44187 26103 44193
rect 26069 44125 26103 44149
rect 26069 44115 26103 44125
rect 26069 44057 26103 44077
rect 26069 44043 26103 44057
rect 26069 43989 26103 44005
rect 26069 43971 26103 43989
rect 26069 43921 26103 43933
rect 26069 43899 26103 43921
rect 26069 43853 26103 43861
rect 26069 43827 26103 43853
rect 26069 43785 26103 43789
rect 26069 43755 26103 43785
rect 26069 43683 26103 43717
rect 26527 44907 26561 44941
rect 26527 44839 26561 44869
rect 26527 44835 26561 44839
rect 26527 44771 26561 44797
rect 26527 44763 26561 44771
rect 26527 44703 26561 44725
rect 26527 44691 26561 44703
rect 26527 44635 26561 44653
rect 26527 44619 26561 44635
rect 26527 44567 26561 44581
rect 26527 44547 26561 44567
rect 26527 44499 26561 44509
rect 26527 44475 26561 44499
rect 26527 44431 26561 44437
rect 26527 44403 26561 44431
rect 26527 44363 26561 44365
rect 26527 44331 26561 44363
rect 26527 44261 26561 44293
rect 26527 44259 26561 44261
rect 26527 44193 26561 44221
rect 26527 44187 26561 44193
rect 26527 44125 26561 44149
rect 26527 44115 26561 44125
rect 26527 44057 26561 44077
rect 26527 44043 26561 44057
rect 26527 43989 26561 44005
rect 26527 43971 26561 43989
rect 26527 43921 26561 43933
rect 26527 43899 26561 43921
rect 26527 43853 26561 43861
rect 26527 43827 26561 43853
rect 26527 43785 26561 43789
rect 26527 43755 26561 43785
rect 26527 43683 26561 43717
rect 26985 44907 27019 44941
rect 26985 44839 27019 44869
rect 26985 44835 27019 44839
rect 26985 44771 27019 44797
rect 26985 44763 27019 44771
rect 26985 44703 27019 44725
rect 26985 44691 27019 44703
rect 26985 44635 27019 44653
rect 26985 44619 27019 44635
rect 26985 44567 27019 44581
rect 26985 44547 27019 44567
rect 26985 44499 27019 44509
rect 26985 44475 27019 44499
rect 26985 44431 27019 44437
rect 26985 44403 27019 44431
rect 26985 44363 27019 44365
rect 26985 44331 27019 44363
rect 26985 44261 27019 44293
rect 26985 44259 27019 44261
rect 26985 44193 27019 44221
rect 26985 44187 27019 44193
rect 26985 44125 27019 44149
rect 26985 44115 27019 44125
rect 26985 44057 27019 44077
rect 26985 44043 27019 44057
rect 26985 43989 27019 44005
rect 26985 43971 27019 43989
rect 26985 43921 27019 43933
rect 26985 43899 27019 43921
rect 26985 43853 27019 43861
rect 26985 43827 27019 43853
rect 26985 43785 27019 43789
rect 26985 43755 27019 43785
rect 26985 43683 27019 43717
rect 27443 44907 27477 44941
rect 27443 44839 27477 44869
rect 27443 44835 27477 44839
rect 27443 44771 27477 44797
rect 27443 44763 27477 44771
rect 27443 44703 27477 44725
rect 27443 44691 27477 44703
rect 27443 44635 27477 44653
rect 27443 44619 27477 44635
rect 27443 44567 27477 44581
rect 27443 44547 27477 44567
rect 27443 44499 27477 44509
rect 27443 44475 27477 44499
rect 27443 44431 27477 44437
rect 27443 44403 27477 44431
rect 27443 44363 27477 44365
rect 27443 44331 27477 44363
rect 27443 44261 27477 44293
rect 27443 44259 27477 44261
rect 27443 44193 27477 44221
rect 27443 44187 27477 44193
rect 27443 44125 27477 44149
rect 27443 44115 27477 44125
rect 27443 44057 27477 44077
rect 27443 44043 27477 44057
rect 27443 43989 27477 44005
rect 27443 43971 27477 43989
rect 27443 43921 27477 43933
rect 27443 43899 27477 43921
rect 27443 43853 27477 43861
rect 27443 43827 27477 43853
rect 27443 43785 27477 43789
rect 27443 43755 27477 43785
rect 27443 43683 27477 43717
rect 27901 44907 27935 44941
rect 27901 44839 27935 44869
rect 27901 44835 27935 44839
rect 27901 44771 27935 44797
rect 27901 44763 27935 44771
rect 27901 44703 27935 44725
rect 27901 44691 27935 44703
rect 27901 44635 27935 44653
rect 27901 44619 27935 44635
rect 27901 44567 27935 44581
rect 27901 44547 27935 44567
rect 27901 44499 27935 44509
rect 27901 44475 27935 44499
rect 27901 44431 27935 44437
rect 27901 44403 27935 44431
rect 27901 44363 27935 44365
rect 27901 44331 27935 44363
rect 27901 44261 27935 44293
rect 27901 44259 27935 44261
rect 27901 44193 27935 44221
rect 27901 44187 27935 44193
rect 27901 44125 27935 44149
rect 27901 44115 27935 44125
rect 27901 44057 27935 44077
rect 27901 44043 27935 44057
rect 27901 43989 27935 44005
rect 27901 43971 27935 43989
rect 27901 43921 27935 43933
rect 27901 43899 27935 43921
rect 27901 43853 27935 43861
rect 27901 43827 27935 43853
rect 27901 43785 27935 43789
rect 27901 43755 27935 43785
rect 27901 43683 27935 43717
rect 28359 44907 28393 44941
rect 28359 44839 28393 44869
rect 28359 44835 28393 44839
rect 28359 44771 28393 44797
rect 28359 44763 28393 44771
rect 28359 44703 28393 44725
rect 28359 44691 28393 44703
rect 28359 44635 28393 44653
rect 28359 44619 28393 44635
rect 28359 44567 28393 44581
rect 28359 44547 28393 44567
rect 28359 44499 28393 44509
rect 28359 44475 28393 44499
rect 28359 44431 28393 44437
rect 28359 44403 28393 44431
rect 28359 44363 28393 44365
rect 28359 44331 28393 44363
rect 28359 44261 28393 44293
rect 28359 44259 28393 44261
rect 28359 44193 28393 44221
rect 28359 44187 28393 44193
rect 28359 44125 28393 44149
rect 28359 44115 28393 44125
rect 28359 44057 28393 44077
rect 28359 44043 28393 44057
rect 28359 43989 28393 44005
rect 28359 43971 28393 43989
rect 28359 43921 28393 43933
rect 28359 43899 28393 43921
rect 28359 43853 28393 43861
rect 28359 43827 28393 43853
rect 28359 43785 28393 43789
rect 28359 43755 28393 43785
rect 28359 43683 28393 43717
rect 28817 44907 28851 44941
rect 28817 44839 28851 44869
rect 28817 44835 28851 44839
rect 28817 44771 28851 44797
rect 28817 44763 28851 44771
rect 28817 44703 28851 44725
rect 28817 44691 28851 44703
rect 28817 44635 28851 44653
rect 28817 44619 28851 44635
rect 28817 44567 28851 44581
rect 28817 44547 28851 44567
rect 28817 44499 28851 44509
rect 28817 44475 28851 44499
rect 28817 44431 28851 44437
rect 28817 44403 28851 44431
rect 28817 44363 28851 44365
rect 28817 44331 28851 44363
rect 28817 44261 28851 44293
rect 28817 44259 28851 44261
rect 28817 44193 28851 44221
rect 28817 44187 28851 44193
rect 28817 44125 28851 44149
rect 28817 44115 28851 44125
rect 28817 44057 28851 44077
rect 28817 44043 28851 44057
rect 28817 43989 28851 44005
rect 28817 43971 28851 43989
rect 28817 43921 28851 43933
rect 28817 43899 28851 43921
rect 28817 43853 28851 43861
rect 28817 43827 28851 43853
rect 28817 43785 28851 43789
rect 28817 43755 28851 43785
rect 28817 43683 28851 43717
rect 29275 44907 29309 44941
rect 29275 44839 29309 44869
rect 29275 44835 29309 44839
rect 29275 44771 29309 44797
rect 29275 44763 29309 44771
rect 29275 44703 29309 44725
rect 29275 44691 29309 44703
rect 29275 44635 29309 44653
rect 29275 44619 29309 44635
rect 29275 44567 29309 44581
rect 29275 44547 29309 44567
rect 29275 44499 29309 44509
rect 29275 44475 29309 44499
rect 29275 44431 29309 44437
rect 29275 44403 29309 44431
rect 29275 44363 29309 44365
rect 29275 44331 29309 44363
rect 29275 44261 29309 44293
rect 29275 44259 29309 44261
rect 29275 44193 29309 44221
rect 29275 44187 29309 44193
rect 29275 44125 29309 44149
rect 29275 44115 29309 44125
rect 29275 44057 29309 44077
rect 29275 44043 29309 44057
rect 29275 43989 29309 44005
rect 29275 43971 29309 43989
rect 29275 43921 29309 43933
rect 29275 43899 29309 43921
rect 29275 43853 29309 43861
rect 29275 43827 29309 43853
rect 29275 43785 29309 43789
rect 29275 43755 29309 43785
rect 29275 43683 29309 43717
rect 29733 44907 29767 44941
rect 29733 44839 29767 44869
rect 29733 44835 29767 44839
rect 29733 44771 29767 44797
rect 29733 44763 29767 44771
rect 29733 44703 29767 44725
rect 29733 44691 29767 44703
rect 29733 44635 29767 44653
rect 29733 44619 29767 44635
rect 29733 44567 29767 44581
rect 29733 44547 29767 44567
rect 29733 44499 29767 44509
rect 29733 44475 29767 44499
rect 29733 44431 29767 44437
rect 29733 44403 29767 44431
rect 29733 44363 29767 44365
rect 29733 44331 29767 44363
rect 29733 44261 29767 44293
rect 29733 44259 29767 44261
rect 29733 44193 29767 44221
rect 29733 44187 29767 44193
rect 29733 44125 29767 44149
rect 29733 44115 29767 44125
rect 29733 44057 29767 44077
rect 29733 44043 29767 44057
rect 29733 43989 29767 44005
rect 29733 43971 29767 43989
rect 29733 43921 29767 43933
rect 29733 43899 29767 43921
rect 29733 43853 29767 43861
rect 29733 43827 29767 43853
rect 29733 43785 29767 43789
rect 29733 43755 29767 43785
rect 29733 43683 29767 43717
rect 30191 44907 30225 44941
rect 30191 44839 30225 44869
rect 30191 44835 30225 44839
rect 30191 44771 30225 44797
rect 30191 44763 30225 44771
rect 30191 44703 30225 44725
rect 30191 44691 30225 44703
rect 30191 44635 30225 44653
rect 30191 44619 30225 44635
rect 30191 44567 30225 44581
rect 30191 44547 30225 44567
rect 30191 44499 30225 44509
rect 30191 44475 30225 44499
rect 30191 44431 30225 44437
rect 30191 44403 30225 44431
rect 30191 44363 30225 44365
rect 30191 44331 30225 44363
rect 30191 44261 30225 44293
rect 30191 44259 30225 44261
rect 30191 44193 30225 44221
rect 30191 44187 30225 44193
rect 30191 44125 30225 44149
rect 30191 44115 30225 44125
rect 30191 44057 30225 44077
rect 30191 44043 30225 44057
rect 30191 43989 30225 44005
rect 30191 43971 30225 43989
rect 30191 43921 30225 43933
rect 30191 43899 30225 43921
rect 30191 43853 30225 43861
rect 30191 43827 30225 43853
rect 30191 43785 30225 43789
rect 30191 43755 30225 43785
rect 30191 43683 30225 43717
rect 30649 44907 30683 44941
rect 30649 44839 30683 44869
rect 30649 44835 30683 44839
rect 30649 44771 30683 44797
rect 30649 44763 30683 44771
rect 30649 44703 30683 44725
rect 30649 44691 30683 44703
rect 30649 44635 30683 44653
rect 30649 44619 30683 44635
rect 30649 44567 30683 44581
rect 30649 44547 30683 44567
rect 30649 44499 30683 44509
rect 30649 44475 30683 44499
rect 30649 44431 30683 44437
rect 30649 44403 30683 44431
rect 30649 44363 30683 44365
rect 30649 44331 30683 44363
rect 30649 44261 30683 44293
rect 30649 44259 30683 44261
rect 30649 44193 30683 44221
rect 30649 44187 30683 44193
rect 30649 44125 30683 44149
rect 30649 44115 30683 44125
rect 30649 44057 30683 44077
rect 30649 44043 30683 44057
rect 30649 43989 30683 44005
rect 30649 43971 30683 43989
rect 30649 43921 30683 43933
rect 30649 43899 30683 43921
rect 30649 43853 30683 43861
rect 30649 43827 30683 43853
rect 30649 43785 30683 43789
rect 30649 43755 30683 43785
rect 30649 43683 30683 43717
rect 31107 44907 31141 44941
rect 31107 44839 31141 44869
rect 31107 44835 31141 44839
rect 31107 44771 31141 44797
rect 31107 44763 31141 44771
rect 31107 44703 31141 44725
rect 31107 44691 31141 44703
rect 31107 44635 31141 44653
rect 31107 44619 31141 44635
rect 31107 44567 31141 44581
rect 31107 44547 31141 44567
rect 31107 44499 31141 44509
rect 31107 44475 31141 44499
rect 31107 44431 31141 44437
rect 31107 44403 31141 44431
rect 31107 44363 31141 44365
rect 31107 44331 31141 44363
rect 31107 44261 31141 44293
rect 31107 44259 31141 44261
rect 31107 44193 31141 44221
rect 31107 44187 31141 44193
rect 31107 44125 31141 44149
rect 31107 44115 31141 44125
rect 31107 44057 31141 44077
rect 31107 44043 31141 44057
rect 31107 43989 31141 44005
rect 31107 43971 31141 43989
rect 31107 43921 31141 43933
rect 31107 43899 31141 43921
rect 31107 43853 31141 43861
rect 31107 43827 31141 43853
rect 31107 43785 31141 43789
rect 31107 43755 31141 43785
rect 31107 43683 31141 43717
rect 31565 44907 31599 44941
rect 31565 44839 31599 44869
rect 31565 44835 31599 44839
rect 31565 44771 31599 44797
rect 31565 44763 31599 44771
rect 31565 44703 31599 44725
rect 31565 44691 31599 44703
rect 31565 44635 31599 44653
rect 31565 44619 31599 44635
rect 31565 44567 31599 44581
rect 31565 44547 31599 44567
rect 31565 44499 31599 44509
rect 31565 44475 31599 44499
rect 31565 44431 31599 44437
rect 31565 44403 31599 44431
rect 31565 44363 31599 44365
rect 31565 44331 31599 44363
rect 31565 44261 31599 44293
rect 31565 44259 31599 44261
rect 31565 44193 31599 44221
rect 31565 44187 31599 44193
rect 31565 44125 31599 44149
rect 31565 44115 31599 44125
rect 31565 44057 31599 44077
rect 31565 44043 31599 44057
rect 31565 43989 31599 44005
rect 31565 43971 31599 43989
rect 31565 43921 31599 43933
rect 31565 43899 31599 43921
rect 31565 43853 31599 43861
rect 31565 43827 31599 43853
rect 31565 43785 31599 43789
rect 31565 43755 31599 43785
rect 31565 43683 31599 43717
rect 32023 44907 32057 44941
rect 32023 44839 32057 44869
rect 32023 44835 32057 44839
rect 32023 44771 32057 44797
rect 32023 44763 32057 44771
rect 32023 44703 32057 44725
rect 32023 44691 32057 44703
rect 32023 44635 32057 44653
rect 32023 44619 32057 44635
rect 32023 44567 32057 44581
rect 32023 44547 32057 44567
rect 32023 44499 32057 44509
rect 32023 44475 32057 44499
rect 32023 44431 32057 44437
rect 32023 44403 32057 44431
rect 32023 44363 32057 44365
rect 32023 44331 32057 44363
rect 32023 44261 32057 44293
rect 32023 44259 32057 44261
rect 32023 44193 32057 44221
rect 32023 44187 32057 44193
rect 32023 44125 32057 44149
rect 32023 44115 32057 44125
rect 32023 44057 32057 44077
rect 32023 44043 32057 44057
rect 32023 43989 32057 44005
rect 32023 43971 32057 43989
rect 32023 43921 32057 43933
rect 32023 43899 32057 43921
rect 32023 43853 32057 43861
rect 32023 43827 32057 43853
rect 32023 43785 32057 43789
rect 32023 43755 32057 43785
rect 32023 43683 32057 43717
rect 32481 44907 32515 44941
rect 32481 44839 32515 44869
rect 32481 44835 32515 44839
rect 32481 44771 32515 44797
rect 32481 44763 32515 44771
rect 32481 44703 32515 44725
rect 32481 44691 32515 44703
rect 32481 44635 32515 44653
rect 32481 44619 32515 44635
rect 32481 44567 32515 44581
rect 32481 44547 32515 44567
rect 32481 44499 32515 44509
rect 32481 44475 32515 44499
rect 32481 44431 32515 44437
rect 32481 44403 32515 44431
rect 32481 44363 32515 44365
rect 32481 44331 32515 44363
rect 32481 44261 32515 44293
rect 32481 44259 32515 44261
rect 32481 44193 32515 44221
rect 32481 44187 32515 44193
rect 32481 44125 32515 44149
rect 32481 44115 32515 44125
rect 32481 44057 32515 44077
rect 32481 44043 32515 44057
rect 32481 43989 32515 44005
rect 32481 43971 32515 43989
rect 32481 43921 32515 43933
rect 32481 43899 32515 43921
rect 32481 43853 32515 43861
rect 32481 43827 32515 43853
rect 32481 43785 32515 43789
rect 32481 43755 32515 43785
rect 32481 43683 32515 43717
rect 32939 44907 32973 44941
rect 32939 44839 32973 44869
rect 32939 44835 32973 44839
rect 32939 44771 32973 44797
rect 32939 44763 32973 44771
rect 32939 44703 32973 44725
rect 32939 44691 32973 44703
rect 32939 44635 32973 44653
rect 32939 44619 32973 44635
rect 32939 44567 32973 44581
rect 32939 44547 32973 44567
rect 32939 44499 32973 44509
rect 32939 44475 32973 44499
rect 32939 44431 32973 44437
rect 32939 44403 32973 44431
rect 32939 44363 32973 44365
rect 32939 44331 32973 44363
rect 32939 44261 32973 44293
rect 32939 44259 32973 44261
rect 32939 44193 32973 44221
rect 32939 44187 32973 44193
rect 32939 44125 32973 44149
rect 32939 44115 32973 44125
rect 32939 44057 32973 44077
rect 32939 44043 32973 44057
rect 32939 43989 32973 44005
rect 32939 43971 32973 43989
rect 32939 43921 32973 43933
rect 32939 43899 32973 43921
rect 32939 43853 32973 43861
rect 32939 43827 32973 43853
rect 32939 43785 32973 43789
rect 32939 43755 32973 43785
rect 32939 43683 32973 43717
rect 33397 44907 33431 44941
rect 33397 44839 33431 44869
rect 33397 44835 33431 44839
rect 33397 44771 33431 44797
rect 33397 44763 33431 44771
rect 33397 44703 33431 44725
rect 33397 44691 33431 44703
rect 33397 44635 33431 44653
rect 33397 44619 33431 44635
rect 33397 44567 33431 44581
rect 33397 44547 33431 44567
rect 33397 44499 33431 44509
rect 33397 44475 33431 44499
rect 33397 44431 33431 44437
rect 33397 44403 33431 44431
rect 33397 44363 33431 44365
rect 33397 44331 33431 44363
rect 33397 44261 33431 44293
rect 33397 44259 33431 44261
rect 33397 44193 33431 44221
rect 33397 44187 33431 44193
rect 33397 44125 33431 44149
rect 33397 44115 33431 44125
rect 33397 44057 33431 44077
rect 33397 44043 33431 44057
rect 33397 43989 33431 44005
rect 33397 43971 33431 43989
rect 33397 43921 33431 43933
rect 33397 43899 33431 43921
rect 33397 43853 33431 43861
rect 33397 43827 33431 43853
rect 33397 43785 33431 43789
rect 33397 43755 33431 43785
rect 33397 43683 33431 43717
rect 33855 44907 33889 44941
rect 33855 44839 33889 44869
rect 33855 44835 33889 44839
rect 33855 44771 33889 44797
rect 33855 44763 33889 44771
rect 33855 44703 33889 44725
rect 33855 44691 33889 44703
rect 33855 44635 33889 44653
rect 33855 44619 33889 44635
rect 33855 44567 33889 44581
rect 33855 44547 33889 44567
rect 33855 44499 33889 44509
rect 33855 44475 33889 44499
rect 33855 44431 33889 44437
rect 33855 44403 33889 44431
rect 33855 44363 33889 44365
rect 33855 44331 33889 44363
rect 33855 44261 33889 44293
rect 33855 44259 33889 44261
rect 33855 44193 33889 44221
rect 33855 44187 33889 44193
rect 33855 44125 33889 44149
rect 33855 44115 33889 44125
rect 33855 44057 33889 44077
rect 33855 44043 33889 44057
rect 33855 43989 33889 44005
rect 33855 43971 33889 43989
rect 33855 43921 33889 43933
rect 33855 43899 33889 43921
rect 33855 43853 33889 43861
rect 33855 43827 33889 43853
rect 33855 43785 33889 43789
rect 33855 43755 33889 43785
rect 33855 43683 33889 43717
rect 34313 44907 34347 44941
rect 34313 44839 34347 44869
rect 34313 44835 34347 44839
rect 34313 44771 34347 44797
rect 34313 44763 34347 44771
rect 34313 44703 34347 44725
rect 34313 44691 34347 44703
rect 34313 44635 34347 44653
rect 34313 44619 34347 44635
rect 34313 44567 34347 44581
rect 34313 44547 34347 44567
rect 34313 44499 34347 44509
rect 34313 44475 34347 44499
rect 34313 44431 34347 44437
rect 34313 44403 34347 44431
rect 34313 44363 34347 44365
rect 34313 44331 34347 44363
rect 34313 44261 34347 44293
rect 34313 44259 34347 44261
rect 34313 44193 34347 44221
rect 34313 44187 34347 44193
rect 34313 44125 34347 44149
rect 34313 44115 34347 44125
rect 34313 44057 34347 44077
rect 34313 44043 34347 44057
rect 34313 43989 34347 44005
rect 34313 43971 34347 43989
rect 34313 43921 34347 43933
rect 34313 43899 34347 43921
rect 34313 43853 34347 43861
rect 34313 43827 34347 43853
rect 34313 43785 34347 43789
rect 34313 43755 34347 43785
rect 34313 43683 34347 43717
rect 34771 44907 34805 44941
rect 34771 44839 34805 44869
rect 34771 44835 34805 44839
rect 34771 44771 34805 44797
rect 34771 44763 34805 44771
rect 34771 44703 34805 44725
rect 34771 44691 34805 44703
rect 34771 44635 34805 44653
rect 34771 44619 34805 44635
rect 34771 44567 34805 44581
rect 34771 44547 34805 44567
rect 34771 44499 34805 44509
rect 34771 44475 34805 44499
rect 34771 44431 34805 44437
rect 34771 44403 34805 44431
rect 34771 44363 34805 44365
rect 34771 44331 34805 44363
rect 34771 44261 34805 44293
rect 34771 44259 34805 44261
rect 34771 44193 34805 44221
rect 34771 44187 34805 44193
rect 34771 44125 34805 44149
rect 34771 44115 34805 44125
rect 34771 44057 34805 44077
rect 34771 44043 34805 44057
rect 34771 43989 34805 44005
rect 34771 43971 34805 43989
rect 34771 43921 34805 43933
rect 34771 43899 34805 43921
rect 34771 43853 34805 43861
rect 34771 43827 34805 43853
rect 34771 43785 34805 43789
rect 34771 43755 34805 43785
rect 34771 43683 34805 43717
rect 35229 44907 35263 44941
rect 35229 44839 35263 44869
rect 35229 44835 35263 44839
rect 35229 44771 35263 44797
rect 35229 44763 35263 44771
rect 35229 44703 35263 44725
rect 35229 44691 35263 44703
rect 35229 44635 35263 44653
rect 35229 44619 35263 44635
rect 35229 44567 35263 44581
rect 35229 44547 35263 44567
rect 35229 44499 35263 44509
rect 35229 44475 35263 44499
rect 35229 44431 35263 44437
rect 35229 44403 35263 44431
rect 35229 44363 35263 44365
rect 35229 44331 35263 44363
rect 35229 44261 35263 44293
rect 35229 44259 35263 44261
rect 35229 44193 35263 44221
rect 35229 44187 35263 44193
rect 35229 44125 35263 44149
rect 35229 44115 35263 44125
rect 35229 44057 35263 44077
rect 35229 44043 35263 44057
rect 35229 43989 35263 44005
rect 35229 43971 35263 43989
rect 35229 43921 35263 43933
rect 35229 43899 35263 43921
rect 35229 43853 35263 43861
rect 35229 43827 35263 43853
rect 35229 43785 35263 43789
rect 35229 43755 35263 43785
rect 35229 43683 35263 43717
rect 35687 44907 35721 44941
rect 35687 44839 35721 44869
rect 35687 44835 35721 44839
rect 35687 44771 35721 44797
rect 35687 44763 35721 44771
rect 35687 44703 35721 44725
rect 35687 44691 35721 44703
rect 35687 44635 35721 44653
rect 35687 44619 35721 44635
rect 35687 44567 35721 44581
rect 35687 44547 35721 44567
rect 35687 44499 35721 44509
rect 35687 44475 35721 44499
rect 35687 44431 35721 44437
rect 35687 44403 35721 44431
rect 35687 44363 35721 44365
rect 35687 44331 35721 44363
rect 35687 44261 35721 44293
rect 35687 44259 35721 44261
rect 35687 44193 35721 44221
rect 35687 44187 35721 44193
rect 35687 44125 35721 44149
rect 35687 44115 35721 44125
rect 35687 44057 35721 44077
rect 35687 44043 35721 44057
rect 35687 43989 35721 44005
rect 35687 43971 35721 43989
rect 35687 43921 35721 43933
rect 35687 43899 35721 43921
rect 35687 43853 35721 43861
rect 35687 43827 35721 43853
rect 35687 43785 35721 43789
rect 35687 43755 35721 43785
rect 35687 43683 35721 43717
rect 36145 44907 36179 44941
rect 36145 44839 36179 44869
rect 36145 44835 36179 44839
rect 36145 44771 36179 44797
rect 36145 44763 36179 44771
rect 36145 44703 36179 44725
rect 36145 44691 36179 44703
rect 36145 44635 36179 44653
rect 36145 44619 36179 44635
rect 36145 44567 36179 44581
rect 36145 44547 36179 44567
rect 36145 44499 36179 44509
rect 36145 44475 36179 44499
rect 36145 44431 36179 44437
rect 36145 44403 36179 44431
rect 36145 44363 36179 44365
rect 36145 44331 36179 44363
rect 36145 44261 36179 44293
rect 36145 44259 36179 44261
rect 36145 44193 36179 44221
rect 36145 44187 36179 44193
rect 36145 44125 36179 44149
rect 36145 44115 36179 44125
rect 36145 44057 36179 44077
rect 36145 44043 36179 44057
rect 36145 43989 36179 44005
rect 36145 43971 36179 43989
rect 36145 43921 36179 43933
rect 36145 43899 36179 43921
rect 36145 43853 36179 43861
rect 36145 43827 36179 43853
rect 36145 43785 36179 43789
rect 36145 43755 36179 43785
rect 36145 43683 36179 43717
rect 36603 44907 36637 44941
rect 36603 44839 36637 44869
rect 36603 44835 36637 44839
rect 36603 44771 36637 44797
rect 36603 44763 36637 44771
rect 36603 44703 36637 44725
rect 36603 44691 36637 44703
rect 36603 44635 36637 44653
rect 36603 44619 36637 44635
rect 36603 44567 36637 44581
rect 36603 44547 36637 44567
rect 36603 44499 36637 44509
rect 36603 44475 36637 44499
rect 36603 44431 36637 44437
rect 36603 44403 36637 44431
rect 36603 44363 36637 44365
rect 36603 44331 36637 44363
rect 36603 44261 36637 44293
rect 36603 44259 36637 44261
rect 36603 44193 36637 44221
rect 36603 44187 36637 44193
rect 36603 44125 36637 44149
rect 36603 44115 36637 44125
rect 36603 44057 36637 44077
rect 36603 44043 36637 44057
rect 36603 43989 36637 44005
rect 36603 43971 36637 43989
rect 36603 43921 36637 43933
rect 36603 43899 36637 43921
rect 36603 43853 36637 43861
rect 36603 43827 36637 43853
rect 36603 43785 36637 43789
rect 36603 43755 36637 43785
rect 36603 43683 36637 43717
rect 37061 44907 37095 44941
rect 37061 44839 37095 44869
rect 37061 44835 37095 44839
rect 37061 44771 37095 44797
rect 37061 44763 37095 44771
rect 37061 44703 37095 44725
rect 37061 44691 37095 44703
rect 37061 44635 37095 44653
rect 37061 44619 37095 44635
rect 37061 44567 37095 44581
rect 37061 44547 37095 44567
rect 37061 44499 37095 44509
rect 37061 44475 37095 44499
rect 37061 44431 37095 44437
rect 37061 44403 37095 44431
rect 37061 44363 37095 44365
rect 37061 44331 37095 44363
rect 37061 44261 37095 44293
rect 37061 44259 37095 44261
rect 37061 44193 37095 44221
rect 37061 44187 37095 44193
rect 37061 44125 37095 44149
rect 37061 44115 37095 44125
rect 37061 44057 37095 44077
rect 37061 44043 37095 44057
rect 37061 43989 37095 44005
rect 37061 43971 37095 43989
rect 37061 43921 37095 43933
rect 37061 43899 37095 43921
rect 37061 43853 37095 43861
rect 37061 43827 37095 43853
rect 37061 43785 37095 43789
rect 37061 43755 37095 43785
rect 37061 43683 37095 43717
rect 37519 44907 37553 44941
rect 37519 44839 37553 44869
rect 37519 44835 37553 44839
rect 37519 44771 37553 44797
rect 37519 44763 37553 44771
rect 37519 44703 37553 44725
rect 37519 44691 37553 44703
rect 37519 44635 37553 44653
rect 37519 44619 37553 44635
rect 37519 44567 37553 44581
rect 37519 44547 37553 44567
rect 37519 44499 37553 44509
rect 37519 44475 37553 44499
rect 37519 44431 37553 44437
rect 37519 44403 37553 44431
rect 37519 44363 37553 44365
rect 37519 44331 37553 44363
rect 37519 44261 37553 44293
rect 37519 44259 37553 44261
rect 37519 44193 37553 44221
rect 37519 44187 37553 44193
rect 37519 44125 37553 44149
rect 37519 44115 37553 44125
rect 37519 44057 37553 44077
rect 37519 44043 37553 44057
rect 37519 43989 37553 44005
rect 37519 43971 37553 43989
rect 37519 43921 37553 43933
rect 37519 43899 37553 43921
rect 37519 43853 37553 43861
rect 37519 43827 37553 43853
rect 37519 43785 37553 43789
rect 37519 43755 37553 43785
rect 37519 43683 37553 43717
rect 37977 44907 38011 44941
rect 37977 44839 38011 44869
rect 37977 44835 38011 44839
rect 37977 44771 38011 44797
rect 37977 44763 38011 44771
rect 37977 44703 38011 44725
rect 37977 44691 38011 44703
rect 37977 44635 38011 44653
rect 37977 44619 38011 44635
rect 37977 44567 38011 44581
rect 37977 44547 38011 44567
rect 37977 44499 38011 44509
rect 37977 44475 38011 44499
rect 37977 44431 38011 44437
rect 37977 44403 38011 44431
rect 37977 44363 38011 44365
rect 37977 44331 38011 44363
rect 37977 44261 38011 44293
rect 37977 44259 38011 44261
rect 37977 44193 38011 44221
rect 37977 44187 38011 44193
rect 37977 44125 38011 44149
rect 37977 44115 38011 44125
rect 37977 44057 38011 44077
rect 37977 44043 38011 44057
rect 37977 43989 38011 44005
rect 37977 43971 38011 43989
rect 37977 43921 38011 43933
rect 37977 43899 38011 43921
rect 37977 43853 38011 43861
rect 37977 43827 38011 43853
rect 37977 43785 38011 43789
rect 37977 43755 38011 43785
rect 37977 43683 38011 43717
rect 38435 44907 38469 44941
rect 38435 44839 38469 44869
rect 38435 44835 38469 44839
rect 38435 44771 38469 44797
rect 38435 44763 38469 44771
rect 38435 44703 38469 44725
rect 38435 44691 38469 44703
rect 38435 44635 38469 44653
rect 38435 44619 38469 44635
rect 38435 44567 38469 44581
rect 38435 44547 38469 44567
rect 38435 44499 38469 44509
rect 38435 44475 38469 44499
rect 38435 44431 38469 44437
rect 38435 44403 38469 44431
rect 38435 44363 38469 44365
rect 38435 44331 38469 44363
rect 38435 44261 38469 44293
rect 38435 44259 38469 44261
rect 38435 44193 38469 44221
rect 38435 44187 38469 44193
rect 38435 44125 38469 44149
rect 38435 44115 38469 44125
rect 38435 44057 38469 44077
rect 38435 44043 38469 44057
rect 38435 43989 38469 44005
rect 38435 43971 38469 43989
rect 38435 43921 38469 43933
rect 38435 43899 38469 43921
rect 38435 43853 38469 43861
rect 38435 43827 38469 43853
rect 38435 43785 38469 43789
rect 38435 43755 38469 43785
rect 38435 43683 38469 43717
rect 38893 44907 38927 44941
rect 38893 44839 38927 44869
rect 38893 44835 38927 44839
rect 38893 44771 38927 44797
rect 38893 44763 38927 44771
rect 38893 44703 38927 44725
rect 38893 44691 38927 44703
rect 38893 44635 38927 44653
rect 38893 44619 38927 44635
rect 38893 44567 38927 44581
rect 38893 44547 38927 44567
rect 38893 44499 38927 44509
rect 38893 44475 38927 44499
rect 38893 44431 38927 44437
rect 38893 44403 38927 44431
rect 38893 44363 38927 44365
rect 38893 44331 38927 44363
rect 38893 44261 38927 44293
rect 38893 44259 38927 44261
rect 38893 44193 38927 44221
rect 38893 44187 38927 44193
rect 38893 44125 38927 44149
rect 38893 44115 38927 44125
rect 38893 44057 38927 44077
rect 38893 44043 38927 44057
rect 38893 43989 38927 44005
rect 38893 43971 38927 43989
rect 38893 43921 38927 43933
rect 38893 43899 38927 43921
rect 38893 43853 38927 43861
rect 38893 43827 38927 43853
rect 38893 43785 38927 43789
rect 38893 43755 38927 43785
rect 38893 43683 38927 43717
rect 39351 44907 39385 44941
rect 39351 44839 39385 44869
rect 39351 44835 39385 44839
rect 39351 44771 39385 44797
rect 39351 44763 39385 44771
rect 39351 44703 39385 44725
rect 39351 44691 39385 44703
rect 39351 44635 39385 44653
rect 39351 44619 39385 44635
rect 39351 44567 39385 44581
rect 39351 44547 39385 44567
rect 39351 44499 39385 44509
rect 39351 44475 39385 44499
rect 39351 44431 39385 44437
rect 39351 44403 39385 44431
rect 39351 44363 39385 44365
rect 39351 44331 39385 44363
rect 39351 44261 39385 44293
rect 39351 44259 39385 44261
rect 39351 44193 39385 44221
rect 39351 44187 39385 44193
rect 39351 44125 39385 44149
rect 39351 44115 39385 44125
rect 39351 44057 39385 44077
rect 39351 44043 39385 44057
rect 39351 43989 39385 44005
rect 39351 43971 39385 43989
rect 39351 43921 39385 43933
rect 39351 43899 39385 43921
rect 39351 43853 39385 43861
rect 39351 43827 39385 43853
rect 39351 43785 39385 43789
rect 39351 43755 39385 43785
rect 39351 43683 39385 43717
rect 39809 44907 39843 44941
rect 39809 44839 39843 44869
rect 39809 44835 39843 44839
rect 39809 44771 39843 44797
rect 39809 44763 39843 44771
rect 39809 44703 39843 44725
rect 39809 44691 39843 44703
rect 39809 44635 39843 44653
rect 39809 44619 39843 44635
rect 39809 44567 39843 44581
rect 39809 44547 39843 44567
rect 39809 44499 39843 44509
rect 39809 44475 39843 44499
rect 39809 44431 39843 44437
rect 39809 44403 39843 44431
rect 39809 44363 39843 44365
rect 39809 44331 39843 44363
rect 39809 44261 39843 44293
rect 39809 44259 39843 44261
rect 39809 44193 39843 44221
rect 39809 44187 39843 44193
rect 39809 44125 39843 44149
rect 39809 44115 39843 44125
rect 39809 44057 39843 44077
rect 39809 44043 39843 44057
rect 39809 43989 39843 44005
rect 39809 43971 39843 43989
rect 39809 43921 39843 43933
rect 39809 43899 39843 43921
rect 39809 43853 39843 43861
rect 39809 43827 39843 43853
rect 39809 43785 39843 43789
rect 39809 43755 39843 43785
rect 39809 43683 39843 43717
rect 40267 44907 40301 44941
rect 40267 44839 40301 44869
rect 40267 44835 40301 44839
rect 40267 44771 40301 44797
rect 40267 44763 40301 44771
rect 40267 44703 40301 44725
rect 40267 44691 40301 44703
rect 40267 44635 40301 44653
rect 40267 44619 40301 44635
rect 40267 44567 40301 44581
rect 40267 44547 40301 44567
rect 40267 44499 40301 44509
rect 40267 44475 40301 44499
rect 40267 44431 40301 44437
rect 40267 44403 40301 44431
rect 40267 44363 40301 44365
rect 40267 44331 40301 44363
rect 40267 44261 40301 44293
rect 40267 44259 40301 44261
rect 40267 44193 40301 44221
rect 40267 44187 40301 44193
rect 40267 44125 40301 44149
rect 40267 44115 40301 44125
rect 40267 44057 40301 44077
rect 40267 44043 40301 44057
rect 40267 43989 40301 44005
rect 40267 43971 40301 43989
rect 40267 43921 40301 43933
rect 40267 43899 40301 43921
rect 40267 43853 40301 43861
rect 40267 43827 40301 43853
rect 40267 43785 40301 43789
rect 40267 43755 40301 43785
rect 40267 43683 40301 43717
rect 40725 44907 40759 44941
rect 40725 44839 40759 44869
rect 40725 44835 40759 44839
rect 40725 44771 40759 44797
rect 40725 44763 40759 44771
rect 40725 44703 40759 44725
rect 40725 44691 40759 44703
rect 40725 44635 40759 44653
rect 40725 44619 40759 44635
rect 40725 44567 40759 44581
rect 40725 44547 40759 44567
rect 40725 44499 40759 44509
rect 40725 44475 40759 44499
rect 40725 44431 40759 44437
rect 40725 44403 40759 44431
rect 40725 44363 40759 44365
rect 40725 44331 40759 44363
rect 40725 44261 40759 44293
rect 40725 44259 40759 44261
rect 40725 44193 40759 44221
rect 40725 44187 40759 44193
rect 40725 44125 40759 44149
rect 40725 44115 40759 44125
rect 40725 44057 40759 44077
rect 40725 44043 40759 44057
rect 40725 43989 40759 44005
rect 40725 43971 40759 43989
rect 40725 43921 40759 43933
rect 40725 43899 40759 43921
rect 40725 43853 40759 43861
rect 40725 43827 40759 43853
rect 40725 43785 40759 43789
rect 40725 43755 40759 43785
rect 40725 43683 40759 43717
rect 41183 44907 41217 44941
rect 41183 44839 41217 44869
rect 41183 44835 41217 44839
rect 41183 44771 41217 44797
rect 41183 44763 41217 44771
rect 41183 44703 41217 44725
rect 41183 44691 41217 44703
rect 41183 44635 41217 44653
rect 41183 44619 41217 44635
rect 41183 44567 41217 44581
rect 41183 44547 41217 44567
rect 41183 44499 41217 44509
rect 41183 44475 41217 44499
rect 41183 44431 41217 44437
rect 41183 44403 41217 44431
rect 41183 44363 41217 44365
rect 41183 44331 41217 44363
rect 41183 44261 41217 44293
rect 41183 44259 41217 44261
rect 41183 44193 41217 44221
rect 41183 44187 41217 44193
rect 41183 44125 41217 44149
rect 41183 44115 41217 44125
rect 41183 44057 41217 44077
rect 41183 44043 41217 44057
rect 41183 43989 41217 44005
rect 41183 43971 41217 43989
rect 41183 43921 41217 43933
rect 41183 43899 41217 43921
rect 41183 43853 41217 43861
rect 41183 43827 41217 43853
rect 41183 43785 41217 43789
rect 41183 43755 41217 43785
rect 41183 43683 41217 43717
rect 41641 44907 41675 44941
rect 41641 44839 41675 44869
rect 41641 44835 41675 44839
rect 41641 44771 41675 44797
rect 41641 44763 41675 44771
rect 41641 44703 41675 44725
rect 41641 44691 41675 44703
rect 41641 44635 41675 44653
rect 41641 44619 41675 44635
rect 41641 44567 41675 44581
rect 41641 44547 41675 44567
rect 41641 44499 41675 44509
rect 41641 44475 41675 44499
rect 41641 44431 41675 44437
rect 41641 44403 41675 44431
rect 41641 44363 41675 44365
rect 41641 44331 41675 44363
rect 41641 44261 41675 44293
rect 41641 44259 41675 44261
rect 41641 44193 41675 44221
rect 41641 44187 41675 44193
rect 41641 44125 41675 44149
rect 41641 44115 41675 44125
rect 41641 44057 41675 44077
rect 41641 44043 41675 44057
rect 41641 43989 41675 44005
rect 41641 43971 41675 43989
rect 41641 43921 41675 43933
rect 41641 43899 41675 43921
rect 41641 43853 41675 43861
rect 41641 43827 41675 43853
rect 41641 43785 41675 43789
rect 41641 43755 41675 43785
rect 41641 43683 41675 43717
rect 42099 44907 42133 44941
rect 42099 44839 42133 44869
rect 42099 44835 42133 44839
rect 42099 44771 42133 44797
rect 42099 44763 42133 44771
rect 42099 44703 42133 44725
rect 42099 44691 42133 44703
rect 42099 44635 42133 44653
rect 42099 44619 42133 44635
rect 42099 44567 42133 44581
rect 42099 44547 42133 44567
rect 42099 44499 42133 44509
rect 42099 44475 42133 44499
rect 42099 44431 42133 44437
rect 42099 44403 42133 44431
rect 42099 44363 42133 44365
rect 42099 44331 42133 44363
rect 42099 44261 42133 44293
rect 42099 44259 42133 44261
rect 42099 44193 42133 44221
rect 42099 44187 42133 44193
rect 42099 44125 42133 44149
rect 42099 44115 42133 44125
rect 42099 44057 42133 44077
rect 42099 44043 42133 44057
rect 42099 43989 42133 44005
rect 42099 43971 42133 43989
rect 42099 43921 42133 43933
rect 42099 43899 42133 43921
rect 42099 43853 42133 43861
rect 42099 43827 42133 43853
rect 42099 43785 42133 43789
rect 42099 43755 42133 43785
rect 42099 43683 42133 43717
rect 42557 44907 42591 44941
rect 42557 44839 42591 44869
rect 42557 44835 42591 44839
rect 42557 44771 42591 44797
rect 42557 44763 42591 44771
rect 42557 44703 42591 44725
rect 42557 44691 42591 44703
rect 42557 44635 42591 44653
rect 42557 44619 42591 44635
rect 42557 44567 42591 44581
rect 42557 44547 42591 44567
rect 42557 44499 42591 44509
rect 42557 44475 42591 44499
rect 42557 44431 42591 44437
rect 42557 44403 42591 44431
rect 42557 44363 42591 44365
rect 42557 44331 42591 44363
rect 42557 44261 42591 44293
rect 42557 44259 42591 44261
rect 42557 44193 42591 44221
rect 42557 44187 42591 44193
rect 42557 44125 42591 44149
rect 42557 44115 42591 44125
rect 42557 44057 42591 44077
rect 42557 44043 42591 44057
rect 42557 43989 42591 44005
rect 42557 43971 42591 43989
rect 42557 43921 42591 43933
rect 42557 43899 42591 43921
rect 42557 43853 42591 43861
rect 42557 43827 42591 43853
rect 42557 43785 42591 43789
rect 42557 43755 42591 43785
rect 42557 43683 42591 43717
rect 43006 44842 43040 44876
rect 43096 44861 43130 44876
rect 43186 44861 43220 44876
rect 43276 44861 43310 44876
rect 43366 44861 43400 44876
rect 43456 44861 43490 44876
rect 43546 44861 43580 44876
rect 43636 44861 43670 44876
rect 43726 44861 43760 44876
rect 43816 44861 43850 44876
rect 43906 44861 43940 44876
rect 43996 44861 44030 44876
rect 44086 44861 44120 44876
rect 43096 44842 43116 44861
rect 43116 44842 43130 44861
rect 43186 44842 43206 44861
rect 43206 44842 43220 44861
rect 43276 44842 43296 44861
rect 43296 44842 43310 44861
rect 43366 44842 43386 44861
rect 43386 44842 43400 44861
rect 43456 44842 43476 44861
rect 43476 44842 43490 44861
rect 43546 44842 43566 44861
rect 43566 44842 43580 44861
rect 43636 44842 43656 44861
rect 43656 44842 43670 44861
rect 43726 44842 43746 44861
rect 43746 44842 43760 44861
rect 43816 44842 43836 44861
rect 43836 44842 43850 44861
rect 43906 44842 43926 44861
rect 43926 44842 43940 44861
rect 43996 44842 44016 44861
rect 44016 44842 44030 44861
rect 44086 44842 44106 44861
rect 44106 44842 44120 44861
rect 44176 44842 44210 44876
rect 44346 44842 44380 44876
rect 44436 44861 44470 44876
rect 44526 44861 44560 44876
rect 44616 44861 44650 44876
rect 44706 44861 44740 44876
rect 44796 44861 44830 44876
rect 44886 44861 44920 44876
rect 44976 44861 45010 44876
rect 45066 44861 45100 44876
rect 45156 44861 45190 44876
rect 45246 44861 45280 44876
rect 45336 44861 45370 44876
rect 45426 44861 45460 44876
rect 44436 44842 44456 44861
rect 44456 44842 44470 44861
rect 44526 44842 44546 44861
rect 44546 44842 44560 44861
rect 44616 44842 44636 44861
rect 44636 44842 44650 44861
rect 44706 44842 44726 44861
rect 44726 44842 44740 44861
rect 44796 44842 44816 44861
rect 44816 44842 44830 44861
rect 44886 44842 44906 44861
rect 44906 44842 44920 44861
rect 44976 44842 44996 44861
rect 44996 44842 45010 44861
rect 45066 44842 45086 44861
rect 45086 44842 45100 44861
rect 45156 44842 45176 44861
rect 45176 44842 45190 44861
rect 45246 44842 45266 44861
rect 45266 44842 45280 44861
rect 45336 44842 45356 44861
rect 45356 44842 45370 44861
rect 45426 44842 45446 44861
rect 45446 44842 45460 44861
rect 45516 44842 45550 44876
rect 45686 44842 45720 44876
rect 45776 44861 45810 44876
rect 45866 44861 45900 44876
rect 45956 44861 45990 44876
rect 46046 44861 46080 44876
rect 46136 44861 46170 44876
rect 46226 44861 46260 44876
rect 46316 44861 46350 44876
rect 46406 44861 46440 44876
rect 46496 44861 46530 44876
rect 46586 44861 46620 44876
rect 46676 44861 46710 44876
rect 46766 44861 46800 44876
rect 45776 44842 45796 44861
rect 45796 44842 45810 44861
rect 45866 44842 45886 44861
rect 45886 44842 45900 44861
rect 45956 44842 45976 44861
rect 45976 44842 45990 44861
rect 46046 44842 46066 44861
rect 46066 44842 46080 44861
rect 46136 44842 46156 44861
rect 46156 44842 46170 44861
rect 46226 44842 46246 44861
rect 46246 44842 46260 44861
rect 46316 44842 46336 44861
rect 46336 44842 46350 44861
rect 46406 44842 46426 44861
rect 46426 44842 46440 44861
rect 46496 44842 46516 44861
rect 46516 44842 46530 44861
rect 46586 44842 46606 44861
rect 46606 44842 46620 44861
rect 46676 44842 46696 44861
rect 46696 44842 46710 44861
rect 46766 44842 46786 44861
rect 46786 44842 46800 44861
rect 46856 44842 46890 44876
rect 47026 44842 47060 44876
rect 47116 44861 47150 44876
rect 47206 44861 47240 44876
rect 47296 44861 47330 44876
rect 47386 44861 47420 44876
rect 47476 44861 47510 44876
rect 47566 44861 47600 44876
rect 47656 44861 47690 44876
rect 47746 44861 47780 44876
rect 47836 44861 47870 44876
rect 47926 44861 47960 44876
rect 48016 44861 48050 44876
rect 48106 44861 48140 44876
rect 47116 44842 47136 44861
rect 47136 44842 47150 44861
rect 47206 44842 47226 44861
rect 47226 44842 47240 44861
rect 47296 44842 47316 44861
rect 47316 44842 47330 44861
rect 47386 44842 47406 44861
rect 47406 44842 47420 44861
rect 47476 44842 47496 44861
rect 47496 44842 47510 44861
rect 47566 44842 47586 44861
rect 47586 44842 47600 44861
rect 47656 44842 47676 44861
rect 47676 44842 47690 44861
rect 47746 44842 47766 44861
rect 47766 44842 47780 44861
rect 47836 44842 47856 44861
rect 47856 44842 47870 44861
rect 47926 44842 47946 44861
rect 47946 44842 47960 44861
rect 48016 44842 48036 44861
rect 48036 44842 48050 44861
rect 48106 44842 48126 44861
rect 48126 44842 48140 44861
rect 48196 44842 48230 44876
rect 48366 44842 48400 44876
rect 48456 44861 48490 44876
rect 48546 44861 48580 44876
rect 48636 44861 48670 44876
rect 48726 44861 48760 44876
rect 48816 44861 48850 44876
rect 48906 44861 48940 44876
rect 48996 44861 49030 44876
rect 49086 44861 49120 44876
rect 49176 44861 49210 44876
rect 49266 44861 49300 44876
rect 49356 44861 49390 44876
rect 49446 44861 49480 44876
rect 48456 44842 48476 44861
rect 48476 44842 48490 44861
rect 48546 44842 48566 44861
rect 48566 44842 48580 44861
rect 48636 44842 48656 44861
rect 48656 44842 48670 44861
rect 48726 44842 48746 44861
rect 48746 44842 48760 44861
rect 48816 44842 48836 44861
rect 48836 44842 48850 44861
rect 48906 44842 48926 44861
rect 48926 44842 48940 44861
rect 48996 44842 49016 44861
rect 49016 44842 49030 44861
rect 49086 44842 49106 44861
rect 49106 44842 49120 44861
rect 49176 44842 49196 44861
rect 49196 44842 49210 44861
rect 49266 44842 49286 44861
rect 49286 44842 49300 44861
rect 49356 44842 49376 44861
rect 49376 44842 49390 44861
rect 49446 44842 49466 44861
rect 49466 44842 49480 44861
rect 49536 44842 49570 44876
rect 49706 44842 49740 44876
rect 49796 44861 49830 44876
rect 49886 44861 49920 44876
rect 49976 44861 50010 44876
rect 50066 44861 50100 44876
rect 50156 44861 50190 44876
rect 50246 44861 50280 44876
rect 50336 44861 50370 44876
rect 50426 44861 50460 44876
rect 50516 44861 50550 44876
rect 50606 44861 50640 44876
rect 50696 44861 50730 44876
rect 50786 44861 50820 44876
rect 49796 44842 49816 44861
rect 49816 44842 49830 44861
rect 49886 44842 49906 44861
rect 49906 44842 49920 44861
rect 49976 44842 49996 44861
rect 49996 44842 50010 44861
rect 50066 44842 50086 44861
rect 50086 44842 50100 44861
rect 50156 44842 50176 44861
rect 50176 44842 50190 44861
rect 50246 44842 50266 44861
rect 50266 44842 50280 44861
rect 50336 44842 50356 44861
rect 50356 44842 50370 44861
rect 50426 44842 50446 44861
rect 50446 44842 50460 44861
rect 50516 44842 50536 44861
rect 50536 44842 50550 44861
rect 50606 44842 50626 44861
rect 50626 44842 50640 44861
rect 50696 44842 50716 44861
rect 50716 44842 50730 44861
rect 50786 44842 50806 44861
rect 50806 44842 50820 44861
rect 50876 44842 50910 44876
rect 51046 44842 51080 44876
rect 51136 44861 51170 44876
rect 51226 44861 51260 44876
rect 51316 44861 51350 44876
rect 51406 44861 51440 44876
rect 51496 44861 51530 44876
rect 51586 44861 51620 44876
rect 51676 44861 51710 44876
rect 51766 44861 51800 44876
rect 51856 44861 51890 44876
rect 51946 44861 51980 44876
rect 52036 44861 52070 44876
rect 52126 44861 52160 44876
rect 51136 44842 51156 44861
rect 51156 44842 51170 44861
rect 51226 44842 51246 44861
rect 51246 44842 51260 44861
rect 51316 44842 51336 44861
rect 51336 44842 51350 44861
rect 51406 44842 51426 44861
rect 51426 44842 51440 44861
rect 51496 44842 51516 44861
rect 51516 44842 51530 44861
rect 51586 44842 51606 44861
rect 51606 44842 51620 44861
rect 51676 44842 51696 44861
rect 51696 44842 51710 44861
rect 51766 44842 51786 44861
rect 51786 44842 51800 44861
rect 51856 44842 51876 44861
rect 51876 44842 51890 44861
rect 51946 44842 51966 44861
rect 51966 44842 51980 44861
rect 52036 44842 52056 44861
rect 52056 44842 52070 44861
rect 52126 44842 52146 44861
rect 52146 44842 52160 44861
rect 52216 44842 52250 44876
rect 43170 44682 43204 44716
rect 43260 44714 43294 44716
rect 43350 44714 43384 44716
rect 43440 44714 43474 44716
rect 43530 44714 43564 44716
rect 43620 44714 43654 44716
rect 43710 44714 43744 44716
rect 43800 44714 43834 44716
rect 43890 44714 43924 44716
rect 43980 44714 44014 44716
rect 43260 44682 43280 44714
rect 43280 44682 43294 44714
rect 43350 44682 43370 44714
rect 43370 44682 43384 44714
rect 43440 44682 43460 44714
rect 43460 44682 43474 44714
rect 43530 44682 43550 44714
rect 43550 44682 43564 44714
rect 43620 44682 43640 44714
rect 43640 44682 43654 44714
rect 43710 44682 43730 44714
rect 43730 44682 43744 44714
rect 43800 44682 43820 44714
rect 43820 44682 43834 44714
rect 43890 44682 43910 44714
rect 43910 44682 43924 44714
rect 43980 44682 44000 44714
rect 44000 44682 44014 44714
rect 44070 44682 44104 44716
rect 43356 44506 43378 44512
rect 43378 44506 43390 44512
rect 43456 44506 43468 44512
rect 43468 44506 43490 44512
rect 43556 44506 43558 44512
rect 43558 44506 43590 44512
rect 43356 44478 43390 44506
rect 43456 44478 43490 44506
rect 43556 44478 43590 44506
rect 43656 44478 43690 44512
rect 43756 44478 43790 44512
rect 43856 44506 43884 44512
rect 43884 44506 43890 44512
rect 43856 44478 43890 44506
rect 43356 44378 43390 44412
rect 43456 44378 43490 44412
rect 43556 44378 43590 44412
rect 43656 44378 43690 44412
rect 43756 44378 43790 44412
rect 43856 44378 43890 44412
rect 43356 44278 43390 44312
rect 43456 44278 43490 44312
rect 43556 44278 43590 44312
rect 43656 44278 43690 44312
rect 43756 44278 43790 44312
rect 43856 44278 43890 44312
rect 43356 44180 43390 44212
rect 43456 44180 43490 44212
rect 43556 44180 43590 44212
rect 43356 44178 43378 44180
rect 43378 44178 43390 44180
rect 43456 44178 43468 44180
rect 43468 44178 43490 44180
rect 43556 44178 43558 44180
rect 43558 44178 43590 44180
rect 43656 44178 43690 44212
rect 43756 44178 43790 44212
rect 43856 44180 43890 44212
rect 43856 44178 43884 44180
rect 43884 44178 43890 44180
rect 43356 44090 43390 44112
rect 43456 44090 43490 44112
rect 43556 44090 43590 44112
rect 43356 44078 43378 44090
rect 43378 44078 43390 44090
rect 43456 44078 43468 44090
rect 43468 44078 43490 44090
rect 43556 44078 43558 44090
rect 43558 44078 43590 44090
rect 43656 44078 43690 44112
rect 43756 44078 43790 44112
rect 43856 44090 43890 44112
rect 43856 44078 43884 44090
rect 43884 44078 43890 44090
rect 43356 44000 43390 44012
rect 43456 44000 43490 44012
rect 43556 44000 43590 44012
rect 43356 43978 43378 44000
rect 43378 43978 43390 44000
rect 43456 43978 43468 44000
rect 43468 43978 43490 44000
rect 43556 43978 43558 44000
rect 43558 43978 43590 44000
rect 43656 43978 43690 44012
rect 43756 43978 43790 44012
rect 43856 44000 43890 44012
rect 43856 43978 43884 44000
rect 43884 43978 43890 44000
rect 44510 44682 44544 44716
rect 44600 44714 44634 44716
rect 44690 44714 44724 44716
rect 44780 44714 44814 44716
rect 44870 44714 44904 44716
rect 44960 44714 44994 44716
rect 45050 44714 45084 44716
rect 45140 44714 45174 44716
rect 45230 44714 45264 44716
rect 45320 44714 45354 44716
rect 44600 44682 44620 44714
rect 44620 44682 44634 44714
rect 44690 44682 44710 44714
rect 44710 44682 44724 44714
rect 44780 44682 44800 44714
rect 44800 44682 44814 44714
rect 44870 44682 44890 44714
rect 44890 44682 44904 44714
rect 44960 44682 44980 44714
rect 44980 44682 44994 44714
rect 45050 44682 45070 44714
rect 45070 44682 45084 44714
rect 45140 44682 45160 44714
rect 45160 44682 45174 44714
rect 45230 44682 45250 44714
rect 45250 44682 45264 44714
rect 45320 44682 45340 44714
rect 45340 44682 45354 44714
rect 45410 44682 45444 44716
rect 44696 44506 44718 44512
rect 44718 44506 44730 44512
rect 44796 44506 44808 44512
rect 44808 44506 44830 44512
rect 44896 44506 44898 44512
rect 44898 44506 44930 44512
rect 44696 44478 44730 44506
rect 44796 44478 44830 44506
rect 44896 44478 44930 44506
rect 44996 44478 45030 44512
rect 45096 44478 45130 44512
rect 45196 44506 45224 44512
rect 45224 44506 45230 44512
rect 45196 44478 45230 44506
rect 44696 44378 44730 44412
rect 44796 44378 44830 44412
rect 44896 44378 44930 44412
rect 44996 44378 45030 44412
rect 45096 44378 45130 44412
rect 45196 44378 45230 44412
rect 44696 44278 44730 44312
rect 44796 44278 44830 44312
rect 44896 44278 44930 44312
rect 44996 44278 45030 44312
rect 45096 44278 45130 44312
rect 45196 44278 45230 44312
rect 44696 44180 44730 44212
rect 44796 44180 44830 44212
rect 44896 44180 44930 44212
rect 44696 44178 44718 44180
rect 44718 44178 44730 44180
rect 44796 44178 44808 44180
rect 44808 44178 44830 44180
rect 44896 44178 44898 44180
rect 44898 44178 44930 44180
rect 44996 44178 45030 44212
rect 45096 44178 45130 44212
rect 45196 44180 45230 44212
rect 45196 44178 45224 44180
rect 45224 44178 45230 44180
rect 44696 44090 44730 44112
rect 44796 44090 44830 44112
rect 44896 44090 44930 44112
rect 44696 44078 44718 44090
rect 44718 44078 44730 44090
rect 44796 44078 44808 44090
rect 44808 44078 44830 44090
rect 44896 44078 44898 44090
rect 44898 44078 44930 44090
rect 44996 44078 45030 44112
rect 45096 44078 45130 44112
rect 45196 44090 45230 44112
rect 45196 44078 45224 44090
rect 45224 44078 45230 44090
rect 44696 44000 44730 44012
rect 44796 44000 44830 44012
rect 44896 44000 44930 44012
rect 44696 43978 44718 44000
rect 44718 43978 44730 44000
rect 44796 43978 44808 44000
rect 44808 43978 44830 44000
rect 44896 43978 44898 44000
rect 44898 43978 44930 44000
rect 44996 43978 45030 44012
rect 45096 43978 45130 44012
rect 45196 44000 45230 44012
rect 45196 43978 45224 44000
rect 45224 43978 45230 44000
rect 45850 44682 45884 44716
rect 45940 44714 45974 44716
rect 46030 44714 46064 44716
rect 46120 44714 46154 44716
rect 46210 44714 46244 44716
rect 46300 44714 46334 44716
rect 46390 44714 46424 44716
rect 46480 44714 46514 44716
rect 46570 44714 46604 44716
rect 46660 44714 46694 44716
rect 45940 44682 45960 44714
rect 45960 44682 45974 44714
rect 46030 44682 46050 44714
rect 46050 44682 46064 44714
rect 46120 44682 46140 44714
rect 46140 44682 46154 44714
rect 46210 44682 46230 44714
rect 46230 44682 46244 44714
rect 46300 44682 46320 44714
rect 46320 44682 46334 44714
rect 46390 44682 46410 44714
rect 46410 44682 46424 44714
rect 46480 44682 46500 44714
rect 46500 44682 46514 44714
rect 46570 44682 46590 44714
rect 46590 44682 46604 44714
rect 46660 44682 46680 44714
rect 46680 44682 46694 44714
rect 46750 44682 46784 44716
rect 46036 44506 46058 44512
rect 46058 44506 46070 44512
rect 46136 44506 46148 44512
rect 46148 44506 46170 44512
rect 46236 44506 46238 44512
rect 46238 44506 46270 44512
rect 46036 44478 46070 44506
rect 46136 44478 46170 44506
rect 46236 44478 46270 44506
rect 46336 44478 46370 44512
rect 46436 44478 46470 44512
rect 46536 44506 46564 44512
rect 46564 44506 46570 44512
rect 46536 44478 46570 44506
rect 46036 44378 46070 44412
rect 46136 44378 46170 44412
rect 46236 44378 46270 44412
rect 46336 44378 46370 44412
rect 46436 44378 46470 44412
rect 46536 44378 46570 44412
rect 46036 44278 46070 44312
rect 46136 44278 46170 44312
rect 46236 44278 46270 44312
rect 46336 44278 46370 44312
rect 46436 44278 46470 44312
rect 46536 44278 46570 44312
rect 46036 44180 46070 44212
rect 46136 44180 46170 44212
rect 46236 44180 46270 44212
rect 46036 44178 46058 44180
rect 46058 44178 46070 44180
rect 46136 44178 46148 44180
rect 46148 44178 46170 44180
rect 46236 44178 46238 44180
rect 46238 44178 46270 44180
rect 46336 44178 46370 44212
rect 46436 44178 46470 44212
rect 46536 44180 46570 44212
rect 46536 44178 46564 44180
rect 46564 44178 46570 44180
rect 46036 44090 46070 44112
rect 46136 44090 46170 44112
rect 46236 44090 46270 44112
rect 46036 44078 46058 44090
rect 46058 44078 46070 44090
rect 46136 44078 46148 44090
rect 46148 44078 46170 44090
rect 46236 44078 46238 44090
rect 46238 44078 46270 44090
rect 46336 44078 46370 44112
rect 46436 44078 46470 44112
rect 46536 44090 46570 44112
rect 46536 44078 46564 44090
rect 46564 44078 46570 44090
rect 46036 44000 46070 44012
rect 46136 44000 46170 44012
rect 46236 44000 46270 44012
rect 46036 43978 46058 44000
rect 46058 43978 46070 44000
rect 46136 43978 46148 44000
rect 46148 43978 46170 44000
rect 46236 43978 46238 44000
rect 46238 43978 46270 44000
rect 46336 43978 46370 44012
rect 46436 43978 46470 44012
rect 46536 44000 46570 44012
rect 46536 43978 46564 44000
rect 46564 43978 46570 44000
rect 47190 44682 47224 44716
rect 47280 44714 47314 44716
rect 47370 44714 47404 44716
rect 47460 44714 47494 44716
rect 47550 44714 47584 44716
rect 47640 44714 47674 44716
rect 47730 44714 47764 44716
rect 47820 44714 47854 44716
rect 47910 44714 47944 44716
rect 48000 44714 48034 44716
rect 47280 44682 47300 44714
rect 47300 44682 47314 44714
rect 47370 44682 47390 44714
rect 47390 44682 47404 44714
rect 47460 44682 47480 44714
rect 47480 44682 47494 44714
rect 47550 44682 47570 44714
rect 47570 44682 47584 44714
rect 47640 44682 47660 44714
rect 47660 44682 47674 44714
rect 47730 44682 47750 44714
rect 47750 44682 47764 44714
rect 47820 44682 47840 44714
rect 47840 44682 47854 44714
rect 47910 44682 47930 44714
rect 47930 44682 47944 44714
rect 48000 44682 48020 44714
rect 48020 44682 48034 44714
rect 48090 44682 48124 44716
rect 47376 44506 47398 44512
rect 47398 44506 47410 44512
rect 47476 44506 47488 44512
rect 47488 44506 47510 44512
rect 47576 44506 47578 44512
rect 47578 44506 47610 44512
rect 47376 44478 47410 44506
rect 47476 44478 47510 44506
rect 47576 44478 47610 44506
rect 47676 44478 47710 44512
rect 47776 44478 47810 44512
rect 47876 44506 47904 44512
rect 47904 44506 47910 44512
rect 47876 44478 47910 44506
rect 47376 44378 47410 44412
rect 47476 44378 47510 44412
rect 47576 44378 47610 44412
rect 47676 44378 47710 44412
rect 47776 44378 47810 44412
rect 47876 44378 47910 44412
rect 47376 44278 47410 44312
rect 47476 44278 47510 44312
rect 47576 44278 47610 44312
rect 47676 44278 47710 44312
rect 47776 44278 47810 44312
rect 47876 44278 47910 44312
rect 47376 44180 47410 44212
rect 47476 44180 47510 44212
rect 47576 44180 47610 44212
rect 47376 44178 47398 44180
rect 47398 44178 47410 44180
rect 47476 44178 47488 44180
rect 47488 44178 47510 44180
rect 47576 44178 47578 44180
rect 47578 44178 47610 44180
rect 47676 44178 47710 44212
rect 47776 44178 47810 44212
rect 47876 44180 47910 44212
rect 47876 44178 47904 44180
rect 47904 44178 47910 44180
rect 47376 44090 47410 44112
rect 47476 44090 47510 44112
rect 47576 44090 47610 44112
rect 47376 44078 47398 44090
rect 47398 44078 47410 44090
rect 47476 44078 47488 44090
rect 47488 44078 47510 44090
rect 47576 44078 47578 44090
rect 47578 44078 47610 44090
rect 47676 44078 47710 44112
rect 47776 44078 47810 44112
rect 47876 44090 47910 44112
rect 47876 44078 47904 44090
rect 47904 44078 47910 44090
rect 47376 44000 47410 44012
rect 47476 44000 47510 44012
rect 47576 44000 47610 44012
rect 47376 43978 47398 44000
rect 47398 43978 47410 44000
rect 47476 43978 47488 44000
rect 47488 43978 47510 44000
rect 47576 43978 47578 44000
rect 47578 43978 47610 44000
rect 47676 43978 47710 44012
rect 47776 43978 47810 44012
rect 47876 44000 47910 44012
rect 47876 43978 47904 44000
rect 47904 43978 47910 44000
rect 48530 44682 48564 44716
rect 48620 44714 48654 44716
rect 48710 44714 48744 44716
rect 48800 44714 48834 44716
rect 48890 44714 48924 44716
rect 48980 44714 49014 44716
rect 49070 44714 49104 44716
rect 49160 44714 49194 44716
rect 49250 44714 49284 44716
rect 49340 44714 49374 44716
rect 48620 44682 48640 44714
rect 48640 44682 48654 44714
rect 48710 44682 48730 44714
rect 48730 44682 48744 44714
rect 48800 44682 48820 44714
rect 48820 44682 48834 44714
rect 48890 44682 48910 44714
rect 48910 44682 48924 44714
rect 48980 44682 49000 44714
rect 49000 44682 49014 44714
rect 49070 44682 49090 44714
rect 49090 44682 49104 44714
rect 49160 44682 49180 44714
rect 49180 44682 49194 44714
rect 49250 44682 49270 44714
rect 49270 44682 49284 44714
rect 49340 44682 49360 44714
rect 49360 44682 49374 44714
rect 49430 44682 49464 44716
rect 48716 44506 48738 44512
rect 48738 44506 48750 44512
rect 48816 44506 48828 44512
rect 48828 44506 48850 44512
rect 48916 44506 48918 44512
rect 48918 44506 48950 44512
rect 48716 44478 48750 44506
rect 48816 44478 48850 44506
rect 48916 44478 48950 44506
rect 49016 44478 49050 44512
rect 49116 44478 49150 44512
rect 49216 44506 49244 44512
rect 49244 44506 49250 44512
rect 49216 44478 49250 44506
rect 48716 44378 48750 44412
rect 48816 44378 48850 44412
rect 48916 44378 48950 44412
rect 49016 44378 49050 44412
rect 49116 44378 49150 44412
rect 49216 44378 49250 44412
rect 48716 44278 48750 44312
rect 48816 44278 48850 44312
rect 48916 44278 48950 44312
rect 49016 44278 49050 44312
rect 49116 44278 49150 44312
rect 49216 44278 49250 44312
rect 48716 44180 48750 44212
rect 48816 44180 48850 44212
rect 48916 44180 48950 44212
rect 48716 44178 48738 44180
rect 48738 44178 48750 44180
rect 48816 44178 48828 44180
rect 48828 44178 48850 44180
rect 48916 44178 48918 44180
rect 48918 44178 48950 44180
rect 49016 44178 49050 44212
rect 49116 44178 49150 44212
rect 49216 44180 49250 44212
rect 49216 44178 49244 44180
rect 49244 44178 49250 44180
rect 48716 44090 48750 44112
rect 48816 44090 48850 44112
rect 48916 44090 48950 44112
rect 48716 44078 48738 44090
rect 48738 44078 48750 44090
rect 48816 44078 48828 44090
rect 48828 44078 48850 44090
rect 48916 44078 48918 44090
rect 48918 44078 48950 44090
rect 49016 44078 49050 44112
rect 49116 44078 49150 44112
rect 49216 44090 49250 44112
rect 49216 44078 49244 44090
rect 49244 44078 49250 44090
rect 48716 44000 48750 44012
rect 48816 44000 48850 44012
rect 48916 44000 48950 44012
rect 48716 43978 48738 44000
rect 48738 43978 48750 44000
rect 48816 43978 48828 44000
rect 48828 43978 48850 44000
rect 48916 43978 48918 44000
rect 48918 43978 48950 44000
rect 49016 43978 49050 44012
rect 49116 43978 49150 44012
rect 49216 44000 49250 44012
rect 49216 43978 49244 44000
rect 49244 43978 49250 44000
rect 49870 44682 49904 44716
rect 49960 44714 49994 44716
rect 50050 44714 50084 44716
rect 50140 44714 50174 44716
rect 50230 44714 50264 44716
rect 50320 44714 50354 44716
rect 50410 44714 50444 44716
rect 50500 44714 50534 44716
rect 50590 44714 50624 44716
rect 50680 44714 50714 44716
rect 49960 44682 49980 44714
rect 49980 44682 49994 44714
rect 50050 44682 50070 44714
rect 50070 44682 50084 44714
rect 50140 44682 50160 44714
rect 50160 44682 50174 44714
rect 50230 44682 50250 44714
rect 50250 44682 50264 44714
rect 50320 44682 50340 44714
rect 50340 44682 50354 44714
rect 50410 44682 50430 44714
rect 50430 44682 50444 44714
rect 50500 44682 50520 44714
rect 50520 44682 50534 44714
rect 50590 44682 50610 44714
rect 50610 44682 50624 44714
rect 50680 44682 50700 44714
rect 50700 44682 50714 44714
rect 50770 44682 50804 44716
rect 50056 44506 50078 44512
rect 50078 44506 50090 44512
rect 50156 44506 50168 44512
rect 50168 44506 50190 44512
rect 50256 44506 50258 44512
rect 50258 44506 50290 44512
rect 50056 44478 50090 44506
rect 50156 44478 50190 44506
rect 50256 44478 50290 44506
rect 50356 44478 50390 44512
rect 50456 44478 50490 44512
rect 50556 44506 50584 44512
rect 50584 44506 50590 44512
rect 50556 44478 50590 44506
rect 50056 44378 50090 44412
rect 50156 44378 50190 44412
rect 50256 44378 50290 44412
rect 50356 44378 50390 44412
rect 50456 44378 50490 44412
rect 50556 44378 50590 44412
rect 50056 44278 50090 44312
rect 50156 44278 50190 44312
rect 50256 44278 50290 44312
rect 50356 44278 50390 44312
rect 50456 44278 50490 44312
rect 50556 44278 50590 44312
rect 50056 44180 50090 44212
rect 50156 44180 50190 44212
rect 50256 44180 50290 44212
rect 50056 44178 50078 44180
rect 50078 44178 50090 44180
rect 50156 44178 50168 44180
rect 50168 44178 50190 44180
rect 50256 44178 50258 44180
rect 50258 44178 50290 44180
rect 50356 44178 50390 44212
rect 50456 44178 50490 44212
rect 50556 44180 50590 44212
rect 50556 44178 50584 44180
rect 50584 44178 50590 44180
rect 50056 44090 50090 44112
rect 50156 44090 50190 44112
rect 50256 44090 50290 44112
rect 50056 44078 50078 44090
rect 50078 44078 50090 44090
rect 50156 44078 50168 44090
rect 50168 44078 50190 44090
rect 50256 44078 50258 44090
rect 50258 44078 50290 44090
rect 50356 44078 50390 44112
rect 50456 44078 50490 44112
rect 50556 44090 50590 44112
rect 50556 44078 50584 44090
rect 50584 44078 50590 44090
rect 50056 44000 50090 44012
rect 50156 44000 50190 44012
rect 50256 44000 50290 44012
rect 50056 43978 50078 44000
rect 50078 43978 50090 44000
rect 50156 43978 50168 44000
rect 50168 43978 50190 44000
rect 50256 43978 50258 44000
rect 50258 43978 50290 44000
rect 50356 43978 50390 44012
rect 50456 43978 50490 44012
rect 50556 44000 50590 44012
rect 50556 43978 50584 44000
rect 50584 43978 50590 44000
rect 51210 44682 51244 44716
rect 51300 44714 51334 44716
rect 51390 44714 51424 44716
rect 51480 44714 51514 44716
rect 51570 44714 51604 44716
rect 51660 44714 51694 44716
rect 51750 44714 51784 44716
rect 51840 44714 51874 44716
rect 51930 44714 51964 44716
rect 52020 44714 52054 44716
rect 51300 44682 51320 44714
rect 51320 44682 51334 44714
rect 51390 44682 51410 44714
rect 51410 44682 51424 44714
rect 51480 44682 51500 44714
rect 51500 44682 51514 44714
rect 51570 44682 51590 44714
rect 51590 44682 51604 44714
rect 51660 44682 51680 44714
rect 51680 44682 51694 44714
rect 51750 44682 51770 44714
rect 51770 44682 51784 44714
rect 51840 44682 51860 44714
rect 51860 44682 51874 44714
rect 51930 44682 51950 44714
rect 51950 44682 51964 44714
rect 52020 44682 52040 44714
rect 52040 44682 52054 44714
rect 52110 44682 52144 44716
rect 51396 44506 51418 44512
rect 51418 44506 51430 44512
rect 51496 44506 51508 44512
rect 51508 44506 51530 44512
rect 51596 44506 51598 44512
rect 51598 44506 51630 44512
rect 51396 44478 51430 44506
rect 51496 44478 51530 44506
rect 51596 44478 51630 44506
rect 51696 44478 51730 44512
rect 51796 44478 51830 44512
rect 51896 44506 51924 44512
rect 51924 44506 51930 44512
rect 51896 44478 51930 44506
rect 51396 44378 51430 44412
rect 51496 44378 51530 44412
rect 51596 44378 51630 44412
rect 51696 44378 51730 44412
rect 51796 44378 51830 44412
rect 51896 44378 51930 44412
rect 51396 44278 51430 44312
rect 51496 44278 51530 44312
rect 51596 44278 51630 44312
rect 51696 44278 51730 44312
rect 51796 44278 51830 44312
rect 51896 44278 51930 44312
rect 51396 44180 51430 44212
rect 51496 44180 51530 44212
rect 51596 44180 51630 44212
rect 51396 44178 51418 44180
rect 51418 44178 51430 44180
rect 51496 44178 51508 44180
rect 51508 44178 51530 44180
rect 51596 44178 51598 44180
rect 51598 44178 51630 44180
rect 51696 44178 51730 44212
rect 51796 44178 51830 44212
rect 51896 44180 51930 44212
rect 51896 44178 51924 44180
rect 51924 44178 51930 44180
rect 51396 44090 51430 44112
rect 51496 44090 51530 44112
rect 51596 44090 51630 44112
rect 51396 44078 51418 44090
rect 51418 44078 51430 44090
rect 51496 44078 51508 44090
rect 51508 44078 51530 44090
rect 51596 44078 51598 44090
rect 51598 44078 51630 44090
rect 51696 44078 51730 44112
rect 51796 44078 51830 44112
rect 51896 44090 51930 44112
rect 51896 44078 51924 44090
rect 51924 44078 51930 44090
rect 51396 44000 51430 44012
rect 51496 44000 51530 44012
rect 51596 44000 51630 44012
rect 51396 43978 51418 44000
rect 51418 43978 51430 44000
rect 51496 43978 51508 44000
rect 51508 43978 51530 44000
rect 51596 43978 51598 44000
rect 51598 43978 51630 44000
rect 51696 43978 51730 44012
rect 51796 43978 51830 44012
rect 51896 44000 51930 44012
rect 51896 43978 51924 44000
rect 51924 43978 51930 44000
rect 15025 43537 15059 43571
rect 14565 43469 14599 43503
rect 29469 43435 29503 43469
rect 6101 43295 6135 43329
rect 6501 43295 6535 43329
rect 6901 43295 6935 43329
rect 7301 43295 7335 43329
rect 7701 43295 7735 43329
rect 8101 43295 8135 43329
rect 8501 43295 8535 43329
rect 8901 43295 8935 43329
rect 9301 43295 9335 43329
rect 9701 43295 9735 43329
rect 10101 43295 10135 43329
rect 10501 43295 10535 43329
rect 10901 43295 10935 43329
rect 11301 43295 11335 43329
rect 11701 43295 11735 43329
rect 12101 43295 12135 43329
rect 12501 43295 12535 43329
rect 12901 43295 12935 43329
rect 14301 43295 14335 43329
rect 15213 43295 15247 43329
rect 15613 43295 15647 43329
rect 16013 43295 16047 43329
rect 16413 43295 16447 43329
rect 16813 43295 16847 43329
rect 17213 43295 17247 43329
rect 17613 43295 17647 43329
rect 18013 43295 18047 43329
rect 18413 43295 18447 43329
rect 18813 43295 18847 43329
rect 19213 43295 19247 43329
rect 19613 43295 19647 43329
rect 20013 43295 20047 43329
rect 20413 43295 20447 43329
rect 20813 43295 20847 43329
rect 21213 43295 21247 43329
rect 21613 43295 21647 43329
rect 22013 43295 22047 43329
rect 22413 43295 22447 43329
rect 22813 43295 22847 43329
rect 23213 43295 23247 43329
rect 23613 43295 23647 43329
rect 24013 43295 24047 43329
rect 24413 43295 24447 43329
rect 24813 43295 24847 43329
rect 25213 43295 25247 43329
rect 25613 43295 25647 43329
rect 26013 43295 26047 43329
rect 26413 43295 26447 43329
rect 26813 43295 26847 43329
rect 27213 43295 27247 43329
rect 27613 43295 27647 43329
rect 28013 43295 28047 43329
rect 28413 43295 28447 43329
rect 28813 43295 28847 43329
rect 29213 43295 29247 43329
rect 29613 43295 29647 43329
rect 30013 43295 30047 43329
rect 30413 43295 30447 43329
rect 30813 43295 30847 43329
rect 31213 43295 31247 43329
rect 31613 43295 31647 43329
rect 32013 43295 32047 43329
rect 32413 43295 32447 43329
rect 32813 43295 32847 43329
rect 33213 43295 33247 43329
rect 33613 43295 33647 43329
rect 34013 43295 34047 43329
rect 34413 43295 34447 43329
rect 34813 43295 34847 43329
rect 35213 43295 35247 43329
rect 35613 43295 35647 43329
rect 36013 43295 36047 43329
rect 36413 43295 36447 43329
rect 36813 43295 36847 43329
rect 37213 43295 37247 43329
rect 37613 43295 37647 43329
rect 38013 43295 38047 43329
rect 38413 43295 38447 43329
rect 38813 43295 38847 43329
rect 39213 43295 39247 43329
rect 39613 43295 39647 43329
rect 40013 43295 40047 43329
rect 40413 43295 40447 43329
rect 40813 43295 40847 43329
rect 41213 43295 41247 43329
rect 41613 43295 41647 43329
rect 42013 43295 42047 43329
rect 42413 43295 42447 43329
rect 43143 43295 43177 43329
rect 43343 43295 43377 43329
rect 43543 43295 43577 43329
rect 43743 43295 43777 43329
rect 43943 43295 43977 43329
rect 44143 43295 44177 43329
rect 44343 43295 44377 43329
rect 44543 43295 44577 43329
rect 44743 43295 44777 43329
rect 44943 43295 44977 43329
rect 45143 43295 45177 43329
rect 45343 43295 45377 43329
rect 45543 43295 45577 43329
rect 45743 43295 45777 43329
rect 45943 43295 45977 43329
rect 46143 43295 46177 43329
rect 46343 43295 46377 43329
rect 46543 43295 46577 43329
rect 46743 43295 46777 43329
rect 46943 43295 46977 43329
rect 47143 43295 47177 43329
rect 47343 43295 47377 43329
rect 47543 43295 47577 43329
rect 47743 43295 47777 43329
rect 47943 43295 47977 43329
rect 48143 43295 48177 43329
rect 48343 43295 48377 43329
rect 48543 43295 48577 43329
rect 48743 43295 48777 43329
rect 48943 43295 48977 43329
rect 49143 43295 49177 43329
rect 49343 43295 49377 43329
rect 49543 43295 49577 43329
rect 49743 43295 49777 43329
rect 49943 43295 49977 43329
rect 50143 43295 50177 43329
rect 50343 43295 50377 43329
rect 50543 43295 50577 43329
rect 50743 43295 50777 43329
rect 50943 43295 50977 43329
rect 51143 43295 51177 43329
rect 51343 43295 51377 43329
rect 51543 43295 51577 43329
rect 51743 43295 51777 43329
rect 51943 43295 51977 43329
rect 52143 43295 52177 43329
rect 6493 41415 6527 41449
rect 6893 41415 6927 41449
rect 7293 41415 7327 41449
rect 7693 41415 7727 41449
rect 8093 41415 8127 41449
rect 8493 41415 8527 41449
rect 8893 41415 8927 41449
rect 9293 41415 9327 41449
rect 9693 41415 9727 41449
rect 10093 41415 10127 41449
rect 10493 41415 10527 41449
rect 10893 41415 10927 41449
rect 11293 41415 11327 41449
rect 11693 41415 11727 41449
rect 12093 41415 12127 41449
rect 12493 41415 12527 41449
rect 12893 41415 12927 41449
rect 13293 41415 13327 41449
rect 15313 41415 15347 41449
rect 15713 41415 15747 41449
rect 16113 41415 16147 41449
rect 16513 41415 16547 41449
rect 16913 41415 16947 41449
rect 17313 41415 17347 41449
rect 17713 41415 17747 41449
rect 18113 41415 18147 41449
rect 18513 41415 18547 41449
rect 18913 41415 18947 41449
rect 19313 41415 19347 41449
rect 19713 41415 19747 41449
rect 20113 41415 20147 41449
rect 20513 41415 20547 41449
rect 20913 41415 20947 41449
rect 21313 41415 21347 41449
rect 21713 41415 21747 41449
rect 22113 41415 22147 41449
rect 22857 41415 22891 41449
rect 23257 41415 23291 41449
rect 23657 41415 23691 41449
rect 24057 41415 24091 41449
rect 24457 41415 24491 41449
rect 24857 41415 24891 41449
rect 25257 41415 25291 41449
rect 25657 41415 25691 41449
rect 26057 41415 26091 41449
rect 26457 41415 26491 41449
rect 26857 41415 26891 41449
rect 27257 41415 27291 41449
rect 27657 41415 27691 41449
rect 28057 41415 28091 41449
rect 29521 41415 29555 41449
rect 29921 41415 29955 41449
rect 30321 41415 30355 41449
rect 30721 41415 30755 41449
rect 31121 41415 31155 41449
rect 31521 41415 31555 41449
rect 31921 41415 31955 41449
rect 32321 41415 32355 41449
rect 32721 41415 32755 41449
rect 33121 41415 33155 41449
rect 33521 41415 33555 41449
rect 33921 41415 33955 41449
rect 34321 41415 34355 41449
rect 34721 41415 34755 41449
rect 37459 41415 37493 41449
rect 37859 41415 37893 41449
rect 38259 41415 38293 41449
rect 38659 41415 38693 41449
rect 39059 41415 39093 41449
rect 39459 41415 39493 41449
rect 39859 41415 39893 41449
rect 40259 41415 40293 41449
rect 40659 41415 40693 41449
rect 41059 41415 41093 41449
rect 41967 41415 42001 41449
rect 42167 41415 42201 41449
rect 42367 41415 42401 41449
rect 42567 41415 42601 41449
rect 42767 41415 42801 41449
rect 42967 41415 43001 41449
rect 43167 41415 43201 41449
rect 43367 41415 43401 41449
rect 43567 41415 43601 41449
rect 43767 41415 43801 41449
rect 43967 41415 44001 41449
rect 44167 41415 44201 41449
rect 44367 41415 44401 41449
rect 44567 41415 44601 41449
rect 44767 41415 44801 41449
rect 44967 41415 45001 41449
rect 45167 41415 45201 41449
rect 45367 41415 45401 41449
rect 45567 41415 45601 41449
rect 45767 41415 45801 41449
rect 45967 41415 46001 41449
rect 46167 41415 46201 41449
rect 46367 41415 46401 41449
rect 46567 41415 46601 41449
rect 46767 41415 46801 41449
rect 46967 41415 47001 41449
rect 47167 41415 47201 41449
rect 47367 41415 47401 41449
rect 47567 41415 47601 41449
rect 47767 41415 47801 41449
rect 47967 41415 48001 41449
rect 48167 41415 48201 41449
rect 48367 41415 48401 41449
rect 48567 41415 48601 41449
rect 48767 41415 48801 41449
rect 48967 41415 49001 41449
rect 49167 41415 49201 41449
rect 49367 41415 49401 41449
rect 49567 41415 49601 41449
rect 49767 41415 49801 41449
rect 49967 41415 50001 41449
rect 50167 41415 50201 41449
rect 50367 41415 50401 41449
rect 50567 41415 50601 41449
rect 50767 41415 50801 41449
rect 50967 41415 51001 41449
rect 51167 41415 51201 41449
rect 51367 41415 51401 41449
rect 51567 41415 51601 41449
rect 51767 41415 51801 41449
rect 51967 41415 52001 41449
rect 52167 41415 52201 41449
rect 52367 41415 52401 41449
rect 22721 41147 22755 41181
rect 22721 41079 22755 41109
rect 22721 41075 22755 41079
rect 22721 41011 22755 41037
rect 22721 41003 22755 41011
rect 22721 40943 22755 40965
rect 22721 40931 22755 40943
rect 22721 40875 22755 40893
rect 22721 40859 22755 40875
rect 22721 40807 22755 40821
rect 22721 40787 22755 40807
rect 22721 40739 22755 40749
rect 22721 40715 22755 40739
rect 22721 40671 22755 40677
rect 22721 40643 22755 40671
rect 22721 40603 22755 40605
rect 22721 40571 22755 40603
rect 22721 40501 22755 40533
rect 22721 40499 22755 40501
rect 22721 40433 22755 40461
rect 22721 40427 22755 40433
rect 22721 40365 22755 40389
rect 22721 40355 22755 40365
rect 22721 40297 22755 40317
rect 22721 40283 22755 40297
rect 22721 40229 22755 40245
rect 22721 40211 22755 40229
rect 22721 40161 22755 40173
rect 22721 40139 22755 40161
rect 22721 40093 22755 40101
rect 22721 40067 22755 40093
rect 22721 40025 22755 40029
rect 22721 39995 22755 40025
rect 22721 39923 22755 39957
rect 23179 41147 23213 41181
rect 23179 41079 23213 41109
rect 23179 41075 23213 41079
rect 23179 41011 23213 41037
rect 23179 41003 23213 41011
rect 23179 40943 23213 40965
rect 23179 40931 23213 40943
rect 23179 40875 23213 40893
rect 23179 40859 23213 40875
rect 23179 40807 23213 40821
rect 23179 40787 23213 40807
rect 23179 40739 23213 40749
rect 23179 40715 23213 40739
rect 23179 40671 23213 40677
rect 23179 40643 23213 40671
rect 23179 40603 23213 40605
rect 23179 40571 23213 40603
rect 23179 40501 23213 40533
rect 23179 40499 23213 40501
rect 23179 40433 23213 40461
rect 23179 40427 23213 40433
rect 23179 40365 23213 40389
rect 23179 40355 23213 40365
rect 23179 40297 23213 40317
rect 23179 40283 23213 40297
rect 23179 40229 23213 40245
rect 23179 40211 23213 40229
rect 23179 40161 23213 40173
rect 23179 40139 23213 40161
rect 23179 40093 23213 40101
rect 23179 40067 23213 40093
rect 23179 40025 23213 40029
rect 23179 39995 23213 40025
rect 23179 39923 23213 39957
rect 23637 41147 23671 41181
rect 23637 41079 23671 41109
rect 23637 41075 23671 41079
rect 23637 41011 23671 41037
rect 23637 41003 23671 41011
rect 23637 40943 23671 40965
rect 23637 40931 23671 40943
rect 23637 40875 23671 40893
rect 23637 40859 23671 40875
rect 23637 40807 23671 40821
rect 23637 40787 23671 40807
rect 23637 40739 23671 40749
rect 23637 40715 23671 40739
rect 23637 40671 23671 40677
rect 23637 40643 23671 40671
rect 23637 40603 23671 40605
rect 23637 40571 23671 40603
rect 23637 40501 23671 40533
rect 23637 40499 23671 40501
rect 23637 40433 23671 40461
rect 23637 40427 23671 40433
rect 23637 40365 23671 40389
rect 23637 40355 23671 40365
rect 23637 40297 23671 40317
rect 23637 40283 23671 40297
rect 23637 40229 23671 40245
rect 23637 40211 23671 40229
rect 23637 40161 23671 40173
rect 23637 40139 23671 40161
rect 23637 40093 23671 40101
rect 23637 40067 23671 40093
rect 23637 40025 23671 40029
rect 23637 39995 23671 40025
rect 23637 39923 23671 39957
rect 22753 39797 22787 39831
rect 24869 41225 24903 41259
rect 24095 41147 24129 41181
rect 24095 41079 24129 41109
rect 24095 41075 24129 41079
rect 24095 41011 24129 41037
rect 24095 41003 24129 41011
rect 24095 40943 24129 40965
rect 24095 40931 24129 40943
rect 24095 40875 24129 40893
rect 24095 40859 24129 40875
rect 24095 40807 24129 40821
rect 24095 40787 24129 40807
rect 24095 40739 24129 40749
rect 24095 40715 24129 40739
rect 24095 40671 24129 40677
rect 24095 40643 24129 40671
rect 24095 40603 24129 40605
rect 24095 40571 24129 40603
rect 24095 40501 24129 40533
rect 24095 40499 24129 40501
rect 24095 40433 24129 40461
rect 24095 40427 24129 40433
rect 24095 40365 24129 40389
rect 24095 40355 24129 40365
rect 24095 40297 24129 40317
rect 24095 40283 24129 40297
rect 24095 40229 24129 40245
rect 24095 40211 24129 40229
rect 24095 40161 24129 40173
rect 24095 40139 24129 40161
rect 24095 40093 24129 40101
rect 24095 40067 24129 40093
rect 24095 40025 24129 40029
rect 24095 39995 24129 40025
rect 24095 39923 24129 39957
rect 24553 41147 24587 41181
rect 24553 41079 24587 41109
rect 24553 41075 24587 41079
rect 24553 41011 24587 41037
rect 24553 41003 24587 41011
rect 24553 40943 24587 40965
rect 24553 40931 24587 40943
rect 24553 40875 24587 40893
rect 24553 40859 24587 40875
rect 24553 40807 24587 40821
rect 24553 40787 24587 40807
rect 24553 40739 24587 40749
rect 24553 40715 24587 40739
rect 24553 40671 24587 40677
rect 24553 40643 24587 40671
rect 24553 40603 24587 40605
rect 24553 40571 24587 40603
rect 24553 40501 24587 40533
rect 24553 40499 24587 40501
rect 24553 40433 24587 40461
rect 24553 40427 24587 40433
rect 24553 40365 24587 40389
rect 24553 40355 24587 40365
rect 24553 40297 24587 40317
rect 24553 40283 24587 40297
rect 24553 40229 24587 40245
rect 24553 40211 24587 40229
rect 24553 40161 24587 40173
rect 24553 40139 24587 40161
rect 24553 40093 24587 40101
rect 24553 40067 24587 40093
rect 24553 40025 24587 40029
rect 24553 39995 24587 40025
rect 24553 39923 24587 39957
rect 25011 41147 25045 41181
rect 25011 41079 25045 41109
rect 25011 41075 25045 41079
rect 25011 41011 25045 41037
rect 25011 41003 25045 41011
rect 25011 40943 25045 40965
rect 25011 40931 25045 40943
rect 25011 40875 25045 40893
rect 25011 40859 25045 40875
rect 25011 40807 25045 40821
rect 25011 40787 25045 40807
rect 25011 40739 25045 40749
rect 25011 40715 25045 40739
rect 25011 40671 25045 40677
rect 25011 40643 25045 40671
rect 25011 40603 25045 40605
rect 25011 40571 25045 40603
rect 25011 40501 25045 40533
rect 25011 40499 25045 40501
rect 25011 40433 25045 40461
rect 25011 40427 25045 40433
rect 25011 40365 25045 40389
rect 25011 40355 25045 40365
rect 25011 40297 25045 40317
rect 25011 40283 25045 40297
rect 25011 40229 25045 40245
rect 25011 40211 25045 40229
rect 25011 40161 25045 40173
rect 25011 40139 25045 40161
rect 25011 40093 25045 40101
rect 25011 40067 25045 40093
rect 25011 40025 25045 40029
rect 25011 39995 25045 40025
rect 25011 39923 25045 39957
rect 25469 41147 25503 41181
rect 25469 41079 25503 41109
rect 25469 41075 25503 41079
rect 25469 41011 25503 41037
rect 25469 41003 25503 41011
rect 25469 40943 25503 40965
rect 25469 40931 25503 40943
rect 25469 40875 25503 40893
rect 25469 40859 25503 40875
rect 25469 40807 25503 40821
rect 25469 40787 25503 40807
rect 25469 40739 25503 40749
rect 25469 40715 25503 40739
rect 25469 40671 25503 40677
rect 25469 40643 25503 40671
rect 25469 40603 25503 40605
rect 25469 40571 25503 40603
rect 25469 40501 25503 40533
rect 25469 40499 25503 40501
rect 25469 40433 25503 40461
rect 25469 40427 25503 40433
rect 25469 40365 25503 40389
rect 25469 40355 25503 40365
rect 25469 40297 25503 40317
rect 25469 40283 25503 40297
rect 25469 40229 25503 40245
rect 25469 40211 25503 40229
rect 25469 40161 25503 40173
rect 25469 40139 25503 40161
rect 25469 40093 25503 40101
rect 25469 40067 25503 40093
rect 25469 40025 25503 40029
rect 25469 39995 25503 40025
rect 25469 39923 25503 39957
rect 25927 41147 25961 41181
rect 25927 41079 25961 41109
rect 25927 41075 25961 41079
rect 25927 41011 25961 41037
rect 25927 41003 25961 41011
rect 25927 40943 25961 40965
rect 25927 40931 25961 40943
rect 25927 40875 25961 40893
rect 25927 40859 25961 40875
rect 25927 40807 25961 40821
rect 25927 40787 25961 40807
rect 25927 40739 25961 40749
rect 25927 40715 25961 40739
rect 25927 40671 25961 40677
rect 25927 40643 25961 40671
rect 25927 40603 25961 40605
rect 25927 40571 25961 40603
rect 25927 40501 25961 40533
rect 25927 40499 25961 40501
rect 25927 40433 25961 40461
rect 25927 40427 25961 40433
rect 25927 40365 25961 40389
rect 25927 40355 25961 40365
rect 25927 40297 25961 40317
rect 25927 40283 25961 40297
rect 25927 40229 25961 40245
rect 25927 40211 25961 40229
rect 25927 40161 25961 40173
rect 25927 40139 25961 40161
rect 25927 40093 25961 40101
rect 25927 40067 25961 40093
rect 25927 40025 25961 40029
rect 25927 39995 25961 40025
rect 25927 39923 25961 39957
rect 26385 41147 26419 41181
rect 26385 41079 26419 41109
rect 26385 41075 26419 41079
rect 26385 41011 26419 41037
rect 26385 41003 26419 41011
rect 26385 40943 26419 40965
rect 26385 40931 26419 40943
rect 26385 40875 26419 40893
rect 26385 40859 26419 40875
rect 26385 40807 26419 40821
rect 26385 40787 26419 40807
rect 26385 40739 26419 40749
rect 26385 40715 26419 40739
rect 26385 40671 26419 40677
rect 26385 40643 26419 40671
rect 26385 40603 26419 40605
rect 26385 40571 26419 40603
rect 26385 40501 26419 40533
rect 26385 40499 26419 40501
rect 26385 40433 26419 40461
rect 26385 40427 26419 40433
rect 26385 40365 26419 40389
rect 26385 40355 26419 40365
rect 26385 40297 26419 40317
rect 26385 40283 26419 40297
rect 26385 40229 26419 40245
rect 26385 40211 26419 40229
rect 26385 40161 26419 40173
rect 26385 40139 26419 40161
rect 26385 40093 26419 40101
rect 26385 40067 26419 40093
rect 26385 40025 26419 40029
rect 26385 39995 26419 40025
rect 26385 39923 26419 39957
rect 26843 41147 26877 41181
rect 26843 41079 26877 41109
rect 26843 41075 26877 41079
rect 26843 41011 26877 41037
rect 26843 41003 26877 41011
rect 26843 40943 26877 40965
rect 26843 40931 26877 40943
rect 26843 40875 26877 40893
rect 26843 40859 26877 40875
rect 26843 40807 26877 40821
rect 26843 40787 26877 40807
rect 26843 40739 26877 40749
rect 26843 40715 26877 40739
rect 26843 40671 26877 40677
rect 26843 40643 26877 40671
rect 26843 40603 26877 40605
rect 26843 40571 26877 40603
rect 26843 40501 26877 40533
rect 26843 40499 26877 40501
rect 26843 40433 26877 40461
rect 26843 40427 26877 40433
rect 26843 40365 26877 40389
rect 26843 40355 26877 40365
rect 26843 40297 26877 40317
rect 26843 40283 26877 40297
rect 26843 40229 26877 40245
rect 26843 40211 26877 40229
rect 26843 40161 26877 40173
rect 26843 40139 26877 40161
rect 26843 40093 26877 40101
rect 26843 40067 26877 40093
rect 26843 40025 26877 40029
rect 26843 39995 26877 40025
rect 26843 39923 26877 39957
rect 27301 41147 27335 41181
rect 27301 41079 27335 41109
rect 27301 41075 27335 41079
rect 27301 41011 27335 41037
rect 27301 41003 27335 41011
rect 27301 40943 27335 40965
rect 27301 40931 27335 40943
rect 27301 40875 27335 40893
rect 27301 40859 27335 40875
rect 27301 40807 27335 40821
rect 27301 40787 27335 40807
rect 27301 40739 27335 40749
rect 27301 40715 27335 40739
rect 27301 40671 27335 40677
rect 27301 40643 27335 40671
rect 27301 40603 27335 40605
rect 27301 40571 27335 40603
rect 27301 40501 27335 40533
rect 27301 40499 27335 40501
rect 27301 40433 27335 40461
rect 27301 40427 27335 40433
rect 27301 40365 27335 40389
rect 27301 40355 27335 40365
rect 27301 40297 27335 40317
rect 27301 40283 27335 40297
rect 27301 40229 27335 40245
rect 27301 40211 27335 40229
rect 27301 40161 27335 40173
rect 27301 40139 27335 40161
rect 27301 40093 27335 40101
rect 27301 40067 27335 40093
rect 27301 40025 27335 40029
rect 27301 39995 27335 40025
rect 27301 39923 27335 39957
rect 27759 41147 27793 41181
rect 27759 41079 27793 41109
rect 27759 41075 27793 41079
rect 27759 41011 27793 41037
rect 27759 41003 27793 41011
rect 27759 40943 27793 40965
rect 27759 40931 27793 40943
rect 27759 40875 27793 40893
rect 27759 40859 27793 40875
rect 27759 40807 27793 40821
rect 27759 40787 27793 40807
rect 27759 40739 27793 40749
rect 27759 40715 27793 40739
rect 27759 40671 27793 40677
rect 27759 40643 27793 40671
rect 27759 40603 27793 40605
rect 27759 40571 27793 40603
rect 27759 40501 27793 40533
rect 27759 40499 27793 40501
rect 27759 40433 27793 40461
rect 27759 40427 27793 40433
rect 27759 40365 27793 40389
rect 27759 40355 27793 40365
rect 27759 40297 27793 40317
rect 27759 40283 27793 40297
rect 27759 40229 27793 40245
rect 27759 40211 27793 40229
rect 27759 40161 27793 40173
rect 27759 40139 27793 40161
rect 27759 40093 27793 40101
rect 27759 40067 27793 40093
rect 27759 40025 27793 40029
rect 27759 39995 27793 40025
rect 27759 39923 27793 39957
rect 28217 41147 28251 41181
rect 28217 41079 28251 41109
rect 28217 41075 28251 41079
rect 28217 41011 28251 41037
rect 28217 41003 28251 41011
rect 28217 40943 28251 40965
rect 28217 40931 28251 40943
rect 28217 40875 28251 40893
rect 28217 40859 28251 40875
rect 28217 40807 28251 40821
rect 28217 40787 28251 40807
rect 28217 40739 28251 40749
rect 28217 40715 28251 40739
rect 28217 40671 28251 40677
rect 28217 40643 28251 40671
rect 28217 40603 28251 40605
rect 28217 40571 28251 40603
rect 28217 40501 28251 40533
rect 28217 40499 28251 40501
rect 28217 40433 28251 40461
rect 28217 40427 28251 40433
rect 28217 40365 28251 40389
rect 28217 40355 28251 40365
rect 28217 40297 28251 40317
rect 28217 40283 28251 40297
rect 28217 40229 28251 40245
rect 28217 40211 28251 40229
rect 28217 40161 28251 40173
rect 28217 40139 28251 40161
rect 28217 40093 28251 40101
rect 28217 40067 28251 40093
rect 28217 40025 28251 40029
rect 28217 39995 28251 40025
rect 28217 39923 28251 39957
rect 28089 39797 28123 39831
rect 29385 41147 29419 41181
rect 29385 41079 29419 41109
rect 29385 41075 29419 41079
rect 29385 41011 29419 41037
rect 29385 41003 29419 41011
rect 29385 40943 29419 40965
rect 29385 40931 29419 40943
rect 29385 40875 29419 40893
rect 29385 40859 29419 40875
rect 29385 40807 29419 40821
rect 29385 40787 29419 40807
rect 29385 40739 29419 40749
rect 29385 40715 29419 40739
rect 29385 40671 29419 40677
rect 29385 40643 29419 40671
rect 29385 40603 29419 40605
rect 29385 40571 29419 40603
rect 29385 40501 29419 40533
rect 29385 40499 29419 40501
rect 29385 40433 29419 40461
rect 29385 40427 29419 40433
rect 29385 40365 29419 40389
rect 29385 40355 29419 40365
rect 29385 40297 29419 40317
rect 29385 40283 29419 40297
rect 29385 40229 29419 40245
rect 29385 40211 29419 40229
rect 29385 40161 29419 40173
rect 29385 40139 29419 40161
rect 29385 40093 29419 40101
rect 29385 40067 29419 40093
rect 29385 40025 29419 40029
rect 29385 39995 29419 40025
rect 29385 39923 29419 39957
rect 29843 41147 29877 41181
rect 29843 41079 29877 41109
rect 29843 41075 29877 41079
rect 29843 41011 29877 41037
rect 29843 41003 29877 41011
rect 29843 40943 29877 40965
rect 29843 40931 29877 40943
rect 29843 40875 29877 40893
rect 29843 40859 29877 40875
rect 29843 40807 29877 40821
rect 29843 40787 29877 40807
rect 29843 40739 29877 40749
rect 29843 40715 29877 40739
rect 29843 40671 29877 40677
rect 29843 40643 29877 40671
rect 29843 40603 29877 40605
rect 29843 40571 29877 40603
rect 29843 40501 29877 40533
rect 29843 40499 29877 40501
rect 29843 40433 29877 40461
rect 29843 40427 29877 40433
rect 29843 40365 29877 40389
rect 29843 40355 29877 40365
rect 29843 40297 29877 40317
rect 29843 40283 29877 40297
rect 29843 40229 29877 40245
rect 29843 40211 29877 40229
rect 29843 40161 29877 40173
rect 29843 40139 29877 40161
rect 29843 40093 29877 40101
rect 29843 40067 29877 40093
rect 29843 40025 29877 40029
rect 29843 39995 29877 40025
rect 29843 39923 29877 39957
rect 30301 41147 30335 41181
rect 30301 41079 30335 41109
rect 30301 41075 30335 41079
rect 30301 41011 30335 41037
rect 30301 41003 30335 41011
rect 30301 40943 30335 40965
rect 30301 40931 30335 40943
rect 30301 40875 30335 40893
rect 30301 40859 30335 40875
rect 30301 40807 30335 40821
rect 30301 40787 30335 40807
rect 30301 40739 30335 40749
rect 30301 40715 30335 40739
rect 30301 40671 30335 40677
rect 30301 40643 30335 40671
rect 30301 40603 30335 40605
rect 30301 40571 30335 40603
rect 30301 40501 30335 40533
rect 30301 40499 30335 40501
rect 30301 40433 30335 40461
rect 30301 40427 30335 40433
rect 30301 40365 30335 40389
rect 30301 40355 30335 40365
rect 30301 40297 30335 40317
rect 30301 40283 30335 40297
rect 30301 40229 30335 40245
rect 30301 40211 30335 40229
rect 30301 40161 30335 40173
rect 30301 40139 30335 40161
rect 30301 40093 30335 40101
rect 30301 40067 30335 40093
rect 30301 40025 30335 40029
rect 30301 39995 30335 40025
rect 30301 39923 30335 39957
rect 30759 41147 30793 41181
rect 30759 41079 30793 41109
rect 30759 41075 30793 41079
rect 30759 41011 30793 41037
rect 30759 41003 30793 41011
rect 30759 40943 30793 40965
rect 30759 40931 30793 40943
rect 30759 40875 30793 40893
rect 30759 40859 30793 40875
rect 30759 40807 30793 40821
rect 30759 40787 30793 40807
rect 30759 40739 30793 40749
rect 30759 40715 30793 40739
rect 30759 40671 30793 40677
rect 30759 40643 30793 40671
rect 30759 40603 30793 40605
rect 30759 40571 30793 40603
rect 30759 40501 30793 40533
rect 30759 40499 30793 40501
rect 30759 40433 30793 40461
rect 30759 40427 30793 40433
rect 30759 40365 30793 40389
rect 30759 40355 30793 40365
rect 30759 40297 30793 40317
rect 30759 40283 30793 40297
rect 30759 40229 30793 40245
rect 30759 40211 30793 40229
rect 30759 40161 30793 40173
rect 30759 40139 30793 40161
rect 30759 40093 30793 40101
rect 30759 40067 30793 40093
rect 30759 40025 30793 40029
rect 30759 39995 30793 40025
rect 30759 39923 30793 39957
rect 31217 41147 31251 41181
rect 31217 41079 31251 41109
rect 31217 41075 31251 41079
rect 31217 41011 31251 41037
rect 31217 41003 31251 41011
rect 31217 40943 31251 40965
rect 31217 40931 31251 40943
rect 31217 40875 31251 40893
rect 31217 40859 31251 40875
rect 31217 40807 31251 40821
rect 31217 40787 31251 40807
rect 31217 40739 31251 40749
rect 31217 40715 31251 40739
rect 31217 40671 31251 40677
rect 31217 40643 31251 40671
rect 31217 40603 31251 40605
rect 31217 40571 31251 40603
rect 31217 40501 31251 40533
rect 31217 40499 31251 40501
rect 31217 40433 31251 40461
rect 31217 40427 31251 40433
rect 31217 40365 31251 40389
rect 31217 40355 31251 40365
rect 31217 40297 31251 40317
rect 31217 40283 31251 40297
rect 31217 40229 31251 40245
rect 31217 40211 31251 40229
rect 31217 40161 31251 40173
rect 31217 40139 31251 40161
rect 31217 40093 31251 40101
rect 31217 40067 31251 40093
rect 31217 40025 31251 40029
rect 31217 39995 31251 40025
rect 31217 39923 31251 39957
rect 31675 41147 31709 41181
rect 31675 41079 31709 41109
rect 31675 41075 31709 41079
rect 31675 41011 31709 41037
rect 31675 41003 31709 41011
rect 31675 40943 31709 40965
rect 31675 40931 31709 40943
rect 31675 40875 31709 40893
rect 31675 40859 31709 40875
rect 31675 40807 31709 40821
rect 31675 40787 31709 40807
rect 31675 40739 31709 40749
rect 31675 40715 31709 40739
rect 31675 40671 31709 40677
rect 31675 40643 31709 40671
rect 31675 40603 31709 40605
rect 31675 40571 31709 40603
rect 31675 40501 31709 40533
rect 31675 40499 31709 40501
rect 31675 40433 31709 40461
rect 31675 40427 31709 40433
rect 31675 40365 31709 40389
rect 31675 40355 31709 40365
rect 31675 40297 31709 40317
rect 31675 40283 31709 40297
rect 31675 40229 31709 40245
rect 31675 40211 31709 40229
rect 31675 40161 31709 40173
rect 31675 40139 31709 40161
rect 31675 40093 31709 40101
rect 31675 40067 31709 40093
rect 31675 40025 31709 40029
rect 31675 39995 31709 40025
rect 31675 39923 31709 39957
rect 32133 41147 32167 41181
rect 32133 41079 32167 41109
rect 32133 41075 32167 41079
rect 32133 41011 32167 41037
rect 32133 41003 32167 41011
rect 32133 40943 32167 40965
rect 32133 40931 32167 40943
rect 32133 40875 32167 40893
rect 32133 40859 32167 40875
rect 32133 40807 32167 40821
rect 32133 40787 32167 40807
rect 32133 40739 32167 40749
rect 32133 40715 32167 40739
rect 32133 40671 32167 40677
rect 32133 40643 32167 40671
rect 32133 40603 32167 40605
rect 32133 40571 32167 40603
rect 32133 40501 32167 40533
rect 32133 40499 32167 40501
rect 32133 40433 32167 40461
rect 32133 40427 32167 40433
rect 32133 40365 32167 40389
rect 32133 40355 32167 40365
rect 32133 40297 32167 40317
rect 32133 40283 32167 40297
rect 32133 40229 32167 40245
rect 32133 40211 32167 40229
rect 32133 40161 32167 40173
rect 32133 40139 32167 40161
rect 32133 40093 32167 40101
rect 32133 40067 32167 40093
rect 32133 40025 32167 40029
rect 32133 39995 32167 40025
rect 32133 39923 32167 39957
rect 32591 41147 32625 41181
rect 32591 41079 32625 41109
rect 32591 41075 32625 41079
rect 32591 41011 32625 41037
rect 32591 41003 32625 41011
rect 32591 40943 32625 40965
rect 32591 40931 32625 40943
rect 32591 40875 32625 40893
rect 32591 40859 32625 40875
rect 32591 40807 32625 40821
rect 32591 40787 32625 40807
rect 32591 40739 32625 40749
rect 32591 40715 32625 40739
rect 32591 40671 32625 40677
rect 32591 40643 32625 40671
rect 32591 40603 32625 40605
rect 32591 40571 32625 40603
rect 32591 40501 32625 40533
rect 32591 40499 32625 40501
rect 32591 40433 32625 40461
rect 32591 40427 32625 40433
rect 32591 40365 32625 40389
rect 32591 40355 32625 40365
rect 32591 40297 32625 40317
rect 32591 40283 32625 40297
rect 32591 40229 32625 40245
rect 32591 40211 32625 40229
rect 32591 40161 32625 40173
rect 32591 40139 32625 40161
rect 32591 40093 32625 40101
rect 32591 40067 32625 40093
rect 32591 40025 32625 40029
rect 32591 39995 32625 40025
rect 32591 39923 32625 39957
rect 33049 41147 33083 41181
rect 33049 41079 33083 41109
rect 33049 41075 33083 41079
rect 33049 41011 33083 41037
rect 33049 41003 33083 41011
rect 33049 40943 33083 40965
rect 33049 40931 33083 40943
rect 33049 40875 33083 40893
rect 33049 40859 33083 40875
rect 33049 40807 33083 40821
rect 33049 40787 33083 40807
rect 33049 40739 33083 40749
rect 33049 40715 33083 40739
rect 33049 40671 33083 40677
rect 33049 40643 33083 40671
rect 33049 40603 33083 40605
rect 33049 40571 33083 40603
rect 33049 40501 33083 40533
rect 33049 40499 33083 40501
rect 33049 40433 33083 40461
rect 33049 40427 33083 40433
rect 33049 40365 33083 40389
rect 33049 40355 33083 40365
rect 33049 40297 33083 40317
rect 33049 40283 33083 40297
rect 33049 40229 33083 40245
rect 33049 40211 33083 40229
rect 33049 40161 33083 40173
rect 33049 40139 33083 40161
rect 33049 40093 33083 40101
rect 33049 40067 33083 40093
rect 33049 40025 33083 40029
rect 33049 39995 33083 40025
rect 33049 39923 33083 39957
rect 33507 41147 33541 41181
rect 33507 41079 33541 41109
rect 33507 41075 33541 41079
rect 33507 41011 33541 41037
rect 33507 41003 33541 41011
rect 33507 40943 33541 40965
rect 33507 40931 33541 40943
rect 33507 40875 33541 40893
rect 33507 40859 33541 40875
rect 33507 40807 33541 40821
rect 33507 40787 33541 40807
rect 33507 40739 33541 40749
rect 33507 40715 33541 40739
rect 33507 40671 33541 40677
rect 33507 40643 33541 40671
rect 33507 40603 33541 40605
rect 33507 40571 33541 40603
rect 33507 40501 33541 40533
rect 33507 40499 33541 40501
rect 33507 40433 33541 40461
rect 33507 40427 33541 40433
rect 33507 40365 33541 40389
rect 33507 40355 33541 40365
rect 33507 40297 33541 40317
rect 33507 40283 33541 40297
rect 33507 40229 33541 40245
rect 33507 40211 33541 40229
rect 33507 40161 33541 40173
rect 33507 40139 33541 40161
rect 33507 40093 33541 40101
rect 33507 40067 33541 40093
rect 33507 40025 33541 40029
rect 33507 39995 33541 40025
rect 33507 39923 33541 39957
rect 33965 41147 33999 41181
rect 33965 41079 33999 41109
rect 33965 41075 33999 41079
rect 33965 41011 33999 41037
rect 33965 41003 33999 41011
rect 33965 40943 33999 40965
rect 33965 40931 33999 40943
rect 33965 40875 33999 40893
rect 33965 40859 33999 40875
rect 33965 40807 33999 40821
rect 33965 40787 33999 40807
rect 33965 40739 33999 40749
rect 33965 40715 33999 40739
rect 33965 40671 33999 40677
rect 33965 40643 33999 40671
rect 33965 40603 33999 40605
rect 33965 40571 33999 40603
rect 33965 40501 33999 40533
rect 33965 40499 33999 40501
rect 33965 40433 33999 40461
rect 33965 40427 33999 40433
rect 33965 40365 33999 40389
rect 33965 40355 33999 40365
rect 33965 40297 33999 40317
rect 33965 40283 33999 40297
rect 33965 40229 33999 40245
rect 33965 40211 33999 40229
rect 33965 40161 33999 40173
rect 33965 40139 33999 40161
rect 33965 40093 33999 40101
rect 33965 40067 33999 40093
rect 33965 40025 33999 40029
rect 33965 39995 33999 40025
rect 33965 39923 33999 39957
rect 34423 41147 34457 41181
rect 34423 41079 34457 41109
rect 34423 41075 34457 41079
rect 34423 41011 34457 41037
rect 34423 41003 34457 41011
rect 34423 40943 34457 40965
rect 34423 40931 34457 40943
rect 34423 40875 34457 40893
rect 34423 40859 34457 40875
rect 34423 40807 34457 40821
rect 34423 40787 34457 40807
rect 34423 40739 34457 40749
rect 34423 40715 34457 40739
rect 34423 40671 34457 40677
rect 34423 40643 34457 40671
rect 34423 40603 34457 40605
rect 34423 40571 34457 40603
rect 34423 40501 34457 40533
rect 34423 40499 34457 40501
rect 34423 40433 34457 40461
rect 34423 40427 34457 40433
rect 34423 40365 34457 40389
rect 34423 40355 34457 40365
rect 34423 40297 34457 40317
rect 34423 40283 34457 40297
rect 34423 40229 34457 40245
rect 34423 40211 34457 40229
rect 34423 40161 34457 40173
rect 34423 40139 34457 40161
rect 34423 40093 34457 40101
rect 34423 40067 34457 40093
rect 34423 40025 34457 40029
rect 34423 39995 34457 40025
rect 34423 39923 34457 39957
rect 34881 41147 34915 41181
rect 34881 41079 34915 41109
rect 34881 41075 34915 41079
rect 34881 41011 34915 41037
rect 34881 41003 34915 41011
rect 34881 40943 34915 40965
rect 41830 41082 41864 41116
rect 41920 41101 41954 41116
rect 42010 41101 42044 41116
rect 42100 41101 42134 41116
rect 42190 41101 42224 41116
rect 42280 41101 42314 41116
rect 42370 41101 42404 41116
rect 42460 41101 42494 41116
rect 42550 41101 42584 41116
rect 42640 41101 42674 41116
rect 42730 41101 42764 41116
rect 42820 41101 42854 41116
rect 42910 41101 42944 41116
rect 41920 41082 41940 41101
rect 41940 41082 41954 41101
rect 42010 41082 42030 41101
rect 42030 41082 42044 41101
rect 42100 41082 42120 41101
rect 42120 41082 42134 41101
rect 42190 41082 42210 41101
rect 42210 41082 42224 41101
rect 42280 41082 42300 41101
rect 42300 41082 42314 41101
rect 42370 41082 42390 41101
rect 42390 41082 42404 41101
rect 42460 41082 42480 41101
rect 42480 41082 42494 41101
rect 42550 41082 42570 41101
rect 42570 41082 42584 41101
rect 42640 41082 42660 41101
rect 42660 41082 42674 41101
rect 42730 41082 42750 41101
rect 42750 41082 42764 41101
rect 42820 41082 42840 41101
rect 42840 41082 42854 41101
rect 42910 41082 42930 41101
rect 42930 41082 42944 41101
rect 43000 41082 43034 41116
rect 43170 41082 43204 41116
rect 43260 41101 43294 41116
rect 43350 41101 43384 41116
rect 43440 41101 43474 41116
rect 43530 41101 43564 41116
rect 43620 41101 43654 41116
rect 43710 41101 43744 41116
rect 43800 41101 43834 41116
rect 43890 41101 43924 41116
rect 43980 41101 44014 41116
rect 44070 41101 44104 41116
rect 44160 41101 44194 41116
rect 44250 41101 44284 41116
rect 43260 41082 43280 41101
rect 43280 41082 43294 41101
rect 43350 41082 43370 41101
rect 43370 41082 43384 41101
rect 43440 41082 43460 41101
rect 43460 41082 43474 41101
rect 43530 41082 43550 41101
rect 43550 41082 43564 41101
rect 43620 41082 43640 41101
rect 43640 41082 43654 41101
rect 43710 41082 43730 41101
rect 43730 41082 43744 41101
rect 43800 41082 43820 41101
rect 43820 41082 43834 41101
rect 43890 41082 43910 41101
rect 43910 41082 43924 41101
rect 43980 41082 44000 41101
rect 44000 41082 44014 41101
rect 44070 41082 44090 41101
rect 44090 41082 44104 41101
rect 44160 41082 44180 41101
rect 44180 41082 44194 41101
rect 44250 41082 44270 41101
rect 44270 41082 44284 41101
rect 44340 41082 44374 41116
rect 44510 41082 44544 41116
rect 44600 41101 44634 41116
rect 44690 41101 44724 41116
rect 44780 41101 44814 41116
rect 44870 41101 44904 41116
rect 44960 41101 44994 41116
rect 45050 41101 45084 41116
rect 45140 41101 45174 41116
rect 45230 41101 45264 41116
rect 45320 41101 45354 41116
rect 45410 41101 45444 41116
rect 45500 41101 45534 41116
rect 45590 41101 45624 41116
rect 44600 41082 44620 41101
rect 44620 41082 44634 41101
rect 44690 41082 44710 41101
rect 44710 41082 44724 41101
rect 44780 41082 44800 41101
rect 44800 41082 44814 41101
rect 44870 41082 44890 41101
rect 44890 41082 44904 41101
rect 44960 41082 44980 41101
rect 44980 41082 44994 41101
rect 45050 41082 45070 41101
rect 45070 41082 45084 41101
rect 45140 41082 45160 41101
rect 45160 41082 45174 41101
rect 45230 41082 45250 41101
rect 45250 41082 45264 41101
rect 45320 41082 45340 41101
rect 45340 41082 45354 41101
rect 45410 41082 45430 41101
rect 45430 41082 45444 41101
rect 45500 41082 45520 41101
rect 45520 41082 45534 41101
rect 45590 41082 45610 41101
rect 45610 41082 45624 41101
rect 45680 41082 45714 41116
rect 45850 41082 45884 41116
rect 45940 41101 45974 41116
rect 46030 41101 46064 41116
rect 46120 41101 46154 41116
rect 46210 41101 46244 41116
rect 46300 41101 46334 41116
rect 46390 41101 46424 41116
rect 46480 41101 46514 41116
rect 46570 41101 46604 41116
rect 46660 41101 46694 41116
rect 46750 41101 46784 41116
rect 46840 41101 46874 41116
rect 46930 41101 46964 41116
rect 45940 41082 45960 41101
rect 45960 41082 45974 41101
rect 46030 41082 46050 41101
rect 46050 41082 46064 41101
rect 46120 41082 46140 41101
rect 46140 41082 46154 41101
rect 46210 41082 46230 41101
rect 46230 41082 46244 41101
rect 46300 41082 46320 41101
rect 46320 41082 46334 41101
rect 46390 41082 46410 41101
rect 46410 41082 46424 41101
rect 46480 41082 46500 41101
rect 46500 41082 46514 41101
rect 46570 41082 46590 41101
rect 46590 41082 46604 41101
rect 46660 41082 46680 41101
rect 46680 41082 46694 41101
rect 46750 41082 46770 41101
rect 46770 41082 46784 41101
rect 46840 41082 46860 41101
rect 46860 41082 46874 41101
rect 46930 41082 46950 41101
rect 46950 41082 46964 41101
rect 47020 41082 47054 41116
rect 47190 41082 47224 41116
rect 47280 41101 47314 41116
rect 47370 41101 47404 41116
rect 47460 41101 47494 41116
rect 47550 41101 47584 41116
rect 47640 41101 47674 41116
rect 47730 41101 47764 41116
rect 47820 41101 47854 41116
rect 47910 41101 47944 41116
rect 48000 41101 48034 41116
rect 48090 41101 48124 41116
rect 48180 41101 48214 41116
rect 48270 41101 48304 41116
rect 47280 41082 47300 41101
rect 47300 41082 47314 41101
rect 47370 41082 47390 41101
rect 47390 41082 47404 41101
rect 47460 41082 47480 41101
rect 47480 41082 47494 41101
rect 47550 41082 47570 41101
rect 47570 41082 47584 41101
rect 47640 41082 47660 41101
rect 47660 41082 47674 41101
rect 47730 41082 47750 41101
rect 47750 41082 47764 41101
rect 47820 41082 47840 41101
rect 47840 41082 47854 41101
rect 47910 41082 47930 41101
rect 47930 41082 47944 41101
rect 48000 41082 48020 41101
rect 48020 41082 48034 41101
rect 48090 41082 48110 41101
rect 48110 41082 48124 41101
rect 48180 41082 48200 41101
rect 48200 41082 48214 41101
rect 48270 41082 48290 41101
rect 48290 41082 48304 41101
rect 48360 41082 48394 41116
rect 48530 41082 48564 41116
rect 48620 41101 48654 41116
rect 48710 41101 48744 41116
rect 48800 41101 48834 41116
rect 48890 41101 48924 41116
rect 48980 41101 49014 41116
rect 49070 41101 49104 41116
rect 49160 41101 49194 41116
rect 49250 41101 49284 41116
rect 49340 41101 49374 41116
rect 49430 41101 49464 41116
rect 49520 41101 49554 41116
rect 49610 41101 49644 41116
rect 48620 41082 48640 41101
rect 48640 41082 48654 41101
rect 48710 41082 48730 41101
rect 48730 41082 48744 41101
rect 48800 41082 48820 41101
rect 48820 41082 48834 41101
rect 48890 41082 48910 41101
rect 48910 41082 48924 41101
rect 48980 41082 49000 41101
rect 49000 41082 49014 41101
rect 49070 41082 49090 41101
rect 49090 41082 49104 41101
rect 49160 41082 49180 41101
rect 49180 41082 49194 41101
rect 49250 41082 49270 41101
rect 49270 41082 49284 41101
rect 49340 41082 49360 41101
rect 49360 41082 49374 41101
rect 49430 41082 49450 41101
rect 49450 41082 49464 41101
rect 49520 41082 49540 41101
rect 49540 41082 49554 41101
rect 49610 41082 49630 41101
rect 49630 41082 49644 41101
rect 49700 41082 49734 41116
rect 49870 41082 49904 41116
rect 49960 41101 49994 41116
rect 50050 41101 50084 41116
rect 50140 41101 50174 41116
rect 50230 41101 50264 41116
rect 50320 41101 50354 41116
rect 50410 41101 50444 41116
rect 50500 41101 50534 41116
rect 50590 41101 50624 41116
rect 50680 41101 50714 41116
rect 50770 41101 50804 41116
rect 50860 41101 50894 41116
rect 50950 41101 50984 41116
rect 49960 41082 49980 41101
rect 49980 41082 49994 41101
rect 50050 41082 50070 41101
rect 50070 41082 50084 41101
rect 50140 41082 50160 41101
rect 50160 41082 50174 41101
rect 50230 41082 50250 41101
rect 50250 41082 50264 41101
rect 50320 41082 50340 41101
rect 50340 41082 50354 41101
rect 50410 41082 50430 41101
rect 50430 41082 50444 41101
rect 50500 41082 50520 41101
rect 50520 41082 50534 41101
rect 50590 41082 50610 41101
rect 50610 41082 50624 41101
rect 50680 41082 50700 41101
rect 50700 41082 50714 41101
rect 50770 41082 50790 41101
rect 50790 41082 50804 41101
rect 50860 41082 50880 41101
rect 50880 41082 50894 41101
rect 50950 41082 50970 41101
rect 50970 41082 50984 41101
rect 51040 41082 51074 41116
rect 51210 41082 51244 41116
rect 51300 41101 51334 41116
rect 51390 41101 51424 41116
rect 51480 41101 51514 41116
rect 51570 41101 51604 41116
rect 51660 41101 51694 41116
rect 51750 41101 51784 41116
rect 51840 41101 51874 41116
rect 51930 41101 51964 41116
rect 52020 41101 52054 41116
rect 52110 41101 52144 41116
rect 52200 41101 52234 41116
rect 52290 41101 52324 41116
rect 51300 41082 51320 41101
rect 51320 41082 51334 41101
rect 51390 41082 51410 41101
rect 51410 41082 51424 41101
rect 51480 41082 51500 41101
rect 51500 41082 51514 41101
rect 51570 41082 51590 41101
rect 51590 41082 51604 41101
rect 51660 41082 51680 41101
rect 51680 41082 51694 41101
rect 51750 41082 51770 41101
rect 51770 41082 51784 41101
rect 51840 41082 51860 41101
rect 51860 41082 51874 41101
rect 51930 41082 51950 41101
rect 51950 41082 51964 41101
rect 52020 41082 52040 41101
rect 52040 41082 52054 41101
rect 52110 41082 52130 41101
rect 52130 41082 52144 41101
rect 52200 41082 52220 41101
rect 52220 41082 52234 41101
rect 52290 41082 52310 41101
rect 52310 41082 52324 41101
rect 52380 41082 52414 41116
rect 34881 40931 34915 40943
rect 34881 40875 34915 40893
rect 34881 40859 34915 40875
rect 34881 40807 34915 40821
rect 34881 40787 34915 40807
rect 34881 40739 34915 40749
rect 34881 40715 34915 40739
rect 34881 40671 34915 40677
rect 34881 40643 34915 40671
rect 34881 40603 34915 40605
rect 34881 40571 34915 40603
rect 34881 40501 34915 40533
rect 34881 40499 34915 40501
rect 34881 40433 34915 40461
rect 34881 40427 34915 40433
rect 34881 40365 34915 40389
rect 34881 40355 34915 40365
rect 34881 40297 34915 40317
rect 34881 40283 34915 40297
rect 34881 40229 34915 40245
rect 34881 40211 34915 40229
rect 37288 40909 37322 40929
rect 37288 40895 37322 40909
rect 37288 40841 37322 40857
rect 37288 40823 37322 40841
rect 37288 40773 37322 40785
rect 37288 40751 37322 40773
rect 37288 40705 37322 40713
rect 37288 40679 37322 40705
rect 37288 40637 37322 40641
rect 37288 40607 37322 40637
rect 37288 40535 37322 40569
rect 37288 40467 37322 40497
rect 37288 40463 37322 40467
rect 37288 40399 37322 40425
rect 37288 40391 37322 40399
rect 37288 40331 37322 40353
rect 37288 40319 37322 40331
rect 37288 40263 37322 40281
rect 37288 40247 37322 40263
rect 34881 40161 34915 40173
rect 34881 40139 34915 40161
rect 34881 40093 34915 40101
rect 34881 40067 34915 40093
rect 37288 40195 37322 40209
rect 37288 40175 37322 40195
rect 37746 40909 37780 40929
rect 37746 40895 37780 40909
rect 37746 40841 37780 40857
rect 37746 40823 37780 40841
rect 37746 40773 37780 40785
rect 37746 40751 37780 40773
rect 37746 40705 37780 40713
rect 37746 40679 37780 40705
rect 37746 40637 37780 40641
rect 37746 40607 37780 40637
rect 37746 40535 37780 40569
rect 37746 40467 37780 40497
rect 37746 40463 37780 40467
rect 37746 40399 37780 40425
rect 37746 40391 37780 40399
rect 37746 40331 37780 40353
rect 37746 40319 37780 40331
rect 37746 40263 37780 40281
rect 37746 40247 37780 40263
rect 37746 40195 37780 40209
rect 38204 40909 38238 40929
rect 38204 40895 38238 40909
rect 38204 40841 38238 40857
rect 38204 40823 38238 40841
rect 38204 40773 38238 40785
rect 38204 40751 38238 40773
rect 38204 40705 38238 40713
rect 38204 40679 38238 40705
rect 38204 40637 38238 40641
rect 38204 40607 38238 40637
rect 38204 40535 38238 40569
rect 38204 40467 38238 40497
rect 38204 40463 38238 40467
rect 38204 40399 38238 40425
rect 38204 40391 38238 40399
rect 38204 40331 38238 40353
rect 38204 40319 38238 40331
rect 38204 40263 38238 40281
rect 38204 40247 38238 40263
rect 37746 40175 37780 40195
rect 38204 40195 38238 40209
rect 38204 40175 38238 40195
rect 38662 40909 38696 40929
rect 38662 40895 38696 40909
rect 38662 40841 38696 40857
rect 38662 40823 38696 40841
rect 38662 40773 38696 40785
rect 38662 40751 38696 40773
rect 38662 40705 38696 40713
rect 38662 40679 38696 40705
rect 38662 40637 38696 40641
rect 38662 40607 38696 40637
rect 38662 40535 38696 40569
rect 38662 40467 38696 40497
rect 38662 40463 38696 40467
rect 38662 40399 38696 40425
rect 38662 40391 38696 40399
rect 38662 40331 38696 40353
rect 38662 40319 38696 40331
rect 38662 40263 38696 40281
rect 38662 40247 38696 40263
rect 38662 40195 38696 40209
rect 39120 40909 39154 40929
rect 39120 40895 39154 40909
rect 39120 40841 39154 40857
rect 39120 40823 39154 40841
rect 39120 40773 39154 40785
rect 39120 40751 39154 40773
rect 39120 40705 39154 40713
rect 39120 40679 39154 40705
rect 39120 40637 39154 40641
rect 39120 40607 39154 40637
rect 39120 40535 39154 40569
rect 39120 40467 39154 40497
rect 39120 40463 39154 40467
rect 39120 40399 39154 40425
rect 39120 40391 39154 40399
rect 39120 40331 39154 40353
rect 39120 40319 39154 40331
rect 39120 40263 39154 40281
rect 39120 40247 39154 40263
rect 38662 40175 38696 40195
rect 39120 40195 39154 40209
rect 39120 40175 39154 40195
rect 39578 40909 39612 40929
rect 39578 40895 39612 40909
rect 39578 40841 39612 40857
rect 39578 40823 39612 40841
rect 39578 40773 39612 40785
rect 39578 40751 39612 40773
rect 39578 40705 39612 40713
rect 39578 40679 39612 40705
rect 39578 40637 39612 40641
rect 39578 40607 39612 40637
rect 39578 40535 39612 40569
rect 39578 40467 39612 40497
rect 39578 40463 39612 40467
rect 39578 40399 39612 40425
rect 39578 40391 39612 40399
rect 39578 40331 39612 40353
rect 39578 40319 39612 40331
rect 39578 40263 39612 40281
rect 39578 40247 39612 40263
rect 39578 40195 39612 40209
rect 40036 40909 40070 40929
rect 40036 40895 40070 40909
rect 40036 40841 40070 40857
rect 40036 40823 40070 40841
rect 40036 40773 40070 40785
rect 40036 40751 40070 40773
rect 40036 40705 40070 40713
rect 40036 40679 40070 40705
rect 40036 40637 40070 40641
rect 40036 40607 40070 40637
rect 40036 40535 40070 40569
rect 40036 40467 40070 40497
rect 40036 40463 40070 40467
rect 40036 40399 40070 40425
rect 40036 40391 40070 40399
rect 40036 40331 40070 40353
rect 40036 40319 40070 40331
rect 40036 40263 40070 40281
rect 40036 40247 40070 40263
rect 39578 40175 39612 40195
rect 40036 40195 40070 40209
rect 40036 40175 40070 40195
rect 40494 40909 40528 40929
rect 40494 40895 40528 40909
rect 40494 40841 40528 40857
rect 40494 40823 40528 40841
rect 40494 40773 40528 40785
rect 40494 40751 40528 40773
rect 40494 40705 40528 40713
rect 40494 40679 40528 40705
rect 40494 40637 40528 40641
rect 40494 40607 40528 40637
rect 40494 40535 40528 40569
rect 40494 40467 40528 40497
rect 40494 40463 40528 40467
rect 40494 40399 40528 40425
rect 40494 40391 40528 40399
rect 40494 40331 40528 40353
rect 40494 40319 40528 40331
rect 40494 40263 40528 40281
rect 40494 40247 40528 40263
rect 40494 40195 40528 40209
rect 40952 40909 40986 40929
rect 40952 40895 40986 40909
rect 40952 40841 40986 40857
rect 40952 40823 40986 40841
rect 40952 40773 40986 40785
rect 40952 40751 40986 40773
rect 40952 40705 40986 40713
rect 40952 40679 40986 40705
rect 40952 40637 40986 40641
rect 40952 40607 40986 40637
rect 40952 40535 40986 40569
rect 40952 40467 40986 40497
rect 40952 40463 40986 40467
rect 40952 40399 40986 40425
rect 40952 40391 40986 40399
rect 40952 40331 40986 40353
rect 40952 40319 40986 40331
rect 40952 40263 40986 40281
rect 40952 40247 40986 40263
rect 40494 40175 40528 40195
rect 40952 40195 40986 40209
rect 40952 40175 40986 40195
rect 41410 40909 41444 40929
rect 41410 40895 41444 40909
rect 41410 40841 41444 40857
rect 41410 40823 41444 40841
rect 41410 40773 41444 40785
rect 41410 40751 41444 40773
rect 41410 40705 41444 40713
rect 41410 40679 41444 40705
rect 41410 40637 41444 40641
rect 41410 40607 41444 40637
rect 41410 40535 41444 40569
rect 41410 40467 41444 40497
rect 41410 40463 41444 40467
rect 41410 40399 41444 40425
rect 41410 40391 41444 40399
rect 41410 40331 41444 40353
rect 41410 40319 41444 40331
rect 41410 40263 41444 40281
rect 41410 40247 41444 40263
rect 41410 40195 41444 40209
rect 41410 40175 41444 40195
rect 34881 40025 34915 40029
rect 34881 39995 34915 40025
rect 34881 39923 34915 39957
rect 41994 40922 42028 40956
rect 42084 40954 42118 40956
rect 42174 40954 42208 40956
rect 42264 40954 42298 40956
rect 42354 40954 42388 40956
rect 42444 40954 42478 40956
rect 42534 40954 42568 40956
rect 42624 40954 42658 40956
rect 42714 40954 42748 40956
rect 42804 40954 42838 40956
rect 42084 40922 42104 40954
rect 42104 40922 42118 40954
rect 42174 40922 42194 40954
rect 42194 40922 42208 40954
rect 42264 40922 42284 40954
rect 42284 40922 42298 40954
rect 42354 40922 42374 40954
rect 42374 40922 42388 40954
rect 42444 40922 42464 40954
rect 42464 40922 42478 40954
rect 42534 40922 42554 40954
rect 42554 40922 42568 40954
rect 42624 40922 42644 40954
rect 42644 40922 42658 40954
rect 42714 40922 42734 40954
rect 42734 40922 42748 40954
rect 42804 40922 42824 40954
rect 42824 40922 42838 40954
rect 42894 40922 42928 40956
rect 42180 40746 42202 40752
rect 42202 40746 42214 40752
rect 42280 40746 42292 40752
rect 42292 40746 42314 40752
rect 42380 40746 42382 40752
rect 42382 40746 42414 40752
rect 42180 40718 42214 40746
rect 42280 40718 42314 40746
rect 42380 40718 42414 40746
rect 42480 40718 42514 40752
rect 42580 40718 42614 40752
rect 42680 40746 42708 40752
rect 42708 40746 42714 40752
rect 42680 40718 42714 40746
rect 42180 40618 42214 40652
rect 42280 40618 42314 40652
rect 42380 40618 42414 40652
rect 42480 40618 42514 40652
rect 42580 40618 42614 40652
rect 42680 40618 42714 40652
rect 42180 40518 42214 40552
rect 42280 40518 42314 40552
rect 42380 40518 42414 40552
rect 42480 40518 42514 40552
rect 42580 40518 42614 40552
rect 42680 40518 42714 40552
rect 42180 40420 42214 40452
rect 42280 40420 42314 40452
rect 42380 40420 42414 40452
rect 42180 40418 42202 40420
rect 42202 40418 42214 40420
rect 42280 40418 42292 40420
rect 42292 40418 42314 40420
rect 42380 40418 42382 40420
rect 42382 40418 42414 40420
rect 42480 40418 42514 40452
rect 42580 40418 42614 40452
rect 42680 40420 42714 40452
rect 42680 40418 42708 40420
rect 42708 40418 42714 40420
rect 42180 40330 42214 40352
rect 42280 40330 42314 40352
rect 42380 40330 42414 40352
rect 42180 40318 42202 40330
rect 42202 40318 42214 40330
rect 42280 40318 42292 40330
rect 42292 40318 42314 40330
rect 42380 40318 42382 40330
rect 42382 40318 42414 40330
rect 42480 40318 42514 40352
rect 42580 40318 42614 40352
rect 42680 40330 42714 40352
rect 42680 40318 42708 40330
rect 42708 40318 42714 40330
rect 42180 40240 42214 40252
rect 42280 40240 42314 40252
rect 42380 40240 42414 40252
rect 42180 40218 42202 40240
rect 42202 40218 42214 40240
rect 42280 40218 42292 40240
rect 42292 40218 42314 40240
rect 42380 40218 42382 40240
rect 42382 40218 42414 40240
rect 42480 40218 42514 40252
rect 42580 40218 42614 40252
rect 42680 40240 42714 40252
rect 42680 40218 42708 40240
rect 42708 40218 42714 40240
rect 43334 40922 43368 40956
rect 43424 40954 43458 40956
rect 43514 40954 43548 40956
rect 43604 40954 43638 40956
rect 43694 40954 43728 40956
rect 43784 40954 43818 40956
rect 43874 40954 43908 40956
rect 43964 40954 43998 40956
rect 44054 40954 44088 40956
rect 44144 40954 44178 40956
rect 43424 40922 43444 40954
rect 43444 40922 43458 40954
rect 43514 40922 43534 40954
rect 43534 40922 43548 40954
rect 43604 40922 43624 40954
rect 43624 40922 43638 40954
rect 43694 40922 43714 40954
rect 43714 40922 43728 40954
rect 43784 40922 43804 40954
rect 43804 40922 43818 40954
rect 43874 40922 43894 40954
rect 43894 40922 43908 40954
rect 43964 40922 43984 40954
rect 43984 40922 43998 40954
rect 44054 40922 44074 40954
rect 44074 40922 44088 40954
rect 44144 40922 44164 40954
rect 44164 40922 44178 40954
rect 44234 40922 44268 40956
rect 43520 40746 43542 40752
rect 43542 40746 43554 40752
rect 43620 40746 43632 40752
rect 43632 40746 43654 40752
rect 43720 40746 43722 40752
rect 43722 40746 43754 40752
rect 43520 40718 43554 40746
rect 43620 40718 43654 40746
rect 43720 40718 43754 40746
rect 43820 40718 43854 40752
rect 43920 40718 43954 40752
rect 44020 40746 44048 40752
rect 44048 40746 44054 40752
rect 44020 40718 44054 40746
rect 43520 40618 43554 40652
rect 43620 40618 43654 40652
rect 43720 40618 43754 40652
rect 43820 40618 43854 40652
rect 43920 40618 43954 40652
rect 44020 40618 44054 40652
rect 43520 40518 43554 40552
rect 43620 40518 43654 40552
rect 43720 40518 43754 40552
rect 43820 40518 43854 40552
rect 43920 40518 43954 40552
rect 44020 40518 44054 40552
rect 43520 40420 43554 40452
rect 43620 40420 43654 40452
rect 43720 40420 43754 40452
rect 43520 40418 43542 40420
rect 43542 40418 43554 40420
rect 43620 40418 43632 40420
rect 43632 40418 43654 40420
rect 43720 40418 43722 40420
rect 43722 40418 43754 40420
rect 43820 40418 43854 40452
rect 43920 40418 43954 40452
rect 44020 40420 44054 40452
rect 44020 40418 44048 40420
rect 44048 40418 44054 40420
rect 43520 40330 43554 40352
rect 43620 40330 43654 40352
rect 43720 40330 43754 40352
rect 43520 40318 43542 40330
rect 43542 40318 43554 40330
rect 43620 40318 43632 40330
rect 43632 40318 43654 40330
rect 43720 40318 43722 40330
rect 43722 40318 43754 40330
rect 43820 40318 43854 40352
rect 43920 40318 43954 40352
rect 44020 40330 44054 40352
rect 44020 40318 44048 40330
rect 44048 40318 44054 40330
rect 43520 40240 43554 40252
rect 43620 40240 43654 40252
rect 43720 40240 43754 40252
rect 43520 40218 43542 40240
rect 43542 40218 43554 40240
rect 43620 40218 43632 40240
rect 43632 40218 43654 40240
rect 43720 40218 43722 40240
rect 43722 40218 43754 40240
rect 43820 40218 43854 40252
rect 43920 40218 43954 40252
rect 44020 40240 44054 40252
rect 44020 40218 44048 40240
rect 44048 40218 44054 40240
rect 44674 40922 44708 40956
rect 44764 40954 44798 40956
rect 44854 40954 44888 40956
rect 44944 40954 44978 40956
rect 45034 40954 45068 40956
rect 45124 40954 45158 40956
rect 45214 40954 45248 40956
rect 45304 40954 45338 40956
rect 45394 40954 45428 40956
rect 45484 40954 45518 40956
rect 44764 40922 44784 40954
rect 44784 40922 44798 40954
rect 44854 40922 44874 40954
rect 44874 40922 44888 40954
rect 44944 40922 44964 40954
rect 44964 40922 44978 40954
rect 45034 40922 45054 40954
rect 45054 40922 45068 40954
rect 45124 40922 45144 40954
rect 45144 40922 45158 40954
rect 45214 40922 45234 40954
rect 45234 40922 45248 40954
rect 45304 40922 45324 40954
rect 45324 40922 45338 40954
rect 45394 40922 45414 40954
rect 45414 40922 45428 40954
rect 45484 40922 45504 40954
rect 45504 40922 45518 40954
rect 45574 40922 45608 40956
rect 44860 40746 44882 40752
rect 44882 40746 44894 40752
rect 44960 40746 44972 40752
rect 44972 40746 44994 40752
rect 45060 40746 45062 40752
rect 45062 40746 45094 40752
rect 44860 40718 44894 40746
rect 44960 40718 44994 40746
rect 45060 40718 45094 40746
rect 45160 40718 45194 40752
rect 45260 40718 45294 40752
rect 45360 40746 45388 40752
rect 45388 40746 45394 40752
rect 45360 40718 45394 40746
rect 44860 40618 44894 40652
rect 44960 40618 44994 40652
rect 45060 40618 45094 40652
rect 45160 40618 45194 40652
rect 45260 40618 45294 40652
rect 45360 40618 45394 40652
rect 44860 40518 44894 40552
rect 44960 40518 44994 40552
rect 45060 40518 45094 40552
rect 45160 40518 45194 40552
rect 45260 40518 45294 40552
rect 45360 40518 45394 40552
rect 44860 40420 44894 40452
rect 44960 40420 44994 40452
rect 45060 40420 45094 40452
rect 44860 40418 44882 40420
rect 44882 40418 44894 40420
rect 44960 40418 44972 40420
rect 44972 40418 44994 40420
rect 45060 40418 45062 40420
rect 45062 40418 45094 40420
rect 45160 40418 45194 40452
rect 45260 40418 45294 40452
rect 45360 40420 45394 40452
rect 45360 40418 45388 40420
rect 45388 40418 45394 40420
rect 44860 40330 44894 40352
rect 44960 40330 44994 40352
rect 45060 40330 45094 40352
rect 44860 40318 44882 40330
rect 44882 40318 44894 40330
rect 44960 40318 44972 40330
rect 44972 40318 44994 40330
rect 45060 40318 45062 40330
rect 45062 40318 45094 40330
rect 45160 40318 45194 40352
rect 45260 40318 45294 40352
rect 45360 40330 45394 40352
rect 45360 40318 45388 40330
rect 45388 40318 45394 40330
rect 44860 40240 44894 40252
rect 44960 40240 44994 40252
rect 45060 40240 45094 40252
rect 44860 40218 44882 40240
rect 44882 40218 44894 40240
rect 44960 40218 44972 40240
rect 44972 40218 44994 40240
rect 45060 40218 45062 40240
rect 45062 40218 45094 40240
rect 45160 40218 45194 40252
rect 45260 40218 45294 40252
rect 45360 40240 45394 40252
rect 45360 40218 45388 40240
rect 45388 40218 45394 40240
rect 46014 40922 46048 40956
rect 46104 40954 46138 40956
rect 46194 40954 46228 40956
rect 46284 40954 46318 40956
rect 46374 40954 46408 40956
rect 46464 40954 46498 40956
rect 46554 40954 46588 40956
rect 46644 40954 46678 40956
rect 46734 40954 46768 40956
rect 46824 40954 46858 40956
rect 46104 40922 46124 40954
rect 46124 40922 46138 40954
rect 46194 40922 46214 40954
rect 46214 40922 46228 40954
rect 46284 40922 46304 40954
rect 46304 40922 46318 40954
rect 46374 40922 46394 40954
rect 46394 40922 46408 40954
rect 46464 40922 46484 40954
rect 46484 40922 46498 40954
rect 46554 40922 46574 40954
rect 46574 40922 46588 40954
rect 46644 40922 46664 40954
rect 46664 40922 46678 40954
rect 46734 40922 46754 40954
rect 46754 40922 46768 40954
rect 46824 40922 46844 40954
rect 46844 40922 46858 40954
rect 46914 40922 46948 40956
rect 46200 40746 46222 40752
rect 46222 40746 46234 40752
rect 46300 40746 46312 40752
rect 46312 40746 46334 40752
rect 46400 40746 46402 40752
rect 46402 40746 46434 40752
rect 46200 40718 46234 40746
rect 46300 40718 46334 40746
rect 46400 40718 46434 40746
rect 46500 40718 46534 40752
rect 46600 40718 46634 40752
rect 46700 40746 46728 40752
rect 46728 40746 46734 40752
rect 46700 40718 46734 40746
rect 46200 40618 46234 40652
rect 46300 40618 46334 40652
rect 46400 40618 46434 40652
rect 46500 40618 46534 40652
rect 46600 40618 46634 40652
rect 46700 40618 46734 40652
rect 46200 40518 46234 40552
rect 46300 40518 46334 40552
rect 46400 40518 46434 40552
rect 46500 40518 46534 40552
rect 46600 40518 46634 40552
rect 46700 40518 46734 40552
rect 46200 40420 46234 40452
rect 46300 40420 46334 40452
rect 46400 40420 46434 40452
rect 46200 40418 46222 40420
rect 46222 40418 46234 40420
rect 46300 40418 46312 40420
rect 46312 40418 46334 40420
rect 46400 40418 46402 40420
rect 46402 40418 46434 40420
rect 46500 40418 46534 40452
rect 46600 40418 46634 40452
rect 46700 40420 46734 40452
rect 46700 40418 46728 40420
rect 46728 40418 46734 40420
rect 46200 40330 46234 40352
rect 46300 40330 46334 40352
rect 46400 40330 46434 40352
rect 46200 40318 46222 40330
rect 46222 40318 46234 40330
rect 46300 40318 46312 40330
rect 46312 40318 46334 40330
rect 46400 40318 46402 40330
rect 46402 40318 46434 40330
rect 46500 40318 46534 40352
rect 46600 40318 46634 40352
rect 46700 40330 46734 40352
rect 46700 40318 46728 40330
rect 46728 40318 46734 40330
rect 46200 40240 46234 40252
rect 46300 40240 46334 40252
rect 46400 40240 46434 40252
rect 46200 40218 46222 40240
rect 46222 40218 46234 40240
rect 46300 40218 46312 40240
rect 46312 40218 46334 40240
rect 46400 40218 46402 40240
rect 46402 40218 46434 40240
rect 46500 40218 46534 40252
rect 46600 40218 46634 40252
rect 46700 40240 46734 40252
rect 46700 40218 46728 40240
rect 46728 40218 46734 40240
rect 47354 40922 47388 40956
rect 47444 40954 47478 40956
rect 47534 40954 47568 40956
rect 47624 40954 47658 40956
rect 47714 40954 47748 40956
rect 47804 40954 47838 40956
rect 47894 40954 47928 40956
rect 47984 40954 48018 40956
rect 48074 40954 48108 40956
rect 48164 40954 48198 40956
rect 47444 40922 47464 40954
rect 47464 40922 47478 40954
rect 47534 40922 47554 40954
rect 47554 40922 47568 40954
rect 47624 40922 47644 40954
rect 47644 40922 47658 40954
rect 47714 40922 47734 40954
rect 47734 40922 47748 40954
rect 47804 40922 47824 40954
rect 47824 40922 47838 40954
rect 47894 40922 47914 40954
rect 47914 40922 47928 40954
rect 47984 40922 48004 40954
rect 48004 40922 48018 40954
rect 48074 40922 48094 40954
rect 48094 40922 48108 40954
rect 48164 40922 48184 40954
rect 48184 40922 48198 40954
rect 48254 40922 48288 40956
rect 47540 40746 47562 40752
rect 47562 40746 47574 40752
rect 47640 40746 47652 40752
rect 47652 40746 47674 40752
rect 47740 40746 47742 40752
rect 47742 40746 47774 40752
rect 47540 40718 47574 40746
rect 47640 40718 47674 40746
rect 47740 40718 47774 40746
rect 47840 40718 47874 40752
rect 47940 40718 47974 40752
rect 48040 40746 48068 40752
rect 48068 40746 48074 40752
rect 48040 40718 48074 40746
rect 47540 40618 47574 40652
rect 47640 40618 47674 40652
rect 47740 40618 47774 40652
rect 47840 40618 47874 40652
rect 47940 40618 47974 40652
rect 48040 40618 48074 40652
rect 47540 40518 47574 40552
rect 47640 40518 47674 40552
rect 47740 40518 47774 40552
rect 47840 40518 47874 40552
rect 47940 40518 47974 40552
rect 48040 40518 48074 40552
rect 47540 40420 47574 40452
rect 47640 40420 47674 40452
rect 47740 40420 47774 40452
rect 47540 40418 47562 40420
rect 47562 40418 47574 40420
rect 47640 40418 47652 40420
rect 47652 40418 47674 40420
rect 47740 40418 47742 40420
rect 47742 40418 47774 40420
rect 47840 40418 47874 40452
rect 47940 40418 47974 40452
rect 48040 40420 48074 40452
rect 48040 40418 48068 40420
rect 48068 40418 48074 40420
rect 47540 40330 47574 40352
rect 47640 40330 47674 40352
rect 47740 40330 47774 40352
rect 47540 40318 47562 40330
rect 47562 40318 47574 40330
rect 47640 40318 47652 40330
rect 47652 40318 47674 40330
rect 47740 40318 47742 40330
rect 47742 40318 47774 40330
rect 47840 40318 47874 40352
rect 47940 40318 47974 40352
rect 48040 40330 48074 40352
rect 48040 40318 48068 40330
rect 48068 40318 48074 40330
rect 47540 40240 47574 40252
rect 47640 40240 47674 40252
rect 47740 40240 47774 40252
rect 47540 40218 47562 40240
rect 47562 40218 47574 40240
rect 47640 40218 47652 40240
rect 47652 40218 47674 40240
rect 47740 40218 47742 40240
rect 47742 40218 47774 40240
rect 47840 40218 47874 40252
rect 47940 40218 47974 40252
rect 48040 40240 48074 40252
rect 48040 40218 48068 40240
rect 48068 40218 48074 40240
rect 48694 40922 48728 40956
rect 48784 40954 48818 40956
rect 48874 40954 48908 40956
rect 48964 40954 48998 40956
rect 49054 40954 49088 40956
rect 49144 40954 49178 40956
rect 49234 40954 49268 40956
rect 49324 40954 49358 40956
rect 49414 40954 49448 40956
rect 49504 40954 49538 40956
rect 48784 40922 48804 40954
rect 48804 40922 48818 40954
rect 48874 40922 48894 40954
rect 48894 40922 48908 40954
rect 48964 40922 48984 40954
rect 48984 40922 48998 40954
rect 49054 40922 49074 40954
rect 49074 40922 49088 40954
rect 49144 40922 49164 40954
rect 49164 40922 49178 40954
rect 49234 40922 49254 40954
rect 49254 40922 49268 40954
rect 49324 40922 49344 40954
rect 49344 40922 49358 40954
rect 49414 40922 49434 40954
rect 49434 40922 49448 40954
rect 49504 40922 49524 40954
rect 49524 40922 49538 40954
rect 49594 40922 49628 40956
rect 48880 40746 48902 40752
rect 48902 40746 48914 40752
rect 48980 40746 48992 40752
rect 48992 40746 49014 40752
rect 49080 40746 49082 40752
rect 49082 40746 49114 40752
rect 48880 40718 48914 40746
rect 48980 40718 49014 40746
rect 49080 40718 49114 40746
rect 49180 40718 49214 40752
rect 49280 40718 49314 40752
rect 49380 40746 49408 40752
rect 49408 40746 49414 40752
rect 49380 40718 49414 40746
rect 48880 40618 48914 40652
rect 48980 40618 49014 40652
rect 49080 40618 49114 40652
rect 49180 40618 49214 40652
rect 49280 40618 49314 40652
rect 49380 40618 49414 40652
rect 48880 40518 48914 40552
rect 48980 40518 49014 40552
rect 49080 40518 49114 40552
rect 49180 40518 49214 40552
rect 49280 40518 49314 40552
rect 49380 40518 49414 40552
rect 48880 40420 48914 40452
rect 48980 40420 49014 40452
rect 49080 40420 49114 40452
rect 48880 40418 48902 40420
rect 48902 40418 48914 40420
rect 48980 40418 48992 40420
rect 48992 40418 49014 40420
rect 49080 40418 49082 40420
rect 49082 40418 49114 40420
rect 49180 40418 49214 40452
rect 49280 40418 49314 40452
rect 49380 40420 49414 40452
rect 49380 40418 49408 40420
rect 49408 40418 49414 40420
rect 48880 40330 48914 40352
rect 48980 40330 49014 40352
rect 49080 40330 49114 40352
rect 48880 40318 48902 40330
rect 48902 40318 48914 40330
rect 48980 40318 48992 40330
rect 48992 40318 49014 40330
rect 49080 40318 49082 40330
rect 49082 40318 49114 40330
rect 49180 40318 49214 40352
rect 49280 40318 49314 40352
rect 49380 40330 49414 40352
rect 49380 40318 49408 40330
rect 49408 40318 49414 40330
rect 48880 40240 48914 40252
rect 48980 40240 49014 40252
rect 49080 40240 49114 40252
rect 48880 40218 48902 40240
rect 48902 40218 48914 40240
rect 48980 40218 48992 40240
rect 48992 40218 49014 40240
rect 49080 40218 49082 40240
rect 49082 40218 49114 40240
rect 49180 40218 49214 40252
rect 49280 40218 49314 40252
rect 49380 40240 49414 40252
rect 49380 40218 49408 40240
rect 49408 40218 49414 40240
rect 50034 40922 50068 40956
rect 50124 40954 50158 40956
rect 50214 40954 50248 40956
rect 50304 40954 50338 40956
rect 50394 40954 50428 40956
rect 50484 40954 50518 40956
rect 50574 40954 50608 40956
rect 50664 40954 50698 40956
rect 50754 40954 50788 40956
rect 50844 40954 50878 40956
rect 50124 40922 50144 40954
rect 50144 40922 50158 40954
rect 50214 40922 50234 40954
rect 50234 40922 50248 40954
rect 50304 40922 50324 40954
rect 50324 40922 50338 40954
rect 50394 40922 50414 40954
rect 50414 40922 50428 40954
rect 50484 40922 50504 40954
rect 50504 40922 50518 40954
rect 50574 40922 50594 40954
rect 50594 40922 50608 40954
rect 50664 40922 50684 40954
rect 50684 40922 50698 40954
rect 50754 40922 50774 40954
rect 50774 40922 50788 40954
rect 50844 40922 50864 40954
rect 50864 40922 50878 40954
rect 50934 40922 50968 40956
rect 50220 40746 50242 40752
rect 50242 40746 50254 40752
rect 50320 40746 50332 40752
rect 50332 40746 50354 40752
rect 50420 40746 50422 40752
rect 50422 40746 50454 40752
rect 50220 40718 50254 40746
rect 50320 40718 50354 40746
rect 50420 40718 50454 40746
rect 50520 40718 50554 40752
rect 50620 40718 50654 40752
rect 50720 40746 50748 40752
rect 50748 40746 50754 40752
rect 50720 40718 50754 40746
rect 50220 40618 50254 40652
rect 50320 40618 50354 40652
rect 50420 40618 50454 40652
rect 50520 40618 50554 40652
rect 50620 40618 50654 40652
rect 50720 40618 50754 40652
rect 50220 40518 50254 40552
rect 50320 40518 50354 40552
rect 50420 40518 50454 40552
rect 50520 40518 50554 40552
rect 50620 40518 50654 40552
rect 50720 40518 50754 40552
rect 50220 40420 50254 40452
rect 50320 40420 50354 40452
rect 50420 40420 50454 40452
rect 50220 40418 50242 40420
rect 50242 40418 50254 40420
rect 50320 40418 50332 40420
rect 50332 40418 50354 40420
rect 50420 40418 50422 40420
rect 50422 40418 50454 40420
rect 50520 40418 50554 40452
rect 50620 40418 50654 40452
rect 50720 40420 50754 40452
rect 50720 40418 50748 40420
rect 50748 40418 50754 40420
rect 50220 40330 50254 40352
rect 50320 40330 50354 40352
rect 50420 40330 50454 40352
rect 50220 40318 50242 40330
rect 50242 40318 50254 40330
rect 50320 40318 50332 40330
rect 50332 40318 50354 40330
rect 50420 40318 50422 40330
rect 50422 40318 50454 40330
rect 50520 40318 50554 40352
rect 50620 40318 50654 40352
rect 50720 40330 50754 40352
rect 50720 40318 50748 40330
rect 50748 40318 50754 40330
rect 50220 40240 50254 40252
rect 50320 40240 50354 40252
rect 50420 40240 50454 40252
rect 50220 40218 50242 40240
rect 50242 40218 50254 40240
rect 50320 40218 50332 40240
rect 50332 40218 50354 40240
rect 50420 40218 50422 40240
rect 50422 40218 50454 40240
rect 50520 40218 50554 40252
rect 50620 40218 50654 40252
rect 50720 40240 50754 40252
rect 50720 40218 50748 40240
rect 50748 40218 50754 40240
rect 51374 40922 51408 40956
rect 51464 40954 51498 40956
rect 51554 40954 51588 40956
rect 51644 40954 51678 40956
rect 51734 40954 51768 40956
rect 51824 40954 51858 40956
rect 51914 40954 51948 40956
rect 52004 40954 52038 40956
rect 52094 40954 52128 40956
rect 52184 40954 52218 40956
rect 51464 40922 51484 40954
rect 51484 40922 51498 40954
rect 51554 40922 51574 40954
rect 51574 40922 51588 40954
rect 51644 40922 51664 40954
rect 51664 40922 51678 40954
rect 51734 40922 51754 40954
rect 51754 40922 51768 40954
rect 51824 40922 51844 40954
rect 51844 40922 51858 40954
rect 51914 40922 51934 40954
rect 51934 40922 51948 40954
rect 52004 40922 52024 40954
rect 52024 40922 52038 40954
rect 52094 40922 52114 40954
rect 52114 40922 52128 40954
rect 52184 40922 52204 40954
rect 52204 40922 52218 40954
rect 52274 40922 52308 40956
rect 51560 40746 51582 40752
rect 51582 40746 51594 40752
rect 51660 40746 51672 40752
rect 51672 40746 51694 40752
rect 51760 40746 51762 40752
rect 51762 40746 51794 40752
rect 51560 40718 51594 40746
rect 51660 40718 51694 40746
rect 51760 40718 51794 40746
rect 51860 40718 51894 40752
rect 51960 40718 51994 40752
rect 52060 40746 52088 40752
rect 52088 40746 52094 40752
rect 52060 40718 52094 40746
rect 51560 40618 51594 40652
rect 51660 40618 51694 40652
rect 51760 40618 51794 40652
rect 51860 40618 51894 40652
rect 51960 40618 51994 40652
rect 52060 40618 52094 40652
rect 51560 40518 51594 40552
rect 51660 40518 51694 40552
rect 51760 40518 51794 40552
rect 51860 40518 51894 40552
rect 51960 40518 51994 40552
rect 52060 40518 52094 40552
rect 51560 40420 51594 40452
rect 51660 40420 51694 40452
rect 51760 40420 51794 40452
rect 51560 40418 51582 40420
rect 51582 40418 51594 40420
rect 51660 40418 51672 40420
rect 51672 40418 51694 40420
rect 51760 40418 51762 40420
rect 51762 40418 51794 40420
rect 51860 40418 51894 40452
rect 51960 40418 51994 40452
rect 52060 40420 52094 40452
rect 52060 40418 52088 40420
rect 52088 40418 52094 40420
rect 51560 40330 51594 40352
rect 51660 40330 51694 40352
rect 51760 40330 51794 40352
rect 51560 40318 51582 40330
rect 51582 40318 51594 40330
rect 51660 40318 51672 40330
rect 51672 40318 51694 40330
rect 51760 40318 51762 40330
rect 51762 40318 51794 40330
rect 51860 40318 51894 40352
rect 51960 40318 51994 40352
rect 52060 40330 52094 40352
rect 52060 40318 52088 40330
rect 52088 40318 52094 40330
rect 51560 40240 51594 40252
rect 51660 40240 51694 40252
rect 51760 40240 51794 40252
rect 51560 40218 51582 40240
rect 51582 40218 51594 40240
rect 51660 40218 51672 40240
rect 51672 40218 51694 40240
rect 51760 40218 51762 40240
rect 51762 40218 51794 40240
rect 51860 40218 51894 40252
rect 51960 40218 51994 40252
rect 52060 40240 52094 40252
rect 52060 40218 52088 40240
rect 52088 40218 52094 40240
rect 41429 39865 41463 39899
rect 28273 39661 28307 39695
rect 29469 39661 29503 39695
rect 6493 39535 6527 39569
rect 6893 39535 6927 39569
rect 7293 39535 7327 39569
rect 7693 39535 7727 39569
rect 8093 39535 8127 39569
rect 8493 39535 8527 39569
rect 8893 39535 8927 39569
rect 9293 39535 9327 39569
rect 9693 39535 9727 39569
rect 10093 39535 10127 39569
rect 10493 39535 10527 39569
rect 10893 39535 10927 39569
rect 11293 39535 11327 39569
rect 11693 39535 11727 39569
rect 12093 39535 12127 39569
rect 12493 39535 12527 39569
rect 12893 39535 12927 39569
rect 13293 39535 13327 39569
rect 15313 39535 15347 39569
rect 15713 39535 15747 39569
rect 16113 39535 16147 39569
rect 16513 39535 16547 39569
rect 16913 39535 16947 39569
rect 17313 39535 17347 39569
rect 17713 39535 17747 39569
rect 18113 39535 18147 39569
rect 18513 39535 18547 39569
rect 18913 39535 18947 39569
rect 19313 39535 19347 39569
rect 19713 39535 19747 39569
rect 20113 39535 20147 39569
rect 20513 39535 20547 39569
rect 20913 39535 20947 39569
rect 21313 39535 21347 39569
rect 21713 39535 21747 39569
rect 22113 39535 22147 39569
rect 22857 39535 22891 39569
rect 23257 39535 23291 39569
rect 23657 39535 23691 39569
rect 24057 39535 24091 39569
rect 24457 39535 24491 39569
rect 24857 39535 24891 39569
rect 25257 39535 25291 39569
rect 25657 39535 25691 39569
rect 26057 39535 26091 39569
rect 26457 39535 26491 39569
rect 26857 39535 26891 39569
rect 27257 39535 27291 39569
rect 27657 39535 27691 39569
rect 28057 39535 28091 39569
rect 29521 39535 29555 39569
rect 29921 39535 29955 39569
rect 30321 39535 30355 39569
rect 30721 39535 30755 39569
rect 31121 39535 31155 39569
rect 31521 39535 31555 39569
rect 31921 39535 31955 39569
rect 32321 39535 32355 39569
rect 32721 39535 32755 39569
rect 33121 39535 33155 39569
rect 33521 39535 33555 39569
rect 33921 39535 33955 39569
rect 34321 39535 34355 39569
rect 34721 39535 34755 39569
rect 37459 39535 37493 39569
rect 37859 39535 37893 39569
rect 38259 39535 38293 39569
rect 38659 39535 38693 39569
rect 39059 39535 39093 39569
rect 39459 39535 39493 39569
rect 39859 39535 39893 39569
rect 40259 39535 40293 39569
rect 40659 39535 40693 39569
rect 41059 39535 41093 39569
rect 41967 39535 42001 39569
rect 42167 39535 42201 39569
rect 42367 39535 42401 39569
rect 42567 39535 42601 39569
rect 42767 39535 42801 39569
rect 42967 39535 43001 39569
rect 43167 39535 43201 39569
rect 43367 39535 43401 39569
rect 43567 39535 43601 39569
rect 43767 39535 43801 39569
rect 43967 39535 44001 39569
rect 44167 39535 44201 39569
rect 44367 39535 44401 39569
rect 44567 39535 44601 39569
rect 44767 39535 44801 39569
rect 44967 39535 45001 39569
rect 45167 39535 45201 39569
rect 45367 39535 45401 39569
rect 45567 39535 45601 39569
rect 45767 39535 45801 39569
rect 45967 39535 46001 39569
rect 46167 39535 46201 39569
rect 46367 39535 46401 39569
rect 46567 39535 46601 39569
rect 46767 39535 46801 39569
rect 46967 39535 47001 39569
rect 47167 39535 47201 39569
rect 47367 39535 47401 39569
rect 47567 39535 47601 39569
rect 47767 39535 47801 39569
rect 47967 39535 48001 39569
rect 48167 39535 48201 39569
rect 48367 39535 48401 39569
rect 48567 39535 48601 39569
rect 48767 39535 48801 39569
rect 48967 39535 49001 39569
rect 49167 39535 49201 39569
rect 49367 39535 49401 39569
rect 49567 39535 49601 39569
rect 49767 39535 49801 39569
rect 49967 39535 50001 39569
rect 50167 39535 50201 39569
rect 50367 39535 50401 39569
rect 50567 39535 50601 39569
rect 50767 39535 50801 39569
rect 50967 39535 51001 39569
rect 51167 39535 51201 39569
rect 51367 39535 51401 39569
rect 51567 39535 51601 39569
rect 51767 39535 51801 39569
rect 51967 39535 52001 39569
rect 52167 39535 52201 39569
rect 52367 39535 52401 39569
rect 12175 37655 12209 37689
rect 12375 37655 12409 37689
rect 12575 37655 12609 37689
rect 12775 37655 12809 37689
rect 12975 37655 13009 37689
rect 13175 37655 13209 37689
rect 13861 37655 13895 37689
rect 14061 37655 14095 37689
rect 14261 37655 14295 37689
rect 14461 37655 14495 37689
rect 14661 37655 14695 37689
rect 14861 37655 14895 37689
rect 15061 37655 15095 37689
rect 15261 37655 15295 37689
rect 15461 37655 15495 37689
rect 15661 37655 15695 37689
rect 15861 37655 15895 37689
rect 16605 37655 16639 37689
rect 16805 37655 16839 37689
rect 17005 37655 17039 37689
rect 17205 37655 17239 37689
rect 17405 37655 17439 37689
rect 17605 37655 17639 37689
rect 17805 37655 17839 37689
rect 18005 37655 18039 37689
rect 18205 37655 18239 37689
rect 18405 37655 18439 37689
rect 18605 37655 18639 37689
rect 19351 37655 19385 37689
rect 19551 37655 19585 37689
rect 19751 37655 19785 37689
rect 19951 37655 19985 37689
rect 20151 37655 20185 37689
rect 20351 37655 20385 37689
rect 20551 37655 20585 37689
rect 20751 37655 20785 37689
rect 20951 37655 20985 37689
rect 21151 37655 21185 37689
rect 21351 37655 21385 37689
rect 21551 37655 21585 37689
rect 21751 37655 21785 37689
rect 21951 37655 21985 37689
rect 22681 37655 22715 37689
rect 22881 37655 22915 37689
rect 23081 37655 23115 37689
rect 23281 37655 23315 37689
rect 23481 37655 23515 37689
rect 23681 37655 23715 37689
rect 23881 37655 23915 37689
rect 24081 37655 24115 37689
rect 24281 37655 24315 37689
rect 24481 37655 24515 37689
rect 24681 37655 24715 37689
rect 25601 37655 25635 37689
rect 26001 37655 26035 37689
rect 26401 37655 26435 37689
rect 26801 37655 26835 37689
rect 27201 37655 27235 37689
rect 27601 37655 27635 37689
rect 28001 37655 28035 37689
rect 28401 37655 28435 37689
rect 28801 37655 28835 37689
rect 29201 37655 29235 37689
rect 30111 37655 30145 37689
rect 30511 37655 30545 37689
rect 30911 37655 30945 37689
rect 31311 37655 31345 37689
rect 31711 37655 31745 37689
rect 32111 37655 32145 37689
rect 32511 37655 32545 37689
rect 32911 37655 32945 37689
rect 33311 37655 33345 37689
rect 33711 37655 33745 37689
rect 34111 37655 34145 37689
rect 34511 37655 34545 37689
rect 34911 37655 34945 37689
rect 35311 37655 35345 37689
rect 35711 37655 35745 37689
rect 36111 37655 36145 37689
rect 36511 37655 36545 37689
rect 36911 37655 36945 37689
rect 37655 37655 37689 37689
rect 38055 37655 38089 37689
rect 38455 37655 38489 37689
rect 38855 37655 38889 37689
rect 39255 37655 39289 37689
rect 39655 37655 39689 37689
rect 40055 37655 40089 37689
rect 41967 37655 42001 37689
rect 42167 37655 42201 37689
rect 42367 37655 42401 37689
rect 42567 37655 42601 37689
rect 42767 37655 42801 37689
rect 42967 37655 43001 37689
rect 43167 37655 43201 37689
rect 43367 37655 43401 37689
rect 43567 37655 43601 37689
rect 43767 37655 43801 37689
rect 43967 37655 44001 37689
rect 44167 37655 44201 37689
rect 44367 37655 44401 37689
rect 44567 37655 44601 37689
rect 44767 37655 44801 37689
rect 44967 37655 45001 37689
rect 45167 37655 45201 37689
rect 45367 37655 45401 37689
rect 45567 37655 45601 37689
rect 45767 37655 45801 37689
rect 45967 37655 46001 37689
rect 46167 37655 46201 37689
rect 46367 37655 46401 37689
rect 46567 37655 46601 37689
rect 46767 37655 46801 37689
rect 46967 37655 47001 37689
rect 47167 37655 47201 37689
rect 47367 37655 47401 37689
rect 47567 37655 47601 37689
rect 47767 37655 47801 37689
rect 47967 37655 48001 37689
rect 48167 37655 48201 37689
rect 48367 37655 48401 37689
rect 48567 37655 48601 37689
rect 48767 37655 48801 37689
rect 48967 37655 49001 37689
rect 49167 37655 49201 37689
rect 49367 37655 49401 37689
rect 49567 37655 49601 37689
rect 49767 37655 49801 37689
rect 49967 37655 50001 37689
rect 50167 37655 50201 37689
rect 50367 37655 50401 37689
rect 50567 37655 50601 37689
rect 50767 37655 50801 37689
rect 50967 37655 51001 37689
rect 51167 37655 51201 37689
rect 51367 37655 51401 37689
rect 51567 37655 51601 37689
rect 51767 37655 51801 37689
rect 51967 37655 52001 37689
rect 52167 37655 52201 37689
rect 52367 37655 52401 37689
rect 12388 36986 12410 36992
rect 12410 36986 12422 36992
rect 12488 36986 12500 36992
rect 12500 36986 12522 36992
rect 12588 36986 12590 36992
rect 12590 36986 12622 36992
rect 12388 36958 12422 36986
rect 12488 36958 12522 36986
rect 12588 36958 12622 36986
rect 12688 36958 12722 36992
rect 12788 36958 12822 36992
rect 12888 36986 12916 36992
rect 12916 36986 12922 36992
rect 12888 36958 12922 36986
rect 12388 36858 12422 36892
rect 12488 36858 12522 36892
rect 12588 36858 12622 36892
rect 12688 36858 12722 36892
rect 12788 36858 12822 36892
rect 12888 36858 12922 36892
rect 12388 36758 12422 36792
rect 12488 36758 12522 36792
rect 12588 36758 12622 36792
rect 12688 36758 12722 36792
rect 12788 36758 12822 36792
rect 12888 36758 12922 36792
rect 12388 36660 12422 36692
rect 12488 36660 12522 36692
rect 12588 36660 12622 36692
rect 12388 36658 12410 36660
rect 12410 36658 12422 36660
rect 12488 36658 12500 36660
rect 12500 36658 12522 36660
rect 12588 36658 12590 36660
rect 12590 36658 12622 36660
rect 12688 36658 12722 36692
rect 12788 36658 12822 36692
rect 12888 36660 12922 36692
rect 12888 36658 12916 36660
rect 12916 36658 12922 36660
rect 12388 36570 12422 36592
rect 12488 36570 12522 36592
rect 12588 36570 12622 36592
rect 12388 36558 12410 36570
rect 12410 36558 12422 36570
rect 12488 36558 12500 36570
rect 12500 36558 12522 36570
rect 12588 36558 12590 36570
rect 12590 36558 12622 36570
rect 12688 36558 12722 36592
rect 12788 36558 12822 36592
rect 12888 36570 12922 36592
rect 12888 36558 12916 36570
rect 12916 36558 12922 36570
rect 12388 36480 12422 36492
rect 12488 36480 12522 36492
rect 12588 36480 12622 36492
rect 12388 36458 12410 36480
rect 12410 36458 12422 36480
rect 12488 36458 12500 36480
rect 12500 36458 12522 36480
rect 12588 36458 12590 36480
rect 12590 36458 12622 36480
rect 12688 36458 12722 36492
rect 12788 36458 12822 36492
rect 12888 36480 12922 36492
rect 12888 36458 12916 36480
rect 12916 36458 12922 36480
rect 13093 36261 13127 36295
rect 13697 36883 14091 37421
rect 15704 36883 16098 37421
rect 16441 36883 16835 37421
rect 18448 36883 18842 37421
rect 19186 36883 19580 37421
rect 21767 36883 22161 37421
rect 22517 36883 22911 37421
rect 24524 36883 24918 37421
rect 37565 37485 37599 37519
rect 37519 37387 37553 37421
rect 37519 37319 37553 37349
rect 37519 37315 37553 37319
rect 37519 37251 37553 37277
rect 37519 37243 37553 37251
rect 13277 36125 13311 36159
rect 13697 35923 14091 36461
rect 15704 35923 16098 36461
rect 16441 35923 16835 36461
rect 18448 35923 18842 36461
rect 19186 35923 19580 36461
rect 21767 35923 22161 36461
rect 22517 35923 22911 36461
rect 24524 35923 24918 36461
rect 25430 37149 25464 37169
rect 25430 37135 25464 37149
rect 25430 37081 25464 37097
rect 25430 37063 25464 37081
rect 25430 37013 25464 37025
rect 25430 36991 25464 37013
rect 25430 36945 25464 36953
rect 25430 36919 25464 36945
rect 25430 36877 25464 36881
rect 25430 36847 25464 36877
rect 25430 36775 25464 36809
rect 25430 36707 25464 36737
rect 25430 36703 25464 36707
rect 25430 36639 25464 36665
rect 25430 36631 25464 36639
rect 25430 36571 25464 36593
rect 25430 36559 25464 36571
rect 25430 36503 25464 36521
rect 25430 36487 25464 36503
rect 25430 36435 25464 36449
rect 25430 36415 25464 36435
rect 25888 37149 25922 37169
rect 25888 37135 25922 37149
rect 25888 37081 25922 37097
rect 25888 37063 25922 37081
rect 25888 37013 25922 37025
rect 25888 36991 25922 37013
rect 25888 36945 25922 36953
rect 25888 36919 25922 36945
rect 25888 36877 25922 36881
rect 25888 36847 25922 36877
rect 25888 36775 25922 36809
rect 25888 36707 25922 36737
rect 25888 36703 25922 36707
rect 25888 36639 25922 36665
rect 25888 36631 25922 36639
rect 25888 36571 25922 36593
rect 25888 36559 25922 36571
rect 25888 36503 25922 36521
rect 25888 36487 25922 36503
rect 25888 36435 25922 36449
rect 26346 37149 26380 37169
rect 26346 37135 26380 37149
rect 26346 37081 26380 37097
rect 26346 37063 26380 37081
rect 26346 37013 26380 37025
rect 26346 36991 26380 37013
rect 26346 36945 26380 36953
rect 26346 36919 26380 36945
rect 26346 36877 26380 36881
rect 26346 36847 26380 36877
rect 26346 36775 26380 36809
rect 26346 36707 26380 36737
rect 26346 36703 26380 36707
rect 26346 36639 26380 36665
rect 26346 36631 26380 36639
rect 26346 36571 26380 36593
rect 26346 36559 26380 36571
rect 26346 36503 26380 36521
rect 26346 36487 26380 36503
rect 25888 36415 25922 36435
rect 26346 36435 26380 36449
rect 26346 36415 26380 36435
rect 26804 37149 26838 37169
rect 26804 37135 26838 37149
rect 26804 37081 26838 37097
rect 26804 37063 26838 37081
rect 26804 37013 26838 37025
rect 26804 36991 26838 37013
rect 26804 36945 26838 36953
rect 26804 36919 26838 36945
rect 26804 36877 26838 36881
rect 26804 36847 26838 36877
rect 26804 36775 26838 36809
rect 26804 36707 26838 36737
rect 26804 36703 26838 36707
rect 26804 36639 26838 36665
rect 26804 36631 26838 36639
rect 26804 36571 26838 36593
rect 26804 36559 26838 36571
rect 26804 36503 26838 36521
rect 26804 36487 26838 36503
rect 26804 36435 26838 36449
rect 27262 37149 27296 37169
rect 27262 37135 27296 37149
rect 27262 37081 27296 37097
rect 27262 37063 27296 37081
rect 27262 37013 27296 37025
rect 27262 36991 27296 37013
rect 27262 36945 27296 36953
rect 27262 36919 27296 36945
rect 27262 36877 27296 36881
rect 27262 36847 27296 36877
rect 27262 36775 27296 36809
rect 27262 36707 27296 36737
rect 27262 36703 27296 36707
rect 27262 36639 27296 36665
rect 27262 36631 27296 36639
rect 27262 36571 27296 36593
rect 27262 36559 27296 36571
rect 27262 36503 27296 36521
rect 27262 36487 27296 36503
rect 26804 36415 26838 36435
rect 27262 36435 27296 36449
rect 27262 36415 27296 36435
rect 27720 37149 27754 37169
rect 27720 37135 27754 37149
rect 27720 37081 27754 37097
rect 27720 37063 27754 37081
rect 27720 37013 27754 37025
rect 27720 36991 27754 37013
rect 27720 36945 27754 36953
rect 27720 36919 27754 36945
rect 27720 36877 27754 36881
rect 27720 36847 27754 36877
rect 27720 36775 27754 36809
rect 27720 36707 27754 36737
rect 27720 36703 27754 36707
rect 27720 36639 27754 36665
rect 27720 36631 27754 36639
rect 27720 36571 27754 36593
rect 27720 36559 27754 36571
rect 27720 36503 27754 36521
rect 27720 36487 27754 36503
rect 27720 36435 27754 36449
rect 28178 37149 28212 37169
rect 28178 37135 28212 37149
rect 28178 37081 28212 37097
rect 28178 37063 28212 37081
rect 28178 37013 28212 37025
rect 28178 36991 28212 37013
rect 28178 36945 28212 36953
rect 28178 36919 28212 36945
rect 28178 36877 28212 36881
rect 28178 36847 28212 36877
rect 28178 36775 28212 36809
rect 28178 36707 28212 36737
rect 28178 36703 28212 36707
rect 28178 36639 28212 36665
rect 28178 36631 28212 36639
rect 28178 36571 28212 36593
rect 28178 36559 28212 36571
rect 28178 36503 28212 36521
rect 28178 36487 28212 36503
rect 27720 36415 27754 36435
rect 28178 36435 28212 36449
rect 28178 36415 28212 36435
rect 28636 37149 28670 37169
rect 28636 37135 28670 37149
rect 28636 37081 28670 37097
rect 28636 37063 28670 37081
rect 28636 37013 28670 37025
rect 28636 36991 28670 37013
rect 28636 36945 28670 36953
rect 28636 36919 28670 36945
rect 28636 36877 28670 36881
rect 28636 36847 28670 36877
rect 28636 36775 28670 36809
rect 28636 36707 28670 36737
rect 28636 36703 28670 36707
rect 28636 36639 28670 36665
rect 28636 36631 28670 36639
rect 28636 36571 28670 36593
rect 28636 36559 28670 36571
rect 28636 36503 28670 36521
rect 28636 36487 28670 36503
rect 28636 36435 28670 36449
rect 29094 37149 29128 37169
rect 29094 37135 29128 37149
rect 29094 37081 29128 37097
rect 29094 37063 29128 37081
rect 29094 37013 29128 37025
rect 29094 36991 29128 37013
rect 29094 36945 29128 36953
rect 29094 36919 29128 36945
rect 29094 36877 29128 36881
rect 29094 36847 29128 36877
rect 29094 36775 29128 36809
rect 29094 36707 29128 36737
rect 29094 36703 29128 36707
rect 29094 36639 29128 36665
rect 29094 36631 29128 36639
rect 29094 36571 29128 36593
rect 29094 36559 29128 36571
rect 29094 36503 29128 36521
rect 29094 36487 29128 36503
rect 28636 36415 28670 36435
rect 29094 36435 29128 36449
rect 29094 36415 29128 36435
rect 29552 37149 29586 37169
rect 29552 37135 29586 37149
rect 29552 37081 29586 37097
rect 29552 37063 29586 37081
rect 29552 37013 29586 37025
rect 29552 36991 29586 37013
rect 29552 36945 29586 36953
rect 29552 36919 29586 36945
rect 29552 36877 29586 36881
rect 29552 36847 29586 36877
rect 29552 36775 29586 36809
rect 29552 36707 29586 36737
rect 29552 36703 29586 36707
rect 29552 36639 29586 36665
rect 29552 36631 29586 36639
rect 29552 36571 29586 36593
rect 29552 36559 29586 36571
rect 29552 36503 29586 36521
rect 29552 36487 29586 36503
rect 29552 36435 29586 36449
rect 29552 36415 29586 36435
rect 37519 37183 37553 37205
rect 37519 37171 37553 37183
rect 37519 37115 37553 37133
rect 37519 37099 37553 37115
rect 37519 37047 37553 37061
rect 37519 37027 37553 37047
rect 37519 36979 37553 36989
rect 37519 36955 37553 36979
rect 37519 36911 37553 36917
rect 37519 36883 37553 36911
rect 37519 36843 37553 36845
rect 37519 36811 37553 36843
rect 37519 36741 37553 36773
rect 37519 36739 37553 36741
rect 37519 36673 37553 36701
rect 37519 36667 37553 36673
rect 37519 36605 37553 36629
rect 37519 36595 37553 36605
rect 37519 36537 37553 36557
rect 37519 36523 37553 36537
rect 37519 36469 37553 36485
rect 37519 36451 37553 36469
rect 37519 36401 37553 36413
rect 37519 36379 37553 36401
rect 37519 36333 37553 36341
rect 37519 36307 37553 36333
rect 37519 36265 37553 36269
rect 37519 36235 37553 36265
rect 37519 36163 37553 36197
rect 28089 36125 28123 36159
rect 37977 37387 38011 37421
rect 37977 37319 38011 37349
rect 37977 37315 38011 37319
rect 37977 37251 38011 37277
rect 37977 37243 38011 37251
rect 37977 37183 38011 37205
rect 37977 37171 38011 37183
rect 37977 37115 38011 37133
rect 37977 37099 38011 37115
rect 37977 37047 38011 37061
rect 37977 37027 38011 37047
rect 37977 36979 38011 36989
rect 37977 36955 38011 36979
rect 37977 36911 38011 36917
rect 37977 36883 38011 36911
rect 37977 36843 38011 36845
rect 37977 36811 38011 36843
rect 37977 36741 38011 36773
rect 37977 36739 38011 36741
rect 37977 36673 38011 36701
rect 37977 36667 38011 36673
rect 37977 36605 38011 36629
rect 37977 36595 38011 36605
rect 37977 36537 38011 36557
rect 37977 36523 38011 36537
rect 37977 36469 38011 36485
rect 37977 36451 38011 36469
rect 37977 36401 38011 36413
rect 37977 36379 38011 36401
rect 37977 36333 38011 36341
rect 37977 36307 38011 36333
rect 37977 36265 38011 36269
rect 37977 36235 38011 36265
rect 37977 36163 38011 36197
rect 38435 37387 38469 37421
rect 38435 37319 38469 37349
rect 38435 37315 38469 37319
rect 38435 37251 38469 37277
rect 38435 37243 38469 37251
rect 38435 37183 38469 37205
rect 38435 37171 38469 37183
rect 38435 37115 38469 37133
rect 38435 37099 38469 37115
rect 38435 37047 38469 37061
rect 38435 37027 38469 37047
rect 38435 36979 38469 36989
rect 38435 36955 38469 36979
rect 38435 36911 38469 36917
rect 38435 36883 38469 36911
rect 38435 36843 38469 36845
rect 38435 36811 38469 36843
rect 38435 36741 38469 36773
rect 38435 36739 38469 36741
rect 38435 36673 38469 36701
rect 38435 36667 38469 36673
rect 38435 36605 38469 36629
rect 38435 36595 38469 36605
rect 38435 36537 38469 36557
rect 38435 36523 38469 36537
rect 38435 36469 38469 36485
rect 38435 36451 38469 36469
rect 38435 36401 38469 36413
rect 38435 36379 38469 36401
rect 38435 36333 38469 36341
rect 38435 36307 38469 36333
rect 38435 36265 38469 36269
rect 38435 36235 38469 36265
rect 38435 36163 38469 36197
rect 38893 37387 38927 37421
rect 38893 37319 38927 37349
rect 38893 37315 38927 37319
rect 38893 37251 38927 37277
rect 38893 37243 38927 37251
rect 38893 37183 38927 37205
rect 38893 37171 38927 37183
rect 38893 37115 38927 37133
rect 38893 37099 38927 37115
rect 38893 37047 38927 37061
rect 38893 37027 38927 37047
rect 38893 36979 38927 36989
rect 38893 36955 38927 36979
rect 38893 36911 38927 36917
rect 38893 36883 38927 36911
rect 38893 36843 38927 36845
rect 38893 36811 38927 36843
rect 38893 36741 38927 36773
rect 38893 36739 38927 36741
rect 38893 36673 38927 36701
rect 38893 36667 38927 36673
rect 38893 36605 38927 36629
rect 38893 36595 38927 36605
rect 38893 36537 38927 36557
rect 38893 36523 38927 36537
rect 38893 36469 38927 36485
rect 38893 36451 38927 36469
rect 38893 36401 38927 36413
rect 38893 36379 38927 36401
rect 38893 36333 38927 36341
rect 38893 36307 38927 36333
rect 38893 36265 38927 36269
rect 38893 36235 38927 36265
rect 38893 36163 38927 36197
rect 39351 37387 39385 37421
rect 39351 37319 39385 37349
rect 39351 37315 39385 37319
rect 39351 37251 39385 37277
rect 39351 37243 39385 37251
rect 39351 37183 39385 37205
rect 39351 37171 39385 37183
rect 39351 37115 39385 37133
rect 39351 37099 39385 37115
rect 39351 37047 39385 37061
rect 39351 37027 39385 37047
rect 39351 36979 39385 36989
rect 39351 36955 39385 36979
rect 39351 36911 39385 36917
rect 39351 36883 39385 36911
rect 39351 36843 39385 36845
rect 39351 36811 39385 36843
rect 39351 36741 39385 36773
rect 39351 36739 39385 36741
rect 39351 36673 39385 36701
rect 39351 36667 39385 36673
rect 39351 36605 39385 36629
rect 39351 36595 39385 36605
rect 39351 36537 39385 36557
rect 39351 36523 39385 36537
rect 39351 36469 39385 36485
rect 39351 36451 39385 36469
rect 39351 36401 39385 36413
rect 39351 36379 39385 36401
rect 39351 36333 39385 36341
rect 39351 36307 39385 36333
rect 39351 36265 39385 36269
rect 39351 36235 39385 36265
rect 39351 36163 39385 36197
rect 39809 37387 39843 37421
rect 39809 37319 39843 37349
rect 39809 37315 39843 37319
rect 39809 37251 39843 37277
rect 39809 37243 39843 37251
rect 39809 37183 39843 37205
rect 39809 37171 39843 37183
rect 39809 37115 39843 37133
rect 39809 37099 39843 37115
rect 39809 37047 39843 37061
rect 39809 37027 39843 37047
rect 39809 36979 39843 36989
rect 39809 36955 39843 36979
rect 39809 36911 39843 36917
rect 39809 36883 39843 36911
rect 39809 36843 39843 36845
rect 39809 36811 39843 36843
rect 39809 36741 39843 36773
rect 39809 36739 39843 36741
rect 39809 36673 39843 36701
rect 39809 36667 39843 36673
rect 39809 36605 39843 36629
rect 39809 36595 39843 36605
rect 39809 36537 39843 36557
rect 39809 36523 39843 36537
rect 39809 36469 39843 36485
rect 39809 36451 39843 36469
rect 39809 36401 39843 36413
rect 39809 36379 39843 36401
rect 39809 36333 39843 36341
rect 39809 36307 39843 36333
rect 39809 36265 39843 36269
rect 39809 36235 39843 36265
rect 39809 36163 39843 36197
rect 40267 37387 40301 37421
rect 40267 37319 40301 37349
rect 40267 37315 40301 37319
rect 40267 37251 40301 37277
rect 40267 37243 40301 37251
rect 40267 37183 40301 37205
rect 40267 37171 40301 37183
rect 40267 37115 40301 37133
rect 40267 37099 40301 37115
rect 40267 37047 40301 37061
rect 40267 37027 40301 37047
rect 40267 36979 40301 36989
rect 40267 36955 40301 36979
rect 40267 36911 40301 36917
rect 40267 36883 40301 36911
rect 40267 36843 40301 36845
rect 40267 36811 40301 36843
rect 40267 36741 40301 36773
rect 40267 36739 40301 36741
rect 40267 36673 40301 36701
rect 40267 36667 40301 36673
rect 40267 36605 40301 36629
rect 40267 36595 40301 36605
rect 40267 36537 40301 36557
rect 40267 36523 40301 36537
rect 40267 36469 40301 36485
rect 40267 36451 40301 36469
rect 40267 36401 40301 36413
rect 40267 36379 40301 36401
rect 40267 36333 40301 36341
rect 40267 36307 40301 36333
rect 40267 36265 40301 36269
rect 40267 36235 40301 36265
rect 40267 36163 40301 36197
rect 41830 37322 41864 37356
rect 41920 37341 41954 37356
rect 42010 37341 42044 37356
rect 42100 37341 42134 37356
rect 42190 37341 42224 37356
rect 42280 37341 42314 37356
rect 42370 37341 42404 37356
rect 42460 37341 42494 37356
rect 42550 37341 42584 37356
rect 42640 37341 42674 37356
rect 42730 37341 42764 37356
rect 42820 37341 42854 37356
rect 42910 37341 42944 37356
rect 41920 37322 41940 37341
rect 41940 37322 41954 37341
rect 42010 37322 42030 37341
rect 42030 37322 42044 37341
rect 42100 37322 42120 37341
rect 42120 37322 42134 37341
rect 42190 37322 42210 37341
rect 42210 37322 42224 37341
rect 42280 37322 42300 37341
rect 42300 37322 42314 37341
rect 42370 37322 42390 37341
rect 42390 37322 42404 37341
rect 42460 37322 42480 37341
rect 42480 37322 42494 37341
rect 42550 37322 42570 37341
rect 42570 37322 42584 37341
rect 42640 37322 42660 37341
rect 42660 37322 42674 37341
rect 42730 37322 42750 37341
rect 42750 37322 42764 37341
rect 42820 37322 42840 37341
rect 42840 37322 42854 37341
rect 42910 37322 42930 37341
rect 42930 37322 42944 37341
rect 43000 37322 43034 37356
rect 43170 37322 43204 37356
rect 43260 37341 43294 37356
rect 43350 37341 43384 37356
rect 43440 37341 43474 37356
rect 43530 37341 43564 37356
rect 43620 37341 43654 37356
rect 43710 37341 43744 37356
rect 43800 37341 43834 37356
rect 43890 37341 43924 37356
rect 43980 37341 44014 37356
rect 44070 37341 44104 37356
rect 44160 37341 44194 37356
rect 44250 37341 44284 37356
rect 43260 37322 43280 37341
rect 43280 37322 43294 37341
rect 43350 37322 43370 37341
rect 43370 37322 43384 37341
rect 43440 37322 43460 37341
rect 43460 37322 43474 37341
rect 43530 37322 43550 37341
rect 43550 37322 43564 37341
rect 43620 37322 43640 37341
rect 43640 37322 43654 37341
rect 43710 37322 43730 37341
rect 43730 37322 43744 37341
rect 43800 37322 43820 37341
rect 43820 37322 43834 37341
rect 43890 37322 43910 37341
rect 43910 37322 43924 37341
rect 43980 37322 44000 37341
rect 44000 37322 44014 37341
rect 44070 37322 44090 37341
rect 44090 37322 44104 37341
rect 44160 37322 44180 37341
rect 44180 37322 44194 37341
rect 44250 37322 44270 37341
rect 44270 37322 44284 37341
rect 44340 37322 44374 37356
rect 44510 37322 44544 37356
rect 44600 37341 44634 37356
rect 44690 37341 44724 37356
rect 44780 37341 44814 37356
rect 44870 37341 44904 37356
rect 44960 37341 44994 37356
rect 45050 37341 45084 37356
rect 45140 37341 45174 37356
rect 45230 37341 45264 37356
rect 45320 37341 45354 37356
rect 45410 37341 45444 37356
rect 45500 37341 45534 37356
rect 45590 37341 45624 37356
rect 44600 37322 44620 37341
rect 44620 37322 44634 37341
rect 44690 37322 44710 37341
rect 44710 37322 44724 37341
rect 44780 37322 44800 37341
rect 44800 37322 44814 37341
rect 44870 37322 44890 37341
rect 44890 37322 44904 37341
rect 44960 37322 44980 37341
rect 44980 37322 44994 37341
rect 45050 37322 45070 37341
rect 45070 37322 45084 37341
rect 45140 37322 45160 37341
rect 45160 37322 45174 37341
rect 45230 37322 45250 37341
rect 45250 37322 45264 37341
rect 45320 37322 45340 37341
rect 45340 37322 45354 37341
rect 45410 37322 45430 37341
rect 45430 37322 45444 37341
rect 45500 37322 45520 37341
rect 45520 37322 45534 37341
rect 45590 37322 45610 37341
rect 45610 37322 45624 37341
rect 45680 37322 45714 37356
rect 45850 37322 45884 37356
rect 45940 37341 45974 37356
rect 46030 37341 46064 37356
rect 46120 37341 46154 37356
rect 46210 37341 46244 37356
rect 46300 37341 46334 37356
rect 46390 37341 46424 37356
rect 46480 37341 46514 37356
rect 46570 37341 46604 37356
rect 46660 37341 46694 37356
rect 46750 37341 46784 37356
rect 46840 37341 46874 37356
rect 46930 37341 46964 37356
rect 45940 37322 45960 37341
rect 45960 37322 45974 37341
rect 46030 37322 46050 37341
rect 46050 37322 46064 37341
rect 46120 37322 46140 37341
rect 46140 37322 46154 37341
rect 46210 37322 46230 37341
rect 46230 37322 46244 37341
rect 46300 37322 46320 37341
rect 46320 37322 46334 37341
rect 46390 37322 46410 37341
rect 46410 37322 46424 37341
rect 46480 37322 46500 37341
rect 46500 37322 46514 37341
rect 46570 37322 46590 37341
rect 46590 37322 46604 37341
rect 46660 37322 46680 37341
rect 46680 37322 46694 37341
rect 46750 37322 46770 37341
rect 46770 37322 46784 37341
rect 46840 37322 46860 37341
rect 46860 37322 46874 37341
rect 46930 37322 46950 37341
rect 46950 37322 46964 37341
rect 47020 37322 47054 37356
rect 47190 37322 47224 37356
rect 47280 37341 47314 37356
rect 47370 37341 47404 37356
rect 47460 37341 47494 37356
rect 47550 37341 47584 37356
rect 47640 37341 47674 37356
rect 47730 37341 47764 37356
rect 47820 37341 47854 37356
rect 47910 37341 47944 37356
rect 48000 37341 48034 37356
rect 48090 37341 48124 37356
rect 48180 37341 48214 37356
rect 48270 37341 48304 37356
rect 47280 37322 47300 37341
rect 47300 37322 47314 37341
rect 47370 37322 47390 37341
rect 47390 37322 47404 37341
rect 47460 37322 47480 37341
rect 47480 37322 47494 37341
rect 47550 37322 47570 37341
rect 47570 37322 47584 37341
rect 47640 37322 47660 37341
rect 47660 37322 47674 37341
rect 47730 37322 47750 37341
rect 47750 37322 47764 37341
rect 47820 37322 47840 37341
rect 47840 37322 47854 37341
rect 47910 37322 47930 37341
rect 47930 37322 47944 37341
rect 48000 37322 48020 37341
rect 48020 37322 48034 37341
rect 48090 37322 48110 37341
rect 48110 37322 48124 37341
rect 48180 37322 48200 37341
rect 48200 37322 48214 37341
rect 48270 37322 48290 37341
rect 48290 37322 48304 37341
rect 48360 37322 48394 37356
rect 48530 37322 48564 37356
rect 48620 37341 48654 37356
rect 48710 37341 48744 37356
rect 48800 37341 48834 37356
rect 48890 37341 48924 37356
rect 48980 37341 49014 37356
rect 49070 37341 49104 37356
rect 49160 37341 49194 37356
rect 49250 37341 49284 37356
rect 49340 37341 49374 37356
rect 49430 37341 49464 37356
rect 49520 37341 49554 37356
rect 49610 37341 49644 37356
rect 48620 37322 48640 37341
rect 48640 37322 48654 37341
rect 48710 37322 48730 37341
rect 48730 37322 48744 37341
rect 48800 37322 48820 37341
rect 48820 37322 48834 37341
rect 48890 37322 48910 37341
rect 48910 37322 48924 37341
rect 48980 37322 49000 37341
rect 49000 37322 49014 37341
rect 49070 37322 49090 37341
rect 49090 37322 49104 37341
rect 49160 37322 49180 37341
rect 49180 37322 49194 37341
rect 49250 37322 49270 37341
rect 49270 37322 49284 37341
rect 49340 37322 49360 37341
rect 49360 37322 49374 37341
rect 49430 37322 49450 37341
rect 49450 37322 49464 37341
rect 49520 37322 49540 37341
rect 49540 37322 49554 37341
rect 49610 37322 49630 37341
rect 49630 37322 49644 37341
rect 49700 37322 49734 37356
rect 49870 37322 49904 37356
rect 49960 37341 49994 37356
rect 50050 37341 50084 37356
rect 50140 37341 50174 37356
rect 50230 37341 50264 37356
rect 50320 37341 50354 37356
rect 50410 37341 50444 37356
rect 50500 37341 50534 37356
rect 50590 37341 50624 37356
rect 50680 37341 50714 37356
rect 50770 37341 50804 37356
rect 50860 37341 50894 37356
rect 50950 37341 50984 37356
rect 49960 37322 49980 37341
rect 49980 37322 49994 37341
rect 50050 37322 50070 37341
rect 50070 37322 50084 37341
rect 50140 37322 50160 37341
rect 50160 37322 50174 37341
rect 50230 37322 50250 37341
rect 50250 37322 50264 37341
rect 50320 37322 50340 37341
rect 50340 37322 50354 37341
rect 50410 37322 50430 37341
rect 50430 37322 50444 37341
rect 50500 37322 50520 37341
rect 50520 37322 50534 37341
rect 50590 37322 50610 37341
rect 50610 37322 50624 37341
rect 50680 37322 50700 37341
rect 50700 37322 50714 37341
rect 50770 37322 50790 37341
rect 50790 37322 50804 37341
rect 50860 37322 50880 37341
rect 50880 37322 50894 37341
rect 50950 37322 50970 37341
rect 50970 37322 50984 37341
rect 51040 37322 51074 37356
rect 51210 37322 51244 37356
rect 51300 37341 51334 37356
rect 51390 37341 51424 37356
rect 51480 37341 51514 37356
rect 51570 37341 51604 37356
rect 51660 37341 51694 37356
rect 51750 37341 51784 37356
rect 51840 37341 51874 37356
rect 51930 37341 51964 37356
rect 52020 37341 52054 37356
rect 52110 37341 52144 37356
rect 52200 37341 52234 37356
rect 52290 37341 52324 37356
rect 51300 37322 51320 37341
rect 51320 37322 51334 37341
rect 51390 37322 51410 37341
rect 51410 37322 51424 37341
rect 51480 37322 51500 37341
rect 51500 37322 51514 37341
rect 51570 37322 51590 37341
rect 51590 37322 51604 37341
rect 51660 37322 51680 37341
rect 51680 37322 51694 37341
rect 51750 37322 51770 37341
rect 51770 37322 51784 37341
rect 51840 37322 51860 37341
rect 51860 37322 51874 37341
rect 51930 37322 51950 37341
rect 51950 37322 51964 37341
rect 52020 37322 52040 37341
rect 52040 37322 52054 37341
rect 52110 37322 52130 37341
rect 52130 37322 52144 37341
rect 52200 37322 52220 37341
rect 52220 37322 52234 37341
rect 52290 37322 52310 37341
rect 52310 37322 52324 37341
rect 52380 37322 52414 37356
rect 41994 37162 42028 37196
rect 42084 37194 42118 37196
rect 42174 37194 42208 37196
rect 42264 37194 42298 37196
rect 42354 37194 42388 37196
rect 42444 37194 42478 37196
rect 42534 37194 42568 37196
rect 42624 37194 42658 37196
rect 42714 37194 42748 37196
rect 42804 37194 42838 37196
rect 42084 37162 42104 37194
rect 42104 37162 42118 37194
rect 42174 37162 42194 37194
rect 42194 37162 42208 37194
rect 42264 37162 42284 37194
rect 42284 37162 42298 37194
rect 42354 37162 42374 37194
rect 42374 37162 42388 37194
rect 42444 37162 42464 37194
rect 42464 37162 42478 37194
rect 42534 37162 42554 37194
rect 42554 37162 42568 37194
rect 42624 37162 42644 37194
rect 42644 37162 42658 37194
rect 42714 37162 42734 37194
rect 42734 37162 42748 37194
rect 42804 37162 42824 37194
rect 42824 37162 42838 37194
rect 42894 37162 42928 37196
rect 42180 36986 42202 36992
rect 42202 36986 42214 36992
rect 42280 36986 42292 36992
rect 42292 36986 42314 36992
rect 42380 36986 42382 36992
rect 42382 36986 42414 36992
rect 42180 36958 42214 36986
rect 42280 36958 42314 36986
rect 42380 36958 42414 36986
rect 42480 36958 42514 36992
rect 42580 36958 42614 36992
rect 42680 36986 42708 36992
rect 42708 36986 42714 36992
rect 42680 36958 42714 36986
rect 42180 36858 42214 36892
rect 42280 36858 42314 36892
rect 42380 36858 42414 36892
rect 42480 36858 42514 36892
rect 42580 36858 42614 36892
rect 42680 36858 42714 36892
rect 42180 36758 42214 36792
rect 42280 36758 42314 36792
rect 42380 36758 42414 36792
rect 42480 36758 42514 36792
rect 42580 36758 42614 36792
rect 42680 36758 42714 36792
rect 42180 36660 42214 36692
rect 42280 36660 42314 36692
rect 42380 36660 42414 36692
rect 42180 36658 42202 36660
rect 42202 36658 42214 36660
rect 42280 36658 42292 36660
rect 42292 36658 42314 36660
rect 42380 36658 42382 36660
rect 42382 36658 42414 36660
rect 42480 36658 42514 36692
rect 42580 36658 42614 36692
rect 42680 36660 42714 36692
rect 42680 36658 42708 36660
rect 42708 36658 42714 36660
rect 42180 36570 42214 36592
rect 42280 36570 42314 36592
rect 42380 36570 42414 36592
rect 42180 36558 42202 36570
rect 42202 36558 42214 36570
rect 42280 36558 42292 36570
rect 42292 36558 42314 36570
rect 42380 36558 42382 36570
rect 42382 36558 42414 36570
rect 42480 36558 42514 36592
rect 42580 36558 42614 36592
rect 42680 36570 42714 36592
rect 42680 36558 42708 36570
rect 42708 36558 42714 36570
rect 42180 36480 42214 36492
rect 42280 36480 42314 36492
rect 42380 36480 42414 36492
rect 42180 36458 42202 36480
rect 42202 36458 42214 36480
rect 42280 36458 42292 36480
rect 42292 36458 42314 36480
rect 42380 36458 42382 36480
rect 42382 36458 42414 36480
rect 42480 36458 42514 36492
rect 42580 36458 42614 36492
rect 42680 36480 42714 36492
rect 42680 36458 42708 36480
rect 42708 36458 42714 36480
rect 43334 37162 43368 37196
rect 43424 37194 43458 37196
rect 43514 37194 43548 37196
rect 43604 37194 43638 37196
rect 43694 37194 43728 37196
rect 43784 37194 43818 37196
rect 43874 37194 43908 37196
rect 43964 37194 43998 37196
rect 44054 37194 44088 37196
rect 44144 37194 44178 37196
rect 43424 37162 43444 37194
rect 43444 37162 43458 37194
rect 43514 37162 43534 37194
rect 43534 37162 43548 37194
rect 43604 37162 43624 37194
rect 43624 37162 43638 37194
rect 43694 37162 43714 37194
rect 43714 37162 43728 37194
rect 43784 37162 43804 37194
rect 43804 37162 43818 37194
rect 43874 37162 43894 37194
rect 43894 37162 43908 37194
rect 43964 37162 43984 37194
rect 43984 37162 43998 37194
rect 44054 37162 44074 37194
rect 44074 37162 44088 37194
rect 44144 37162 44164 37194
rect 44164 37162 44178 37194
rect 44234 37162 44268 37196
rect 43520 36986 43542 36992
rect 43542 36986 43554 36992
rect 43620 36986 43632 36992
rect 43632 36986 43654 36992
rect 43720 36986 43722 36992
rect 43722 36986 43754 36992
rect 43520 36958 43554 36986
rect 43620 36958 43654 36986
rect 43720 36958 43754 36986
rect 43820 36958 43854 36992
rect 43920 36958 43954 36992
rect 44020 36986 44048 36992
rect 44048 36986 44054 36992
rect 44020 36958 44054 36986
rect 43520 36858 43554 36892
rect 43620 36858 43654 36892
rect 43720 36858 43754 36892
rect 43820 36858 43854 36892
rect 43920 36858 43954 36892
rect 44020 36858 44054 36892
rect 43520 36758 43554 36792
rect 43620 36758 43654 36792
rect 43720 36758 43754 36792
rect 43820 36758 43854 36792
rect 43920 36758 43954 36792
rect 44020 36758 44054 36792
rect 43520 36660 43554 36692
rect 43620 36660 43654 36692
rect 43720 36660 43754 36692
rect 43520 36658 43542 36660
rect 43542 36658 43554 36660
rect 43620 36658 43632 36660
rect 43632 36658 43654 36660
rect 43720 36658 43722 36660
rect 43722 36658 43754 36660
rect 43820 36658 43854 36692
rect 43920 36658 43954 36692
rect 44020 36660 44054 36692
rect 44020 36658 44048 36660
rect 44048 36658 44054 36660
rect 43520 36570 43554 36592
rect 43620 36570 43654 36592
rect 43720 36570 43754 36592
rect 43520 36558 43542 36570
rect 43542 36558 43554 36570
rect 43620 36558 43632 36570
rect 43632 36558 43654 36570
rect 43720 36558 43722 36570
rect 43722 36558 43754 36570
rect 43820 36558 43854 36592
rect 43920 36558 43954 36592
rect 44020 36570 44054 36592
rect 44020 36558 44048 36570
rect 44048 36558 44054 36570
rect 43520 36480 43554 36492
rect 43620 36480 43654 36492
rect 43720 36480 43754 36492
rect 43520 36458 43542 36480
rect 43542 36458 43554 36480
rect 43620 36458 43632 36480
rect 43632 36458 43654 36480
rect 43720 36458 43722 36480
rect 43722 36458 43754 36480
rect 43820 36458 43854 36492
rect 43920 36458 43954 36492
rect 44020 36480 44054 36492
rect 44020 36458 44048 36480
rect 44048 36458 44054 36480
rect 44674 37162 44708 37196
rect 44764 37194 44798 37196
rect 44854 37194 44888 37196
rect 44944 37194 44978 37196
rect 45034 37194 45068 37196
rect 45124 37194 45158 37196
rect 45214 37194 45248 37196
rect 45304 37194 45338 37196
rect 45394 37194 45428 37196
rect 45484 37194 45518 37196
rect 44764 37162 44784 37194
rect 44784 37162 44798 37194
rect 44854 37162 44874 37194
rect 44874 37162 44888 37194
rect 44944 37162 44964 37194
rect 44964 37162 44978 37194
rect 45034 37162 45054 37194
rect 45054 37162 45068 37194
rect 45124 37162 45144 37194
rect 45144 37162 45158 37194
rect 45214 37162 45234 37194
rect 45234 37162 45248 37194
rect 45304 37162 45324 37194
rect 45324 37162 45338 37194
rect 45394 37162 45414 37194
rect 45414 37162 45428 37194
rect 45484 37162 45504 37194
rect 45504 37162 45518 37194
rect 45574 37162 45608 37196
rect 44860 36986 44882 36992
rect 44882 36986 44894 36992
rect 44960 36986 44972 36992
rect 44972 36986 44994 36992
rect 45060 36986 45062 36992
rect 45062 36986 45094 36992
rect 44860 36958 44894 36986
rect 44960 36958 44994 36986
rect 45060 36958 45094 36986
rect 45160 36958 45194 36992
rect 45260 36958 45294 36992
rect 45360 36986 45388 36992
rect 45388 36986 45394 36992
rect 45360 36958 45394 36986
rect 44860 36858 44894 36892
rect 44960 36858 44994 36892
rect 45060 36858 45094 36892
rect 45160 36858 45194 36892
rect 45260 36858 45294 36892
rect 45360 36858 45394 36892
rect 44860 36758 44894 36792
rect 44960 36758 44994 36792
rect 45060 36758 45094 36792
rect 45160 36758 45194 36792
rect 45260 36758 45294 36792
rect 45360 36758 45394 36792
rect 44860 36660 44894 36692
rect 44960 36660 44994 36692
rect 45060 36660 45094 36692
rect 44860 36658 44882 36660
rect 44882 36658 44894 36660
rect 44960 36658 44972 36660
rect 44972 36658 44994 36660
rect 45060 36658 45062 36660
rect 45062 36658 45094 36660
rect 45160 36658 45194 36692
rect 45260 36658 45294 36692
rect 45360 36660 45394 36692
rect 45360 36658 45388 36660
rect 45388 36658 45394 36660
rect 44860 36570 44894 36592
rect 44960 36570 44994 36592
rect 45060 36570 45094 36592
rect 44860 36558 44882 36570
rect 44882 36558 44894 36570
rect 44960 36558 44972 36570
rect 44972 36558 44994 36570
rect 45060 36558 45062 36570
rect 45062 36558 45094 36570
rect 45160 36558 45194 36592
rect 45260 36558 45294 36592
rect 45360 36570 45394 36592
rect 45360 36558 45388 36570
rect 45388 36558 45394 36570
rect 44860 36480 44894 36492
rect 44960 36480 44994 36492
rect 45060 36480 45094 36492
rect 44860 36458 44882 36480
rect 44882 36458 44894 36480
rect 44960 36458 44972 36480
rect 44972 36458 44994 36480
rect 45060 36458 45062 36480
rect 45062 36458 45094 36480
rect 45160 36458 45194 36492
rect 45260 36458 45294 36492
rect 45360 36480 45394 36492
rect 45360 36458 45388 36480
rect 45388 36458 45394 36480
rect 46014 37162 46048 37196
rect 46104 37194 46138 37196
rect 46194 37194 46228 37196
rect 46284 37194 46318 37196
rect 46374 37194 46408 37196
rect 46464 37194 46498 37196
rect 46554 37194 46588 37196
rect 46644 37194 46678 37196
rect 46734 37194 46768 37196
rect 46824 37194 46858 37196
rect 46104 37162 46124 37194
rect 46124 37162 46138 37194
rect 46194 37162 46214 37194
rect 46214 37162 46228 37194
rect 46284 37162 46304 37194
rect 46304 37162 46318 37194
rect 46374 37162 46394 37194
rect 46394 37162 46408 37194
rect 46464 37162 46484 37194
rect 46484 37162 46498 37194
rect 46554 37162 46574 37194
rect 46574 37162 46588 37194
rect 46644 37162 46664 37194
rect 46664 37162 46678 37194
rect 46734 37162 46754 37194
rect 46754 37162 46768 37194
rect 46824 37162 46844 37194
rect 46844 37162 46858 37194
rect 46914 37162 46948 37196
rect 46200 36986 46222 36992
rect 46222 36986 46234 36992
rect 46300 36986 46312 36992
rect 46312 36986 46334 36992
rect 46400 36986 46402 36992
rect 46402 36986 46434 36992
rect 46200 36958 46234 36986
rect 46300 36958 46334 36986
rect 46400 36958 46434 36986
rect 46500 36958 46534 36992
rect 46600 36958 46634 36992
rect 46700 36986 46728 36992
rect 46728 36986 46734 36992
rect 46700 36958 46734 36986
rect 46200 36858 46234 36892
rect 46300 36858 46334 36892
rect 46400 36858 46434 36892
rect 46500 36858 46534 36892
rect 46600 36858 46634 36892
rect 46700 36858 46734 36892
rect 46200 36758 46234 36792
rect 46300 36758 46334 36792
rect 46400 36758 46434 36792
rect 46500 36758 46534 36792
rect 46600 36758 46634 36792
rect 46700 36758 46734 36792
rect 46200 36660 46234 36692
rect 46300 36660 46334 36692
rect 46400 36660 46434 36692
rect 46200 36658 46222 36660
rect 46222 36658 46234 36660
rect 46300 36658 46312 36660
rect 46312 36658 46334 36660
rect 46400 36658 46402 36660
rect 46402 36658 46434 36660
rect 46500 36658 46534 36692
rect 46600 36658 46634 36692
rect 46700 36660 46734 36692
rect 46700 36658 46728 36660
rect 46728 36658 46734 36660
rect 46200 36570 46234 36592
rect 46300 36570 46334 36592
rect 46400 36570 46434 36592
rect 46200 36558 46222 36570
rect 46222 36558 46234 36570
rect 46300 36558 46312 36570
rect 46312 36558 46334 36570
rect 46400 36558 46402 36570
rect 46402 36558 46434 36570
rect 46500 36558 46534 36592
rect 46600 36558 46634 36592
rect 46700 36570 46734 36592
rect 46700 36558 46728 36570
rect 46728 36558 46734 36570
rect 46200 36480 46234 36492
rect 46300 36480 46334 36492
rect 46400 36480 46434 36492
rect 46200 36458 46222 36480
rect 46222 36458 46234 36480
rect 46300 36458 46312 36480
rect 46312 36458 46334 36480
rect 46400 36458 46402 36480
rect 46402 36458 46434 36480
rect 46500 36458 46534 36492
rect 46600 36458 46634 36492
rect 46700 36480 46734 36492
rect 46700 36458 46728 36480
rect 46728 36458 46734 36480
rect 47354 37162 47388 37196
rect 47444 37194 47478 37196
rect 47534 37194 47568 37196
rect 47624 37194 47658 37196
rect 47714 37194 47748 37196
rect 47804 37194 47838 37196
rect 47894 37194 47928 37196
rect 47984 37194 48018 37196
rect 48074 37194 48108 37196
rect 48164 37194 48198 37196
rect 47444 37162 47464 37194
rect 47464 37162 47478 37194
rect 47534 37162 47554 37194
rect 47554 37162 47568 37194
rect 47624 37162 47644 37194
rect 47644 37162 47658 37194
rect 47714 37162 47734 37194
rect 47734 37162 47748 37194
rect 47804 37162 47824 37194
rect 47824 37162 47838 37194
rect 47894 37162 47914 37194
rect 47914 37162 47928 37194
rect 47984 37162 48004 37194
rect 48004 37162 48018 37194
rect 48074 37162 48094 37194
rect 48094 37162 48108 37194
rect 48164 37162 48184 37194
rect 48184 37162 48198 37194
rect 48254 37162 48288 37196
rect 47540 36986 47562 36992
rect 47562 36986 47574 36992
rect 47640 36986 47652 36992
rect 47652 36986 47674 36992
rect 47740 36986 47742 36992
rect 47742 36986 47774 36992
rect 47540 36958 47574 36986
rect 47640 36958 47674 36986
rect 47740 36958 47774 36986
rect 47840 36958 47874 36992
rect 47940 36958 47974 36992
rect 48040 36986 48068 36992
rect 48068 36986 48074 36992
rect 48040 36958 48074 36986
rect 47540 36858 47574 36892
rect 47640 36858 47674 36892
rect 47740 36858 47774 36892
rect 47840 36858 47874 36892
rect 47940 36858 47974 36892
rect 48040 36858 48074 36892
rect 47540 36758 47574 36792
rect 47640 36758 47674 36792
rect 47740 36758 47774 36792
rect 47840 36758 47874 36792
rect 47940 36758 47974 36792
rect 48040 36758 48074 36792
rect 47540 36660 47574 36692
rect 47640 36660 47674 36692
rect 47740 36660 47774 36692
rect 47540 36658 47562 36660
rect 47562 36658 47574 36660
rect 47640 36658 47652 36660
rect 47652 36658 47674 36660
rect 47740 36658 47742 36660
rect 47742 36658 47774 36660
rect 47840 36658 47874 36692
rect 47940 36658 47974 36692
rect 48040 36660 48074 36692
rect 48040 36658 48068 36660
rect 48068 36658 48074 36660
rect 47540 36570 47574 36592
rect 47640 36570 47674 36592
rect 47740 36570 47774 36592
rect 47540 36558 47562 36570
rect 47562 36558 47574 36570
rect 47640 36558 47652 36570
rect 47652 36558 47674 36570
rect 47740 36558 47742 36570
rect 47742 36558 47774 36570
rect 47840 36558 47874 36592
rect 47940 36558 47974 36592
rect 48040 36570 48074 36592
rect 48040 36558 48068 36570
rect 48068 36558 48074 36570
rect 47540 36480 47574 36492
rect 47640 36480 47674 36492
rect 47740 36480 47774 36492
rect 47540 36458 47562 36480
rect 47562 36458 47574 36480
rect 47640 36458 47652 36480
rect 47652 36458 47674 36480
rect 47740 36458 47742 36480
rect 47742 36458 47774 36480
rect 47840 36458 47874 36492
rect 47940 36458 47974 36492
rect 48040 36480 48074 36492
rect 48040 36458 48068 36480
rect 48068 36458 48074 36480
rect 48694 37162 48728 37196
rect 48784 37194 48818 37196
rect 48874 37194 48908 37196
rect 48964 37194 48998 37196
rect 49054 37194 49088 37196
rect 49144 37194 49178 37196
rect 49234 37194 49268 37196
rect 49324 37194 49358 37196
rect 49414 37194 49448 37196
rect 49504 37194 49538 37196
rect 48784 37162 48804 37194
rect 48804 37162 48818 37194
rect 48874 37162 48894 37194
rect 48894 37162 48908 37194
rect 48964 37162 48984 37194
rect 48984 37162 48998 37194
rect 49054 37162 49074 37194
rect 49074 37162 49088 37194
rect 49144 37162 49164 37194
rect 49164 37162 49178 37194
rect 49234 37162 49254 37194
rect 49254 37162 49268 37194
rect 49324 37162 49344 37194
rect 49344 37162 49358 37194
rect 49414 37162 49434 37194
rect 49434 37162 49448 37194
rect 49504 37162 49524 37194
rect 49524 37162 49538 37194
rect 49594 37162 49628 37196
rect 48880 36986 48902 36992
rect 48902 36986 48914 36992
rect 48980 36986 48992 36992
rect 48992 36986 49014 36992
rect 49080 36986 49082 36992
rect 49082 36986 49114 36992
rect 48880 36958 48914 36986
rect 48980 36958 49014 36986
rect 49080 36958 49114 36986
rect 49180 36958 49214 36992
rect 49280 36958 49314 36992
rect 49380 36986 49408 36992
rect 49408 36986 49414 36992
rect 49380 36958 49414 36986
rect 48880 36858 48914 36892
rect 48980 36858 49014 36892
rect 49080 36858 49114 36892
rect 49180 36858 49214 36892
rect 49280 36858 49314 36892
rect 49380 36858 49414 36892
rect 48880 36758 48914 36792
rect 48980 36758 49014 36792
rect 49080 36758 49114 36792
rect 49180 36758 49214 36792
rect 49280 36758 49314 36792
rect 49380 36758 49414 36792
rect 48880 36660 48914 36692
rect 48980 36660 49014 36692
rect 49080 36660 49114 36692
rect 48880 36658 48902 36660
rect 48902 36658 48914 36660
rect 48980 36658 48992 36660
rect 48992 36658 49014 36660
rect 49080 36658 49082 36660
rect 49082 36658 49114 36660
rect 49180 36658 49214 36692
rect 49280 36658 49314 36692
rect 49380 36660 49414 36692
rect 49380 36658 49408 36660
rect 49408 36658 49414 36660
rect 48880 36570 48914 36592
rect 48980 36570 49014 36592
rect 49080 36570 49114 36592
rect 48880 36558 48902 36570
rect 48902 36558 48914 36570
rect 48980 36558 48992 36570
rect 48992 36558 49014 36570
rect 49080 36558 49082 36570
rect 49082 36558 49114 36570
rect 49180 36558 49214 36592
rect 49280 36558 49314 36592
rect 49380 36570 49414 36592
rect 49380 36558 49408 36570
rect 49408 36558 49414 36570
rect 48880 36480 48914 36492
rect 48980 36480 49014 36492
rect 49080 36480 49114 36492
rect 48880 36458 48902 36480
rect 48902 36458 48914 36480
rect 48980 36458 48992 36480
rect 48992 36458 49014 36480
rect 49080 36458 49082 36480
rect 49082 36458 49114 36480
rect 49180 36458 49214 36492
rect 49280 36458 49314 36492
rect 49380 36480 49414 36492
rect 49380 36458 49408 36480
rect 49408 36458 49414 36480
rect 50034 37162 50068 37196
rect 50124 37194 50158 37196
rect 50214 37194 50248 37196
rect 50304 37194 50338 37196
rect 50394 37194 50428 37196
rect 50484 37194 50518 37196
rect 50574 37194 50608 37196
rect 50664 37194 50698 37196
rect 50754 37194 50788 37196
rect 50844 37194 50878 37196
rect 50124 37162 50144 37194
rect 50144 37162 50158 37194
rect 50214 37162 50234 37194
rect 50234 37162 50248 37194
rect 50304 37162 50324 37194
rect 50324 37162 50338 37194
rect 50394 37162 50414 37194
rect 50414 37162 50428 37194
rect 50484 37162 50504 37194
rect 50504 37162 50518 37194
rect 50574 37162 50594 37194
rect 50594 37162 50608 37194
rect 50664 37162 50684 37194
rect 50684 37162 50698 37194
rect 50754 37162 50774 37194
rect 50774 37162 50788 37194
rect 50844 37162 50864 37194
rect 50864 37162 50878 37194
rect 50934 37162 50968 37196
rect 50220 36986 50242 36992
rect 50242 36986 50254 36992
rect 50320 36986 50332 36992
rect 50332 36986 50354 36992
rect 50420 36986 50422 36992
rect 50422 36986 50454 36992
rect 50220 36958 50254 36986
rect 50320 36958 50354 36986
rect 50420 36958 50454 36986
rect 50520 36958 50554 36992
rect 50620 36958 50654 36992
rect 50720 36986 50748 36992
rect 50748 36986 50754 36992
rect 50720 36958 50754 36986
rect 50220 36858 50254 36892
rect 50320 36858 50354 36892
rect 50420 36858 50454 36892
rect 50520 36858 50554 36892
rect 50620 36858 50654 36892
rect 50720 36858 50754 36892
rect 50220 36758 50254 36792
rect 50320 36758 50354 36792
rect 50420 36758 50454 36792
rect 50520 36758 50554 36792
rect 50620 36758 50654 36792
rect 50720 36758 50754 36792
rect 50220 36660 50254 36692
rect 50320 36660 50354 36692
rect 50420 36660 50454 36692
rect 50220 36658 50242 36660
rect 50242 36658 50254 36660
rect 50320 36658 50332 36660
rect 50332 36658 50354 36660
rect 50420 36658 50422 36660
rect 50422 36658 50454 36660
rect 50520 36658 50554 36692
rect 50620 36658 50654 36692
rect 50720 36660 50754 36692
rect 50720 36658 50748 36660
rect 50748 36658 50754 36660
rect 50220 36570 50254 36592
rect 50320 36570 50354 36592
rect 50420 36570 50454 36592
rect 50220 36558 50242 36570
rect 50242 36558 50254 36570
rect 50320 36558 50332 36570
rect 50332 36558 50354 36570
rect 50420 36558 50422 36570
rect 50422 36558 50454 36570
rect 50520 36558 50554 36592
rect 50620 36558 50654 36592
rect 50720 36570 50754 36592
rect 50720 36558 50748 36570
rect 50748 36558 50754 36570
rect 50220 36480 50254 36492
rect 50320 36480 50354 36492
rect 50420 36480 50454 36492
rect 50220 36458 50242 36480
rect 50242 36458 50254 36480
rect 50320 36458 50332 36480
rect 50332 36458 50354 36480
rect 50420 36458 50422 36480
rect 50422 36458 50454 36480
rect 50520 36458 50554 36492
rect 50620 36458 50654 36492
rect 50720 36480 50754 36492
rect 50720 36458 50748 36480
rect 50748 36458 50754 36480
rect 51374 37162 51408 37196
rect 51464 37194 51498 37196
rect 51554 37194 51588 37196
rect 51644 37194 51678 37196
rect 51734 37194 51768 37196
rect 51824 37194 51858 37196
rect 51914 37194 51948 37196
rect 52004 37194 52038 37196
rect 52094 37194 52128 37196
rect 52184 37194 52218 37196
rect 51464 37162 51484 37194
rect 51484 37162 51498 37194
rect 51554 37162 51574 37194
rect 51574 37162 51588 37194
rect 51644 37162 51664 37194
rect 51664 37162 51678 37194
rect 51734 37162 51754 37194
rect 51754 37162 51768 37194
rect 51824 37162 51844 37194
rect 51844 37162 51858 37194
rect 51914 37162 51934 37194
rect 51934 37162 51948 37194
rect 52004 37162 52024 37194
rect 52024 37162 52038 37194
rect 52094 37162 52114 37194
rect 52114 37162 52128 37194
rect 52184 37162 52204 37194
rect 52204 37162 52218 37194
rect 52274 37162 52308 37196
rect 51560 36986 51582 36992
rect 51582 36986 51594 36992
rect 51660 36986 51672 36992
rect 51672 36986 51694 36992
rect 51760 36986 51762 36992
rect 51762 36986 51794 36992
rect 51560 36958 51594 36986
rect 51660 36958 51694 36986
rect 51760 36958 51794 36986
rect 51860 36958 51894 36992
rect 51960 36958 51994 36992
rect 52060 36986 52088 36992
rect 52088 36986 52094 36992
rect 52060 36958 52094 36986
rect 51560 36858 51594 36892
rect 51660 36858 51694 36892
rect 51760 36858 51794 36892
rect 51860 36858 51894 36892
rect 51960 36858 51994 36892
rect 52060 36858 52094 36892
rect 51560 36758 51594 36792
rect 51660 36758 51694 36792
rect 51760 36758 51794 36792
rect 51860 36758 51894 36792
rect 51960 36758 51994 36792
rect 52060 36758 52094 36792
rect 51560 36660 51594 36692
rect 51660 36660 51694 36692
rect 51760 36660 51794 36692
rect 51560 36658 51582 36660
rect 51582 36658 51594 36660
rect 51660 36658 51672 36660
rect 51672 36658 51694 36660
rect 51760 36658 51762 36660
rect 51762 36658 51794 36660
rect 51860 36658 51894 36692
rect 51960 36658 51994 36692
rect 52060 36660 52094 36692
rect 52060 36658 52088 36660
rect 52088 36658 52094 36660
rect 51560 36570 51594 36592
rect 51660 36570 51694 36592
rect 51760 36570 51794 36592
rect 51560 36558 51582 36570
rect 51582 36558 51594 36570
rect 51660 36558 51672 36570
rect 51672 36558 51694 36570
rect 51760 36558 51762 36570
rect 51762 36558 51794 36570
rect 51860 36558 51894 36592
rect 51960 36558 51994 36592
rect 52060 36570 52094 36592
rect 52060 36558 52088 36570
rect 52088 36558 52094 36570
rect 51560 36480 51594 36492
rect 51660 36480 51694 36492
rect 51760 36480 51794 36492
rect 51560 36458 51582 36480
rect 51582 36458 51594 36480
rect 51660 36458 51672 36480
rect 51672 36458 51694 36480
rect 51760 36458 51762 36480
rect 51762 36458 51794 36480
rect 51860 36458 51894 36492
rect 51960 36458 51994 36492
rect 52060 36480 52094 36492
rect 52060 36458 52088 36480
rect 52088 36458 52094 36480
rect 37565 36023 37599 36057
rect 38577 35921 38611 35955
rect 12175 35775 12209 35809
rect 12375 35775 12409 35809
rect 12575 35775 12609 35809
rect 12775 35775 12809 35809
rect 12975 35775 13009 35809
rect 13175 35775 13209 35809
rect 13861 35775 13895 35809
rect 14061 35775 14095 35809
rect 14261 35775 14295 35809
rect 14461 35775 14495 35809
rect 14661 35775 14695 35809
rect 14861 35775 14895 35809
rect 15061 35775 15095 35809
rect 15261 35775 15295 35809
rect 15461 35775 15495 35809
rect 15661 35775 15695 35809
rect 15861 35775 15895 35809
rect 16605 35775 16639 35809
rect 16805 35775 16839 35809
rect 17005 35775 17039 35809
rect 17205 35775 17239 35809
rect 17405 35775 17439 35809
rect 17605 35775 17639 35809
rect 17805 35775 17839 35809
rect 18005 35775 18039 35809
rect 18205 35775 18239 35809
rect 18405 35775 18439 35809
rect 18605 35775 18639 35809
rect 19351 35775 19385 35809
rect 19551 35775 19585 35809
rect 19751 35775 19785 35809
rect 19951 35775 19985 35809
rect 20151 35775 20185 35809
rect 20351 35775 20385 35809
rect 20551 35775 20585 35809
rect 20751 35775 20785 35809
rect 20951 35775 20985 35809
rect 21151 35775 21185 35809
rect 21351 35775 21385 35809
rect 21551 35775 21585 35809
rect 21751 35775 21785 35809
rect 21951 35775 21985 35809
rect 22681 35775 22715 35809
rect 22881 35775 22915 35809
rect 23081 35775 23115 35809
rect 23281 35775 23315 35809
rect 23481 35775 23515 35809
rect 23681 35775 23715 35809
rect 23881 35775 23915 35809
rect 24081 35775 24115 35809
rect 24281 35775 24315 35809
rect 24481 35775 24515 35809
rect 24681 35775 24715 35809
rect 25601 35775 25635 35809
rect 26001 35775 26035 35809
rect 26401 35775 26435 35809
rect 26801 35775 26835 35809
rect 27201 35775 27235 35809
rect 27601 35775 27635 35809
rect 28001 35775 28035 35809
rect 28401 35775 28435 35809
rect 28801 35775 28835 35809
rect 29201 35775 29235 35809
rect 30111 35775 30145 35809
rect 30511 35775 30545 35809
rect 30911 35775 30945 35809
rect 31311 35775 31345 35809
rect 31711 35775 31745 35809
rect 32111 35775 32145 35809
rect 32511 35775 32545 35809
rect 32911 35775 32945 35809
rect 33311 35775 33345 35809
rect 33711 35775 33745 35809
rect 34111 35775 34145 35809
rect 34511 35775 34545 35809
rect 34911 35775 34945 35809
rect 35311 35775 35345 35809
rect 35711 35775 35745 35809
rect 36111 35775 36145 35809
rect 36511 35775 36545 35809
rect 36911 35775 36945 35809
rect 37655 35775 37689 35809
rect 38055 35775 38089 35809
rect 38455 35775 38489 35809
rect 38855 35775 38889 35809
rect 39255 35775 39289 35809
rect 39655 35775 39689 35809
rect 40055 35775 40089 35809
rect 41967 35775 42001 35809
rect 42167 35775 42201 35809
rect 42367 35775 42401 35809
rect 42567 35775 42601 35809
rect 42767 35775 42801 35809
rect 42967 35775 43001 35809
rect 43167 35775 43201 35809
rect 43367 35775 43401 35809
rect 43567 35775 43601 35809
rect 43767 35775 43801 35809
rect 43967 35775 44001 35809
rect 44167 35775 44201 35809
rect 44367 35775 44401 35809
rect 44567 35775 44601 35809
rect 44767 35775 44801 35809
rect 44967 35775 45001 35809
rect 45167 35775 45201 35809
rect 45367 35775 45401 35809
rect 45567 35775 45601 35809
rect 45767 35775 45801 35809
rect 45967 35775 46001 35809
rect 46167 35775 46201 35809
rect 46367 35775 46401 35809
rect 46567 35775 46601 35809
rect 46767 35775 46801 35809
rect 46967 35775 47001 35809
rect 47167 35775 47201 35809
rect 47367 35775 47401 35809
rect 47567 35775 47601 35809
rect 47767 35775 47801 35809
rect 47967 35775 48001 35809
rect 48167 35775 48201 35809
rect 48367 35775 48401 35809
rect 48567 35775 48601 35809
rect 48767 35775 48801 35809
rect 48967 35775 49001 35809
rect 49167 35775 49201 35809
rect 49367 35775 49401 35809
rect 49567 35775 49601 35809
rect 49767 35775 49801 35809
rect 49967 35775 50001 35809
rect 50167 35775 50201 35809
rect 50367 35775 50401 35809
rect 50567 35775 50601 35809
rect 50767 35775 50801 35809
rect 50967 35775 51001 35809
rect 51167 35775 51201 35809
rect 51367 35775 51401 35809
rect 51567 35775 51601 35809
rect 51767 35775 51801 35809
rect 51967 35775 52001 35809
rect 52167 35775 52201 35809
rect 52367 35775 52401 35809
rect 19447 33895 19481 33929
rect 19647 33895 19681 33929
rect 19847 33895 19881 33929
rect 20047 33895 20081 33929
rect 20247 33895 20281 33929
rect 20447 33895 20481 33929
rect 20647 33895 20681 33929
rect 20847 33895 20881 33929
rect 21047 33895 21081 33929
rect 21247 33895 21281 33929
rect 21447 33895 21481 33929
rect 22193 33895 22227 33929
rect 22393 33895 22427 33929
rect 22593 33895 22627 33929
rect 22793 33895 22827 33929
rect 22993 33895 23027 33929
rect 23193 33895 23227 33929
rect 23393 33895 23427 33929
rect 23593 33895 23627 33929
rect 23793 33895 23827 33929
rect 23993 33895 24027 33929
rect 24193 33895 24227 33929
rect 24393 33895 24427 33929
rect 24593 33895 24627 33929
rect 24793 33895 24827 33929
rect 26387 33895 26421 33929
rect 26787 33895 26821 33929
rect 27187 33895 27221 33929
rect 27587 33895 27621 33929
rect 27987 33895 28021 33929
rect 28387 33895 28421 33929
rect 28787 33895 28821 33929
rect 29187 33895 29221 33929
rect 29587 33895 29621 33929
rect 29987 33895 30021 33929
rect 30387 33895 30421 33929
rect 30787 33895 30821 33929
rect 31187 33895 31221 33929
rect 31587 33895 31621 33929
rect 31987 33895 32021 33929
rect 32387 33895 32421 33929
rect 32787 33895 32821 33929
rect 33187 33895 33221 33929
rect 33835 33895 33869 33929
rect 34235 33895 34269 33929
rect 34635 33895 34669 33929
rect 35035 33895 35069 33929
rect 35435 33895 35469 33929
rect 35835 33895 35869 33929
rect 36235 33895 36269 33929
rect 36635 33895 36669 33929
rect 37035 33895 37069 33929
rect 37435 33895 37469 33929
rect 37835 33895 37869 33929
rect 38235 33895 38269 33929
rect 38635 33895 38669 33929
rect 39035 33895 39069 33929
rect 39435 33895 39469 33929
rect 39835 33895 39869 33929
rect 40235 33895 40269 33929
rect 40635 33895 40669 33929
rect 41967 33895 42001 33929
rect 42167 33895 42201 33929
rect 42367 33895 42401 33929
rect 42567 33895 42601 33929
rect 42767 33895 42801 33929
rect 42967 33895 43001 33929
rect 43167 33895 43201 33929
rect 43367 33895 43401 33929
rect 43567 33895 43601 33929
rect 43767 33895 43801 33929
rect 43967 33895 44001 33929
rect 44167 33895 44201 33929
rect 44367 33895 44401 33929
rect 44567 33895 44601 33929
rect 44767 33895 44801 33929
rect 44967 33895 45001 33929
rect 45167 33895 45201 33929
rect 45367 33895 45401 33929
rect 45567 33895 45601 33929
rect 45767 33895 45801 33929
rect 45967 33895 46001 33929
rect 46167 33895 46201 33929
rect 46367 33895 46401 33929
rect 46567 33895 46601 33929
rect 46767 33895 46801 33929
rect 46967 33895 47001 33929
rect 47167 33895 47201 33929
rect 47367 33895 47401 33929
rect 47567 33895 47601 33929
rect 47767 33895 47801 33929
rect 47967 33895 48001 33929
rect 48167 33895 48201 33929
rect 48367 33895 48401 33929
rect 48567 33895 48601 33929
rect 48767 33895 48801 33929
rect 48967 33895 49001 33929
rect 49167 33895 49201 33929
rect 49367 33895 49401 33929
rect 49567 33895 49601 33929
rect 49767 33895 49801 33929
rect 49967 33895 50001 33929
rect 50167 33895 50201 33929
rect 50367 33895 50401 33929
rect 50567 33895 50601 33929
rect 50767 33895 50801 33929
rect 50967 33895 51001 33929
rect 51167 33895 51201 33929
rect 51367 33895 51401 33929
rect 51567 33895 51601 33929
rect 51767 33895 51801 33929
rect 51967 33895 52001 33929
rect 52167 33895 52201 33929
rect 52367 33895 52401 33929
rect 19283 33123 19677 33661
rect 21290 33123 21684 33661
rect 22028 33123 22422 33661
rect 24609 33123 25003 33661
rect 19283 32163 19677 32701
rect 21290 32163 21684 32701
rect 22028 32163 22422 32701
rect 24609 32163 25003 32701
rect 41830 33562 41864 33596
rect 41920 33581 41954 33596
rect 42010 33581 42044 33596
rect 42100 33581 42134 33596
rect 42190 33581 42224 33596
rect 42280 33581 42314 33596
rect 42370 33581 42404 33596
rect 42460 33581 42494 33596
rect 42550 33581 42584 33596
rect 42640 33581 42674 33596
rect 42730 33581 42764 33596
rect 42820 33581 42854 33596
rect 42910 33581 42944 33596
rect 41920 33562 41940 33581
rect 41940 33562 41954 33581
rect 42010 33562 42030 33581
rect 42030 33562 42044 33581
rect 42100 33562 42120 33581
rect 42120 33562 42134 33581
rect 42190 33562 42210 33581
rect 42210 33562 42224 33581
rect 42280 33562 42300 33581
rect 42300 33562 42314 33581
rect 42370 33562 42390 33581
rect 42390 33562 42404 33581
rect 42460 33562 42480 33581
rect 42480 33562 42494 33581
rect 42550 33562 42570 33581
rect 42570 33562 42584 33581
rect 42640 33562 42660 33581
rect 42660 33562 42674 33581
rect 42730 33562 42750 33581
rect 42750 33562 42764 33581
rect 42820 33562 42840 33581
rect 42840 33562 42854 33581
rect 42910 33562 42930 33581
rect 42930 33562 42944 33581
rect 43000 33562 43034 33596
rect 43170 33562 43204 33596
rect 43260 33581 43294 33596
rect 43350 33581 43384 33596
rect 43440 33581 43474 33596
rect 43530 33581 43564 33596
rect 43620 33581 43654 33596
rect 43710 33581 43744 33596
rect 43800 33581 43834 33596
rect 43890 33581 43924 33596
rect 43980 33581 44014 33596
rect 44070 33581 44104 33596
rect 44160 33581 44194 33596
rect 44250 33581 44284 33596
rect 43260 33562 43280 33581
rect 43280 33562 43294 33581
rect 43350 33562 43370 33581
rect 43370 33562 43384 33581
rect 43440 33562 43460 33581
rect 43460 33562 43474 33581
rect 43530 33562 43550 33581
rect 43550 33562 43564 33581
rect 43620 33562 43640 33581
rect 43640 33562 43654 33581
rect 43710 33562 43730 33581
rect 43730 33562 43744 33581
rect 43800 33562 43820 33581
rect 43820 33562 43834 33581
rect 43890 33562 43910 33581
rect 43910 33562 43924 33581
rect 43980 33562 44000 33581
rect 44000 33562 44014 33581
rect 44070 33562 44090 33581
rect 44090 33562 44104 33581
rect 44160 33562 44180 33581
rect 44180 33562 44194 33581
rect 44250 33562 44270 33581
rect 44270 33562 44284 33581
rect 44340 33562 44374 33596
rect 44510 33562 44544 33596
rect 44600 33581 44634 33596
rect 44690 33581 44724 33596
rect 44780 33581 44814 33596
rect 44870 33581 44904 33596
rect 44960 33581 44994 33596
rect 45050 33581 45084 33596
rect 45140 33581 45174 33596
rect 45230 33581 45264 33596
rect 45320 33581 45354 33596
rect 45410 33581 45444 33596
rect 45500 33581 45534 33596
rect 45590 33581 45624 33596
rect 44600 33562 44620 33581
rect 44620 33562 44634 33581
rect 44690 33562 44710 33581
rect 44710 33562 44724 33581
rect 44780 33562 44800 33581
rect 44800 33562 44814 33581
rect 44870 33562 44890 33581
rect 44890 33562 44904 33581
rect 44960 33562 44980 33581
rect 44980 33562 44994 33581
rect 45050 33562 45070 33581
rect 45070 33562 45084 33581
rect 45140 33562 45160 33581
rect 45160 33562 45174 33581
rect 45230 33562 45250 33581
rect 45250 33562 45264 33581
rect 45320 33562 45340 33581
rect 45340 33562 45354 33581
rect 45410 33562 45430 33581
rect 45430 33562 45444 33581
rect 45500 33562 45520 33581
rect 45520 33562 45534 33581
rect 45590 33562 45610 33581
rect 45610 33562 45624 33581
rect 45680 33562 45714 33596
rect 45850 33562 45884 33596
rect 45940 33581 45974 33596
rect 46030 33581 46064 33596
rect 46120 33581 46154 33596
rect 46210 33581 46244 33596
rect 46300 33581 46334 33596
rect 46390 33581 46424 33596
rect 46480 33581 46514 33596
rect 46570 33581 46604 33596
rect 46660 33581 46694 33596
rect 46750 33581 46784 33596
rect 46840 33581 46874 33596
rect 46930 33581 46964 33596
rect 45940 33562 45960 33581
rect 45960 33562 45974 33581
rect 46030 33562 46050 33581
rect 46050 33562 46064 33581
rect 46120 33562 46140 33581
rect 46140 33562 46154 33581
rect 46210 33562 46230 33581
rect 46230 33562 46244 33581
rect 46300 33562 46320 33581
rect 46320 33562 46334 33581
rect 46390 33562 46410 33581
rect 46410 33562 46424 33581
rect 46480 33562 46500 33581
rect 46500 33562 46514 33581
rect 46570 33562 46590 33581
rect 46590 33562 46604 33581
rect 46660 33562 46680 33581
rect 46680 33562 46694 33581
rect 46750 33562 46770 33581
rect 46770 33562 46784 33581
rect 46840 33562 46860 33581
rect 46860 33562 46874 33581
rect 46930 33562 46950 33581
rect 46950 33562 46964 33581
rect 47020 33562 47054 33596
rect 47190 33562 47224 33596
rect 47280 33581 47314 33596
rect 47370 33581 47404 33596
rect 47460 33581 47494 33596
rect 47550 33581 47584 33596
rect 47640 33581 47674 33596
rect 47730 33581 47764 33596
rect 47820 33581 47854 33596
rect 47910 33581 47944 33596
rect 48000 33581 48034 33596
rect 48090 33581 48124 33596
rect 48180 33581 48214 33596
rect 48270 33581 48304 33596
rect 47280 33562 47300 33581
rect 47300 33562 47314 33581
rect 47370 33562 47390 33581
rect 47390 33562 47404 33581
rect 47460 33562 47480 33581
rect 47480 33562 47494 33581
rect 47550 33562 47570 33581
rect 47570 33562 47584 33581
rect 47640 33562 47660 33581
rect 47660 33562 47674 33581
rect 47730 33562 47750 33581
rect 47750 33562 47764 33581
rect 47820 33562 47840 33581
rect 47840 33562 47854 33581
rect 47910 33562 47930 33581
rect 47930 33562 47944 33581
rect 48000 33562 48020 33581
rect 48020 33562 48034 33581
rect 48090 33562 48110 33581
rect 48110 33562 48124 33581
rect 48180 33562 48200 33581
rect 48200 33562 48214 33581
rect 48270 33562 48290 33581
rect 48290 33562 48304 33581
rect 48360 33562 48394 33596
rect 48530 33562 48564 33596
rect 48620 33581 48654 33596
rect 48710 33581 48744 33596
rect 48800 33581 48834 33596
rect 48890 33581 48924 33596
rect 48980 33581 49014 33596
rect 49070 33581 49104 33596
rect 49160 33581 49194 33596
rect 49250 33581 49284 33596
rect 49340 33581 49374 33596
rect 49430 33581 49464 33596
rect 49520 33581 49554 33596
rect 49610 33581 49644 33596
rect 48620 33562 48640 33581
rect 48640 33562 48654 33581
rect 48710 33562 48730 33581
rect 48730 33562 48744 33581
rect 48800 33562 48820 33581
rect 48820 33562 48834 33581
rect 48890 33562 48910 33581
rect 48910 33562 48924 33581
rect 48980 33562 49000 33581
rect 49000 33562 49014 33581
rect 49070 33562 49090 33581
rect 49090 33562 49104 33581
rect 49160 33562 49180 33581
rect 49180 33562 49194 33581
rect 49250 33562 49270 33581
rect 49270 33562 49284 33581
rect 49340 33562 49360 33581
rect 49360 33562 49374 33581
rect 49430 33562 49450 33581
rect 49450 33562 49464 33581
rect 49520 33562 49540 33581
rect 49540 33562 49554 33581
rect 49610 33562 49630 33581
rect 49630 33562 49644 33581
rect 49700 33562 49734 33596
rect 49870 33562 49904 33596
rect 49960 33581 49994 33596
rect 50050 33581 50084 33596
rect 50140 33581 50174 33596
rect 50230 33581 50264 33596
rect 50320 33581 50354 33596
rect 50410 33581 50444 33596
rect 50500 33581 50534 33596
rect 50590 33581 50624 33596
rect 50680 33581 50714 33596
rect 50770 33581 50804 33596
rect 50860 33581 50894 33596
rect 50950 33581 50984 33596
rect 49960 33562 49980 33581
rect 49980 33562 49994 33581
rect 50050 33562 50070 33581
rect 50070 33562 50084 33581
rect 50140 33562 50160 33581
rect 50160 33562 50174 33581
rect 50230 33562 50250 33581
rect 50250 33562 50264 33581
rect 50320 33562 50340 33581
rect 50340 33562 50354 33581
rect 50410 33562 50430 33581
rect 50430 33562 50444 33581
rect 50500 33562 50520 33581
rect 50520 33562 50534 33581
rect 50590 33562 50610 33581
rect 50610 33562 50624 33581
rect 50680 33562 50700 33581
rect 50700 33562 50714 33581
rect 50770 33562 50790 33581
rect 50790 33562 50804 33581
rect 50860 33562 50880 33581
rect 50880 33562 50894 33581
rect 50950 33562 50970 33581
rect 50970 33562 50984 33581
rect 51040 33562 51074 33596
rect 51210 33562 51244 33596
rect 51300 33581 51334 33596
rect 51390 33581 51424 33596
rect 51480 33581 51514 33596
rect 51570 33581 51604 33596
rect 51660 33581 51694 33596
rect 51750 33581 51784 33596
rect 51840 33581 51874 33596
rect 51930 33581 51964 33596
rect 52020 33581 52054 33596
rect 52110 33581 52144 33596
rect 52200 33581 52234 33596
rect 52290 33581 52324 33596
rect 51300 33562 51320 33581
rect 51320 33562 51334 33581
rect 51390 33562 51410 33581
rect 51410 33562 51424 33581
rect 51480 33562 51500 33581
rect 51500 33562 51514 33581
rect 51570 33562 51590 33581
rect 51590 33562 51604 33581
rect 51660 33562 51680 33581
rect 51680 33562 51694 33581
rect 51750 33562 51770 33581
rect 51770 33562 51784 33581
rect 51840 33562 51860 33581
rect 51860 33562 51874 33581
rect 51930 33562 51950 33581
rect 51950 33562 51964 33581
rect 52020 33562 52040 33581
rect 52040 33562 52054 33581
rect 52110 33562 52130 33581
rect 52130 33562 52144 33581
rect 52200 33562 52220 33581
rect 52220 33562 52234 33581
rect 52290 33562 52310 33581
rect 52310 33562 52324 33581
rect 52380 33562 52414 33596
rect 41994 33402 42028 33436
rect 42084 33434 42118 33436
rect 42174 33434 42208 33436
rect 42264 33434 42298 33436
rect 42354 33434 42388 33436
rect 42444 33434 42478 33436
rect 42534 33434 42568 33436
rect 42624 33434 42658 33436
rect 42714 33434 42748 33436
rect 42804 33434 42838 33436
rect 42084 33402 42104 33434
rect 42104 33402 42118 33434
rect 42174 33402 42194 33434
rect 42194 33402 42208 33434
rect 42264 33402 42284 33434
rect 42284 33402 42298 33434
rect 42354 33402 42374 33434
rect 42374 33402 42388 33434
rect 42444 33402 42464 33434
rect 42464 33402 42478 33434
rect 42534 33402 42554 33434
rect 42554 33402 42568 33434
rect 42624 33402 42644 33434
rect 42644 33402 42658 33434
rect 42714 33402 42734 33434
rect 42734 33402 42748 33434
rect 42804 33402 42824 33434
rect 42824 33402 42838 33434
rect 42894 33402 42928 33436
rect 42180 33226 42202 33232
rect 42202 33226 42214 33232
rect 42280 33226 42292 33232
rect 42292 33226 42314 33232
rect 42380 33226 42382 33232
rect 42382 33226 42414 33232
rect 42180 33198 42214 33226
rect 42280 33198 42314 33226
rect 42380 33198 42414 33226
rect 42480 33198 42514 33232
rect 42580 33198 42614 33232
rect 42680 33226 42708 33232
rect 42708 33226 42714 33232
rect 42680 33198 42714 33226
rect 42180 33098 42214 33132
rect 42280 33098 42314 33132
rect 42380 33098 42414 33132
rect 42480 33098 42514 33132
rect 42580 33098 42614 33132
rect 42680 33098 42714 33132
rect 42180 32998 42214 33032
rect 42280 32998 42314 33032
rect 42380 32998 42414 33032
rect 42480 32998 42514 33032
rect 42580 32998 42614 33032
rect 42680 32998 42714 33032
rect 42180 32900 42214 32932
rect 42280 32900 42314 32932
rect 42380 32900 42414 32932
rect 42180 32898 42202 32900
rect 42202 32898 42214 32900
rect 42280 32898 42292 32900
rect 42292 32898 42314 32900
rect 42380 32898 42382 32900
rect 42382 32898 42414 32900
rect 42480 32898 42514 32932
rect 42580 32898 42614 32932
rect 42680 32900 42714 32932
rect 42680 32898 42708 32900
rect 42708 32898 42714 32900
rect 42180 32810 42214 32832
rect 42280 32810 42314 32832
rect 42380 32810 42414 32832
rect 42180 32798 42202 32810
rect 42202 32798 42214 32810
rect 42280 32798 42292 32810
rect 42292 32798 42314 32810
rect 42380 32798 42382 32810
rect 42382 32798 42414 32810
rect 42480 32798 42514 32832
rect 42580 32798 42614 32832
rect 42680 32810 42714 32832
rect 42680 32798 42708 32810
rect 42708 32798 42714 32810
rect 42180 32720 42214 32732
rect 42280 32720 42314 32732
rect 42380 32720 42414 32732
rect 42180 32698 42202 32720
rect 42202 32698 42214 32720
rect 42280 32698 42292 32720
rect 42292 32698 42314 32720
rect 42380 32698 42382 32720
rect 42382 32698 42414 32720
rect 42480 32698 42514 32732
rect 42580 32698 42614 32732
rect 42680 32720 42714 32732
rect 42680 32698 42708 32720
rect 42708 32698 42714 32720
rect 43334 33402 43368 33436
rect 43424 33434 43458 33436
rect 43514 33434 43548 33436
rect 43604 33434 43638 33436
rect 43694 33434 43728 33436
rect 43784 33434 43818 33436
rect 43874 33434 43908 33436
rect 43964 33434 43998 33436
rect 44054 33434 44088 33436
rect 44144 33434 44178 33436
rect 43424 33402 43444 33434
rect 43444 33402 43458 33434
rect 43514 33402 43534 33434
rect 43534 33402 43548 33434
rect 43604 33402 43624 33434
rect 43624 33402 43638 33434
rect 43694 33402 43714 33434
rect 43714 33402 43728 33434
rect 43784 33402 43804 33434
rect 43804 33402 43818 33434
rect 43874 33402 43894 33434
rect 43894 33402 43908 33434
rect 43964 33402 43984 33434
rect 43984 33402 43998 33434
rect 44054 33402 44074 33434
rect 44074 33402 44088 33434
rect 44144 33402 44164 33434
rect 44164 33402 44178 33434
rect 44234 33402 44268 33436
rect 43520 33226 43542 33232
rect 43542 33226 43554 33232
rect 43620 33226 43632 33232
rect 43632 33226 43654 33232
rect 43720 33226 43722 33232
rect 43722 33226 43754 33232
rect 43520 33198 43554 33226
rect 43620 33198 43654 33226
rect 43720 33198 43754 33226
rect 43820 33198 43854 33232
rect 43920 33198 43954 33232
rect 44020 33226 44048 33232
rect 44048 33226 44054 33232
rect 44020 33198 44054 33226
rect 43520 33098 43554 33132
rect 43620 33098 43654 33132
rect 43720 33098 43754 33132
rect 43820 33098 43854 33132
rect 43920 33098 43954 33132
rect 44020 33098 44054 33132
rect 43520 32998 43554 33032
rect 43620 32998 43654 33032
rect 43720 32998 43754 33032
rect 43820 32998 43854 33032
rect 43920 32998 43954 33032
rect 44020 32998 44054 33032
rect 43520 32900 43554 32932
rect 43620 32900 43654 32932
rect 43720 32900 43754 32932
rect 43520 32898 43542 32900
rect 43542 32898 43554 32900
rect 43620 32898 43632 32900
rect 43632 32898 43654 32900
rect 43720 32898 43722 32900
rect 43722 32898 43754 32900
rect 43820 32898 43854 32932
rect 43920 32898 43954 32932
rect 44020 32900 44054 32932
rect 44020 32898 44048 32900
rect 44048 32898 44054 32900
rect 43520 32810 43554 32832
rect 43620 32810 43654 32832
rect 43720 32810 43754 32832
rect 43520 32798 43542 32810
rect 43542 32798 43554 32810
rect 43620 32798 43632 32810
rect 43632 32798 43654 32810
rect 43720 32798 43722 32810
rect 43722 32798 43754 32810
rect 43820 32798 43854 32832
rect 43920 32798 43954 32832
rect 44020 32810 44054 32832
rect 44020 32798 44048 32810
rect 44048 32798 44054 32810
rect 43520 32720 43554 32732
rect 43620 32720 43654 32732
rect 43720 32720 43754 32732
rect 43520 32698 43542 32720
rect 43542 32698 43554 32720
rect 43620 32698 43632 32720
rect 43632 32698 43654 32720
rect 43720 32698 43722 32720
rect 43722 32698 43754 32720
rect 43820 32698 43854 32732
rect 43920 32698 43954 32732
rect 44020 32720 44054 32732
rect 44020 32698 44048 32720
rect 44048 32698 44054 32720
rect 44674 33402 44708 33436
rect 44764 33434 44798 33436
rect 44854 33434 44888 33436
rect 44944 33434 44978 33436
rect 45034 33434 45068 33436
rect 45124 33434 45158 33436
rect 45214 33434 45248 33436
rect 45304 33434 45338 33436
rect 45394 33434 45428 33436
rect 45484 33434 45518 33436
rect 44764 33402 44784 33434
rect 44784 33402 44798 33434
rect 44854 33402 44874 33434
rect 44874 33402 44888 33434
rect 44944 33402 44964 33434
rect 44964 33402 44978 33434
rect 45034 33402 45054 33434
rect 45054 33402 45068 33434
rect 45124 33402 45144 33434
rect 45144 33402 45158 33434
rect 45214 33402 45234 33434
rect 45234 33402 45248 33434
rect 45304 33402 45324 33434
rect 45324 33402 45338 33434
rect 45394 33402 45414 33434
rect 45414 33402 45428 33434
rect 45484 33402 45504 33434
rect 45504 33402 45518 33434
rect 45574 33402 45608 33436
rect 44860 33226 44882 33232
rect 44882 33226 44894 33232
rect 44960 33226 44972 33232
rect 44972 33226 44994 33232
rect 45060 33226 45062 33232
rect 45062 33226 45094 33232
rect 44860 33198 44894 33226
rect 44960 33198 44994 33226
rect 45060 33198 45094 33226
rect 45160 33198 45194 33232
rect 45260 33198 45294 33232
rect 45360 33226 45388 33232
rect 45388 33226 45394 33232
rect 45360 33198 45394 33226
rect 44860 33098 44894 33132
rect 44960 33098 44994 33132
rect 45060 33098 45094 33132
rect 45160 33098 45194 33132
rect 45260 33098 45294 33132
rect 45360 33098 45394 33132
rect 44860 32998 44894 33032
rect 44960 32998 44994 33032
rect 45060 32998 45094 33032
rect 45160 32998 45194 33032
rect 45260 32998 45294 33032
rect 45360 32998 45394 33032
rect 44860 32900 44894 32932
rect 44960 32900 44994 32932
rect 45060 32900 45094 32932
rect 44860 32898 44882 32900
rect 44882 32898 44894 32900
rect 44960 32898 44972 32900
rect 44972 32898 44994 32900
rect 45060 32898 45062 32900
rect 45062 32898 45094 32900
rect 45160 32898 45194 32932
rect 45260 32898 45294 32932
rect 45360 32900 45394 32932
rect 45360 32898 45388 32900
rect 45388 32898 45394 32900
rect 44860 32810 44894 32832
rect 44960 32810 44994 32832
rect 45060 32810 45094 32832
rect 44860 32798 44882 32810
rect 44882 32798 44894 32810
rect 44960 32798 44972 32810
rect 44972 32798 44994 32810
rect 45060 32798 45062 32810
rect 45062 32798 45094 32810
rect 45160 32798 45194 32832
rect 45260 32798 45294 32832
rect 45360 32810 45394 32832
rect 45360 32798 45388 32810
rect 45388 32798 45394 32810
rect 44860 32720 44894 32732
rect 44960 32720 44994 32732
rect 45060 32720 45094 32732
rect 44860 32698 44882 32720
rect 44882 32698 44894 32720
rect 44960 32698 44972 32720
rect 44972 32698 44994 32720
rect 45060 32698 45062 32720
rect 45062 32698 45094 32720
rect 45160 32698 45194 32732
rect 45260 32698 45294 32732
rect 45360 32720 45394 32732
rect 45360 32698 45388 32720
rect 45388 32698 45394 32720
rect 46014 33402 46048 33436
rect 46104 33434 46138 33436
rect 46194 33434 46228 33436
rect 46284 33434 46318 33436
rect 46374 33434 46408 33436
rect 46464 33434 46498 33436
rect 46554 33434 46588 33436
rect 46644 33434 46678 33436
rect 46734 33434 46768 33436
rect 46824 33434 46858 33436
rect 46104 33402 46124 33434
rect 46124 33402 46138 33434
rect 46194 33402 46214 33434
rect 46214 33402 46228 33434
rect 46284 33402 46304 33434
rect 46304 33402 46318 33434
rect 46374 33402 46394 33434
rect 46394 33402 46408 33434
rect 46464 33402 46484 33434
rect 46484 33402 46498 33434
rect 46554 33402 46574 33434
rect 46574 33402 46588 33434
rect 46644 33402 46664 33434
rect 46664 33402 46678 33434
rect 46734 33402 46754 33434
rect 46754 33402 46768 33434
rect 46824 33402 46844 33434
rect 46844 33402 46858 33434
rect 46914 33402 46948 33436
rect 46200 33226 46222 33232
rect 46222 33226 46234 33232
rect 46300 33226 46312 33232
rect 46312 33226 46334 33232
rect 46400 33226 46402 33232
rect 46402 33226 46434 33232
rect 46200 33198 46234 33226
rect 46300 33198 46334 33226
rect 46400 33198 46434 33226
rect 46500 33198 46534 33232
rect 46600 33198 46634 33232
rect 46700 33226 46728 33232
rect 46728 33226 46734 33232
rect 46700 33198 46734 33226
rect 46200 33098 46234 33132
rect 46300 33098 46334 33132
rect 46400 33098 46434 33132
rect 46500 33098 46534 33132
rect 46600 33098 46634 33132
rect 46700 33098 46734 33132
rect 46200 32998 46234 33032
rect 46300 32998 46334 33032
rect 46400 32998 46434 33032
rect 46500 32998 46534 33032
rect 46600 32998 46634 33032
rect 46700 32998 46734 33032
rect 46200 32900 46234 32932
rect 46300 32900 46334 32932
rect 46400 32900 46434 32932
rect 46200 32898 46222 32900
rect 46222 32898 46234 32900
rect 46300 32898 46312 32900
rect 46312 32898 46334 32900
rect 46400 32898 46402 32900
rect 46402 32898 46434 32900
rect 46500 32898 46534 32932
rect 46600 32898 46634 32932
rect 46700 32900 46734 32932
rect 46700 32898 46728 32900
rect 46728 32898 46734 32900
rect 46200 32810 46234 32832
rect 46300 32810 46334 32832
rect 46400 32810 46434 32832
rect 46200 32798 46222 32810
rect 46222 32798 46234 32810
rect 46300 32798 46312 32810
rect 46312 32798 46334 32810
rect 46400 32798 46402 32810
rect 46402 32798 46434 32810
rect 46500 32798 46534 32832
rect 46600 32798 46634 32832
rect 46700 32810 46734 32832
rect 46700 32798 46728 32810
rect 46728 32798 46734 32810
rect 46200 32720 46234 32732
rect 46300 32720 46334 32732
rect 46400 32720 46434 32732
rect 46200 32698 46222 32720
rect 46222 32698 46234 32720
rect 46300 32698 46312 32720
rect 46312 32698 46334 32720
rect 46400 32698 46402 32720
rect 46402 32698 46434 32720
rect 46500 32698 46534 32732
rect 46600 32698 46634 32732
rect 46700 32720 46734 32732
rect 46700 32698 46728 32720
rect 46728 32698 46734 32720
rect 47354 33402 47388 33436
rect 47444 33434 47478 33436
rect 47534 33434 47568 33436
rect 47624 33434 47658 33436
rect 47714 33434 47748 33436
rect 47804 33434 47838 33436
rect 47894 33434 47928 33436
rect 47984 33434 48018 33436
rect 48074 33434 48108 33436
rect 48164 33434 48198 33436
rect 47444 33402 47464 33434
rect 47464 33402 47478 33434
rect 47534 33402 47554 33434
rect 47554 33402 47568 33434
rect 47624 33402 47644 33434
rect 47644 33402 47658 33434
rect 47714 33402 47734 33434
rect 47734 33402 47748 33434
rect 47804 33402 47824 33434
rect 47824 33402 47838 33434
rect 47894 33402 47914 33434
rect 47914 33402 47928 33434
rect 47984 33402 48004 33434
rect 48004 33402 48018 33434
rect 48074 33402 48094 33434
rect 48094 33402 48108 33434
rect 48164 33402 48184 33434
rect 48184 33402 48198 33434
rect 48254 33402 48288 33436
rect 47540 33226 47562 33232
rect 47562 33226 47574 33232
rect 47640 33226 47652 33232
rect 47652 33226 47674 33232
rect 47740 33226 47742 33232
rect 47742 33226 47774 33232
rect 47540 33198 47574 33226
rect 47640 33198 47674 33226
rect 47740 33198 47774 33226
rect 47840 33198 47874 33232
rect 47940 33198 47974 33232
rect 48040 33226 48068 33232
rect 48068 33226 48074 33232
rect 48040 33198 48074 33226
rect 47540 33098 47574 33132
rect 47640 33098 47674 33132
rect 47740 33098 47774 33132
rect 47840 33098 47874 33132
rect 47940 33098 47974 33132
rect 48040 33098 48074 33132
rect 47540 32998 47574 33032
rect 47640 32998 47674 33032
rect 47740 32998 47774 33032
rect 47840 32998 47874 33032
rect 47940 32998 47974 33032
rect 48040 32998 48074 33032
rect 47540 32900 47574 32932
rect 47640 32900 47674 32932
rect 47740 32900 47774 32932
rect 47540 32898 47562 32900
rect 47562 32898 47574 32900
rect 47640 32898 47652 32900
rect 47652 32898 47674 32900
rect 47740 32898 47742 32900
rect 47742 32898 47774 32900
rect 47840 32898 47874 32932
rect 47940 32898 47974 32932
rect 48040 32900 48074 32932
rect 48040 32898 48068 32900
rect 48068 32898 48074 32900
rect 47540 32810 47574 32832
rect 47640 32810 47674 32832
rect 47740 32810 47774 32832
rect 47540 32798 47562 32810
rect 47562 32798 47574 32810
rect 47640 32798 47652 32810
rect 47652 32798 47674 32810
rect 47740 32798 47742 32810
rect 47742 32798 47774 32810
rect 47840 32798 47874 32832
rect 47940 32798 47974 32832
rect 48040 32810 48074 32832
rect 48040 32798 48068 32810
rect 48068 32798 48074 32810
rect 47540 32720 47574 32732
rect 47640 32720 47674 32732
rect 47740 32720 47774 32732
rect 47540 32698 47562 32720
rect 47562 32698 47574 32720
rect 47640 32698 47652 32720
rect 47652 32698 47674 32720
rect 47740 32698 47742 32720
rect 47742 32698 47774 32720
rect 47840 32698 47874 32732
rect 47940 32698 47974 32732
rect 48040 32720 48074 32732
rect 48040 32698 48068 32720
rect 48068 32698 48074 32720
rect 48694 33402 48728 33436
rect 48784 33434 48818 33436
rect 48874 33434 48908 33436
rect 48964 33434 48998 33436
rect 49054 33434 49088 33436
rect 49144 33434 49178 33436
rect 49234 33434 49268 33436
rect 49324 33434 49358 33436
rect 49414 33434 49448 33436
rect 49504 33434 49538 33436
rect 48784 33402 48804 33434
rect 48804 33402 48818 33434
rect 48874 33402 48894 33434
rect 48894 33402 48908 33434
rect 48964 33402 48984 33434
rect 48984 33402 48998 33434
rect 49054 33402 49074 33434
rect 49074 33402 49088 33434
rect 49144 33402 49164 33434
rect 49164 33402 49178 33434
rect 49234 33402 49254 33434
rect 49254 33402 49268 33434
rect 49324 33402 49344 33434
rect 49344 33402 49358 33434
rect 49414 33402 49434 33434
rect 49434 33402 49448 33434
rect 49504 33402 49524 33434
rect 49524 33402 49538 33434
rect 49594 33402 49628 33436
rect 48880 33226 48902 33232
rect 48902 33226 48914 33232
rect 48980 33226 48992 33232
rect 48992 33226 49014 33232
rect 49080 33226 49082 33232
rect 49082 33226 49114 33232
rect 48880 33198 48914 33226
rect 48980 33198 49014 33226
rect 49080 33198 49114 33226
rect 49180 33198 49214 33232
rect 49280 33198 49314 33232
rect 49380 33226 49408 33232
rect 49408 33226 49414 33232
rect 49380 33198 49414 33226
rect 48880 33098 48914 33132
rect 48980 33098 49014 33132
rect 49080 33098 49114 33132
rect 49180 33098 49214 33132
rect 49280 33098 49314 33132
rect 49380 33098 49414 33132
rect 48880 32998 48914 33032
rect 48980 32998 49014 33032
rect 49080 32998 49114 33032
rect 49180 32998 49214 33032
rect 49280 32998 49314 33032
rect 49380 32998 49414 33032
rect 48880 32900 48914 32932
rect 48980 32900 49014 32932
rect 49080 32900 49114 32932
rect 48880 32898 48902 32900
rect 48902 32898 48914 32900
rect 48980 32898 48992 32900
rect 48992 32898 49014 32900
rect 49080 32898 49082 32900
rect 49082 32898 49114 32900
rect 49180 32898 49214 32932
rect 49280 32898 49314 32932
rect 49380 32900 49414 32932
rect 49380 32898 49408 32900
rect 49408 32898 49414 32900
rect 48880 32810 48914 32832
rect 48980 32810 49014 32832
rect 49080 32810 49114 32832
rect 48880 32798 48902 32810
rect 48902 32798 48914 32810
rect 48980 32798 48992 32810
rect 48992 32798 49014 32810
rect 49080 32798 49082 32810
rect 49082 32798 49114 32810
rect 49180 32798 49214 32832
rect 49280 32798 49314 32832
rect 49380 32810 49414 32832
rect 49380 32798 49408 32810
rect 49408 32798 49414 32810
rect 48880 32720 48914 32732
rect 48980 32720 49014 32732
rect 49080 32720 49114 32732
rect 48880 32698 48902 32720
rect 48902 32698 48914 32720
rect 48980 32698 48992 32720
rect 48992 32698 49014 32720
rect 49080 32698 49082 32720
rect 49082 32698 49114 32720
rect 49180 32698 49214 32732
rect 49280 32698 49314 32732
rect 49380 32720 49414 32732
rect 49380 32698 49408 32720
rect 49408 32698 49414 32720
rect 50034 33402 50068 33436
rect 50124 33434 50158 33436
rect 50214 33434 50248 33436
rect 50304 33434 50338 33436
rect 50394 33434 50428 33436
rect 50484 33434 50518 33436
rect 50574 33434 50608 33436
rect 50664 33434 50698 33436
rect 50754 33434 50788 33436
rect 50844 33434 50878 33436
rect 50124 33402 50144 33434
rect 50144 33402 50158 33434
rect 50214 33402 50234 33434
rect 50234 33402 50248 33434
rect 50304 33402 50324 33434
rect 50324 33402 50338 33434
rect 50394 33402 50414 33434
rect 50414 33402 50428 33434
rect 50484 33402 50504 33434
rect 50504 33402 50518 33434
rect 50574 33402 50594 33434
rect 50594 33402 50608 33434
rect 50664 33402 50684 33434
rect 50684 33402 50698 33434
rect 50754 33402 50774 33434
rect 50774 33402 50788 33434
rect 50844 33402 50864 33434
rect 50864 33402 50878 33434
rect 50934 33402 50968 33436
rect 50220 33226 50242 33232
rect 50242 33226 50254 33232
rect 50320 33226 50332 33232
rect 50332 33226 50354 33232
rect 50420 33226 50422 33232
rect 50422 33226 50454 33232
rect 50220 33198 50254 33226
rect 50320 33198 50354 33226
rect 50420 33198 50454 33226
rect 50520 33198 50554 33232
rect 50620 33198 50654 33232
rect 50720 33226 50748 33232
rect 50748 33226 50754 33232
rect 50720 33198 50754 33226
rect 50220 33098 50254 33132
rect 50320 33098 50354 33132
rect 50420 33098 50454 33132
rect 50520 33098 50554 33132
rect 50620 33098 50654 33132
rect 50720 33098 50754 33132
rect 50220 32998 50254 33032
rect 50320 32998 50354 33032
rect 50420 32998 50454 33032
rect 50520 32998 50554 33032
rect 50620 32998 50654 33032
rect 50720 32998 50754 33032
rect 50220 32900 50254 32932
rect 50320 32900 50354 32932
rect 50420 32900 50454 32932
rect 50220 32898 50242 32900
rect 50242 32898 50254 32900
rect 50320 32898 50332 32900
rect 50332 32898 50354 32900
rect 50420 32898 50422 32900
rect 50422 32898 50454 32900
rect 50520 32898 50554 32932
rect 50620 32898 50654 32932
rect 50720 32900 50754 32932
rect 50720 32898 50748 32900
rect 50748 32898 50754 32900
rect 50220 32810 50254 32832
rect 50320 32810 50354 32832
rect 50420 32810 50454 32832
rect 50220 32798 50242 32810
rect 50242 32798 50254 32810
rect 50320 32798 50332 32810
rect 50332 32798 50354 32810
rect 50420 32798 50422 32810
rect 50422 32798 50454 32810
rect 50520 32798 50554 32832
rect 50620 32798 50654 32832
rect 50720 32810 50754 32832
rect 50720 32798 50748 32810
rect 50748 32798 50754 32810
rect 50220 32720 50254 32732
rect 50320 32720 50354 32732
rect 50420 32720 50454 32732
rect 50220 32698 50242 32720
rect 50242 32698 50254 32720
rect 50320 32698 50332 32720
rect 50332 32698 50354 32720
rect 50420 32698 50422 32720
rect 50422 32698 50454 32720
rect 50520 32698 50554 32732
rect 50620 32698 50654 32732
rect 50720 32720 50754 32732
rect 50720 32698 50748 32720
rect 50748 32698 50754 32720
rect 51374 33402 51408 33436
rect 51464 33434 51498 33436
rect 51554 33434 51588 33436
rect 51644 33434 51678 33436
rect 51734 33434 51768 33436
rect 51824 33434 51858 33436
rect 51914 33434 51948 33436
rect 52004 33434 52038 33436
rect 52094 33434 52128 33436
rect 52184 33434 52218 33436
rect 51464 33402 51484 33434
rect 51484 33402 51498 33434
rect 51554 33402 51574 33434
rect 51574 33402 51588 33434
rect 51644 33402 51664 33434
rect 51664 33402 51678 33434
rect 51734 33402 51754 33434
rect 51754 33402 51768 33434
rect 51824 33402 51844 33434
rect 51844 33402 51858 33434
rect 51914 33402 51934 33434
rect 51934 33402 51948 33434
rect 52004 33402 52024 33434
rect 52024 33402 52038 33434
rect 52094 33402 52114 33434
rect 52114 33402 52128 33434
rect 52184 33402 52204 33434
rect 52204 33402 52218 33434
rect 52274 33402 52308 33436
rect 51560 33226 51582 33232
rect 51582 33226 51594 33232
rect 51660 33226 51672 33232
rect 51672 33226 51694 33232
rect 51760 33226 51762 33232
rect 51762 33226 51794 33232
rect 51560 33198 51594 33226
rect 51660 33198 51694 33226
rect 51760 33198 51794 33226
rect 51860 33198 51894 33232
rect 51960 33198 51994 33232
rect 52060 33226 52088 33232
rect 52088 33226 52094 33232
rect 52060 33198 52094 33226
rect 51560 33098 51594 33132
rect 51660 33098 51694 33132
rect 51760 33098 51794 33132
rect 51860 33098 51894 33132
rect 51960 33098 51994 33132
rect 52060 33098 52094 33132
rect 51560 32998 51594 33032
rect 51660 32998 51694 33032
rect 51760 32998 51794 33032
rect 51860 32998 51894 33032
rect 51960 32998 51994 33032
rect 52060 32998 52094 33032
rect 51560 32900 51594 32932
rect 51660 32900 51694 32932
rect 51760 32900 51794 32932
rect 51560 32898 51582 32900
rect 51582 32898 51594 32900
rect 51660 32898 51672 32900
rect 51672 32898 51694 32900
rect 51760 32898 51762 32900
rect 51762 32898 51794 32900
rect 51860 32898 51894 32932
rect 51960 32898 51994 32932
rect 52060 32900 52094 32932
rect 52060 32898 52088 32900
rect 52088 32898 52094 32900
rect 51560 32810 51594 32832
rect 51660 32810 51694 32832
rect 51760 32810 51794 32832
rect 51560 32798 51582 32810
rect 51582 32798 51594 32810
rect 51660 32798 51672 32810
rect 51672 32798 51694 32810
rect 51760 32798 51762 32810
rect 51762 32798 51794 32810
rect 51860 32798 51894 32832
rect 51960 32798 51994 32832
rect 52060 32810 52094 32832
rect 52060 32798 52088 32810
rect 52088 32798 52094 32810
rect 51560 32720 51594 32732
rect 51660 32720 51694 32732
rect 51760 32720 51794 32732
rect 51560 32698 51582 32720
rect 51582 32698 51594 32720
rect 51660 32698 51672 32720
rect 51672 32698 51694 32720
rect 51760 32698 51762 32720
rect 51762 32698 51794 32720
rect 51860 32698 51894 32732
rect 51960 32698 51994 32732
rect 52060 32720 52094 32732
rect 52060 32698 52088 32720
rect 52088 32698 52094 32720
rect 19447 32015 19481 32049
rect 19647 32015 19681 32049
rect 19847 32015 19881 32049
rect 20047 32015 20081 32049
rect 20247 32015 20281 32049
rect 20447 32015 20481 32049
rect 20647 32015 20681 32049
rect 20847 32015 20881 32049
rect 21047 32015 21081 32049
rect 21247 32015 21281 32049
rect 21447 32015 21481 32049
rect 22193 32015 22227 32049
rect 22393 32015 22427 32049
rect 22593 32015 22627 32049
rect 22793 32015 22827 32049
rect 22993 32015 23027 32049
rect 23193 32015 23227 32049
rect 23393 32015 23427 32049
rect 23593 32015 23627 32049
rect 23793 32015 23827 32049
rect 23993 32015 24027 32049
rect 24193 32015 24227 32049
rect 24393 32015 24427 32049
rect 24593 32015 24627 32049
rect 24793 32015 24827 32049
rect 26387 32015 26421 32049
rect 26787 32015 26821 32049
rect 27187 32015 27221 32049
rect 27587 32015 27621 32049
rect 27987 32015 28021 32049
rect 28387 32015 28421 32049
rect 28787 32015 28821 32049
rect 29187 32015 29221 32049
rect 29587 32015 29621 32049
rect 29987 32015 30021 32049
rect 30387 32015 30421 32049
rect 30787 32015 30821 32049
rect 31187 32015 31221 32049
rect 31587 32015 31621 32049
rect 31987 32015 32021 32049
rect 32387 32015 32421 32049
rect 32787 32015 32821 32049
rect 33187 32015 33221 32049
rect 33835 32015 33869 32049
rect 34235 32015 34269 32049
rect 34635 32015 34669 32049
rect 35035 32015 35069 32049
rect 35435 32015 35469 32049
rect 35835 32015 35869 32049
rect 36235 32015 36269 32049
rect 36635 32015 36669 32049
rect 37035 32015 37069 32049
rect 37435 32015 37469 32049
rect 37835 32015 37869 32049
rect 38235 32015 38269 32049
rect 38635 32015 38669 32049
rect 39035 32015 39069 32049
rect 39435 32015 39469 32049
rect 39835 32015 39869 32049
rect 40235 32015 40269 32049
rect 40635 32015 40669 32049
rect 41967 32015 42001 32049
rect 42167 32015 42201 32049
rect 42367 32015 42401 32049
rect 42567 32015 42601 32049
rect 42767 32015 42801 32049
rect 42967 32015 43001 32049
rect 43167 32015 43201 32049
rect 43367 32015 43401 32049
rect 43567 32015 43601 32049
rect 43767 32015 43801 32049
rect 43967 32015 44001 32049
rect 44167 32015 44201 32049
rect 44367 32015 44401 32049
rect 44567 32015 44601 32049
rect 44767 32015 44801 32049
rect 44967 32015 45001 32049
rect 45167 32015 45201 32049
rect 45367 32015 45401 32049
rect 45567 32015 45601 32049
rect 45767 32015 45801 32049
rect 45967 32015 46001 32049
rect 46167 32015 46201 32049
rect 46367 32015 46401 32049
rect 46567 32015 46601 32049
rect 46767 32015 46801 32049
rect 46967 32015 47001 32049
rect 47167 32015 47201 32049
rect 47367 32015 47401 32049
rect 47567 32015 47601 32049
rect 47767 32015 47801 32049
rect 47967 32015 48001 32049
rect 48167 32015 48201 32049
rect 48367 32015 48401 32049
rect 48567 32015 48601 32049
rect 48767 32015 48801 32049
rect 48967 32015 49001 32049
rect 49167 32015 49201 32049
rect 49367 32015 49401 32049
rect 49567 32015 49601 32049
rect 49767 32015 49801 32049
rect 49967 32015 50001 32049
rect 50167 32015 50201 32049
rect 50367 32015 50401 32049
rect 50567 32015 50601 32049
rect 50767 32015 50801 32049
rect 50967 32015 51001 32049
rect 51167 32015 51201 32049
rect 51367 32015 51401 32049
rect 51567 32015 51601 32049
rect 51767 32015 51801 32049
rect 51967 32015 52001 32049
rect 52167 32015 52201 32049
rect 52367 32015 52401 32049
rect 16703 30135 16737 30169
rect 16903 30135 16937 30169
rect 17103 30135 17137 30169
rect 17303 30135 17337 30169
rect 17503 30135 17537 30169
rect 17703 30135 17737 30169
rect 17903 30135 17937 30169
rect 18103 30135 18137 30169
rect 18303 30135 18337 30169
rect 18503 30135 18537 30169
rect 18703 30135 18737 30169
rect 19447 30135 19481 30169
rect 19647 30135 19681 30169
rect 19847 30135 19881 30169
rect 20047 30135 20081 30169
rect 20247 30135 20281 30169
rect 20447 30135 20481 30169
rect 20647 30135 20681 30169
rect 20847 30135 20881 30169
rect 21047 30135 21081 30169
rect 21247 30135 21281 30169
rect 21447 30135 21481 30169
rect 22191 30135 22225 30169
rect 22391 30135 22425 30169
rect 22591 30135 22625 30169
rect 22791 30135 22825 30169
rect 22991 30135 23025 30169
rect 23191 30135 23225 30169
rect 23391 30135 23425 30169
rect 23591 30135 23625 30169
rect 23791 30135 23825 30169
rect 23991 30135 24025 30169
rect 24191 30135 24225 30169
rect 27385 30135 27419 30169
rect 27585 30135 27619 30169
rect 27785 30135 27819 30169
rect 27985 30135 28019 30169
rect 28185 30135 28219 30169
rect 28385 30135 28419 30169
rect 28585 30135 28619 30169
rect 28785 30135 28819 30169
rect 28985 30135 29019 30169
rect 29185 30135 29219 30169
rect 29385 30135 29419 30169
rect 30111 30135 30145 30169
rect 30511 30135 30545 30169
rect 30911 30135 30945 30169
rect 31311 30135 31345 30169
rect 31711 30135 31745 30169
rect 32111 30135 32145 30169
rect 32511 30135 32545 30169
rect 32911 30135 32945 30169
rect 33311 30135 33345 30169
rect 33711 30135 33745 30169
rect 34111 30135 34145 30169
rect 34511 30135 34545 30169
rect 34911 30135 34945 30169
rect 35311 30135 35345 30169
rect 35711 30135 35745 30169
rect 36111 30135 36145 30169
rect 36511 30135 36545 30169
rect 36911 30135 36945 30169
rect 37655 30135 37689 30169
rect 38055 30135 38089 30169
rect 38455 30135 38489 30169
rect 38855 30135 38889 30169
rect 39255 30135 39289 30169
rect 39655 30135 39689 30169
rect 40055 30135 40089 30169
rect 41967 30135 42001 30169
rect 42167 30135 42201 30169
rect 42367 30135 42401 30169
rect 42567 30135 42601 30169
rect 42767 30135 42801 30169
rect 42967 30135 43001 30169
rect 43167 30135 43201 30169
rect 43367 30135 43401 30169
rect 43567 30135 43601 30169
rect 43767 30135 43801 30169
rect 43967 30135 44001 30169
rect 44167 30135 44201 30169
rect 44367 30135 44401 30169
rect 44567 30135 44601 30169
rect 44767 30135 44801 30169
rect 44967 30135 45001 30169
rect 45167 30135 45201 30169
rect 45367 30135 45401 30169
rect 45567 30135 45601 30169
rect 45767 30135 45801 30169
rect 45967 30135 46001 30169
rect 46167 30135 46201 30169
rect 46367 30135 46401 30169
rect 46567 30135 46601 30169
rect 46767 30135 46801 30169
rect 46967 30135 47001 30169
rect 47167 30135 47201 30169
rect 47367 30135 47401 30169
rect 47567 30135 47601 30169
rect 47767 30135 47801 30169
rect 47967 30135 48001 30169
rect 48167 30135 48201 30169
rect 48367 30135 48401 30169
rect 48567 30135 48601 30169
rect 48767 30135 48801 30169
rect 48967 30135 49001 30169
rect 49167 30135 49201 30169
rect 49367 30135 49401 30169
rect 49567 30135 49601 30169
rect 49767 30135 49801 30169
rect 49967 30135 50001 30169
rect 50167 30135 50201 30169
rect 50367 30135 50401 30169
rect 50567 30135 50601 30169
rect 50767 30135 50801 30169
rect 50967 30135 51001 30169
rect 51167 30135 51201 30169
rect 51367 30135 51401 30169
rect 51567 30135 51601 30169
rect 51767 30135 51801 30169
rect 51967 30135 52001 30169
rect 52167 30135 52201 30169
rect 52367 30135 52401 30169
rect 16539 29363 16933 29901
rect 18546 29363 18940 29901
rect 19283 29363 19677 29901
rect 21290 29363 21684 29901
rect 22027 29363 22421 29901
rect 24034 29363 24428 29901
rect 27221 29363 27615 29901
rect 40325 29965 40359 29999
rect 29228 29363 29622 29901
rect 16539 28403 16933 28941
rect 18546 28403 18940 28941
rect 19283 28403 19677 28941
rect 21290 28403 21684 28941
rect 22027 28403 22421 28941
rect 24034 28403 24428 28941
rect 27221 28403 27615 28941
rect 29228 28403 29622 28941
rect 37519 29867 37553 29901
rect 37519 29799 37553 29829
rect 37519 29795 37553 29799
rect 37519 29731 37553 29757
rect 37519 29723 37553 29731
rect 37519 29663 37553 29685
rect 37519 29651 37553 29663
rect 37519 29595 37553 29613
rect 37519 29579 37553 29595
rect 37519 29527 37553 29541
rect 37519 29507 37553 29527
rect 37519 29459 37553 29469
rect 37519 29435 37553 29459
rect 37519 29391 37553 29397
rect 37519 29363 37553 29391
rect 37519 29323 37553 29325
rect 37519 29291 37553 29323
rect 37519 29221 37553 29253
rect 37519 29219 37553 29221
rect 37519 29153 37553 29181
rect 37519 29147 37553 29153
rect 37519 29085 37553 29109
rect 37519 29075 37553 29085
rect 37519 29017 37553 29037
rect 37519 29003 37553 29017
rect 37519 28949 37553 28965
rect 37519 28931 37553 28949
rect 37519 28881 37553 28893
rect 37519 28859 37553 28881
rect 37519 28813 37553 28821
rect 37519 28787 37553 28813
rect 37519 28745 37553 28749
rect 37519 28715 37553 28745
rect 37519 28643 37553 28677
rect 37977 29867 38011 29901
rect 37977 29799 38011 29829
rect 37977 29795 38011 29799
rect 37977 29731 38011 29757
rect 37977 29723 38011 29731
rect 37977 29663 38011 29685
rect 37977 29651 38011 29663
rect 37977 29595 38011 29613
rect 37977 29579 38011 29595
rect 37977 29527 38011 29541
rect 37977 29507 38011 29527
rect 37977 29459 38011 29469
rect 37977 29435 38011 29459
rect 37977 29391 38011 29397
rect 37977 29363 38011 29391
rect 37977 29323 38011 29325
rect 37977 29291 38011 29323
rect 37977 29221 38011 29253
rect 37977 29219 38011 29221
rect 37977 29153 38011 29181
rect 37977 29147 38011 29153
rect 37977 29085 38011 29109
rect 37977 29075 38011 29085
rect 37977 29017 38011 29037
rect 37977 29003 38011 29017
rect 37977 28949 38011 28965
rect 37977 28931 38011 28949
rect 37977 28881 38011 28893
rect 37977 28859 38011 28881
rect 37977 28813 38011 28821
rect 37977 28787 38011 28813
rect 37977 28745 38011 28749
rect 37977 28715 38011 28745
rect 37977 28643 38011 28677
rect 38435 29867 38469 29901
rect 38435 29799 38469 29829
rect 38435 29795 38469 29799
rect 38435 29731 38469 29757
rect 38435 29723 38469 29731
rect 38435 29663 38469 29685
rect 38435 29651 38469 29663
rect 38435 29595 38469 29613
rect 38435 29579 38469 29595
rect 38435 29527 38469 29541
rect 38435 29507 38469 29527
rect 38435 29459 38469 29469
rect 38435 29435 38469 29459
rect 38435 29391 38469 29397
rect 38435 29363 38469 29391
rect 38435 29323 38469 29325
rect 38435 29291 38469 29323
rect 38435 29221 38469 29253
rect 38435 29219 38469 29221
rect 38435 29153 38469 29181
rect 38435 29147 38469 29153
rect 38435 29085 38469 29109
rect 38435 29075 38469 29085
rect 38435 29017 38469 29037
rect 38435 29003 38469 29017
rect 38435 28949 38469 28965
rect 38435 28931 38469 28949
rect 38435 28881 38469 28893
rect 38435 28859 38469 28881
rect 38435 28813 38469 28821
rect 38435 28787 38469 28813
rect 38435 28745 38469 28749
rect 38435 28715 38469 28745
rect 38435 28643 38469 28677
rect 38893 29867 38927 29901
rect 38893 29799 38927 29829
rect 38893 29795 38927 29799
rect 38893 29731 38927 29757
rect 38893 29723 38927 29731
rect 38893 29663 38927 29685
rect 38893 29651 38927 29663
rect 38893 29595 38927 29613
rect 38893 29579 38927 29595
rect 38893 29527 38927 29541
rect 38893 29507 38927 29527
rect 38893 29459 38927 29469
rect 38893 29435 38927 29459
rect 38893 29391 38927 29397
rect 38893 29363 38927 29391
rect 38893 29323 38927 29325
rect 38893 29291 38927 29323
rect 38893 29221 38927 29253
rect 38893 29219 38927 29221
rect 38893 29153 38927 29181
rect 38893 29147 38927 29153
rect 38893 29085 38927 29109
rect 38893 29075 38927 29085
rect 38893 29017 38927 29037
rect 38893 29003 38927 29017
rect 38893 28949 38927 28965
rect 38893 28931 38927 28949
rect 38893 28881 38927 28893
rect 38893 28859 38927 28881
rect 38893 28813 38927 28821
rect 38893 28787 38927 28813
rect 38893 28745 38927 28749
rect 38893 28715 38927 28745
rect 38893 28643 38927 28677
rect 39351 29867 39385 29901
rect 39351 29799 39385 29829
rect 39351 29795 39385 29799
rect 39351 29731 39385 29757
rect 39351 29723 39385 29731
rect 39351 29663 39385 29685
rect 39351 29651 39385 29663
rect 39351 29595 39385 29613
rect 39351 29579 39385 29595
rect 39351 29527 39385 29541
rect 39351 29507 39385 29527
rect 39351 29459 39385 29469
rect 39351 29435 39385 29459
rect 39351 29391 39385 29397
rect 39351 29363 39385 29391
rect 39351 29323 39385 29325
rect 39351 29291 39385 29323
rect 39351 29221 39385 29253
rect 39351 29219 39385 29221
rect 39351 29153 39385 29181
rect 39351 29147 39385 29153
rect 39351 29085 39385 29109
rect 39351 29075 39385 29085
rect 39351 29017 39385 29037
rect 39351 29003 39385 29017
rect 39351 28949 39385 28965
rect 39351 28931 39385 28949
rect 39351 28881 39385 28893
rect 39351 28859 39385 28881
rect 39351 28813 39385 28821
rect 39351 28787 39385 28813
rect 39351 28745 39385 28749
rect 39351 28715 39385 28745
rect 39351 28643 39385 28677
rect 38577 28509 38611 28543
rect 39809 29867 39843 29901
rect 39809 29799 39843 29829
rect 39809 29795 39843 29799
rect 39809 29731 39843 29757
rect 39809 29723 39843 29731
rect 39809 29663 39843 29685
rect 39809 29651 39843 29663
rect 39809 29595 39843 29613
rect 39809 29579 39843 29595
rect 39809 29527 39843 29541
rect 39809 29507 39843 29527
rect 39809 29459 39843 29469
rect 39809 29435 39843 29459
rect 39809 29391 39843 29397
rect 39809 29363 39843 29391
rect 39809 29323 39843 29325
rect 39809 29291 39843 29323
rect 39809 29221 39843 29253
rect 39809 29219 39843 29221
rect 39809 29153 39843 29181
rect 39809 29147 39843 29153
rect 39809 29085 39843 29109
rect 39809 29075 39843 29085
rect 39809 29017 39843 29037
rect 39809 29003 39843 29017
rect 39809 28949 39843 28965
rect 39809 28931 39843 28949
rect 39809 28881 39843 28893
rect 39809 28859 39843 28881
rect 39809 28813 39843 28821
rect 39809 28787 39843 28813
rect 39809 28745 39843 28749
rect 39809 28715 39843 28745
rect 39809 28643 39843 28677
rect 40267 29867 40301 29901
rect 40267 29799 40301 29829
rect 40267 29795 40301 29799
rect 40267 29731 40301 29757
rect 40267 29723 40301 29731
rect 40267 29663 40301 29685
rect 40267 29651 40301 29663
rect 40267 29595 40301 29613
rect 40267 29579 40301 29595
rect 40267 29527 40301 29541
rect 40267 29507 40301 29527
rect 40267 29459 40301 29469
rect 40267 29435 40301 29459
rect 40267 29391 40301 29397
rect 40267 29363 40301 29391
rect 40267 29323 40301 29325
rect 40267 29291 40301 29323
rect 40267 29221 40301 29253
rect 40267 29219 40301 29221
rect 40267 29153 40301 29181
rect 40267 29147 40301 29153
rect 40267 29085 40301 29109
rect 40267 29075 40301 29085
rect 40267 29017 40301 29037
rect 40267 29003 40301 29017
rect 40267 28949 40301 28965
rect 40267 28931 40301 28949
rect 40267 28881 40301 28893
rect 40267 28859 40301 28881
rect 40267 28813 40301 28821
rect 40267 28787 40301 28813
rect 40267 28745 40301 28749
rect 40267 28715 40301 28745
rect 40267 28643 40301 28677
rect 41830 29802 41864 29836
rect 41920 29821 41954 29836
rect 42010 29821 42044 29836
rect 42100 29821 42134 29836
rect 42190 29821 42224 29836
rect 42280 29821 42314 29836
rect 42370 29821 42404 29836
rect 42460 29821 42494 29836
rect 42550 29821 42584 29836
rect 42640 29821 42674 29836
rect 42730 29821 42764 29836
rect 42820 29821 42854 29836
rect 42910 29821 42944 29836
rect 41920 29802 41940 29821
rect 41940 29802 41954 29821
rect 42010 29802 42030 29821
rect 42030 29802 42044 29821
rect 42100 29802 42120 29821
rect 42120 29802 42134 29821
rect 42190 29802 42210 29821
rect 42210 29802 42224 29821
rect 42280 29802 42300 29821
rect 42300 29802 42314 29821
rect 42370 29802 42390 29821
rect 42390 29802 42404 29821
rect 42460 29802 42480 29821
rect 42480 29802 42494 29821
rect 42550 29802 42570 29821
rect 42570 29802 42584 29821
rect 42640 29802 42660 29821
rect 42660 29802 42674 29821
rect 42730 29802 42750 29821
rect 42750 29802 42764 29821
rect 42820 29802 42840 29821
rect 42840 29802 42854 29821
rect 42910 29802 42930 29821
rect 42930 29802 42944 29821
rect 43000 29802 43034 29836
rect 43170 29802 43204 29836
rect 43260 29821 43294 29836
rect 43350 29821 43384 29836
rect 43440 29821 43474 29836
rect 43530 29821 43564 29836
rect 43620 29821 43654 29836
rect 43710 29821 43744 29836
rect 43800 29821 43834 29836
rect 43890 29821 43924 29836
rect 43980 29821 44014 29836
rect 44070 29821 44104 29836
rect 44160 29821 44194 29836
rect 44250 29821 44284 29836
rect 43260 29802 43280 29821
rect 43280 29802 43294 29821
rect 43350 29802 43370 29821
rect 43370 29802 43384 29821
rect 43440 29802 43460 29821
rect 43460 29802 43474 29821
rect 43530 29802 43550 29821
rect 43550 29802 43564 29821
rect 43620 29802 43640 29821
rect 43640 29802 43654 29821
rect 43710 29802 43730 29821
rect 43730 29802 43744 29821
rect 43800 29802 43820 29821
rect 43820 29802 43834 29821
rect 43890 29802 43910 29821
rect 43910 29802 43924 29821
rect 43980 29802 44000 29821
rect 44000 29802 44014 29821
rect 44070 29802 44090 29821
rect 44090 29802 44104 29821
rect 44160 29802 44180 29821
rect 44180 29802 44194 29821
rect 44250 29802 44270 29821
rect 44270 29802 44284 29821
rect 44340 29802 44374 29836
rect 44510 29802 44544 29836
rect 44600 29821 44634 29836
rect 44690 29821 44724 29836
rect 44780 29821 44814 29836
rect 44870 29821 44904 29836
rect 44960 29821 44994 29836
rect 45050 29821 45084 29836
rect 45140 29821 45174 29836
rect 45230 29821 45264 29836
rect 45320 29821 45354 29836
rect 45410 29821 45444 29836
rect 45500 29821 45534 29836
rect 45590 29821 45624 29836
rect 44600 29802 44620 29821
rect 44620 29802 44634 29821
rect 44690 29802 44710 29821
rect 44710 29802 44724 29821
rect 44780 29802 44800 29821
rect 44800 29802 44814 29821
rect 44870 29802 44890 29821
rect 44890 29802 44904 29821
rect 44960 29802 44980 29821
rect 44980 29802 44994 29821
rect 45050 29802 45070 29821
rect 45070 29802 45084 29821
rect 45140 29802 45160 29821
rect 45160 29802 45174 29821
rect 45230 29802 45250 29821
rect 45250 29802 45264 29821
rect 45320 29802 45340 29821
rect 45340 29802 45354 29821
rect 45410 29802 45430 29821
rect 45430 29802 45444 29821
rect 45500 29802 45520 29821
rect 45520 29802 45534 29821
rect 45590 29802 45610 29821
rect 45610 29802 45624 29821
rect 45680 29802 45714 29836
rect 45850 29802 45884 29836
rect 45940 29821 45974 29836
rect 46030 29821 46064 29836
rect 46120 29821 46154 29836
rect 46210 29821 46244 29836
rect 46300 29821 46334 29836
rect 46390 29821 46424 29836
rect 46480 29821 46514 29836
rect 46570 29821 46604 29836
rect 46660 29821 46694 29836
rect 46750 29821 46784 29836
rect 46840 29821 46874 29836
rect 46930 29821 46964 29836
rect 45940 29802 45960 29821
rect 45960 29802 45974 29821
rect 46030 29802 46050 29821
rect 46050 29802 46064 29821
rect 46120 29802 46140 29821
rect 46140 29802 46154 29821
rect 46210 29802 46230 29821
rect 46230 29802 46244 29821
rect 46300 29802 46320 29821
rect 46320 29802 46334 29821
rect 46390 29802 46410 29821
rect 46410 29802 46424 29821
rect 46480 29802 46500 29821
rect 46500 29802 46514 29821
rect 46570 29802 46590 29821
rect 46590 29802 46604 29821
rect 46660 29802 46680 29821
rect 46680 29802 46694 29821
rect 46750 29802 46770 29821
rect 46770 29802 46784 29821
rect 46840 29802 46860 29821
rect 46860 29802 46874 29821
rect 46930 29802 46950 29821
rect 46950 29802 46964 29821
rect 47020 29802 47054 29836
rect 47190 29802 47224 29836
rect 47280 29821 47314 29836
rect 47370 29821 47404 29836
rect 47460 29821 47494 29836
rect 47550 29821 47584 29836
rect 47640 29821 47674 29836
rect 47730 29821 47764 29836
rect 47820 29821 47854 29836
rect 47910 29821 47944 29836
rect 48000 29821 48034 29836
rect 48090 29821 48124 29836
rect 48180 29821 48214 29836
rect 48270 29821 48304 29836
rect 47280 29802 47300 29821
rect 47300 29802 47314 29821
rect 47370 29802 47390 29821
rect 47390 29802 47404 29821
rect 47460 29802 47480 29821
rect 47480 29802 47494 29821
rect 47550 29802 47570 29821
rect 47570 29802 47584 29821
rect 47640 29802 47660 29821
rect 47660 29802 47674 29821
rect 47730 29802 47750 29821
rect 47750 29802 47764 29821
rect 47820 29802 47840 29821
rect 47840 29802 47854 29821
rect 47910 29802 47930 29821
rect 47930 29802 47944 29821
rect 48000 29802 48020 29821
rect 48020 29802 48034 29821
rect 48090 29802 48110 29821
rect 48110 29802 48124 29821
rect 48180 29802 48200 29821
rect 48200 29802 48214 29821
rect 48270 29802 48290 29821
rect 48290 29802 48304 29821
rect 48360 29802 48394 29836
rect 48530 29802 48564 29836
rect 48620 29821 48654 29836
rect 48710 29821 48744 29836
rect 48800 29821 48834 29836
rect 48890 29821 48924 29836
rect 48980 29821 49014 29836
rect 49070 29821 49104 29836
rect 49160 29821 49194 29836
rect 49250 29821 49284 29836
rect 49340 29821 49374 29836
rect 49430 29821 49464 29836
rect 49520 29821 49554 29836
rect 49610 29821 49644 29836
rect 48620 29802 48640 29821
rect 48640 29802 48654 29821
rect 48710 29802 48730 29821
rect 48730 29802 48744 29821
rect 48800 29802 48820 29821
rect 48820 29802 48834 29821
rect 48890 29802 48910 29821
rect 48910 29802 48924 29821
rect 48980 29802 49000 29821
rect 49000 29802 49014 29821
rect 49070 29802 49090 29821
rect 49090 29802 49104 29821
rect 49160 29802 49180 29821
rect 49180 29802 49194 29821
rect 49250 29802 49270 29821
rect 49270 29802 49284 29821
rect 49340 29802 49360 29821
rect 49360 29802 49374 29821
rect 49430 29802 49450 29821
rect 49450 29802 49464 29821
rect 49520 29802 49540 29821
rect 49540 29802 49554 29821
rect 49610 29802 49630 29821
rect 49630 29802 49644 29821
rect 49700 29802 49734 29836
rect 49870 29802 49904 29836
rect 49960 29821 49994 29836
rect 50050 29821 50084 29836
rect 50140 29821 50174 29836
rect 50230 29821 50264 29836
rect 50320 29821 50354 29836
rect 50410 29821 50444 29836
rect 50500 29821 50534 29836
rect 50590 29821 50624 29836
rect 50680 29821 50714 29836
rect 50770 29821 50804 29836
rect 50860 29821 50894 29836
rect 50950 29821 50984 29836
rect 49960 29802 49980 29821
rect 49980 29802 49994 29821
rect 50050 29802 50070 29821
rect 50070 29802 50084 29821
rect 50140 29802 50160 29821
rect 50160 29802 50174 29821
rect 50230 29802 50250 29821
rect 50250 29802 50264 29821
rect 50320 29802 50340 29821
rect 50340 29802 50354 29821
rect 50410 29802 50430 29821
rect 50430 29802 50444 29821
rect 50500 29802 50520 29821
rect 50520 29802 50534 29821
rect 50590 29802 50610 29821
rect 50610 29802 50624 29821
rect 50680 29802 50700 29821
rect 50700 29802 50714 29821
rect 50770 29802 50790 29821
rect 50790 29802 50804 29821
rect 50860 29802 50880 29821
rect 50880 29802 50894 29821
rect 50950 29802 50970 29821
rect 50970 29802 50984 29821
rect 51040 29802 51074 29836
rect 51210 29802 51244 29836
rect 51300 29821 51334 29836
rect 51390 29821 51424 29836
rect 51480 29821 51514 29836
rect 51570 29821 51604 29836
rect 51660 29821 51694 29836
rect 51750 29821 51784 29836
rect 51840 29821 51874 29836
rect 51930 29821 51964 29836
rect 52020 29821 52054 29836
rect 52110 29821 52144 29836
rect 52200 29821 52234 29836
rect 52290 29821 52324 29836
rect 51300 29802 51320 29821
rect 51320 29802 51334 29821
rect 51390 29802 51410 29821
rect 51410 29802 51424 29821
rect 51480 29802 51500 29821
rect 51500 29802 51514 29821
rect 51570 29802 51590 29821
rect 51590 29802 51604 29821
rect 51660 29802 51680 29821
rect 51680 29802 51694 29821
rect 51750 29802 51770 29821
rect 51770 29802 51784 29821
rect 51840 29802 51860 29821
rect 51860 29802 51874 29821
rect 51930 29802 51950 29821
rect 51950 29802 51964 29821
rect 52020 29802 52040 29821
rect 52040 29802 52054 29821
rect 52110 29802 52130 29821
rect 52130 29802 52144 29821
rect 52200 29802 52220 29821
rect 52220 29802 52234 29821
rect 52290 29802 52310 29821
rect 52310 29802 52324 29821
rect 52380 29802 52414 29836
rect 41994 29642 42028 29676
rect 42084 29674 42118 29676
rect 42174 29674 42208 29676
rect 42264 29674 42298 29676
rect 42354 29674 42388 29676
rect 42444 29674 42478 29676
rect 42534 29674 42568 29676
rect 42624 29674 42658 29676
rect 42714 29674 42748 29676
rect 42804 29674 42838 29676
rect 42084 29642 42104 29674
rect 42104 29642 42118 29674
rect 42174 29642 42194 29674
rect 42194 29642 42208 29674
rect 42264 29642 42284 29674
rect 42284 29642 42298 29674
rect 42354 29642 42374 29674
rect 42374 29642 42388 29674
rect 42444 29642 42464 29674
rect 42464 29642 42478 29674
rect 42534 29642 42554 29674
rect 42554 29642 42568 29674
rect 42624 29642 42644 29674
rect 42644 29642 42658 29674
rect 42714 29642 42734 29674
rect 42734 29642 42748 29674
rect 42804 29642 42824 29674
rect 42824 29642 42838 29674
rect 42894 29642 42928 29676
rect 42180 29466 42202 29472
rect 42202 29466 42214 29472
rect 42280 29466 42292 29472
rect 42292 29466 42314 29472
rect 42380 29466 42382 29472
rect 42382 29466 42414 29472
rect 42180 29438 42214 29466
rect 42280 29438 42314 29466
rect 42380 29438 42414 29466
rect 42480 29438 42514 29472
rect 42580 29438 42614 29472
rect 42680 29466 42708 29472
rect 42708 29466 42714 29472
rect 42680 29438 42714 29466
rect 42180 29338 42214 29372
rect 42280 29338 42314 29372
rect 42380 29338 42414 29372
rect 42480 29338 42514 29372
rect 42580 29338 42614 29372
rect 42680 29338 42714 29372
rect 42180 29238 42214 29272
rect 42280 29238 42314 29272
rect 42380 29238 42414 29272
rect 42480 29238 42514 29272
rect 42580 29238 42614 29272
rect 42680 29238 42714 29272
rect 42180 29140 42214 29172
rect 42280 29140 42314 29172
rect 42380 29140 42414 29172
rect 42180 29138 42202 29140
rect 42202 29138 42214 29140
rect 42280 29138 42292 29140
rect 42292 29138 42314 29140
rect 42380 29138 42382 29140
rect 42382 29138 42414 29140
rect 42480 29138 42514 29172
rect 42580 29138 42614 29172
rect 42680 29140 42714 29172
rect 42680 29138 42708 29140
rect 42708 29138 42714 29140
rect 42180 29050 42214 29072
rect 42280 29050 42314 29072
rect 42380 29050 42414 29072
rect 42180 29038 42202 29050
rect 42202 29038 42214 29050
rect 42280 29038 42292 29050
rect 42292 29038 42314 29050
rect 42380 29038 42382 29050
rect 42382 29038 42414 29050
rect 42480 29038 42514 29072
rect 42580 29038 42614 29072
rect 42680 29050 42714 29072
rect 42680 29038 42708 29050
rect 42708 29038 42714 29050
rect 42180 28960 42214 28972
rect 42280 28960 42314 28972
rect 42380 28960 42414 28972
rect 42180 28938 42202 28960
rect 42202 28938 42214 28960
rect 42280 28938 42292 28960
rect 42292 28938 42314 28960
rect 42380 28938 42382 28960
rect 42382 28938 42414 28960
rect 42480 28938 42514 28972
rect 42580 28938 42614 28972
rect 42680 28960 42714 28972
rect 42680 28938 42708 28960
rect 42708 28938 42714 28960
rect 43334 29642 43368 29676
rect 43424 29674 43458 29676
rect 43514 29674 43548 29676
rect 43604 29674 43638 29676
rect 43694 29674 43728 29676
rect 43784 29674 43818 29676
rect 43874 29674 43908 29676
rect 43964 29674 43998 29676
rect 44054 29674 44088 29676
rect 44144 29674 44178 29676
rect 43424 29642 43444 29674
rect 43444 29642 43458 29674
rect 43514 29642 43534 29674
rect 43534 29642 43548 29674
rect 43604 29642 43624 29674
rect 43624 29642 43638 29674
rect 43694 29642 43714 29674
rect 43714 29642 43728 29674
rect 43784 29642 43804 29674
rect 43804 29642 43818 29674
rect 43874 29642 43894 29674
rect 43894 29642 43908 29674
rect 43964 29642 43984 29674
rect 43984 29642 43998 29674
rect 44054 29642 44074 29674
rect 44074 29642 44088 29674
rect 44144 29642 44164 29674
rect 44164 29642 44178 29674
rect 44234 29642 44268 29676
rect 43520 29466 43542 29472
rect 43542 29466 43554 29472
rect 43620 29466 43632 29472
rect 43632 29466 43654 29472
rect 43720 29466 43722 29472
rect 43722 29466 43754 29472
rect 43520 29438 43554 29466
rect 43620 29438 43654 29466
rect 43720 29438 43754 29466
rect 43820 29438 43854 29472
rect 43920 29438 43954 29472
rect 44020 29466 44048 29472
rect 44048 29466 44054 29472
rect 44020 29438 44054 29466
rect 43520 29338 43554 29372
rect 43620 29338 43654 29372
rect 43720 29338 43754 29372
rect 43820 29338 43854 29372
rect 43920 29338 43954 29372
rect 44020 29338 44054 29372
rect 43520 29238 43554 29272
rect 43620 29238 43654 29272
rect 43720 29238 43754 29272
rect 43820 29238 43854 29272
rect 43920 29238 43954 29272
rect 44020 29238 44054 29272
rect 43520 29140 43554 29172
rect 43620 29140 43654 29172
rect 43720 29140 43754 29172
rect 43520 29138 43542 29140
rect 43542 29138 43554 29140
rect 43620 29138 43632 29140
rect 43632 29138 43654 29140
rect 43720 29138 43722 29140
rect 43722 29138 43754 29140
rect 43820 29138 43854 29172
rect 43920 29138 43954 29172
rect 44020 29140 44054 29172
rect 44020 29138 44048 29140
rect 44048 29138 44054 29140
rect 43520 29050 43554 29072
rect 43620 29050 43654 29072
rect 43720 29050 43754 29072
rect 43520 29038 43542 29050
rect 43542 29038 43554 29050
rect 43620 29038 43632 29050
rect 43632 29038 43654 29050
rect 43720 29038 43722 29050
rect 43722 29038 43754 29050
rect 43820 29038 43854 29072
rect 43920 29038 43954 29072
rect 44020 29050 44054 29072
rect 44020 29038 44048 29050
rect 44048 29038 44054 29050
rect 43520 28960 43554 28972
rect 43620 28960 43654 28972
rect 43720 28960 43754 28972
rect 43520 28938 43542 28960
rect 43542 28938 43554 28960
rect 43620 28938 43632 28960
rect 43632 28938 43654 28960
rect 43720 28938 43722 28960
rect 43722 28938 43754 28960
rect 43820 28938 43854 28972
rect 43920 28938 43954 28972
rect 44020 28960 44054 28972
rect 44020 28938 44048 28960
rect 44048 28938 44054 28960
rect 44674 29642 44708 29676
rect 44764 29674 44798 29676
rect 44854 29674 44888 29676
rect 44944 29674 44978 29676
rect 45034 29674 45068 29676
rect 45124 29674 45158 29676
rect 45214 29674 45248 29676
rect 45304 29674 45338 29676
rect 45394 29674 45428 29676
rect 45484 29674 45518 29676
rect 44764 29642 44784 29674
rect 44784 29642 44798 29674
rect 44854 29642 44874 29674
rect 44874 29642 44888 29674
rect 44944 29642 44964 29674
rect 44964 29642 44978 29674
rect 45034 29642 45054 29674
rect 45054 29642 45068 29674
rect 45124 29642 45144 29674
rect 45144 29642 45158 29674
rect 45214 29642 45234 29674
rect 45234 29642 45248 29674
rect 45304 29642 45324 29674
rect 45324 29642 45338 29674
rect 45394 29642 45414 29674
rect 45414 29642 45428 29674
rect 45484 29642 45504 29674
rect 45504 29642 45518 29674
rect 45574 29642 45608 29676
rect 44860 29466 44882 29472
rect 44882 29466 44894 29472
rect 44960 29466 44972 29472
rect 44972 29466 44994 29472
rect 45060 29466 45062 29472
rect 45062 29466 45094 29472
rect 44860 29438 44894 29466
rect 44960 29438 44994 29466
rect 45060 29438 45094 29466
rect 45160 29438 45194 29472
rect 45260 29438 45294 29472
rect 45360 29466 45388 29472
rect 45388 29466 45394 29472
rect 45360 29438 45394 29466
rect 44860 29338 44894 29372
rect 44960 29338 44994 29372
rect 45060 29338 45094 29372
rect 45160 29338 45194 29372
rect 45260 29338 45294 29372
rect 45360 29338 45394 29372
rect 44860 29238 44894 29272
rect 44960 29238 44994 29272
rect 45060 29238 45094 29272
rect 45160 29238 45194 29272
rect 45260 29238 45294 29272
rect 45360 29238 45394 29272
rect 44860 29140 44894 29172
rect 44960 29140 44994 29172
rect 45060 29140 45094 29172
rect 44860 29138 44882 29140
rect 44882 29138 44894 29140
rect 44960 29138 44972 29140
rect 44972 29138 44994 29140
rect 45060 29138 45062 29140
rect 45062 29138 45094 29140
rect 45160 29138 45194 29172
rect 45260 29138 45294 29172
rect 45360 29140 45394 29172
rect 45360 29138 45388 29140
rect 45388 29138 45394 29140
rect 44860 29050 44894 29072
rect 44960 29050 44994 29072
rect 45060 29050 45094 29072
rect 44860 29038 44882 29050
rect 44882 29038 44894 29050
rect 44960 29038 44972 29050
rect 44972 29038 44994 29050
rect 45060 29038 45062 29050
rect 45062 29038 45094 29050
rect 45160 29038 45194 29072
rect 45260 29038 45294 29072
rect 45360 29050 45394 29072
rect 45360 29038 45388 29050
rect 45388 29038 45394 29050
rect 44860 28960 44894 28972
rect 44960 28960 44994 28972
rect 45060 28960 45094 28972
rect 44860 28938 44882 28960
rect 44882 28938 44894 28960
rect 44960 28938 44972 28960
rect 44972 28938 44994 28960
rect 45060 28938 45062 28960
rect 45062 28938 45094 28960
rect 45160 28938 45194 28972
rect 45260 28938 45294 28972
rect 45360 28960 45394 28972
rect 45360 28938 45388 28960
rect 45388 28938 45394 28960
rect 46014 29642 46048 29676
rect 46104 29674 46138 29676
rect 46194 29674 46228 29676
rect 46284 29674 46318 29676
rect 46374 29674 46408 29676
rect 46464 29674 46498 29676
rect 46554 29674 46588 29676
rect 46644 29674 46678 29676
rect 46734 29674 46768 29676
rect 46824 29674 46858 29676
rect 46104 29642 46124 29674
rect 46124 29642 46138 29674
rect 46194 29642 46214 29674
rect 46214 29642 46228 29674
rect 46284 29642 46304 29674
rect 46304 29642 46318 29674
rect 46374 29642 46394 29674
rect 46394 29642 46408 29674
rect 46464 29642 46484 29674
rect 46484 29642 46498 29674
rect 46554 29642 46574 29674
rect 46574 29642 46588 29674
rect 46644 29642 46664 29674
rect 46664 29642 46678 29674
rect 46734 29642 46754 29674
rect 46754 29642 46768 29674
rect 46824 29642 46844 29674
rect 46844 29642 46858 29674
rect 46914 29642 46948 29676
rect 46200 29466 46222 29472
rect 46222 29466 46234 29472
rect 46300 29466 46312 29472
rect 46312 29466 46334 29472
rect 46400 29466 46402 29472
rect 46402 29466 46434 29472
rect 46200 29438 46234 29466
rect 46300 29438 46334 29466
rect 46400 29438 46434 29466
rect 46500 29438 46534 29472
rect 46600 29438 46634 29472
rect 46700 29466 46728 29472
rect 46728 29466 46734 29472
rect 46700 29438 46734 29466
rect 46200 29338 46234 29372
rect 46300 29338 46334 29372
rect 46400 29338 46434 29372
rect 46500 29338 46534 29372
rect 46600 29338 46634 29372
rect 46700 29338 46734 29372
rect 46200 29238 46234 29272
rect 46300 29238 46334 29272
rect 46400 29238 46434 29272
rect 46500 29238 46534 29272
rect 46600 29238 46634 29272
rect 46700 29238 46734 29272
rect 46200 29140 46234 29172
rect 46300 29140 46334 29172
rect 46400 29140 46434 29172
rect 46200 29138 46222 29140
rect 46222 29138 46234 29140
rect 46300 29138 46312 29140
rect 46312 29138 46334 29140
rect 46400 29138 46402 29140
rect 46402 29138 46434 29140
rect 46500 29138 46534 29172
rect 46600 29138 46634 29172
rect 46700 29140 46734 29172
rect 46700 29138 46728 29140
rect 46728 29138 46734 29140
rect 46200 29050 46234 29072
rect 46300 29050 46334 29072
rect 46400 29050 46434 29072
rect 46200 29038 46222 29050
rect 46222 29038 46234 29050
rect 46300 29038 46312 29050
rect 46312 29038 46334 29050
rect 46400 29038 46402 29050
rect 46402 29038 46434 29050
rect 46500 29038 46534 29072
rect 46600 29038 46634 29072
rect 46700 29050 46734 29072
rect 46700 29038 46728 29050
rect 46728 29038 46734 29050
rect 46200 28960 46234 28972
rect 46300 28960 46334 28972
rect 46400 28960 46434 28972
rect 46200 28938 46222 28960
rect 46222 28938 46234 28960
rect 46300 28938 46312 28960
rect 46312 28938 46334 28960
rect 46400 28938 46402 28960
rect 46402 28938 46434 28960
rect 46500 28938 46534 28972
rect 46600 28938 46634 28972
rect 46700 28960 46734 28972
rect 46700 28938 46728 28960
rect 46728 28938 46734 28960
rect 47354 29642 47388 29676
rect 47444 29674 47478 29676
rect 47534 29674 47568 29676
rect 47624 29674 47658 29676
rect 47714 29674 47748 29676
rect 47804 29674 47838 29676
rect 47894 29674 47928 29676
rect 47984 29674 48018 29676
rect 48074 29674 48108 29676
rect 48164 29674 48198 29676
rect 47444 29642 47464 29674
rect 47464 29642 47478 29674
rect 47534 29642 47554 29674
rect 47554 29642 47568 29674
rect 47624 29642 47644 29674
rect 47644 29642 47658 29674
rect 47714 29642 47734 29674
rect 47734 29642 47748 29674
rect 47804 29642 47824 29674
rect 47824 29642 47838 29674
rect 47894 29642 47914 29674
rect 47914 29642 47928 29674
rect 47984 29642 48004 29674
rect 48004 29642 48018 29674
rect 48074 29642 48094 29674
rect 48094 29642 48108 29674
rect 48164 29642 48184 29674
rect 48184 29642 48198 29674
rect 48254 29642 48288 29676
rect 47540 29466 47562 29472
rect 47562 29466 47574 29472
rect 47640 29466 47652 29472
rect 47652 29466 47674 29472
rect 47740 29466 47742 29472
rect 47742 29466 47774 29472
rect 47540 29438 47574 29466
rect 47640 29438 47674 29466
rect 47740 29438 47774 29466
rect 47840 29438 47874 29472
rect 47940 29438 47974 29472
rect 48040 29466 48068 29472
rect 48068 29466 48074 29472
rect 48040 29438 48074 29466
rect 47540 29338 47574 29372
rect 47640 29338 47674 29372
rect 47740 29338 47774 29372
rect 47840 29338 47874 29372
rect 47940 29338 47974 29372
rect 48040 29338 48074 29372
rect 47540 29238 47574 29272
rect 47640 29238 47674 29272
rect 47740 29238 47774 29272
rect 47840 29238 47874 29272
rect 47940 29238 47974 29272
rect 48040 29238 48074 29272
rect 47540 29140 47574 29172
rect 47640 29140 47674 29172
rect 47740 29140 47774 29172
rect 47540 29138 47562 29140
rect 47562 29138 47574 29140
rect 47640 29138 47652 29140
rect 47652 29138 47674 29140
rect 47740 29138 47742 29140
rect 47742 29138 47774 29140
rect 47840 29138 47874 29172
rect 47940 29138 47974 29172
rect 48040 29140 48074 29172
rect 48040 29138 48068 29140
rect 48068 29138 48074 29140
rect 47540 29050 47574 29072
rect 47640 29050 47674 29072
rect 47740 29050 47774 29072
rect 47540 29038 47562 29050
rect 47562 29038 47574 29050
rect 47640 29038 47652 29050
rect 47652 29038 47674 29050
rect 47740 29038 47742 29050
rect 47742 29038 47774 29050
rect 47840 29038 47874 29072
rect 47940 29038 47974 29072
rect 48040 29050 48074 29072
rect 48040 29038 48068 29050
rect 48068 29038 48074 29050
rect 47540 28960 47574 28972
rect 47640 28960 47674 28972
rect 47740 28960 47774 28972
rect 47540 28938 47562 28960
rect 47562 28938 47574 28960
rect 47640 28938 47652 28960
rect 47652 28938 47674 28960
rect 47740 28938 47742 28960
rect 47742 28938 47774 28960
rect 47840 28938 47874 28972
rect 47940 28938 47974 28972
rect 48040 28960 48074 28972
rect 48040 28938 48068 28960
rect 48068 28938 48074 28960
rect 48694 29642 48728 29676
rect 48784 29674 48818 29676
rect 48874 29674 48908 29676
rect 48964 29674 48998 29676
rect 49054 29674 49088 29676
rect 49144 29674 49178 29676
rect 49234 29674 49268 29676
rect 49324 29674 49358 29676
rect 49414 29674 49448 29676
rect 49504 29674 49538 29676
rect 48784 29642 48804 29674
rect 48804 29642 48818 29674
rect 48874 29642 48894 29674
rect 48894 29642 48908 29674
rect 48964 29642 48984 29674
rect 48984 29642 48998 29674
rect 49054 29642 49074 29674
rect 49074 29642 49088 29674
rect 49144 29642 49164 29674
rect 49164 29642 49178 29674
rect 49234 29642 49254 29674
rect 49254 29642 49268 29674
rect 49324 29642 49344 29674
rect 49344 29642 49358 29674
rect 49414 29642 49434 29674
rect 49434 29642 49448 29674
rect 49504 29642 49524 29674
rect 49524 29642 49538 29674
rect 49594 29642 49628 29676
rect 48880 29466 48902 29472
rect 48902 29466 48914 29472
rect 48980 29466 48992 29472
rect 48992 29466 49014 29472
rect 49080 29466 49082 29472
rect 49082 29466 49114 29472
rect 48880 29438 48914 29466
rect 48980 29438 49014 29466
rect 49080 29438 49114 29466
rect 49180 29438 49214 29472
rect 49280 29438 49314 29472
rect 49380 29466 49408 29472
rect 49408 29466 49414 29472
rect 49380 29438 49414 29466
rect 48880 29338 48914 29372
rect 48980 29338 49014 29372
rect 49080 29338 49114 29372
rect 49180 29338 49214 29372
rect 49280 29338 49314 29372
rect 49380 29338 49414 29372
rect 48880 29238 48914 29272
rect 48980 29238 49014 29272
rect 49080 29238 49114 29272
rect 49180 29238 49214 29272
rect 49280 29238 49314 29272
rect 49380 29238 49414 29272
rect 48880 29140 48914 29172
rect 48980 29140 49014 29172
rect 49080 29140 49114 29172
rect 48880 29138 48902 29140
rect 48902 29138 48914 29140
rect 48980 29138 48992 29140
rect 48992 29138 49014 29140
rect 49080 29138 49082 29140
rect 49082 29138 49114 29140
rect 49180 29138 49214 29172
rect 49280 29138 49314 29172
rect 49380 29140 49414 29172
rect 49380 29138 49408 29140
rect 49408 29138 49414 29140
rect 48880 29050 48914 29072
rect 48980 29050 49014 29072
rect 49080 29050 49114 29072
rect 48880 29038 48902 29050
rect 48902 29038 48914 29050
rect 48980 29038 48992 29050
rect 48992 29038 49014 29050
rect 49080 29038 49082 29050
rect 49082 29038 49114 29050
rect 49180 29038 49214 29072
rect 49280 29038 49314 29072
rect 49380 29050 49414 29072
rect 49380 29038 49408 29050
rect 49408 29038 49414 29050
rect 48880 28960 48914 28972
rect 48980 28960 49014 28972
rect 49080 28960 49114 28972
rect 48880 28938 48902 28960
rect 48902 28938 48914 28960
rect 48980 28938 48992 28960
rect 48992 28938 49014 28960
rect 49080 28938 49082 28960
rect 49082 28938 49114 28960
rect 49180 28938 49214 28972
rect 49280 28938 49314 28972
rect 49380 28960 49414 28972
rect 49380 28938 49408 28960
rect 49408 28938 49414 28960
rect 50034 29642 50068 29676
rect 50124 29674 50158 29676
rect 50214 29674 50248 29676
rect 50304 29674 50338 29676
rect 50394 29674 50428 29676
rect 50484 29674 50518 29676
rect 50574 29674 50608 29676
rect 50664 29674 50698 29676
rect 50754 29674 50788 29676
rect 50844 29674 50878 29676
rect 50124 29642 50144 29674
rect 50144 29642 50158 29674
rect 50214 29642 50234 29674
rect 50234 29642 50248 29674
rect 50304 29642 50324 29674
rect 50324 29642 50338 29674
rect 50394 29642 50414 29674
rect 50414 29642 50428 29674
rect 50484 29642 50504 29674
rect 50504 29642 50518 29674
rect 50574 29642 50594 29674
rect 50594 29642 50608 29674
rect 50664 29642 50684 29674
rect 50684 29642 50698 29674
rect 50754 29642 50774 29674
rect 50774 29642 50788 29674
rect 50844 29642 50864 29674
rect 50864 29642 50878 29674
rect 50934 29642 50968 29676
rect 50220 29466 50242 29472
rect 50242 29466 50254 29472
rect 50320 29466 50332 29472
rect 50332 29466 50354 29472
rect 50420 29466 50422 29472
rect 50422 29466 50454 29472
rect 50220 29438 50254 29466
rect 50320 29438 50354 29466
rect 50420 29438 50454 29466
rect 50520 29438 50554 29472
rect 50620 29438 50654 29472
rect 50720 29466 50748 29472
rect 50748 29466 50754 29472
rect 50720 29438 50754 29466
rect 50220 29338 50254 29372
rect 50320 29338 50354 29372
rect 50420 29338 50454 29372
rect 50520 29338 50554 29372
rect 50620 29338 50654 29372
rect 50720 29338 50754 29372
rect 50220 29238 50254 29272
rect 50320 29238 50354 29272
rect 50420 29238 50454 29272
rect 50520 29238 50554 29272
rect 50620 29238 50654 29272
rect 50720 29238 50754 29272
rect 50220 29140 50254 29172
rect 50320 29140 50354 29172
rect 50420 29140 50454 29172
rect 50220 29138 50242 29140
rect 50242 29138 50254 29140
rect 50320 29138 50332 29140
rect 50332 29138 50354 29140
rect 50420 29138 50422 29140
rect 50422 29138 50454 29140
rect 50520 29138 50554 29172
rect 50620 29138 50654 29172
rect 50720 29140 50754 29172
rect 50720 29138 50748 29140
rect 50748 29138 50754 29140
rect 50220 29050 50254 29072
rect 50320 29050 50354 29072
rect 50420 29050 50454 29072
rect 50220 29038 50242 29050
rect 50242 29038 50254 29050
rect 50320 29038 50332 29050
rect 50332 29038 50354 29050
rect 50420 29038 50422 29050
rect 50422 29038 50454 29050
rect 50520 29038 50554 29072
rect 50620 29038 50654 29072
rect 50720 29050 50754 29072
rect 50720 29038 50748 29050
rect 50748 29038 50754 29050
rect 50220 28960 50254 28972
rect 50320 28960 50354 28972
rect 50420 28960 50454 28972
rect 50220 28938 50242 28960
rect 50242 28938 50254 28960
rect 50320 28938 50332 28960
rect 50332 28938 50354 28960
rect 50420 28938 50422 28960
rect 50422 28938 50454 28960
rect 50520 28938 50554 28972
rect 50620 28938 50654 28972
rect 50720 28960 50754 28972
rect 50720 28938 50748 28960
rect 50748 28938 50754 28960
rect 51374 29642 51408 29676
rect 51464 29674 51498 29676
rect 51554 29674 51588 29676
rect 51644 29674 51678 29676
rect 51734 29674 51768 29676
rect 51824 29674 51858 29676
rect 51914 29674 51948 29676
rect 52004 29674 52038 29676
rect 52094 29674 52128 29676
rect 52184 29674 52218 29676
rect 51464 29642 51484 29674
rect 51484 29642 51498 29674
rect 51554 29642 51574 29674
rect 51574 29642 51588 29674
rect 51644 29642 51664 29674
rect 51664 29642 51678 29674
rect 51734 29642 51754 29674
rect 51754 29642 51768 29674
rect 51824 29642 51844 29674
rect 51844 29642 51858 29674
rect 51914 29642 51934 29674
rect 51934 29642 51948 29674
rect 52004 29642 52024 29674
rect 52024 29642 52038 29674
rect 52094 29642 52114 29674
rect 52114 29642 52128 29674
rect 52184 29642 52204 29674
rect 52204 29642 52218 29674
rect 52274 29642 52308 29676
rect 51560 29466 51582 29472
rect 51582 29466 51594 29472
rect 51660 29466 51672 29472
rect 51672 29466 51694 29472
rect 51760 29466 51762 29472
rect 51762 29466 51794 29472
rect 51560 29438 51594 29466
rect 51660 29438 51694 29466
rect 51760 29438 51794 29466
rect 51860 29438 51894 29472
rect 51960 29438 51994 29472
rect 52060 29466 52088 29472
rect 52088 29466 52094 29472
rect 52060 29438 52094 29466
rect 51560 29338 51594 29372
rect 51660 29338 51694 29372
rect 51760 29338 51794 29372
rect 51860 29338 51894 29372
rect 51960 29338 51994 29372
rect 52060 29338 52094 29372
rect 51560 29238 51594 29272
rect 51660 29238 51694 29272
rect 51760 29238 51794 29272
rect 51860 29238 51894 29272
rect 51960 29238 51994 29272
rect 52060 29238 52094 29272
rect 51560 29140 51594 29172
rect 51660 29140 51694 29172
rect 51760 29140 51794 29172
rect 51560 29138 51582 29140
rect 51582 29138 51594 29140
rect 51660 29138 51672 29140
rect 51672 29138 51694 29140
rect 51760 29138 51762 29140
rect 51762 29138 51794 29140
rect 51860 29138 51894 29172
rect 51960 29138 51994 29172
rect 52060 29140 52094 29172
rect 52060 29138 52088 29140
rect 52088 29138 52094 29140
rect 51560 29050 51594 29072
rect 51660 29050 51694 29072
rect 51760 29050 51794 29072
rect 51560 29038 51582 29050
rect 51582 29038 51594 29050
rect 51660 29038 51672 29050
rect 51672 29038 51694 29050
rect 51760 29038 51762 29050
rect 51762 29038 51794 29050
rect 51860 29038 51894 29072
rect 51960 29038 51994 29072
rect 52060 29050 52094 29072
rect 52060 29038 52088 29050
rect 52088 29038 52094 29050
rect 51560 28960 51594 28972
rect 51660 28960 51694 28972
rect 51760 28960 51794 28972
rect 51560 28938 51582 28960
rect 51582 28938 51594 28960
rect 51660 28938 51672 28960
rect 51672 28938 51694 28960
rect 51760 28938 51762 28960
rect 51762 28938 51794 28960
rect 51860 28938 51894 28972
rect 51960 28938 51994 28972
rect 52060 28960 52094 28972
rect 52060 28938 52088 28960
rect 52088 28938 52094 28960
rect 38577 28373 38611 28407
rect 16703 28255 16737 28289
rect 16903 28255 16937 28289
rect 17103 28255 17137 28289
rect 17303 28255 17337 28289
rect 17503 28255 17537 28289
rect 17703 28255 17737 28289
rect 17903 28255 17937 28289
rect 18103 28255 18137 28289
rect 18303 28255 18337 28289
rect 18503 28255 18537 28289
rect 18703 28255 18737 28289
rect 19447 28255 19481 28289
rect 19647 28255 19681 28289
rect 19847 28255 19881 28289
rect 20047 28255 20081 28289
rect 20247 28255 20281 28289
rect 20447 28255 20481 28289
rect 20647 28255 20681 28289
rect 20847 28255 20881 28289
rect 21047 28255 21081 28289
rect 21247 28255 21281 28289
rect 21447 28255 21481 28289
rect 22191 28255 22225 28289
rect 22391 28255 22425 28289
rect 22591 28255 22625 28289
rect 22791 28255 22825 28289
rect 22991 28255 23025 28289
rect 23191 28255 23225 28289
rect 23391 28255 23425 28289
rect 23591 28255 23625 28289
rect 23791 28255 23825 28289
rect 23991 28255 24025 28289
rect 24191 28255 24225 28289
rect 27385 28255 27419 28289
rect 27585 28255 27619 28289
rect 27785 28255 27819 28289
rect 27985 28255 28019 28289
rect 28185 28255 28219 28289
rect 28385 28255 28419 28289
rect 28585 28255 28619 28289
rect 28785 28255 28819 28289
rect 28985 28255 29019 28289
rect 29185 28255 29219 28289
rect 29385 28255 29419 28289
rect 30111 28255 30145 28289
rect 30511 28255 30545 28289
rect 30911 28255 30945 28289
rect 31311 28255 31345 28289
rect 31711 28255 31745 28289
rect 32111 28255 32145 28289
rect 32511 28255 32545 28289
rect 32911 28255 32945 28289
rect 33311 28255 33345 28289
rect 33711 28255 33745 28289
rect 34111 28255 34145 28289
rect 34511 28255 34545 28289
rect 34911 28255 34945 28289
rect 35311 28255 35345 28289
rect 35711 28255 35745 28289
rect 36111 28255 36145 28289
rect 36511 28255 36545 28289
rect 36911 28255 36945 28289
rect 37655 28255 37689 28289
rect 38055 28255 38089 28289
rect 38455 28255 38489 28289
rect 38855 28255 38889 28289
rect 39255 28255 39289 28289
rect 39655 28255 39689 28289
rect 40055 28255 40089 28289
rect 41967 28255 42001 28289
rect 42167 28255 42201 28289
rect 42367 28255 42401 28289
rect 42567 28255 42601 28289
rect 42767 28255 42801 28289
rect 42967 28255 43001 28289
rect 43167 28255 43201 28289
rect 43367 28255 43401 28289
rect 43567 28255 43601 28289
rect 43767 28255 43801 28289
rect 43967 28255 44001 28289
rect 44167 28255 44201 28289
rect 44367 28255 44401 28289
rect 44567 28255 44601 28289
rect 44767 28255 44801 28289
rect 44967 28255 45001 28289
rect 45167 28255 45201 28289
rect 45367 28255 45401 28289
rect 45567 28255 45601 28289
rect 45767 28255 45801 28289
rect 45967 28255 46001 28289
rect 46167 28255 46201 28289
rect 46367 28255 46401 28289
rect 46567 28255 46601 28289
rect 46767 28255 46801 28289
rect 46967 28255 47001 28289
rect 47167 28255 47201 28289
rect 47367 28255 47401 28289
rect 47567 28255 47601 28289
rect 47767 28255 47801 28289
rect 47967 28255 48001 28289
rect 48167 28255 48201 28289
rect 48367 28255 48401 28289
rect 48567 28255 48601 28289
rect 48767 28255 48801 28289
rect 48967 28255 49001 28289
rect 49167 28255 49201 28289
rect 49367 28255 49401 28289
rect 49567 28255 49601 28289
rect 49767 28255 49801 28289
rect 49967 28255 50001 28289
rect 50167 28255 50201 28289
rect 50367 28255 50401 28289
rect 50567 28255 50601 28289
rect 50767 28255 50801 28289
rect 50967 28255 51001 28289
rect 51167 28255 51201 28289
rect 51367 28255 51401 28289
rect 51567 28255 51601 28289
rect 51767 28255 51801 28289
rect 51967 28255 52001 28289
rect 52167 28255 52201 28289
rect 52367 28255 52401 28289
rect 22583 26375 22617 26409
rect 22783 26375 22817 26409
rect 22983 26375 23017 26409
rect 23183 26375 23217 26409
rect 23383 26375 23417 26409
rect 23583 26375 23617 26409
rect 23783 26375 23817 26409
rect 23983 26375 24017 26409
rect 24183 26375 24217 26409
rect 24383 26375 24417 26409
rect 24583 26375 24617 26409
rect 25601 26375 25635 26409
rect 26001 26375 26035 26409
rect 26401 26375 26435 26409
rect 26801 26375 26835 26409
rect 27201 26375 27235 26409
rect 27601 26375 27635 26409
rect 28001 26375 28035 26409
rect 28401 26375 28435 26409
rect 28801 26375 28835 26409
rect 29201 26375 29235 26409
rect 30111 26375 30145 26409
rect 30511 26375 30545 26409
rect 30911 26375 30945 26409
rect 31311 26375 31345 26409
rect 31711 26375 31745 26409
rect 32111 26375 32145 26409
rect 32511 26375 32545 26409
rect 32911 26375 32945 26409
rect 33311 26375 33345 26409
rect 33711 26375 33745 26409
rect 34111 26375 34145 26409
rect 34511 26375 34545 26409
rect 34911 26375 34945 26409
rect 35311 26375 35345 26409
rect 35711 26375 35745 26409
rect 36111 26375 36145 26409
rect 36511 26375 36545 26409
rect 36911 26375 36945 26409
rect 37577 26375 37611 26409
rect 37777 26375 37811 26409
rect 37977 26375 38011 26409
rect 38177 26375 38211 26409
rect 38377 26375 38411 26409
rect 38577 26375 38611 26409
rect 38777 26375 38811 26409
rect 38977 26375 39011 26409
rect 39177 26375 39211 26409
rect 39377 26375 39411 26409
rect 39577 26375 39611 26409
rect 40321 26375 40355 26409
rect 40521 26375 40555 26409
rect 40721 26375 40755 26409
rect 40921 26375 40955 26409
rect 41121 26375 41155 26409
rect 41321 26375 41355 26409
rect 41521 26375 41555 26409
rect 41721 26375 41755 26409
rect 41921 26375 41955 26409
rect 42121 26375 42155 26409
rect 42321 26375 42355 26409
rect 43065 26375 43099 26409
rect 43265 26375 43299 26409
rect 43465 26375 43499 26409
rect 43665 26375 43699 26409
rect 43865 26375 43899 26409
rect 44065 26375 44099 26409
rect 44265 26375 44299 26409
rect 44465 26375 44499 26409
rect 44665 26375 44699 26409
rect 44865 26375 44899 26409
rect 45065 26375 45099 26409
rect 45809 26375 45843 26409
rect 46009 26375 46043 26409
rect 46209 26375 46243 26409
rect 46409 26375 46443 26409
rect 46609 26375 46643 26409
rect 46809 26375 46843 26409
rect 47009 26375 47043 26409
rect 47209 26375 47243 26409
rect 47409 26375 47443 26409
rect 47609 26375 47643 26409
rect 47809 26375 47843 26409
rect 48553 26375 48587 26409
rect 48753 26375 48787 26409
rect 48953 26375 48987 26409
rect 49153 26375 49187 26409
rect 49353 26375 49387 26409
rect 49553 26375 49587 26409
rect 49753 26375 49787 26409
rect 49953 26375 49987 26409
rect 50153 26375 50187 26409
rect 50353 26375 50387 26409
rect 50553 26375 50587 26409
rect 22419 25603 22813 26141
rect 24426 25603 24820 26141
rect 22419 24643 22813 25181
rect 24426 24643 24820 25181
rect 25430 25869 25464 25889
rect 25430 25855 25464 25869
rect 25430 25801 25464 25817
rect 25430 25783 25464 25801
rect 25430 25733 25464 25745
rect 25430 25711 25464 25733
rect 25430 25665 25464 25673
rect 25430 25639 25464 25665
rect 25430 25597 25464 25601
rect 25430 25567 25464 25597
rect 25430 25495 25464 25529
rect 25430 25427 25464 25457
rect 25430 25423 25464 25427
rect 25430 25359 25464 25385
rect 25430 25351 25464 25359
rect 25430 25291 25464 25313
rect 25430 25279 25464 25291
rect 25430 25223 25464 25241
rect 25430 25207 25464 25223
rect 25430 25155 25464 25169
rect 25430 25135 25464 25155
rect 25888 25869 25922 25889
rect 25888 25855 25922 25869
rect 25888 25801 25922 25817
rect 25888 25783 25922 25801
rect 25888 25733 25922 25745
rect 25888 25711 25922 25733
rect 25888 25665 25922 25673
rect 25888 25639 25922 25665
rect 25888 25597 25922 25601
rect 25888 25567 25922 25597
rect 25888 25495 25922 25529
rect 25888 25427 25922 25457
rect 25888 25423 25922 25427
rect 25888 25359 25922 25385
rect 25888 25351 25922 25359
rect 25888 25291 25922 25313
rect 25888 25279 25922 25291
rect 25888 25223 25922 25241
rect 25888 25207 25922 25223
rect 25888 25155 25922 25169
rect 26346 25869 26380 25889
rect 26346 25855 26380 25869
rect 26346 25801 26380 25817
rect 26346 25783 26380 25801
rect 26346 25733 26380 25745
rect 26346 25711 26380 25733
rect 26346 25665 26380 25673
rect 26346 25639 26380 25665
rect 26346 25597 26380 25601
rect 26346 25567 26380 25597
rect 26346 25495 26380 25529
rect 26346 25427 26380 25457
rect 26346 25423 26380 25427
rect 26346 25359 26380 25385
rect 26346 25351 26380 25359
rect 26346 25291 26380 25313
rect 26346 25279 26380 25291
rect 26346 25223 26380 25241
rect 26346 25207 26380 25223
rect 25888 25135 25922 25155
rect 26346 25155 26380 25169
rect 26346 25135 26380 25155
rect 26804 25869 26838 25889
rect 26804 25855 26838 25869
rect 26804 25801 26838 25817
rect 26804 25783 26838 25801
rect 26804 25733 26838 25745
rect 26804 25711 26838 25733
rect 26804 25665 26838 25673
rect 26804 25639 26838 25665
rect 26804 25597 26838 25601
rect 26804 25567 26838 25597
rect 26804 25495 26838 25529
rect 26804 25427 26838 25457
rect 26804 25423 26838 25427
rect 26804 25359 26838 25385
rect 26804 25351 26838 25359
rect 26804 25291 26838 25313
rect 26804 25279 26838 25291
rect 26804 25223 26838 25241
rect 26804 25207 26838 25223
rect 26804 25155 26838 25169
rect 27262 25869 27296 25889
rect 27262 25855 27296 25869
rect 27262 25801 27296 25817
rect 27262 25783 27296 25801
rect 27262 25733 27296 25745
rect 27262 25711 27296 25733
rect 27262 25665 27296 25673
rect 27262 25639 27296 25665
rect 27262 25597 27296 25601
rect 27262 25567 27296 25597
rect 27262 25495 27296 25529
rect 27262 25427 27296 25457
rect 27262 25423 27296 25427
rect 27262 25359 27296 25385
rect 27262 25351 27296 25359
rect 27262 25291 27296 25313
rect 27262 25279 27296 25291
rect 27262 25223 27296 25241
rect 27262 25207 27296 25223
rect 26804 25135 26838 25155
rect 27262 25155 27296 25169
rect 27262 25135 27296 25155
rect 27720 25869 27754 25889
rect 27720 25855 27754 25869
rect 27720 25801 27754 25817
rect 27720 25783 27754 25801
rect 27720 25733 27754 25745
rect 27720 25711 27754 25733
rect 27720 25665 27754 25673
rect 27720 25639 27754 25665
rect 27720 25597 27754 25601
rect 27720 25567 27754 25597
rect 27720 25495 27754 25529
rect 27720 25427 27754 25457
rect 27720 25423 27754 25427
rect 27720 25359 27754 25385
rect 27720 25351 27754 25359
rect 27720 25291 27754 25313
rect 27720 25279 27754 25291
rect 27720 25223 27754 25241
rect 27720 25207 27754 25223
rect 27720 25155 27754 25169
rect 28178 25869 28212 25889
rect 28178 25855 28212 25869
rect 28178 25801 28212 25817
rect 28178 25783 28212 25801
rect 28178 25733 28212 25745
rect 28178 25711 28212 25733
rect 28178 25665 28212 25673
rect 28178 25639 28212 25665
rect 28178 25597 28212 25601
rect 28178 25567 28212 25597
rect 28178 25495 28212 25529
rect 28178 25427 28212 25457
rect 28178 25423 28212 25427
rect 28178 25359 28212 25385
rect 28178 25351 28212 25359
rect 28178 25291 28212 25313
rect 28178 25279 28212 25291
rect 28178 25223 28212 25241
rect 28178 25207 28212 25223
rect 27720 25135 27754 25155
rect 28178 25155 28212 25169
rect 28178 25135 28212 25155
rect 28636 25869 28670 25889
rect 28636 25855 28670 25869
rect 28636 25801 28670 25817
rect 28636 25783 28670 25801
rect 28636 25733 28670 25745
rect 28636 25711 28670 25733
rect 28636 25665 28670 25673
rect 28636 25639 28670 25665
rect 28636 25597 28670 25601
rect 28636 25567 28670 25597
rect 28636 25495 28670 25529
rect 28636 25427 28670 25457
rect 28636 25423 28670 25427
rect 28636 25359 28670 25385
rect 28636 25351 28670 25359
rect 28636 25291 28670 25313
rect 28636 25279 28670 25291
rect 28636 25223 28670 25241
rect 28636 25207 28670 25223
rect 28636 25155 28670 25169
rect 29094 25869 29128 25889
rect 29094 25855 29128 25869
rect 29094 25801 29128 25817
rect 29094 25783 29128 25801
rect 29094 25733 29128 25745
rect 29094 25711 29128 25733
rect 29094 25665 29128 25673
rect 29094 25639 29128 25665
rect 29094 25597 29128 25601
rect 29094 25567 29128 25597
rect 29094 25495 29128 25529
rect 29094 25427 29128 25457
rect 29094 25423 29128 25427
rect 29094 25359 29128 25385
rect 29094 25351 29128 25359
rect 29094 25291 29128 25313
rect 29094 25279 29128 25291
rect 29094 25223 29128 25241
rect 29094 25207 29128 25223
rect 28636 25135 28670 25155
rect 29094 25155 29128 25169
rect 29094 25135 29128 25155
rect 29552 25869 29586 25889
rect 29552 25855 29586 25869
rect 29552 25801 29586 25817
rect 29552 25783 29586 25801
rect 29552 25733 29586 25745
rect 29552 25711 29586 25733
rect 29552 25665 29586 25673
rect 29552 25639 29586 25665
rect 29552 25597 29586 25601
rect 29552 25567 29586 25597
rect 37413 25603 37807 26141
rect 39420 25603 39814 26141
rect 40157 25603 40551 26141
rect 42164 25603 42558 26141
rect 42901 25603 43295 26141
rect 44908 25603 45302 26141
rect 45645 25603 46039 26141
rect 47652 25603 48046 26141
rect 48389 25603 48783 26141
rect 50396 25603 50790 26141
rect 29552 25495 29586 25529
rect 29552 25427 29586 25457
rect 29552 25423 29586 25427
rect 29552 25359 29586 25385
rect 29552 25351 29586 25359
rect 29552 25291 29586 25313
rect 29552 25279 29586 25291
rect 29552 25223 29586 25241
rect 29552 25207 29586 25223
rect 29552 25155 29586 25169
rect 29552 25135 29586 25155
rect 27537 24837 27571 24871
rect 37413 24643 37807 25181
rect 39420 24643 39814 25181
rect 40157 24643 40551 25181
rect 42164 24643 42558 25181
rect 42901 24643 43295 25181
rect 44908 24643 45302 25181
rect 45645 24643 46039 25181
rect 47652 24643 48046 25181
rect 48389 24643 48783 25181
rect 50396 24643 50790 25181
rect 22583 24495 22617 24529
rect 22783 24495 22817 24529
rect 22983 24495 23017 24529
rect 23183 24495 23217 24529
rect 23383 24495 23417 24529
rect 23583 24495 23617 24529
rect 23783 24495 23817 24529
rect 23983 24495 24017 24529
rect 24183 24495 24217 24529
rect 24383 24495 24417 24529
rect 24583 24495 24617 24529
rect 25601 24495 25635 24529
rect 26001 24495 26035 24529
rect 26401 24495 26435 24529
rect 26801 24495 26835 24529
rect 27201 24495 27235 24529
rect 27601 24495 27635 24529
rect 28001 24495 28035 24529
rect 28401 24495 28435 24529
rect 28801 24495 28835 24529
rect 29201 24495 29235 24529
rect 30111 24495 30145 24529
rect 30511 24495 30545 24529
rect 30911 24495 30945 24529
rect 31311 24495 31345 24529
rect 31711 24495 31745 24529
rect 32111 24495 32145 24529
rect 32511 24495 32545 24529
rect 32911 24495 32945 24529
rect 33311 24495 33345 24529
rect 33711 24495 33745 24529
rect 34111 24495 34145 24529
rect 34511 24495 34545 24529
rect 34911 24495 34945 24529
rect 35311 24495 35345 24529
rect 35711 24495 35745 24529
rect 36111 24495 36145 24529
rect 36511 24495 36545 24529
rect 36911 24495 36945 24529
rect 37577 24495 37611 24529
rect 37777 24495 37811 24529
rect 37977 24495 38011 24529
rect 38177 24495 38211 24529
rect 38377 24495 38411 24529
rect 38577 24495 38611 24529
rect 38777 24495 38811 24529
rect 38977 24495 39011 24529
rect 39177 24495 39211 24529
rect 39377 24495 39411 24529
rect 39577 24495 39611 24529
rect 40321 24495 40355 24529
rect 40521 24495 40555 24529
rect 40721 24495 40755 24529
rect 40921 24495 40955 24529
rect 41121 24495 41155 24529
rect 41321 24495 41355 24529
rect 41521 24495 41555 24529
rect 41721 24495 41755 24529
rect 41921 24495 41955 24529
rect 42121 24495 42155 24529
rect 42321 24495 42355 24529
rect 43065 24495 43099 24529
rect 43265 24495 43299 24529
rect 43465 24495 43499 24529
rect 43665 24495 43699 24529
rect 43865 24495 43899 24529
rect 44065 24495 44099 24529
rect 44265 24495 44299 24529
rect 44465 24495 44499 24529
rect 44665 24495 44699 24529
rect 44865 24495 44899 24529
rect 45065 24495 45099 24529
rect 45809 24495 45843 24529
rect 46009 24495 46043 24529
rect 46209 24495 46243 24529
rect 46409 24495 46443 24529
rect 46609 24495 46643 24529
rect 46809 24495 46843 24529
rect 47009 24495 47043 24529
rect 47209 24495 47243 24529
rect 47409 24495 47443 24529
rect 47609 24495 47643 24529
rect 47809 24495 47843 24529
rect 48553 24495 48587 24529
rect 48753 24495 48787 24529
rect 48953 24495 48987 24529
rect 49153 24495 49187 24529
rect 49353 24495 49387 24529
rect 49553 24495 49587 24529
rect 49753 24495 49787 24529
rect 49953 24495 49987 24529
rect 50153 24495 50187 24529
rect 50353 24495 50387 24529
rect 50553 24495 50587 24529
rect 24053 22615 24087 22649
rect 24253 22615 24287 22649
rect 24453 22615 24487 22649
rect 24653 22615 24687 22649
rect 24853 22615 24887 22649
rect 25053 22615 25087 22649
rect 25253 22615 25287 22649
rect 25453 22615 25487 22649
rect 25653 22615 25687 22649
rect 25853 22615 25887 22649
rect 26053 22615 26087 22649
rect 27385 22615 27419 22649
rect 27585 22615 27619 22649
rect 27785 22615 27819 22649
rect 27985 22615 28019 22649
rect 28185 22615 28219 22649
rect 28385 22615 28419 22649
rect 28585 22615 28619 22649
rect 28785 22615 28819 22649
rect 28985 22615 29019 22649
rect 29185 22615 29219 22649
rect 29385 22615 29419 22649
rect 30129 22615 30163 22649
rect 30329 22615 30363 22649
rect 30529 22615 30563 22649
rect 30729 22615 30763 22649
rect 30929 22615 30963 22649
rect 31129 22615 31163 22649
rect 31329 22615 31363 22649
rect 31529 22615 31563 22649
rect 31729 22615 31763 22649
rect 31929 22615 31963 22649
rect 32129 22615 32163 22649
rect 33363 22615 33397 22649
rect 33563 22615 33597 22649
rect 33763 22615 33797 22649
rect 33963 22615 33997 22649
rect 34163 22615 34197 22649
rect 34363 22615 34397 22649
rect 34563 22615 34597 22649
rect 34763 22615 34797 22649
rect 34963 22615 34997 22649
rect 35163 22615 35197 22649
rect 35363 22615 35397 22649
rect 37577 22615 37611 22649
rect 37777 22615 37811 22649
rect 37977 22615 38011 22649
rect 38177 22615 38211 22649
rect 38377 22615 38411 22649
rect 38577 22615 38611 22649
rect 38777 22615 38811 22649
rect 38977 22615 39011 22649
rect 39177 22615 39211 22649
rect 39377 22615 39411 22649
rect 39577 22615 39611 22649
rect 40321 22615 40355 22649
rect 40521 22615 40555 22649
rect 40721 22615 40755 22649
rect 40921 22615 40955 22649
rect 41121 22615 41155 22649
rect 41321 22615 41355 22649
rect 41521 22615 41555 22649
rect 41721 22615 41755 22649
rect 41921 22615 41955 22649
rect 42121 22615 42155 22649
rect 42321 22615 42355 22649
rect 48553 22615 48587 22649
rect 48753 22615 48787 22649
rect 48953 22615 48987 22649
rect 49153 22615 49187 22649
rect 49353 22615 49387 22649
rect 49553 22615 49587 22649
rect 49753 22615 49787 22649
rect 49953 22615 49987 22649
rect 50153 22615 50187 22649
rect 50353 22615 50387 22649
rect 50553 22615 50587 22649
rect 23889 21843 24283 22381
rect 25896 21843 26290 22381
rect 27221 21843 27615 22381
rect 29228 21843 29622 22381
rect 29965 21843 30359 22381
rect 31972 21843 32366 22381
rect 33199 21843 33593 22381
rect 35206 21843 35600 22381
rect 37413 21843 37807 22381
rect 39420 21843 39814 22381
rect 40157 21843 40551 22381
rect 42164 21843 42558 22381
rect 48389 21843 48783 22381
rect 50396 21843 50790 22381
rect 23889 20883 24283 21421
rect 25896 20883 26290 21421
rect 27221 20883 27615 21421
rect 29228 20883 29622 21421
rect 29965 20883 30359 21421
rect 31972 20883 32366 21421
rect 33199 20883 33593 21421
rect 35206 20883 35600 21421
rect 37413 20883 37807 21421
rect 39420 20883 39814 21421
rect 40157 20883 40551 21421
rect 42164 20883 42558 21421
rect 48389 20883 48783 21421
rect 50396 20883 50790 21421
rect 24053 20735 24087 20769
rect 24253 20735 24287 20769
rect 24453 20735 24487 20769
rect 24653 20735 24687 20769
rect 24853 20735 24887 20769
rect 25053 20735 25087 20769
rect 25253 20735 25287 20769
rect 25453 20735 25487 20769
rect 25653 20735 25687 20769
rect 25853 20735 25887 20769
rect 26053 20735 26087 20769
rect 27385 20735 27419 20769
rect 27585 20735 27619 20769
rect 27785 20735 27819 20769
rect 27985 20735 28019 20769
rect 28185 20735 28219 20769
rect 28385 20735 28419 20769
rect 28585 20735 28619 20769
rect 28785 20735 28819 20769
rect 28985 20735 29019 20769
rect 29185 20735 29219 20769
rect 29385 20735 29419 20769
rect 30129 20735 30163 20769
rect 30329 20735 30363 20769
rect 30529 20735 30563 20769
rect 30729 20735 30763 20769
rect 30929 20735 30963 20769
rect 31129 20735 31163 20769
rect 31329 20735 31363 20769
rect 31529 20735 31563 20769
rect 31729 20735 31763 20769
rect 31929 20735 31963 20769
rect 32129 20735 32163 20769
rect 33363 20735 33397 20769
rect 33563 20735 33597 20769
rect 33763 20735 33797 20769
rect 33963 20735 33997 20769
rect 34163 20735 34197 20769
rect 34363 20735 34397 20769
rect 34563 20735 34597 20769
rect 34763 20735 34797 20769
rect 34963 20735 34997 20769
rect 35163 20735 35197 20769
rect 35363 20735 35397 20769
rect 37577 20735 37611 20769
rect 37777 20735 37811 20769
rect 37977 20735 38011 20769
rect 38177 20735 38211 20769
rect 38377 20735 38411 20769
rect 38577 20735 38611 20769
rect 38777 20735 38811 20769
rect 38977 20735 39011 20769
rect 39177 20735 39211 20769
rect 39377 20735 39411 20769
rect 39577 20735 39611 20769
rect 40321 20735 40355 20769
rect 40521 20735 40555 20769
rect 40721 20735 40755 20769
rect 40921 20735 40955 20769
rect 41121 20735 41155 20769
rect 41321 20735 41355 20769
rect 41521 20735 41555 20769
rect 41721 20735 41755 20769
rect 41921 20735 41955 20769
rect 42121 20735 42155 20769
rect 42321 20735 42355 20769
rect 48553 20735 48587 20769
rect 48753 20735 48787 20769
rect 48953 20735 48987 20769
rect 49153 20735 49187 20769
rect 49353 20735 49387 20769
rect 49553 20735 49587 20769
rect 49753 20735 49787 20769
rect 49953 20735 49987 20769
rect 50153 20735 50187 20769
rect 50353 20735 50387 20769
rect 50553 20735 50587 20769
rect 25013 18855 25047 18889
rect 25413 18855 25447 18889
rect 25813 18855 25847 18889
rect 26213 18855 26247 18889
rect 26613 18855 26647 18889
rect 27013 18855 27047 18889
rect 27413 18855 27447 18889
rect 27813 18855 27847 18889
rect 28213 18855 28247 18889
rect 28613 18855 28647 18889
rect 29013 18855 29047 18889
rect 29413 18855 29447 18889
rect 29813 18855 29847 18889
rect 30213 18855 30247 18889
rect 30613 18855 30647 18889
rect 31013 18855 31047 18889
rect 31413 18855 31447 18889
rect 31813 18855 31847 18889
rect 32213 18855 32247 18889
rect 32613 18855 32647 18889
rect 33013 18855 33047 18889
rect 33413 18855 33447 18889
rect 33813 18855 33847 18889
rect 34213 18855 34247 18889
rect 34613 18855 34647 18889
rect 35013 18855 35047 18889
rect 35413 18855 35447 18889
rect 35813 18855 35847 18889
rect 36213 18855 36247 18889
rect 36613 18855 36647 18889
rect 37013 18855 37047 18889
rect 37413 18855 37447 18889
rect 37813 18855 37847 18889
rect 38213 18855 38247 18889
rect 38613 18855 38647 18889
rect 39013 18855 39047 18889
rect 39413 18855 39447 18889
rect 39813 18855 39847 18889
rect 40213 18855 40247 18889
rect 40613 18855 40647 18889
rect 41013 18855 41047 18889
rect 41413 18855 41447 18889
rect 41813 18855 41847 18889
rect 42213 18855 42247 18889
rect 42613 18855 42647 18889
rect 43013 18855 43047 18889
rect 43413 18855 43447 18889
rect 43813 18855 43847 18889
rect 44213 18855 44247 18889
rect 44613 18855 44647 18889
rect 45013 18855 45047 18889
rect 45413 18855 45447 18889
rect 45813 18855 45847 18889
rect 46213 18855 46247 18889
rect 46613 18855 46647 18889
rect 47013 18855 47047 18889
rect 47413 18855 47447 18889
rect 47813 18855 47847 18889
rect 48213 18855 48247 18889
rect 48613 18855 48647 18889
rect 49013 18855 49047 18889
rect 49413 18855 49447 18889
rect 49813 18855 49847 18889
rect 50213 18855 50247 18889
rect 50613 18855 50647 18889
rect 51013 18855 51047 18889
rect 51413 18855 51447 18889
rect 51813 18855 51847 18889
rect 52213 18855 52247 18889
rect 24877 18587 24911 18621
rect 24877 18519 24911 18549
rect 24877 18515 24911 18519
rect 24877 18451 24911 18477
rect 24877 18443 24911 18451
rect 24877 18383 24911 18405
rect 24877 18371 24911 18383
rect 24877 18315 24911 18333
rect 24877 18299 24911 18315
rect 24877 18247 24911 18261
rect 24877 18227 24911 18247
rect 24877 18179 24911 18189
rect 24877 18155 24911 18179
rect 24877 18111 24911 18117
rect 24877 18083 24911 18111
rect 24877 18043 24911 18045
rect 24877 18011 24911 18043
rect 24877 17941 24911 17973
rect 24877 17939 24911 17941
rect 24877 17873 24911 17901
rect 24877 17867 24911 17873
rect 24877 17805 24911 17829
rect 24877 17795 24911 17805
rect 24877 17737 24911 17757
rect 24877 17723 24911 17737
rect 24877 17669 24911 17685
rect 24877 17651 24911 17669
rect 24877 17601 24911 17613
rect 24877 17579 24911 17601
rect 24877 17533 24911 17541
rect 24877 17507 24911 17533
rect 24877 17465 24911 17469
rect 24877 17435 24911 17465
rect 24877 17363 24911 17397
rect 25335 18587 25369 18621
rect 25335 18519 25369 18549
rect 25335 18515 25369 18519
rect 25335 18451 25369 18477
rect 25335 18443 25369 18451
rect 25335 18383 25369 18405
rect 25335 18371 25369 18383
rect 25335 18315 25369 18333
rect 25335 18299 25369 18315
rect 25335 18247 25369 18261
rect 25335 18227 25369 18247
rect 25335 18179 25369 18189
rect 25335 18155 25369 18179
rect 25335 18111 25369 18117
rect 25335 18083 25369 18111
rect 25335 18043 25369 18045
rect 25335 18011 25369 18043
rect 25335 17941 25369 17973
rect 25335 17939 25369 17941
rect 25335 17873 25369 17901
rect 25335 17867 25369 17873
rect 25335 17805 25369 17829
rect 25335 17795 25369 17805
rect 25335 17737 25369 17757
rect 25335 17723 25369 17737
rect 25335 17669 25369 17685
rect 25335 17651 25369 17669
rect 25335 17601 25369 17613
rect 25335 17579 25369 17601
rect 25335 17533 25369 17541
rect 25335 17507 25369 17533
rect 25335 17465 25369 17469
rect 25335 17435 25369 17465
rect 25335 17363 25369 17397
rect 25793 18587 25827 18621
rect 25793 18519 25827 18549
rect 25793 18515 25827 18519
rect 25793 18451 25827 18477
rect 25793 18443 25827 18451
rect 25793 18383 25827 18405
rect 25793 18371 25827 18383
rect 25793 18315 25827 18333
rect 25793 18299 25827 18315
rect 25793 18247 25827 18261
rect 25793 18227 25827 18247
rect 25793 18179 25827 18189
rect 25793 18155 25827 18179
rect 25793 18111 25827 18117
rect 25793 18083 25827 18111
rect 25793 18043 25827 18045
rect 25793 18011 25827 18043
rect 25793 17941 25827 17973
rect 25793 17939 25827 17941
rect 25793 17873 25827 17901
rect 25793 17867 25827 17873
rect 25793 17805 25827 17829
rect 25793 17795 25827 17805
rect 25793 17737 25827 17757
rect 25793 17723 25827 17737
rect 25793 17669 25827 17685
rect 25793 17651 25827 17669
rect 25793 17601 25827 17613
rect 25793 17579 25827 17601
rect 25793 17533 25827 17541
rect 25793 17507 25827 17533
rect 25793 17465 25827 17469
rect 25793 17435 25827 17465
rect 25793 17363 25827 17397
rect 26251 18587 26285 18621
rect 26251 18519 26285 18549
rect 26251 18515 26285 18519
rect 26251 18451 26285 18477
rect 26251 18443 26285 18451
rect 26251 18383 26285 18405
rect 26251 18371 26285 18383
rect 26251 18315 26285 18333
rect 26251 18299 26285 18315
rect 26251 18247 26285 18261
rect 26251 18227 26285 18247
rect 26251 18179 26285 18189
rect 26251 18155 26285 18179
rect 26251 18111 26285 18117
rect 26251 18083 26285 18111
rect 26251 18043 26285 18045
rect 26251 18011 26285 18043
rect 26251 17941 26285 17973
rect 26251 17939 26285 17941
rect 26251 17873 26285 17901
rect 26251 17867 26285 17873
rect 26251 17805 26285 17829
rect 26251 17795 26285 17805
rect 26251 17737 26285 17757
rect 26251 17723 26285 17737
rect 26251 17669 26285 17685
rect 26251 17651 26285 17669
rect 26251 17601 26285 17613
rect 26251 17579 26285 17601
rect 26251 17533 26285 17541
rect 26251 17507 26285 17533
rect 26251 17465 26285 17469
rect 26251 17435 26285 17465
rect 26251 17363 26285 17397
rect 26709 18587 26743 18621
rect 26709 18519 26743 18549
rect 26709 18515 26743 18519
rect 26709 18451 26743 18477
rect 26709 18443 26743 18451
rect 26709 18383 26743 18405
rect 26709 18371 26743 18383
rect 26709 18315 26743 18333
rect 26709 18299 26743 18315
rect 26709 18247 26743 18261
rect 26709 18227 26743 18247
rect 26709 18179 26743 18189
rect 26709 18155 26743 18179
rect 26709 18111 26743 18117
rect 26709 18083 26743 18111
rect 26709 18043 26743 18045
rect 26709 18011 26743 18043
rect 26709 17941 26743 17973
rect 26709 17939 26743 17941
rect 26709 17873 26743 17901
rect 26709 17867 26743 17873
rect 26709 17805 26743 17829
rect 26709 17795 26743 17805
rect 26709 17737 26743 17757
rect 26709 17723 26743 17737
rect 26709 17669 26743 17685
rect 26709 17651 26743 17669
rect 26709 17601 26743 17613
rect 26709 17579 26743 17601
rect 26709 17533 26743 17541
rect 26709 17507 26743 17533
rect 26709 17465 26743 17469
rect 26709 17435 26743 17465
rect 26709 17363 26743 17397
rect 27167 18587 27201 18621
rect 27167 18519 27201 18549
rect 27167 18515 27201 18519
rect 27167 18451 27201 18477
rect 27167 18443 27201 18451
rect 27167 18383 27201 18405
rect 27167 18371 27201 18383
rect 27167 18315 27201 18333
rect 27167 18299 27201 18315
rect 27167 18247 27201 18261
rect 27167 18227 27201 18247
rect 27167 18179 27201 18189
rect 27167 18155 27201 18179
rect 27167 18111 27201 18117
rect 27167 18083 27201 18111
rect 27167 18043 27201 18045
rect 27167 18011 27201 18043
rect 27167 17941 27201 17973
rect 27167 17939 27201 17941
rect 27167 17873 27201 17901
rect 27167 17867 27201 17873
rect 27167 17805 27201 17829
rect 27167 17795 27201 17805
rect 27167 17737 27201 17757
rect 27167 17723 27201 17737
rect 27167 17669 27201 17685
rect 27167 17651 27201 17669
rect 27167 17601 27201 17613
rect 27167 17579 27201 17601
rect 27167 17533 27201 17541
rect 27167 17507 27201 17533
rect 27167 17465 27201 17469
rect 27167 17435 27201 17465
rect 27167 17363 27201 17397
rect 27625 18587 27659 18621
rect 27625 18519 27659 18549
rect 27625 18515 27659 18519
rect 27625 18451 27659 18477
rect 27625 18443 27659 18451
rect 27625 18383 27659 18405
rect 27625 18371 27659 18383
rect 27625 18315 27659 18333
rect 27625 18299 27659 18315
rect 27625 18247 27659 18261
rect 27625 18227 27659 18247
rect 27625 18179 27659 18189
rect 27625 18155 27659 18179
rect 27625 18111 27659 18117
rect 27625 18083 27659 18111
rect 27625 18043 27659 18045
rect 27625 18011 27659 18043
rect 27625 17941 27659 17973
rect 27625 17939 27659 17941
rect 27625 17873 27659 17901
rect 27625 17867 27659 17873
rect 27625 17805 27659 17829
rect 27625 17795 27659 17805
rect 27625 17737 27659 17757
rect 27625 17723 27659 17737
rect 27625 17669 27659 17685
rect 27625 17651 27659 17669
rect 27625 17601 27659 17613
rect 27625 17579 27659 17601
rect 27625 17533 27659 17541
rect 27625 17507 27659 17533
rect 27625 17465 27659 17469
rect 27625 17435 27659 17465
rect 27625 17363 27659 17397
rect 28083 18587 28117 18621
rect 28083 18519 28117 18549
rect 28083 18515 28117 18519
rect 28083 18451 28117 18477
rect 28083 18443 28117 18451
rect 28083 18383 28117 18405
rect 28083 18371 28117 18383
rect 28083 18315 28117 18333
rect 28083 18299 28117 18315
rect 28083 18247 28117 18261
rect 28083 18227 28117 18247
rect 28083 18179 28117 18189
rect 28083 18155 28117 18179
rect 28083 18111 28117 18117
rect 28083 18083 28117 18111
rect 28083 18043 28117 18045
rect 28083 18011 28117 18043
rect 28083 17941 28117 17973
rect 28083 17939 28117 17941
rect 28083 17873 28117 17901
rect 28083 17867 28117 17873
rect 28083 17805 28117 17829
rect 28083 17795 28117 17805
rect 28083 17737 28117 17757
rect 28083 17723 28117 17737
rect 28083 17669 28117 17685
rect 28083 17651 28117 17669
rect 28083 17601 28117 17613
rect 28083 17579 28117 17601
rect 28083 17533 28117 17541
rect 28083 17507 28117 17533
rect 28083 17465 28117 17469
rect 28083 17435 28117 17465
rect 28083 17363 28117 17397
rect 28541 18587 28575 18621
rect 28541 18519 28575 18549
rect 28541 18515 28575 18519
rect 28541 18451 28575 18477
rect 28541 18443 28575 18451
rect 28541 18383 28575 18405
rect 28541 18371 28575 18383
rect 28541 18315 28575 18333
rect 28541 18299 28575 18315
rect 28541 18247 28575 18261
rect 28541 18227 28575 18247
rect 28541 18179 28575 18189
rect 28541 18155 28575 18179
rect 28541 18111 28575 18117
rect 28541 18083 28575 18111
rect 28541 18043 28575 18045
rect 28541 18011 28575 18043
rect 28541 17941 28575 17973
rect 28541 17939 28575 17941
rect 28541 17873 28575 17901
rect 28541 17867 28575 17873
rect 28541 17805 28575 17829
rect 28541 17795 28575 17805
rect 28541 17737 28575 17757
rect 28541 17723 28575 17737
rect 28541 17669 28575 17685
rect 28541 17651 28575 17669
rect 28541 17601 28575 17613
rect 28541 17579 28575 17601
rect 28541 17533 28575 17541
rect 28541 17507 28575 17533
rect 28541 17465 28575 17469
rect 28541 17435 28575 17465
rect 28541 17363 28575 17397
rect 28999 18587 29033 18621
rect 28999 18519 29033 18549
rect 28999 18515 29033 18519
rect 28999 18451 29033 18477
rect 28999 18443 29033 18451
rect 28999 18383 29033 18405
rect 28999 18371 29033 18383
rect 28999 18315 29033 18333
rect 28999 18299 29033 18315
rect 28999 18247 29033 18261
rect 28999 18227 29033 18247
rect 28999 18179 29033 18189
rect 28999 18155 29033 18179
rect 28999 18111 29033 18117
rect 28999 18083 29033 18111
rect 28999 18043 29033 18045
rect 28999 18011 29033 18043
rect 28999 17941 29033 17973
rect 28999 17939 29033 17941
rect 28999 17873 29033 17901
rect 28999 17867 29033 17873
rect 28999 17805 29033 17829
rect 28999 17795 29033 17805
rect 28999 17737 29033 17757
rect 28999 17723 29033 17737
rect 28999 17669 29033 17685
rect 28999 17651 29033 17669
rect 28999 17601 29033 17613
rect 28999 17579 29033 17601
rect 28999 17533 29033 17541
rect 28999 17507 29033 17533
rect 28999 17465 29033 17469
rect 28999 17435 29033 17465
rect 28999 17363 29033 17397
rect 29457 18587 29491 18621
rect 29457 18519 29491 18549
rect 29457 18515 29491 18519
rect 29457 18451 29491 18477
rect 29457 18443 29491 18451
rect 29457 18383 29491 18405
rect 29457 18371 29491 18383
rect 29457 18315 29491 18333
rect 29457 18299 29491 18315
rect 29457 18247 29491 18261
rect 29457 18227 29491 18247
rect 29457 18179 29491 18189
rect 29457 18155 29491 18179
rect 29457 18111 29491 18117
rect 29457 18083 29491 18111
rect 29457 18043 29491 18045
rect 29457 18011 29491 18043
rect 29457 17941 29491 17973
rect 29457 17939 29491 17941
rect 29457 17873 29491 17901
rect 29457 17867 29491 17873
rect 29457 17805 29491 17829
rect 29457 17795 29491 17805
rect 29457 17737 29491 17757
rect 29457 17723 29491 17737
rect 29457 17669 29491 17685
rect 29457 17651 29491 17669
rect 29457 17601 29491 17613
rect 29457 17579 29491 17601
rect 29457 17533 29491 17541
rect 29457 17507 29491 17533
rect 29457 17465 29491 17469
rect 29457 17435 29491 17465
rect 29457 17363 29491 17397
rect 29915 18587 29949 18621
rect 29915 18519 29949 18549
rect 29915 18515 29949 18519
rect 29915 18451 29949 18477
rect 29915 18443 29949 18451
rect 29915 18383 29949 18405
rect 29915 18371 29949 18383
rect 29915 18315 29949 18333
rect 29915 18299 29949 18315
rect 29915 18247 29949 18261
rect 29915 18227 29949 18247
rect 29915 18179 29949 18189
rect 29915 18155 29949 18179
rect 29915 18111 29949 18117
rect 29915 18083 29949 18111
rect 29915 18043 29949 18045
rect 29915 18011 29949 18043
rect 29915 17941 29949 17973
rect 29915 17939 29949 17941
rect 29915 17873 29949 17901
rect 29915 17867 29949 17873
rect 29915 17805 29949 17829
rect 29915 17795 29949 17805
rect 29915 17737 29949 17757
rect 29915 17723 29949 17737
rect 29915 17669 29949 17685
rect 29915 17651 29949 17669
rect 29915 17601 29949 17613
rect 29915 17579 29949 17601
rect 29915 17533 29949 17541
rect 29915 17507 29949 17533
rect 29915 17465 29949 17469
rect 29915 17435 29949 17465
rect 29915 17363 29949 17397
rect 30373 18587 30407 18621
rect 30373 18519 30407 18549
rect 30373 18515 30407 18519
rect 30373 18451 30407 18477
rect 30373 18443 30407 18451
rect 30373 18383 30407 18405
rect 30373 18371 30407 18383
rect 30373 18315 30407 18333
rect 30373 18299 30407 18315
rect 30373 18247 30407 18261
rect 30373 18227 30407 18247
rect 30373 18179 30407 18189
rect 30373 18155 30407 18179
rect 30373 18111 30407 18117
rect 30373 18083 30407 18111
rect 30373 18043 30407 18045
rect 30373 18011 30407 18043
rect 30373 17941 30407 17973
rect 30373 17939 30407 17941
rect 30373 17873 30407 17901
rect 30373 17867 30407 17873
rect 30373 17805 30407 17829
rect 30373 17795 30407 17805
rect 30373 17737 30407 17757
rect 30373 17723 30407 17737
rect 30373 17669 30407 17685
rect 30373 17651 30407 17669
rect 30373 17601 30407 17613
rect 30373 17579 30407 17601
rect 30373 17533 30407 17541
rect 30373 17507 30407 17533
rect 30373 17465 30407 17469
rect 30373 17435 30407 17465
rect 30373 17363 30407 17397
rect 30831 18587 30865 18621
rect 30831 18519 30865 18549
rect 30831 18515 30865 18519
rect 30831 18451 30865 18477
rect 30831 18443 30865 18451
rect 30831 18383 30865 18405
rect 30831 18371 30865 18383
rect 30831 18315 30865 18333
rect 30831 18299 30865 18315
rect 30831 18247 30865 18261
rect 30831 18227 30865 18247
rect 30831 18179 30865 18189
rect 30831 18155 30865 18179
rect 30831 18111 30865 18117
rect 30831 18083 30865 18111
rect 30831 18043 30865 18045
rect 30831 18011 30865 18043
rect 30831 17941 30865 17973
rect 30831 17939 30865 17941
rect 30831 17873 30865 17901
rect 30831 17867 30865 17873
rect 30831 17805 30865 17829
rect 30831 17795 30865 17805
rect 30831 17737 30865 17757
rect 30831 17723 30865 17737
rect 30831 17669 30865 17685
rect 30831 17651 30865 17669
rect 30831 17601 30865 17613
rect 30831 17579 30865 17601
rect 30831 17533 30865 17541
rect 30831 17507 30865 17533
rect 30831 17465 30865 17469
rect 30831 17435 30865 17465
rect 30831 17363 30865 17397
rect 31289 18587 31323 18621
rect 31289 18519 31323 18549
rect 31289 18515 31323 18519
rect 31289 18451 31323 18477
rect 31289 18443 31323 18451
rect 31289 18383 31323 18405
rect 31289 18371 31323 18383
rect 31289 18315 31323 18333
rect 31289 18299 31323 18315
rect 31289 18247 31323 18261
rect 31289 18227 31323 18247
rect 31289 18179 31323 18189
rect 31289 18155 31323 18179
rect 31289 18111 31323 18117
rect 31289 18083 31323 18111
rect 31289 18043 31323 18045
rect 31289 18011 31323 18043
rect 31289 17941 31323 17973
rect 31289 17939 31323 17941
rect 31289 17873 31323 17901
rect 31289 17867 31323 17873
rect 31289 17805 31323 17829
rect 31289 17795 31323 17805
rect 31289 17737 31323 17757
rect 31289 17723 31323 17737
rect 31289 17669 31323 17685
rect 31289 17651 31323 17669
rect 31289 17601 31323 17613
rect 31289 17579 31323 17601
rect 31289 17533 31323 17541
rect 31289 17507 31323 17533
rect 31289 17465 31323 17469
rect 31289 17435 31323 17465
rect 31289 17363 31323 17397
rect 31747 18587 31781 18621
rect 31747 18519 31781 18549
rect 31747 18515 31781 18519
rect 31747 18451 31781 18477
rect 31747 18443 31781 18451
rect 31747 18383 31781 18405
rect 31747 18371 31781 18383
rect 31747 18315 31781 18333
rect 31747 18299 31781 18315
rect 31747 18247 31781 18261
rect 31747 18227 31781 18247
rect 31747 18179 31781 18189
rect 31747 18155 31781 18179
rect 31747 18111 31781 18117
rect 31747 18083 31781 18111
rect 31747 18043 31781 18045
rect 31747 18011 31781 18043
rect 31747 17941 31781 17973
rect 31747 17939 31781 17941
rect 31747 17873 31781 17901
rect 31747 17867 31781 17873
rect 31747 17805 31781 17829
rect 31747 17795 31781 17805
rect 31747 17737 31781 17757
rect 31747 17723 31781 17737
rect 31747 17669 31781 17685
rect 31747 17651 31781 17669
rect 31747 17601 31781 17613
rect 31747 17579 31781 17601
rect 31747 17533 31781 17541
rect 31747 17507 31781 17533
rect 31747 17465 31781 17469
rect 31747 17435 31781 17465
rect 31747 17363 31781 17397
rect 32205 18587 32239 18621
rect 32205 18519 32239 18549
rect 32205 18515 32239 18519
rect 32205 18451 32239 18477
rect 32205 18443 32239 18451
rect 32205 18383 32239 18405
rect 32205 18371 32239 18383
rect 32205 18315 32239 18333
rect 32205 18299 32239 18315
rect 32205 18247 32239 18261
rect 32205 18227 32239 18247
rect 32205 18179 32239 18189
rect 32205 18155 32239 18179
rect 32205 18111 32239 18117
rect 32205 18083 32239 18111
rect 32205 18043 32239 18045
rect 32205 18011 32239 18043
rect 32205 17941 32239 17973
rect 32205 17939 32239 17941
rect 32205 17873 32239 17901
rect 32205 17867 32239 17873
rect 32205 17805 32239 17829
rect 32205 17795 32239 17805
rect 32205 17737 32239 17757
rect 32205 17723 32239 17737
rect 32205 17669 32239 17685
rect 32205 17651 32239 17669
rect 32205 17601 32239 17613
rect 32205 17579 32239 17601
rect 32205 17533 32239 17541
rect 32205 17507 32239 17533
rect 32205 17465 32239 17469
rect 32205 17435 32239 17465
rect 32205 17363 32239 17397
rect 32663 18587 32697 18621
rect 32663 18519 32697 18549
rect 32663 18515 32697 18519
rect 32663 18451 32697 18477
rect 32663 18443 32697 18451
rect 32663 18383 32697 18405
rect 32663 18371 32697 18383
rect 32663 18315 32697 18333
rect 32663 18299 32697 18315
rect 32663 18247 32697 18261
rect 32663 18227 32697 18247
rect 32663 18179 32697 18189
rect 32663 18155 32697 18179
rect 32663 18111 32697 18117
rect 32663 18083 32697 18111
rect 32663 18043 32697 18045
rect 32663 18011 32697 18043
rect 32663 17941 32697 17973
rect 32663 17939 32697 17941
rect 32663 17873 32697 17901
rect 32663 17867 32697 17873
rect 32663 17805 32697 17829
rect 32663 17795 32697 17805
rect 32663 17737 32697 17757
rect 32663 17723 32697 17737
rect 32663 17669 32697 17685
rect 32663 17651 32697 17669
rect 32663 17601 32697 17613
rect 32663 17579 32697 17601
rect 32663 17533 32697 17541
rect 32663 17507 32697 17533
rect 32663 17465 32697 17469
rect 32663 17435 32697 17465
rect 32663 17363 32697 17397
rect 33121 18587 33155 18621
rect 33121 18519 33155 18549
rect 33121 18515 33155 18519
rect 33121 18451 33155 18477
rect 33121 18443 33155 18451
rect 33121 18383 33155 18405
rect 33121 18371 33155 18383
rect 33121 18315 33155 18333
rect 33121 18299 33155 18315
rect 33121 18247 33155 18261
rect 33121 18227 33155 18247
rect 33121 18179 33155 18189
rect 33121 18155 33155 18179
rect 33121 18111 33155 18117
rect 33121 18083 33155 18111
rect 33121 18043 33155 18045
rect 33121 18011 33155 18043
rect 33121 17941 33155 17973
rect 33121 17939 33155 17941
rect 33121 17873 33155 17901
rect 33121 17867 33155 17873
rect 33121 17805 33155 17829
rect 33121 17795 33155 17805
rect 33121 17737 33155 17757
rect 33121 17723 33155 17737
rect 33121 17669 33155 17685
rect 33121 17651 33155 17669
rect 33121 17601 33155 17613
rect 33121 17579 33155 17601
rect 33121 17533 33155 17541
rect 33121 17507 33155 17533
rect 33121 17465 33155 17469
rect 33121 17435 33155 17465
rect 33121 17363 33155 17397
rect 33579 18587 33613 18621
rect 33579 18519 33613 18549
rect 33579 18515 33613 18519
rect 33579 18451 33613 18477
rect 33579 18443 33613 18451
rect 33579 18383 33613 18405
rect 33579 18371 33613 18383
rect 33579 18315 33613 18333
rect 33579 18299 33613 18315
rect 33579 18247 33613 18261
rect 33579 18227 33613 18247
rect 33579 18179 33613 18189
rect 33579 18155 33613 18179
rect 33579 18111 33613 18117
rect 33579 18083 33613 18111
rect 33579 18043 33613 18045
rect 33579 18011 33613 18043
rect 33579 17941 33613 17973
rect 33579 17939 33613 17941
rect 33579 17873 33613 17901
rect 33579 17867 33613 17873
rect 33579 17805 33613 17829
rect 33579 17795 33613 17805
rect 33579 17737 33613 17757
rect 33579 17723 33613 17737
rect 33579 17669 33613 17685
rect 33579 17651 33613 17669
rect 33579 17601 33613 17613
rect 33579 17579 33613 17601
rect 33579 17533 33613 17541
rect 33579 17507 33613 17533
rect 33579 17465 33613 17469
rect 33579 17435 33613 17465
rect 33579 17363 33613 17397
rect 34037 18587 34071 18621
rect 34037 18519 34071 18549
rect 34037 18515 34071 18519
rect 34037 18451 34071 18477
rect 34037 18443 34071 18451
rect 34037 18383 34071 18405
rect 34037 18371 34071 18383
rect 34037 18315 34071 18333
rect 34037 18299 34071 18315
rect 34037 18247 34071 18261
rect 34037 18227 34071 18247
rect 34037 18179 34071 18189
rect 34037 18155 34071 18179
rect 34037 18111 34071 18117
rect 34037 18083 34071 18111
rect 34037 18043 34071 18045
rect 34037 18011 34071 18043
rect 34037 17941 34071 17973
rect 34037 17939 34071 17941
rect 34037 17873 34071 17901
rect 34037 17867 34071 17873
rect 34037 17805 34071 17829
rect 34037 17795 34071 17805
rect 34037 17737 34071 17757
rect 34037 17723 34071 17737
rect 34037 17669 34071 17685
rect 34037 17651 34071 17669
rect 34037 17601 34071 17613
rect 34037 17579 34071 17601
rect 34037 17533 34071 17541
rect 34037 17507 34071 17533
rect 34037 17465 34071 17469
rect 34037 17435 34071 17465
rect 34037 17363 34071 17397
rect 34495 18587 34529 18621
rect 34495 18519 34529 18549
rect 34495 18515 34529 18519
rect 34495 18451 34529 18477
rect 34495 18443 34529 18451
rect 34495 18383 34529 18405
rect 34495 18371 34529 18383
rect 34495 18315 34529 18333
rect 34495 18299 34529 18315
rect 34495 18247 34529 18261
rect 34495 18227 34529 18247
rect 34495 18179 34529 18189
rect 34495 18155 34529 18179
rect 34495 18111 34529 18117
rect 34495 18083 34529 18111
rect 34495 18043 34529 18045
rect 34495 18011 34529 18043
rect 34495 17941 34529 17973
rect 34495 17939 34529 17941
rect 34495 17873 34529 17901
rect 34495 17867 34529 17873
rect 34495 17805 34529 17829
rect 34495 17795 34529 17805
rect 34495 17737 34529 17757
rect 34495 17723 34529 17737
rect 34495 17669 34529 17685
rect 34495 17651 34529 17669
rect 34495 17601 34529 17613
rect 34495 17579 34529 17601
rect 34495 17533 34529 17541
rect 34495 17507 34529 17533
rect 34495 17465 34529 17469
rect 34495 17435 34529 17465
rect 34495 17363 34529 17397
rect 34953 18587 34987 18621
rect 34953 18519 34987 18549
rect 34953 18515 34987 18519
rect 34953 18451 34987 18477
rect 34953 18443 34987 18451
rect 34953 18383 34987 18405
rect 34953 18371 34987 18383
rect 34953 18315 34987 18333
rect 34953 18299 34987 18315
rect 34953 18247 34987 18261
rect 34953 18227 34987 18247
rect 34953 18179 34987 18189
rect 34953 18155 34987 18179
rect 34953 18111 34987 18117
rect 34953 18083 34987 18111
rect 34953 18043 34987 18045
rect 34953 18011 34987 18043
rect 34953 17941 34987 17973
rect 34953 17939 34987 17941
rect 34953 17873 34987 17901
rect 34953 17867 34987 17873
rect 34953 17805 34987 17829
rect 34953 17795 34987 17805
rect 34953 17737 34987 17757
rect 34953 17723 34987 17737
rect 34953 17669 34987 17685
rect 34953 17651 34987 17669
rect 34953 17601 34987 17613
rect 34953 17579 34987 17601
rect 34953 17533 34987 17541
rect 34953 17507 34987 17533
rect 34953 17465 34987 17469
rect 34953 17435 34987 17465
rect 34953 17363 34987 17397
rect 35411 18587 35445 18621
rect 35411 18519 35445 18549
rect 35411 18515 35445 18519
rect 35411 18451 35445 18477
rect 35411 18443 35445 18451
rect 35411 18383 35445 18405
rect 35411 18371 35445 18383
rect 35411 18315 35445 18333
rect 35411 18299 35445 18315
rect 35411 18247 35445 18261
rect 35411 18227 35445 18247
rect 35411 18179 35445 18189
rect 35411 18155 35445 18179
rect 35411 18111 35445 18117
rect 35411 18083 35445 18111
rect 35411 18043 35445 18045
rect 35411 18011 35445 18043
rect 35411 17941 35445 17973
rect 35411 17939 35445 17941
rect 35411 17873 35445 17901
rect 35411 17867 35445 17873
rect 35411 17805 35445 17829
rect 35411 17795 35445 17805
rect 35411 17737 35445 17757
rect 35411 17723 35445 17737
rect 35411 17669 35445 17685
rect 35411 17651 35445 17669
rect 35411 17601 35445 17613
rect 35411 17579 35445 17601
rect 35411 17533 35445 17541
rect 35411 17507 35445 17533
rect 35411 17465 35445 17469
rect 35411 17435 35445 17465
rect 35411 17363 35445 17397
rect 35869 18587 35903 18621
rect 35869 18519 35903 18549
rect 35869 18515 35903 18519
rect 35869 18451 35903 18477
rect 35869 18443 35903 18451
rect 35869 18383 35903 18405
rect 35869 18371 35903 18383
rect 35869 18315 35903 18333
rect 35869 18299 35903 18315
rect 35869 18247 35903 18261
rect 35869 18227 35903 18247
rect 35869 18179 35903 18189
rect 35869 18155 35903 18179
rect 35869 18111 35903 18117
rect 35869 18083 35903 18111
rect 35869 18043 35903 18045
rect 35869 18011 35903 18043
rect 35869 17941 35903 17973
rect 35869 17939 35903 17941
rect 35869 17873 35903 17901
rect 35869 17867 35903 17873
rect 35869 17805 35903 17829
rect 35869 17795 35903 17805
rect 35869 17737 35903 17757
rect 35869 17723 35903 17737
rect 35869 17669 35903 17685
rect 35869 17651 35903 17669
rect 35869 17601 35903 17613
rect 35869 17579 35903 17601
rect 35869 17533 35903 17541
rect 35869 17507 35903 17533
rect 35869 17465 35903 17469
rect 35869 17435 35903 17465
rect 35869 17363 35903 17397
rect 36327 18587 36361 18621
rect 36327 18519 36361 18549
rect 36327 18515 36361 18519
rect 36327 18451 36361 18477
rect 36327 18443 36361 18451
rect 36327 18383 36361 18405
rect 36327 18371 36361 18383
rect 36327 18315 36361 18333
rect 36327 18299 36361 18315
rect 36327 18247 36361 18261
rect 36327 18227 36361 18247
rect 36327 18179 36361 18189
rect 36327 18155 36361 18179
rect 36327 18111 36361 18117
rect 36327 18083 36361 18111
rect 36327 18043 36361 18045
rect 36327 18011 36361 18043
rect 36327 17941 36361 17973
rect 36327 17939 36361 17941
rect 36327 17873 36361 17901
rect 36327 17867 36361 17873
rect 36327 17805 36361 17829
rect 36327 17795 36361 17805
rect 36327 17737 36361 17757
rect 36327 17723 36361 17737
rect 36327 17669 36361 17685
rect 36327 17651 36361 17669
rect 36327 17601 36361 17613
rect 36327 17579 36361 17601
rect 36327 17533 36361 17541
rect 36327 17507 36361 17533
rect 36327 17465 36361 17469
rect 36327 17435 36361 17465
rect 36327 17363 36361 17397
rect 36785 18587 36819 18621
rect 36785 18519 36819 18549
rect 36785 18515 36819 18519
rect 36785 18451 36819 18477
rect 36785 18443 36819 18451
rect 36785 18383 36819 18405
rect 36785 18371 36819 18383
rect 36785 18315 36819 18333
rect 36785 18299 36819 18315
rect 36785 18247 36819 18261
rect 36785 18227 36819 18247
rect 36785 18179 36819 18189
rect 36785 18155 36819 18179
rect 36785 18111 36819 18117
rect 36785 18083 36819 18111
rect 36785 18043 36819 18045
rect 36785 18011 36819 18043
rect 36785 17941 36819 17973
rect 36785 17939 36819 17941
rect 36785 17873 36819 17901
rect 36785 17867 36819 17873
rect 36785 17805 36819 17829
rect 36785 17795 36819 17805
rect 36785 17737 36819 17757
rect 36785 17723 36819 17737
rect 36785 17669 36819 17685
rect 36785 17651 36819 17669
rect 36785 17601 36819 17613
rect 36785 17579 36819 17601
rect 36785 17533 36819 17541
rect 36785 17507 36819 17533
rect 36785 17465 36819 17469
rect 36785 17435 36819 17465
rect 36785 17363 36819 17397
rect 37243 18587 37277 18621
rect 37243 18519 37277 18549
rect 37243 18515 37277 18519
rect 37243 18451 37277 18477
rect 37243 18443 37277 18451
rect 37243 18383 37277 18405
rect 37243 18371 37277 18383
rect 37243 18315 37277 18333
rect 37243 18299 37277 18315
rect 37243 18247 37277 18261
rect 37243 18227 37277 18247
rect 37243 18179 37277 18189
rect 37243 18155 37277 18179
rect 37243 18111 37277 18117
rect 37243 18083 37277 18111
rect 37243 18043 37277 18045
rect 37243 18011 37277 18043
rect 37243 17941 37277 17973
rect 37243 17939 37277 17941
rect 37243 17873 37277 17901
rect 37243 17867 37277 17873
rect 37243 17805 37277 17829
rect 37243 17795 37277 17805
rect 37243 17737 37277 17757
rect 37243 17723 37277 17737
rect 37243 17669 37277 17685
rect 37243 17651 37277 17669
rect 37243 17601 37277 17613
rect 37243 17579 37277 17601
rect 37243 17533 37277 17541
rect 37243 17507 37277 17533
rect 37243 17465 37277 17469
rect 37243 17435 37277 17465
rect 37243 17363 37277 17397
rect 37701 18587 37735 18621
rect 37701 18519 37735 18549
rect 37701 18515 37735 18519
rect 37701 18451 37735 18477
rect 37701 18443 37735 18451
rect 37701 18383 37735 18405
rect 37701 18371 37735 18383
rect 37701 18315 37735 18333
rect 37701 18299 37735 18315
rect 37701 18247 37735 18261
rect 37701 18227 37735 18247
rect 37701 18179 37735 18189
rect 37701 18155 37735 18179
rect 37701 18111 37735 18117
rect 37701 18083 37735 18111
rect 37701 18043 37735 18045
rect 37701 18011 37735 18043
rect 37701 17941 37735 17973
rect 37701 17939 37735 17941
rect 37701 17873 37735 17901
rect 37701 17867 37735 17873
rect 37701 17805 37735 17829
rect 37701 17795 37735 17805
rect 37701 17737 37735 17757
rect 37701 17723 37735 17737
rect 37701 17669 37735 17685
rect 37701 17651 37735 17669
rect 37701 17601 37735 17613
rect 37701 17579 37735 17601
rect 37701 17533 37735 17541
rect 37701 17507 37735 17533
rect 37701 17465 37735 17469
rect 37701 17435 37735 17465
rect 37701 17363 37735 17397
rect 38159 18587 38193 18621
rect 38159 18519 38193 18549
rect 38159 18515 38193 18519
rect 38159 18451 38193 18477
rect 38159 18443 38193 18451
rect 38159 18383 38193 18405
rect 38159 18371 38193 18383
rect 38159 18315 38193 18333
rect 38159 18299 38193 18315
rect 38159 18247 38193 18261
rect 38159 18227 38193 18247
rect 38159 18179 38193 18189
rect 38159 18155 38193 18179
rect 38159 18111 38193 18117
rect 38159 18083 38193 18111
rect 38159 18043 38193 18045
rect 38159 18011 38193 18043
rect 38159 17941 38193 17973
rect 38159 17939 38193 17941
rect 38159 17873 38193 17901
rect 38159 17867 38193 17873
rect 38159 17805 38193 17829
rect 38159 17795 38193 17805
rect 38159 17737 38193 17757
rect 38159 17723 38193 17737
rect 38159 17669 38193 17685
rect 38159 17651 38193 17669
rect 38159 17601 38193 17613
rect 38159 17579 38193 17601
rect 38159 17533 38193 17541
rect 38159 17507 38193 17533
rect 38159 17465 38193 17469
rect 38159 17435 38193 17465
rect 38159 17363 38193 17397
rect 38617 18587 38651 18621
rect 38617 18519 38651 18549
rect 38617 18515 38651 18519
rect 38617 18451 38651 18477
rect 38617 18443 38651 18451
rect 38617 18383 38651 18405
rect 38617 18371 38651 18383
rect 38617 18315 38651 18333
rect 38617 18299 38651 18315
rect 38617 18247 38651 18261
rect 38617 18227 38651 18247
rect 38617 18179 38651 18189
rect 38617 18155 38651 18179
rect 38617 18111 38651 18117
rect 38617 18083 38651 18111
rect 38617 18043 38651 18045
rect 38617 18011 38651 18043
rect 38617 17941 38651 17973
rect 38617 17939 38651 17941
rect 38617 17873 38651 17901
rect 38617 17867 38651 17873
rect 38617 17805 38651 17829
rect 38617 17795 38651 17805
rect 38617 17737 38651 17757
rect 38617 17723 38651 17737
rect 38617 17669 38651 17685
rect 38617 17651 38651 17669
rect 38617 17601 38651 17613
rect 38617 17579 38651 17601
rect 38617 17533 38651 17541
rect 38617 17507 38651 17533
rect 38617 17465 38651 17469
rect 38617 17435 38651 17465
rect 38617 17363 38651 17397
rect 39075 18587 39109 18621
rect 39075 18519 39109 18549
rect 39075 18515 39109 18519
rect 39075 18451 39109 18477
rect 39075 18443 39109 18451
rect 39075 18383 39109 18405
rect 39075 18371 39109 18383
rect 39075 18315 39109 18333
rect 39075 18299 39109 18315
rect 39075 18247 39109 18261
rect 39075 18227 39109 18247
rect 39075 18179 39109 18189
rect 39075 18155 39109 18179
rect 39075 18111 39109 18117
rect 39075 18083 39109 18111
rect 39075 18043 39109 18045
rect 39075 18011 39109 18043
rect 39075 17941 39109 17973
rect 39075 17939 39109 17941
rect 39075 17873 39109 17901
rect 39075 17867 39109 17873
rect 39075 17805 39109 17829
rect 39075 17795 39109 17805
rect 39075 17737 39109 17757
rect 39075 17723 39109 17737
rect 39075 17669 39109 17685
rect 39075 17651 39109 17669
rect 39075 17601 39109 17613
rect 39075 17579 39109 17601
rect 39075 17533 39109 17541
rect 39075 17507 39109 17533
rect 39075 17465 39109 17469
rect 39075 17435 39109 17465
rect 39075 17363 39109 17397
rect 39533 18587 39567 18621
rect 39533 18519 39567 18549
rect 39533 18515 39567 18519
rect 39533 18451 39567 18477
rect 39533 18443 39567 18451
rect 39533 18383 39567 18405
rect 39533 18371 39567 18383
rect 39533 18315 39567 18333
rect 39533 18299 39567 18315
rect 39533 18247 39567 18261
rect 39533 18227 39567 18247
rect 39533 18179 39567 18189
rect 39533 18155 39567 18179
rect 39533 18111 39567 18117
rect 39533 18083 39567 18111
rect 39533 18043 39567 18045
rect 39533 18011 39567 18043
rect 39533 17941 39567 17973
rect 39533 17939 39567 17941
rect 39533 17873 39567 17901
rect 39533 17867 39567 17873
rect 39533 17805 39567 17829
rect 39533 17795 39567 17805
rect 39533 17737 39567 17757
rect 39533 17723 39567 17737
rect 39533 17669 39567 17685
rect 39533 17651 39567 17669
rect 39533 17601 39567 17613
rect 39533 17579 39567 17601
rect 39533 17533 39567 17541
rect 39533 17507 39567 17533
rect 39533 17465 39567 17469
rect 39533 17435 39567 17465
rect 39533 17363 39567 17397
rect 39991 18587 40025 18621
rect 39991 18519 40025 18549
rect 39991 18515 40025 18519
rect 39991 18451 40025 18477
rect 39991 18443 40025 18451
rect 39991 18383 40025 18405
rect 39991 18371 40025 18383
rect 39991 18315 40025 18333
rect 39991 18299 40025 18315
rect 39991 18247 40025 18261
rect 39991 18227 40025 18247
rect 39991 18179 40025 18189
rect 39991 18155 40025 18179
rect 39991 18111 40025 18117
rect 39991 18083 40025 18111
rect 39991 18043 40025 18045
rect 39991 18011 40025 18043
rect 39991 17941 40025 17973
rect 39991 17939 40025 17941
rect 39991 17873 40025 17901
rect 39991 17867 40025 17873
rect 39991 17805 40025 17829
rect 39991 17795 40025 17805
rect 39991 17737 40025 17757
rect 39991 17723 40025 17737
rect 39991 17669 40025 17685
rect 39991 17651 40025 17669
rect 39991 17601 40025 17613
rect 39991 17579 40025 17601
rect 39991 17533 40025 17541
rect 39991 17507 40025 17533
rect 39991 17465 40025 17469
rect 39991 17435 40025 17465
rect 39991 17363 40025 17397
rect 40449 18587 40483 18621
rect 40449 18519 40483 18549
rect 40449 18515 40483 18519
rect 40449 18451 40483 18477
rect 40449 18443 40483 18451
rect 40449 18383 40483 18405
rect 40449 18371 40483 18383
rect 40449 18315 40483 18333
rect 40449 18299 40483 18315
rect 40449 18247 40483 18261
rect 40449 18227 40483 18247
rect 40449 18179 40483 18189
rect 40449 18155 40483 18179
rect 40449 18111 40483 18117
rect 40449 18083 40483 18111
rect 40449 18043 40483 18045
rect 40449 18011 40483 18043
rect 40449 17941 40483 17973
rect 40449 17939 40483 17941
rect 40449 17873 40483 17901
rect 40449 17867 40483 17873
rect 40449 17805 40483 17829
rect 40449 17795 40483 17805
rect 40449 17737 40483 17757
rect 40449 17723 40483 17737
rect 40449 17669 40483 17685
rect 40449 17651 40483 17669
rect 40449 17601 40483 17613
rect 40449 17579 40483 17601
rect 40449 17533 40483 17541
rect 40449 17507 40483 17533
rect 40449 17465 40483 17469
rect 40449 17435 40483 17465
rect 40449 17363 40483 17397
rect 40907 18587 40941 18621
rect 40907 18519 40941 18549
rect 40907 18515 40941 18519
rect 40907 18451 40941 18477
rect 40907 18443 40941 18451
rect 40907 18383 40941 18405
rect 40907 18371 40941 18383
rect 40907 18315 40941 18333
rect 40907 18299 40941 18315
rect 40907 18247 40941 18261
rect 40907 18227 40941 18247
rect 40907 18179 40941 18189
rect 40907 18155 40941 18179
rect 40907 18111 40941 18117
rect 40907 18083 40941 18111
rect 40907 18043 40941 18045
rect 40907 18011 40941 18043
rect 40907 17941 40941 17973
rect 40907 17939 40941 17941
rect 40907 17873 40941 17901
rect 40907 17867 40941 17873
rect 40907 17805 40941 17829
rect 40907 17795 40941 17805
rect 40907 17737 40941 17757
rect 40907 17723 40941 17737
rect 40907 17669 40941 17685
rect 40907 17651 40941 17669
rect 40907 17601 40941 17613
rect 40907 17579 40941 17601
rect 40907 17533 40941 17541
rect 40907 17507 40941 17533
rect 40907 17465 40941 17469
rect 40907 17435 40941 17465
rect 40907 17363 40941 17397
rect 41365 18587 41399 18621
rect 41365 18519 41399 18549
rect 41365 18515 41399 18519
rect 41365 18451 41399 18477
rect 41365 18443 41399 18451
rect 41365 18383 41399 18405
rect 41365 18371 41399 18383
rect 41365 18315 41399 18333
rect 41365 18299 41399 18315
rect 41365 18247 41399 18261
rect 41365 18227 41399 18247
rect 41365 18179 41399 18189
rect 41365 18155 41399 18179
rect 41365 18111 41399 18117
rect 41365 18083 41399 18111
rect 41365 18043 41399 18045
rect 41365 18011 41399 18043
rect 41365 17941 41399 17973
rect 41365 17939 41399 17941
rect 41365 17873 41399 17901
rect 41365 17867 41399 17873
rect 41365 17805 41399 17829
rect 41365 17795 41399 17805
rect 41365 17737 41399 17757
rect 41365 17723 41399 17737
rect 41365 17669 41399 17685
rect 41365 17651 41399 17669
rect 41365 17601 41399 17613
rect 41365 17579 41399 17601
rect 41365 17533 41399 17541
rect 41365 17507 41399 17533
rect 41365 17465 41399 17469
rect 41365 17435 41399 17465
rect 41365 17363 41399 17397
rect 41823 18587 41857 18621
rect 41823 18519 41857 18549
rect 41823 18515 41857 18519
rect 41823 18451 41857 18477
rect 41823 18443 41857 18451
rect 41823 18383 41857 18405
rect 41823 18371 41857 18383
rect 41823 18315 41857 18333
rect 41823 18299 41857 18315
rect 41823 18247 41857 18261
rect 41823 18227 41857 18247
rect 41823 18179 41857 18189
rect 41823 18155 41857 18179
rect 41823 18111 41857 18117
rect 41823 18083 41857 18111
rect 41823 18043 41857 18045
rect 41823 18011 41857 18043
rect 41823 17941 41857 17973
rect 41823 17939 41857 17941
rect 41823 17873 41857 17901
rect 41823 17867 41857 17873
rect 41823 17805 41857 17829
rect 41823 17795 41857 17805
rect 41823 17737 41857 17757
rect 41823 17723 41857 17737
rect 41823 17669 41857 17685
rect 41823 17651 41857 17669
rect 41823 17601 41857 17613
rect 41823 17579 41857 17601
rect 41823 17533 41857 17541
rect 41823 17507 41857 17533
rect 41823 17465 41857 17469
rect 41823 17435 41857 17465
rect 41823 17363 41857 17397
rect 42281 18587 42315 18621
rect 42281 18519 42315 18549
rect 42281 18515 42315 18519
rect 42281 18451 42315 18477
rect 42281 18443 42315 18451
rect 42281 18383 42315 18405
rect 42281 18371 42315 18383
rect 42281 18315 42315 18333
rect 42281 18299 42315 18315
rect 42281 18247 42315 18261
rect 42281 18227 42315 18247
rect 42281 18179 42315 18189
rect 42281 18155 42315 18179
rect 42281 18111 42315 18117
rect 42281 18083 42315 18111
rect 42281 18043 42315 18045
rect 42281 18011 42315 18043
rect 42281 17941 42315 17973
rect 42281 17939 42315 17941
rect 42281 17873 42315 17901
rect 42281 17867 42315 17873
rect 42281 17805 42315 17829
rect 42281 17795 42315 17805
rect 42281 17737 42315 17757
rect 42281 17723 42315 17737
rect 42281 17669 42315 17685
rect 42281 17651 42315 17669
rect 42281 17601 42315 17613
rect 42281 17579 42315 17601
rect 42281 17533 42315 17541
rect 42281 17507 42315 17533
rect 42281 17465 42315 17469
rect 42281 17435 42315 17465
rect 42281 17363 42315 17397
rect 42739 18587 42773 18621
rect 42739 18519 42773 18549
rect 42739 18515 42773 18519
rect 42739 18451 42773 18477
rect 42739 18443 42773 18451
rect 42739 18383 42773 18405
rect 42739 18371 42773 18383
rect 42739 18315 42773 18333
rect 42739 18299 42773 18315
rect 42739 18247 42773 18261
rect 42739 18227 42773 18247
rect 42739 18179 42773 18189
rect 42739 18155 42773 18179
rect 42739 18111 42773 18117
rect 42739 18083 42773 18111
rect 42739 18043 42773 18045
rect 42739 18011 42773 18043
rect 42739 17941 42773 17973
rect 42739 17939 42773 17941
rect 42739 17873 42773 17901
rect 42739 17867 42773 17873
rect 42739 17805 42773 17829
rect 42739 17795 42773 17805
rect 42739 17737 42773 17757
rect 42739 17723 42773 17737
rect 42739 17669 42773 17685
rect 42739 17651 42773 17669
rect 42739 17601 42773 17613
rect 42739 17579 42773 17601
rect 42739 17533 42773 17541
rect 42739 17507 42773 17533
rect 42739 17465 42773 17469
rect 42739 17435 42773 17465
rect 42739 17363 42773 17397
rect 43197 18587 43231 18621
rect 43197 18519 43231 18549
rect 43197 18515 43231 18519
rect 43197 18451 43231 18477
rect 43197 18443 43231 18451
rect 43197 18383 43231 18405
rect 43197 18371 43231 18383
rect 43197 18315 43231 18333
rect 43197 18299 43231 18315
rect 43197 18247 43231 18261
rect 43197 18227 43231 18247
rect 43197 18179 43231 18189
rect 43197 18155 43231 18179
rect 43197 18111 43231 18117
rect 43197 18083 43231 18111
rect 43197 18043 43231 18045
rect 43197 18011 43231 18043
rect 43197 17941 43231 17973
rect 43197 17939 43231 17941
rect 43197 17873 43231 17901
rect 43197 17867 43231 17873
rect 43197 17805 43231 17829
rect 43197 17795 43231 17805
rect 43197 17737 43231 17757
rect 43197 17723 43231 17737
rect 43197 17669 43231 17685
rect 43197 17651 43231 17669
rect 43197 17601 43231 17613
rect 43197 17579 43231 17601
rect 43197 17533 43231 17541
rect 43197 17507 43231 17533
rect 43197 17465 43231 17469
rect 43197 17435 43231 17465
rect 43197 17363 43231 17397
rect 43655 18587 43689 18621
rect 43655 18519 43689 18549
rect 43655 18515 43689 18519
rect 43655 18451 43689 18477
rect 43655 18443 43689 18451
rect 43655 18383 43689 18405
rect 43655 18371 43689 18383
rect 43655 18315 43689 18333
rect 43655 18299 43689 18315
rect 43655 18247 43689 18261
rect 43655 18227 43689 18247
rect 43655 18179 43689 18189
rect 43655 18155 43689 18179
rect 43655 18111 43689 18117
rect 43655 18083 43689 18111
rect 43655 18043 43689 18045
rect 43655 18011 43689 18043
rect 43655 17941 43689 17973
rect 43655 17939 43689 17941
rect 43655 17873 43689 17901
rect 43655 17867 43689 17873
rect 43655 17805 43689 17829
rect 43655 17795 43689 17805
rect 43655 17737 43689 17757
rect 43655 17723 43689 17737
rect 43655 17669 43689 17685
rect 43655 17651 43689 17669
rect 43655 17601 43689 17613
rect 43655 17579 43689 17601
rect 43655 17533 43689 17541
rect 43655 17507 43689 17533
rect 43655 17465 43689 17469
rect 43655 17435 43689 17465
rect 43655 17363 43689 17397
rect 44113 18587 44147 18621
rect 44113 18519 44147 18549
rect 44113 18515 44147 18519
rect 44113 18451 44147 18477
rect 44113 18443 44147 18451
rect 44113 18383 44147 18405
rect 44113 18371 44147 18383
rect 44113 18315 44147 18333
rect 44113 18299 44147 18315
rect 44113 18247 44147 18261
rect 44113 18227 44147 18247
rect 44113 18179 44147 18189
rect 44113 18155 44147 18179
rect 44113 18111 44147 18117
rect 44113 18083 44147 18111
rect 44113 18043 44147 18045
rect 44113 18011 44147 18043
rect 44113 17941 44147 17973
rect 44113 17939 44147 17941
rect 44113 17873 44147 17901
rect 44113 17867 44147 17873
rect 44113 17805 44147 17829
rect 44113 17795 44147 17805
rect 44113 17737 44147 17757
rect 44113 17723 44147 17737
rect 44113 17669 44147 17685
rect 44113 17651 44147 17669
rect 44113 17601 44147 17613
rect 44113 17579 44147 17601
rect 44113 17533 44147 17541
rect 44113 17507 44147 17533
rect 44113 17465 44147 17469
rect 44113 17435 44147 17465
rect 44113 17363 44147 17397
rect 44571 18587 44605 18621
rect 44571 18519 44605 18549
rect 44571 18515 44605 18519
rect 44571 18451 44605 18477
rect 44571 18443 44605 18451
rect 44571 18383 44605 18405
rect 44571 18371 44605 18383
rect 44571 18315 44605 18333
rect 44571 18299 44605 18315
rect 44571 18247 44605 18261
rect 44571 18227 44605 18247
rect 44571 18179 44605 18189
rect 44571 18155 44605 18179
rect 44571 18111 44605 18117
rect 44571 18083 44605 18111
rect 44571 18043 44605 18045
rect 44571 18011 44605 18043
rect 44571 17941 44605 17973
rect 44571 17939 44605 17941
rect 44571 17873 44605 17901
rect 44571 17867 44605 17873
rect 44571 17805 44605 17829
rect 44571 17795 44605 17805
rect 44571 17737 44605 17757
rect 44571 17723 44605 17737
rect 44571 17669 44605 17685
rect 44571 17651 44605 17669
rect 44571 17601 44605 17613
rect 44571 17579 44605 17601
rect 44571 17533 44605 17541
rect 44571 17507 44605 17533
rect 44571 17465 44605 17469
rect 44571 17435 44605 17465
rect 44571 17363 44605 17397
rect 45029 18587 45063 18621
rect 45029 18519 45063 18549
rect 45029 18515 45063 18519
rect 45029 18451 45063 18477
rect 45029 18443 45063 18451
rect 45029 18383 45063 18405
rect 45029 18371 45063 18383
rect 45029 18315 45063 18333
rect 45029 18299 45063 18315
rect 45029 18247 45063 18261
rect 45029 18227 45063 18247
rect 45029 18179 45063 18189
rect 45029 18155 45063 18179
rect 45029 18111 45063 18117
rect 45029 18083 45063 18111
rect 45029 18043 45063 18045
rect 45029 18011 45063 18043
rect 45029 17941 45063 17973
rect 45029 17939 45063 17941
rect 45029 17873 45063 17901
rect 45029 17867 45063 17873
rect 45029 17805 45063 17829
rect 45029 17795 45063 17805
rect 45029 17737 45063 17757
rect 45029 17723 45063 17737
rect 45029 17669 45063 17685
rect 45029 17651 45063 17669
rect 45029 17601 45063 17613
rect 45029 17579 45063 17601
rect 45029 17533 45063 17541
rect 45029 17507 45063 17533
rect 45029 17465 45063 17469
rect 45029 17435 45063 17465
rect 45029 17363 45063 17397
rect 45487 18587 45521 18621
rect 45487 18519 45521 18549
rect 45487 18515 45521 18519
rect 45487 18451 45521 18477
rect 45487 18443 45521 18451
rect 45487 18383 45521 18405
rect 45487 18371 45521 18383
rect 45487 18315 45521 18333
rect 45487 18299 45521 18315
rect 45487 18247 45521 18261
rect 45487 18227 45521 18247
rect 45487 18179 45521 18189
rect 45487 18155 45521 18179
rect 45487 18111 45521 18117
rect 45487 18083 45521 18111
rect 45487 18043 45521 18045
rect 45487 18011 45521 18043
rect 45487 17941 45521 17973
rect 45487 17939 45521 17941
rect 45487 17873 45521 17901
rect 45487 17867 45521 17873
rect 45487 17805 45521 17829
rect 45487 17795 45521 17805
rect 45487 17737 45521 17757
rect 45487 17723 45521 17737
rect 45487 17669 45521 17685
rect 45487 17651 45521 17669
rect 45487 17601 45521 17613
rect 45487 17579 45521 17601
rect 45487 17533 45521 17541
rect 45487 17507 45521 17533
rect 45487 17465 45521 17469
rect 45487 17435 45521 17465
rect 45487 17363 45521 17397
rect 45945 18587 45979 18621
rect 45945 18519 45979 18549
rect 45945 18515 45979 18519
rect 45945 18451 45979 18477
rect 45945 18443 45979 18451
rect 45945 18383 45979 18405
rect 45945 18371 45979 18383
rect 45945 18315 45979 18333
rect 45945 18299 45979 18315
rect 45945 18247 45979 18261
rect 45945 18227 45979 18247
rect 45945 18179 45979 18189
rect 45945 18155 45979 18179
rect 45945 18111 45979 18117
rect 45945 18083 45979 18111
rect 45945 18043 45979 18045
rect 45945 18011 45979 18043
rect 45945 17941 45979 17973
rect 45945 17939 45979 17941
rect 45945 17873 45979 17901
rect 45945 17867 45979 17873
rect 45945 17805 45979 17829
rect 45945 17795 45979 17805
rect 45945 17737 45979 17757
rect 45945 17723 45979 17737
rect 45945 17669 45979 17685
rect 45945 17651 45979 17669
rect 45945 17601 45979 17613
rect 45945 17579 45979 17601
rect 45945 17533 45979 17541
rect 45945 17507 45979 17533
rect 45945 17465 45979 17469
rect 45945 17435 45979 17465
rect 45945 17363 45979 17397
rect 46403 18587 46437 18621
rect 46403 18519 46437 18549
rect 46403 18515 46437 18519
rect 46403 18451 46437 18477
rect 46403 18443 46437 18451
rect 46403 18383 46437 18405
rect 46403 18371 46437 18383
rect 46403 18315 46437 18333
rect 46403 18299 46437 18315
rect 46403 18247 46437 18261
rect 46403 18227 46437 18247
rect 46403 18179 46437 18189
rect 46403 18155 46437 18179
rect 46403 18111 46437 18117
rect 46403 18083 46437 18111
rect 46403 18043 46437 18045
rect 46403 18011 46437 18043
rect 46403 17941 46437 17973
rect 46403 17939 46437 17941
rect 46403 17873 46437 17901
rect 46403 17867 46437 17873
rect 46403 17805 46437 17829
rect 46403 17795 46437 17805
rect 46403 17737 46437 17757
rect 46403 17723 46437 17737
rect 46403 17669 46437 17685
rect 46403 17651 46437 17669
rect 46403 17601 46437 17613
rect 46403 17579 46437 17601
rect 46403 17533 46437 17541
rect 46403 17507 46437 17533
rect 46403 17465 46437 17469
rect 46403 17435 46437 17465
rect 46403 17363 46437 17397
rect 46861 18587 46895 18621
rect 46861 18519 46895 18549
rect 46861 18515 46895 18519
rect 46861 18451 46895 18477
rect 46861 18443 46895 18451
rect 46861 18383 46895 18405
rect 46861 18371 46895 18383
rect 46861 18315 46895 18333
rect 46861 18299 46895 18315
rect 46861 18247 46895 18261
rect 46861 18227 46895 18247
rect 46861 18179 46895 18189
rect 46861 18155 46895 18179
rect 46861 18111 46895 18117
rect 46861 18083 46895 18111
rect 46861 18043 46895 18045
rect 46861 18011 46895 18043
rect 46861 17941 46895 17973
rect 46861 17939 46895 17941
rect 46861 17873 46895 17901
rect 46861 17867 46895 17873
rect 46861 17805 46895 17829
rect 46861 17795 46895 17805
rect 46861 17737 46895 17757
rect 46861 17723 46895 17737
rect 46861 17669 46895 17685
rect 46861 17651 46895 17669
rect 46861 17601 46895 17613
rect 46861 17579 46895 17601
rect 46861 17533 46895 17541
rect 46861 17507 46895 17533
rect 46861 17465 46895 17469
rect 46861 17435 46895 17465
rect 46861 17363 46895 17397
rect 47319 18587 47353 18621
rect 47319 18519 47353 18549
rect 47319 18515 47353 18519
rect 47319 18451 47353 18477
rect 47319 18443 47353 18451
rect 47319 18383 47353 18405
rect 47319 18371 47353 18383
rect 47319 18315 47353 18333
rect 47319 18299 47353 18315
rect 47319 18247 47353 18261
rect 47319 18227 47353 18247
rect 47319 18179 47353 18189
rect 47319 18155 47353 18179
rect 47319 18111 47353 18117
rect 47319 18083 47353 18111
rect 47319 18043 47353 18045
rect 47319 18011 47353 18043
rect 47319 17941 47353 17973
rect 47319 17939 47353 17941
rect 47319 17873 47353 17901
rect 47319 17867 47353 17873
rect 47319 17805 47353 17829
rect 47319 17795 47353 17805
rect 47319 17737 47353 17757
rect 47319 17723 47353 17737
rect 47319 17669 47353 17685
rect 47319 17651 47353 17669
rect 47319 17601 47353 17613
rect 47319 17579 47353 17601
rect 47319 17533 47353 17541
rect 47319 17507 47353 17533
rect 47319 17465 47353 17469
rect 47319 17435 47353 17465
rect 47319 17363 47353 17397
rect 47777 18587 47811 18621
rect 47777 18519 47811 18549
rect 47777 18515 47811 18519
rect 47777 18451 47811 18477
rect 47777 18443 47811 18451
rect 47777 18383 47811 18405
rect 47777 18371 47811 18383
rect 47777 18315 47811 18333
rect 47777 18299 47811 18315
rect 47777 18247 47811 18261
rect 47777 18227 47811 18247
rect 47777 18179 47811 18189
rect 47777 18155 47811 18179
rect 47777 18111 47811 18117
rect 47777 18083 47811 18111
rect 47777 18043 47811 18045
rect 47777 18011 47811 18043
rect 47777 17941 47811 17973
rect 47777 17939 47811 17941
rect 47777 17873 47811 17901
rect 47777 17867 47811 17873
rect 47777 17805 47811 17829
rect 47777 17795 47811 17805
rect 47777 17737 47811 17757
rect 47777 17723 47811 17737
rect 47777 17669 47811 17685
rect 47777 17651 47811 17669
rect 47777 17601 47811 17613
rect 47777 17579 47811 17601
rect 47777 17533 47811 17541
rect 47777 17507 47811 17533
rect 47777 17465 47811 17469
rect 47777 17435 47811 17465
rect 47777 17363 47811 17397
rect 48235 18587 48269 18621
rect 48235 18519 48269 18549
rect 48235 18515 48269 18519
rect 48235 18451 48269 18477
rect 48235 18443 48269 18451
rect 48235 18383 48269 18405
rect 48235 18371 48269 18383
rect 48235 18315 48269 18333
rect 48235 18299 48269 18315
rect 48235 18247 48269 18261
rect 48235 18227 48269 18247
rect 48235 18179 48269 18189
rect 48235 18155 48269 18179
rect 48235 18111 48269 18117
rect 48235 18083 48269 18111
rect 48235 18043 48269 18045
rect 48235 18011 48269 18043
rect 48235 17941 48269 17973
rect 48235 17939 48269 17941
rect 48235 17873 48269 17901
rect 48235 17867 48269 17873
rect 48235 17805 48269 17829
rect 48235 17795 48269 17805
rect 48235 17737 48269 17757
rect 48235 17723 48269 17737
rect 48235 17669 48269 17685
rect 48235 17651 48269 17669
rect 48235 17601 48269 17613
rect 48235 17579 48269 17601
rect 48235 17533 48269 17541
rect 48235 17507 48269 17533
rect 48235 17465 48269 17469
rect 48235 17435 48269 17465
rect 48235 17363 48269 17397
rect 48693 18587 48727 18621
rect 48693 18519 48727 18549
rect 48693 18515 48727 18519
rect 48693 18451 48727 18477
rect 48693 18443 48727 18451
rect 48693 18383 48727 18405
rect 48693 18371 48727 18383
rect 48693 18315 48727 18333
rect 48693 18299 48727 18315
rect 48693 18247 48727 18261
rect 48693 18227 48727 18247
rect 48693 18179 48727 18189
rect 48693 18155 48727 18179
rect 48693 18111 48727 18117
rect 48693 18083 48727 18111
rect 48693 18043 48727 18045
rect 48693 18011 48727 18043
rect 48693 17941 48727 17973
rect 48693 17939 48727 17941
rect 48693 17873 48727 17901
rect 48693 17867 48727 17873
rect 48693 17805 48727 17829
rect 48693 17795 48727 17805
rect 48693 17737 48727 17757
rect 48693 17723 48727 17737
rect 48693 17669 48727 17685
rect 48693 17651 48727 17669
rect 48693 17601 48727 17613
rect 48693 17579 48727 17601
rect 48693 17533 48727 17541
rect 48693 17507 48727 17533
rect 48693 17465 48727 17469
rect 48693 17435 48727 17465
rect 48693 17363 48727 17397
rect 49151 18587 49185 18621
rect 49151 18519 49185 18549
rect 49151 18515 49185 18519
rect 49151 18451 49185 18477
rect 49151 18443 49185 18451
rect 49151 18383 49185 18405
rect 49151 18371 49185 18383
rect 49151 18315 49185 18333
rect 49151 18299 49185 18315
rect 49151 18247 49185 18261
rect 49151 18227 49185 18247
rect 49151 18179 49185 18189
rect 49151 18155 49185 18179
rect 49151 18111 49185 18117
rect 49151 18083 49185 18111
rect 49151 18043 49185 18045
rect 49151 18011 49185 18043
rect 49151 17941 49185 17973
rect 49151 17939 49185 17941
rect 49151 17873 49185 17901
rect 49151 17867 49185 17873
rect 49151 17805 49185 17829
rect 49151 17795 49185 17805
rect 49151 17737 49185 17757
rect 49151 17723 49185 17737
rect 49151 17669 49185 17685
rect 49151 17651 49185 17669
rect 49151 17601 49185 17613
rect 49151 17579 49185 17601
rect 49151 17533 49185 17541
rect 49151 17507 49185 17533
rect 49151 17465 49185 17469
rect 49151 17435 49185 17465
rect 49151 17363 49185 17397
rect 49609 18587 49643 18621
rect 49609 18519 49643 18549
rect 49609 18515 49643 18519
rect 49609 18451 49643 18477
rect 49609 18443 49643 18451
rect 49609 18383 49643 18405
rect 49609 18371 49643 18383
rect 49609 18315 49643 18333
rect 49609 18299 49643 18315
rect 49609 18247 49643 18261
rect 49609 18227 49643 18247
rect 49609 18179 49643 18189
rect 49609 18155 49643 18179
rect 49609 18111 49643 18117
rect 49609 18083 49643 18111
rect 49609 18043 49643 18045
rect 49609 18011 49643 18043
rect 49609 17941 49643 17973
rect 49609 17939 49643 17941
rect 49609 17873 49643 17901
rect 49609 17867 49643 17873
rect 49609 17805 49643 17829
rect 49609 17795 49643 17805
rect 49609 17737 49643 17757
rect 49609 17723 49643 17737
rect 49609 17669 49643 17685
rect 49609 17651 49643 17669
rect 49609 17601 49643 17613
rect 49609 17579 49643 17601
rect 49609 17533 49643 17541
rect 49609 17507 49643 17533
rect 49609 17465 49643 17469
rect 49609 17435 49643 17465
rect 49609 17363 49643 17397
rect 50067 18587 50101 18621
rect 50067 18519 50101 18549
rect 50067 18515 50101 18519
rect 50067 18451 50101 18477
rect 50067 18443 50101 18451
rect 50067 18383 50101 18405
rect 50067 18371 50101 18383
rect 50067 18315 50101 18333
rect 50067 18299 50101 18315
rect 50067 18247 50101 18261
rect 50067 18227 50101 18247
rect 50067 18179 50101 18189
rect 50067 18155 50101 18179
rect 50067 18111 50101 18117
rect 50067 18083 50101 18111
rect 50067 18043 50101 18045
rect 50067 18011 50101 18043
rect 50067 17941 50101 17973
rect 50067 17939 50101 17941
rect 50067 17873 50101 17901
rect 50067 17867 50101 17873
rect 50067 17805 50101 17829
rect 50067 17795 50101 17805
rect 50067 17737 50101 17757
rect 50067 17723 50101 17737
rect 50067 17669 50101 17685
rect 50067 17651 50101 17669
rect 50067 17601 50101 17613
rect 50067 17579 50101 17601
rect 50067 17533 50101 17541
rect 50067 17507 50101 17533
rect 50067 17465 50101 17469
rect 50067 17435 50101 17465
rect 50067 17363 50101 17397
rect 50525 18587 50559 18621
rect 50525 18519 50559 18549
rect 50525 18515 50559 18519
rect 50525 18451 50559 18477
rect 50525 18443 50559 18451
rect 50525 18383 50559 18405
rect 50525 18371 50559 18383
rect 50525 18315 50559 18333
rect 50525 18299 50559 18315
rect 50525 18247 50559 18261
rect 50525 18227 50559 18247
rect 50525 18179 50559 18189
rect 50525 18155 50559 18179
rect 50525 18111 50559 18117
rect 50525 18083 50559 18111
rect 50525 18043 50559 18045
rect 50525 18011 50559 18043
rect 50525 17941 50559 17973
rect 50525 17939 50559 17941
rect 50525 17873 50559 17901
rect 50525 17867 50559 17873
rect 50525 17805 50559 17829
rect 50525 17795 50559 17805
rect 50525 17737 50559 17757
rect 50525 17723 50559 17737
rect 50525 17669 50559 17685
rect 50525 17651 50559 17669
rect 50525 17601 50559 17613
rect 50525 17579 50559 17601
rect 50525 17533 50559 17541
rect 50525 17507 50559 17533
rect 50525 17465 50559 17469
rect 50525 17435 50559 17465
rect 50525 17363 50559 17397
rect 50983 18587 51017 18621
rect 50983 18519 51017 18549
rect 50983 18515 51017 18519
rect 50983 18451 51017 18477
rect 50983 18443 51017 18451
rect 50983 18383 51017 18405
rect 50983 18371 51017 18383
rect 50983 18315 51017 18333
rect 50983 18299 51017 18315
rect 50983 18247 51017 18261
rect 50983 18227 51017 18247
rect 50983 18179 51017 18189
rect 50983 18155 51017 18179
rect 50983 18111 51017 18117
rect 50983 18083 51017 18111
rect 50983 18043 51017 18045
rect 50983 18011 51017 18043
rect 50983 17941 51017 17973
rect 50983 17939 51017 17941
rect 50983 17873 51017 17901
rect 50983 17867 51017 17873
rect 50983 17805 51017 17829
rect 50983 17795 51017 17805
rect 50983 17737 51017 17757
rect 50983 17723 51017 17737
rect 50983 17669 51017 17685
rect 50983 17651 51017 17669
rect 50983 17601 51017 17613
rect 50983 17579 51017 17601
rect 50983 17533 51017 17541
rect 50983 17507 51017 17533
rect 50983 17465 51017 17469
rect 50983 17435 51017 17465
rect 50983 17363 51017 17397
rect 51441 18587 51475 18621
rect 51441 18519 51475 18549
rect 51441 18515 51475 18519
rect 51441 18451 51475 18477
rect 51441 18443 51475 18451
rect 51441 18383 51475 18405
rect 51441 18371 51475 18383
rect 51441 18315 51475 18333
rect 51441 18299 51475 18315
rect 51441 18247 51475 18261
rect 51441 18227 51475 18247
rect 51441 18179 51475 18189
rect 51441 18155 51475 18179
rect 51441 18111 51475 18117
rect 51441 18083 51475 18111
rect 51441 18043 51475 18045
rect 51441 18011 51475 18043
rect 51441 17941 51475 17973
rect 51441 17939 51475 17941
rect 51441 17873 51475 17901
rect 51441 17867 51475 17873
rect 51441 17805 51475 17829
rect 51441 17795 51475 17805
rect 51441 17737 51475 17757
rect 51441 17723 51475 17737
rect 51441 17669 51475 17685
rect 51441 17651 51475 17669
rect 51441 17601 51475 17613
rect 51441 17579 51475 17601
rect 51441 17533 51475 17541
rect 51441 17507 51475 17533
rect 51441 17465 51475 17469
rect 51441 17435 51475 17465
rect 51441 17363 51475 17397
rect 51899 18587 51933 18621
rect 51899 18519 51933 18549
rect 51899 18515 51933 18519
rect 51899 18451 51933 18477
rect 51899 18443 51933 18451
rect 51899 18383 51933 18405
rect 51899 18371 51933 18383
rect 51899 18315 51933 18333
rect 51899 18299 51933 18315
rect 51899 18247 51933 18261
rect 51899 18227 51933 18247
rect 51899 18179 51933 18189
rect 51899 18155 51933 18179
rect 51899 18111 51933 18117
rect 51899 18083 51933 18111
rect 51899 18043 51933 18045
rect 51899 18011 51933 18043
rect 51899 17941 51933 17973
rect 51899 17939 51933 17941
rect 51899 17873 51933 17901
rect 51899 17867 51933 17873
rect 51899 17805 51933 17829
rect 51899 17795 51933 17805
rect 51899 17737 51933 17757
rect 51899 17723 51933 17737
rect 51899 17669 51933 17685
rect 51899 17651 51933 17669
rect 51899 17601 51933 17613
rect 51899 17579 51933 17601
rect 51899 17533 51933 17541
rect 51899 17507 51933 17533
rect 51899 17465 51933 17469
rect 51899 17435 51933 17465
rect 51899 17363 51933 17397
rect 52357 18587 52391 18621
rect 52357 18519 52391 18549
rect 52357 18515 52391 18519
rect 52357 18451 52391 18477
rect 52357 18443 52391 18451
rect 52357 18383 52391 18405
rect 52357 18371 52391 18383
rect 52357 18315 52391 18333
rect 52357 18299 52391 18315
rect 52357 18247 52391 18261
rect 52357 18227 52391 18247
rect 52357 18179 52391 18189
rect 52357 18155 52391 18179
rect 52357 18111 52391 18117
rect 52357 18083 52391 18111
rect 52357 18043 52391 18045
rect 52357 18011 52391 18043
rect 52357 17941 52391 17973
rect 52357 17939 52391 17941
rect 52357 17873 52391 17901
rect 52357 17867 52391 17873
rect 52357 17805 52391 17829
rect 52357 17795 52391 17805
rect 52357 17737 52391 17757
rect 52357 17723 52391 17737
rect 52357 17669 52391 17685
rect 52357 17651 52391 17669
rect 52357 17601 52391 17613
rect 52357 17579 52391 17601
rect 52357 17533 52391 17541
rect 52357 17507 52391 17533
rect 52357 17465 52391 17469
rect 52357 17435 52391 17465
rect 52357 17363 52391 17397
rect 34345 17221 34379 17255
rect 25421 17143 25455 17153
rect 25421 17119 25447 17143
rect 25447 17119 25455 17143
rect 25013 16975 25047 17009
rect 25413 16975 25447 17009
rect 25813 16975 25847 17009
rect 26213 16975 26247 17009
rect 26613 16975 26647 17009
rect 27013 16975 27047 17009
rect 27413 16975 27447 17009
rect 27813 16975 27847 17009
rect 28213 16975 28247 17009
rect 28613 16975 28647 17009
rect 29013 16975 29047 17009
rect 29413 16975 29447 17009
rect 29813 16975 29847 17009
rect 30213 16975 30247 17009
rect 30613 16975 30647 17009
rect 31013 16975 31047 17009
rect 31413 16975 31447 17009
rect 31813 16975 31847 17009
rect 32213 16975 32247 17009
rect 32613 16975 32647 17009
rect 33013 16975 33047 17009
rect 33413 16975 33447 17009
rect 33813 16975 33847 17009
rect 34213 16975 34247 17009
rect 34613 16975 34647 17009
rect 35013 16975 35047 17009
rect 35413 16975 35447 17009
rect 35813 16975 35847 17009
rect 36213 16975 36247 17009
rect 36613 16975 36647 17009
rect 37013 16975 37047 17009
rect 37413 16975 37447 17009
rect 37813 16975 37847 17009
rect 38213 16975 38247 17009
rect 38613 16975 38647 17009
rect 39013 16975 39047 17009
rect 39413 16975 39447 17009
rect 39813 16975 39847 17009
rect 40213 16975 40247 17009
rect 40613 16975 40647 17009
rect 41013 16975 41047 17009
rect 41413 16975 41447 17009
rect 41813 16975 41847 17009
rect 42213 16975 42247 17009
rect 42613 16975 42647 17009
rect 43013 16975 43047 17009
rect 43413 16975 43447 17009
rect 43813 16975 43847 17009
rect 44213 16975 44247 17009
rect 44613 16975 44647 17009
rect 45013 16975 45047 17009
rect 45413 16975 45447 17009
rect 45813 16975 45847 17009
rect 46213 16975 46247 17009
rect 46613 16975 46647 17009
rect 47013 16975 47047 17009
rect 47413 16975 47447 17009
rect 47813 16975 47847 17009
rect 48213 16975 48247 17009
rect 48613 16975 48647 17009
rect 49013 16975 49047 17009
rect 49413 16975 49447 17009
rect 49813 16975 49847 17009
rect 50213 16975 50247 17009
rect 50613 16975 50647 17009
rect 51013 16975 51047 17009
rect 51413 16975 51447 17009
rect 51813 16975 51847 17009
rect 52213 16975 52247 17009
rect 44045 15095 44079 15129
rect 44245 15095 44279 15129
rect 44445 15095 44479 15129
rect 44645 15095 44679 15129
rect 44845 15095 44879 15129
rect 45045 15095 45079 15129
rect 45245 15095 45279 15129
rect 45445 15095 45479 15129
rect 45645 15095 45679 15129
rect 45845 15095 45879 15129
rect 46045 15095 46079 15129
rect 46789 15095 46823 15129
rect 46989 15095 47023 15129
rect 47189 15095 47223 15129
rect 47389 15095 47423 15129
rect 47589 15095 47623 15129
rect 47789 15095 47823 15129
rect 47989 15095 48023 15129
rect 48189 15095 48223 15129
rect 48389 15095 48423 15129
rect 48589 15095 48623 15129
rect 48789 15095 48823 15129
rect 49533 15095 49567 15129
rect 49733 15095 49767 15129
rect 49933 15095 49967 15129
rect 50133 15095 50167 15129
rect 50333 15095 50367 15129
rect 50533 15095 50567 15129
rect 50733 15095 50767 15129
rect 50933 15095 50967 15129
rect 51133 15095 51167 15129
rect 51333 15095 51367 15129
rect 51533 15095 51567 15129
rect 43881 14323 44275 14861
rect 45888 14323 46282 14861
rect 46625 14323 47019 14861
rect 48632 14323 49026 14861
rect 49369 14323 49763 14861
rect 51376 14323 51770 14861
rect 43881 13363 44275 13901
rect 45888 13363 46282 13901
rect 46625 13363 47019 13901
rect 48632 13363 49026 13901
rect 49369 13363 49763 13901
rect 51376 13363 51770 13901
rect 44045 13215 44079 13249
rect 44245 13215 44279 13249
rect 44445 13215 44479 13249
rect 44645 13215 44679 13249
rect 44845 13215 44879 13249
rect 45045 13215 45079 13249
rect 45245 13215 45279 13249
rect 45445 13215 45479 13249
rect 45645 13215 45679 13249
rect 45845 13215 45879 13249
rect 46045 13215 46079 13249
rect 46789 13215 46823 13249
rect 46989 13215 47023 13249
rect 47189 13215 47223 13249
rect 47389 13215 47423 13249
rect 47589 13215 47623 13249
rect 47789 13215 47823 13249
rect 47989 13215 48023 13249
rect 48189 13215 48223 13249
rect 48389 13215 48423 13249
rect 48589 13215 48623 13249
rect 48789 13215 48823 13249
rect 49533 13215 49567 13249
rect 49733 13215 49767 13249
rect 49933 13215 49967 13249
rect 50133 13215 50167 13249
rect 50333 13215 50367 13249
rect 50533 13215 50567 13249
rect 50733 13215 50767 13249
rect 50933 13215 50967 13249
rect 51133 13215 51167 13249
rect 51333 13215 51367 13249
rect 51533 13215 51567 13249
rect 43947 11335 43981 11369
rect 44147 11335 44181 11369
rect 44347 11335 44381 11369
rect 44547 11335 44581 11369
rect 44747 11335 44781 11369
rect 44947 11335 44981 11369
rect 45147 11335 45181 11369
rect 45347 11335 45381 11369
rect 45547 11335 45581 11369
rect 45747 11335 45781 11369
rect 45947 11335 45981 11369
rect 46691 11335 46725 11369
rect 46891 11335 46925 11369
rect 47091 11335 47125 11369
rect 47291 11335 47325 11369
rect 47491 11335 47525 11369
rect 47691 11335 47725 11369
rect 47891 11335 47925 11369
rect 48091 11335 48125 11369
rect 48291 11335 48325 11369
rect 48491 11335 48525 11369
rect 48691 11335 48725 11369
rect 49435 11335 49469 11369
rect 49635 11335 49669 11369
rect 49835 11335 49869 11369
rect 50035 11335 50069 11369
rect 50235 11335 50269 11369
rect 50435 11335 50469 11369
rect 50635 11335 50669 11369
rect 50835 11335 50869 11369
rect 51035 11335 51069 11369
rect 51235 11335 51269 11369
rect 51435 11335 51469 11369
rect 43783 10563 44177 11101
rect 45790 10563 46184 11101
rect 46527 10563 46921 11101
rect 48534 10563 48928 11101
rect 49271 10563 49665 11101
rect 51278 10563 51672 11101
rect 43783 9603 44177 10141
rect 45790 9603 46184 10141
rect 46527 9603 46921 10141
rect 48534 9603 48928 10141
rect 49271 9603 49665 10141
rect 51278 9603 51672 10141
rect 43947 9455 43981 9489
rect 44147 9455 44181 9489
rect 44347 9455 44381 9489
rect 44547 9455 44581 9489
rect 44747 9455 44781 9489
rect 44947 9455 44981 9489
rect 45147 9455 45181 9489
rect 45347 9455 45381 9489
rect 45547 9455 45581 9489
rect 45747 9455 45781 9489
rect 45947 9455 45981 9489
rect 46691 9455 46725 9489
rect 46891 9455 46925 9489
rect 47091 9455 47125 9489
rect 47291 9455 47325 9489
rect 47491 9455 47525 9489
rect 47691 9455 47725 9489
rect 47891 9455 47925 9489
rect 48091 9455 48125 9489
rect 48291 9455 48325 9489
rect 48491 9455 48525 9489
rect 48691 9455 48725 9489
rect 49435 9455 49469 9489
rect 49635 9455 49669 9489
rect 49835 9455 49869 9489
rect 50035 9455 50069 9489
rect 50235 9455 50269 9489
rect 50435 9455 50469 9489
rect 50635 9455 50669 9489
rect 50835 9455 50869 9489
rect 51035 9455 51069 9489
rect 51235 9455 51269 9489
rect 51435 9455 51469 9489
rect 44731 7575 44765 7609
rect 44931 7575 44965 7609
rect 45131 7575 45165 7609
rect 45331 7575 45365 7609
rect 45531 7575 45565 7609
rect 45731 7575 45765 7609
rect 45931 7575 45965 7609
rect 46131 7575 46165 7609
rect 46331 7575 46365 7609
rect 46531 7575 46565 7609
rect 46731 7575 46765 7609
rect 47475 7575 47509 7609
rect 47675 7575 47709 7609
rect 47875 7575 47909 7609
rect 48075 7575 48109 7609
rect 48275 7575 48309 7609
rect 48475 7575 48509 7609
rect 48675 7575 48709 7609
rect 48875 7575 48909 7609
rect 49075 7575 49109 7609
rect 49275 7575 49309 7609
rect 49475 7575 49509 7609
rect 50219 7575 50253 7609
rect 50419 7575 50453 7609
rect 50619 7575 50653 7609
rect 50819 7575 50853 7609
rect 51019 7575 51053 7609
rect 51219 7575 51253 7609
rect 51419 7575 51453 7609
rect 51619 7575 51653 7609
rect 51819 7575 51853 7609
rect 52019 7575 52053 7609
rect 52219 7575 52253 7609
rect 44567 6803 44961 7341
rect 46574 6803 46968 7341
rect 47311 6803 47705 7341
rect 49318 6803 49712 7341
rect 50055 6803 50449 7341
rect 52062 6803 52456 7341
rect 44567 5843 44961 6381
rect 46574 5843 46968 6381
rect 47311 5843 47705 6381
rect 49318 5843 49712 6381
rect 50055 5843 50449 6381
rect 52062 5843 52456 6381
rect 44731 5695 44765 5729
rect 44931 5695 44965 5729
rect 45131 5695 45165 5729
rect 45331 5695 45365 5729
rect 45531 5695 45565 5729
rect 45731 5695 45765 5729
rect 45931 5695 45965 5729
rect 46131 5695 46165 5729
rect 46331 5695 46365 5729
rect 46531 5695 46565 5729
rect 46731 5695 46765 5729
rect 47475 5695 47509 5729
rect 47675 5695 47709 5729
rect 47875 5695 47909 5729
rect 48075 5695 48109 5729
rect 48275 5695 48309 5729
rect 48475 5695 48509 5729
rect 48675 5695 48709 5729
rect 48875 5695 48909 5729
rect 49075 5695 49109 5729
rect 49275 5695 49309 5729
rect 49475 5695 49509 5729
rect 50219 5695 50253 5729
rect 50419 5695 50453 5729
rect 50619 5695 50653 5729
rect 50819 5695 50853 5729
rect 51019 5695 51053 5729
rect 51219 5695 51253 5729
rect 51419 5695 51453 5729
rect 51619 5695 51653 5729
rect 51819 5695 51853 5729
rect 52019 5695 52053 5729
rect 52219 5695 52253 5729
<< metal1 >>
rect 900 50890 57536 50892
rect 900 50774 922 50890
rect 2510 50774 55926 50890
rect 57514 50774 57536 50890
rect 900 50772 57536 50774
rect 3348 49010 55088 49012
rect 3348 48894 3370 49010
rect 4958 48969 53478 49010
rect 4958 48935 6101 48969
rect 6135 48935 6501 48969
rect 6535 48935 6901 48969
rect 6935 48935 7301 48969
rect 7335 48935 7701 48969
rect 7735 48935 8101 48969
rect 8135 48935 8501 48969
rect 8535 48935 8901 48969
rect 8935 48935 9301 48969
rect 9335 48935 9701 48969
rect 9735 48935 10101 48969
rect 10135 48935 10501 48969
rect 10535 48935 10901 48969
rect 10935 48935 11301 48969
rect 11335 48935 11701 48969
rect 11735 48935 12101 48969
rect 12135 48935 12501 48969
rect 12535 48935 12901 48969
rect 12935 48935 13549 48969
rect 13583 48935 13949 48969
rect 13983 48935 14349 48969
rect 14383 48935 14749 48969
rect 14783 48935 15149 48969
rect 15183 48935 15549 48969
rect 15583 48935 15949 48969
rect 15983 48935 16349 48969
rect 16383 48935 16749 48969
rect 16783 48935 17149 48969
rect 17183 48935 17549 48969
rect 17583 48935 17949 48969
rect 17983 48935 18349 48969
rect 18383 48935 18749 48969
rect 18783 48935 19149 48969
rect 19183 48935 19549 48969
rect 19583 48935 19949 48969
rect 19983 48935 20349 48969
rect 20383 48935 21015 48969
rect 21049 48935 21215 48969
rect 21249 48935 21415 48969
rect 21449 48935 21615 48969
rect 21649 48935 21815 48969
rect 21849 48935 22015 48969
rect 22049 48935 22215 48969
rect 22249 48935 22415 48969
rect 22449 48935 22615 48969
rect 22649 48935 22815 48969
rect 22849 48935 23015 48969
rect 23049 48935 24101 48969
rect 24135 48935 25013 48969
rect 25047 48935 25413 48969
rect 25447 48935 25813 48969
rect 25847 48935 26213 48969
rect 26247 48935 26613 48969
rect 26647 48935 27013 48969
rect 27047 48935 27413 48969
rect 27447 48935 27813 48969
rect 27847 48935 28213 48969
rect 28247 48935 28613 48969
rect 28647 48935 29013 48969
rect 29047 48935 29413 48969
rect 29447 48935 29813 48969
rect 29847 48935 30213 48969
rect 30247 48935 30613 48969
rect 30647 48935 31013 48969
rect 31047 48935 31413 48969
rect 31447 48935 31813 48969
rect 31847 48935 32213 48969
rect 32247 48935 32613 48969
rect 32647 48935 33013 48969
rect 33047 48935 33413 48969
rect 33447 48935 33813 48969
rect 33847 48935 34213 48969
rect 34247 48935 34613 48969
rect 34647 48935 35013 48969
rect 35047 48935 35413 48969
rect 35447 48935 35813 48969
rect 35847 48935 36213 48969
rect 36247 48935 36613 48969
rect 36647 48935 37013 48969
rect 37047 48935 37413 48969
rect 37447 48935 37813 48969
rect 37847 48935 38213 48969
rect 38247 48935 38613 48969
rect 38647 48935 39013 48969
rect 39047 48935 39413 48969
rect 39447 48935 39813 48969
rect 39847 48935 40213 48969
rect 40247 48935 40613 48969
rect 40647 48935 41013 48969
rect 41047 48935 41413 48969
rect 41447 48935 41813 48969
rect 41847 48935 42213 48969
rect 42247 48935 42613 48969
rect 42647 48935 43013 48969
rect 43047 48935 43413 48969
rect 43447 48935 43813 48969
rect 43847 48935 44213 48969
rect 44247 48935 44613 48969
rect 44647 48935 45013 48969
rect 45047 48935 45413 48969
rect 45447 48935 45813 48969
rect 45847 48935 46213 48969
rect 46247 48935 46613 48969
rect 46647 48935 47013 48969
rect 47047 48935 47413 48969
rect 47447 48935 47813 48969
rect 47847 48935 48213 48969
rect 48247 48935 48613 48969
rect 48647 48935 49013 48969
rect 49047 48935 49413 48969
rect 49447 48935 49813 48969
rect 49847 48935 50213 48969
rect 50247 48935 50613 48969
rect 50647 48935 51013 48969
rect 51047 48935 51413 48969
rect 51447 48935 51813 48969
rect 51847 48935 52213 48969
rect 52247 48935 53478 48969
rect 4958 48894 53478 48935
rect 55066 48894 55088 49010
rect 3348 48892 55088 48894
rect 25332 48717 25360 48892
rect 20843 48701 21253 48713
rect 20843 48163 20851 48701
rect 21245 48163 21253 48701
rect 20843 48151 21253 48163
rect 22851 48701 23261 48713
rect 22851 48163 22858 48701
rect 23252 48163 23261 48701
rect 24871 48701 24917 48717
rect 24871 48667 24877 48701
rect 24911 48667 24917 48701
rect 24871 48629 24917 48667
rect 24871 48595 24877 48629
rect 24911 48595 24917 48629
rect 24871 48557 24917 48595
rect 24871 48523 24877 48557
rect 24911 48523 24917 48557
rect 24871 48485 24917 48523
rect 22851 48151 23261 48163
rect 23924 48449 23970 48472
rect 23924 48415 23930 48449
rect 23964 48415 23970 48449
rect 23924 48377 23970 48415
rect 23924 48343 23930 48377
rect 23964 48343 23970 48377
rect 23924 48305 23970 48343
rect 23924 48271 23930 48305
rect 23964 48271 23970 48305
rect 23924 48233 23970 48271
rect 23924 48199 23930 48233
rect 23964 48199 23970 48233
rect 23924 48161 23970 48199
rect 21008 48068 21036 48151
rect 20990 48016 20996 48068
rect 21048 48016 21054 48068
rect 20843 47741 21253 47753
rect 19426 47268 19432 47320
rect 19484 47308 19490 47320
rect 20843 47308 20851 47741
rect 19484 47280 20851 47308
rect 19484 47268 19490 47280
rect 20843 47203 20851 47280
rect 21245 47203 21253 47741
rect 20843 47191 21253 47203
rect 22840 47741 23272 48151
rect 22840 47203 22858 47741
rect 23252 47203 23272 47741
rect 23924 48127 23930 48161
rect 23964 48127 23970 48161
rect 23924 48089 23970 48127
rect 23924 48055 23930 48089
rect 23964 48055 23970 48089
rect 23924 48017 23970 48055
rect 23924 47983 23930 48017
rect 23964 47983 23970 48017
rect 23924 47945 23970 47983
rect 23924 47911 23930 47945
rect 23964 47911 23970 47945
rect 23924 47873 23970 47911
rect 23924 47839 23930 47873
rect 23964 47839 23970 47873
rect 23924 47801 23970 47839
rect 23924 47767 23930 47801
rect 23964 47767 23970 47801
rect 23924 47729 23970 47767
rect 23924 47695 23930 47729
rect 23964 47716 23970 47729
rect 24382 48449 24428 48472
rect 24382 48415 24388 48449
rect 24422 48415 24428 48449
rect 24382 48377 24428 48415
rect 24382 48343 24388 48377
rect 24422 48343 24428 48377
rect 24382 48305 24428 48343
rect 24382 48271 24388 48305
rect 24422 48271 24428 48305
rect 24382 48233 24428 48271
rect 24382 48199 24388 48233
rect 24422 48199 24428 48233
rect 24382 48161 24428 48199
rect 24382 48127 24388 48161
rect 24422 48127 24428 48161
rect 24382 48089 24428 48127
rect 24382 48055 24388 48089
rect 24422 48055 24428 48089
rect 24382 48017 24428 48055
rect 24382 47983 24388 48017
rect 24422 47983 24428 48017
rect 24382 47945 24428 47983
rect 24382 47911 24388 47945
rect 24422 47911 24428 47945
rect 24382 47873 24428 47911
rect 24382 47839 24388 47873
rect 24422 47839 24428 47873
rect 24382 47801 24428 47839
rect 24382 47767 24388 47801
rect 24422 47767 24428 47801
rect 24382 47729 24428 47767
rect 24382 47716 24388 47729
rect 23964 47695 24072 47716
rect 23924 47688 24072 47695
rect 23924 47672 23970 47688
rect 22840 47187 23272 47203
rect 23750 47200 23756 47252
rect 23808 47240 23814 47252
rect 24044 47249 24072 47688
rect 24320 47695 24388 47716
rect 24422 47695 24428 47729
rect 24320 47688 24428 47695
rect 24029 47243 24087 47249
rect 24029 47240 24041 47243
rect 23808 47212 24041 47240
rect 23808 47200 23814 47212
rect 24029 47209 24041 47212
rect 24075 47209 24087 47243
rect 24029 47203 24087 47209
rect 24320 47132 24348 47688
rect 24382 47672 24428 47688
rect 24871 48451 24877 48485
rect 24911 48451 24917 48485
rect 24871 48413 24917 48451
rect 24871 48379 24877 48413
rect 24911 48379 24917 48413
rect 24871 48341 24917 48379
rect 24871 48307 24877 48341
rect 24911 48307 24917 48341
rect 24871 48269 24917 48307
rect 24871 48235 24877 48269
rect 24911 48235 24917 48269
rect 24871 48197 24917 48235
rect 24871 48163 24877 48197
rect 24911 48163 24917 48197
rect 24871 48125 24917 48163
rect 24871 48091 24877 48125
rect 24911 48091 24917 48125
rect 24871 48053 24917 48091
rect 24871 48019 24877 48053
rect 24911 48019 24917 48053
rect 24871 47981 24917 48019
rect 24871 47947 24877 47981
rect 24911 47947 24917 47981
rect 24871 47909 24917 47947
rect 24871 47875 24877 47909
rect 24911 47875 24917 47909
rect 24871 47837 24917 47875
rect 24871 47803 24877 47837
rect 24911 47803 24917 47837
rect 24871 47765 24917 47803
rect 24871 47731 24877 47765
rect 24911 47731 24917 47765
rect 24871 47693 24917 47731
rect 24871 47659 24877 47693
rect 24911 47659 24917 47693
rect 24871 47621 24917 47659
rect 24871 47587 24877 47621
rect 24911 47587 24917 47621
rect 24871 47549 24917 47587
rect 24871 47515 24877 47549
rect 24911 47515 24917 47549
rect 24871 47477 24917 47515
rect 24871 47443 24877 47477
rect 24911 47443 24917 47477
rect 24871 47427 24917 47443
rect 25329 48701 25375 48717
rect 25329 48667 25335 48701
rect 25369 48667 25375 48701
rect 25329 48629 25375 48667
rect 25329 48595 25335 48629
rect 25369 48595 25375 48629
rect 25329 48557 25375 48595
rect 25329 48523 25335 48557
rect 25369 48523 25375 48557
rect 25329 48485 25375 48523
rect 25329 48451 25335 48485
rect 25369 48451 25375 48485
rect 25329 48413 25375 48451
rect 25329 48379 25335 48413
rect 25369 48379 25375 48413
rect 25329 48341 25375 48379
rect 25329 48307 25335 48341
rect 25369 48307 25375 48341
rect 25329 48269 25375 48307
rect 25329 48235 25335 48269
rect 25369 48235 25375 48269
rect 25329 48197 25375 48235
rect 25329 48163 25335 48197
rect 25369 48163 25375 48197
rect 25329 48125 25375 48163
rect 25329 48091 25335 48125
rect 25369 48091 25375 48125
rect 25329 48053 25375 48091
rect 25329 48019 25335 48053
rect 25369 48019 25375 48053
rect 25329 47981 25375 48019
rect 25329 47947 25335 47981
rect 25369 47947 25375 47981
rect 25329 47909 25375 47947
rect 25329 47875 25335 47909
rect 25369 47875 25375 47909
rect 25329 47837 25375 47875
rect 25329 47803 25335 47837
rect 25369 47803 25375 47837
rect 25329 47765 25375 47803
rect 25329 47731 25335 47765
rect 25369 47731 25375 47765
rect 25329 47693 25375 47731
rect 25329 47659 25335 47693
rect 25369 47659 25375 47693
rect 25329 47621 25375 47659
rect 25329 47587 25335 47621
rect 25369 47587 25375 47621
rect 25329 47549 25375 47587
rect 25329 47515 25335 47549
rect 25369 47515 25375 47549
rect 25329 47477 25375 47515
rect 25329 47443 25335 47477
rect 25369 47443 25375 47477
rect 25329 47427 25375 47443
rect 25787 48701 25833 48717
rect 25787 48667 25793 48701
rect 25827 48667 25833 48701
rect 25787 48629 25833 48667
rect 25787 48595 25793 48629
rect 25827 48595 25833 48629
rect 25787 48557 25833 48595
rect 25787 48523 25793 48557
rect 25827 48523 25833 48557
rect 25787 48485 25833 48523
rect 25787 48451 25793 48485
rect 25827 48451 25833 48485
rect 25787 48413 25833 48451
rect 25787 48379 25793 48413
rect 25827 48379 25833 48413
rect 25787 48341 25833 48379
rect 25787 48307 25793 48341
rect 25827 48307 25833 48341
rect 25787 48269 25833 48307
rect 25787 48235 25793 48269
rect 25827 48235 25833 48269
rect 25787 48197 25833 48235
rect 25787 48163 25793 48197
rect 25827 48163 25833 48197
rect 25787 48125 25833 48163
rect 25787 48091 25793 48125
rect 25827 48091 25833 48125
rect 25787 48053 25833 48091
rect 25787 48019 25793 48053
rect 25827 48019 25833 48053
rect 25787 47981 25833 48019
rect 25787 47947 25793 47981
rect 25827 47947 25833 47981
rect 25787 47909 25833 47947
rect 25787 47875 25793 47909
rect 25827 47875 25833 47909
rect 25787 47837 25833 47875
rect 25787 47803 25793 47837
rect 25827 47803 25833 47837
rect 25787 47765 25833 47803
rect 25787 47731 25793 47765
rect 25827 47731 25833 47765
rect 25787 47693 25833 47731
rect 25787 47659 25793 47693
rect 25827 47659 25833 47693
rect 25787 47621 25833 47659
rect 25787 47587 25793 47621
rect 25827 47587 25833 47621
rect 25787 47549 25833 47587
rect 25787 47515 25793 47549
rect 25827 47515 25833 47549
rect 25787 47477 25833 47515
rect 25787 47443 25793 47477
rect 25827 47443 25833 47477
rect 25787 47427 25833 47443
rect 26245 48701 26291 48717
rect 26245 48667 26251 48701
rect 26285 48667 26291 48701
rect 26245 48629 26291 48667
rect 26245 48595 26251 48629
rect 26285 48595 26291 48629
rect 26245 48557 26291 48595
rect 26245 48523 26251 48557
rect 26285 48523 26291 48557
rect 26245 48485 26291 48523
rect 26245 48451 26251 48485
rect 26285 48451 26291 48485
rect 26245 48413 26291 48451
rect 26245 48379 26251 48413
rect 26285 48379 26291 48413
rect 26245 48341 26291 48379
rect 26245 48307 26251 48341
rect 26285 48307 26291 48341
rect 26245 48269 26291 48307
rect 26245 48235 26251 48269
rect 26285 48235 26291 48269
rect 26245 48197 26291 48235
rect 26245 48163 26251 48197
rect 26285 48163 26291 48197
rect 26245 48125 26291 48163
rect 26245 48091 26251 48125
rect 26285 48091 26291 48125
rect 26245 48053 26291 48091
rect 26245 48019 26251 48053
rect 26285 48019 26291 48053
rect 26245 47981 26291 48019
rect 26245 47947 26251 47981
rect 26285 47947 26291 47981
rect 26245 47909 26291 47947
rect 26245 47875 26251 47909
rect 26285 47875 26291 47909
rect 26245 47837 26291 47875
rect 26245 47803 26251 47837
rect 26285 47803 26291 47837
rect 26245 47765 26291 47803
rect 26245 47731 26251 47765
rect 26285 47731 26291 47765
rect 26245 47693 26291 47731
rect 26245 47659 26251 47693
rect 26285 47659 26291 47693
rect 26245 47621 26291 47659
rect 26245 47587 26251 47621
rect 26285 47587 26291 47621
rect 26245 47549 26291 47587
rect 26245 47515 26251 47549
rect 26285 47515 26291 47549
rect 26245 47477 26291 47515
rect 26245 47443 26251 47477
rect 26285 47443 26291 47477
rect 26245 47427 26291 47443
rect 26703 48701 26749 48717
rect 26703 48667 26709 48701
rect 26743 48667 26749 48701
rect 26703 48629 26749 48667
rect 26703 48595 26709 48629
rect 26743 48595 26749 48629
rect 26703 48557 26749 48595
rect 26703 48523 26709 48557
rect 26743 48523 26749 48557
rect 26703 48485 26749 48523
rect 26703 48451 26709 48485
rect 26743 48451 26749 48485
rect 26703 48413 26749 48451
rect 26703 48379 26709 48413
rect 26743 48379 26749 48413
rect 26703 48341 26749 48379
rect 26703 48307 26709 48341
rect 26743 48307 26749 48341
rect 26703 48269 26749 48307
rect 26703 48235 26709 48269
rect 26743 48235 26749 48269
rect 26703 48197 26749 48235
rect 26703 48163 26709 48197
rect 26743 48163 26749 48197
rect 26703 48125 26749 48163
rect 26703 48091 26709 48125
rect 26743 48091 26749 48125
rect 26703 48053 26749 48091
rect 26703 48019 26709 48053
rect 26743 48019 26749 48053
rect 26703 47981 26749 48019
rect 26703 47947 26709 47981
rect 26743 47947 26749 47981
rect 26703 47909 26749 47947
rect 26703 47875 26709 47909
rect 26743 47875 26749 47909
rect 26703 47837 26749 47875
rect 26703 47803 26709 47837
rect 26743 47803 26749 47837
rect 26703 47765 26749 47803
rect 26703 47731 26709 47765
rect 26743 47731 26749 47765
rect 26703 47693 26749 47731
rect 26703 47659 26709 47693
rect 26743 47659 26749 47693
rect 26703 47621 26749 47659
rect 26703 47587 26709 47621
rect 26743 47587 26749 47621
rect 26703 47549 26749 47587
rect 26703 47515 26709 47549
rect 26743 47515 26749 47549
rect 26703 47477 26749 47515
rect 26703 47443 26709 47477
rect 26743 47443 26749 47477
rect 26703 47427 26749 47443
rect 27161 48701 27207 48717
rect 27161 48667 27167 48701
rect 27201 48667 27207 48701
rect 27161 48629 27207 48667
rect 27161 48595 27167 48629
rect 27201 48595 27207 48629
rect 27161 48557 27207 48595
rect 27161 48523 27167 48557
rect 27201 48523 27207 48557
rect 27161 48485 27207 48523
rect 27161 48451 27167 48485
rect 27201 48451 27207 48485
rect 27161 48413 27207 48451
rect 27161 48379 27167 48413
rect 27201 48379 27207 48413
rect 27161 48341 27207 48379
rect 27161 48307 27167 48341
rect 27201 48307 27207 48341
rect 27161 48269 27207 48307
rect 27161 48235 27167 48269
rect 27201 48235 27207 48269
rect 27161 48197 27207 48235
rect 27161 48163 27167 48197
rect 27201 48163 27207 48197
rect 27161 48125 27207 48163
rect 27161 48091 27167 48125
rect 27201 48091 27207 48125
rect 27161 48053 27207 48091
rect 27161 48019 27167 48053
rect 27201 48019 27207 48053
rect 27161 47981 27207 48019
rect 27161 47947 27167 47981
rect 27201 47947 27207 47981
rect 27161 47909 27207 47947
rect 27161 47875 27167 47909
rect 27201 47875 27207 47909
rect 27161 47837 27207 47875
rect 27161 47803 27167 47837
rect 27201 47803 27207 47837
rect 27161 47765 27207 47803
rect 27161 47731 27167 47765
rect 27201 47731 27207 47765
rect 27161 47693 27207 47731
rect 27161 47659 27167 47693
rect 27201 47659 27207 47693
rect 27161 47621 27207 47659
rect 27161 47587 27167 47621
rect 27201 47587 27207 47621
rect 27161 47549 27207 47587
rect 27161 47515 27167 47549
rect 27201 47515 27207 47549
rect 27161 47477 27207 47515
rect 27161 47443 27167 47477
rect 27201 47443 27207 47477
rect 27161 47427 27207 47443
rect 27619 48701 27665 48717
rect 27619 48667 27625 48701
rect 27659 48667 27665 48701
rect 27619 48629 27665 48667
rect 27619 48595 27625 48629
rect 27659 48595 27665 48629
rect 27619 48557 27665 48595
rect 27619 48523 27625 48557
rect 27659 48523 27665 48557
rect 27619 48485 27665 48523
rect 27619 48451 27625 48485
rect 27659 48451 27665 48485
rect 27619 48413 27665 48451
rect 27619 48379 27625 48413
rect 27659 48379 27665 48413
rect 27619 48341 27665 48379
rect 27619 48307 27625 48341
rect 27659 48307 27665 48341
rect 27619 48269 27665 48307
rect 27619 48235 27625 48269
rect 27659 48235 27665 48269
rect 27619 48197 27665 48235
rect 27619 48163 27625 48197
rect 27659 48163 27665 48197
rect 27619 48125 27665 48163
rect 27619 48091 27625 48125
rect 27659 48091 27665 48125
rect 27619 48053 27665 48091
rect 27619 48019 27625 48053
rect 27659 48019 27665 48053
rect 27619 47981 27665 48019
rect 27619 47947 27625 47981
rect 27659 47947 27665 47981
rect 27619 47909 27665 47947
rect 27619 47875 27625 47909
rect 27659 47875 27665 47909
rect 27619 47837 27665 47875
rect 27619 47803 27625 47837
rect 27659 47803 27665 47837
rect 27619 47765 27665 47803
rect 27619 47731 27625 47765
rect 27659 47731 27665 47765
rect 27619 47693 27665 47731
rect 27619 47659 27625 47693
rect 27659 47659 27665 47693
rect 27619 47621 27665 47659
rect 27619 47587 27625 47621
rect 27659 47587 27665 47621
rect 27619 47549 27665 47587
rect 27619 47515 27625 47549
rect 27659 47515 27665 47549
rect 27619 47477 27665 47515
rect 27619 47443 27625 47477
rect 27659 47443 27665 47477
rect 27619 47427 27665 47443
rect 28077 48701 28123 48717
rect 28077 48667 28083 48701
rect 28117 48667 28123 48701
rect 28077 48629 28123 48667
rect 28077 48595 28083 48629
rect 28117 48595 28123 48629
rect 28077 48557 28123 48595
rect 28077 48523 28083 48557
rect 28117 48523 28123 48557
rect 28077 48485 28123 48523
rect 28077 48451 28083 48485
rect 28117 48451 28123 48485
rect 28077 48413 28123 48451
rect 28077 48379 28083 48413
rect 28117 48379 28123 48413
rect 28077 48341 28123 48379
rect 28077 48307 28083 48341
rect 28117 48307 28123 48341
rect 28077 48269 28123 48307
rect 28077 48235 28083 48269
rect 28117 48235 28123 48269
rect 28077 48197 28123 48235
rect 28077 48163 28083 48197
rect 28117 48163 28123 48197
rect 28077 48125 28123 48163
rect 28077 48091 28083 48125
rect 28117 48091 28123 48125
rect 28077 48053 28123 48091
rect 28077 48019 28083 48053
rect 28117 48019 28123 48053
rect 28077 47981 28123 48019
rect 28077 47947 28083 47981
rect 28117 47947 28123 47981
rect 28077 47909 28123 47947
rect 28077 47875 28083 47909
rect 28117 47875 28123 47909
rect 28077 47837 28123 47875
rect 28077 47803 28083 47837
rect 28117 47803 28123 47837
rect 28077 47765 28123 47803
rect 28077 47731 28083 47765
rect 28117 47731 28123 47765
rect 28077 47693 28123 47731
rect 28077 47659 28083 47693
rect 28117 47659 28123 47693
rect 28077 47621 28123 47659
rect 28077 47587 28083 47621
rect 28117 47587 28123 47621
rect 28077 47549 28123 47587
rect 28077 47515 28083 47549
rect 28117 47515 28123 47549
rect 28077 47477 28123 47515
rect 28077 47443 28083 47477
rect 28117 47443 28123 47477
rect 28077 47427 28123 47443
rect 28535 48701 28581 48717
rect 28535 48667 28541 48701
rect 28575 48667 28581 48701
rect 28535 48629 28581 48667
rect 28535 48595 28541 48629
rect 28575 48595 28581 48629
rect 28535 48557 28581 48595
rect 28535 48523 28541 48557
rect 28575 48523 28581 48557
rect 28535 48485 28581 48523
rect 28535 48451 28541 48485
rect 28575 48451 28581 48485
rect 28535 48413 28581 48451
rect 28535 48379 28541 48413
rect 28575 48379 28581 48413
rect 28535 48341 28581 48379
rect 28535 48307 28541 48341
rect 28575 48307 28581 48341
rect 28535 48269 28581 48307
rect 28535 48235 28541 48269
rect 28575 48235 28581 48269
rect 28535 48197 28581 48235
rect 28535 48163 28541 48197
rect 28575 48163 28581 48197
rect 28535 48125 28581 48163
rect 28535 48091 28541 48125
rect 28575 48091 28581 48125
rect 28535 48053 28581 48091
rect 28535 48019 28541 48053
rect 28575 48019 28581 48053
rect 28535 47981 28581 48019
rect 28535 47947 28541 47981
rect 28575 47947 28581 47981
rect 28535 47909 28581 47947
rect 28535 47875 28541 47909
rect 28575 47875 28581 47909
rect 28535 47837 28581 47875
rect 28535 47803 28541 47837
rect 28575 47803 28581 47837
rect 28535 47765 28581 47803
rect 28535 47731 28541 47765
rect 28575 47731 28581 47765
rect 28535 47693 28581 47731
rect 28535 47659 28541 47693
rect 28575 47659 28581 47693
rect 28535 47621 28581 47659
rect 28535 47587 28541 47621
rect 28575 47587 28581 47621
rect 28535 47549 28581 47587
rect 28535 47515 28541 47549
rect 28575 47515 28581 47549
rect 28535 47477 28581 47515
rect 28535 47443 28541 47477
rect 28575 47443 28581 47477
rect 28535 47427 28581 47443
rect 28993 48701 29039 48717
rect 28993 48667 28999 48701
rect 29033 48667 29039 48701
rect 28993 48629 29039 48667
rect 28993 48595 28999 48629
rect 29033 48595 29039 48629
rect 28993 48557 29039 48595
rect 28993 48523 28999 48557
rect 29033 48523 29039 48557
rect 28993 48485 29039 48523
rect 28993 48451 28999 48485
rect 29033 48451 29039 48485
rect 28993 48413 29039 48451
rect 28993 48379 28999 48413
rect 29033 48379 29039 48413
rect 28993 48341 29039 48379
rect 28993 48307 28999 48341
rect 29033 48307 29039 48341
rect 28993 48269 29039 48307
rect 28993 48235 28999 48269
rect 29033 48235 29039 48269
rect 28993 48197 29039 48235
rect 28993 48163 28999 48197
rect 29033 48163 29039 48197
rect 28993 48125 29039 48163
rect 28993 48091 28999 48125
rect 29033 48091 29039 48125
rect 28993 48053 29039 48091
rect 28993 48019 28999 48053
rect 29033 48019 29039 48053
rect 28993 47981 29039 48019
rect 28993 47947 28999 47981
rect 29033 47947 29039 47981
rect 28993 47909 29039 47947
rect 28993 47875 28999 47909
rect 29033 47875 29039 47909
rect 28993 47837 29039 47875
rect 28993 47803 28999 47837
rect 29033 47803 29039 47837
rect 28993 47765 29039 47803
rect 28993 47731 28999 47765
rect 29033 47731 29039 47765
rect 28993 47693 29039 47731
rect 28993 47659 28999 47693
rect 29033 47659 29039 47693
rect 28993 47621 29039 47659
rect 28993 47587 28999 47621
rect 29033 47587 29039 47621
rect 28993 47549 29039 47587
rect 28993 47515 28999 47549
rect 29033 47515 29039 47549
rect 28993 47477 29039 47515
rect 28993 47443 28999 47477
rect 29033 47443 29039 47477
rect 28993 47427 29039 47443
rect 29451 48701 29497 48717
rect 29451 48667 29457 48701
rect 29491 48667 29497 48701
rect 29451 48629 29497 48667
rect 29451 48595 29457 48629
rect 29491 48595 29497 48629
rect 29451 48557 29497 48595
rect 29451 48523 29457 48557
rect 29491 48523 29497 48557
rect 29451 48485 29497 48523
rect 29451 48451 29457 48485
rect 29491 48451 29497 48485
rect 29451 48413 29497 48451
rect 29451 48379 29457 48413
rect 29491 48379 29497 48413
rect 29451 48341 29497 48379
rect 29451 48307 29457 48341
rect 29491 48307 29497 48341
rect 29451 48269 29497 48307
rect 29451 48235 29457 48269
rect 29491 48235 29497 48269
rect 29451 48197 29497 48235
rect 29451 48163 29457 48197
rect 29491 48163 29497 48197
rect 29451 48125 29497 48163
rect 29451 48091 29457 48125
rect 29491 48091 29497 48125
rect 29451 48053 29497 48091
rect 29451 48019 29457 48053
rect 29491 48019 29497 48053
rect 29451 47981 29497 48019
rect 29451 47947 29457 47981
rect 29491 47947 29497 47981
rect 29451 47909 29497 47947
rect 29451 47875 29457 47909
rect 29491 47875 29497 47909
rect 29451 47837 29497 47875
rect 29451 47803 29457 47837
rect 29491 47803 29497 47837
rect 29451 47765 29497 47803
rect 29451 47731 29457 47765
rect 29491 47731 29497 47765
rect 29451 47693 29497 47731
rect 29451 47659 29457 47693
rect 29491 47659 29497 47693
rect 29451 47621 29497 47659
rect 29451 47587 29457 47621
rect 29491 47587 29497 47621
rect 29451 47549 29497 47587
rect 29451 47515 29457 47549
rect 29491 47515 29497 47549
rect 29451 47477 29497 47515
rect 29451 47443 29457 47477
rect 29491 47443 29497 47477
rect 29451 47427 29497 47443
rect 29909 48701 29955 48717
rect 29909 48667 29915 48701
rect 29949 48667 29955 48701
rect 29909 48629 29955 48667
rect 29909 48595 29915 48629
rect 29949 48595 29955 48629
rect 29909 48557 29955 48595
rect 29909 48523 29915 48557
rect 29949 48523 29955 48557
rect 29909 48485 29955 48523
rect 29909 48451 29915 48485
rect 29949 48451 29955 48485
rect 29909 48413 29955 48451
rect 29909 48379 29915 48413
rect 29949 48379 29955 48413
rect 29909 48341 29955 48379
rect 29909 48307 29915 48341
rect 29949 48307 29955 48341
rect 29909 48269 29955 48307
rect 29909 48235 29915 48269
rect 29949 48235 29955 48269
rect 29909 48197 29955 48235
rect 29909 48163 29915 48197
rect 29949 48163 29955 48197
rect 29909 48125 29955 48163
rect 29909 48091 29915 48125
rect 29949 48091 29955 48125
rect 29909 48053 29955 48091
rect 29909 48019 29915 48053
rect 29949 48019 29955 48053
rect 29909 47981 29955 48019
rect 29909 47947 29915 47981
rect 29949 47947 29955 47981
rect 29909 47909 29955 47947
rect 29909 47875 29915 47909
rect 29949 47875 29955 47909
rect 29909 47837 29955 47875
rect 29909 47803 29915 47837
rect 29949 47803 29955 47837
rect 29909 47765 29955 47803
rect 29909 47731 29915 47765
rect 29949 47731 29955 47765
rect 29909 47693 29955 47731
rect 29909 47659 29915 47693
rect 29949 47659 29955 47693
rect 29909 47621 29955 47659
rect 29909 47587 29915 47621
rect 29949 47587 29955 47621
rect 29909 47549 29955 47587
rect 29909 47515 29915 47549
rect 29949 47515 29955 47549
rect 29909 47477 29955 47515
rect 29909 47443 29915 47477
rect 29949 47443 29955 47477
rect 29909 47427 29955 47443
rect 30367 48701 30413 48717
rect 30367 48667 30373 48701
rect 30407 48667 30413 48701
rect 30367 48629 30413 48667
rect 30367 48595 30373 48629
rect 30407 48595 30413 48629
rect 30367 48557 30413 48595
rect 30367 48523 30373 48557
rect 30407 48523 30413 48557
rect 30367 48485 30413 48523
rect 30367 48451 30373 48485
rect 30407 48451 30413 48485
rect 30367 48413 30413 48451
rect 30367 48379 30373 48413
rect 30407 48379 30413 48413
rect 30367 48341 30413 48379
rect 30367 48307 30373 48341
rect 30407 48307 30413 48341
rect 30367 48269 30413 48307
rect 30367 48235 30373 48269
rect 30407 48235 30413 48269
rect 30367 48197 30413 48235
rect 30367 48163 30373 48197
rect 30407 48163 30413 48197
rect 30367 48125 30413 48163
rect 30367 48091 30373 48125
rect 30407 48091 30413 48125
rect 30367 48053 30413 48091
rect 30367 48019 30373 48053
rect 30407 48019 30413 48053
rect 30367 47981 30413 48019
rect 30367 47947 30373 47981
rect 30407 47947 30413 47981
rect 30367 47909 30413 47947
rect 30367 47875 30373 47909
rect 30407 47875 30413 47909
rect 30367 47837 30413 47875
rect 30367 47803 30373 47837
rect 30407 47803 30413 47837
rect 30367 47765 30413 47803
rect 30367 47731 30373 47765
rect 30407 47731 30413 47765
rect 30367 47693 30413 47731
rect 30367 47659 30373 47693
rect 30407 47659 30413 47693
rect 30367 47621 30413 47659
rect 30367 47587 30373 47621
rect 30407 47587 30413 47621
rect 30367 47549 30413 47587
rect 30367 47515 30373 47549
rect 30407 47515 30413 47549
rect 30367 47477 30413 47515
rect 30367 47443 30373 47477
rect 30407 47443 30413 47477
rect 30367 47427 30413 47443
rect 30825 48701 30871 48717
rect 30825 48667 30831 48701
rect 30865 48667 30871 48701
rect 30825 48629 30871 48667
rect 30825 48595 30831 48629
rect 30865 48595 30871 48629
rect 30825 48557 30871 48595
rect 30825 48523 30831 48557
rect 30865 48523 30871 48557
rect 30825 48485 30871 48523
rect 30825 48451 30831 48485
rect 30865 48451 30871 48485
rect 30825 48413 30871 48451
rect 30825 48379 30831 48413
rect 30865 48379 30871 48413
rect 30825 48341 30871 48379
rect 30825 48307 30831 48341
rect 30865 48307 30871 48341
rect 30825 48269 30871 48307
rect 30825 48235 30831 48269
rect 30865 48235 30871 48269
rect 30825 48197 30871 48235
rect 30825 48163 30831 48197
rect 30865 48163 30871 48197
rect 30825 48125 30871 48163
rect 30825 48091 30831 48125
rect 30865 48091 30871 48125
rect 30825 48053 30871 48091
rect 30825 48019 30831 48053
rect 30865 48019 30871 48053
rect 30825 47981 30871 48019
rect 30825 47947 30831 47981
rect 30865 47947 30871 47981
rect 30825 47909 30871 47947
rect 30825 47875 30831 47909
rect 30865 47875 30871 47909
rect 30825 47837 30871 47875
rect 30825 47803 30831 47837
rect 30865 47803 30871 47837
rect 30825 47765 30871 47803
rect 30825 47731 30831 47765
rect 30865 47731 30871 47765
rect 30825 47693 30871 47731
rect 30825 47659 30831 47693
rect 30865 47659 30871 47693
rect 30825 47621 30871 47659
rect 30825 47587 30831 47621
rect 30865 47587 30871 47621
rect 30825 47549 30871 47587
rect 30825 47515 30831 47549
rect 30865 47515 30871 47549
rect 30825 47477 30871 47515
rect 30825 47443 30831 47477
rect 30865 47443 30871 47477
rect 30825 47427 30871 47443
rect 31283 48701 31329 48717
rect 31283 48667 31289 48701
rect 31323 48667 31329 48701
rect 31283 48629 31329 48667
rect 31283 48595 31289 48629
rect 31323 48595 31329 48629
rect 31283 48557 31329 48595
rect 31283 48523 31289 48557
rect 31323 48523 31329 48557
rect 31283 48485 31329 48523
rect 31283 48451 31289 48485
rect 31323 48451 31329 48485
rect 31283 48413 31329 48451
rect 31283 48379 31289 48413
rect 31323 48379 31329 48413
rect 31283 48341 31329 48379
rect 31283 48307 31289 48341
rect 31323 48307 31329 48341
rect 31283 48269 31329 48307
rect 31283 48235 31289 48269
rect 31323 48235 31329 48269
rect 31283 48197 31329 48235
rect 31283 48163 31289 48197
rect 31323 48163 31329 48197
rect 31283 48125 31329 48163
rect 31283 48091 31289 48125
rect 31323 48091 31329 48125
rect 31283 48053 31329 48091
rect 31283 48019 31289 48053
rect 31323 48019 31329 48053
rect 31283 47981 31329 48019
rect 31283 47947 31289 47981
rect 31323 47947 31329 47981
rect 31283 47909 31329 47947
rect 31283 47875 31289 47909
rect 31323 47875 31329 47909
rect 31283 47837 31329 47875
rect 31283 47803 31289 47837
rect 31323 47803 31329 47837
rect 31283 47765 31329 47803
rect 31283 47731 31289 47765
rect 31323 47731 31329 47765
rect 31283 47693 31329 47731
rect 31283 47659 31289 47693
rect 31323 47659 31329 47693
rect 31283 47621 31329 47659
rect 31283 47587 31289 47621
rect 31323 47587 31329 47621
rect 31283 47549 31329 47587
rect 31283 47515 31289 47549
rect 31323 47515 31329 47549
rect 31283 47477 31329 47515
rect 31283 47443 31289 47477
rect 31323 47443 31329 47477
rect 31283 47427 31329 47443
rect 31741 48701 31787 48717
rect 31741 48667 31747 48701
rect 31781 48667 31787 48701
rect 31741 48629 31787 48667
rect 31741 48595 31747 48629
rect 31781 48595 31787 48629
rect 31741 48557 31787 48595
rect 31741 48523 31747 48557
rect 31781 48523 31787 48557
rect 31741 48485 31787 48523
rect 31741 48451 31747 48485
rect 31781 48451 31787 48485
rect 31741 48413 31787 48451
rect 31741 48379 31747 48413
rect 31781 48379 31787 48413
rect 31741 48341 31787 48379
rect 31741 48307 31747 48341
rect 31781 48307 31787 48341
rect 31741 48269 31787 48307
rect 31741 48235 31747 48269
rect 31781 48235 31787 48269
rect 31741 48197 31787 48235
rect 31741 48163 31747 48197
rect 31781 48163 31787 48197
rect 31741 48125 31787 48163
rect 31741 48091 31747 48125
rect 31781 48091 31787 48125
rect 31741 48053 31787 48091
rect 31741 48019 31747 48053
rect 31781 48019 31787 48053
rect 31741 47981 31787 48019
rect 31741 47947 31747 47981
rect 31781 47947 31787 47981
rect 31741 47909 31787 47947
rect 31741 47875 31747 47909
rect 31781 47875 31787 47909
rect 31741 47837 31787 47875
rect 31741 47803 31747 47837
rect 31781 47803 31787 47837
rect 31741 47765 31787 47803
rect 31741 47731 31747 47765
rect 31781 47731 31787 47765
rect 31741 47693 31787 47731
rect 31741 47659 31747 47693
rect 31781 47659 31787 47693
rect 31741 47621 31787 47659
rect 31741 47587 31747 47621
rect 31781 47587 31787 47621
rect 31741 47549 31787 47587
rect 31741 47515 31747 47549
rect 31781 47515 31787 47549
rect 31741 47477 31787 47515
rect 31741 47443 31747 47477
rect 31781 47443 31787 47477
rect 31741 47427 31787 47443
rect 32199 48701 32245 48717
rect 32199 48667 32205 48701
rect 32239 48667 32245 48701
rect 32199 48629 32245 48667
rect 32199 48595 32205 48629
rect 32239 48595 32245 48629
rect 32199 48557 32245 48595
rect 32199 48523 32205 48557
rect 32239 48523 32245 48557
rect 32199 48485 32245 48523
rect 32199 48451 32205 48485
rect 32239 48451 32245 48485
rect 32199 48413 32245 48451
rect 32199 48379 32205 48413
rect 32239 48379 32245 48413
rect 32199 48341 32245 48379
rect 32199 48307 32205 48341
rect 32239 48307 32245 48341
rect 32199 48269 32245 48307
rect 32199 48235 32205 48269
rect 32239 48235 32245 48269
rect 32199 48197 32245 48235
rect 32199 48163 32205 48197
rect 32239 48163 32245 48197
rect 32199 48125 32245 48163
rect 32199 48091 32205 48125
rect 32239 48091 32245 48125
rect 32199 48053 32245 48091
rect 32199 48019 32205 48053
rect 32239 48019 32245 48053
rect 32199 47981 32245 48019
rect 32199 47947 32205 47981
rect 32239 47947 32245 47981
rect 32199 47909 32245 47947
rect 32199 47875 32205 47909
rect 32239 47875 32245 47909
rect 32199 47837 32245 47875
rect 32199 47803 32205 47837
rect 32239 47803 32245 47837
rect 32199 47765 32245 47803
rect 32199 47731 32205 47765
rect 32239 47731 32245 47765
rect 32199 47693 32245 47731
rect 32199 47659 32205 47693
rect 32239 47659 32245 47693
rect 32199 47621 32245 47659
rect 32199 47587 32205 47621
rect 32239 47587 32245 47621
rect 32199 47549 32245 47587
rect 32199 47515 32205 47549
rect 32239 47515 32245 47549
rect 32199 47477 32245 47515
rect 32199 47443 32205 47477
rect 32239 47443 32245 47477
rect 32199 47427 32245 47443
rect 32657 48701 32703 48717
rect 32657 48667 32663 48701
rect 32697 48667 32703 48701
rect 32657 48629 32703 48667
rect 32657 48595 32663 48629
rect 32697 48595 32703 48629
rect 32657 48557 32703 48595
rect 32657 48523 32663 48557
rect 32697 48523 32703 48557
rect 32657 48485 32703 48523
rect 32657 48451 32663 48485
rect 32697 48451 32703 48485
rect 32657 48413 32703 48451
rect 32657 48379 32663 48413
rect 32697 48379 32703 48413
rect 32657 48341 32703 48379
rect 32657 48307 32663 48341
rect 32697 48307 32703 48341
rect 32657 48269 32703 48307
rect 32657 48235 32663 48269
rect 32697 48235 32703 48269
rect 32657 48197 32703 48235
rect 32657 48163 32663 48197
rect 32697 48163 32703 48197
rect 32657 48125 32703 48163
rect 32657 48091 32663 48125
rect 32697 48091 32703 48125
rect 32657 48053 32703 48091
rect 32657 48019 32663 48053
rect 32697 48019 32703 48053
rect 32657 47981 32703 48019
rect 32657 47947 32663 47981
rect 32697 47947 32703 47981
rect 32657 47909 32703 47947
rect 32657 47875 32663 47909
rect 32697 47875 32703 47909
rect 32657 47837 32703 47875
rect 32657 47803 32663 47837
rect 32697 47803 32703 47837
rect 32657 47765 32703 47803
rect 32657 47731 32663 47765
rect 32697 47731 32703 47765
rect 32657 47693 32703 47731
rect 32657 47659 32663 47693
rect 32697 47659 32703 47693
rect 32657 47621 32703 47659
rect 32657 47587 32663 47621
rect 32697 47587 32703 47621
rect 32657 47549 32703 47587
rect 32657 47515 32663 47549
rect 32697 47515 32703 47549
rect 32657 47477 32703 47515
rect 32657 47443 32663 47477
rect 32697 47443 32703 47477
rect 32657 47427 32703 47443
rect 33115 48701 33161 48717
rect 33115 48667 33121 48701
rect 33155 48667 33161 48701
rect 33115 48629 33161 48667
rect 33115 48595 33121 48629
rect 33155 48595 33161 48629
rect 33115 48557 33161 48595
rect 33115 48523 33121 48557
rect 33155 48523 33161 48557
rect 33115 48485 33161 48523
rect 33115 48451 33121 48485
rect 33155 48451 33161 48485
rect 33115 48413 33161 48451
rect 33115 48379 33121 48413
rect 33155 48379 33161 48413
rect 33115 48341 33161 48379
rect 33115 48307 33121 48341
rect 33155 48307 33161 48341
rect 33115 48269 33161 48307
rect 33115 48235 33121 48269
rect 33155 48235 33161 48269
rect 33115 48197 33161 48235
rect 33115 48163 33121 48197
rect 33155 48163 33161 48197
rect 33115 48125 33161 48163
rect 33115 48091 33121 48125
rect 33155 48091 33161 48125
rect 33115 48053 33161 48091
rect 33115 48019 33121 48053
rect 33155 48019 33161 48053
rect 33115 47981 33161 48019
rect 33115 47947 33121 47981
rect 33155 47947 33161 47981
rect 33115 47909 33161 47947
rect 33115 47875 33121 47909
rect 33155 47875 33161 47909
rect 33115 47837 33161 47875
rect 33115 47803 33121 47837
rect 33155 47803 33161 47837
rect 33115 47765 33161 47803
rect 33115 47731 33121 47765
rect 33155 47731 33161 47765
rect 33115 47693 33161 47731
rect 33115 47659 33121 47693
rect 33155 47659 33161 47693
rect 33115 47621 33161 47659
rect 33115 47587 33121 47621
rect 33155 47587 33161 47621
rect 33115 47549 33161 47587
rect 33115 47515 33121 47549
rect 33155 47515 33161 47549
rect 33115 47477 33161 47515
rect 33115 47443 33121 47477
rect 33155 47443 33161 47477
rect 33115 47427 33161 47443
rect 33573 48701 33619 48717
rect 33573 48667 33579 48701
rect 33613 48667 33619 48701
rect 33573 48629 33619 48667
rect 33573 48595 33579 48629
rect 33613 48595 33619 48629
rect 33573 48557 33619 48595
rect 33573 48523 33579 48557
rect 33613 48523 33619 48557
rect 33573 48485 33619 48523
rect 33573 48451 33579 48485
rect 33613 48451 33619 48485
rect 33573 48413 33619 48451
rect 33573 48379 33579 48413
rect 33613 48379 33619 48413
rect 33573 48341 33619 48379
rect 33573 48307 33579 48341
rect 33613 48307 33619 48341
rect 33573 48269 33619 48307
rect 33573 48235 33579 48269
rect 33613 48235 33619 48269
rect 33573 48197 33619 48235
rect 33573 48163 33579 48197
rect 33613 48163 33619 48197
rect 33573 48125 33619 48163
rect 33573 48091 33579 48125
rect 33613 48091 33619 48125
rect 33573 48053 33619 48091
rect 33573 48019 33579 48053
rect 33613 48019 33619 48053
rect 33573 47981 33619 48019
rect 33573 47947 33579 47981
rect 33613 47947 33619 47981
rect 33573 47909 33619 47947
rect 33573 47875 33579 47909
rect 33613 47875 33619 47909
rect 33573 47837 33619 47875
rect 33573 47803 33579 47837
rect 33613 47803 33619 47837
rect 33573 47765 33619 47803
rect 33573 47731 33579 47765
rect 33613 47731 33619 47765
rect 33573 47693 33619 47731
rect 33573 47659 33579 47693
rect 33613 47659 33619 47693
rect 33573 47621 33619 47659
rect 33573 47587 33579 47621
rect 33613 47587 33619 47621
rect 33573 47549 33619 47587
rect 33573 47515 33579 47549
rect 33613 47515 33619 47549
rect 33573 47477 33619 47515
rect 33573 47443 33579 47477
rect 33613 47443 33619 47477
rect 33573 47427 33619 47443
rect 34031 48701 34077 48717
rect 34031 48667 34037 48701
rect 34071 48667 34077 48701
rect 34031 48629 34077 48667
rect 34031 48595 34037 48629
rect 34071 48595 34077 48629
rect 34031 48557 34077 48595
rect 34031 48523 34037 48557
rect 34071 48523 34077 48557
rect 34031 48485 34077 48523
rect 34031 48451 34037 48485
rect 34071 48451 34077 48485
rect 34031 48413 34077 48451
rect 34031 48379 34037 48413
rect 34071 48379 34077 48413
rect 34031 48341 34077 48379
rect 34031 48307 34037 48341
rect 34071 48307 34077 48341
rect 34031 48269 34077 48307
rect 34031 48235 34037 48269
rect 34071 48235 34077 48269
rect 34031 48197 34077 48235
rect 34031 48163 34037 48197
rect 34071 48163 34077 48197
rect 34031 48125 34077 48163
rect 34031 48091 34037 48125
rect 34071 48091 34077 48125
rect 34031 48053 34077 48091
rect 34031 48019 34037 48053
rect 34071 48019 34077 48053
rect 34031 47981 34077 48019
rect 34031 47947 34037 47981
rect 34071 47947 34077 47981
rect 34031 47909 34077 47947
rect 34031 47875 34037 47909
rect 34071 47875 34077 47909
rect 34031 47837 34077 47875
rect 34031 47803 34037 47837
rect 34071 47803 34077 47837
rect 34031 47765 34077 47803
rect 34031 47731 34037 47765
rect 34071 47731 34077 47765
rect 34031 47693 34077 47731
rect 34031 47659 34037 47693
rect 34071 47659 34077 47693
rect 34031 47621 34077 47659
rect 34031 47587 34037 47621
rect 34071 47587 34077 47621
rect 34031 47549 34077 47587
rect 34031 47515 34037 47549
rect 34071 47515 34077 47549
rect 34031 47477 34077 47515
rect 34031 47443 34037 47477
rect 34071 47443 34077 47477
rect 34031 47427 34077 47443
rect 34489 48701 34535 48717
rect 34489 48667 34495 48701
rect 34529 48667 34535 48701
rect 34489 48629 34535 48667
rect 34489 48595 34495 48629
rect 34529 48595 34535 48629
rect 34489 48557 34535 48595
rect 34489 48523 34495 48557
rect 34529 48523 34535 48557
rect 34489 48485 34535 48523
rect 34489 48451 34495 48485
rect 34529 48451 34535 48485
rect 34489 48413 34535 48451
rect 34489 48379 34495 48413
rect 34529 48379 34535 48413
rect 34489 48341 34535 48379
rect 34489 48307 34495 48341
rect 34529 48307 34535 48341
rect 34489 48269 34535 48307
rect 34489 48235 34495 48269
rect 34529 48235 34535 48269
rect 34489 48197 34535 48235
rect 34489 48163 34495 48197
rect 34529 48163 34535 48197
rect 34489 48125 34535 48163
rect 34489 48091 34495 48125
rect 34529 48091 34535 48125
rect 34489 48053 34535 48091
rect 34489 48019 34495 48053
rect 34529 48019 34535 48053
rect 34489 47981 34535 48019
rect 34489 47947 34495 47981
rect 34529 47947 34535 47981
rect 34489 47909 34535 47947
rect 34489 47875 34495 47909
rect 34529 47875 34535 47909
rect 34489 47837 34535 47875
rect 34489 47803 34495 47837
rect 34529 47803 34535 47837
rect 34489 47765 34535 47803
rect 34489 47731 34495 47765
rect 34529 47731 34535 47765
rect 34489 47693 34535 47731
rect 34489 47659 34495 47693
rect 34529 47659 34535 47693
rect 34489 47621 34535 47659
rect 34489 47587 34495 47621
rect 34529 47587 34535 47621
rect 34489 47549 34535 47587
rect 34489 47515 34495 47549
rect 34529 47515 34535 47549
rect 34489 47477 34535 47515
rect 34489 47443 34495 47477
rect 34529 47443 34535 47477
rect 34489 47427 34535 47443
rect 34947 48701 34993 48717
rect 34947 48667 34953 48701
rect 34987 48667 34993 48701
rect 34947 48629 34993 48667
rect 34947 48595 34953 48629
rect 34987 48595 34993 48629
rect 34947 48557 34993 48595
rect 34947 48523 34953 48557
rect 34987 48523 34993 48557
rect 34947 48485 34993 48523
rect 34947 48451 34953 48485
rect 34987 48451 34993 48485
rect 34947 48413 34993 48451
rect 34947 48379 34953 48413
rect 34987 48379 34993 48413
rect 34947 48341 34993 48379
rect 34947 48307 34953 48341
rect 34987 48307 34993 48341
rect 34947 48269 34993 48307
rect 34947 48235 34953 48269
rect 34987 48235 34993 48269
rect 34947 48197 34993 48235
rect 34947 48163 34953 48197
rect 34987 48163 34993 48197
rect 34947 48125 34993 48163
rect 34947 48091 34953 48125
rect 34987 48091 34993 48125
rect 34947 48053 34993 48091
rect 34947 48019 34953 48053
rect 34987 48019 34993 48053
rect 34947 47981 34993 48019
rect 34947 47947 34953 47981
rect 34987 47947 34993 47981
rect 34947 47909 34993 47947
rect 34947 47875 34953 47909
rect 34987 47875 34993 47909
rect 34947 47837 34993 47875
rect 34947 47803 34953 47837
rect 34987 47803 34993 47837
rect 34947 47765 34993 47803
rect 34947 47731 34953 47765
rect 34987 47731 34993 47765
rect 34947 47693 34993 47731
rect 34947 47659 34953 47693
rect 34987 47659 34993 47693
rect 34947 47621 34993 47659
rect 34947 47587 34953 47621
rect 34987 47587 34993 47621
rect 34947 47549 34993 47587
rect 34947 47515 34953 47549
rect 34987 47515 34993 47549
rect 34947 47477 34993 47515
rect 34947 47443 34953 47477
rect 34987 47443 34993 47477
rect 34947 47427 34993 47443
rect 35405 48701 35451 48717
rect 35405 48667 35411 48701
rect 35445 48667 35451 48701
rect 35405 48629 35451 48667
rect 35405 48595 35411 48629
rect 35445 48595 35451 48629
rect 35405 48557 35451 48595
rect 35405 48523 35411 48557
rect 35445 48523 35451 48557
rect 35405 48485 35451 48523
rect 35405 48451 35411 48485
rect 35445 48451 35451 48485
rect 35405 48413 35451 48451
rect 35405 48379 35411 48413
rect 35445 48379 35451 48413
rect 35405 48341 35451 48379
rect 35405 48307 35411 48341
rect 35445 48307 35451 48341
rect 35405 48269 35451 48307
rect 35405 48235 35411 48269
rect 35445 48235 35451 48269
rect 35405 48197 35451 48235
rect 35405 48163 35411 48197
rect 35445 48163 35451 48197
rect 35405 48125 35451 48163
rect 35405 48091 35411 48125
rect 35445 48091 35451 48125
rect 35405 48053 35451 48091
rect 35405 48019 35411 48053
rect 35445 48019 35451 48053
rect 35405 47981 35451 48019
rect 35405 47947 35411 47981
rect 35445 47947 35451 47981
rect 35405 47909 35451 47947
rect 35405 47875 35411 47909
rect 35445 47875 35451 47909
rect 35405 47837 35451 47875
rect 35405 47803 35411 47837
rect 35445 47803 35451 47837
rect 35405 47765 35451 47803
rect 35405 47731 35411 47765
rect 35445 47731 35451 47765
rect 35405 47693 35451 47731
rect 35405 47659 35411 47693
rect 35445 47659 35451 47693
rect 35405 47621 35451 47659
rect 35405 47587 35411 47621
rect 35445 47587 35451 47621
rect 35405 47549 35451 47587
rect 35405 47515 35411 47549
rect 35445 47515 35451 47549
rect 35405 47477 35451 47515
rect 35405 47443 35411 47477
rect 35445 47443 35451 47477
rect 35405 47427 35451 47443
rect 35863 48701 35909 48717
rect 35863 48667 35869 48701
rect 35903 48667 35909 48701
rect 35863 48629 35909 48667
rect 35863 48595 35869 48629
rect 35903 48595 35909 48629
rect 35863 48557 35909 48595
rect 35863 48523 35869 48557
rect 35903 48523 35909 48557
rect 35863 48485 35909 48523
rect 35863 48451 35869 48485
rect 35903 48451 35909 48485
rect 35863 48413 35909 48451
rect 35863 48379 35869 48413
rect 35903 48379 35909 48413
rect 35863 48341 35909 48379
rect 35863 48307 35869 48341
rect 35903 48307 35909 48341
rect 35863 48269 35909 48307
rect 35863 48235 35869 48269
rect 35903 48235 35909 48269
rect 35863 48197 35909 48235
rect 35863 48163 35869 48197
rect 35903 48163 35909 48197
rect 35863 48125 35909 48163
rect 35863 48091 35869 48125
rect 35903 48091 35909 48125
rect 35863 48053 35909 48091
rect 35863 48019 35869 48053
rect 35903 48019 35909 48053
rect 35863 47981 35909 48019
rect 35863 47947 35869 47981
rect 35903 47947 35909 47981
rect 35863 47909 35909 47947
rect 35863 47875 35869 47909
rect 35903 47875 35909 47909
rect 35863 47837 35909 47875
rect 35863 47803 35869 47837
rect 35903 47803 35909 47837
rect 35863 47765 35909 47803
rect 35863 47731 35869 47765
rect 35903 47731 35909 47765
rect 35863 47693 35909 47731
rect 35863 47659 35869 47693
rect 35903 47659 35909 47693
rect 35863 47621 35909 47659
rect 35863 47587 35869 47621
rect 35903 47587 35909 47621
rect 35863 47549 35909 47587
rect 35863 47515 35869 47549
rect 35903 47515 35909 47549
rect 35863 47477 35909 47515
rect 35863 47443 35869 47477
rect 35903 47443 35909 47477
rect 35863 47427 35909 47443
rect 36321 48701 36367 48717
rect 36321 48667 36327 48701
rect 36361 48667 36367 48701
rect 36321 48629 36367 48667
rect 36321 48595 36327 48629
rect 36361 48595 36367 48629
rect 36321 48557 36367 48595
rect 36321 48523 36327 48557
rect 36361 48523 36367 48557
rect 36321 48485 36367 48523
rect 36321 48451 36327 48485
rect 36361 48451 36367 48485
rect 36321 48413 36367 48451
rect 36321 48379 36327 48413
rect 36361 48379 36367 48413
rect 36321 48341 36367 48379
rect 36321 48307 36327 48341
rect 36361 48307 36367 48341
rect 36321 48269 36367 48307
rect 36321 48235 36327 48269
rect 36361 48235 36367 48269
rect 36321 48197 36367 48235
rect 36321 48163 36327 48197
rect 36361 48163 36367 48197
rect 36321 48125 36367 48163
rect 36321 48091 36327 48125
rect 36361 48091 36367 48125
rect 36321 48053 36367 48091
rect 36321 48019 36327 48053
rect 36361 48019 36367 48053
rect 36321 47981 36367 48019
rect 36321 47947 36327 47981
rect 36361 47947 36367 47981
rect 36321 47909 36367 47947
rect 36321 47875 36327 47909
rect 36361 47875 36367 47909
rect 36321 47837 36367 47875
rect 36321 47803 36327 47837
rect 36361 47803 36367 47837
rect 36321 47765 36367 47803
rect 36321 47731 36327 47765
rect 36361 47731 36367 47765
rect 36321 47693 36367 47731
rect 36321 47659 36327 47693
rect 36361 47659 36367 47693
rect 36321 47621 36367 47659
rect 36321 47587 36327 47621
rect 36361 47587 36367 47621
rect 36321 47549 36367 47587
rect 36321 47515 36327 47549
rect 36361 47515 36367 47549
rect 36321 47477 36367 47515
rect 36321 47443 36327 47477
rect 36361 47443 36367 47477
rect 36321 47427 36367 47443
rect 36779 48701 36825 48717
rect 36779 48667 36785 48701
rect 36819 48667 36825 48701
rect 36779 48629 36825 48667
rect 36779 48595 36785 48629
rect 36819 48595 36825 48629
rect 36779 48557 36825 48595
rect 36779 48523 36785 48557
rect 36819 48523 36825 48557
rect 36779 48485 36825 48523
rect 36779 48451 36785 48485
rect 36819 48451 36825 48485
rect 36779 48413 36825 48451
rect 36779 48379 36785 48413
rect 36819 48379 36825 48413
rect 36779 48341 36825 48379
rect 36779 48307 36785 48341
rect 36819 48307 36825 48341
rect 36779 48269 36825 48307
rect 36779 48235 36785 48269
rect 36819 48235 36825 48269
rect 36779 48197 36825 48235
rect 36779 48163 36785 48197
rect 36819 48163 36825 48197
rect 36779 48125 36825 48163
rect 36779 48091 36785 48125
rect 36819 48091 36825 48125
rect 36779 48053 36825 48091
rect 36779 48019 36785 48053
rect 36819 48019 36825 48053
rect 36779 47981 36825 48019
rect 36779 47947 36785 47981
rect 36819 47947 36825 47981
rect 36779 47909 36825 47947
rect 36779 47875 36785 47909
rect 36819 47875 36825 47909
rect 36779 47837 36825 47875
rect 36779 47803 36785 47837
rect 36819 47803 36825 47837
rect 36779 47765 36825 47803
rect 36779 47731 36785 47765
rect 36819 47731 36825 47765
rect 36779 47693 36825 47731
rect 36779 47659 36785 47693
rect 36819 47659 36825 47693
rect 36779 47621 36825 47659
rect 36779 47587 36785 47621
rect 36819 47587 36825 47621
rect 36779 47549 36825 47587
rect 36779 47515 36785 47549
rect 36819 47515 36825 47549
rect 36779 47477 36825 47515
rect 36779 47443 36785 47477
rect 36819 47443 36825 47477
rect 36779 47427 36825 47443
rect 37237 48701 37283 48717
rect 37237 48667 37243 48701
rect 37277 48667 37283 48701
rect 37237 48629 37283 48667
rect 37237 48595 37243 48629
rect 37277 48595 37283 48629
rect 37237 48557 37283 48595
rect 37237 48523 37243 48557
rect 37277 48523 37283 48557
rect 37237 48485 37283 48523
rect 37237 48451 37243 48485
rect 37277 48451 37283 48485
rect 37237 48413 37283 48451
rect 37237 48379 37243 48413
rect 37277 48379 37283 48413
rect 37237 48341 37283 48379
rect 37237 48307 37243 48341
rect 37277 48307 37283 48341
rect 37237 48269 37283 48307
rect 37237 48235 37243 48269
rect 37277 48235 37283 48269
rect 37237 48197 37283 48235
rect 37237 48163 37243 48197
rect 37277 48163 37283 48197
rect 37237 48125 37283 48163
rect 37237 48091 37243 48125
rect 37277 48091 37283 48125
rect 37237 48053 37283 48091
rect 37237 48019 37243 48053
rect 37277 48019 37283 48053
rect 37237 47981 37283 48019
rect 37237 47947 37243 47981
rect 37277 47947 37283 47981
rect 37237 47909 37283 47947
rect 37237 47875 37243 47909
rect 37277 47875 37283 47909
rect 37237 47837 37283 47875
rect 37237 47803 37243 47837
rect 37277 47803 37283 47837
rect 37237 47765 37283 47803
rect 37237 47731 37243 47765
rect 37277 47731 37283 47765
rect 37237 47693 37283 47731
rect 37237 47659 37243 47693
rect 37277 47659 37283 47693
rect 37237 47621 37283 47659
rect 37237 47587 37243 47621
rect 37277 47587 37283 47621
rect 37237 47549 37283 47587
rect 37237 47515 37243 47549
rect 37277 47515 37283 47549
rect 37237 47477 37283 47515
rect 37237 47443 37243 47477
rect 37277 47443 37283 47477
rect 37237 47427 37283 47443
rect 37695 48701 37741 48717
rect 37695 48667 37701 48701
rect 37735 48667 37741 48701
rect 37695 48629 37741 48667
rect 37695 48595 37701 48629
rect 37735 48595 37741 48629
rect 37695 48557 37741 48595
rect 37695 48523 37701 48557
rect 37735 48523 37741 48557
rect 37695 48485 37741 48523
rect 37695 48451 37701 48485
rect 37735 48451 37741 48485
rect 37695 48413 37741 48451
rect 37695 48379 37701 48413
rect 37735 48379 37741 48413
rect 37695 48341 37741 48379
rect 37695 48307 37701 48341
rect 37735 48307 37741 48341
rect 37695 48269 37741 48307
rect 37695 48235 37701 48269
rect 37735 48235 37741 48269
rect 37695 48197 37741 48235
rect 37695 48163 37701 48197
rect 37735 48163 37741 48197
rect 37695 48125 37741 48163
rect 37695 48091 37701 48125
rect 37735 48091 37741 48125
rect 37695 48053 37741 48091
rect 37695 48019 37701 48053
rect 37735 48019 37741 48053
rect 37695 47981 37741 48019
rect 37695 47947 37701 47981
rect 37735 47947 37741 47981
rect 37695 47909 37741 47947
rect 37695 47875 37701 47909
rect 37735 47875 37741 47909
rect 37695 47837 37741 47875
rect 37695 47803 37701 47837
rect 37735 47803 37741 47837
rect 37695 47765 37741 47803
rect 37695 47731 37701 47765
rect 37735 47731 37741 47765
rect 37695 47693 37741 47731
rect 37695 47659 37701 47693
rect 37735 47659 37741 47693
rect 37695 47621 37741 47659
rect 37695 47587 37701 47621
rect 37735 47587 37741 47621
rect 37695 47549 37741 47587
rect 37695 47515 37701 47549
rect 37735 47515 37741 47549
rect 37695 47477 37741 47515
rect 37695 47443 37701 47477
rect 37735 47443 37741 47477
rect 37695 47427 37741 47443
rect 38153 48701 38199 48717
rect 38153 48667 38159 48701
rect 38193 48667 38199 48701
rect 38153 48629 38199 48667
rect 38153 48595 38159 48629
rect 38193 48595 38199 48629
rect 38153 48557 38199 48595
rect 38153 48523 38159 48557
rect 38193 48523 38199 48557
rect 38153 48485 38199 48523
rect 38153 48451 38159 48485
rect 38193 48451 38199 48485
rect 38153 48413 38199 48451
rect 38153 48379 38159 48413
rect 38193 48379 38199 48413
rect 38153 48341 38199 48379
rect 38153 48307 38159 48341
rect 38193 48307 38199 48341
rect 38153 48269 38199 48307
rect 38153 48235 38159 48269
rect 38193 48235 38199 48269
rect 38153 48197 38199 48235
rect 38153 48163 38159 48197
rect 38193 48163 38199 48197
rect 38153 48125 38199 48163
rect 38153 48091 38159 48125
rect 38193 48091 38199 48125
rect 38153 48053 38199 48091
rect 38153 48019 38159 48053
rect 38193 48019 38199 48053
rect 38153 47981 38199 48019
rect 38153 47947 38159 47981
rect 38193 47947 38199 47981
rect 38153 47909 38199 47947
rect 38153 47875 38159 47909
rect 38193 47875 38199 47909
rect 38153 47837 38199 47875
rect 38153 47803 38159 47837
rect 38193 47803 38199 47837
rect 38153 47765 38199 47803
rect 38153 47731 38159 47765
rect 38193 47731 38199 47765
rect 38153 47693 38199 47731
rect 38153 47659 38159 47693
rect 38193 47659 38199 47693
rect 38153 47621 38199 47659
rect 38153 47587 38159 47621
rect 38193 47587 38199 47621
rect 38153 47549 38199 47587
rect 38153 47515 38159 47549
rect 38193 47515 38199 47549
rect 38153 47477 38199 47515
rect 38153 47443 38159 47477
rect 38193 47443 38199 47477
rect 38153 47427 38199 47443
rect 38611 48701 38657 48717
rect 38611 48667 38617 48701
rect 38651 48667 38657 48701
rect 38611 48629 38657 48667
rect 38611 48595 38617 48629
rect 38651 48595 38657 48629
rect 38611 48557 38657 48595
rect 38611 48523 38617 48557
rect 38651 48523 38657 48557
rect 38611 48485 38657 48523
rect 38611 48451 38617 48485
rect 38651 48451 38657 48485
rect 38611 48413 38657 48451
rect 38611 48379 38617 48413
rect 38651 48379 38657 48413
rect 38611 48341 38657 48379
rect 38611 48307 38617 48341
rect 38651 48307 38657 48341
rect 38611 48269 38657 48307
rect 38611 48235 38617 48269
rect 38651 48235 38657 48269
rect 38611 48197 38657 48235
rect 38611 48163 38617 48197
rect 38651 48163 38657 48197
rect 38611 48125 38657 48163
rect 38611 48091 38617 48125
rect 38651 48091 38657 48125
rect 38611 48053 38657 48091
rect 38611 48019 38617 48053
rect 38651 48019 38657 48053
rect 38611 47981 38657 48019
rect 38611 47947 38617 47981
rect 38651 47947 38657 47981
rect 38611 47909 38657 47947
rect 38611 47875 38617 47909
rect 38651 47875 38657 47909
rect 38611 47837 38657 47875
rect 38611 47803 38617 47837
rect 38651 47803 38657 47837
rect 38611 47765 38657 47803
rect 38611 47731 38617 47765
rect 38651 47731 38657 47765
rect 38611 47693 38657 47731
rect 38611 47659 38617 47693
rect 38651 47659 38657 47693
rect 38611 47621 38657 47659
rect 38611 47587 38617 47621
rect 38651 47587 38657 47621
rect 38611 47549 38657 47587
rect 38611 47515 38617 47549
rect 38651 47515 38657 47549
rect 38611 47477 38657 47515
rect 38611 47443 38617 47477
rect 38651 47443 38657 47477
rect 38611 47427 38657 47443
rect 39069 48701 39115 48717
rect 39069 48667 39075 48701
rect 39109 48667 39115 48701
rect 39069 48629 39115 48667
rect 39069 48595 39075 48629
rect 39109 48595 39115 48629
rect 39069 48557 39115 48595
rect 39069 48523 39075 48557
rect 39109 48523 39115 48557
rect 39069 48485 39115 48523
rect 39069 48451 39075 48485
rect 39109 48451 39115 48485
rect 39069 48413 39115 48451
rect 39069 48379 39075 48413
rect 39109 48379 39115 48413
rect 39069 48341 39115 48379
rect 39069 48307 39075 48341
rect 39109 48307 39115 48341
rect 39069 48269 39115 48307
rect 39069 48235 39075 48269
rect 39109 48235 39115 48269
rect 39069 48197 39115 48235
rect 39069 48163 39075 48197
rect 39109 48163 39115 48197
rect 39069 48125 39115 48163
rect 39069 48091 39075 48125
rect 39109 48091 39115 48125
rect 39069 48053 39115 48091
rect 39069 48019 39075 48053
rect 39109 48019 39115 48053
rect 39069 47981 39115 48019
rect 39069 47947 39075 47981
rect 39109 47947 39115 47981
rect 39069 47909 39115 47947
rect 39069 47875 39075 47909
rect 39109 47875 39115 47909
rect 39069 47837 39115 47875
rect 39069 47803 39075 47837
rect 39109 47803 39115 47837
rect 39069 47765 39115 47803
rect 39069 47731 39075 47765
rect 39109 47731 39115 47765
rect 39069 47693 39115 47731
rect 39069 47659 39075 47693
rect 39109 47659 39115 47693
rect 39069 47621 39115 47659
rect 39069 47587 39075 47621
rect 39109 47587 39115 47621
rect 39069 47549 39115 47587
rect 39069 47515 39075 47549
rect 39109 47515 39115 47549
rect 39069 47477 39115 47515
rect 39069 47443 39075 47477
rect 39109 47443 39115 47477
rect 39069 47427 39115 47443
rect 39527 48701 39573 48717
rect 39527 48667 39533 48701
rect 39567 48667 39573 48701
rect 39527 48629 39573 48667
rect 39527 48595 39533 48629
rect 39567 48595 39573 48629
rect 39527 48557 39573 48595
rect 39527 48523 39533 48557
rect 39567 48523 39573 48557
rect 39527 48485 39573 48523
rect 39527 48451 39533 48485
rect 39567 48451 39573 48485
rect 39527 48413 39573 48451
rect 39527 48379 39533 48413
rect 39567 48379 39573 48413
rect 39527 48341 39573 48379
rect 39527 48307 39533 48341
rect 39567 48307 39573 48341
rect 39527 48269 39573 48307
rect 39527 48235 39533 48269
rect 39567 48235 39573 48269
rect 39527 48197 39573 48235
rect 39527 48163 39533 48197
rect 39567 48163 39573 48197
rect 39527 48125 39573 48163
rect 39527 48091 39533 48125
rect 39567 48091 39573 48125
rect 39527 48053 39573 48091
rect 39527 48019 39533 48053
rect 39567 48019 39573 48053
rect 39527 47981 39573 48019
rect 39527 47947 39533 47981
rect 39567 47947 39573 47981
rect 39527 47909 39573 47947
rect 39527 47875 39533 47909
rect 39567 47875 39573 47909
rect 39527 47837 39573 47875
rect 39527 47803 39533 47837
rect 39567 47803 39573 47837
rect 39527 47765 39573 47803
rect 39527 47731 39533 47765
rect 39567 47731 39573 47765
rect 39527 47693 39573 47731
rect 39527 47659 39533 47693
rect 39567 47659 39573 47693
rect 39527 47621 39573 47659
rect 39527 47587 39533 47621
rect 39567 47587 39573 47621
rect 39527 47549 39573 47587
rect 39527 47515 39533 47549
rect 39567 47515 39573 47549
rect 39527 47477 39573 47515
rect 39527 47443 39533 47477
rect 39567 47443 39573 47477
rect 39527 47427 39573 47443
rect 39985 48701 40031 48717
rect 39985 48667 39991 48701
rect 40025 48667 40031 48701
rect 39985 48629 40031 48667
rect 39985 48595 39991 48629
rect 40025 48595 40031 48629
rect 39985 48557 40031 48595
rect 39985 48523 39991 48557
rect 40025 48523 40031 48557
rect 39985 48485 40031 48523
rect 39985 48451 39991 48485
rect 40025 48451 40031 48485
rect 39985 48413 40031 48451
rect 39985 48379 39991 48413
rect 40025 48379 40031 48413
rect 39985 48341 40031 48379
rect 39985 48307 39991 48341
rect 40025 48307 40031 48341
rect 39985 48269 40031 48307
rect 39985 48235 39991 48269
rect 40025 48235 40031 48269
rect 39985 48197 40031 48235
rect 39985 48163 39991 48197
rect 40025 48163 40031 48197
rect 39985 48125 40031 48163
rect 39985 48091 39991 48125
rect 40025 48091 40031 48125
rect 39985 48053 40031 48091
rect 39985 48019 39991 48053
rect 40025 48019 40031 48053
rect 39985 47981 40031 48019
rect 39985 47947 39991 47981
rect 40025 47947 40031 47981
rect 39985 47909 40031 47947
rect 39985 47875 39991 47909
rect 40025 47875 40031 47909
rect 39985 47837 40031 47875
rect 39985 47803 39991 47837
rect 40025 47803 40031 47837
rect 39985 47765 40031 47803
rect 39985 47731 39991 47765
rect 40025 47731 40031 47765
rect 39985 47693 40031 47731
rect 39985 47659 39991 47693
rect 40025 47659 40031 47693
rect 39985 47621 40031 47659
rect 39985 47587 39991 47621
rect 40025 47587 40031 47621
rect 39985 47549 40031 47587
rect 39985 47515 39991 47549
rect 40025 47515 40031 47549
rect 39985 47477 40031 47515
rect 39985 47443 39991 47477
rect 40025 47443 40031 47477
rect 39985 47427 40031 47443
rect 40443 48701 40489 48717
rect 40443 48667 40449 48701
rect 40483 48667 40489 48701
rect 40443 48629 40489 48667
rect 40443 48595 40449 48629
rect 40483 48595 40489 48629
rect 40443 48557 40489 48595
rect 40443 48523 40449 48557
rect 40483 48523 40489 48557
rect 40443 48485 40489 48523
rect 40443 48451 40449 48485
rect 40483 48451 40489 48485
rect 40443 48413 40489 48451
rect 40443 48379 40449 48413
rect 40483 48379 40489 48413
rect 40443 48341 40489 48379
rect 40443 48307 40449 48341
rect 40483 48307 40489 48341
rect 40443 48269 40489 48307
rect 40443 48235 40449 48269
rect 40483 48235 40489 48269
rect 40443 48197 40489 48235
rect 40443 48163 40449 48197
rect 40483 48163 40489 48197
rect 40443 48125 40489 48163
rect 40443 48091 40449 48125
rect 40483 48091 40489 48125
rect 40443 48053 40489 48091
rect 40443 48019 40449 48053
rect 40483 48019 40489 48053
rect 40443 47981 40489 48019
rect 40443 47947 40449 47981
rect 40483 47947 40489 47981
rect 40443 47909 40489 47947
rect 40443 47875 40449 47909
rect 40483 47875 40489 47909
rect 40443 47837 40489 47875
rect 40443 47803 40449 47837
rect 40483 47803 40489 47837
rect 40443 47765 40489 47803
rect 40443 47731 40449 47765
rect 40483 47731 40489 47765
rect 40443 47693 40489 47731
rect 40443 47659 40449 47693
rect 40483 47659 40489 47693
rect 40443 47621 40489 47659
rect 40443 47587 40449 47621
rect 40483 47587 40489 47621
rect 40443 47549 40489 47587
rect 40443 47515 40449 47549
rect 40483 47515 40489 47549
rect 40443 47477 40489 47515
rect 40443 47443 40449 47477
rect 40483 47443 40489 47477
rect 40443 47427 40489 47443
rect 40901 48701 40947 48717
rect 40901 48667 40907 48701
rect 40941 48667 40947 48701
rect 40901 48629 40947 48667
rect 40901 48595 40907 48629
rect 40941 48595 40947 48629
rect 40901 48557 40947 48595
rect 40901 48523 40907 48557
rect 40941 48523 40947 48557
rect 40901 48485 40947 48523
rect 40901 48451 40907 48485
rect 40941 48451 40947 48485
rect 40901 48413 40947 48451
rect 40901 48379 40907 48413
rect 40941 48379 40947 48413
rect 40901 48341 40947 48379
rect 40901 48307 40907 48341
rect 40941 48307 40947 48341
rect 40901 48269 40947 48307
rect 40901 48235 40907 48269
rect 40941 48235 40947 48269
rect 40901 48197 40947 48235
rect 40901 48163 40907 48197
rect 40941 48163 40947 48197
rect 40901 48125 40947 48163
rect 40901 48091 40907 48125
rect 40941 48091 40947 48125
rect 40901 48053 40947 48091
rect 40901 48019 40907 48053
rect 40941 48019 40947 48053
rect 40901 47981 40947 48019
rect 40901 47947 40907 47981
rect 40941 47947 40947 47981
rect 40901 47909 40947 47947
rect 40901 47875 40907 47909
rect 40941 47875 40947 47909
rect 40901 47837 40947 47875
rect 40901 47803 40907 47837
rect 40941 47803 40947 47837
rect 40901 47765 40947 47803
rect 40901 47731 40907 47765
rect 40941 47731 40947 47765
rect 40901 47693 40947 47731
rect 40901 47659 40907 47693
rect 40941 47659 40947 47693
rect 40901 47621 40947 47659
rect 40901 47587 40907 47621
rect 40941 47587 40947 47621
rect 40901 47549 40947 47587
rect 40901 47515 40907 47549
rect 40941 47515 40947 47549
rect 40901 47477 40947 47515
rect 40901 47443 40907 47477
rect 40941 47443 40947 47477
rect 40901 47427 40947 47443
rect 41359 48701 41405 48717
rect 41359 48667 41365 48701
rect 41399 48667 41405 48701
rect 41359 48629 41405 48667
rect 41359 48595 41365 48629
rect 41399 48595 41405 48629
rect 41359 48557 41405 48595
rect 41359 48523 41365 48557
rect 41399 48523 41405 48557
rect 41359 48485 41405 48523
rect 41359 48451 41365 48485
rect 41399 48451 41405 48485
rect 41359 48413 41405 48451
rect 41359 48379 41365 48413
rect 41399 48379 41405 48413
rect 41359 48341 41405 48379
rect 41359 48307 41365 48341
rect 41399 48307 41405 48341
rect 41359 48269 41405 48307
rect 41359 48235 41365 48269
rect 41399 48235 41405 48269
rect 41359 48197 41405 48235
rect 41359 48163 41365 48197
rect 41399 48163 41405 48197
rect 41359 48125 41405 48163
rect 41359 48091 41365 48125
rect 41399 48091 41405 48125
rect 41359 48053 41405 48091
rect 41359 48019 41365 48053
rect 41399 48019 41405 48053
rect 41359 47981 41405 48019
rect 41359 47947 41365 47981
rect 41399 47947 41405 47981
rect 41359 47909 41405 47947
rect 41359 47875 41365 47909
rect 41399 47875 41405 47909
rect 41359 47837 41405 47875
rect 41359 47803 41365 47837
rect 41399 47803 41405 47837
rect 41359 47765 41405 47803
rect 41359 47731 41365 47765
rect 41399 47731 41405 47765
rect 41359 47693 41405 47731
rect 41359 47659 41365 47693
rect 41399 47659 41405 47693
rect 41359 47621 41405 47659
rect 41359 47587 41365 47621
rect 41399 47587 41405 47621
rect 41359 47549 41405 47587
rect 41359 47515 41365 47549
rect 41399 47515 41405 47549
rect 41359 47477 41405 47515
rect 41359 47443 41365 47477
rect 41399 47443 41405 47477
rect 41359 47427 41405 47443
rect 41817 48701 41863 48717
rect 41817 48667 41823 48701
rect 41857 48667 41863 48701
rect 41817 48629 41863 48667
rect 41817 48595 41823 48629
rect 41857 48595 41863 48629
rect 41817 48557 41863 48595
rect 41817 48523 41823 48557
rect 41857 48523 41863 48557
rect 41817 48485 41863 48523
rect 41817 48451 41823 48485
rect 41857 48451 41863 48485
rect 41817 48413 41863 48451
rect 41817 48379 41823 48413
rect 41857 48379 41863 48413
rect 41817 48341 41863 48379
rect 41817 48307 41823 48341
rect 41857 48307 41863 48341
rect 41817 48269 41863 48307
rect 41817 48235 41823 48269
rect 41857 48235 41863 48269
rect 41817 48197 41863 48235
rect 41817 48163 41823 48197
rect 41857 48163 41863 48197
rect 41817 48125 41863 48163
rect 41817 48091 41823 48125
rect 41857 48091 41863 48125
rect 41817 48053 41863 48091
rect 41817 48019 41823 48053
rect 41857 48019 41863 48053
rect 41817 47981 41863 48019
rect 41817 47947 41823 47981
rect 41857 47947 41863 47981
rect 41817 47909 41863 47947
rect 41817 47875 41823 47909
rect 41857 47875 41863 47909
rect 41817 47837 41863 47875
rect 41817 47803 41823 47837
rect 41857 47803 41863 47837
rect 41817 47765 41863 47803
rect 41817 47731 41823 47765
rect 41857 47731 41863 47765
rect 41817 47693 41863 47731
rect 41817 47659 41823 47693
rect 41857 47659 41863 47693
rect 41817 47621 41863 47659
rect 41817 47587 41823 47621
rect 41857 47587 41863 47621
rect 41817 47549 41863 47587
rect 41817 47515 41823 47549
rect 41857 47515 41863 47549
rect 41817 47477 41863 47515
rect 41817 47443 41823 47477
rect 41857 47443 41863 47477
rect 41817 47427 41863 47443
rect 42275 48701 42321 48717
rect 42275 48667 42281 48701
rect 42315 48667 42321 48701
rect 42275 48629 42321 48667
rect 42275 48595 42281 48629
rect 42315 48595 42321 48629
rect 42275 48557 42321 48595
rect 42275 48523 42281 48557
rect 42315 48523 42321 48557
rect 42275 48485 42321 48523
rect 42275 48451 42281 48485
rect 42315 48451 42321 48485
rect 42275 48413 42321 48451
rect 42275 48379 42281 48413
rect 42315 48379 42321 48413
rect 42275 48341 42321 48379
rect 42275 48307 42281 48341
rect 42315 48307 42321 48341
rect 42275 48269 42321 48307
rect 42275 48235 42281 48269
rect 42315 48235 42321 48269
rect 42275 48197 42321 48235
rect 42275 48163 42281 48197
rect 42315 48163 42321 48197
rect 42275 48125 42321 48163
rect 42275 48091 42281 48125
rect 42315 48091 42321 48125
rect 42275 48053 42321 48091
rect 42275 48019 42281 48053
rect 42315 48019 42321 48053
rect 42275 47981 42321 48019
rect 42275 47947 42281 47981
rect 42315 47947 42321 47981
rect 42275 47909 42321 47947
rect 42275 47875 42281 47909
rect 42315 47875 42321 47909
rect 42275 47837 42321 47875
rect 42275 47803 42281 47837
rect 42315 47803 42321 47837
rect 42275 47765 42321 47803
rect 42275 47731 42281 47765
rect 42315 47731 42321 47765
rect 42275 47693 42321 47731
rect 42275 47659 42281 47693
rect 42315 47659 42321 47693
rect 42275 47621 42321 47659
rect 42275 47587 42281 47621
rect 42315 47587 42321 47621
rect 42275 47549 42321 47587
rect 42275 47515 42281 47549
rect 42315 47515 42321 47549
rect 42275 47477 42321 47515
rect 42275 47443 42281 47477
rect 42315 47443 42321 47477
rect 42275 47427 42321 47443
rect 42733 48701 42779 48717
rect 42733 48667 42739 48701
rect 42773 48667 42779 48701
rect 42733 48629 42779 48667
rect 42733 48595 42739 48629
rect 42773 48595 42779 48629
rect 42733 48557 42779 48595
rect 42733 48523 42739 48557
rect 42773 48523 42779 48557
rect 42733 48485 42779 48523
rect 42733 48451 42739 48485
rect 42773 48451 42779 48485
rect 42733 48413 42779 48451
rect 42733 48379 42739 48413
rect 42773 48379 42779 48413
rect 42733 48341 42779 48379
rect 42733 48307 42739 48341
rect 42773 48307 42779 48341
rect 42733 48269 42779 48307
rect 42733 48235 42739 48269
rect 42773 48235 42779 48269
rect 42733 48197 42779 48235
rect 42733 48163 42739 48197
rect 42773 48163 42779 48197
rect 42733 48125 42779 48163
rect 42733 48091 42739 48125
rect 42773 48091 42779 48125
rect 42733 48053 42779 48091
rect 42733 48019 42739 48053
rect 42773 48019 42779 48053
rect 42733 47981 42779 48019
rect 42733 47947 42739 47981
rect 42773 47947 42779 47981
rect 42733 47909 42779 47947
rect 42733 47875 42739 47909
rect 42773 47875 42779 47909
rect 42733 47837 42779 47875
rect 42733 47803 42739 47837
rect 42773 47803 42779 47837
rect 42733 47765 42779 47803
rect 42733 47731 42739 47765
rect 42773 47731 42779 47765
rect 42733 47693 42779 47731
rect 42733 47659 42739 47693
rect 42773 47659 42779 47693
rect 42733 47621 42779 47659
rect 42733 47587 42739 47621
rect 42773 47587 42779 47621
rect 42733 47549 42779 47587
rect 42733 47515 42739 47549
rect 42773 47515 42779 47549
rect 42733 47477 42779 47515
rect 42733 47443 42739 47477
rect 42773 47443 42779 47477
rect 42733 47427 42779 47443
rect 43191 48701 43237 48717
rect 43191 48667 43197 48701
rect 43231 48667 43237 48701
rect 43191 48629 43237 48667
rect 43191 48595 43197 48629
rect 43231 48595 43237 48629
rect 43191 48557 43237 48595
rect 43191 48523 43197 48557
rect 43231 48523 43237 48557
rect 43191 48485 43237 48523
rect 43191 48451 43197 48485
rect 43231 48451 43237 48485
rect 43191 48413 43237 48451
rect 43191 48379 43197 48413
rect 43231 48379 43237 48413
rect 43191 48341 43237 48379
rect 43191 48307 43197 48341
rect 43231 48307 43237 48341
rect 43191 48269 43237 48307
rect 43191 48235 43197 48269
rect 43231 48235 43237 48269
rect 43191 48197 43237 48235
rect 43191 48163 43197 48197
rect 43231 48163 43237 48197
rect 43191 48125 43237 48163
rect 43191 48091 43197 48125
rect 43231 48091 43237 48125
rect 43191 48053 43237 48091
rect 43191 48019 43197 48053
rect 43231 48019 43237 48053
rect 43191 47981 43237 48019
rect 43191 47947 43197 47981
rect 43231 47947 43237 47981
rect 43191 47909 43237 47947
rect 43191 47875 43197 47909
rect 43231 47875 43237 47909
rect 43191 47837 43237 47875
rect 43191 47803 43197 47837
rect 43231 47803 43237 47837
rect 43191 47765 43237 47803
rect 43191 47731 43197 47765
rect 43231 47731 43237 47765
rect 43191 47693 43237 47731
rect 43191 47659 43197 47693
rect 43231 47659 43237 47693
rect 43191 47621 43237 47659
rect 43191 47587 43197 47621
rect 43231 47587 43237 47621
rect 43191 47549 43237 47587
rect 43191 47515 43197 47549
rect 43231 47515 43237 47549
rect 43191 47477 43237 47515
rect 43191 47443 43197 47477
rect 43231 47443 43237 47477
rect 43191 47427 43237 47443
rect 43649 48701 43695 48717
rect 43649 48667 43655 48701
rect 43689 48667 43695 48701
rect 43649 48629 43695 48667
rect 43649 48595 43655 48629
rect 43689 48595 43695 48629
rect 43649 48557 43695 48595
rect 43649 48523 43655 48557
rect 43689 48523 43695 48557
rect 43649 48485 43695 48523
rect 43649 48451 43655 48485
rect 43689 48451 43695 48485
rect 43649 48413 43695 48451
rect 43649 48379 43655 48413
rect 43689 48379 43695 48413
rect 43649 48341 43695 48379
rect 43649 48307 43655 48341
rect 43689 48307 43695 48341
rect 43649 48269 43695 48307
rect 43649 48235 43655 48269
rect 43689 48235 43695 48269
rect 43649 48197 43695 48235
rect 43649 48163 43655 48197
rect 43689 48163 43695 48197
rect 43649 48125 43695 48163
rect 43649 48091 43655 48125
rect 43689 48091 43695 48125
rect 43649 48053 43695 48091
rect 43649 48019 43655 48053
rect 43689 48019 43695 48053
rect 43649 47981 43695 48019
rect 43649 47947 43655 47981
rect 43689 47947 43695 47981
rect 43649 47909 43695 47947
rect 43649 47875 43655 47909
rect 43689 47875 43695 47909
rect 43649 47837 43695 47875
rect 43649 47803 43655 47837
rect 43689 47803 43695 47837
rect 43649 47765 43695 47803
rect 43649 47731 43655 47765
rect 43689 47731 43695 47765
rect 43649 47693 43695 47731
rect 43649 47659 43655 47693
rect 43689 47659 43695 47693
rect 43649 47621 43695 47659
rect 43649 47587 43655 47621
rect 43689 47587 43695 47621
rect 43649 47549 43695 47587
rect 43649 47515 43655 47549
rect 43689 47515 43695 47549
rect 43649 47477 43695 47515
rect 43649 47443 43655 47477
rect 43689 47443 43695 47477
rect 43649 47427 43695 47443
rect 44107 48701 44153 48717
rect 44107 48667 44113 48701
rect 44147 48667 44153 48701
rect 44107 48629 44153 48667
rect 44107 48595 44113 48629
rect 44147 48595 44153 48629
rect 44107 48557 44153 48595
rect 44107 48523 44113 48557
rect 44147 48523 44153 48557
rect 44107 48485 44153 48523
rect 44107 48451 44113 48485
rect 44147 48451 44153 48485
rect 44107 48413 44153 48451
rect 44107 48379 44113 48413
rect 44147 48379 44153 48413
rect 44107 48341 44153 48379
rect 44107 48307 44113 48341
rect 44147 48307 44153 48341
rect 44107 48269 44153 48307
rect 44107 48235 44113 48269
rect 44147 48235 44153 48269
rect 44107 48197 44153 48235
rect 44107 48163 44113 48197
rect 44147 48163 44153 48197
rect 44107 48125 44153 48163
rect 44107 48091 44113 48125
rect 44147 48091 44153 48125
rect 44107 48053 44153 48091
rect 44107 48019 44113 48053
rect 44147 48019 44153 48053
rect 44107 47981 44153 48019
rect 44107 47947 44113 47981
rect 44147 47947 44153 47981
rect 44107 47909 44153 47947
rect 44107 47875 44113 47909
rect 44147 47875 44153 47909
rect 44107 47837 44153 47875
rect 44107 47803 44113 47837
rect 44147 47803 44153 47837
rect 44107 47765 44153 47803
rect 44107 47731 44113 47765
rect 44147 47731 44153 47765
rect 44107 47693 44153 47731
rect 44107 47659 44113 47693
rect 44147 47659 44153 47693
rect 44107 47621 44153 47659
rect 44107 47587 44113 47621
rect 44147 47587 44153 47621
rect 44107 47549 44153 47587
rect 44107 47515 44113 47549
rect 44147 47515 44153 47549
rect 44107 47477 44153 47515
rect 44107 47443 44113 47477
rect 44147 47443 44153 47477
rect 44107 47427 44153 47443
rect 44565 48701 44611 48717
rect 44565 48667 44571 48701
rect 44605 48667 44611 48701
rect 44565 48629 44611 48667
rect 44565 48595 44571 48629
rect 44605 48595 44611 48629
rect 44565 48557 44611 48595
rect 44565 48523 44571 48557
rect 44605 48523 44611 48557
rect 44565 48485 44611 48523
rect 44565 48451 44571 48485
rect 44605 48451 44611 48485
rect 44565 48413 44611 48451
rect 44565 48379 44571 48413
rect 44605 48379 44611 48413
rect 44565 48341 44611 48379
rect 44565 48307 44571 48341
rect 44605 48307 44611 48341
rect 44565 48269 44611 48307
rect 44565 48235 44571 48269
rect 44605 48235 44611 48269
rect 44565 48197 44611 48235
rect 44565 48163 44571 48197
rect 44605 48163 44611 48197
rect 44565 48125 44611 48163
rect 44565 48091 44571 48125
rect 44605 48091 44611 48125
rect 44565 48053 44611 48091
rect 44565 48019 44571 48053
rect 44605 48019 44611 48053
rect 44565 47981 44611 48019
rect 44565 47947 44571 47981
rect 44605 47947 44611 47981
rect 44565 47909 44611 47947
rect 44565 47875 44571 47909
rect 44605 47875 44611 47909
rect 44565 47837 44611 47875
rect 44565 47803 44571 47837
rect 44605 47803 44611 47837
rect 44565 47765 44611 47803
rect 44565 47731 44571 47765
rect 44605 47731 44611 47765
rect 44565 47693 44611 47731
rect 44565 47659 44571 47693
rect 44605 47659 44611 47693
rect 44565 47621 44611 47659
rect 44565 47587 44571 47621
rect 44605 47587 44611 47621
rect 44565 47549 44611 47587
rect 44565 47515 44571 47549
rect 44605 47515 44611 47549
rect 44565 47477 44611 47515
rect 44565 47443 44571 47477
rect 44605 47443 44611 47477
rect 44565 47427 44611 47443
rect 45023 48701 45069 48717
rect 45023 48667 45029 48701
rect 45063 48667 45069 48701
rect 45023 48629 45069 48667
rect 45023 48595 45029 48629
rect 45063 48595 45069 48629
rect 45023 48557 45069 48595
rect 45023 48523 45029 48557
rect 45063 48523 45069 48557
rect 45023 48485 45069 48523
rect 45023 48451 45029 48485
rect 45063 48451 45069 48485
rect 45023 48413 45069 48451
rect 45023 48379 45029 48413
rect 45063 48379 45069 48413
rect 45023 48341 45069 48379
rect 45023 48307 45029 48341
rect 45063 48307 45069 48341
rect 45023 48269 45069 48307
rect 45023 48235 45029 48269
rect 45063 48235 45069 48269
rect 45023 48197 45069 48235
rect 45023 48163 45029 48197
rect 45063 48163 45069 48197
rect 45023 48125 45069 48163
rect 45023 48091 45029 48125
rect 45063 48091 45069 48125
rect 45023 48053 45069 48091
rect 45023 48019 45029 48053
rect 45063 48019 45069 48053
rect 45023 47981 45069 48019
rect 45023 47947 45029 47981
rect 45063 47947 45069 47981
rect 45023 47909 45069 47947
rect 45023 47875 45029 47909
rect 45063 47875 45069 47909
rect 45023 47837 45069 47875
rect 45023 47803 45029 47837
rect 45063 47803 45069 47837
rect 45023 47765 45069 47803
rect 45023 47731 45029 47765
rect 45063 47731 45069 47765
rect 45023 47693 45069 47731
rect 45023 47659 45029 47693
rect 45063 47659 45069 47693
rect 45023 47621 45069 47659
rect 45023 47587 45029 47621
rect 45063 47587 45069 47621
rect 45023 47549 45069 47587
rect 45023 47515 45029 47549
rect 45063 47515 45069 47549
rect 45023 47477 45069 47515
rect 45023 47443 45029 47477
rect 45063 47443 45069 47477
rect 45023 47427 45069 47443
rect 45481 48701 45527 48717
rect 45481 48667 45487 48701
rect 45521 48667 45527 48701
rect 45481 48629 45527 48667
rect 45481 48595 45487 48629
rect 45521 48595 45527 48629
rect 45481 48557 45527 48595
rect 45481 48523 45487 48557
rect 45521 48523 45527 48557
rect 45481 48485 45527 48523
rect 45481 48451 45487 48485
rect 45521 48451 45527 48485
rect 45481 48413 45527 48451
rect 45481 48379 45487 48413
rect 45521 48379 45527 48413
rect 45481 48341 45527 48379
rect 45481 48307 45487 48341
rect 45521 48307 45527 48341
rect 45481 48269 45527 48307
rect 45481 48235 45487 48269
rect 45521 48235 45527 48269
rect 45481 48197 45527 48235
rect 45481 48163 45487 48197
rect 45521 48163 45527 48197
rect 45481 48125 45527 48163
rect 45481 48091 45487 48125
rect 45521 48091 45527 48125
rect 45481 48053 45527 48091
rect 45481 48019 45487 48053
rect 45521 48019 45527 48053
rect 45481 47981 45527 48019
rect 45481 47947 45487 47981
rect 45521 47947 45527 47981
rect 45481 47909 45527 47947
rect 45481 47875 45487 47909
rect 45521 47875 45527 47909
rect 45481 47837 45527 47875
rect 45481 47803 45487 47837
rect 45521 47803 45527 47837
rect 45481 47765 45527 47803
rect 45481 47731 45487 47765
rect 45521 47731 45527 47765
rect 45481 47693 45527 47731
rect 45481 47659 45487 47693
rect 45521 47659 45527 47693
rect 45481 47621 45527 47659
rect 45481 47587 45487 47621
rect 45521 47587 45527 47621
rect 45481 47549 45527 47587
rect 45481 47515 45487 47549
rect 45521 47515 45527 47549
rect 45481 47477 45527 47515
rect 45481 47443 45487 47477
rect 45521 47443 45527 47477
rect 45481 47427 45527 47443
rect 45939 48701 45985 48717
rect 45939 48667 45945 48701
rect 45979 48667 45985 48701
rect 45939 48629 45985 48667
rect 45939 48595 45945 48629
rect 45979 48595 45985 48629
rect 45939 48557 45985 48595
rect 45939 48523 45945 48557
rect 45979 48523 45985 48557
rect 45939 48485 45985 48523
rect 45939 48451 45945 48485
rect 45979 48451 45985 48485
rect 45939 48413 45985 48451
rect 45939 48379 45945 48413
rect 45979 48379 45985 48413
rect 45939 48341 45985 48379
rect 45939 48307 45945 48341
rect 45979 48307 45985 48341
rect 45939 48269 45985 48307
rect 45939 48235 45945 48269
rect 45979 48235 45985 48269
rect 45939 48197 45985 48235
rect 45939 48163 45945 48197
rect 45979 48163 45985 48197
rect 45939 48125 45985 48163
rect 45939 48091 45945 48125
rect 45979 48091 45985 48125
rect 45939 48053 45985 48091
rect 45939 48019 45945 48053
rect 45979 48019 45985 48053
rect 45939 47981 45985 48019
rect 45939 47947 45945 47981
rect 45979 47947 45985 47981
rect 45939 47909 45985 47947
rect 45939 47875 45945 47909
rect 45979 47875 45985 47909
rect 45939 47837 45985 47875
rect 45939 47803 45945 47837
rect 45979 47803 45985 47837
rect 45939 47765 45985 47803
rect 45939 47731 45945 47765
rect 45979 47731 45985 47765
rect 45939 47693 45985 47731
rect 45939 47659 45945 47693
rect 45979 47659 45985 47693
rect 45939 47621 45985 47659
rect 45939 47587 45945 47621
rect 45979 47587 45985 47621
rect 45939 47549 45985 47587
rect 45939 47515 45945 47549
rect 45979 47515 45985 47549
rect 45939 47477 45985 47515
rect 45939 47443 45945 47477
rect 45979 47443 45985 47477
rect 45939 47427 45985 47443
rect 46397 48701 46443 48717
rect 46397 48667 46403 48701
rect 46437 48667 46443 48701
rect 46397 48629 46443 48667
rect 46397 48595 46403 48629
rect 46437 48595 46443 48629
rect 46397 48557 46443 48595
rect 46397 48523 46403 48557
rect 46437 48523 46443 48557
rect 46397 48485 46443 48523
rect 46397 48451 46403 48485
rect 46437 48451 46443 48485
rect 46397 48413 46443 48451
rect 46397 48379 46403 48413
rect 46437 48379 46443 48413
rect 46397 48341 46443 48379
rect 46397 48307 46403 48341
rect 46437 48307 46443 48341
rect 46397 48269 46443 48307
rect 46397 48235 46403 48269
rect 46437 48235 46443 48269
rect 46397 48197 46443 48235
rect 46397 48163 46403 48197
rect 46437 48163 46443 48197
rect 46397 48125 46443 48163
rect 46397 48091 46403 48125
rect 46437 48091 46443 48125
rect 46397 48053 46443 48091
rect 46397 48019 46403 48053
rect 46437 48019 46443 48053
rect 46397 47981 46443 48019
rect 46397 47947 46403 47981
rect 46437 47947 46443 47981
rect 46397 47909 46443 47947
rect 46397 47875 46403 47909
rect 46437 47875 46443 47909
rect 46397 47837 46443 47875
rect 46397 47803 46403 47837
rect 46437 47803 46443 47837
rect 46397 47765 46443 47803
rect 46397 47731 46403 47765
rect 46437 47731 46443 47765
rect 46397 47693 46443 47731
rect 46397 47659 46403 47693
rect 46437 47659 46443 47693
rect 46397 47621 46443 47659
rect 46397 47587 46403 47621
rect 46437 47587 46443 47621
rect 46397 47549 46443 47587
rect 46397 47515 46403 47549
rect 46437 47515 46443 47549
rect 46397 47477 46443 47515
rect 46397 47443 46403 47477
rect 46437 47443 46443 47477
rect 46397 47427 46443 47443
rect 46855 48701 46901 48717
rect 46855 48667 46861 48701
rect 46895 48667 46901 48701
rect 46855 48629 46901 48667
rect 46855 48595 46861 48629
rect 46895 48595 46901 48629
rect 46855 48557 46901 48595
rect 46855 48523 46861 48557
rect 46895 48523 46901 48557
rect 46855 48485 46901 48523
rect 46855 48451 46861 48485
rect 46895 48451 46901 48485
rect 46855 48413 46901 48451
rect 46855 48379 46861 48413
rect 46895 48379 46901 48413
rect 46855 48341 46901 48379
rect 46855 48307 46861 48341
rect 46895 48307 46901 48341
rect 46855 48269 46901 48307
rect 46855 48235 46861 48269
rect 46895 48235 46901 48269
rect 46855 48197 46901 48235
rect 46855 48163 46861 48197
rect 46895 48163 46901 48197
rect 46855 48125 46901 48163
rect 46855 48091 46861 48125
rect 46895 48091 46901 48125
rect 46855 48053 46901 48091
rect 46855 48019 46861 48053
rect 46895 48019 46901 48053
rect 46855 47981 46901 48019
rect 46855 47947 46861 47981
rect 46895 47947 46901 47981
rect 46855 47909 46901 47947
rect 46855 47875 46861 47909
rect 46895 47875 46901 47909
rect 46855 47837 46901 47875
rect 46855 47803 46861 47837
rect 46895 47803 46901 47837
rect 46855 47765 46901 47803
rect 46855 47731 46861 47765
rect 46895 47731 46901 47765
rect 46855 47693 46901 47731
rect 46855 47659 46861 47693
rect 46895 47659 46901 47693
rect 46855 47621 46901 47659
rect 46855 47587 46861 47621
rect 46895 47587 46901 47621
rect 46855 47549 46901 47587
rect 46855 47515 46861 47549
rect 46895 47515 46901 47549
rect 46855 47477 46901 47515
rect 46855 47443 46861 47477
rect 46895 47443 46901 47477
rect 46855 47427 46901 47443
rect 47313 48701 47359 48717
rect 47313 48667 47319 48701
rect 47353 48667 47359 48701
rect 47313 48629 47359 48667
rect 47313 48595 47319 48629
rect 47353 48595 47359 48629
rect 47313 48557 47359 48595
rect 47313 48523 47319 48557
rect 47353 48523 47359 48557
rect 47313 48485 47359 48523
rect 47313 48451 47319 48485
rect 47353 48451 47359 48485
rect 47313 48413 47359 48451
rect 47313 48379 47319 48413
rect 47353 48379 47359 48413
rect 47313 48341 47359 48379
rect 47313 48307 47319 48341
rect 47353 48307 47359 48341
rect 47313 48269 47359 48307
rect 47313 48235 47319 48269
rect 47353 48235 47359 48269
rect 47313 48197 47359 48235
rect 47313 48163 47319 48197
rect 47353 48163 47359 48197
rect 47313 48125 47359 48163
rect 47313 48091 47319 48125
rect 47353 48091 47359 48125
rect 47313 48053 47359 48091
rect 47313 48019 47319 48053
rect 47353 48019 47359 48053
rect 47313 47981 47359 48019
rect 47313 47947 47319 47981
rect 47353 47947 47359 47981
rect 47313 47909 47359 47947
rect 47313 47875 47319 47909
rect 47353 47875 47359 47909
rect 47313 47837 47359 47875
rect 47313 47803 47319 47837
rect 47353 47803 47359 47837
rect 47313 47765 47359 47803
rect 47313 47731 47319 47765
rect 47353 47731 47359 47765
rect 47313 47693 47359 47731
rect 47313 47659 47319 47693
rect 47353 47659 47359 47693
rect 47313 47621 47359 47659
rect 47313 47587 47319 47621
rect 47353 47587 47359 47621
rect 47313 47549 47359 47587
rect 47313 47515 47319 47549
rect 47353 47515 47359 47549
rect 47313 47477 47359 47515
rect 47313 47443 47319 47477
rect 47353 47443 47359 47477
rect 47313 47427 47359 47443
rect 47771 48701 47817 48717
rect 47771 48667 47777 48701
rect 47811 48667 47817 48701
rect 47771 48629 47817 48667
rect 47771 48595 47777 48629
rect 47811 48595 47817 48629
rect 47771 48557 47817 48595
rect 47771 48523 47777 48557
rect 47811 48523 47817 48557
rect 47771 48485 47817 48523
rect 47771 48451 47777 48485
rect 47811 48451 47817 48485
rect 47771 48413 47817 48451
rect 47771 48379 47777 48413
rect 47811 48379 47817 48413
rect 47771 48341 47817 48379
rect 47771 48307 47777 48341
rect 47811 48307 47817 48341
rect 47771 48269 47817 48307
rect 47771 48235 47777 48269
rect 47811 48235 47817 48269
rect 47771 48197 47817 48235
rect 47771 48163 47777 48197
rect 47811 48163 47817 48197
rect 47771 48125 47817 48163
rect 47771 48091 47777 48125
rect 47811 48091 47817 48125
rect 47771 48053 47817 48091
rect 47771 48019 47777 48053
rect 47811 48019 47817 48053
rect 47771 47981 47817 48019
rect 47771 47947 47777 47981
rect 47811 47947 47817 47981
rect 47771 47909 47817 47947
rect 47771 47875 47777 47909
rect 47811 47875 47817 47909
rect 47771 47837 47817 47875
rect 47771 47803 47777 47837
rect 47811 47803 47817 47837
rect 47771 47765 47817 47803
rect 47771 47731 47777 47765
rect 47811 47731 47817 47765
rect 47771 47693 47817 47731
rect 47771 47659 47777 47693
rect 47811 47659 47817 47693
rect 47771 47621 47817 47659
rect 47771 47587 47777 47621
rect 47811 47587 47817 47621
rect 47771 47549 47817 47587
rect 47771 47515 47777 47549
rect 47811 47515 47817 47549
rect 47771 47477 47817 47515
rect 47771 47443 47777 47477
rect 47811 47443 47817 47477
rect 47771 47427 47817 47443
rect 48229 48701 48275 48717
rect 48229 48667 48235 48701
rect 48269 48667 48275 48701
rect 48229 48629 48275 48667
rect 48229 48595 48235 48629
rect 48269 48595 48275 48629
rect 48229 48557 48275 48595
rect 48229 48523 48235 48557
rect 48269 48523 48275 48557
rect 48229 48485 48275 48523
rect 48229 48451 48235 48485
rect 48269 48451 48275 48485
rect 48229 48413 48275 48451
rect 48229 48379 48235 48413
rect 48269 48379 48275 48413
rect 48229 48341 48275 48379
rect 48229 48307 48235 48341
rect 48269 48307 48275 48341
rect 48229 48269 48275 48307
rect 48229 48235 48235 48269
rect 48269 48235 48275 48269
rect 48229 48197 48275 48235
rect 48229 48163 48235 48197
rect 48269 48163 48275 48197
rect 48229 48125 48275 48163
rect 48229 48091 48235 48125
rect 48269 48091 48275 48125
rect 48229 48053 48275 48091
rect 48229 48019 48235 48053
rect 48269 48019 48275 48053
rect 48229 47981 48275 48019
rect 48229 47947 48235 47981
rect 48269 47947 48275 47981
rect 48229 47909 48275 47947
rect 48229 47875 48235 47909
rect 48269 47875 48275 47909
rect 48229 47837 48275 47875
rect 48229 47803 48235 47837
rect 48269 47803 48275 47837
rect 48229 47765 48275 47803
rect 48229 47731 48235 47765
rect 48269 47731 48275 47765
rect 48229 47693 48275 47731
rect 48229 47659 48235 47693
rect 48269 47659 48275 47693
rect 48229 47621 48275 47659
rect 48229 47587 48235 47621
rect 48269 47587 48275 47621
rect 48229 47549 48275 47587
rect 48229 47515 48235 47549
rect 48269 47515 48275 47549
rect 48687 48701 48733 48717
rect 48687 48667 48693 48701
rect 48727 48667 48733 48701
rect 48687 48629 48733 48667
rect 48687 48595 48693 48629
rect 48727 48595 48733 48629
rect 48687 48557 48733 48595
rect 48687 48523 48693 48557
rect 48727 48523 48733 48557
rect 48687 48485 48733 48523
rect 48687 48451 48693 48485
rect 48727 48451 48733 48485
rect 48687 48413 48733 48451
rect 48687 48379 48693 48413
rect 48727 48379 48733 48413
rect 48687 48341 48733 48379
rect 48687 48307 48693 48341
rect 48727 48307 48733 48341
rect 48687 48269 48733 48307
rect 48687 48235 48693 48269
rect 48727 48235 48733 48269
rect 48687 48197 48733 48235
rect 48687 48163 48693 48197
rect 48727 48163 48733 48197
rect 48687 48125 48733 48163
rect 48687 48091 48693 48125
rect 48727 48091 48733 48125
rect 48687 48053 48733 48091
rect 48687 48019 48693 48053
rect 48727 48019 48733 48053
rect 48687 47981 48733 48019
rect 48687 47947 48693 47981
rect 48727 47947 48733 47981
rect 48687 47909 48733 47947
rect 48687 47875 48693 47909
rect 48727 47875 48733 47909
rect 48687 47837 48733 47875
rect 48687 47803 48693 47837
rect 48727 47803 48733 47837
rect 48687 47765 48733 47803
rect 48687 47731 48693 47765
rect 48727 47731 48733 47765
rect 48687 47693 48733 47731
rect 48687 47659 48693 47693
rect 48727 47659 48733 47693
rect 48687 47621 48733 47659
rect 48687 47587 48693 47621
rect 48727 47587 48733 47621
rect 48687 47549 48733 47587
rect 48229 47477 48275 47515
rect 48229 47443 48235 47477
rect 48269 47443 48275 47477
rect 48314 47472 48320 47524
rect 48372 47512 48378 47524
rect 48687 47515 48693 47549
rect 48727 47515 48733 47549
rect 48687 47512 48733 47515
rect 48372 47484 48733 47512
rect 48372 47472 48378 47484
rect 48687 47477 48733 47484
rect 48229 47427 48275 47443
rect 48687 47443 48693 47477
rect 48727 47443 48733 47477
rect 48687 47427 48733 47443
rect 49145 48701 49191 48717
rect 49145 48667 49151 48701
rect 49185 48667 49191 48701
rect 49145 48629 49191 48667
rect 49145 48595 49151 48629
rect 49185 48595 49191 48629
rect 49145 48557 49191 48595
rect 49145 48523 49151 48557
rect 49185 48523 49191 48557
rect 49145 48485 49191 48523
rect 49145 48451 49151 48485
rect 49185 48451 49191 48485
rect 49145 48413 49191 48451
rect 49145 48379 49151 48413
rect 49185 48379 49191 48413
rect 49145 48341 49191 48379
rect 49145 48307 49151 48341
rect 49185 48307 49191 48341
rect 49145 48269 49191 48307
rect 49145 48235 49151 48269
rect 49185 48235 49191 48269
rect 49145 48197 49191 48235
rect 49145 48163 49151 48197
rect 49185 48163 49191 48197
rect 49145 48125 49191 48163
rect 49145 48091 49151 48125
rect 49185 48091 49191 48125
rect 49145 48053 49191 48091
rect 49145 48019 49151 48053
rect 49185 48019 49191 48053
rect 49145 47981 49191 48019
rect 49145 47947 49151 47981
rect 49185 47947 49191 47981
rect 49145 47909 49191 47947
rect 49145 47875 49151 47909
rect 49185 47875 49191 47909
rect 49145 47837 49191 47875
rect 49145 47803 49151 47837
rect 49185 47803 49191 47837
rect 49145 47765 49191 47803
rect 49145 47731 49151 47765
rect 49185 47731 49191 47765
rect 49145 47693 49191 47731
rect 49145 47659 49151 47693
rect 49185 47659 49191 47693
rect 49145 47621 49191 47659
rect 49145 47587 49151 47621
rect 49185 47587 49191 47621
rect 49145 47549 49191 47587
rect 49145 47515 49151 47549
rect 49185 47515 49191 47549
rect 49145 47477 49191 47515
rect 49145 47443 49151 47477
rect 49185 47443 49191 47477
rect 49145 47427 49191 47443
rect 49603 48701 49649 48717
rect 49603 48667 49609 48701
rect 49643 48667 49649 48701
rect 49603 48629 49649 48667
rect 49603 48595 49609 48629
rect 49643 48595 49649 48629
rect 49603 48557 49649 48595
rect 49603 48523 49609 48557
rect 49643 48523 49649 48557
rect 49603 48485 49649 48523
rect 49603 48451 49609 48485
rect 49643 48451 49649 48485
rect 49603 48413 49649 48451
rect 49603 48379 49609 48413
rect 49643 48379 49649 48413
rect 49603 48341 49649 48379
rect 49603 48307 49609 48341
rect 49643 48307 49649 48341
rect 49603 48269 49649 48307
rect 49603 48235 49609 48269
rect 49643 48235 49649 48269
rect 49603 48197 49649 48235
rect 49603 48163 49609 48197
rect 49643 48163 49649 48197
rect 49603 48125 49649 48163
rect 49603 48091 49609 48125
rect 49643 48091 49649 48125
rect 49603 48053 49649 48091
rect 49603 48019 49609 48053
rect 49643 48019 49649 48053
rect 49603 47981 49649 48019
rect 49603 47947 49609 47981
rect 49643 47947 49649 47981
rect 49603 47909 49649 47947
rect 49603 47875 49609 47909
rect 49643 47875 49649 47909
rect 49603 47837 49649 47875
rect 49603 47803 49609 47837
rect 49643 47803 49649 47837
rect 49603 47765 49649 47803
rect 49603 47731 49609 47765
rect 49643 47731 49649 47765
rect 49603 47693 49649 47731
rect 49603 47659 49609 47693
rect 49643 47659 49649 47693
rect 49603 47621 49649 47659
rect 49603 47587 49609 47621
rect 49643 47587 49649 47621
rect 49603 47549 49649 47587
rect 49603 47515 49609 47549
rect 49643 47515 49649 47549
rect 49603 47477 49649 47515
rect 49603 47443 49609 47477
rect 49643 47443 49649 47477
rect 49603 47427 49649 47443
rect 50061 48701 50107 48717
rect 50061 48667 50067 48701
rect 50101 48667 50107 48701
rect 50061 48629 50107 48667
rect 50061 48595 50067 48629
rect 50101 48595 50107 48629
rect 50061 48557 50107 48595
rect 50061 48523 50067 48557
rect 50101 48523 50107 48557
rect 50061 48485 50107 48523
rect 50061 48451 50067 48485
rect 50101 48451 50107 48485
rect 50061 48413 50107 48451
rect 50061 48379 50067 48413
rect 50101 48379 50107 48413
rect 50061 48341 50107 48379
rect 50061 48307 50067 48341
rect 50101 48307 50107 48341
rect 50061 48269 50107 48307
rect 50061 48235 50067 48269
rect 50101 48235 50107 48269
rect 50061 48197 50107 48235
rect 50061 48163 50067 48197
rect 50101 48163 50107 48197
rect 50061 48125 50107 48163
rect 50061 48091 50067 48125
rect 50101 48091 50107 48125
rect 50061 48053 50107 48091
rect 50061 48019 50067 48053
rect 50101 48019 50107 48053
rect 50061 47981 50107 48019
rect 50061 47947 50067 47981
rect 50101 47947 50107 47981
rect 50061 47909 50107 47947
rect 50061 47875 50067 47909
rect 50101 47875 50107 47909
rect 50061 47837 50107 47875
rect 50061 47803 50067 47837
rect 50101 47803 50107 47837
rect 50061 47765 50107 47803
rect 50061 47731 50067 47765
rect 50101 47731 50107 47765
rect 50061 47693 50107 47731
rect 50061 47659 50067 47693
rect 50101 47659 50107 47693
rect 50061 47621 50107 47659
rect 50061 47587 50067 47621
rect 50101 47587 50107 47621
rect 50061 47549 50107 47587
rect 50061 47515 50067 47549
rect 50101 47515 50107 47549
rect 50061 47477 50107 47515
rect 50061 47443 50067 47477
rect 50101 47443 50107 47477
rect 50061 47427 50107 47443
rect 50519 48701 50565 48717
rect 50519 48667 50525 48701
rect 50559 48667 50565 48701
rect 50519 48629 50565 48667
rect 50519 48595 50525 48629
rect 50559 48595 50565 48629
rect 50519 48557 50565 48595
rect 50519 48523 50525 48557
rect 50559 48523 50565 48557
rect 50519 48485 50565 48523
rect 50519 48451 50525 48485
rect 50559 48451 50565 48485
rect 50519 48413 50565 48451
rect 50519 48379 50525 48413
rect 50559 48379 50565 48413
rect 50519 48341 50565 48379
rect 50519 48307 50525 48341
rect 50559 48307 50565 48341
rect 50519 48269 50565 48307
rect 50519 48235 50525 48269
rect 50559 48235 50565 48269
rect 50519 48197 50565 48235
rect 50519 48163 50525 48197
rect 50559 48163 50565 48197
rect 50519 48125 50565 48163
rect 50519 48091 50525 48125
rect 50559 48091 50565 48125
rect 50519 48053 50565 48091
rect 50519 48019 50525 48053
rect 50559 48019 50565 48053
rect 50519 47981 50565 48019
rect 50519 47947 50525 47981
rect 50559 47947 50565 47981
rect 50519 47909 50565 47947
rect 50519 47875 50525 47909
rect 50559 47875 50565 47909
rect 50519 47837 50565 47875
rect 50519 47803 50525 47837
rect 50559 47803 50565 47837
rect 50519 47765 50565 47803
rect 50519 47731 50525 47765
rect 50559 47731 50565 47765
rect 50519 47693 50565 47731
rect 50519 47659 50525 47693
rect 50559 47659 50565 47693
rect 50519 47621 50565 47659
rect 50519 47587 50525 47621
rect 50559 47587 50565 47621
rect 50519 47549 50565 47587
rect 50519 47515 50525 47549
rect 50559 47515 50565 47549
rect 50519 47477 50565 47515
rect 50519 47443 50525 47477
rect 50559 47443 50565 47477
rect 50519 47427 50565 47443
rect 50977 48701 51023 48717
rect 50977 48667 50983 48701
rect 51017 48667 51023 48701
rect 50977 48629 51023 48667
rect 50977 48595 50983 48629
rect 51017 48595 51023 48629
rect 50977 48557 51023 48595
rect 50977 48523 50983 48557
rect 51017 48523 51023 48557
rect 50977 48485 51023 48523
rect 50977 48451 50983 48485
rect 51017 48451 51023 48485
rect 50977 48413 51023 48451
rect 50977 48379 50983 48413
rect 51017 48379 51023 48413
rect 50977 48341 51023 48379
rect 50977 48307 50983 48341
rect 51017 48307 51023 48341
rect 50977 48269 51023 48307
rect 50977 48235 50983 48269
rect 51017 48235 51023 48269
rect 50977 48197 51023 48235
rect 50977 48163 50983 48197
rect 51017 48163 51023 48197
rect 50977 48125 51023 48163
rect 50977 48091 50983 48125
rect 51017 48091 51023 48125
rect 50977 48053 51023 48091
rect 50977 48019 50983 48053
rect 51017 48019 51023 48053
rect 50977 47981 51023 48019
rect 50977 47947 50983 47981
rect 51017 47947 51023 47981
rect 50977 47909 51023 47947
rect 50977 47875 50983 47909
rect 51017 47875 51023 47909
rect 50977 47837 51023 47875
rect 50977 47803 50983 47837
rect 51017 47803 51023 47837
rect 50977 47765 51023 47803
rect 50977 47731 50983 47765
rect 51017 47731 51023 47765
rect 50977 47693 51023 47731
rect 50977 47659 50983 47693
rect 51017 47659 51023 47693
rect 50977 47621 51023 47659
rect 50977 47587 50983 47621
rect 51017 47587 51023 47621
rect 50977 47549 51023 47587
rect 50977 47515 50983 47549
rect 51017 47515 51023 47549
rect 50977 47477 51023 47515
rect 50977 47443 50983 47477
rect 51017 47443 51023 47477
rect 50977 47427 51023 47443
rect 51435 48701 51481 48717
rect 51435 48667 51441 48701
rect 51475 48667 51481 48701
rect 51435 48629 51481 48667
rect 51435 48595 51441 48629
rect 51475 48595 51481 48629
rect 51435 48557 51481 48595
rect 51435 48523 51441 48557
rect 51475 48523 51481 48557
rect 51435 48485 51481 48523
rect 51435 48451 51441 48485
rect 51475 48451 51481 48485
rect 51435 48413 51481 48451
rect 51435 48379 51441 48413
rect 51475 48379 51481 48413
rect 51435 48341 51481 48379
rect 51435 48307 51441 48341
rect 51475 48307 51481 48341
rect 51435 48269 51481 48307
rect 51435 48235 51441 48269
rect 51475 48235 51481 48269
rect 51435 48197 51481 48235
rect 51435 48163 51441 48197
rect 51475 48163 51481 48197
rect 51435 48125 51481 48163
rect 51435 48091 51441 48125
rect 51475 48091 51481 48125
rect 51435 48053 51481 48091
rect 51435 48019 51441 48053
rect 51475 48019 51481 48053
rect 51435 47981 51481 48019
rect 51435 47947 51441 47981
rect 51475 47947 51481 47981
rect 51435 47909 51481 47947
rect 51435 47875 51441 47909
rect 51475 47875 51481 47909
rect 51435 47837 51481 47875
rect 51435 47803 51441 47837
rect 51475 47803 51481 47837
rect 51435 47765 51481 47803
rect 51435 47731 51441 47765
rect 51475 47731 51481 47765
rect 51435 47693 51481 47731
rect 51435 47659 51441 47693
rect 51475 47659 51481 47693
rect 51435 47621 51481 47659
rect 51435 47587 51441 47621
rect 51475 47587 51481 47621
rect 51435 47549 51481 47587
rect 51435 47515 51441 47549
rect 51475 47515 51481 47549
rect 51435 47477 51481 47515
rect 51435 47443 51441 47477
rect 51475 47443 51481 47477
rect 51435 47427 51481 47443
rect 51893 48701 51939 48717
rect 51893 48667 51899 48701
rect 51933 48667 51939 48701
rect 51893 48629 51939 48667
rect 51893 48595 51899 48629
rect 51933 48595 51939 48629
rect 51893 48557 51939 48595
rect 51893 48523 51899 48557
rect 51933 48523 51939 48557
rect 51893 48485 51939 48523
rect 51893 48451 51899 48485
rect 51933 48451 51939 48485
rect 51893 48413 51939 48451
rect 51893 48379 51899 48413
rect 51933 48379 51939 48413
rect 51893 48341 51939 48379
rect 51893 48307 51899 48341
rect 51933 48307 51939 48341
rect 51893 48269 51939 48307
rect 51893 48235 51899 48269
rect 51933 48235 51939 48269
rect 51893 48197 51939 48235
rect 51893 48163 51899 48197
rect 51933 48163 51939 48197
rect 51893 48125 51939 48163
rect 51893 48091 51899 48125
rect 51933 48091 51939 48125
rect 51893 48053 51939 48091
rect 51893 48019 51899 48053
rect 51933 48019 51939 48053
rect 51893 47981 51939 48019
rect 51893 47947 51899 47981
rect 51933 47947 51939 47981
rect 51893 47909 51939 47947
rect 51893 47875 51899 47909
rect 51933 47875 51939 47909
rect 51893 47837 51939 47875
rect 51893 47803 51899 47837
rect 51933 47803 51939 47837
rect 51893 47765 51939 47803
rect 51893 47731 51899 47765
rect 51933 47731 51939 47765
rect 51893 47693 51939 47731
rect 51893 47659 51899 47693
rect 51933 47659 51939 47693
rect 51893 47621 51939 47659
rect 51893 47587 51899 47621
rect 51933 47587 51939 47621
rect 51893 47549 51939 47587
rect 51893 47515 51899 47549
rect 51933 47515 51939 47549
rect 51893 47477 51939 47515
rect 51893 47443 51899 47477
rect 51933 47443 51939 47477
rect 51893 47427 51939 47443
rect 52351 48701 52397 48717
rect 52351 48667 52357 48701
rect 52391 48667 52397 48701
rect 52351 48629 52397 48667
rect 52351 48595 52357 48629
rect 52391 48595 52397 48629
rect 52351 48557 52397 48595
rect 52351 48523 52357 48557
rect 52391 48523 52397 48557
rect 52351 48485 52397 48523
rect 52351 48451 52357 48485
rect 52391 48451 52397 48485
rect 52351 48413 52397 48451
rect 52351 48379 52357 48413
rect 52391 48379 52397 48413
rect 52351 48341 52397 48379
rect 52351 48307 52357 48341
rect 52391 48307 52397 48341
rect 52351 48269 52397 48307
rect 52351 48235 52357 48269
rect 52391 48235 52397 48269
rect 52351 48197 52397 48235
rect 52351 48163 52357 48197
rect 52391 48163 52397 48197
rect 52351 48125 52397 48163
rect 52351 48091 52357 48125
rect 52391 48091 52397 48125
rect 52351 48053 52397 48091
rect 52351 48019 52357 48053
rect 52391 48019 52397 48053
rect 52351 47981 52397 48019
rect 52351 47947 52357 47981
rect 52391 47947 52397 47981
rect 52351 47909 52397 47947
rect 52351 47875 52357 47909
rect 52391 47875 52397 47909
rect 52351 47837 52397 47875
rect 52351 47803 52357 47837
rect 52391 47803 52397 47837
rect 52351 47765 52397 47803
rect 52351 47731 52357 47765
rect 52391 47731 52397 47765
rect 52351 47693 52397 47731
rect 52351 47659 52357 47693
rect 52391 47659 52397 47693
rect 52351 47621 52397 47659
rect 52351 47587 52357 47621
rect 52391 47587 52397 47621
rect 52351 47549 52397 47587
rect 52351 47515 52357 47549
rect 52391 47515 52397 47549
rect 52351 47477 52397 47515
rect 52351 47443 52357 47477
rect 52391 47443 52397 47477
rect 52351 47427 52397 47443
rect 29454 47240 29460 47252
rect 29399 47212 29460 47240
rect 29454 47200 29460 47212
rect 29512 47200 29518 47252
rect 900 47130 57536 47132
rect 900 47014 922 47130
rect 2510 47116 55926 47130
rect 2510 47089 17684 47116
rect 2510 47055 6101 47089
rect 6135 47055 6501 47089
rect 6535 47055 6901 47089
rect 6935 47055 7301 47089
rect 7335 47055 7701 47089
rect 7735 47055 8101 47089
rect 8135 47055 8501 47089
rect 8535 47055 8901 47089
rect 8935 47055 9301 47089
rect 9335 47055 9701 47089
rect 9735 47055 10101 47089
rect 10135 47055 10501 47089
rect 10535 47055 10901 47089
rect 10935 47055 11301 47089
rect 11335 47055 11701 47089
rect 11735 47055 12101 47089
rect 12135 47055 12501 47089
rect 12535 47055 12901 47089
rect 12935 47055 13549 47089
rect 13583 47055 13949 47089
rect 13983 47055 14349 47089
rect 14383 47055 14749 47089
rect 14783 47055 15149 47089
rect 15183 47055 15549 47089
rect 15583 47055 15949 47089
rect 15983 47055 16349 47089
rect 16383 47055 16749 47089
rect 16783 47055 17149 47089
rect 17183 47055 17549 47089
rect 17583 47064 17684 47089
rect 17736 47089 55926 47116
rect 17736 47064 17949 47089
rect 17583 47055 17949 47064
rect 17983 47055 18349 47089
rect 18383 47055 18749 47089
rect 18783 47055 19149 47089
rect 19183 47055 19549 47089
rect 19583 47055 19949 47089
rect 19983 47055 20349 47089
rect 20383 47055 21015 47089
rect 21049 47055 21215 47089
rect 21249 47055 21415 47089
rect 21449 47055 21615 47089
rect 21649 47055 21815 47089
rect 21849 47055 22015 47089
rect 22049 47055 22215 47089
rect 22249 47055 22415 47089
rect 22449 47055 22615 47089
rect 22649 47055 22815 47089
rect 22849 47055 23015 47089
rect 23049 47055 24101 47089
rect 24135 47055 25013 47089
rect 25047 47055 25413 47089
rect 25447 47055 25813 47089
rect 25847 47055 26213 47089
rect 26247 47055 26613 47089
rect 26647 47055 27013 47089
rect 27047 47055 27413 47089
rect 27447 47055 27813 47089
rect 27847 47055 28213 47089
rect 28247 47055 28613 47089
rect 28647 47055 29013 47089
rect 29047 47055 29413 47089
rect 29447 47055 29813 47089
rect 29847 47055 30213 47089
rect 30247 47055 30613 47089
rect 30647 47055 31013 47089
rect 31047 47055 31413 47089
rect 31447 47055 31813 47089
rect 31847 47055 32213 47089
rect 32247 47055 32613 47089
rect 32647 47055 33013 47089
rect 33047 47055 33413 47089
rect 33447 47055 33813 47089
rect 33847 47055 34213 47089
rect 34247 47055 34613 47089
rect 34647 47055 35013 47089
rect 35047 47055 35413 47089
rect 35447 47055 35813 47089
rect 35847 47055 36213 47089
rect 36247 47055 36613 47089
rect 36647 47055 37013 47089
rect 37047 47055 37413 47089
rect 37447 47055 37813 47089
rect 37847 47055 38213 47089
rect 38247 47055 38613 47089
rect 38647 47055 39013 47089
rect 39047 47055 39413 47089
rect 39447 47055 39813 47089
rect 39847 47055 40213 47089
rect 40247 47055 40613 47089
rect 40647 47055 41013 47089
rect 41047 47055 41413 47089
rect 41447 47055 41813 47089
rect 41847 47055 42213 47089
rect 42247 47055 42613 47089
rect 42647 47055 43013 47089
rect 43047 47055 43413 47089
rect 43447 47055 43813 47089
rect 43847 47055 44213 47089
rect 44247 47055 44613 47089
rect 44647 47055 45013 47089
rect 45047 47055 45413 47089
rect 45447 47055 45813 47089
rect 45847 47055 46213 47089
rect 46247 47055 46613 47089
rect 46647 47055 47013 47089
rect 47047 47055 47413 47089
rect 47447 47055 47813 47089
rect 47847 47055 48213 47089
rect 48247 47055 48613 47089
rect 48647 47055 49013 47089
rect 49047 47055 49413 47089
rect 49447 47055 49813 47089
rect 49847 47055 50213 47089
rect 50247 47055 50613 47089
rect 50647 47055 51013 47089
rect 51047 47055 51413 47089
rect 51447 47055 51813 47089
rect 51847 47055 52213 47089
rect 52247 47055 55926 47089
rect 2510 47014 55926 47055
rect 57514 47014 57536 47130
rect 900 47012 57536 47014
rect 3348 45250 55088 45252
rect 3348 45134 3370 45250
rect 4958 45209 53478 45250
rect 4958 45175 6101 45209
rect 6135 45175 6501 45209
rect 6535 45175 6901 45209
rect 6935 45175 7301 45209
rect 7335 45175 7701 45209
rect 7735 45175 8101 45209
rect 8135 45175 8501 45209
rect 8535 45175 8901 45209
rect 8935 45175 9301 45209
rect 9335 45175 9701 45209
rect 9735 45175 10101 45209
rect 10135 45175 10501 45209
rect 10535 45175 10901 45209
rect 10935 45175 11301 45209
rect 11335 45175 11701 45209
rect 11735 45175 12101 45209
rect 12135 45175 12501 45209
rect 12535 45175 12901 45209
rect 12935 45175 14301 45209
rect 14335 45175 15213 45209
rect 15247 45175 15613 45209
rect 15647 45175 16013 45209
rect 16047 45175 16413 45209
rect 16447 45175 16813 45209
rect 16847 45175 17213 45209
rect 17247 45175 17613 45209
rect 17647 45175 18013 45209
rect 18047 45175 18413 45209
rect 18447 45175 18813 45209
rect 18847 45175 19213 45209
rect 19247 45175 19613 45209
rect 19647 45175 20013 45209
rect 20047 45175 20413 45209
rect 20447 45175 20813 45209
rect 20847 45175 21213 45209
rect 21247 45175 21613 45209
rect 21647 45175 22013 45209
rect 22047 45175 22413 45209
rect 22447 45175 22813 45209
rect 22847 45175 23213 45209
rect 23247 45175 23613 45209
rect 23647 45175 24013 45209
rect 24047 45175 24413 45209
rect 24447 45175 24813 45209
rect 24847 45175 25213 45209
rect 25247 45175 25613 45209
rect 25647 45175 26013 45209
rect 26047 45175 26413 45209
rect 26447 45175 26813 45209
rect 26847 45175 27213 45209
rect 27247 45175 27613 45209
rect 27647 45175 28013 45209
rect 28047 45175 28413 45209
rect 28447 45175 28813 45209
rect 28847 45175 29213 45209
rect 29247 45175 29613 45209
rect 29647 45175 30013 45209
rect 30047 45175 30413 45209
rect 30447 45175 30813 45209
rect 30847 45175 31213 45209
rect 31247 45175 31613 45209
rect 31647 45175 32013 45209
rect 32047 45175 32413 45209
rect 32447 45175 32813 45209
rect 32847 45175 33213 45209
rect 33247 45175 33613 45209
rect 33647 45175 34013 45209
rect 34047 45175 34413 45209
rect 34447 45175 34813 45209
rect 34847 45175 35213 45209
rect 35247 45175 35613 45209
rect 35647 45175 36013 45209
rect 36047 45175 36413 45209
rect 36447 45175 36813 45209
rect 36847 45175 37213 45209
rect 37247 45175 37613 45209
rect 37647 45175 38013 45209
rect 38047 45175 38413 45209
rect 38447 45175 38813 45209
rect 38847 45175 39213 45209
rect 39247 45175 39613 45209
rect 39647 45175 40013 45209
rect 40047 45175 40413 45209
rect 40447 45175 40813 45209
rect 40847 45175 41213 45209
rect 41247 45175 41613 45209
rect 41647 45175 42013 45209
rect 42047 45175 42413 45209
rect 42447 45175 43143 45209
rect 43177 45175 43343 45209
rect 43377 45175 43543 45209
rect 43577 45175 43743 45209
rect 43777 45175 43943 45209
rect 43977 45175 44143 45209
rect 44177 45175 44343 45209
rect 44377 45175 44543 45209
rect 44577 45175 44743 45209
rect 44777 45175 44943 45209
rect 44977 45175 45143 45209
rect 45177 45175 45343 45209
rect 45377 45175 45543 45209
rect 45577 45175 45743 45209
rect 45777 45175 45943 45209
rect 45977 45175 46143 45209
rect 46177 45175 46343 45209
rect 46377 45175 46543 45209
rect 46577 45175 46743 45209
rect 46777 45175 46943 45209
rect 46977 45175 47143 45209
rect 47177 45175 47343 45209
rect 47377 45175 47543 45209
rect 47577 45175 47743 45209
rect 47777 45175 47943 45209
rect 47977 45175 48143 45209
rect 48177 45175 48343 45209
rect 48377 45175 48543 45209
rect 48577 45175 48743 45209
rect 48777 45175 48943 45209
rect 48977 45175 49143 45209
rect 49177 45175 49343 45209
rect 49377 45175 49543 45209
rect 49577 45175 49743 45209
rect 49777 45175 49943 45209
rect 49977 45175 50143 45209
rect 50177 45175 50343 45209
rect 50377 45175 50543 45209
rect 50577 45175 50743 45209
rect 50777 45175 50943 45209
rect 50977 45175 51143 45209
rect 51177 45175 51343 45209
rect 51377 45175 51543 45209
rect 51577 45175 51743 45209
rect 51777 45175 51943 45209
rect 51977 45175 52143 45209
rect 52177 45175 53478 45209
rect 4958 45134 53478 45175
rect 55066 45134 55088 45250
rect 3348 45132 55088 45134
rect 25608 44957 25636 45132
rect 15071 44941 15117 44957
rect 15071 44907 15077 44941
rect 15111 44907 15117 44941
rect 15071 44869 15117 44907
rect 15071 44835 15077 44869
rect 15111 44835 15117 44869
rect 15071 44797 15117 44835
rect 15071 44763 15077 44797
rect 15111 44763 15117 44797
rect 15071 44725 15117 44763
rect 14124 44689 14170 44712
rect 14124 44655 14130 44689
rect 14164 44655 14170 44689
rect 14124 44617 14170 44655
rect 14124 44583 14130 44617
rect 14164 44583 14170 44617
rect 14124 44545 14170 44583
rect 14124 44511 14130 44545
rect 14164 44511 14170 44545
rect 14124 44473 14170 44511
rect 14124 44439 14130 44473
rect 14164 44439 14170 44473
rect 14124 44401 14170 44439
rect 14124 44367 14130 44401
rect 14164 44367 14170 44401
rect 14124 44329 14170 44367
rect 14124 44295 14130 44329
rect 14164 44295 14170 44329
rect 14124 44257 14170 44295
rect 14124 44223 14130 44257
rect 14164 44223 14170 44257
rect 14124 44185 14170 44223
rect 14124 44151 14130 44185
rect 14164 44151 14170 44185
rect 14124 44113 14170 44151
rect 14124 44079 14130 44113
rect 14164 44079 14170 44113
rect 14124 44041 14170 44079
rect 14124 44007 14130 44041
rect 14164 44007 14170 44041
rect 14124 43969 14170 44007
rect 14124 43935 14130 43969
rect 14164 43935 14170 43969
rect 14124 43912 14170 43935
rect 14582 44689 14628 44712
rect 14582 44655 14588 44689
rect 14622 44655 14628 44689
rect 14582 44617 14628 44655
rect 14582 44583 14588 44617
rect 14622 44583 14628 44617
rect 14582 44545 14628 44583
rect 14582 44511 14588 44545
rect 14622 44511 14628 44545
rect 14582 44473 14628 44511
rect 14582 44439 14588 44473
rect 14622 44439 14628 44473
rect 14582 44401 14628 44439
rect 14582 44367 14588 44401
rect 14622 44367 14628 44401
rect 14582 44329 14628 44367
rect 14582 44295 14588 44329
rect 14622 44295 14628 44329
rect 14582 44257 14628 44295
rect 14582 44223 14588 44257
rect 14622 44223 14628 44257
rect 14582 44185 14628 44223
rect 14582 44151 14588 44185
rect 14622 44151 14628 44185
rect 14582 44113 14628 44151
rect 14582 44079 14588 44113
rect 14622 44079 14628 44113
rect 14582 44041 14628 44079
rect 14582 44007 14588 44041
rect 14622 44007 14628 44041
rect 14582 43976 14628 44007
rect 15071 44691 15077 44725
rect 15111 44691 15117 44725
rect 15071 44653 15117 44691
rect 15071 44619 15077 44653
rect 15111 44619 15117 44653
rect 15071 44581 15117 44619
rect 15071 44547 15077 44581
rect 15111 44547 15117 44581
rect 15071 44509 15117 44547
rect 15071 44475 15077 44509
rect 15111 44475 15117 44509
rect 15071 44437 15117 44475
rect 15071 44403 15077 44437
rect 15111 44403 15117 44437
rect 15071 44365 15117 44403
rect 15071 44331 15077 44365
rect 15111 44331 15117 44365
rect 15071 44293 15117 44331
rect 15071 44259 15077 44293
rect 15111 44259 15117 44293
rect 15071 44221 15117 44259
rect 15071 44187 15077 44221
rect 15111 44187 15117 44221
rect 15071 44149 15117 44187
rect 15071 44115 15077 44149
rect 15111 44115 15117 44149
rect 15071 44077 15117 44115
rect 15071 44043 15077 44077
rect 15111 44043 15117 44077
rect 15071 44005 15117 44043
rect 14582 43969 14688 43976
rect 14582 43935 14588 43969
rect 14622 43948 14688 43969
rect 14622 43935 14628 43948
rect 14582 43912 14628 43935
rect 14366 43704 14372 43716
rect 14311 43676 14372 43704
rect 14366 43664 14372 43676
rect 14424 43664 14430 43716
rect 14550 43500 14556 43512
rect 14495 43472 14556 43500
rect 14550 43460 14556 43472
rect 14608 43460 14614 43512
rect 14660 43372 14688 43948
rect 15071 43971 15077 44005
rect 15111 43971 15117 44005
rect 15071 43933 15117 43971
rect 15071 43899 15077 43933
rect 15111 43899 15117 43933
rect 15071 43861 15117 43899
rect 15071 43827 15077 43861
rect 15111 43827 15117 43861
rect 15071 43789 15117 43827
rect 15071 43755 15077 43789
rect 15111 43755 15117 43789
rect 15071 43717 15117 43755
rect 15071 43683 15077 43717
rect 15111 43683 15117 43717
rect 15071 43667 15117 43683
rect 15529 44941 15575 44957
rect 15529 44907 15535 44941
rect 15569 44907 15575 44941
rect 15529 44869 15575 44907
rect 15529 44835 15535 44869
rect 15569 44835 15575 44869
rect 15529 44797 15575 44835
rect 15529 44763 15535 44797
rect 15569 44763 15575 44797
rect 15529 44725 15575 44763
rect 15529 44691 15535 44725
rect 15569 44691 15575 44725
rect 15529 44653 15575 44691
rect 15529 44619 15535 44653
rect 15569 44619 15575 44653
rect 15529 44581 15575 44619
rect 15529 44547 15535 44581
rect 15569 44547 15575 44581
rect 15529 44509 15575 44547
rect 15529 44475 15535 44509
rect 15569 44475 15575 44509
rect 15529 44437 15575 44475
rect 15529 44403 15535 44437
rect 15569 44403 15575 44437
rect 15529 44365 15575 44403
rect 15529 44331 15535 44365
rect 15569 44331 15575 44365
rect 15529 44293 15575 44331
rect 15529 44259 15535 44293
rect 15569 44259 15575 44293
rect 15529 44221 15575 44259
rect 15529 44187 15535 44221
rect 15569 44187 15575 44221
rect 15529 44149 15575 44187
rect 15529 44115 15535 44149
rect 15569 44115 15575 44149
rect 15529 44077 15575 44115
rect 15529 44043 15535 44077
rect 15569 44043 15575 44077
rect 15529 44005 15575 44043
rect 15529 43971 15535 44005
rect 15569 43971 15575 44005
rect 15529 43933 15575 43971
rect 15529 43899 15535 43933
rect 15569 43899 15575 43933
rect 15529 43861 15575 43899
rect 15529 43827 15535 43861
rect 15569 43827 15575 43861
rect 15529 43789 15575 43827
rect 15529 43755 15535 43789
rect 15569 43755 15575 43789
rect 15529 43717 15575 43755
rect 15529 43683 15535 43717
rect 15569 43683 15575 43717
rect 15529 43667 15575 43683
rect 15987 44941 16033 44957
rect 15987 44907 15993 44941
rect 16027 44907 16033 44941
rect 15987 44869 16033 44907
rect 15987 44835 15993 44869
rect 16027 44835 16033 44869
rect 15987 44797 16033 44835
rect 15987 44763 15993 44797
rect 16027 44763 16033 44797
rect 15987 44725 16033 44763
rect 15987 44691 15993 44725
rect 16027 44691 16033 44725
rect 15987 44653 16033 44691
rect 15987 44619 15993 44653
rect 16027 44619 16033 44653
rect 15987 44581 16033 44619
rect 15987 44547 15993 44581
rect 16027 44547 16033 44581
rect 15987 44509 16033 44547
rect 15987 44475 15993 44509
rect 16027 44475 16033 44509
rect 15987 44437 16033 44475
rect 15987 44403 15993 44437
rect 16027 44403 16033 44437
rect 15987 44365 16033 44403
rect 15987 44331 15993 44365
rect 16027 44331 16033 44365
rect 15987 44293 16033 44331
rect 15987 44259 15993 44293
rect 16027 44259 16033 44293
rect 15987 44221 16033 44259
rect 15987 44187 15993 44221
rect 16027 44187 16033 44221
rect 15987 44149 16033 44187
rect 15987 44115 15993 44149
rect 16027 44115 16033 44149
rect 15987 44077 16033 44115
rect 15987 44043 15993 44077
rect 16027 44043 16033 44077
rect 15987 44005 16033 44043
rect 15987 43971 15993 44005
rect 16027 43971 16033 44005
rect 15987 43933 16033 43971
rect 15987 43899 15993 43933
rect 16027 43899 16033 43933
rect 15987 43861 16033 43899
rect 15987 43827 15993 43861
rect 16027 43827 16033 43861
rect 15987 43789 16033 43827
rect 15987 43755 15993 43789
rect 16027 43755 16033 43789
rect 15987 43717 16033 43755
rect 15987 43683 15993 43717
rect 16027 43683 16033 43717
rect 15987 43667 16033 43683
rect 16445 44941 16491 44957
rect 16445 44907 16451 44941
rect 16485 44907 16491 44941
rect 16445 44869 16491 44907
rect 16445 44835 16451 44869
rect 16485 44835 16491 44869
rect 16445 44797 16491 44835
rect 16445 44763 16451 44797
rect 16485 44763 16491 44797
rect 16445 44725 16491 44763
rect 16445 44691 16451 44725
rect 16485 44691 16491 44725
rect 16445 44653 16491 44691
rect 16445 44619 16451 44653
rect 16485 44619 16491 44653
rect 16445 44581 16491 44619
rect 16445 44547 16451 44581
rect 16485 44547 16491 44581
rect 16445 44509 16491 44547
rect 16445 44475 16451 44509
rect 16485 44475 16491 44509
rect 16445 44437 16491 44475
rect 16445 44403 16451 44437
rect 16485 44403 16491 44437
rect 16445 44365 16491 44403
rect 16445 44331 16451 44365
rect 16485 44331 16491 44365
rect 16445 44293 16491 44331
rect 16445 44259 16451 44293
rect 16485 44259 16491 44293
rect 16445 44221 16491 44259
rect 16445 44187 16451 44221
rect 16485 44187 16491 44221
rect 16445 44149 16491 44187
rect 16445 44115 16451 44149
rect 16485 44115 16491 44149
rect 16445 44077 16491 44115
rect 16445 44043 16451 44077
rect 16485 44043 16491 44077
rect 16445 44005 16491 44043
rect 16445 43971 16451 44005
rect 16485 43971 16491 44005
rect 16445 43933 16491 43971
rect 16445 43899 16451 43933
rect 16485 43899 16491 43933
rect 16445 43861 16491 43899
rect 16445 43827 16451 43861
rect 16485 43827 16491 43861
rect 16445 43789 16491 43827
rect 16445 43755 16451 43789
rect 16485 43755 16491 43789
rect 16445 43717 16491 43755
rect 16445 43683 16451 43717
rect 16485 43683 16491 43717
rect 16445 43667 16491 43683
rect 16903 44941 16949 44957
rect 16903 44907 16909 44941
rect 16943 44907 16949 44941
rect 16903 44869 16949 44907
rect 16903 44835 16909 44869
rect 16943 44835 16949 44869
rect 16903 44797 16949 44835
rect 16903 44763 16909 44797
rect 16943 44763 16949 44797
rect 16903 44725 16949 44763
rect 16903 44691 16909 44725
rect 16943 44691 16949 44725
rect 16903 44653 16949 44691
rect 16903 44619 16909 44653
rect 16943 44619 16949 44653
rect 16903 44581 16949 44619
rect 16903 44547 16909 44581
rect 16943 44547 16949 44581
rect 16903 44509 16949 44547
rect 16903 44475 16909 44509
rect 16943 44475 16949 44509
rect 16903 44437 16949 44475
rect 16903 44403 16909 44437
rect 16943 44403 16949 44437
rect 16903 44365 16949 44403
rect 16903 44331 16909 44365
rect 16943 44331 16949 44365
rect 16903 44293 16949 44331
rect 16903 44259 16909 44293
rect 16943 44259 16949 44293
rect 16903 44221 16949 44259
rect 16903 44187 16909 44221
rect 16943 44187 16949 44221
rect 16903 44149 16949 44187
rect 16903 44115 16909 44149
rect 16943 44115 16949 44149
rect 16903 44077 16949 44115
rect 16903 44043 16909 44077
rect 16943 44043 16949 44077
rect 16903 44005 16949 44043
rect 16903 43971 16909 44005
rect 16943 43971 16949 44005
rect 16903 43933 16949 43971
rect 16903 43899 16909 43933
rect 16943 43899 16949 43933
rect 16903 43861 16949 43899
rect 16903 43827 16909 43861
rect 16943 43827 16949 43861
rect 16903 43789 16949 43827
rect 16903 43755 16909 43789
rect 16943 43755 16949 43789
rect 16903 43717 16949 43755
rect 16903 43683 16909 43717
rect 16943 43683 16949 43717
rect 16903 43667 16949 43683
rect 17361 44941 17407 44957
rect 17361 44907 17367 44941
rect 17401 44907 17407 44941
rect 17361 44869 17407 44907
rect 17361 44835 17367 44869
rect 17401 44835 17407 44869
rect 17361 44797 17407 44835
rect 17361 44763 17367 44797
rect 17401 44763 17407 44797
rect 17361 44725 17407 44763
rect 17361 44691 17367 44725
rect 17401 44691 17407 44725
rect 17361 44653 17407 44691
rect 17361 44619 17367 44653
rect 17401 44619 17407 44653
rect 17361 44581 17407 44619
rect 17361 44547 17367 44581
rect 17401 44547 17407 44581
rect 17361 44509 17407 44547
rect 17361 44475 17367 44509
rect 17401 44475 17407 44509
rect 17361 44437 17407 44475
rect 17361 44403 17367 44437
rect 17401 44403 17407 44437
rect 17361 44365 17407 44403
rect 17361 44331 17367 44365
rect 17401 44331 17407 44365
rect 17361 44293 17407 44331
rect 17361 44259 17367 44293
rect 17401 44259 17407 44293
rect 17361 44221 17407 44259
rect 17361 44187 17367 44221
rect 17401 44187 17407 44221
rect 17361 44149 17407 44187
rect 17361 44115 17367 44149
rect 17401 44115 17407 44149
rect 17361 44077 17407 44115
rect 17361 44043 17367 44077
rect 17401 44043 17407 44077
rect 17361 44005 17407 44043
rect 17361 43971 17367 44005
rect 17401 43971 17407 44005
rect 17361 43933 17407 43971
rect 17361 43899 17367 43933
rect 17401 43899 17407 43933
rect 17361 43861 17407 43899
rect 17361 43827 17367 43861
rect 17401 43827 17407 43861
rect 17361 43789 17407 43827
rect 17361 43755 17367 43789
rect 17401 43755 17407 43789
rect 17361 43717 17407 43755
rect 17361 43683 17367 43717
rect 17401 43683 17407 43717
rect 17361 43667 17407 43683
rect 17819 44941 17865 44957
rect 17819 44907 17825 44941
rect 17859 44907 17865 44941
rect 17819 44869 17865 44907
rect 17819 44835 17825 44869
rect 17859 44835 17865 44869
rect 17819 44797 17865 44835
rect 17819 44763 17825 44797
rect 17859 44763 17865 44797
rect 17819 44725 17865 44763
rect 17819 44691 17825 44725
rect 17859 44691 17865 44725
rect 17819 44653 17865 44691
rect 17819 44619 17825 44653
rect 17859 44619 17865 44653
rect 17819 44581 17865 44619
rect 17819 44547 17825 44581
rect 17859 44547 17865 44581
rect 17819 44509 17865 44547
rect 17819 44475 17825 44509
rect 17859 44475 17865 44509
rect 17819 44437 17865 44475
rect 17819 44403 17825 44437
rect 17859 44403 17865 44437
rect 17819 44365 17865 44403
rect 17819 44331 17825 44365
rect 17859 44331 17865 44365
rect 17819 44293 17865 44331
rect 17819 44259 17825 44293
rect 17859 44259 17865 44293
rect 17819 44221 17865 44259
rect 17819 44187 17825 44221
rect 17859 44187 17865 44221
rect 17819 44149 17865 44187
rect 17819 44115 17825 44149
rect 17859 44115 17865 44149
rect 17819 44077 17865 44115
rect 17819 44043 17825 44077
rect 17859 44043 17865 44077
rect 17819 44005 17865 44043
rect 17819 43971 17825 44005
rect 17859 43971 17865 44005
rect 17819 43933 17865 43971
rect 17819 43899 17825 43933
rect 17859 43899 17865 43933
rect 17819 43861 17865 43899
rect 17819 43827 17825 43861
rect 17859 43827 17865 43861
rect 17819 43789 17865 43827
rect 17819 43755 17825 43789
rect 17859 43755 17865 43789
rect 17819 43717 17865 43755
rect 17819 43683 17825 43717
rect 17859 43683 17865 43717
rect 17819 43667 17865 43683
rect 18277 44941 18323 44957
rect 18277 44907 18283 44941
rect 18317 44907 18323 44941
rect 18277 44869 18323 44907
rect 18277 44835 18283 44869
rect 18317 44835 18323 44869
rect 18277 44797 18323 44835
rect 18277 44763 18283 44797
rect 18317 44763 18323 44797
rect 18277 44725 18323 44763
rect 18277 44691 18283 44725
rect 18317 44691 18323 44725
rect 18277 44653 18323 44691
rect 18277 44619 18283 44653
rect 18317 44619 18323 44653
rect 18277 44581 18323 44619
rect 18277 44547 18283 44581
rect 18317 44547 18323 44581
rect 18277 44509 18323 44547
rect 18277 44475 18283 44509
rect 18317 44475 18323 44509
rect 18277 44437 18323 44475
rect 18277 44403 18283 44437
rect 18317 44403 18323 44437
rect 18277 44365 18323 44403
rect 18277 44331 18283 44365
rect 18317 44331 18323 44365
rect 18277 44293 18323 44331
rect 18277 44259 18283 44293
rect 18317 44259 18323 44293
rect 18277 44221 18323 44259
rect 18277 44187 18283 44221
rect 18317 44187 18323 44221
rect 18277 44149 18323 44187
rect 18277 44115 18283 44149
rect 18317 44115 18323 44149
rect 18277 44077 18323 44115
rect 18277 44043 18283 44077
rect 18317 44043 18323 44077
rect 18277 44005 18323 44043
rect 18277 43971 18283 44005
rect 18317 43971 18323 44005
rect 18277 43933 18323 43971
rect 18277 43899 18283 43933
rect 18317 43899 18323 43933
rect 18277 43861 18323 43899
rect 18277 43827 18283 43861
rect 18317 43827 18323 43861
rect 18277 43789 18323 43827
rect 18277 43755 18283 43789
rect 18317 43755 18323 43789
rect 18277 43717 18323 43755
rect 18277 43683 18283 43717
rect 18317 43683 18323 43717
rect 18277 43667 18323 43683
rect 18735 44941 18781 44957
rect 18735 44907 18741 44941
rect 18775 44907 18781 44941
rect 18735 44869 18781 44907
rect 18735 44835 18741 44869
rect 18775 44835 18781 44869
rect 18735 44797 18781 44835
rect 18735 44763 18741 44797
rect 18775 44763 18781 44797
rect 18735 44725 18781 44763
rect 18735 44691 18741 44725
rect 18775 44691 18781 44725
rect 18735 44653 18781 44691
rect 18735 44619 18741 44653
rect 18775 44619 18781 44653
rect 18735 44581 18781 44619
rect 18735 44547 18741 44581
rect 18775 44547 18781 44581
rect 18735 44509 18781 44547
rect 18735 44475 18741 44509
rect 18775 44475 18781 44509
rect 18735 44437 18781 44475
rect 18735 44403 18741 44437
rect 18775 44403 18781 44437
rect 18735 44365 18781 44403
rect 18735 44331 18741 44365
rect 18775 44331 18781 44365
rect 18735 44293 18781 44331
rect 18735 44259 18741 44293
rect 18775 44259 18781 44293
rect 18735 44221 18781 44259
rect 18735 44187 18741 44221
rect 18775 44187 18781 44221
rect 18735 44149 18781 44187
rect 18735 44115 18741 44149
rect 18775 44115 18781 44149
rect 18735 44077 18781 44115
rect 18735 44043 18741 44077
rect 18775 44043 18781 44077
rect 18735 44005 18781 44043
rect 18735 43971 18741 44005
rect 18775 43971 18781 44005
rect 18735 43933 18781 43971
rect 18735 43899 18741 43933
rect 18775 43899 18781 43933
rect 18735 43861 18781 43899
rect 18735 43827 18741 43861
rect 18775 43827 18781 43861
rect 18735 43789 18781 43827
rect 18735 43755 18741 43789
rect 18775 43755 18781 43789
rect 18735 43717 18781 43755
rect 18735 43683 18741 43717
rect 18775 43683 18781 43717
rect 18735 43667 18781 43683
rect 19193 44941 19239 44957
rect 19193 44907 19199 44941
rect 19233 44907 19239 44941
rect 19193 44869 19239 44907
rect 19193 44835 19199 44869
rect 19233 44835 19239 44869
rect 19193 44797 19239 44835
rect 19193 44763 19199 44797
rect 19233 44763 19239 44797
rect 19193 44725 19239 44763
rect 19193 44691 19199 44725
rect 19233 44691 19239 44725
rect 19193 44653 19239 44691
rect 19193 44619 19199 44653
rect 19233 44619 19239 44653
rect 19193 44581 19239 44619
rect 19193 44547 19199 44581
rect 19233 44547 19239 44581
rect 19193 44509 19239 44547
rect 19193 44475 19199 44509
rect 19233 44475 19239 44509
rect 19193 44437 19239 44475
rect 19193 44403 19199 44437
rect 19233 44403 19239 44437
rect 19193 44365 19239 44403
rect 19193 44331 19199 44365
rect 19233 44331 19239 44365
rect 19193 44293 19239 44331
rect 19193 44259 19199 44293
rect 19233 44259 19239 44293
rect 19193 44221 19239 44259
rect 19193 44187 19199 44221
rect 19233 44187 19239 44221
rect 19193 44149 19239 44187
rect 19193 44115 19199 44149
rect 19233 44115 19239 44149
rect 19193 44077 19239 44115
rect 19193 44043 19199 44077
rect 19233 44043 19239 44077
rect 19193 44005 19239 44043
rect 19193 43971 19199 44005
rect 19233 43971 19239 44005
rect 19193 43933 19239 43971
rect 19193 43899 19199 43933
rect 19233 43899 19239 43933
rect 19193 43861 19239 43899
rect 19193 43827 19199 43861
rect 19233 43827 19239 43861
rect 19193 43789 19239 43827
rect 19193 43755 19199 43789
rect 19233 43755 19239 43789
rect 19193 43717 19239 43755
rect 19193 43683 19199 43717
rect 19233 43683 19239 43717
rect 19193 43667 19239 43683
rect 19651 44941 19697 44957
rect 19651 44907 19657 44941
rect 19691 44907 19697 44941
rect 19651 44869 19697 44907
rect 19651 44835 19657 44869
rect 19691 44835 19697 44869
rect 19651 44797 19697 44835
rect 19651 44763 19657 44797
rect 19691 44763 19697 44797
rect 19651 44725 19697 44763
rect 19651 44691 19657 44725
rect 19691 44691 19697 44725
rect 19651 44653 19697 44691
rect 19651 44619 19657 44653
rect 19691 44619 19697 44653
rect 19651 44581 19697 44619
rect 19651 44547 19657 44581
rect 19691 44547 19697 44581
rect 19651 44509 19697 44547
rect 19651 44475 19657 44509
rect 19691 44475 19697 44509
rect 19651 44437 19697 44475
rect 19651 44403 19657 44437
rect 19691 44403 19697 44437
rect 19651 44365 19697 44403
rect 19651 44331 19657 44365
rect 19691 44331 19697 44365
rect 19651 44293 19697 44331
rect 19651 44259 19657 44293
rect 19691 44259 19697 44293
rect 19651 44221 19697 44259
rect 19651 44187 19657 44221
rect 19691 44187 19697 44221
rect 19651 44149 19697 44187
rect 19651 44115 19657 44149
rect 19691 44115 19697 44149
rect 19651 44077 19697 44115
rect 19651 44043 19657 44077
rect 19691 44043 19697 44077
rect 19651 44005 19697 44043
rect 19651 43971 19657 44005
rect 19691 43971 19697 44005
rect 19651 43933 19697 43971
rect 19651 43899 19657 43933
rect 19691 43899 19697 43933
rect 19651 43861 19697 43899
rect 19651 43827 19657 43861
rect 19691 43827 19697 43861
rect 19651 43789 19697 43827
rect 19651 43755 19657 43789
rect 19691 43755 19697 43789
rect 19651 43717 19697 43755
rect 19651 43683 19657 43717
rect 19691 43683 19697 43717
rect 19651 43667 19697 43683
rect 20109 44941 20155 44957
rect 20109 44907 20115 44941
rect 20149 44907 20155 44941
rect 20109 44869 20155 44907
rect 20109 44835 20115 44869
rect 20149 44835 20155 44869
rect 20109 44797 20155 44835
rect 20109 44763 20115 44797
rect 20149 44763 20155 44797
rect 20109 44725 20155 44763
rect 20109 44691 20115 44725
rect 20149 44691 20155 44725
rect 20109 44653 20155 44691
rect 20109 44619 20115 44653
rect 20149 44619 20155 44653
rect 20109 44581 20155 44619
rect 20109 44547 20115 44581
rect 20149 44547 20155 44581
rect 20109 44509 20155 44547
rect 20109 44475 20115 44509
rect 20149 44475 20155 44509
rect 20109 44437 20155 44475
rect 20109 44403 20115 44437
rect 20149 44403 20155 44437
rect 20109 44365 20155 44403
rect 20109 44331 20115 44365
rect 20149 44331 20155 44365
rect 20109 44293 20155 44331
rect 20109 44259 20115 44293
rect 20149 44259 20155 44293
rect 20109 44221 20155 44259
rect 20109 44187 20115 44221
rect 20149 44187 20155 44221
rect 20109 44149 20155 44187
rect 20109 44115 20115 44149
rect 20149 44115 20155 44149
rect 20109 44077 20155 44115
rect 20109 44043 20115 44077
rect 20149 44043 20155 44077
rect 20109 44005 20155 44043
rect 20109 43971 20115 44005
rect 20149 43971 20155 44005
rect 20109 43933 20155 43971
rect 20109 43899 20115 43933
rect 20149 43899 20155 43933
rect 20109 43861 20155 43899
rect 20109 43827 20115 43861
rect 20149 43827 20155 43861
rect 20109 43789 20155 43827
rect 20109 43755 20115 43789
rect 20149 43755 20155 43789
rect 20109 43717 20155 43755
rect 20109 43683 20115 43717
rect 20149 43683 20155 43717
rect 20109 43667 20155 43683
rect 20567 44941 20613 44957
rect 20567 44907 20573 44941
rect 20607 44907 20613 44941
rect 20567 44869 20613 44907
rect 20567 44835 20573 44869
rect 20607 44835 20613 44869
rect 20567 44797 20613 44835
rect 20567 44763 20573 44797
rect 20607 44763 20613 44797
rect 20567 44725 20613 44763
rect 20567 44691 20573 44725
rect 20607 44691 20613 44725
rect 20567 44653 20613 44691
rect 20567 44619 20573 44653
rect 20607 44619 20613 44653
rect 20567 44581 20613 44619
rect 20567 44547 20573 44581
rect 20607 44547 20613 44581
rect 20567 44509 20613 44547
rect 20567 44475 20573 44509
rect 20607 44475 20613 44509
rect 20567 44437 20613 44475
rect 20567 44403 20573 44437
rect 20607 44403 20613 44437
rect 20567 44365 20613 44403
rect 20567 44331 20573 44365
rect 20607 44331 20613 44365
rect 20567 44293 20613 44331
rect 20567 44259 20573 44293
rect 20607 44259 20613 44293
rect 20567 44221 20613 44259
rect 20567 44187 20573 44221
rect 20607 44187 20613 44221
rect 20567 44149 20613 44187
rect 20567 44115 20573 44149
rect 20607 44115 20613 44149
rect 20567 44077 20613 44115
rect 20567 44043 20573 44077
rect 20607 44043 20613 44077
rect 20567 44005 20613 44043
rect 20567 43971 20573 44005
rect 20607 43971 20613 44005
rect 20567 43933 20613 43971
rect 20567 43899 20573 43933
rect 20607 43899 20613 43933
rect 20567 43861 20613 43899
rect 20567 43827 20573 43861
rect 20607 43827 20613 43861
rect 20567 43789 20613 43827
rect 20567 43755 20573 43789
rect 20607 43755 20613 43789
rect 20567 43717 20613 43755
rect 20567 43683 20573 43717
rect 20607 43683 20613 43717
rect 20567 43667 20613 43683
rect 21025 44941 21071 44957
rect 21025 44907 21031 44941
rect 21065 44907 21071 44941
rect 21025 44869 21071 44907
rect 21025 44835 21031 44869
rect 21065 44835 21071 44869
rect 21025 44797 21071 44835
rect 21025 44763 21031 44797
rect 21065 44763 21071 44797
rect 21025 44725 21071 44763
rect 21025 44691 21031 44725
rect 21065 44691 21071 44725
rect 21025 44653 21071 44691
rect 21025 44619 21031 44653
rect 21065 44619 21071 44653
rect 21025 44581 21071 44619
rect 21025 44547 21031 44581
rect 21065 44547 21071 44581
rect 21025 44509 21071 44547
rect 21025 44475 21031 44509
rect 21065 44475 21071 44509
rect 21025 44437 21071 44475
rect 21025 44403 21031 44437
rect 21065 44403 21071 44437
rect 21025 44365 21071 44403
rect 21025 44331 21031 44365
rect 21065 44331 21071 44365
rect 21025 44293 21071 44331
rect 21025 44259 21031 44293
rect 21065 44259 21071 44293
rect 21025 44221 21071 44259
rect 21025 44187 21031 44221
rect 21065 44187 21071 44221
rect 21025 44149 21071 44187
rect 21025 44115 21031 44149
rect 21065 44115 21071 44149
rect 21025 44077 21071 44115
rect 21025 44043 21031 44077
rect 21065 44043 21071 44077
rect 21025 44005 21071 44043
rect 21025 43971 21031 44005
rect 21065 43971 21071 44005
rect 21025 43933 21071 43971
rect 21025 43899 21031 43933
rect 21065 43899 21071 43933
rect 21025 43861 21071 43899
rect 21025 43827 21031 43861
rect 21065 43827 21071 43861
rect 21025 43789 21071 43827
rect 21025 43755 21031 43789
rect 21065 43755 21071 43789
rect 21025 43717 21071 43755
rect 21025 43683 21031 43717
rect 21065 43683 21071 43717
rect 21025 43667 21071 43683
rect 21483 44941 21529 44957
rect 21483 44907 21489 44941
rect 21523 44907 21529 44941
rect 21483 44869 21529 44907
rect 21483 44835 21489 44869
rect 21523 44835 21529 44869
rect 21483 44797 21529 44835
rect 21483 44763 21489 44797
rect 21523 44763 21529 44797
rect 21483 44725 21529 44763
rect 21483 44691 21489 44725
rect 21523 44691 21529 44725
rect 21483 44653 21529 44691
rect 21483 44619 21489 44653
rect 21523 44619 21529 44653
rect 21483 44581 21529 44619
rect 21483 44547 21489 44581
rect 21523 44547 21529 44581
rect 21483 44509 21529 44547
rect 21483 44475 21489 44509
rect 21523 44475 21529 44509
rect 21483 44437 21529 44475
rect 21483 44403 21489 44437
rect 21523 44403 21529 44437
rect 21483 44365 21529 44403
rect 21483 44331 21489 44365
rect 21523 44331 21529 44365
rect 21483 44293 21529 44331
rect 21483 44259 21489 44293
rect 21523 44259 21529 44293
rect 21483 44221 21529 44259
rect 21483 44187 21489 44221
rect 21523 44187 21529 44221
rect 21483 44149 21529 44187
rect 21483 44115 21489 44149
rect 21523 44115 21529 44149
rect 21483 44077 21529 44115
rect 21483 44043 21489 44077
rect 21523 44043 21529 44077
rect 21483 44005 21529 44043
rect 21483 43971 21489 44005
rect 21523 43971 21529 44005
rect 21483 43933 21529 43971
rect 21483 43899 21489 43933
rect 21523 43899 21529 43933
rect 21483 43861 21529 43899
rect 21483 43827 21489 43861
rect 21523 43827 21529 43861
rect 21483 43789 21529 43827
rect 21483 43755 21489 43789
rect 21523 43755 21529 43789
rect 21483 43717 21529 43755
rect 21483 43683 21489 43717
rect 21523 43683 21529 43717
rect 21483 43667 21529 43683
rect 21941 44941 21987 44957
rect 21941 44907 21947 44941
rect 21981 44907 21987 44941
rect 21941 44869 21987 44907
rect 21941 44835 21947 44869
rect 21981 44835 21987 44869
rect 21941 44797 21987 44835
rect 21941 44763 21947 44797
rect 21981 44763 21987 44797
rect 21941 44725 21987 44763
rect 21941 44691 21947 44725
rect 21981 44691 21987 44725
rect 21941 44653 21987 44691
rect 21941 44619 21947 44653
rect 21981 44619 21987 44653
rect 21941 44581 21987 44619
rect 21941 44547 21947 44581
rect 21981 44547 21987 44581
rect 21941 44509 21987 44547
rect 21941 44475 21947 44509
rect 21981 44475 21987 44509
rect 21941 44437 21987 44475
rect 21941 44403 21947 44437
rect 21981 44403 21987 44437
rect 21941 44365 21987 44403
rect 21941 44331 21947 44365
rect 21981 44331 21987 44365
rect 21941 44293 21987 44331
rect 21941 44259 21947 44293
rect 21981 44259 21987 44293
rect 21941 44221 21987 44259
rect 21941 44187 21947 44221
rect 21981 44187 21987 44221
rect 21941 44149 21987 44187
rect 21941 44115 21947 44149
rect 21981 44115 21987 44149
rect 21941 44077 21987 44115
rect 21941 44043 21947 44077
rect 21981 44043 21987 44077
rect 21941 44005 21987 44043
rect 21941 43971 21947 44005
rect 21981 43971 21987 44005
rect 21941 43933 21987 43971
rect 21941 43899 21947 43933
rect 21981 43899 21987 43933
rect 21941 43861 21987 43899
rect 21941 43827 21947 43861
rect 21981 43827 21987 43861
rect 21941 43789 21987 43827
rect 21941 43755 21947 43789
rect 21981 43755 21987 43789
rect 21941 43717 21987 43755
rect 21941 43683 21947 43717
rect 21981 43683 21987 43717
rect 22399 44941 22445 44957
rect 22399 44907 22405 44941
rect 22439 44907 22445 44941
rect 22399 44869 22445 44907
rect 22399 44835 22405 44869
rect 22439 44835 22445 44869
rect 22399 44797 22445 44835
rect 22399 44763 22405 44797
rect 22439 44763 22445 44797
rect 22399 44725 22445 44763
rect 22399 44691 22405 44725
rect 22439 44691 22445 44725
rect 22399 44653 22445 44691
rect 22399 44619 22405 44653
rect 22439 44619 22445 44653
rect 22399 44581 22445 44619
rect 22399 44547 22405 44581
rect 22439 44547 22445 44581
rect 22399 44509 22445 44547
rect 22399 44475 22405 44509
rect 22439 44475 22445 44509
rect 22399 44437 22445 44475
rect 22399 44403 22405 44437
rect 22439 44403 22445 44437
rect 22399 44365 22445 44403
rect 22399 44331 22405 44365
rect 22439 44331 22445 44365
rect 22399 44293 22445 44331
rect 22399 44259 22405 44293
rect 22439 44259 22445 44293
rect 22399 44221 22445 44259
rect 22399 44187 22405 44221
rect 22439 44187 22445 44221
rect 22399 44149 22445 44187
rect 22399 44115 22405 44149
rect 22439 44115 22445 44149
rect 22399 44077 22445 44115
rect 22399 44043 22405 44077
rect 22439 44043 22445 44077
rect 22399 44005 22445 44043
rect 22399 43971 22405 44005
rect 22439 43971 22445 44005
rect 22399 43933 22445 43971
rect 22399 43899 22405 43933
rect 22439 43899 22445 43933
rect 22399 43861 22445 43899
rect 22399 43827 22405 43861
rect 22439 43827 22445 43861
rect 22399 43789 22445 43827
rect 22399 43755 22405 43789
rect 22439 43755 22445 43789
rect 22399 43717 22445 43755
rect 21941 43667 21987 43683
rect 22186 43664 22192 43716
rect 22244 43704 22250 43716
rect 22399 43704 22405 43717
rect 22244 43683 22405 43704
rect 22439 43683 22445 43717
rect 22244 43676 22445 43683
rect 22244 43664 22250 43676
rect 22399 43667 22445 43676
rect 22857 44941 22903 44957
rect 22857 44907 22863 44941
rect 22897 44907 22903 44941
rect 22857 44869 22903 44907
rect 22857 44835 22863 44869
rect 22897 44835 22903 44869
rect 22857 44797 22903 44835
rect 22857 44763 22863 44797
rect 22897 44763 22903 44797
rect 22857 44725 22903 44763
rect 22857 44691 22863 44725
rect 22897 44691 22903 44725
rect 22857 44653 22903 44691
rect 22857 44619 22863 44653
rect 22897 44619 22903 44653
rect 22857 44581 22903 44619
rect 22857 44547 22863 44581
rect 22897 44547 22903 44581
rect 22857 44509 22903 44547
rect 22857 44475 22863 44509
rect 22897 44475 22903 44509
rect 22857 44437 22903 44475
rect 22857 44403 22863 44437
rect 22897 44403 22903 44437
rect 22857 44365 22903 44403
rect 22857 44331 22863 44365
rect 22897 44331 22903 44365
rect 22857 44293 22903 44331
rect 22857 44259 22863 44293
rect 22897 44259 22903 44293
rect 22857 44221 22903 44259
rect 22857 44187 22863 44221
rect 22897 44187 22903 44221
rect 22857 44149 22903 44187
rect 22857 44115 22863 44149
rect 22897 44115 22903 44149
rect 22857 44077 22903 44115
rect 22857 44043 22863 44077
rect 22897 44043 22903 44077
rect 22857 44005 22903 44043
rect 22857 43971 22863 44005
rect 22897 43971 22903 44005
rect 22857 43933 22903 43971
rect 22857 43899 22863 43933
rect 22897 43899 22903 43933
rect 22857 43861 22903 43899
rect 22857 43827 22863 43861
rect 22897 43827 22903 43861
rect 22857 43789 22903 43827
rect 22857 43755 22863 43789
rect 22897 43755 22903 43789
rect 22857 43717 22903 43755
rect 22857 43683 22863 43717
rect 22897 43683 22903 43717
rect 22857 43667 22903 43683
rect 23315 44941 23361 44957
rect 23315 44907 23321 44941
rect 23355 44907 23361 44941
rect 23315 44869 23361 44907
rect 23315 44835 23321 44869
rect 23355 44835 23361 44869
rect 23315 44797 23361 44835
rect 23315 44763 23321 44797
rect 23355 44763 23361 44797
rect 23315 44725 23361 44763
rect 23315 44691 23321 44725
rect 23355 44691 23361 44725
rect 23315 44653 23361 44691
rect 23315 44619 23321 44653
rect 23355 44619 23361 44653
rect 23315 44581 23361 44619
rect 23315 44547 23321 44581
rect 23355 44547 23361 44581
rect 23315 44509 23361 44547
rect 23315 44475 23321 44509
rect 23355 44475 23361 44509
rect 23315 44437 23361 44475
rect 23315 44403 23321 44437
rect 23355 44403 23361 44437
rect 23315 44365 23361 44403
rect 23315 44331 23321 44365
rect 23355 44331 23361 44365
rect 23315 44293 23361 44331
rect 23315 44259 23321 44293
rect 23355 44259 23361 44293
rect 23315 44221 23361 44259
rect 23315 44187 23321 44221
rect 23355 44187 23361 44221
rect 23315 44149 23361 44187
rect 23315 44115 23321 44149
rect 23355 44115 23361 44149
rect 23315 44077 23361 44115
rect 23315 44043 23321 44077
rect 23355 44043 23361 44077
rect 23315 44005 23361 44043
rect 23315 43971 23321 44005
rect 23355 43971 23361 44005
rect 23315 43933 23361 43971
rect 23315 43899 23321 43933
rect 23355 43899 23361 43933
rect 23315 43861 23361 43899
rect 23315 43827 23321 43861
rect 23355 43827 23361 43861
rect 23315 43789 23361 43827
rect 23315 43755 23321 43789
rect 23355 43755 23361 43789
rect 23315 43717 23361 43755
rect 23315 43683 23321 43717
rect 23355 43683 23361 43717
rect 23315 43667 23361 43683
rect 23773 44941 23819 44957
rect 23773 44907 23779 44941
rect 23813 44907 23819 44941
rect 23773 44869 23819 44907
rect 23773 44835 23779 44869
rect 23813 44835 23819 44869
rect 23773 44797 23819 44835
rect 23773 44763 23779 44797
rect 23813 44763 23819 44797
rect 23773 44725 23819 44763
rect 23773 44691 23779 44725
rect 23813 44691 23819 44725
rect 23773 44653 23819 44691
rect 23773 44619 23779 44653
rect 23813 44619 23819 44653
rect 23773 44581 23819 44619
rect 23773 44547 23779 44581
rect 23813 44547 23819 44581
rect 23773 44509 23819 44547
rect 23773 44475 23779 44509
rect 23813 44475 23819 44509
rect 23773 44437 23819 44475
rect 23773 44403 23779 44437
rect 23813 44403 23819 44437
rect 23773 44365 23819 44403
rect 23773 44331 23779 44365
rect 23813 44331 23819 44365
rect 23773 44293 23819 44331
rect 23773 44259 23779 44293
rect 23813 44259 23819 44293
rect 23773 44221 23819 44259
rect 23773 44187 23779 44221
rect 23813 44187 23819 44221
rect 23773 44149 23819 44187
rect 23773 44115 23779 44149
rect 23813 44115 23819 44149
rect 23773 44077 23819 44115
rect 23773 44043 23779 44077
rect 23813 44043 23819 44077
rect 23773 44005 23819 44043
rect 23773 43971 23779 44005
rect 23813 43971 23819 44005
rect 23773 43933 23819 43971
rect 23773 43899 23779 43933
rect 23813 43899 23819 43933
rect 23773 43861 23819 43899
rect 23773 43827 23779 43861
rect 23813 43827 23819 43861
rect 23773 43789 23819 43827
rect 23773 43755 23779 43789
rect 23813 43755 23819 43789
rect 23773 43717 23819 43755
rect 23773 43683 23779 43717
rect 23813 43683 23819 43717
rect 23773 43667 23819 43683
rect 24231 44941 24277 44957
rect 24231 44907 24237 44941
rect 24271 44907 24277 44941
rect 24231 44869 24277 44907
rect 24231 44835 24237 44869
rect 24271 44835 24277 44869
rect 24231 44797 24277 44835
rect 24231 44763 24237 44797
rect 24271 44763 24277 44797
rect 24231 44725 24277 44763
rect 24231 44691 24237 44725
rect 24271 44691 24277 44725
rect 24231 44653 24277 44691
rect 24231 44619 24237 44653
rect 24271 44619 24277 44653
rect 24231 44581 24277 44619
rect 24231 44547 24237 44581
rect 24271 44547 24277 44581
rect 24231 44509 24277 44547
rect 24231 44475 24237 44509
rect 24271 44475 24277 44509
rect 24231 44437 24277 44475
rect 24231 44403 24237 44437
rect 24271 44403 24277 44437
rect 24231 44365 24277 44403
rect 24231 44331 24237 44365
rect 24271 44331 24277 44365
rect 24231 44293 24277 44331
rect 24231 44259 24237 44293
rect 24271 44259 24277 44293
rect 24231 44221 24277 44259
rect 24231 44187 24237 44221
rect 24271 44187 24277 44221
rect 24231 44149 24277 44187
rect 24231 44115 24237 44149
rect 24271 44115 24277 44149
rect 24231 44077 24277 44115
rect 24231 44043 24237 44077
rect 24271 44043 24277 44077
rect 24231 44005 24277 44043
rect 24231 43971 24237 44005
rect 24271 43971 24277 44005
rect 24231 43933 24277 43971
rect 24231 43899 24237 43933
rect 24271 43899 24277 43933
rect 24231 43861 24277 43899
rect 24231 43827 24237 43861
rect 24271 43827 24277 43861
rect 24231 43789 24277 43827
rect 24231 43755 24237 43789
rect 24271 43755 24277 43789
rect 24231 43717 24277 43755
rect 24231 43683 24237 43717
rect 24271 43683 24277 43717
rect 24231 43667 24277 43683
rect 24689 44941 24735 44957
rect 24689 44907 24695 44941
rect 24729 44907 24735 44941
rect 24689 44869 24735 44907
rect 24689 44835 24695 44869
rect 24729 44835 24735 44869
rect 24689 44797 24735 44835
rect 24689 44763 24695 44797
rect 24729 44763 24735 44797
rect 24689 44725 24735 44763
rect 24689 44691 24695 44725
rect 24729 44691 24735 44725
rect 24689 44653 24735 44691
rect 24689 44619 24695 44653
rect 24729 44619 24735 44653
rect 24689 44581 24735 44619
rect 24689 44547 24695 44581
rect 24729 44547 24735 44581
rect 24689 44509 24735 44547
rect 24689 44475 24695 44509
rect 24729 44475 24735 44509
rect 24689 44437 24735 44475
rect 24689 44403 24695 44437
rect 24729 44403 24735 44437
rect 24689 44365 24735 44403
rect 24689 44331 24695 44365
rect 24729 44331 24735 44365
rect 24689 44293 24735 44331
rect 24689 44259 24695 44293
rect 24729 44259 24735 44293
rect 24689 44221 24735 44259
rect 24689 44187 24695 44221
rect 24729 44187 24735 44221
rect 24689 44149 24735 44187
rect 24689 44115 24695 44149
rect 24729 44115 24735 44149
rect 24689 44077 24735 44115
rect 24689 44043 24695 44077
rect 24729 44043 24735 44077
rect 24689 44005 24735 44043
rect 24689 43971 24695 44005
rect 24729 43971 24735 44005
rect 24689 43933 24735 43971
rect 24689 43899 24695 43933
rect 24729 43899 24735 43933
rect 24689 43861 24735 43899
rect 24689 43827 24695 43861
rect 24729 43827 24735 43861
rect 24689 43789 24735 43827
rect 24689 43755 24695 43789
rect 24729 43755 24735 43789
rect 24689 43717 24735 43755
rect 24689 43683 24695 43717
rect 24729 43683 24735 43717
rect 24689 43667 24735 43683
rect 25147 44941 25193 44957
rect 25147 44907 25153 44941
rect 25187 44907 25193 44941
rect 25147 44869 25193 44907
rect 25147 44835 25153 44869
rect 25187 44835 25193 44869
rect 25147 44797 25193 44835
rect 25147 44763 25153 44797
rect 25187 44763 25193 44797
rect 25147 44725 25193 44763
rect 25147 44691 25153 44725
rect 25187 44691 25193 44725
rect 25147 44653 25193 44691
rect 25147 44619 25153 44653
rect 25187 44619 25193 44653
rect 25147 44581 25193 44619
rect 25147 44547 25153 44581
rect 25187 44547 25193 44581
rect 25147 44509 25193 44547
rect 25147 44475 25153 44509
rect 25187 44475 25193 44509
rect 25147 44437 25193 44475
rect 25147 44403 25153 44437
rect 25187 44403 25193 44437
rect 25147 44365 25193 44403
rect 25147 44331 25153 44365
rect 25187 44331 25193 44365
rect 25147 44293 25193 44331
rect 25147 44259 25153 44293
rect 25187 44259 25193 44293
rect 25147 44221 25193 44259
rect 25147 44187 25153 44221
rect 25187 44187 25193 44221
rect 25147 44149 25193 44187
rect 25147 44115 25153 44149
rect 25187 44115 25193 44149
rect 25147 44077 25193 44115
rect 25147 44043 25153 44077
rect 25187 44043 25193 44077
rect 25147 44005 25193 44043
rect 25147 43971 25153 44005
rect 25187 43971 25193 44005
rect 25147 43933 25193 43971
rect 25147 43899 25153 43933
rect 25187 43899 25193 43933
rect 25147 43861 25193 43899
rect 25147 43827 25153 43861
rect 25187 43827 25193 43861
rect 25147 43789 25193 43827
rect 25147 43755 25153 43789
rect 25187 43755 25193 43789
rect 25147 43717 25193 43755
rect 25147 43683 25153 43717
rect 25187 43683 25193 43717
rect 25147 43667 25193 43683
rect 25605 44941 25651 44957
rect 25605 44907 25611 44941
rect 25645 44907 25651 44941
rect 25605 44869 25651 44907
rect 25605 44835 25611 44869
rect 25645 44835 25651 44869
rect 25605 44797 25651 44835
rect 25605 44763 25611 44797
rect 25645 44763 25651 44797
rect 25605 44725 25651 44763
rect 25605 44691 25611 44725
rect 25645 44691 25651 44725
rect 25605 44653 25651 44691
rect 25605 44619 25611 44653
rect 25645 44619 25651 44653
rect 25605 44581 25651 44619
rect 25605 44547 25611 44581
rect 25645 44547 25651 44581
rect 25605 44509 25651 44547
rect 25605 44475 25611 44509
rect 25645 44475 25651 44509
rect 25605 44437 25651 44475
rect 25605 44403 25611 44437
rect 25645 44403 25651 44437
rect 25605 44365 25651 44403
rect 25605 44331 25611 44365
rect 25645 44331 25651 44365
rect 25605 44293 25651 44331
rect 25605 44259 25611 44293
rect 25645 44259 25651 44293
rect 25605 44221 25651 44259
rect 25605 44187 25611 44221
rect 25645 44187 25651 44221
rect 25605 44149 25651 44187
rect 25605 44115 25611 44149
rect 25645 44115 25651 44149
rect 25605 44077 25651 44115
rect 25605 44043 25611 44077
rect 25645 44043 25651 44077
rect 25605 44005 25651 44043
rect 25605 43971 25611 44005
rect 25645 43971 25651 44005
rect 25605 43933 25651 43971
rect 25605 43899 25611 43933
rect 25645 43899 25651 43933
rect 25605 43861 25651 43899
rect 25605 43827 25611 43861
rect 25645 43827 25651 43861
rect 25605 43789 25651 43827
rect 25605 43755 25611 43789
rect 25645 43755 25651 43789
rect 25605 43717 25651 43755
rect 25605 43683 25611 43717
rect 25645 43683 25651 43717
rect 25605 43667 25651 43683
rect 26063 44941 26109 44957
rect 26063 44907 26069 44941
rect 26103 44907 26109 44941
rect 26063 44869 26109 44907
rect 26063 44835 26069 44869
rect 26103 44835 26109 44869
rect 26063 44797 26109 44835
rect 26063 44763 26069 44797
rect 26103 44763 26109 44797
rect 26063 44725 26109 44763
rect 26063 44691 26069 44725
rect 26103 44691 26109 44725
rect 26063 44653 26109 44691
rect 26063 44619 26069 44653
rect 26103 44619 26109 44653
rect 26063 44581 26109 44619
rect 26063 44547 26069 44581
rect 26103 44547 26109 44581
rect 26063 44509 26109 44547
rect 26063 44475 26069 44509
rect 26103 44475 26109 44509
rect 26063 44437 26109 44475
rect 26063 44403 26069 44437
rect 26103 44403 26109 44437
rect 26063 44365 26109 44403
rect 26063 44331 26069 44365
rect 26103 44331 26109 44365
rect 26063 44293 26109 44331
rect 26063 44259 26069 44293
rect 26103 44259 26109 44293
rect 26063 44221 26109 44259
rect 26063 44187 26069 44221
rect 26103 44187 26109 44221
rect 26063 44149 26109 44187
rect 26063 44115 26069 44149
rect 26103 44115 26109 44149
rect 26063 44077 26109 44115
rect 26063 44043 26069 44077
rect 26103 44043 26109 44077
rect 26063 44005 26109 44043
rect 26063 43971 26069 44005
rect 26103 43971 26109 44005
rect 26063 43933 26109 43971
rect 26063 43899 26069 43933
rect 26103 43899 26109 43933
rect 26063 43861 26109 43899
rect 26063 43827 26069 43861
rect 26103 43827 26109 43861
rect 26063 43789 26109 43827
rect 26063 43755 26069 43789
rect 26103 43755 26109 43789
rect 26063 43717 26109 43755
rect 26063 43683 26069 43717
rect 26103 43683 26109 43717
rect 26063 43667 26109 43683
rect 26521 44941 26567 44957
rect 26521 44907 26527 44941
rect 26561 44907 26567 44941
rect 26521 44869 26567 44907
rect 26521 44835 26527 44869
rect 26561 44835 26567 44869
rect 26521 44797 26567 44835
rect 26521 44763 26527 44797
rect 26561 44763 26567 44797
rect 26521 44725 26567 44763
rect 26521 44691 26527 44725
rect 26561 44691 26567 44725
rect 26521 44653 26567 44691
rect 26521 44619 26527 44653
rect 26561 44619 26567 44653
rect 26521 44581 26567 44619
rect 26521 44547 26527 44581
rect 26561 44547 26567 44581
rect 26521 44509 26567 44547
rect 26521 44475 26527 44509
rect 26561 44475 26567 44509
rect 26521 44437 26567 44475
rect 26521 44403 26527 44437
rect 26561 44403 26567 44437
rect 26521 44365 26567 44403
rect 26521 44331 26527 44365
rect 26561 44331 26567 44365
rect 26521 44293 26567 44331
rect 26521 44259 26527 44293
rect 26561 44259 26567 44293
rect 26521 44221 26567 44259
rect 26521 44187 26527 44221
rect 26561 44187 26567 44221
rect 26521 44149 26567 44187
rect 26521 44115 26527 44149
rect 26561 44115 26567 44149
rect 26521 44077 26567 44115
rect 26521 44043 26527 44077
rect 26561 44043 26567 44077
rect 26521 44005 26567 44043
rect 26521 43971 26527 44005
rect 26561 43971 26567 44005
rect 26521 43933 26567 43971
rect 26521 43899 26527 43933
rect 26561 43899 26567 43933
rect 26521 43861 26567 43899
rect 26521 43827 26527 43861
rect 26561 43827 26567 43861
rect 26521 43789 26567 43827
rect 26521 43755 26527 43789
rect 26561 43755 26567 43789
rect 26521 43717 26567 43755
rect 26521 43683 26527 43717
rect 26561 43683 26567 43717
rect 26521 43667 26567 43683
rect 26979 44941 27025 44957
rect 26979 44907 26985 44941
rect 27019 44907 27025 44941
rect 26979 44869 27025 44907
rect 26979 44835 26985 44869
rect 27019 44835 27025 44869
rect 26979 44797 27025 44835
rect 26979 44763 26985 44797
rect 27019 44763 27025 44797
rect 26979 44725 27025 44763
rect 26979 44691 26985 44725
rect 27019 44691 27025 44725
rect 26979 44653 27025 44691
rect 26979 44619 26985 44653
rect 27019 44619 27025 44653
rect 26979 44581 27025 44619
rect 26979 44547 26985 44581
rect 27019 44547 27025 44581
rect 26979 44509 27025 44547
rect 26979 44475 26985 44509
rect 27019 44475 27025 44509
rect 26979 44437 27025 44475
rect 26979 44403 26985 44437
rect 27019 44403 27025 44437
rect 26979 44365 27025 44403
rect 26979 44331 26985 44365
rect 27019 44331 27025 44365
rect 26979 44293 27025 44331
rect 26979 44259 26985 44293
rect 27019 44259 27025 44293
rect 26979 44221 27025 44259
rect 26979 44187 26985 44221
rect 27019 44187 27025 44221
rect 26979 44149 27025 44187
rect 26979 44115 26985 44149
rect 27019 44115 27025 44149
rect 26979 44077 27025 44115
rect 26979 44043 26985 44077
rect 27019 44043 27025 44077
rect 26979 44005 27025 44043
rect 26979 43971 26985 44005
rect 27019 43971 27025 44005
rect 26979 43933 27025 43971
rect 26979 43899 26985 43933
rect 27019 43899 27025 43933
rect 26979 43861 27025 43899
rect 26979 43827 26985 43861
rect 27019 43827 27025 43861
rect 26979 43789 27025 43827
rect 26979 43755 26985 43789
rect 27019 43755 27025 43789
rect 26979 43717 27025 43755
rect 26979 43683 26985 43717
rect 27019 43683 27025 43717
rect 26979 43667 27025 43683
rect 27437 44941 27483 44957
rect 27437 44907 27443 44941
rect 27477 44907 27483 44941
rect 27437 44869 27483 44907
rect 27437 44835 27443 44869
rect 27477 44835 27483 44869
rect 27437 44797 27483 44835
rect 27437 44763 27443 44797
rect 27477 44763 27483 44797
rect 27437 44725 27483 44763
rect 27437 44691 27443 44725
rect 27477 44691 27483 44725
rect 27437 44653 27483 44691
rect 27437 44619 27443 44653
rect 27477 44619 27483 44653
rect 27437 44581 27483 44619
rect 27437 44547 27443 44581
rect 27477 44547 27483 44581
rect 27437 44509 27483 44547
rect 27437 44475 27443 44509
rect 27477 44475 27483 44509
rect 27437 44437 27483 44475
rect 27437 44403 27443 44437
rect 27477 44403 27483 44437
rect 27437 44365 27483 44403
rect 27437 44331 27443 44365
rect 27477 44331 27483 44365
rect 27437 44293 27483 44331
rect 27437 44259 27443 44293
rect 27477 44259 27483 44293
rect 27437 44221 27483 44259
rect 27437 44187 27443 44221
rect 27477 44187 27483 44221
rect 27437 44149 27483 44187
rect 27437 44115 27443 44149
rect 27477 44115 27483 44149
rect 27437 44077 27483 44115
rect 27437 44043 27443 44077
rect 27477 44043 27483 44077
rect 27437 44005 27483 44043
rect 27437 43971 27443 44005
rect 27477 43971 27483 44005
rect 27437 43933 27483 43971
rect 27437 43899 27443 43933
rect 27477 43899 27483 43933
rect 27437 43861 27483 43899
rect 27437 43827 27443 43861
rect 27477 43827 27483 43861
rect 27437 43789 27483 43827
rect 27437 43755 27443 43789
rect 27477 43755 27483 43789
rect 27437 43717 27483 43755
rect 27437 43683 27443 43717
rect 27477 43683 27483 43717
rect 27437 43667 27483 43683
rect 27895 44941 27941 44957
rect 27895 44907 27901 44941
rect 27935 44907 27941 44941
rect 27895 44869 27941 44907
rect 27895 44835 27901 44869
rect 27935 44835 27941 44869
rect 27895 44797 27941 44835
rect 27895 44763 27901 44797
rect 27935 44763 27941 44797
rect 27895 44725 27941 44763
rect 27895 44691 27901 44725
rect 27935 44691 27941 44725
rect 27895 44653 27941 44691
rect 27895 44619 27901 44653
rect 27935 44619 27941 44653
rect 27895 44581 27941 44619
rect 27895 44547 27901 44581
rect 27935 44547 27941 44581
rect 27895 44509 27941 44547
rect 27895 44475 27901 44509
rect 27935 44475 27941 44509
rect 27895 44437 27941 44475
rect 27895 44403 27901 44437
rect 27935 44403 27941 44437
rect 27895 44365 27941 44403
rect 27895 44331 27901 44365
rect 27935 44331 27941 44365
rect 27895 44293 27941 44331
rect 27895 44259 27901 44293
rect 27935 44259 27941 44293
rect 27895 44221 27941 44259
rect 27895 44187 27901 44221
rect 27935 44187 27941 44221
rect 27895 44149 27941 44187
rect 27895 44115 27901 44149
rect 27935 44115 27941 44149
rect 27895 44077 27941 44115
rect 27895 44043 27901 44077
rect 27935 44043 27941 44077
rect 27895 44005 27941 44043
rect 27895 43971 27901 44005
rect 27935 43971 27941 44005
rect 27895 43933 27941 43971
rect 27895 43899 27901 43933
rect 27935 43899 27941 43933
rect 27895 43861 27941 43899
rect 27895 43827 27901 43861
rect 27935 43827 27941 43861
rect 27895 43789 27941 43827
rect 27895 43755 27901 43789
rect 27935 43755 27941 43789
rect 27895 43717 27941 43755
rect 27895 43683 27901 43717
rect 27935 43683 27941 43717
rect 27895 43667 27941 43683
rect 28353 44941 28399 44957
rect 28353 44907 28359 44941
rect 28393 44907 28399 44941
rect 28353 44869 28399 44907
rect 28353 44835 28359 44869
rect 28393 44835 28399 44869
rect 28353 44797 28399 44835
rect 28353 44763 28359 44797
rect 28393 44763 28399 44797
rect 28353 44725 28399 44763
rect 28353 44691 28359 44725
rect 28393 44691 28399 44725
rect 28353 44653 28399 44691
rect 28353 44619 28359 44653
rect 28393 44619 28399 44653
rect 28353 44581 28399 44619
rect 28353 44547 28359 44581
rect 28393 44547 28399 44581
rect 28353 44509 28399 44547
rect 28353 44475 28359 44509
rect 28393 44475 28399 44509
rect 28353 44437 28399 44475
rect 28353 44403 28359 44437
rect 28393 44403 28399 44437
rect 28353 44365 28399 44403
rect 28353 44331 28359 44365
rect 28393 44331 28399 44365
rect 28353 44293 28399 44331
rect 28353 44259 28359 44293
rect 28393 44259 28399 44293
rect 28353 44221 28399 44259
rect 28353 44187 28359 44221
rect 28393 44187 28399 44221
rect 28353 44149 28399 44187
rect 28353 44115 28359 44149
rect 28393 44115 28399 44149
rect 28353 44077 28399 44115
rect 28353 44043 28359 44077
rect 28393 44043 28399 44077
rect 28353 44005 28399 44043
rect 28353 43971 28359 44005
rect 28393 43971 28399 44005
rect 28353 43933 28399 43971
rect 28353 43899 28359 43933
rect 28393 43899 28399 43933
rect 28353 43861 28399 43899
rect 28353 43827 28359 43861
rect 28393 43827 28399 43861
rect 28353 43789 28399 43827
rect 28353 43755 28359 43789
rect 28393 43755 28399 43789
rect 28353 43717 28399 43755
rect 28353 43683 28359 43717
rect 28393 43683 28399 43717
rect 28353 43667 28399 43683
rect 28811 44941 28857 44957
rect 28811 44907 28817 44941
rect 28851 44907 28857 44941
rect 28811 44869 28857 44907
rect 28811 44835 28817 44869
rect 28851 44835 28857 44869
rect 28811 44797 28857 44835
rect 28811 44763 28817 44797
rect 28851 44763 28857 44797
rect 28811 44725 28857 44763
rect 28811 44691 28817 44725
rect 28851 44691 28857 44725
rect 28811 44653 28857 44691
rect 28811 44619 28817 44653
rect 28851 44619 28857 44653
rect 28811 44581 28857 44619
rect 28811 44547 28817 44581
rect 28851 44547 28857 44581
rect 28811 44509 28857 44547
rect 28811 44475 28817 44509
rect 28851 44475 28857 44509
rect 28811 44437 28857 44475
rect 28811 44403 28817 44437
rect 28851 44403 28857 44437
rect 28811 44365 28857 44403
rect 28811 44331 28817 44365
rect 28851 44331 28857 44365
rect 28811 44293 28857 44331
rect 28811 44259 28817 44293
rect 28851 44259 28857 44293
rect 28811 44221 28857 44259
rect 28811 44187 28817 44221
rect 28851 44187 28857 44221
rect 28811 44149 28857 44187
rect 28811 44115 28817 44149
rect 28851 44115 28857 44149
rect 28811 44077 28857 44115
rect 28811 44043 28817 44077
rect 28851 44043 28857 44077
rect 28811 44005 28857 44043
rect 28811 43971 28817 44005
rect 28851 43971 28857 44005
rect 28811 43933 28857 43971
rect 28811 43899 28817 43933
rect 28851 43899 28857 43933
rect 28811 43861 28857 43899
rect 28811 43827 28817 43861
rect 28851 43827 28857 43861
rect 28811 43789 28857 43827
rect 28811 43755 28817 43789
rect 28851 43755 28857 43789
rect 28811 43717 28857 43755
rect 28811 43683 28817 43717
rect 28851 43683 28857 43717
rect 28811 43667 28857 43683
rect 29269 44941 29315 44957
rect 29269 44907 29275 44941
rect 29309 44907 29315 44941
rect 29269 44869 29315 44907
rect 29269 44835 29275 44869
rect 29309 44835 29315 44869
rect 29269 44797 29315 44835
rect 29269 44763 29275 44797
rect 29309 44763 29315 44797
rect 29269 44725 29315 44763
rect 29269 44691 29275 44725
rect 29309 44691 29315 44725
rect 29269 44653 29315 44691
rect 29269 44619 29275 44653
rect 29309 44619 29315 44653
rect 29269 44581 29315 44619
rect 29269 44547 29275 44581
rect 29309 44547 29315 44581
rect 29269 44509 29315 44547
rect 29269 44475 29275 44509
rect 29309 44475 29315 44509
rect 29269 44437 29315 44475
rect 29269 44403 29275 44437
rect 29309 44403 29315 44437
rect 29269 44365 29315 44403
rect 29269 44331 29275 44365
rect 29309 44331 29315 44365
rect 29269 44293 29315 44331
rect 29269 44259 29275 44293
rect 29309 44259 29315 44293
rect 29269 44221 29315 44259
rect 29269 44187 29275 44221
rect 29309 44187 29315 44221
rect 29269 44149 29315 44187
rect 29269 44115 29275 44149
rect 29309 44115 29315 44149
rect 29269 44077 29315 44115
rect 29269 44043 29275 44077
rect 29309 44043 29315 44077
rect 29269 44005 29315 44043
rect 29269 43971 29275 44005
rect 29309 43971 29315 44005
rect 29269 43933 29315 43971
rect 29269 43899 29275 43933
rect 29309 43899 29315 43933
rect 29269 43861 29315 43899
rect 29269 43827 29275 43861
rect 29309 43827 29315 43861
rect 29269 43789 29315 43827
rect 29269 43755 29275 43789
rect 29309 43755 29315 43789
rect 29269 43717 29315 43755
rect 29269 43683 29275 43717
rect 29309 43683 29315 43717
rect 29269 43667 29315 43683
rect 29727 44941 29773 44957
rect 29727 44907 29733 44941
rect 29767 44907 29773 44941
rect 29727 44869 29773 44907
rect 29727 44835 29733 44869
rect 29767 44835 29773 44869
rect 29727 44797 29773 44835
rect 29727 44763 29733 44797
rect 29767 44763 29773 44797
rect 29727 44725 29773 44763
rect 29727 44691 29733 44725
rect 29767 44691 29773 44725
rect 29727 44653 29773 44691
rect 29727 44619 29733 44653
rect 29767 44619 29773 44653
rect 29727 44581 29773 44619
rect 29727 44547 29733 44581
rect 29767 44547 29773 44581
rect 29727 44509 29773 44547
rect 29727 44475 29733 44509
rect 29767 44475 29773 44509
rect 29727 44437 29773 44475
rect 29727 44403 29733 44437
rect 29767 44403 29773 44437
rect 29727 44365 29773 44403
rect 29727 44331 29733 44365
rect 29767 44331 29773 44365
rect 29727 44293 29773 44331
rect 29727 44259 29733 44293
rect 29767 44259 29773 44293
rect 29727 44221 29773 44259
rect 29727 44187 29733 44221
rect 29767 44187 29773 44221
rect 29727 44149 29773 44187
rect 29727 44115 29733 44149
rect 29767 44115 29773 44149
rect 29727 44077 29773 44115
rect 29727 44043 29733 44077
rect 29767 44043 29773 44077
rect 29727 44005 29773 44043
rect 29727 43971 29733 44005
rect 29767 43971 29773 44005
rect 29727 43933 29773 43971
rect 29727 43899 29733 43933
rect 29767 43899 29773 43933
rect 29727 43861 29773 43899
rect 29727 43827 29733 43861
rect 29767 43827 29773 43861
rect 29727 43789 29773 43827
rect 29727 43755 29733 43789
rect 29767 43755 29773 43789
rect 29727 43717 29773 43755
rect 29727 43683 29733 43717
rect 29767 43683 29773 43717
rect 29727 43667 29773 43683
rect 30185 44941 30231 44957
rect 30185 44907 30191 44941
rect 30225 44907 30231 44941
rect 30185 44869 30231 44907
rect 30185 44835 30191 44869
rect 30225 44835 30231 44869
rect 30185 44797 30231 44835
rect 30185 44763 30191 44797
rect 30225 44763 30231 44797
rect 30185 44725 30231 44763
rect 30185 44691 30191 44725
rect 30225 44691 30231 44725
rect 30185 44653 30231 44691
rect 30185 44619 30191 44653
rect 30225 44619 30231 44653
rect 30185 44581 30231 44619
rect 30185 44547 30191 44581
rect 30225 44547 30231 44581
rect 30185 44509 30231 44547
rect 30185 44475 30191 44509
rect 30225 44475 30231 44509
rect 30185 44437 30231 44475
rect 30185 44403 30191 44437
rect 30225 44403 30231 44437
rect 30185 44365 30231 44403
rect 30185 44331 30191 44365
rect 30225 44331 30231 44365
rect 30185 44293 30231 44331
rect 30185 44259 30191 44293
rect 30225 44259 30231 44293
rect 30185 44221 30231 44259
rect 30185 44187 30191 44221
rect 30225 44187 30231 44221
rect 30185 44149 30231 44187
rect 30185 44115 30191 44149
rect 30225 44115 30231 44149
rect 30185 44077 30231 44115
rect 30185 44043 30191 44077
rect 30225 44043 30231 44077
rect 30185 44005 30231 44043
rect 30185 43971 30191 44005
rect 30225 43971 30231 44005
rect 30185 43933 30231 43971
rect 30185 43899 30191 43933
rect 30225 43899 30231 43933
rect 30185 43861 30231 43899
rect 30185 43827 30191 43861
rect 30225 43827 30231 43861
rect 30185 43789 30231 43827
rect 30185 43755 30191 43789
rect 30225 43755 30231 43789
rect 30185 43717 30231 43755
rect 30185 43683 30191 43717
rect 30225 43683 30231 43717
rect 30185 43667 30231 43683
rect 30643 44941 30689 44957
rect 30643 44907 30649 44941
rect 30683 44907 30689 44941
rect 30643 44869 30689 44907
rect 30643 44835 30649 44869
rect 30683 44835 30689 44869
rect 30643 44797 30689 44835
rect 30643 44763 30649 44797
rect 30683 44763 30689 44797
rect 30643 44725 30689 44763
rect 30643 44691 30649 44725
rect 30683 44691 30689 44725
rect 30643 44653 30689 44691
rect 30643 44619 30649 44653
rect 30683 44619 30689 44653
rect 30643 44581 30689 44619
rect 30643 44547 30649 44581
rect 30683 44547 30689 44581
rect 30643 44509 30689 44547
rect 30643 44475 30649 44509
rect 30683 44475 30689 44509
rect 30643 44437 30689 44475
rect 30643 44403 30649 44437
rect 30683 44403 30689 44437
rect 30643 44365 30689 44403
rect 30643 44331 30649 44365
rect 30683 44331 30689 44365
rect 30643 44293 30689 44331
rect 30643 44259 30649 44293
rect 30683 44259 30689 44293
rect 30643 44221 30689 44259
rect 30643 44187 30649 44221
rect 30683 44187 30689 44221
rect 30643 44149 30689 44187
rect 30643 44115 30649 44149
rect 30683 44115 30689 44149
rect 30643 44077 30689 44115
rect 30643 44043 30649 44077
rect 30683 44043 30689 44077
rect 30643 44005 30689 44043
rect 30643 43971 30649 44005
rect 30683 43971 30689 44005
rect 30643 43933 30689 43971
rect 30643 43899 30649 43933
rect 30683 43899 30689 43933
rect 30643 43861 30689 43899
rect 30643 43827 30649 43861
rect 30683 43827 30689 43861
rect 30643 43789 30689 43827
rect 30643 43755 30649 43789
rect 30683 43755 30689 43789
rect 30643 43717 30689 43755
rect 30643 43683 30649 43717
rect 30683 43683 30689 43717
rect 30643 43667 30689 43683
rect 31101 44941 31147 44957
rect 31101 44907 31107 44941
rect 31141 44907 31147 44941
rect 31101 44869 31147 44907
rect 31101 44835 31107 44869
rect 31141 44835 31147 44869
rect 31101 44797 31147 44835
rect 31101 44763 31107 44797
rect 31141 44763 31147 44797
rect 31101 44725 31147 44763
rect 31101 44691 31107 44725
rect 31141 44691 31147 44725
rect 31101 44653 31147 44691
rect 31101 44619 31107 44653
rect 31141 44619 31147 44653
rect 31101 44581 31147 44619
rect 31101 44547 31107 44581
rect 31141 44547 31147 44581
rect 31101 44509 31147 44547
rect 31101 44475 31107 44509
rect 31141 44475 31147 44509
rect 31101 44437 31147 44475
rect 31101 44403 31107 44437
rect 31141 44403 31147 44437
rect 31101 44365 31147 44403
rect 31101 44331 31107 44365
rect 31141 44331 31147 44365
rect 31101 44293 31147 44331
rect 31101 44259 31107 44293
rect 31141 44259 31147 44293
rect 31101 44221 31147 44259
rect 31101 44187 31107 44221
rect 31141 44187 31147 44221
rect 31101 44149 31147 44187
rect 31101 44115 31107 44149
rect 31141 44115 31147 44149
rect 31101 44077 31147 44115
rect 31101 44043 31107 44077
rect 31141 44043 31147 44077
rect 31101 44005 31147 44043
rect 31101 43971 31107 44005
rect 31141 43971 31147 44005
rect 31101 43933 31147 43971
rect 31101 43899 31107 43933
rect 31141 43899 31147 43933
rect 31101 43861 31147 43899
rect 31101 43827 31107 43861
rect 31141 43827 31147 43861
rect 31101 43789 31147 43827
rect 31101 43755 31107 43789
rect 31141 43755 31147 43789
rect 31101 43717 31147 43755
rect 31101 43683 31107 43717
rect 31141 43683 31147 43717
rect 31101 43667 31147 43683
rect 31559 44941 31605 44957
rect 31559 44907 31565 44941
rect 31599 44907 31605 44941
rect 31559 44869 31605 44907
rect 31559 44835 31565 44869
rect 31599 44835 31605 44869
rect 31559 44797 31605 44835
rect 31559 44763 31565 44797
rect 31599 44763 31605 44797
rect 31559 44725 31605 44763
rect 31559 44691 31565 44725
rect 31599 44691 31605 44725
rect 31559 44653 31605 44691
rect 31559 44619 31565 44653
rect 31599 44619 31605 44653
rect 31559 44581 31605 44619
rect 31559 44547 31565 44581
rect 31599 44547 31605 44581
rect 31559 44509 31605 44547
rect 31559 44475 31565 44509
rect 31599 44475 31605 44509
rect 31559 44437 31605 44475
rect 31559 44403 31565 44437
rect 31599 44403 31605 44437
rect 31559 44365 31605 44403
rect 31559 44331 31565 44365
rect 31599 44331 31605 44365
rect 31559 44293 31605 44331
rect 31559 44259 31565 44293
rect 31599 44259 31605 44293
rect 31559 44221 31605 44259
rect 31559 44187 31565 44221
rect 31599 44187 31605 44221
rect 31559 44149 31605 44187
rect 31559 44115 31565 44149
rect 31599 44115 31605 44149
rect 31559 44077 31605 44115
rect 31559 44043 31565 44077
rect 31599 44043 31605 44077
rect 31559 44005 31605 44043
rect 31559 43971 31565 44005
rect 31599 43971 31605 44005
rect 31559 43933 31605 43971
rect 31559 43899 31565 43933
rect 31599 43899 31605 43933
rect 31559 43861 31605 43899
rect 31559 43827 31565 43861
rect 31599 43827 31605 43861
rect 31559 43789 31605 43827
rect 31559 43755 31565 43789
rect 31599 43755 31605 43789
rect 31559 43717 31605 43755
rect 31559 43683 31565 43717
rect 31599 43683 31605 43717
rect 31559 43667 31605 43683
rect 32017 44941 32063 44957
rect 32017 44907 32023 44941
rect 32057 44907 32063 44941
rect 32017 44869 32063 44907
rect 32017 44835 32023 44869
rect 32057 44835 32063 44869
rect 32017 44797 32063 44835
rect 32017 44763 32023 44797
rect 32057 44763 32063 44797
rect 32017 44725 32063 44763
rect 32017 44691 32023 44725
rect 32057 44691 32063 44725
rect 32017 44653 32063 44691
rect 32017 44619 32023 44653
rect 32057 44619 32063 44653
rect 32017 44581 32063 44619
rect 32017 44547 32023 44581
rect 32057 44547 32063 44581
rect 32017 44509 32063 44547
rect 32017 44475 32023 44509
rect 32057 44475 32063 44509
rect 32017 44437 32063 44475
rect 32017 44403 32023 44437
rect 32057 44403 32063 44437
rect 32017 44365 32063 44403
rect 32017 44331 32023 44365
rect 32057 44331 32063 44365
rect 32017 44293 32063 44331
rect 32017 44259 32023 44293
rect 32057 44259 32063 44293
rect 32017 44221 32063 44259
rect 32017 44187 32023 44221
rect 32057 44187 32063 44221
rect 32017 44149 32063 44187
rect 32017 44115 32023 44149
rect 32057 44115 32063 44149
rect 32017 44077 32063 44115
rect 32017 44043 32023 44077
rect 32057 44043 32063 44077
rect 32017 44005 32063 44043
rect 32017 43971 32023 44005
rect 32057 43971 32063 44005
rect 32017 43933 32063 43971
rect 32017 43899 32023 43933
rect 32057 43899 32063 43933
rect 32017 43861 32063 43899
rect 32017 43827 32023 43861
rect 32057 43827 32063 43861
rect 32017 43789 32063 43827
rect 32017 43755 32023 43789
rect 32057 43755 32063 43789
rect 32017 43717 32063 43755
rect 32017 43683 32023 43717
rect 32057 43683 32063 43717
rect 32017 43667 32063 43683
rect 32475 44941 32521 44957
rect 32475 44907 32481 44941
rect 32515 44907 32521 44941
rect 32475 44869 32521 44907
rect 32475 44835 32481 44869
rect 32515 44835 32521 44869
rect 32475 44797 32521 44835
rect 32475 44763 32481 44797
rect 32515 44763 32521 44797
rect 32475 44725 32521 44763
rect 32475 44691 32481 44725
rect 32515 44691 32521 44725
rect 32475 44653 32521 44691
rect 32475 44619 32481 44653
rect 32515 44619 32521 44653
rect 32475 44581 32521 44619
rect 32475 44547 32481 44581
rect 32515 44547 32521 44581
rect 32475 44509 32521 44547
rect 32475 44475 32481 44509
rect 32515 44475 32521 44509
rect 32475 44437 32521 44475
rect 32475 44403 32481 44437
rect 32515 44403 32521 44437
rect 32475 44365 32521 44403
rect 32475 44331 32481 44365
rect 32515 44331 32521 44365
rect 32475 44293 32521 44331
rect 32475 44259 32481 44293
rect 32515 44259 32521 44293
rect 32475 44221 32521 44259
rect 32475 44187 32481 44221
rect 32515 44187 32521 44221
rect 32475 44149 32521 44187
rect 32475 44115 32481 44149
rect 32515 44115 32521 44149
rect 32475 44077 32521 44115
rect 32475 44043 32481 44077
rect 32515 44043 32521 44077
rect 32475 44005 32521 44043
rect 32475 43971 32481 44005
rect 32515 43971 32521 44005
rect 32475 43933 32521 43971
rect 32475 43899 32481 43933
rect 32515 43899 32521 43933
rect 32475 43861 32521 43899
rect 32475 43827 32481 43861
rect 32515 43827 32521 43861
rect 32475 43789 32521 43827
rect 32475 43755 32481 43789
rect 32515 43755 32521 43789
rect 32475 43717 32521 43755
rect 32475 43683 32481 43717
rect 32515 43683 32521 43717
rect 32475 43667 32521 43683
rect 32933 44941 32979 44957
rect 32933 44907 32939 44941
rect 32973 44907 32979 44941
rect 32933 44869 32979 44907
rect 32933 44835 32939 44869
rect 32973 44835 32979 44869
rect 32933 44797 32979 44835
rect 32933 44763 32939 44797
rect 32973 44763 32979 44797
rect 32933 44725 32979 44763
rect 32933 44691 32939 44725
rect 32973 44691 32979 44725
rect 32933 44653 32979 44691
rect 32933 44619 32939 44653
rect 32973 44619 32979 44653
rect 32933 44581 32979 44619
rect 32933 44547 32939 44581
rect 32973 44547 32979 44581
rect 32933 44509 32979 44547
rect 32933 44475 32939 44509
rect 32973 44475 32979 44509
rect 32933 44437 32979 44475
rect 32933 44403 32939 44437
rect 32973 44403 32979 44437
rect 32933 44365 32979 44403
rect 32933 44331 32939 44365
rect 32973 44331 32979 44365
rect 32933 44293 32979 44331
rect 32933 44259 32939 44293
rect 32973 44259 32979 44293
rect 32933 44221 32979 44259
rect 32933 44187 32939 44221
rect 32973 44187 32979 44221
rect 32933 44149 32979 44187
rect 32933 44115 32939 44149
rect 32973 44115 32979 44149
rect 32933 44077 32979 44115
rect 32933 44043 32939 44077
rect 32973 44043 32979 44077
rect 32933 44005 32979 44043
rect 32933 43971 32939 44005
rect 32973 43971 32979 44005
rect 32933 43933 32979 43971
rect 32933 43899 32939 43933
rect 32973 43899 32979 43933
rect 32933 43861 32979 43899
rect 32933 43827 32939 43861
rect 32973 43827 32979 43861
rect 32933 43789 32979 43827
rect 32933 43755 32939 43789
rect 32973 43755 32979 43789
rect 32933 43717 32979 43755
rect 32933 43683 32939 43717
rect 32973 43683 32979 43717
rect 32933 43667 32979 43683
rect 33391 44941 33437 44957
rect 33391 44907 33397 44941
rect 33431 44907 33437 44941
rect 33391 44869 33437 44907
rect 33391 44835 33397 44869
rect 33431 44835 33437 44869
rect 33391 44797 33437 44835
rect 33391 44763 33397 44797
rect 33431 44763 33437 44797
rect 33391 44725 33437 44763
rect 33391 44691 33397 44725
rect 33431 44691 33437 44725
rect 33391 44653 33437 44691
rect 33391 44619 33397 44653
rect 33431 44619 33437 44653
rect 33391 44581 33437 44619
rect 33391 44547 33397 44581
rect 33431 44547 33437 44581
rect 33391 44509 33437 44547
rect 33391 44475 33397 44509
rect 33431 44475 33437 44509
rect 33391 44437 33437 44475
rect 33391 44403 33397 44437
rect 33431 44403 33437 44437
rect 33391 44365 33437 44403
rect 33391 44331 33397 44365
rect 33431 44331 33437 44365
rect 33391 44293 33437 44331
rect 33391 44259 33397 44293
rect 33431 44259 33437 44293
rect 33391 44221 33437 44259
rect 33391 44187 33397 44221
rect 33431 44187 33437 44221
rect 33391 44149 33437 44187
rect 33391 44115 33397 44149
rect 33431 44115 33437 44149
rect 33391 44077 33437 44115
rect 33391 44043 33397 44077
rect 33431 44043 33437 44077
rect 33391 44005 33437 44043
rect 33391 43971 33397 44005
rect 33431 43971 33437 44005
rect 33391 43933 33437 43971
rect 33391 43899 33397 43933
rect 33431 43899 33437 43933
rect 33391 43861 33437 43899
rect 33391 43827 33397 43861
rect 33431 43827 33437 43861
rect 33391 43789 33437 43827
rect 33391 43755 33397 43789
rect 33431 43755 33437 43789
rect 33391 43717 33437 43755
rect 33391 43683 33397 43717
rect 33431 43683 33437 43717
rect 33391 43667 33437 43683
rect 33849 44941 33895 44957
rect 33849 44907 33855 44941
rect 33889 44907 33895 44941
rect 33849 44869 33895 44907
rect 33849 44835 33855 44869
rect 33889 44835 33895 44869
rect 33849 44797 33895 44835
rect 33849 44763 33855 44797
rect 33889 44763 33895 44797
rect 33849 44725 33895 44763
rect 33849 44691 33855 44725
rect 33889 44691 33895 44725
rect 33849 44653 33895 44691
rect 33849 44619 33855 44653
rect 33889 44619 33895 44653
rect 33849 44581 33895 44619
rect 33849 44547 33855 44581
rect 33889 44547 33895 44581
rect 33849 44509 33895 44547
rect 33849 44475 33855 44509
rect 33889 44475 33895 44509
rect 33849 44437 33895 44475
rect 33849 44403 33855 44437
rect 33889 44403 33895 44437
rect 33849 44365 33895 44403
rect 33849 44331 33855 44365
rect 33889 44331 33895 44365
rect 33849 44293 33895 44331
rect 33849 44259 33855 44293
rect 33889 44259 33895 44293
rect 33849 44221 33895 44259
rect 33849 44187 33855 44221
rect 33889 44187 33895 44221
rect 33849 44149 33895 44187
rect 33849 44115 33855 44149
rect 33889 44115 33895 44149
rect 33849 44077 33895 44115
rect 33849 44043 33855 44077
rect 33889 44043 33895 44077
rect 33849 44005 33895 44043
rect 33849 43971 33855 44005
rect 33889 43971 33895 44005
rect 33849 43933 33895 43971
rect 33849 43899 33855 43933
rect 33889 43899 33895 43933
rect 33849 43861 33895 43899
rect 33849 43827 33855 43861
rect 33889 43827 33895 43861
rect 33849 43789 33895 43827
rect 33849 43755 33855 43789
rect 33889 43755 33895 43789
rect 33849 43717 33895 43755
rect 33849 43683 33855 43717
rect 33889 43683 33895 43717
rect 33849 43667 33895 43683
rect 34307 44941 34353 44957
rect 34307 44907 34313 44941
rect 34347 44907 34353 44941
rect 34307 44869 34353 44907
rect 34307 44835 34313 44869
rect 34347 44835 34353 44869
rect 34307 44797 34353 44835
rect 34307 44763 34313 44797
rect 34347 44763 34353 44797
rect 34307 44725 34353 44763
rect 34307 44691 34313 44725
rect 34347 44691 34353 44725
rect 34307 44653 34353 44691
rect 34307 44619 34313 44653
rect 34347 44619 34353 44653
rect 34307 44581 34353 44619
rect 34307 44547 34313 44581
rect 34347 44547 34353 44581
rect 34307 44509 34353 44547
rect 34307 44475 34313 44509
rect 34347 44475 34353 44509
rect 34307 44437 34353 44475
rect 34307 44403 34313 44437
rect 34347 44403 34353 44437
rect 34307 44365 34353 44403
rect 34307 44331 34313 44365
rect 34347 44331 34353 44365
rect 34307 44293 34353 44331
rect 34307 44259 34313 44293
rect 34347 44259 34353 44293
rect 34307 44221 34353 44259
rect 34307 44187 34313 44221
rect 34347 44187 34353 44221
rect 34307 44149 34353 44187
rect 34307 44115 34313 44149
rect 34347 44115 34353 44149
rect 34307 44077 34353 44115
rect 34307 44043 34313 44077
rect 34347 44043 34353 44077
rect 34307 44005 34353 44043
rect 34307 43971 34313 44005
rect 34347 43971 34353 44005
rect 34307 43933 34353 43971
rect 34307 43899 34313 43933
rect 34347 43899 34353 43933
rect 34307 43861 34353 43899
rect 34307 43827 34313 43861
rect 34347 43827 34353 43861
rect 34307 43789 34353 43827
rect 34307 43755 34313 43789
rect 34347 43755 34353 43789
rect 34307 43717 34353 43755
rect 34307 43683 34313 43717
rect 34347 43683 34353 43717
rect 34307 43667 34353 43683
rect 34765 44941 34811 44957
rect 34765 44907 34771 44941
rect 34805 44907 34811 44941
rect 34765 44869 34811 44907
rect 34765 44835 34771 44869
rect 34805 44835 34811 44869
rect 34765 44797 34811 44835
rect 34765 44763 34771 44797
rect 34805 44763 34811 44797
rect 34765 44725 34811 44763
rect 34765 44691 34771 44725
rect 34805 44691 34811 44725
rect 34765 44653 34811 44691
rect 34765 44619 34771 44653
rect 34805 44619 34811 44653
rect 34765 44581 34811 44619
rect 34765 44547 34771 44581
rect 34805 44547 34811 44581
rect 34765 44509 34811 44547
rect 34765 44475 34771 44509
rect 34805 44475 34811 44509
rect 34765 44437 34811 44475
rect 34765 44403 34771 44437
rect 34805 44403 34811 44437
rect 34765 44365 34811 44403
rect 34765 44331 34771 44365
rect 34805 44331 34811 44365
rect 34765 44293 34811 44331
rect 34765 44259 34771 44293
rect 34805 44259 34811 44293
rect 34765 44221 34811 44259
rect 34765 44187 34771 44221
rect 34805 44187 34811 44221
rect 34765 44149 34811 44187
rect 34765 44115 34771 44149
rect 34805 44115 34811 44149
rect 34765 44077 34811 44115
rect 34765 44043 34771 44077
rect 34805 44043 34811 44077
rect 34765 44005 34811 44043
rect 34765 43971 34771 44005
rect 34805 43971 34811 44005
rect 34765 43933 34811 43971
rect 34765 43899 34771 43933
rect 34805 43899 34811 43933
rect 34765 43861 34811 43899
rect 34765 43827 34771 43861
rect 34805 43827 34811 43861
rect 34765 43789 34811 43827
rect 34765 43755 34771 43789
rect 34805 43755 34811 43789
rect 34765 43717 34811 43755
rect 34765 43683 34771 43717
rect 34805 43683 34811 43717
rect 34765 43667 34811 43683
rect 35223 44941 35269 44957
rect 35223 44907 35229 44941
rect 35263 44907 35269 44941
rect 35223 44869 35269 44907
rect 35223 44835 35229 44869
rect 35263 44835 35269 44869
rect 35223 44797 35269 44835
rect 35223 44763 35229 44797
rect 35263 44763 35269 44797
rect 35223 44725 35269 44763
rect 35223 44691 35229 44725
rect 35263 44691 35269 44725
rect 35223 44653 35269 44691
rect 35223 44619 35229 44653
rect 35263 44619 35269 44653
rect 35223 44581 35269 44619
rect 35223 44547 35229 44581
rect 35263 44547 35269 44581
rect 35223 44509 35269 44547
rect 35223 44475 35229 44509
rect 35263 44475 35269 44509
rect 35223 44437 35269 44475
rect 35223 44403 35229 44437
rect 35263 44403 35269 44437
rect 35223 44365 35269 44403
rect 35223 44331 35229 44365
rect 35263 44331 35269 44365
rect 35223 44293 35269 44331
rect 35223 44259 35229 44293
rect 35263 44259 35269 44293
rect 35223 44221 35269 44259
rect 35223 44187 35229 44221
rect 35263 44187 35269 44221
rect 35223 44149 35269 44187
rect 35223 44115 35229 44149
rect 35263 44115 35269 44149
rect 35223 44077 35269 44115
rect 35223 44043 35229 44077
rect 35263 44043 35269 44077
rect 35223 44005 35269 44043
rect 35223 43971 35229 44005
rect 35263 43971 35269 44005
rect 35223 43933 35269 43971
rect 35223 43899 35229 43933
rect 35263 43899 35269 43933
rect 35223 43861 35269 43899
rect 35223 43827 35229 43861
rect 35263 43827 35269 43861
rect 35223 43789 35269 43827
rect 35223 43755 35229 43789
rect 35263 43755 35269 43789
rect 35223 43717 35269 43755
rect 35223 43683 35229 43717
rect 35263 43683 35269 43717
rect 35223 43667 35269 43683
rect 35681 44941 35727 44957
rect 35681 44907 35687 44941
rect 35721 44907 35727 44941
rect 35681 44869 35727 44907
rect 35681 44835 35687 44869
rect 35721 44835 35727 44869
rect 35681 44797 35727 44835
rect 35681 44763 35687 44797
rect 35721 44763 35727 44797
rect 35681 44725 35727 44763
rect 35681 44691 35687 44725
rect 35721 44691 35727 44725
rect 35681 44653 35727 44691
rect 35681 44619 35687 44653
rect 35721 44619 35727 44653
rect 35681 44581 35727 44619
rect 35681 44547 35687 44581
rect 35721 44547 35727 44581
rect 35681 44509 35727 44547
rect 35681 44475 35687 44509
rect 35721 44475 35727 44509
rect 35681 44437 35727 44475
rect 35681 44403 35687 44437
rect 35721 44403 35727 44437
rect 35681 44365 35727 44403
rect 35681 44331 35687 44365
rect 35721 44331 35727 44365
rect 35681 44293 35727 44331
rect 35681 44259 35687 44293
rect 35721 44259 35727 44293
rect 35681 44221 35727 44259
rect 35681 44187 35687 44221
rect 35721 44187 35727 44221
rect 35681 44149 35727 44187
rect 35681 44115 35687 44149
rect 35721 44115 35727 44149
rect 35681 44077 35727 44115
rect 35681 44043 35687 44077
rect 35721 44043 35727 44077
rect 35681 44005 35727 44043
rect 35681 43971 35687 44005
rect 35721 43971 35727 44005
rect 35681 43933 35727 43971
rect 35681 43899 35687 43933
rect 35721 43899 35727 43933
rect 35681 43861 35727 43899
rect 35681 43827 35687 43861
rect 35721 43827 35727 43861
rect 35681 43789 35727 43827
rect 35681 43755 35687 43789
rect 35721 43755 35727 43789
rect 35681 43717 35727 43755
rect 35681 43683 35687 43717
rect 35721 43683 35727 43717
rect 35681 43667 35727 43683
rect 36139 44941 36185 44957
rect 36139 44907 36145 44941
rect 36179 44907 36185 44941
rect 36139 44869 36185 44907
rect 36139 44835 36145 44869
rect 36179 44835 36185 44869
rect 36139 44797 36185 44835
rect 36139 44763 36145 44797
rect 36179 44763 36185 44797
rect 36139 44725 36185 44763
rect 36139 44691 36145 44725
rect 36179 44691 36185 44725
rect 36139 44653 36185 44691
rect 36139 44619 36145 44653
rect 36179 44619 36185 44653
rect 36139 44581 36185 44619
rect 36139 44547 36145 44581
rect 36179 44547 36185 44581
rect 36139 44509 36185 44547
rect 36139 44475 36145 44509
rect 36179 44475 36185 44509
rect 36139 44437 36185 44475
rect 36139 44403 36145 44437
rect 36179 44403 36185 44437
rect 36139 44365 36185 44403
rect 36139 44331 36145 44365
rect 36179 44331 36185 44365
rect 36139 44293 36185 44331
rect 36139 44259 36145 44293
rect 36179 44259 36185 44293
rect 36139 44221 36185 44259
rect 36139 44187 36145 44221
rect 36179 44187 36185 44221
rect 36139 44149 36185 44187
rect 36139 44115 36145 44149
rect 36179 44115 36185 44149
rect 36139 44077 36185 44115
rect 36139 44043 36145 44077
rect 36179 44043 36185 44077
rect 36139 44005 36185 44043
rect 36139 43971 36145 44005
rect 36179 43971 36185 44005
rect 36139 43933 36185 43971
rect 36139 43899 36145 43933
rect 36179 43899 36185 43933
rect 36139 43861 36185 43899
rect 36139 43827 36145 43861
rect 36179 43827 36185 43861
rect 36139 43789 36185 43827
rect 36139 43755 36145 43789
rect 36179 43755 36185 43789
rect 36139 43717 36185 43755
rect 36139 43683 36145 43717
rect 36179 43683 36185 43717
rect 36139 43667 36185 43683
rect 36597 44941 36643 44957
rect 36597 44907 36603 44941
rect 36637 44907 36643 44941
rect 36597 44869 36643 44907
rect 36597 44835 36603 44869
rect 36637 44835 36643 44869
rect 36597 44797 36643 44835
rect 36597 44763 36603 44797
rect 36637 44763 36643 44797
rect 36597 44725 36643 44763
rect 36597 44691 36603 44725
rect 36637 44691 36643 44725
rect 36597 44653 36643 44691
rect 36597 44619 36603 44653
rect 36637 44619 36643 44653
rect 36597 44581 36643 44619
rect 36597 44547 36603 44581
rect 36637 44547 36643 44581
rect 36597 44509 36643 44547
rect 36597 44475 36603 44509
rect 36637 44475 36643 44509
rect 36597 44437 36643 44475
rect 36597 44403 36603 44437
rect 36637 44403 36643 44437
rect 36597 44365 36643 44403
rect 36597 44331 36603 44365
rect 36637 44331 36643 44365
rect 36597 44293 36643 44331
rect 36597 44259 36603 44293
rect 36637 44259 36643 44293
rect 36597 44221 36643 44259
rect 36597 44187 36603 44221
rect 36637 44187 36643 44221
rect 36597 44149 36643 44187
rect 36597 44115 36603 44149
rect 36637 44115 36643 44149
rect 36597 44077 36643 44115
rect 36597 44043 36603 44077
rect 36637 44043 36643 44077
rect 36597 44005 36643 44043
rect 36597 43971 36603 44005
rect 36637 43971 36643 44005
rect 36597 43933 36643 43971
rect 36597 43899 36603 43933
rect 36637 43899 36643 43933
rect 36597 43861 36643 43899
rect 36597 43827 36603 43861
rect 36637 43827 36643 43861
rect 36597 43789 36643 43827
rect 36597 43755 36603 43789
rect 36637 43755 36643 43789
rect 36597 43717 36643 43755
rect 36597 43683 36603 43717
rect 36637 43683 36643 43717
rect 36597 43667 36643 43683
rect 37055 44941 37101 44957
rect 37055 44907 37061 44941
rect 37095 44907 37101 44941
rect 37055 44869 37101 44907
rect 37055 44835 37061 44869
rect 37095 44835 37101 44869
rect 37055 44797 37101 44835
rect 37055 44763 37061 44797
rect 37095 44763 37101 44797
rect 37055 44725 37101 44763
rect 37055 44691 37061 44725
rect 37095 44691 37101 44725
rect 37055 44653 37101 44691
rect 37055 44619 37061 44653
rect 37095 44619 37101 44653
rect 37055 44581 37101 44619
rect 37055 44547 37061 44581
rect 37095 44547 37101 44581
rect 37055 44509 37101 44547
rect 37055 44475 37061 44509
rect 37095 44475 37101 44509
rect 37055 44437 37101 44475
rect 37055 44403 37061 44437
rect 37095 44403 37101 44437
rect 37055 44365 37101 44403
rect 37055 44331 37061 44365
rect 37095 44331 37101 44365
rect 37055 44293 37101 44331
rect 37055 44259 37061 44293
rect 37095 44259 37101 44293
rect 37055 44221 37101 44259
rect 37055 44187 37061 44221
rect 37095 44187 37101 44221
rect 37055 44149 37101 44187
rect 37055 44115 37061 44149
rect 37095 44115 37101 44149
rect 37055 44077 37101 44115
rect 37055 44043 37061 44077
rect 37095 44043 37101 44077
rect 37055 44005 37101 44043
rect 37055 43971 37061 44005
rect 37095 43971 37101 44005
rect 37055 43933 37101 43971
rect 37055 43899 37061 43933
rect 37095 43899 37101 43933
rect 37055 43861 37101 43899
rect 37055 43827 37061 43861
rect 37095 43827 37101 43861
rect 37055 43789 37101 43827
rect 37055 43755 37061 43789
rect 37095 43755 37101 43789
rect 37055 43717 37101 43755
rect 37055 43683 37061 43717
rect 37095 43683 37101 43717
rect 37055 43667 37101 43683
rect 37513 44941 37559 44957
rect 37513 44907 37519 44941
rect 37553 44907 37559 44941
rect 37513 44869 37559 44907
rect 37513 44835 37519 44869
rect 37553 44835 37559 44869
rect 37513 44797 37559 44835
rect 37513 44763 37519 44797
rect 37553 44763 37559 44797
rect 37513 44725 37559 44763
rect 37513 44691 37519 44725
rect 37553 44691 37559 44725
rect 37513 44653 37559 44691
rect 37513 44619 37519 44653
rect 37553 44619 37559 44653
rect 37513 44581 37559 44619
rect 37513 44547 37519 44581
rect 37553 44547 37559 44581
rect 37513 44509 37559 44547
rect 37513 44475 37519 44509
rect 37553 44475 37559 44509
rect 37513 44437 37559 44475
rect 37513 44403 37519 44437
rect 37553 44403 37559 44437
rect 37513 44365 37559 44403
rect 37513 44331 37519 44365
rect 37553 44331 37559 44365
rect 37513 44293 37559 44331
rect 37513 44259 37519 44293
rect 37553 44259 37559 44293
rect 37513 44221 37559 44259
rect 37513 44187 37519 44221
rect 37553 44187 37559 44221
rect 37513 44149 37559 44187
rect 37513 44115 37519 44149
rect 37553 44115 37559 44149
rect 37513 44077 37559 44115
rect 37513 44043 37519 44077
rect 37553 44043 37559 44077
rect 37513 44005 37559 44043
rect 37513 43971 37519 44005
rect 37553 43971 37559 44005
rect 37513 43933 37559 43971
rect 37513 43899 37519 43933
rect 37553 43899 37559 43933
rect 37513 43861 37559 43899
rect 37513 43827 37519 43861
rect 37553 43827 37559 43861
rect 37513 43789 37559 43827
rect 37513 43755 37519 43789
rect 37553 43755 37559 43789
rect 37513 43717 37559 43755
rect 37513 43683 37519 43717
rect 37553 43683 37559 43717
rect 37513 43667 37559 43683
rect 37971 44941 38017 44957
rect 37971 44907 37977 44941
rect 38011 44907 38017 44941
rect 37971 44869 38017 44907
rect 37971 44835 37977 44869
rect 38011 44835 38017 44869
rect 37971 44797 38017 44835
rect 37971 44763 37977 44797
rect 38011 44763 38017 44797
rect 37971 44725 38017 44763
rect 37971 44691 37977 44725
rect 38011 44691 38017 44725
rect 37971 44653 38017 44691
rect 37971 44619 37977 44653
rect 38011 44619 38017 44653
rect 37971 44581 38017 44619
rect 37971 44547 37977 44581
rect 38011 44547 38017 44581
rect 37971 44509 38017 44547
rect 37971 44475 37977 44509
rect 38011 44475 38017 44509
rect 37971 44437 38017 44475
rect 37971 44403 37977 44437
rect 38011 44403 38017 44437
rect 37971 44365 38017 44403
rect 37971 44331 37977 44365
rect 38011 44331 38017 44365
rect 37971 44293 38017 44331
rect 37971 44259 37977 44293
rect 38011 44259 38017 44293
rect 37971 44221 38017 44259
rect 37971 44187 37977 44221
rect 38011 44187 38017 44221
rect 37971 44149 38017 44187
rect 37971 44115 37977 44149
rect 38011 44115 38017 44149
rect 37971 44077 38017 44115
rect 37971 44043 37977 44077
rect 38011 44043 38017 44077
rect 37971 44005 38017 44043
rect 37971 43971 37977 44005
rect 38011 43971 38017 44005
rect 37971 43933 38017 43971
rect 37971 43899 37977 43933
rect 38011 43899 38017 43933
rect 37971 43861 38017 43899
rect 37971 43827 37977 43861
rect 38011 43827 38017 43861
rect 37971 43789 38017 43827
rect 37971 43755 37977 43789
rect 38011 43755 38017 43789
rect 37971 43717 38017 43755
rect 37971 43683 37977 43717
rect 38011 43683 38017 43717
rect 37971 43667 38017 43683
rect 38429 44941 38475 44957
rect 38429 44907 38435 44941
rect 38469 44907 38475 44941
rect 38429 44869 38475 44907
rect 38429 44835 38435 44869
rect 38469 44835 38475 44869
rect 38429 44797 38475 44835
rect 38429 44763 38435 44797
rect 38469 44763 38475 44797
rect 38429 44725 38475 44763
rect 38429 44691 38435 44725
rect 38469 44691 38475 44725
rect 38429 44653 38475 44691
rect 38429 44619 38435 44653
rect 38469 44619 38475 44653
rect 38429 44581 38475 44619
rect 38429 44547 38435 44581
rect 38469 44547 38475 44581
rect 38429 44509 38475 44547
rect 38429 44475 38435 44509
rect 38469 44475 38475 44509
rect 38429 44437 38475 44475
rect 38429 44403 38435 44437
rect 38469 44403 38475 44437
rect 38429 44365 38475 44403
rect 38429 44331 38435 44365
rect 38469 44331 38475 44365
rect 38429 44293 38475 44331
rect 38429 44259 38435 44293
rect 38469 44259 38475 44293
rect 38429 44221 38475 44259
rect 38429 44187 38435 44221
rect 38469 44187 38475 44221
rect 38429 44149 38475 44187
rect 38429 44115 38435 44149
rect 38469 44115 38475 44149
rect 38429 44077 38475 44115
rect 38429 44043 38435 44077
rect 38469 44043 38475 44077
rect 38429 44005 38475 44043
rect 38429 43971 38435 44005
rect 38469 43971 38475 44005
rect 38429 43933 38475 43971
rect 38429 43899 38435 43933
rect 38469 43899 38475 43933
rect 38429 43861 38475 43899
rect 38429 43827 38435 43861
rect 38469 43827 38475 43861
rect 38429 43789 38475 43827
rect 38429 43755 38435 43789
rect 38469 43755 38475 43789
rect 38429 43717 38475 43755
rect 38429 43683 38435 43717
rect 38469 43683 38475 43717
rect 38429 43667 38475 43683
rect 38887 44941 38933 44957
rect 38887 44907 38893 44941
rect 38927 44907 38933 44941
rect 38887 44869 38933 44907
rect 38887 44835 38893 44869
rect 38927 44835 38933 44869
rect 38887 44797 38933 44835
rect 38887 44763 38893 44797
rect 38927 44763 38933 44797
rect 38887 44725 38933 44763
rect 38887 44691 38893 44725
rect 38927 44691 38933 44725
rect 38887 44653 38933 44691
rect 38887 44619 38893 44653
rect 38927 44619 38933 44653
rect 38887 44581 38933 44619
rect 38887 44547 38893 44581
rect 38927 44547 38933 44581
rect 38887 44509 38933 44547
rect 38887 44475 38893 44509
rect 38927 44475 38933 44509
rect 38887 44437 38933 44475
rect 38887 44403 38893 44437
rect 38927 44403 38933 44437
rect 38887 44365 38933 44403
rect 38887 44331 38893 44365
rect 38927 44331 38933 44365
rect 38887 44293 38933 44331
rect 38887 44259 38893 44293
rect 38927 44259 38933 44293
rect 38887 44221 38933 44259
rect 38887 44187 38893 44221
rect 38927 44187 38933 44221
rect 38887 44149 38933 44187
rect 38887 44115 38893 44149
rect 38927 44115 38933 44149
rect 38887 44077 38933 44115
rect 38887 44043 38893 44077
rect 38927 44043 38933 44077
rect 38887 44005 38933 44043
rect 38887 43971 38893 44005
rect 38927 43971 38933 44005
rect 38887 43933 38933 43971
rect 38887 43899 38893 43933
rect 38927 43899 38933 43933
rect 38887 43861 38933 43899
rect 38887 43827 38893 43861
rect 38927 43827 38933 43861
rect 38887 43789 38933 43827
rect 38887 43755 38893 43789
rect 38927 43755 38933 43789
rect 38887 43717 38933 43755
rect 38887 43683 38893 43717
rect 38927 43683 38933 43717
rect 38887 43667 38933 43683
rect 39345 44941 39391 44957
rect 39345 44907 39351 44941
rect 39385 44907 39391 44941
rect 39345 44869 39391 44907
rect 39345 44835 39351 44869
rect 39385 44835 39391 44869
rect 39345 44797 39391 44835
rect 39345 44763 39351 44797
rect 39385 44763 39391 44797
rect 39345 44725 39391 44763
rect 39345 44691 39351 44725
rect 39385 44691 39391 44725
rect 39345 44653 39391 44691
rect 39345 44619 39351 44653
rect 39385 44619 39391 44653
rect 39345 44581 39391 44619
rect 39345 44547 39351 44581
rect 39385 44547 39391 44581
rect 39345 44509 39391 44547
rect 39345 44475 39351 44509
rect 39385 44475 39391 44509
rect 39345 44437 39391 44475
rect 39345 44403 39351 44437
rect 39385 44403 39391 44437
rect 39345 44365 39391 44403
rect 39345 44331 39351 44365
rect 39385 44331 39391 44365
rect 39345 44293 39391 44331
rect 39345 44259 39351 44293
rect 39385 44259 39391 44293
rect 39345 44221 39391 44259
rect 39345 44187 39351 44221
rect 39385 44187 39391 44221
rect 39345 44149 39391 44187
rect 39345 44115 39351 44149
rect 39385 44115 39391 44149
rect 39345 44077 39391 44115
rect 39345 44043 39351 44077
rect 39385 44043 39391 44077
rect 39345 44005 39391 44043
rect 39345 43971 39351 44005
rect 39385 43971 39391 44005
rect 39345 43933 39391 43971
rect 39345 43899 39351 43933
rect 39385 43899 39391 43933
rect 39345 43861 39391 43899
rect 39345 43827 39351 43861
rect 39385 43827 39391 43861
rect 39345 43789 39391 43827
rect 39345 43755 39351 43789
rect 39385 43755 39391 43789
rect 39345 43717 39391 43755
rect 39345 43683 39351 43717
rect 39385 43683 39391 43717
rect 39345 43667 39391 43683
rect 39803 44941 39849 44957
rect 39803 44907 39809 44941
rect 39843 44907 39849 44941
rect 39803 44869 39849 44907
rect 39803 44835 39809 44869
rect 39843 44835 39849 44869
rect 39803 44797 39849 44835
rect 39803 44763 39809 44797
rect 39843 44763 39849 44797
rect 39803 44725 39849 44763
rect 39803 44691 39809 44725
rect 39843 44691 39849 44725
rect 39803 44653 39849 44691
rect 39803 44619 39809 44653
rect 39843 44619 39849 44653
rect 39803 44581 39849 44619
rect 39803 44547 39809 44581
rect 39843 44547 39849 44581
rect 39803 44509 39849 44547
rect 39803 44475 39809 44509
rect 39843 44475 39849 44509
rect 39803 44437 39849 44475
rect 39803 44403 39809 44437
rect 39843 44403 39849 44437
rect 39803 44365 39849 44403
rect 39803 44331 39809 44365
rect 39843 44331 39849 44365
rect 39803 44293 39849 44331
rect 39803 44259 39809 44293
rect 39843 44259 39849 44293
rect 39803 44221 39849 44259
rect 39803 44187 39809 44221
rect 39843 44187 39849 44221
rect 39803 44149 39849 44187
rect 39803 44115 39809 44149
rect 39843 44115 39849 44149
rect 39803 44077 39849 44115
rect 39803 44043 39809 44077
rect 39843 44043 39849 44077
rect 39803 44005 39849 44043
rect 39803 43971 39809 44005
rect 39843 43971 39849 44005
rect 39803 43933 39849 43971
rect 39803 43899 39809 43933
rect 39843 43899 39849 43933
rect 39803 43861 39849 43899
rect 39803 43827 39809 43861
rect 39843 43827 39849 43861
rect 39803 43789 39849 43827
rect 39803 43755 39809 43789
rect 39843 43755 39849 43789
rect 39803 43717 39849 43755
rect 39803 43683 39809 43717
rect 39843 43683 39849 43717
rect 39803 43667 39849 43683
rect 40261 44941 40307 44957
rect 40261 44907 40267 44941
rect 40301 44907 40307 44941
rect 40261 44869 40307 44907
rect 40261 44835 40267 44869
rect 40301 44835 40307 44869
rect 40261 44797 40307 44835
rect 40261 44763 40267 44797
rect 40301 44763 40307 44797
rect 40261 44725 40307 44763
rect 40261 44691 40267 44725
rect 40301 44691 40307 44725
rect 40261 44653 40307 44691
rect 40261 44619 40267 44653
rect 40301 44619 40307 44653
rect 40261 44581 40307 44619
rect 40261 44547 40267 44581
rect 40301 44547 40307 44581
rect 40261 44509 40307 44547
rect 40261 44475 40267 44509
rect 40301 44475 40307 44509
rect 40261 44437 40307 44475
rect 40261 44403 40267 44437
rect 40301 44403 40307 44437
rect 40261 44365 40307 44403
rect 40261 44331 40267 44365
rect 40301 44331 40307 44365
rect 40261 44293 40307 44331
rect 40261 44259 40267 44293
rect 40301 44259 40307 44293
rect 40261 44221 40307 44259
rect 40261 44187 40267 44221
rect 40301 44187 40307 44221
rect 40261 44149 40307 44187
rect 40261 44115 40267 44149
rect 40301 44115 40307 44149
rect 40261 44077 40307 44115
rect 40261 44043 40267 44077
rect 40301 44043 40307 44077
rect 40261 44005 40307 44043
rect 40261 43971 40267 44005
rect 40301 43971 40307 44005
rect 40261 43933 40307 43971
rect 40261 43899 40267 43933
rect 40301 43899 40307 43933
rect 40261 43861 40307 43899
rect 40261 43827 40267 43861
rect 40301 43827 40307 43861
rect 40261 43789 40307 43827
rect 40261 43755 40267 43789
rect 40301 43755 40307 43789
rect 40261 43717 40307 43755
rect 40261 43683 40267 43717
rect 40301 43683 40307 43717
rect 40261 43667 40307 43683
rect 40719 44941 40765 44957
rect 40719 44907 40725 44941
rect 40759 44907 40765 44941
rect 40719 44869 40765 44907
rect 40719 44835 40725 44869
rect 40759 44835 40765 44869
rect 40719 44797 40765 44835
rect 40719 44763 40725 44797
rect 40759 44763 40765 44797
rect 40719 44725 40765 44763
rect 40719 44691 40725 44725
rect 40759 44691 40765 44725
rect 40719 44653 40765 44691
rect 40719 44619 40725 44653
rect 40759 44619 40765 44653
rect 40719 44581 40765 44619
rect 40719 44547 40725 44581
rect 40759 44547 40765 44581
rect 40719 44509 40765 44547
rect 40719 44475 40725 44509
rect 40759 44475 40765 44509
rect 40719 44437 40765 44475
rect 40719 44403 40725 44437
rect 40759 44403 40765 44437
rect 40719 44365 40765 44403
rect 40719 44331 40725 44365
rect 40759 44331 40765 44365
rect 40719 44293 40765 44331
rect 40719 44259 40725 44293
rect 40759 44259 40765 44293
rect 40719 44221 40765 44259
rect 40719 44187 40725 44221
rect 40759 44187 40765 44221
rect 40719 44149 40765 44187
rect 40719 44115 40725 44149
rect 40759 44115 40765 44149
rect 40719 44077 40765 44115
rect 40719 44043 40725 44077
rect 40759 44043 40765 44077
rect 40719 44005 40765 44043
rect 40719 43971 40725 44005
rect 40759 43971 40765 44005
rect 40719 43933 40765 43971
rect 40719 43899 40725 43933
rect 40759 43899 40765 43933
rect 40719 43861 40765 43899
rect 40719 43827 40725 43861
rect 40759 43827 40765 43861
rect 40719 43789 40765 43827
rect 40719 43755 40725 43789
rect 40759 43755 40765 43789
rect 40719 43717 40765 43755
rect 40719 43683 40725 43717
rect 40759 43683 40765 43717
rect 40719 43667 40765 43683
rect 41177 44941 41223 44957
rect 41177 44907 41183 44941
rect 41217 44907 41223 44941
rect 41177 44869 41223 44907
rect 41177 44835 41183 44869
rect 41217 44835 41223 44869
rect 41177 44797 41223 44835
rect 41177 44763 41183 44797
rect 41217 44763 41223 44797
rect 41177 44725 41223 44763
rect 41177 44691 41183 44725
rect 41217 44691 41223 44725
rect 41177 44653 41223 44691
rect 41177 44619 41183 44653
rect 41217 44619 41223 44653
rect 41177 44581 41223 44619
rect 41177 44547 41183 44581
rect 41217 44547 41223 44581
rect 41177 44509 41223 44547
rect 41177 44475 41183 44509
rect 41217 44475 41223 44509
rect 41177 44437 41223 44475
rect 41177 44403 41183 44437
rect 41217 44403 41223 44437
rect 41177 44365 41223 44403
rect 41177 44331 41183 44365
rect 41217 44331 41223 44365
rect 41177 44293 41223 44331
rect 41177 44259 41183 44293
rect 41217 44259 41223 44293
rect 41177 44221 41223 44259
rect 41177 44187 41183 44221
rect 41217 44187 41223 44221
rect 41177 44149 41223 44187
rect 41177 44115 41183 44149
rect 41217 44115 41223 44149
rect 41177 44077 41223 44115
rect 41177 44043 41183 44077
rect 41217 44043 41223 44077
rect 41177 44005 41223 44043
rect 41177 43971 41183 44005
rect 41217 43971 41223 44005
rect 41177 43933 41223 43971
rect 41177 43899 41183 43933
rect 41217 43899 41223 43933
rect 41177 43861 41223 43899
rect 41177 43827 41183 43861
rect 41217 43827 41223 43861
rect 41177 43789 41223 43827
rect 41177 43755 41183 43789
rect 41217 43755 41223 43789
rect 41177 43717 41223 43755
rect 41177 43683 41183 43717
rect 41217 43683 41223 43717
rect 41177 43667 41223 43683
rect 41635 44941 41681 44957
rect 41635 44907 41641 44941
rect 41675 44907 41681 44941
rect 41635 44869 41681 44907
rect 41635 44835 41641 44869
rect 41675 44835 41681 44869
rect 41635 44797 41681 44835
rect 41635 44763 41641 44797
rect 41675 44763 41681 44797
rect 41635 44725 41681 44763
rect 41635 44691 41641 44725
rect 41675 44691 41681 44725
rect 41635 44653 41681 44691
rect 41635 44619 41641 44653
rect 41675 44619 41681 44653
rect 41635 44581 41681 44619
rect 41635 44547 41641 44581
rect 41675 44547 41681 44581
rect 41635 44509 41681 44547
rect 41635 44475 41641 44509
rect 41675 44475 41681 44509
rect 41635 44437 41681 44475
rect 41635 44403 41641 44437
rect 41675 44403 41681 44437
rect 41635 44365 41681 44403
rect 41635 44331 41641 44365
rect 41675 44331 41681 44365
rect 41635 44293 41681 44331
rect 41635 44259 41641 44293
rect 41675 44259 41681 44293
rect 41635 44221 41681 44259
rect 41635 44187 41641 44221
rect 41675 44187 41681 44221
rect 41635 44149 41681 44187
rect 41635 44115 41641 44149
rect 41675 44115 41681 44149
rect 41635 44077 41681 44115
rect 41635 44043 41641 44077
rect 41675 44043 41681 44077
rect 41635 44005 41681 44043
rect 41635 43971 41641 44005
rect 41675 43971 41681 44005
rect 41635 43933 41681 43971
rect 41635 43899 41641 43933
rect 41675 43899 41681 43933
rect 41635 43861 41681 43899
rect 41635 43827 41641 43861
rect 41675 43827 41681 43861
rect 41635 43789 41681 43827
rect 41635 43755 41641 43789
rect 41675 43755 41681 43789
rect 41635 43717 41681 43755
rect 41635 43683 41641 43717
rect 41675 43683 41681 43717
rect 41635 43667 41681 43683
rect 42093 44941 42139 44957
rect 42093 44907 42099 44941
rect 42133 44907 42139 44941
rect 42093 44869 42139 44907
rect 42093 44835 42099 44869
rect 42133 44835 42139 44869
rect 42093 44797 42139 44835
rect 42093 44763 42099 44797
rect 42133 44763 42139 44797
rect 42093 44725 42139 44763
rect 42093 44691 42099 44725
rect 42133 44691 42139 44725
rect 42093 44653 42139 44691
rect 42093 44619 42099 44653
rect 42133 44619 42139 44653
rect 42093 44581 42139 44619
rect 42093 44547 42099 44581
rect 42133 44547 42139 44581
rect 42093 44509 42139 44547
rect 42093 44475 42099 44509
rect 42133 44475 42139 44509
rect 42093 44437 42139 44475
rect 42093 44403 42099 44437
rect 42133 44403 42139 44437
rect 42093 44365 42139 44403
rect 42093 44331 42099 44365
rect 42133 44331 42139 44365
rect 42093 44293 42139 44331
rect 42093 44259 42099 44293
rect 42133 44259 42139 44293
rect 42093 44221 42139 44259
rect 42093 44187 42099 44221
rect 42133 44187 42139 44221
rect 42093 44149 42139 44187
rect 42093 44115 42099 44149
rect 42133 44115 42139 44149
rect 42093 44077 42139 44115
rect 42093 44043 42099 44077
rect 42133 44043 42139 44077
rect 42093 44005 42139 44043
rect 42093 43971 42099 44005
rect 42133 43971 42139 44005
rect 42093 43933 42139 43971
rect 42093 43899 42099 43933
rect 42133 43899 42139 43933
rect 42093 43861 42139 43899
rect 42093 43827 42099 43861
rect 42133 43827 42139 43861
rect 42093 43789 42139 43827
rect 42093 43755 42099 43789
rect 42133 43755 42139 43789
rect 42093 43717 42139 43755
rect 42093 43683 42099 43717
rect 42133 43683 42139 43717
rect 42093 43667 42139 43683
rect 42551 44941 42597 44957
rect 42551 44907 42557 44941
rect 42591 44907 42597 44941
rect 42551 44869 42597 44907
rect 42551 44835 42557 44869
rect 42591 44835 42597 44869
rect 42551 44797 42597 44835
rect 42986 44876 52314 44882
rect 42986 44842 43006 44876
rect 43040 44842 43096 44876
rect 43130 44842 43186 44876
rect 43220 44842 43276 44876
rect 43310 44842 43366 44876
rect 43400 44842 43456 44876
rect 43490 44842 43546 44876
rect 43580 44842 43636 44876
rect 43670 44842 43726 44876
rect 43760 44842 43816 44876
rect 43850 44842 43906 44876
rect 43940 44842 43996 44876
rect 44030 44842 44086 44876
rect 44120 44842 44176 44876
rect 44210 44842 44346 44876
rect 44380 44842 44436 44876
rect 44470 44842 44526 44876
rect 44560 44842 44616 44876
rect 44650 44842 44706 44876
rect 44740 44842 44796 44876
rect 44830 44842 44886 44876
rect 44920 44842 44976 44876
rect 45010 44842 45066 44876
rect 45100 44842 45156 44876
rect 45190 44842 45246 44876
rect 45280 44842 45336 44876
rect 45370 44842 45426 44876
rect 45460 44842 45516 44876
rect 45550 44842 45686 44876
rect 45720 44842 45776 44876
rect 45810 44842 45866 44876
rect 45900 44842 45956 44876
rect 45990 44842 46046 44876
rect 46080 44842 46136 44876
rect 46170 44842 46226 44876
rect 46260 44842 46316 44876
rect 46350 44842 46406 44876
rect 46440 44842 46496 44876
rect 46530 44842 46586 44876
rect 46620 44842 46676 44876
rect 46710 44842 46766 44876
rect 46800 44842 46856 44876
rect 46890 44842 47026 44876
rect 47060 44842 47116 44876
rect 47150 44842 47206 44876
rect 47240 44842 47296 44876
rect 47330 44842 47386 44876
rect 47420 44842 47476 44876
rect 47510 44842 47566 44876
rect 47600 44842 47656 44876
rect 47690 44842 47746 44876
rect 47780 44842 47836 44876
rect 47870 44842 47926 44876
rect 47960 44842 48016 44876
rect 48050 44842 48106 44876
rect 48140 44842 48196 44876
rect 48230 44842 48366 44876
rect 48400 44842 48456 44876
rect 48490 44842 48546 44876
rect 48580 44842 48636 44876
rect 48670 44842 48726 44876
rect 48760 44842 48816 44876
rect 48850 44842 48906 44876
rect 48940 44842 48996 44876
rect 49030 44842 49086 44876
rect 49120 44842 49176 44876
rect 49210 44842 49266 44876
rect 49300 44842 49356 44876
rect 49390 44842 49446 44876
rect 49480 44842 49536 44876
rect 49570 44842 49706 44876
rect 49740 44842 49796 44876
rect 49830 44842 49886 44876
rect 49920 44842 49976 44876
rect 50010 44842 50066 44876
rect 50100 44842 50156 44876
rect 50190 44842 50246 44876
rect 50280 44842 50336 44876
rect 50370 44842 50426 44876
rect 50460 44842 50516 44876
rect 50550 44842 50606 44876
rect 50640 44842 50696 44876
rect 50730 44842 50786 44876
rect 50820 44842 50876 44876
rect 50910 44842 51046 44876
rect 51080 44842 51136 44876
rect 51170 44842 51226 44876
rect 51260 44842 51316 44876
rect 51350 44842 51406 44876
rect 51440 44842 51496 44876
rect 51530 44842 51586 44876
rect 51620 44842 51676 44876
rect 51710 44842 51766 44876
rect 51800 44842 51856 44876
rect 51890 44842 51946 44876
rect 51980 44842 52036 44876
rect 52070 44842 52126 44876
rect 52160 44842 52216 44876
rect 52250 44842 52314 44876
rect 42986 44812 52314 44842
rect 42551 44763 42557 44797
rect 42591 44763 42597 44797
rect 42551 44725 42597 44763
rect 43272 44736 43300 44812
rect 43254 44732 43260 44736
rect 42551 44691 42557 44725
rect 42591 44691 42597 44725
rect 42551 44653 42597 44691
rect 43150 44716 43260 44732
rect 43312 44732 43318 44736
rect 43312 44716 52150 44732
rect 43150 44682 43170 44716
rect 43204 44682 43260 44716
rect 43312 44684 43350 44716
rect 43294 44682 43350 44684
rect 43384 44682 43440 44716
rect 43474 44682 43530 44716
rect 43564 44682 43620 44716
rect 43654 44682 43710 44716
rect 43744 44682 43800 44716
rect 43834 44682 43890 44716
rect 43924 44682 43980 44716
rect 44014 44682 44070 44716
rect 44104 44682 44510 44716
rect 44544 44682 44600 44716
rect 44634 44682 44690 44716
rect 44724 44682 44780 44716
rect 44814 44682 44870 44716
rect 44904 44682 44960 44716
rect 44994 44682 45050 44716
rect 45084 44682 45140 44716
rect 45174 44682 45230 44716
rect 45264 44682 45320 44716
rect 45354 44682 45410 44716
rect 45444 44682 45850 44716
rect 45884 44682 45940 44716
rect 45974 44682 46030 44716
rect 46064 44682 46120 44716
rect 46154 44682 46210 44716
rect 46244 44682 46300 44716
rect 46334 44682 46390 44716
rect 46424 44682 46480 44716
rect 46514 44682 46570 44716
rect 46604 44682 46660 44716
rect 46694 44682 46750 44716
rect 46784 44682 47190 44716
rect 47224 44682 47280 44716
rect 47314 44682 47370 44716
rect 47404 44682 47460 44716
rect 47494 44682 47550 44716
rect 47584 44682 47640 44716
rect 47674 44682 47730 44716
rect 47764 44682 47820 44716
rect 47854 44682 47910 44716
rect 47944 44682 48000 44716
rect 48034 44682 48090 44716
rect 48124 44682 48530 44716
rect 48564 44682 48620 44716
rect 48654 44682 48710 44716
rect 48744 44682 48800 44716
rect 48834 44682 48890 44716
rect 48924 44682 48980 44716
rect 49014 44682 49070 44716
rect 49104 44682 49160 44716
rect 49194 44682 49250 44716
rect 49284 44682 49340 44716
rect 49374 44682 49430 44716
rect 49464 44682 49870 44716
rect 49904 44682 49960 44716
rect 49994 44682 50050 44716
rect 50084 44682 50140 44716
rect 50174 44682 50230 44716
rect 50264 44682 50320 44716
rect 50354 44682 50410 44716
rect 50444 44682 50500 44716
rect 50534 44682 50590 44716
rect 50624 44682 50680 44716
rect 50714 44682 50770 44716
rect 50804 44682 51210 44716
rect 51244 44682 51300 44716
rect 51334 44682 51390 44716
rect 51424 44682 51480 44716
rect 51514 44682 51570 44716
rect 51604 44682 51660 44716
rect 51694 44682 51750 44716
rect 51784 44682 51840 44716
rect 51874 44682 51930 44716
rect 51964 44682 52020 44716
rect 52054 44682 52110 44716
rect 52144 44682 52150 44716
rect 43150 44662 52150 44682
rect 42551 44619 42557 44653
rect 42591 44619 42597 44653
rect 42551 44581 42597 44619
rect 42551 44547 42557 44581
rect 42591 44547 42597 44581
rect 42551 44509 42597 44547
rect 42551 44475 42557 44509
rect 42591 44475 42597 44509
rect 42551 44437 42597 44475
rect 42551 44403 42557 44437
rect 42591 44403 42597 44437
rect 42551 44365 42597 44403
rect 42551 44331 42557 44365
rect 42591 44331 42597 44365
rect 42551 44293 42597 44331
rect 42551 44259 42557 44293
rect 42591 44259 42597 44293
rect 42551 44221 42597 44259
rect 42551 44187 42557 44221
rect 42591 44187 42597 44221
rect 42551 44149 42597 44187
rect 42551 44115 42557 44149
rect 42591 44115 42597 44149
rect 42551 44077 42597 44115
rect 42551 44043 42557 44077
rect 42591 44043 42597 44077
rect 42551 44005 42597 44043
rect 42551 43971 42557 44005
rect 42591 43971 42597 44005
rect 42551 43933 42597 43971
rect 43324 44512 51976 44558
rect 43324 44478 43356 44512
rect 43390 44478 43456 44512
rect 43490 44478 43556 44512
rect 43590 44478 43656 44512
rect 43690 44478 43756 44512
rect 43790 44478 43856 44512
rect 43890 44478 44696 44512
rect 44730 44478 44796 44512
rect 44830 44478 44896 44512
rect 44930 44478 44996 44512
rect 45030 44478 45096 44512
rect 45130 44478 45196 44512
rect 45230 44478 46036 44512
rect 46070 44478 46136 44512
rect 46170 44478 46236 44512
rect 46270 44478 46336 44512
rect 46370 44478 46436 44512
rect 46470 44478 46536 44512
rect 46570 44478 47376 44512
rect 47410 44478 47476 44512
rect 47510 44478 47576 44512
rect 47610 44478 47676 44512
rect 47710 44478 47776 44512
rect 47810 44478 47876 44512
rect 47910 44478 48716 44512
rect 48750 44478 48816 44512
rect 48850 44478 48916 44512
rect 48950 44478 49016 44512
rect 49050 44478 49116 44512
rect 49150 44478 49216 44512
rect 49250 44478 50056 44512
rect 50090 44478 50156 44512
rect 50190 44478 50256 44512
rect 50290 44478 50356 44512
rect 50390 44478 50456 44512
rect 50490 44478 50556 44512
rect 50590 44478 51396 44512
rect 51430 44478 51496 44512
rect 51530 44478 51596 44512
rect 51630 44478 51696 44512
rect 51730 44478 51796 44512
rect 51830 44478 51896 44512
rect 51930 44478 51976 44512
rect 43324 44412 51976 44478
rect 43324 44378 43356 44412
rect 43390 44378 43456 44412
rect 43490 44378 43556 44412
rect 43590 44378 43656 44412
rect 43690 44378 43756 44412
rect 43790 44378 43856 44412
rect 43890 44378 44696 44412
rect 44730 44378 44796 44412
rect 44830 44378 44896 44412
rect 44930 44378 44996 44412
rect 45030 44378 45096 44412
rect 45130 44378 45196 44412
rect 45230 44378 46036 44412
rect 46070 44378 46136 44412
rect 46170 44378 46236 44412
rect 46270 44378 46336 44412
rect 46370 44378 46436 44412
rect 46470 44378 46536 44412
rect 46570 44378 47376 44412
rect 47410 44378 47476 44412
rect 47510 44378 47576 44412
rect 47610 44378 47676 44412
rect 47710 44378 47776 44412
rect 47810 44378 47876 44412
rect 47910 44378 48716 44412
rect 48750 44378 48816 44412
rect 48850 44378 48916 44412
rect 48950 44378 49016 44412
rect 49050 44378 49116 44412
rect 49150 44378 49216 44412
rect 49250 44378 50056 44412
rect 50090 44378 50156 44412
rect 50190 44378 50256 44412
rect 50290 44378 50356 44412
rect 50390 44378 50456 44412
rect 50490 44378 50556 44412
rect 50590 44378 51396 44412
rect 51430 44378 51496 44412
rect 51530 44378 51596 44412
rect 51630 44378 51696 44412
rect 51730 44378 51796 44412
rect 51830 44378 51896 44412
rect 51930 44378 51976 44412
rect 43324 44312 51976 44378
rect 43324 44278 43356 44312
rect 43390 44278 43456 44312
rect 43490 44278 43556 44312
rect 43590 44278 43656 44312
rect 43690 44278 43756 44312
rect 43790 44278 43856 44312
rect 43890 44278 44696 44312
rect 44730 44278 44796 44312
rect 44830 44278 44896 44312
rect 44930 44278 44996 44312
rect 45030 44278 45096 44312
rect 45130 44278 45196 44312
rect 45230 44278 46036 44312
rect 46070 44278 46136 44312
rect 46170 44278 46236 44312
rect 46270 44278 46336 44312
rect 46370 44278 46436 44312
rect 46470 44278 46536 44312
rect 46570 44278 47376 44312
rect 47410 44278 47476 44312
rect 47510 44278 47576 44312
rect 47610 44278 47676 44312
rect 47710 44278 47776 44312
rect 47810 44278 47876 44312
rect 47910 44278 48716 44312
rect 48750 44278 48816 44312
rect 48850 44278 48916 44312
rect 48950 44278 49016 44312
rect 49050 44278 49116 44312
rect 49150 44278 49216 44312
rect 49250 44278 50056 44312
rect 50090 44278 50156 44312
rect 50190 44278 50256 44312
rect 50290 44278 50356 44312
rect 50390 44278 50456 44312
rect 50490 44278 50556 44312
rect 50590 44278 51396 44312
rect 51430 44278 51496 44312
rect 51530 44278 51596 44312
rect 51630 44278 51696 44312
rect 51730 44278 51796 44312
rect 51830 44278 51896 44312
rect 51930 44278 51976 44312
rect 43324 44212 51976 44278
rect 43324 44178 43356 44212
rect 43390 44178 43456 44212
rect 43490 44178 43556 44212
rect 43590 44178 43656 44212
rect 43690 44178 43756 44212
rect 43790 44178 43856 44212
rect 43890 44178 44696 44212
rect 44730 44178 44796 44212
rect 44830 44178 44896 44212
rect 44930 44178 44996 44212
rect 45030 44178 45096 44212
rect 45130 44178 45196 44212
rect 45230 44178 46036 44212
rect 46070 44178 46136 44212
rect 46170 44178 46236 44212
rect 46270 44178 46336 44212
rect 46370 44178 46436 44212
rect 46470 44178 46536 44212
rect 46570 44178 47376 44212
rect 47410 44178 47476 44212
rect 47510 44178 47576 44212
rect 47610 44178 47676 44212
rect 47710 44178 47776 44212
rect 47810 44178 47876 44212
rect 47910 44178 48716 44212
rect 48750 44178 48816 44212
rect 48850 44178 48916 44212
rect 48950 44178 49016 44212
rect 49050 44178 49116 44212
rect 49150 44178 49216 44212
rect 49250 44178 50056 44212
rect 50090 44178 50156 44212
rect 50190 44178 50256 44212
rect 50290 44178 50356 44212
rect 50390 44178 50456 44212
rect 50490 44178 50556 44212
rect 50590 44178 51396 44212
rect 51430 44178 51496 44212
rect 51530 44178 51596 44212
rect 51630 44178 51696 44212
rect 51730 44178 51796 44212
rect 51830 44178 51896 44212
rect 51930 44178 51976 44212
rect 43324 44112 51976 44178
rect 43324 44078 43356 44112
rect 43390 44078 43456 44112
rect 43490 44078 43556 44112
rect 43590 44078 43656 44112
rect 43690 44078 43756 44112
rect 43790 44078 43856 44112
rect 43890 44078 44696 44112
rect 44730 44078 44796 44112
rect 44830 44078 44896 44112
rect 44930 44078 44996 44112
rect 45030 44078 45096 44112
rect 45130 44078 45196 44112
rect 45230 44078 46036 44112
rect 46070 44078 46136 44112
rect 46170 44078 46236 44112
rect 46270 44078 46336 44112
rect 46370 44078 46436 44112
rect 46470 44078 46536 44112
rect 46570 44078 47376 44112
rect 47410 44078 47476 44112
rect 47510 44078 47576 44112
rect 47610 44078 47676 44112
rect 47710 44078 47776 44112
rect 47810 44078 47876 44112
rect 47910 44078 48716 44112
rect 48750 44078 48816 44112
rect 48850 44078 48916 44112
rect 48950 44078 49016 44112
rect 49050 44078 49116 44112
rect 49150 44078 49216 44112
rect 49250 44078 50056 44112
rect 50090 44078 50156 44112
rect 50190 44078 50256 44112
rect 50290 44078 50356 44112
rect 50390 44078 50456 44112
rect 50490 44078 50556 44112
rect 50590 44078 51396 44112
rect 51430 44078 51496 44112
rect 51530 44078 51596 44112
rect 51630 44078 51696 44112
rect 51730 44078 51796 44112
rect 51830 44078 51896 44112
rect 51930 44078 51976 44112
rect 43324 44012 51976 44078
rect 43324 43978 43356 44012
rect 43390 43978 43456 44012
rect 43490 43978 43556 44012
rect 43590 43978 43656 44012
rect 43690 43978 43756 44012
rect 43790 43978 43856 44012
rect 43890 43978 44696 44012
rect 44730 43978 44796 44012
rect 44830 43978 44896 44012
rect 44930 43978 44996 44012
rect 45030 43978 45096 44012
rect 45130 43978 45196 44012
rect 45230 43978 46036 44012
rect 46070 43978 46136 44012
rect 46170 43978 46236 44012
rect 46270 43978 46336 44012
rect 46370 43978 46436 44012
rect 46470 43978 46536 44012
rect 46570 43978 47376 44012
rect 47410 43978 47476 44012
rect 47510 43978 47576 44012
rect 47610 43978 47676 44012
rect 47710 43978 47776 44012
rect 47810 43978 47876 44012
rect 47910 43978 48716 44012
rect 48750 43978 48816 44012
rect 48850 43978 48916 44012
rect 48950 43978 49016 44012
rect 49050 43978 49116 44012
rect 49150 43978 49216 44012
rect 49250 43978 50056 44012
rect 50090 43978 50156 44012
rect 50190 43978 50256 44012
rect 50290 43978 50356 44012
rect 50390 43978 50456 44012
rect 50490 43978 50556 44012
rect 50590 43978 51396 44012
rect 51430 43978 51496 44012
rect 51530 43978 51596 44012
rect 51630 43978 51696 44012
rect 51730 43978 51796 44012
rect 51830 43978 51896 44012
rect 51930 43978 51976 44012
rect 43324 43946 51976 43978
rect 42551 43899 42557 43933
rect 42591 43899 42597 43933
rect 42551 43861 42597 43899
rect 42551 43827 42557 43861
rect 42591 43827 42597 43861
rect 44100 43852 44128 43946
rect 42551 43789 42597 43827
rect 44082 43800 44088 43852
rect 44140 43800 44146 43852
rect 42551 43755 42557 43789
rect 42591 43755 42597 43789
rect 42551 43717 42597 43755
rect 42551 43683 42557 43717
rect 42591 43683 42597 43717
rect 42551 43667 42597 43683
rect 15010 43568 15016 43580
rect 14955 43540 15016 43568
rect 15010 43528 15016 43540
rect 15068 43528 15074 43580
rect 29454 43466 29460 43478
rect 29399 43438 29460 43466
rect 29454 43426 29460 43438
rect 29512 43426 29518 43478
rect 900 43370 57536 43372
rect 900 43254 922 43370
rect 2510 43329 55926 43370
rect 2510 43295 6101 43329
rect 6135 43295 6501 43329
rect 6535 43295 6901 43329
rect 6935 43295 7301 43329
rect 7335 43295 7701 43329
rect 7735 43295 8101 43329
rect 8135 43308 8501 43329
rect 8135 43295 8300 43308
rect 2510 43256 8300 43295
rect 8352 43295 8501 43308
rect 8535 43295 8901 43329
rect 8935 43295 9301 43329
rect 9335 43295 9701 43329
rect 9735 43295 10101 43329
rect 10135 43295 10501 43329
rect 10535 43295 10901 43329
rect 10935 43295 11301 43329
rect 11335 43295 11701 43329
rect 11735 43295 12101 43329
rect 12135 43295 12501 43329
rect 12535 43295 12901 43329
rect 12935 43295 14301 43329
rect 14335 43295 15213 43329
rect 15247 43295 15613 43329
rect 15647 43295 16013 43329
rect 16047 43295 16413 43329
rect 16447 43295 16813 43329
rect 16847 43295 17213 43329
rect 17247 43295 17613 43329
rect 17647 43295 18013 43329
rect 18047 43295 18413 43329
rect 18447 43295 18813 43329
rect 18847 43295 19213 43329
rect 19247 43295 19613 43329
rect 19647 43295 20013 43329
rect 20047 43295 20413 43329
rect 20447 43295 20813 43329
rect 20847 43295 21213 43329
rect 21247 43295 21613 43329
rect 21647 43295 22013 43329
rect 22047 43295 22413 43329
rect 22447 43295 22813 43329
rect 22847 43295 23213 43329
rect 23247 43295 23613 43329
rect 23647 43295 24013 43329
rect 24047 43295 24413 43329
rect 24447 43295 24813 43329
rect 24847 43295 25213 43329
rect 25247 43295 25613 43329
rect 25647 43295 26013 43329
rect 26047 43295 26413 43329
rect 26447 43295 26813 43329
rect 26847 43295 27213 43329
rect 27247 43295 27613 43329
rect 27647 43295 28013 43329
rect 28047 43295 28413 43329
rect 28447 43295 28813 43329
rect 28847 43295 29213 43329
rect 29247 43295 29613 43329
rect 29647 43295 30013 43329
rect 30047 43295 30413 43329
rect 30447 43295 30813 43329
rect 30847 43295 31213 43329
rect 31247 43295 31613 43329
rect 31647 43295 32013 43329
rect 32047 43295 32413 43329
rect 32447 43295 32813 43329
rect 32847 43295 33213 43329
rect 33247 43295 33613 43329
rect 33647 43295 34013 43329
rect 34047 43295 34413 43329
rect 34447 43295 34813 43329
rect 34847 43295 35213 43329
rect 35247 43295 35613 43329
rect 35647 43295 36013 43329
rect 36047 43295 36413 43329
rect 36447 43295 36813 43329
rect 36847 43295 37213 43329
rect 37247 43295 37613 43329
rect 37647 43295 38013 43329
rect 38047 43295 38413 43329
rect 38447 43295 38813 43329
rect 38847 43295 39213 43329
rect 39247 43295 39613 43329
rect 39647 43295 40013 43329
rect 40047 43295 40413 43329
rect 40447 43295 40813 43329
rect 40847 43295 41213 43329
rect 41247 43295 41613 43329
rect 41647 43295 42013 43329
rect 42047 43295 42413 43329
rect 42447 43295 43143 43329
rect 43177 43308 43343 43329
rect 43177 43295 43260 43308
rect 8352 43256 43260 43295
rect 43312 43295 43343 43308
rect 43377 43295 43543 43329
rect 43577 43295 43743 43329
rect 43777 43295 43943 43329
rect 43977 43295 44143 43329
rect 44177 43295 44343 43329
rect 44377 43295 44543 43329
rect 44577 43295 44743 43329
rect 44777 43295 44943 43329
rect 44977 43295 45143 43329
rect 45177 43295 45343 43329
rect 45377 43295 45543 43329
rect 45577 43295 45743 43329
rect 45777 43295 45943 43329
rect 45977 43295 46143 43329
rect 46177 43295 46343 43329
rect 46377 43295 46543 43329
rect 46577 43295 46743 43329
rect 46777 43295 46943 43329
rect 46977 43295 47143 43329
rect 47177 43295 47343 43329
rect 47377 43295 47543 43329
rect 47577 43295 47743 43329
rect 47777 43295 47943 43329
rect 47977 43295 48143 43329
rect 48177 43295 48343 43329
rect 48377 43295 48543 43329
rect 48577 43295 48743 43329
rect 48777 43295 48943 43329
rect 48977 43295 49143 43329
rect 49177 43295 49343 43329
rect 49377 43295 49543 43329
rect 49577 43295 49743 43329
rect 49777 43295 49943 43329
rect 49977 43295 50143 43329
rect 50177 43295 50343 43329
rect 50377 43295 50543 43329
rect 50577 43295 50743 43329
rect 50777 43295 50943 43329
rect 50977 43295 51143 43329
rect 51177 43295 51343 43329
rect 51377 43295 51543 43329
rect 51577 43295 51743 43329
rect 51777 43295 51943 43329
rect 51977 43295 52143 43329
rect 52177 43295 55926 43329
rect 43312 43256 55926 43295
rect 2510 43254 55926 43256
rect 57514 43254 57536 43370
rect 900 43252 57536 43254
rect 3348 41490 55088 41492
rect 3348 41374 3370 41490
rect 4958 41449 53478 41490
rect 4958 41415 6493 41449
rect 6527 41415 6893 41449
rect 6927 41415 7293 41449
rect 7327 41415 7693 41449
rect 7727 41415 8093 41449
rect 8127 41415 8493 41449
rect 8527 41415 8893 41449
rect 8927 41415 9293 41449
rect 9327 41415 9693 41449
rect 9727 41415 10093 41449
rect 10127 41415 10493 41449
rect 10527 41415 10893 41449
rect 10927 41415 11293 41449
rect 11327 41415 11693 41449
rect 11727 41415 12093 41449
rect 12127 41415 12493 41449
rect 12527 41415 12893 41449
rect 12927 41415 13293 41449
rect 13327 41415 15313 41449
rect 15347 41415 15713 41449
rect 15747 41415 16113 41449
rect 16147 41415 16513 41449
rect 16547 41415 16913 41449
rect 16947 41415 17313 41449
rect 17347 41415 17713 41449
rect 17747 41415 18113 41449
rect 18147 41415 18513 41449
rect 18547 41415 18913 41449
rect 18947 41415 19313 41449
rect 19347 41415 19713 41449
rect 19747 41415 20113 41449
rect 20147 41415 20513 41449
rect 20547 41415 20913 41449
rect 20947 41415 21313 41449
rect 21347 41415 21713 41449
rect 21747 41415 22113 41449
rect 22147 41415 22857 41449
rect 22891 41415 23257 41449
rect 23291 41415 23657 41449
rect 23691 41415 24057 41449
rect 24091 41415 24457 41449
rect 24491 41415 24857 41449
rect 24891 41415 25257 41449
rect 25291 41415 25657 41449
rect 25691 41415 26057 41449
rect 26091 41415 26457 41449
rect 26491 41415 26857 41449
rect 26891 41415 27257 41449
rect 27291 41415 27657 41449
rect 27691 41415 28057 41449
rect 28091 41415 29521 41449
rect 29555 41415 29921 41449
rect 29955 41415 30321 41449
rect 30355 41415 30721 41449
rect 30755 41415 31121 41449
rect 31155 41415 31521 41449
rect 31555 41415 31921 41449
rect 31955 41415 32321 41449
rect 32355 41415 32721 41449
rect 32755 41415 33121 41449
rect 33155 41415 33521 41449
rect 33555 41415 33921 41449
rect 33955 41415 34321 41449
rect 34355 41415 34721 41449
rect 34755 41415 37459 41449
rect 37493 41415 37859 41449
rect 37893 41415 38259 41449
rect 38293 41415 38659 41449
rect 38693 41415 39059 41449
rect 39093 41415 39459 41449
rect 39493 41415 39859 41449
rect 39893 41415 40259 41449
rect 40293 41415 40659 41449
rect 40693 41415 41059 41449
rect 41093 41415 41967 41449
rect 42001 41415 42167 41449
rect 42201 41415 42367 41449
rect 42401 41415 42567 41449
rect 42601 41415 42767 41449
rect 42801 41415 42967 41449
rect 43001 41415 43167 41449
rect 43201 41415 43367 41449
rect 43401 41415 43567 41449
rect 43601 41415 43767 41449
rect 43801 41415 43967 41449
rect 44001 41415 44167 41449
rect 44201 41415 44367 41449
rect 44401 41415 44567 41449
rect 44601 41415 44767 41449
rect 44801 41415 44967 41449
rect 45001 41415 45167 41449
rect 45201 41415 45367 41449
rect 45401 41415 45567 41449
rect 45601 41415 45767 41449
rect 45801 41415 45967 41449
rect 46001 41415 46167 41449
rect 46201 41415 46367 41449
rect 46401 41415 46567 41449
rect 46601 41415 46767 41449
rect 46801 41415 46967 41449
rect 47001 41415 47167 41449
rect 47201 41415 47367 41449
rect 47401 41415 47567 41449
rect 47601 41415 47767 41449
rect 47801 41415 47967 41449
rect 48001 41415 48167 41449
rect 48201 41415 48367 41449
rect 48401 41415 48567 41449
rect 48601 41415 48767 41449
rect 48801 41415 48967 41449
rect 49001 41415 49167 41449
rect 49201 41415 49367 41449
rect 49401 41415 49567 41449
rect 49601 41415 49767 41449
rect 49801 41415 49967 41449
rect 50001 41415 50167 41449
rect 50201 41415 50367 41449
rect 50401 41415 50567 41449
rect 50601 41415 50767 41449
rect 50801 41415 50967 41449
rect 51001 41415 51167 41449
rect 51201 41415 51367 41449
rect 51401 41415 51567 41449
rect 51601 41415 51767 41449
rect 51801 41415 51967 41449
rect 52001 41415 52167 41449
rect 52201 41415 52367 41449
rect 52401 41415 53478 41449
rect 4958 41374 53478 41415
rect 55066 41374 55088 41490
rect 3348 41372 55088 41374
rect 24872 41265 24900 41372
rect 24857 41259 24915 41265
rect 24857 41225 24869 41259
rect 24903 41225 24915 41259
rect 24857 41219 24915 41225
rect 32600 41197 32628 41372
rect 22715 41181 22761 41197
rect 22715 41147 22721 41181
rect 22755 41147 22761 41181
rect 22715 41109 22761 41147
rect 22715 41075 22721 41109
rect 22755 41075 22761 41109
rect 22715 41037 22761 41075
rect 22715 41003 22721 41037
rect 22755 41003 22761 41037
rect 22715 40965 22761 41003
rect 22715 40931 22721 40965
rect 22755 40931 22761 40965
rect 22715 40893 22761 40931
rect 22715 40859 22721 40893
rect 22755 40859 22761 40893
rect 22715 40821 22761 40859
rect 22715 40787 22721 40821
rect 22755 40787 22761 40821
rect 22715 40749 22761 40787
rect 22715 40715 22721 40749
rect 22755 40715 22761 40749
rect 22715 40677 22761 40715
rect 22715 40643 22721 40677
rect 22755 40643 22761 40677
rect 22715 40605 22761 40643
rect 22715 40571 22721 40605
rect 22755 40571 22761 40605
rect 22715 40533 22761 40571
rect 22715 40499 22721 40533
rect 22755 40499 22761 40533
rect 22715 40461 22761 40499
rect 22715 40427 22721 40461
rect 22755 40427 22761 40461
rect 22715 40389 22761 40427
rect 22715 40355 22721 40389
rect 22755 40355 22761 40389
rect 22715 40317 22761 40355
rect 22715 40283 22721 40317
rect 22755 40283 22761 40317
rect 22715 40245 22761 40283
rect 22715 40211 22721 40245
rect 22755 40211 22761 40245
rect 22715 40173 22761 40211
rect 22715 40139 22721 40173
rect 22755 40139 22761 40173
rect 22715 40101 22761 40139
rect 22715 40067 22721 40101
rect 22755 40067 22761 40101
rect 22715 40029 22761 40067
rect 22715 39995 22721 40029
rect 22755 39995 22761 40029
rect 22715 39957 22761 39995
rect 22715 39923 22721 39957
rect 22755 39923 22761 39957
rect 22715 39907 22761 39923
rect 23173 41181 23219 41197
rect 23173 41147 23179 41181
rect 23213 41147 23219 41181
rect 23173 41109 23219 41147
rect 23173 41075 23179 41109
rect 23213 41075 23219 41109
rect 23173 41037 23219 41075
rect 23173 41003 23179 41037
rect 23213 41003 23219 41037
rect 23173 40965 23219 41003
rect 23173 40931 23179 40965
rect 23213 40931 23219 40965
rect 23173 40893 23219 40931
rect 23173 40859 23179 40893
rect 23213 40859 23219 40893
rect 23173 40821 23219 40859
rect 23173 40787 23179 40821
rect 23213 40787 23219 40821
rect 23173 40749 23219 40787
rect 23173 40715 23179 40749
rect 23213 40715 23219 40749
rect 23173 40677 23219 40715
rect 23173 40643 23179 40677
rect 23213 40643 23219 40677
rect 23173 40605 23219 40643
rect 23173 40571 23179 40605
rect 23213 40571 23219 40605
rect 23173 40533 23219 40571
rect 23173 40499 23179 40533
rect 23213 40499 23219 40533
rect 23173 40461 23219 40499
rect 23173 40427 23179 40461
rect 23213 40427 23219 40461
rect 23173 40389 23219 40427
rect 23173 40355 23179 40389
rect 23213 40355 23219 40389
rect 23173 40317 23219 40355
rect 23173 40283 23179 40317
rect 23213 40283 23219 40317
rect 23173 40245 23219 40283
rect 23173 40211 23179 40245
rect 23213 40211 23219 40245
rect 23173 40173 23219 40211
rect 23173 40139 23179 40173
rect 23213 40139 23219 40173
rect 23173 40101 23219 40139
rect 23173 40067 23179 40101
rect 23213 40067 23219 40101
rect 23173 40029 23219 40067
rect 23173 39995 23179 40029
rect 23213 39995 23219 40029
rect 23173 39957 23219 39995
rect 23173 39923 23179 39957
rect 23213 39923 23219 39957
rect 23173 39907 23219 39923
rect 23631 41181 23677 41197
rect 23631 41147 23637 41181
rect 23671 41147 23677 41181
rect 23631 41109 23677 41147
rect 23631 41075 23637 41109
rect 23671 41075 23677 41109
rect 23631 41037 23677 41075
rect 23631 41003 23637 41037
rect 23671 41003 23677 41037
rect 23631 40965 23677 41003
rect 23631 40931 23637 40965
rect 23671 40931 23677 40965
rect 23631 40893 23677 40931
rect 23631 40859 23637 40893
rect 23671 40859 23677 40893
rect 23631 40821 23677 40859
rect 23631 40787 23637 40821
rect 23671 40787 23677 40821
rect 23631 40749 23677 40787
rect 23631 40715 23637 40749
rect 23671 40715 23677 40749
rect 23631 40677 23677 40715
rect 23631 40643 23637 40677
rect 23671 40643 23677 40677
rect 23631 40605 23677 40643
rect 23631 40571 23637 40605
rect 23671 40571 23677 40605
rect 23631 40533 23677 40571
rect 23631 40499 23637 40533
rect 23671 40499 23677 40533
rect 23631 40461 23677 40499
rect 23631 40427 23637 40461
rect 23671 40427 23677 40461
rect 23631 40389 23677 40427
rect 23631 40355 23637 40389
rect 23671 40355 23677 40389
rect 23631 40317 23677 40355
rect 23631 40283 23637 40317
rect 23671 40283 23677 40317
rect 23631 40245 23677 40283
rect 23631 40211 23637 40245
rect 23671 40211 23677 40245
rect 23631 40173 23677 40211
rect 23631 40139 23637 40173
rect 23671 40139 23677 40173
rect 23631 40101 23677 40139
rect 23631 40067 23637 40101
rect 23671 40067 23677 40101
rect 23631 40029 23677 40067
rect 23631 39995 23637 40029
rect 23671 39995 23677 40029
rect 23631 39957 23677 39995
rect 23631 39923 23637 39957
rect 23671 39923 23677 39957
rect 23631 39907 23677 39923
rect 24089 41181 24135 41197
rect 24089 41147 24095 41181
rect 24129 41147 24135 41181
rect 24089 41109 24135 41147
rect 24089 41075 24095 41109
rect 24129 41075 24135 41109
rect 24089 41037 24135 41075
rect 24089 41003 24095 41037
rect 24129 41003 24135 41037
rect 24089 40965 24135 41003
rect 24089 40931 24095 40965
rect 24129 40931 24135 40965
rect 24089 40893 24135 40931
rect 24089 40859 24095 40893
rect 24129 40859 24135 40893
rect 24089 40821 24135 40859
rect 24089 40787 24095 40821
rect 24129 40787 24135 40821
rect 24089 40749 24135 40787
rect 24089 40715 24095 40749
rect 24129 40715 24135 40749
rect 24089 40677 24135 40715
rect 24089 40643 24095 40677
rect 24129 40643 24135 40677
rect 24089 40605 24135 40643
rect 24089 40571 24095 40605
rect 24129 40571 24135 40605
rect 24089 40533 24135 40571
rect 24089 40499 24095 40533
rect 24129 40499 24135 40533
rect 24089 40461 24135 40499
rect 24089 40427 24095 40461
rect 24129 40427 24135 40461
rect 24089 40389 24135 40427
rect 24089 40355 24095 40389
rect 24129 40355 24135 40389
rect 24089 40317 24135 40355
rect 24089 40283 24095 40317
rect 24129 40283 24135 40317
rect 24089 40245 24135 40283
rect 24089 40211 24095 40245
rect 24129 40211 24135 40245
rect 24089 40173 24135 40211
rect 24089 40139 24095 40173
rect 24129 40139 24135 40173
rect 24089 40101 24135 40139
rect 24089 40067 24095 40101
rect 24129 40067 24135 40101
rect 24089 40029 24135 40067
rect 24089 39995 24095 40029
rect 24129 39995 24135 40029
rect 24089 39957 24135 39995
rect 24089 39923 24095 39957
rect 24129 39923 24135 39957
rect 24089 39907 24135 39923
rect 24547 41181 24593 41197
rect 24547 41147 24553 41181
rect 24587 41147 24593 41181
rect 24547 41109 24593 41147
rect 24547 41075 24553 41109
rect 24587 41075 24593 41109
rect 24547 41037 24593 41075
rect 24547 41003 24553 41037
rect 24587 41003 24593 41037
rect 24547 40965 24593 41003
rect 24547 40931 24553 40965
rect 24587 40931 24593 40965
rect 24547 40893 24593 40931
rect 24547 40859 24553 40893
rect 24587 40859 24593 40893
rect 24547 40821 24593 40859
rect 24547 40787 24553 40821
rect 24587 40787 24593 40821
rect 24547 40749 24593 40787
rect 24547 40715 24553 40749
rect 24587 40715 24593 40749
rect 24547 40677 24593 40715
rect 24547 40643 24553 40677
rect 24587 40643 24593 40677
rect 24547 40605 24593 40643
rect 24547 40571 24553 40605
rect 24587 40571 24593 40605
rect 24547 40533 24593 40571
rect 24547 40499 24553 40533
rect 24587 40499 24593 40533
rect 24547 40461 24593 40499
rect 24547 40427 24553 40461
rect 24587 40427 24593 40461
rect 24547 40389 24593 40427
rect 24547 40355 24553 40389
rect 24587 40355 24593 40389
rect 24547 40317 24593 40355
rect 24547 40283 24553 40317
rect 24587 40283 24593 40317
rect 24547 40245 24593 40283
rect 24547 40211 24553 40245
rect 24587 40211 24593 40245
rect 24547 40173 24593 40211
rect 24547 40139 24553 40173
rect 24587 40139 24593 40173
rect 24547 40101 24593 40139
rect 24547 40067 24553 40101
rect 24587 40067 24593 40101
rect 24547 40029 24593 40067
rect 24547 39995 24553 40029
rect 24587 39995 24593 40029
rect 24547 39957 24593 39995
rect 24547 39923 24553 39957
rect 24587 39923 24593 39957
rect 24547 39907 24593 39923
rect 25005 41181 25051 41197
rect 25005 41147 25011 41181
rect 25045 41147 25051 41181
rect 25005 41109 25051 41147
rect 25005 41075 25011 41109
rect 25045 41075 25051 41109
rect 25005 41037 25051 41075
rect 25005 41003 25011 41037
rect 25045 41003 25051 41037
rect 25005 40965 25051 41003
rect 25005 40931 25011 40965
rect 25045 40931 25051 40965
rect 25005 40893 25051 40931
rect 25005 40859 25011 40893
rect 25045 40859 25051 40893
rect 25005 40821 25051 40859
rect 25005 40787 25011 40821
rect 25045 40787 25051 40821
rect 25005 40749 25051 40787
rect 25005 40715 25011 40749
rect 25045 40715 25051 40749
rect 25005 40677 25051 40715
rect 25005 40643 25011 40677
rect 25045 40643 25051 40677
rect 25005 40605 25051 40643
rect 25005 40571 25011 40605
rect 25045 40571 25051 40605
rect 25005 40533 25051 40571
rect 25005 40499 25011 40533
rect 25045 40499 25051 40533
rect 25005 40461 25051 40499
rect 25005 40427 25011 40461
rect 25045 40427 25051 40461
rect 25005 40389 25051 40427
rect 25005 40355 25011 40389
rect 25045 40355 25051 40389
rect 25005 40317 25051 40355
rect 25005 40283 25011 40317
rect 25045 40283 25051 40317
rect 25005 40245 25051 40283
rect 25005 40211 25011 40245
rect 25045 40211 25051 40245
rect 25005 40173 25051 40211
rect 25005 40139 25011 40173
rect 25045 40139 25051 40173
rect 25005 40101 25051 40139
rect 25005 40067 25011 40101
rect 25045 40067 25051 40101
rect 25005 40029 25051 40067
rect 25005 39995 25011 40029
rect 25045 39995 25051 40029
rect 25005 39957 25051 39995
rect 25005 39923 25011 39957
rect 25045 39923 25051 39957
rect 25005 39907 25051 39923
rect 25463 41181 25509 41197
rect 25463 41147 25469 41181
rect 25503 41147 25509 41181
rect 25463 41109 25509 41147
rect 25463 41075 25469 41109
rect 25503 41075 25509 41109
rect 25463 41037 25509 41075
rect 25463 41003 25469 41037
rect 25503 41003 25509 41037
rect 25463 40965 25509 41003
rect 25463 40931 25469 40965
rect 25503 40931 25509 40965
rect 25463 40893 25509 40931
rect 25463 40859 25469 40893
rect 25503 40859 25509 40893
rect 25463 40821 25509 40859
rect 25463 40787 25469 40821
rect 25503 40787 25509 40821
rect 25463 40749 25509 40787
rect 25463 40715 25469 40749
rect 25503 40715 25509 40749
rect 25463 40677 25509 40715
rect 25463 40643 25469 40677
rect 25503 40643 25509 40677
rect 25463 40605 25509 40643
rect 25463 40571 25469 40605
rect 25503 40571 25509 40605
rect 25463 40533 25509 40571
rect 25463 40499 25469 40533
rect 25503 40499 25509 40533
rect 25463 40461 25509 40499
rect 25463 40427 25469 40461
rect 25503 40427 25509 40461
rect 25463 40389 25509 40427
rect 25463 40355 25469 40389
rect 25503 40355 25509 40389
rect 25463 40317 25509 40355
rect 25463 40283 25469 40317
rect 25503 40283 25509 40317
rect 25463 40245 25509 40283
rect 25463 40211 25469 40245
rect 25503 40211 25509 40245
rect 25463 40173 25509 40211
rect 25463 40139 25469 40173
rect 25503 40139 25509 40173
rect 25463 40101 25509 40139
rect 25463 40067 25469 40101
rect 25503 40067 25509 40101
rect 25463 40029 25509 40067
rect 25463 39995 25469 40029
rect 25503 39995 25509 40029
rect 25463 39957 25509 39995
rect 25463 39923 25469 39957
rect 25503 39923 25509 39957
rect 25463 39907 25509 39923
rect 25921 41181 25967 41197
rect 25921 41147 25927 41181
rect 25961 41147 25967 41181
rect 25921 41109 25967 41147
rect 25921 41075 25927 41109
rect 25961 41075 25967 41109
rect 25921 41037 25967 41075
rect 25921 41003 25927 41037
rect 25961 41003 25967 41037
rect 25921 40965 25967 41003
rect 25921 40931 25927 40965
rect 25961 40931 25967 40965
rect 25921 40893 25967 40931
rect 25921 40859 25927 40893
rect 25961 40859 25967 40893
rect 25921 40821 25967 40859
rect 25921 40787 25927 40821
rect 25961 40787 25967 40821
rect 25921 40749 25967 40787
rect 25921 40715 25927 40749
rect 25961 40715 25967 40749
rect 25921 40677 25967 40715
rect 25921 40643 25927 40677
rect 25961 40643 25967 40677
rect 25921 40605 25967 40643
rect 25921 40571 25927 40605
rect 25961 40571 25967 40605
rect 25921 40533 25967 40571
rect 25921 40499 25927 40533
rect 25961 40499 25967 40533
rect 25921 40461 25967 40499
rect 25921 40427 25927 40461
rect 25961 40427 25967 40461
rect 25921 40389 25967 40427
rect 25921 40355 25927 40389
rect 25961 40355 25967 40389
rect 25921 40317 25967 40355
rect 25921 40283 25927 40317
rect 25961 40283 25967 40317
rect 25921 40245 25967 40283
rect 25921 40211 25927 40245
rect 25961 40211 25967 40245
rect 25921 40173 25967 40211
rect 25921 40139 25927 40173
rect 25961 40139 25967 40173
rect 25921 40101 25967 40139
rect 25921 40067 25927 40101
rect 25961 40067 25967 40101
rect 25921 40029 25967 40067
rect 25921 39995 25927 40029
rect 25961 39995 25967 40029
rect 25921 39957 25967 39995
rect 25921 39923 25927 39957
rect 25961 39923 25967 39957
rect 25921 39907 25967 39923
rect 26379 41181 26425 41197
rect 26379 41147 26385 41181
rect 26419 41147 26425 41181
rect 26379 41109 26425 41147
rect 26379 41075 26385 41109
rect 26419 41075 26425 41109
rect 26379 41037 26425 41075
rect 26379 41003 26385 41037
rect 26419 41003 26425 41037
rect 26379 40965 26425 41003
rect 26379 40931 26385 40965
rect 26419 40931 26425 40965
rect 26379 40893 26425 40931
rect 26379 40859 26385 40893
rect 26419 40859 26425 40893
rect 26379 40821 26425 40859
rect 26379 40787 26385 40821
rect 26419 40787 26425 40821
rect 26379 40749 26425 40787
rect 26379 40715 26385 40749
rect 26419 40715 26425 40749
rect 26379 40677 26425 40715
rect 26379 40643 26385 40677
rect 26419 40643 26425 40677
rect 26379 40605 26425 40643
rect 26379 40571 26385 40605
rect 26419 40571 26425 40605
rect 26379 40533 26425 40571
rect 26379 40499 26385 40533
rect 26419 40499 26425 40533
rect 26379 40461 26425 40499
rect 26379 40427 26385 40461
rect 26419 40427 26425 40461
rect 26379 40389 26425 40427
rect 26379 40355 26385 40389
rect 26419 40355 26425 40389
rect 26379 40317 26425 40355
rect 26379 40283 26385 40317
rect 26419 40283 26425 40317
rect 26379 40245 26425 40283
rect 26379 40211 26385 40245
rect 26419 40211 26425 40245
rect 26379 40173 26425 40211
rect 26379 40139 26385 40173
rect 26419 40139 26425 40173
rect 26379 40101 26425 40139
rect 26379 40067 26385 40101
rect 26419 40067 26425 40101
rect 26379 40029 26425 40067
rect 26379 39995 26385 40029
rect 26419 39995 26425 40029
rect 26379 39957 26425 39995
rect 26379 39923 26385 39957
rect 26419 39923 26425 39957
rect 26379 39907 26425 39923
rect 26837 41181 26883 41197
rect 26837 41147 26843 41181
rect 26877 41147 26883 41181
rect 26837 41109 26883 41147
rect 26837 41075 26843 41109
rect 26877 41075 26883 41109
rect 26837 41037 26883 41075
rect 26837 41003 26843 41037
rect 26877 41003 26883 41037
rect 26837 40965 26883 41003
rect 26837 40931 26843 40965
rect 26877 40931 26883 40965
rect 26837 40893 26883 40931
rect 26837 40859 26843 40893
rect 26877 40859 26883 40893
rect 26837 40821 26883 40859
rect 26837 40787 26843 40821
rect 26877 40787 26883 40821
rect 26837 40749 26883 40787
rect 26837 40715 26843 40749
rect 26877 40715 26883 40749
rect 26837 40677 26883 40715
rect 26837 40643 26843 40677
rect 26877 40643 26883 40677
rect 26837 40605 26883 40643
rect 26837 40571 26843 40605
rect 26877 40571 26883 40605
rect 26837 40533 26883 40571
rect 26837 40499 26843 40533
rect 26877 40499 26883 40533
rect 26837 40461 26883 40499
rect 26837 40427 26843 40461
rect 26877 40427 26883 40461
rect 26837 40389 26883 40427
rect 26837 40355 26843 40389
rect 26877 40355 26883 40389
rect 26837 40317 26883 40355
rect 26837 40283 26843 40317
rect 26877 40283 26883 40317
rect 26837 40245 26883 40283
rect 26837 40211 26843 40245
rect 26877 40211 26883 40245
rect 26837 40173 26883 40211
rect 26837 40139 26843 40173
rect 26877 40139 26883 40173
rect 26837 40101 26883 40139
rect 26837 40067 26843 40101
rect 26877 40067 26883 40101
rect 26837 40029 26883 40067
rect 26837 39995 26843 40029
rect 26877 39995 26883 40029
rect 26837 39957 26883 39995
rect 26837 39923 26843 39957
rect 26877 39923 26883 39957
rect 26837 39907 26883 39923
rect 27295 41181 27341 41197
rect 27295 41147 27301 41181
rect 27335 41147 27341 41181
rect 27295 41109 27341 41147
rect 27295 41075 27301 41109
rect 27335 41075 27341 41109
rect 27295 41037 27341 41075
rect 27295 41003 27301 41037
rect 27335 41003 27341 41037
rect 27295 40965 27341 41003
rect 27295 40931 27301 40965
rect 27335 40931 27341 40965
rect 27295 40893 27341 40931
rect 27295 40859 27301 40893
rect 27335 40859 27341 40893
rect 27295 40821 27341 40859
rect 27295 40787 27301 40821
rect 27335 40787 27341 40821
rect 27295 40749 27341 40787
rect 27295 40715 27301 40749
rect 27335 40715 27341 40749
rect 27295 40677 27341 40715
rect 27295 40643 27301 40677
rect 27335 40643 27341 40677
rect 27295 40605 27341 40643
rect 27295 40571 27301 40605
rect 27335 40571 27341 40605
rect 27295 40533 27341 40571
rect 27295 40499 27301 40533
rect 27335 40499 27341 40533
rect 27295 40461 27341 40499
rect 27295 40427 27301 40461
rect 27335 40427 27341 40461
rect 27295 40389 27341 40427
rect 27295 40355 27301 40389
rect 27335 40355 27341 40389
rect 27295 40317 27341 40355
rect 27295 40283 27301 40317
rect 27335 40283 27341 40317
rect 27295 40245 27341 40283
rect 27295 40211 27301 40245
rect 27335 40211 27341 40245
rect 27295 40173 27341 40211
rect 27295 40139 27301 40173
rect 27335 40139 27341 40173
rect 27295 40101 27341 40139
rect 27295 40067 27301 40101
rect 27335 40067 27341 40101
rect 27295 40029 27341 40067
rect 27295 39995 27301 40029
rect 27335 39995 27341 40029
rect 27295 39957 27341 39995
rect 27295 39923 27301 39957
rect 27335 39923 27341 39957
rect 27295 39907 27341 39923
rect 27753 41181 27799 41197
rect 27753 41147 27759 41181
rect 27793 41147 27799 41181
rect 27753 41109 27799 41147
rect 27753 41075 27759 41109
rect 27793 41075 27799 41109
rect 27753 41037 27799 41075
rect 27753 41003 27759 41037
rect 27793 41003 27799 41037
rect 27753 40965 27799 41003
rect 27753 40931 27759 40965
rect 27793 40931 27799 40965
rect 27753 40893 27799 40931
rect 27753 40859 27759 40893
rect 27793 40859 27799 40893
rect 27753 40821 27799 40859
rect 27753 40787 27759 40821
rect 27793 40787 27799 40821
rect 27753 40749 27799 40787
rect 27753 40715 27759 40749
rect 27793 40715 27799 40749
rect 27753 40677 27799 40715
rect 27753 40643 27759 40677
rect 27793 40643 27799 40677
rect 27753 40605 27799 40643
rect 27753 40571 27759 40605
rect 27793 40571 27799 40605
rect 27753 40533 27799 40571
rect 27753 40499 27759 40533
rect 27793 40499 27799 40533
rect 27753 40461 27799 40499
rect 27753 40427 27759 40461
rect 27793 40427 27799 40461
rect 27753 40389 27799 40427
rect 27753 40355 27759 40389
rect 27793 40355 27799 40389
rect 27753 40317 27799 40355
rect 27753 40283 27759 40317
rect 27793 40283 27799 40317
rect 27753 40245 27799 40283
rect 27753 40211 27759 40245
rect 27793 40211 27799 40245
rect 27753 40173 27799 40211
rect 27753 40139 27759 40173
rect 27793 40139 27799 40173
rect 27753 40101 27799 40139
rect 27753 40067 27759 40101
rect 27793 40067 27799 40101
rect 27753 40029 27799 40067
rect 27753 39995 27759 40029
rect 27793 39995 27799 40029
rect 27753 39957 27799 39995
rect 27753 39923 27759 39957
rect 27793 39923 27799 39957
rect 27753 39907 27799 39923
rect 28211 41181 28257 41197
rect 28211 41147 28217 41181
rect 28251 41147 28257 41181
rect 28211 41109 28257 41147
rect 28211 41075 28217 41109
rect 28251 41075 28257 41109
rect 28211 41037 28257 41075
rect 28211 41003 28217 41037
rect 28251 41003 28257 41037
rect 28211 40965 28257 41003
rect 28211 40931 28217 40965
rect 28251 40931 28257 40965
rect 28211 40893 28257 40931
rect 28211 40859 28217 40893
rect 28251 40859 28257 40893
rect 28211 40821 28257 40859
rect 28211 40787 28217 40821
rect 28251 40787 28257 40821
rect 28211 40749 28257 40787
rect 28211 40715 28217 40749
rect 28251 40715 28257 40749
rect 28211 40677 28257 40715
rect 28211 40643 28217 40677
rect 28251 40643 28257 40677
rect 28211 40605 28257 40643
rect 28211 40571 28217 40605
rect 28251 40571 28257 40605
rect 28211 40533 28257 40571
rect 28211 40499 28217 40533
rect 28251 40499 28257 40533
rect 28211 40461 28257 40499
rect 28211 40427 28217 40461
rect 28251 40427 28257 40461
rect 28211 40389 28257 40427
rect 28211 40355 28217 40389
rect 28251 40355 28257 40389
rect 28211 40317 28257 40355
rect 28211 40283 28217 40317
rect 28251 40283 28257 40317
rect 28211 40245 28257 40283
rect 28211 40211 28217 40245
rect 28251 40211 28257 40245
rect 28211 40173 28257 40211
rect 28211 40139 28217 40173
rect 28251 40139 28257 40173
rect 28211 40101 28257 40139
rect 28211 40067 28217 40101
rect 28251 40067 28257 40101
rect 28211 40029 28257 40067
rect 28211 39995 28217 40029
rect 28251 39995 28257 40029
rect 28211 39957 28257 39995
rect 29379 41181 29425 41197
rect 29379 41147 29385 41181
rect 29419 41147 29425 41181
rect 29379 41109 29425 41147
rect 29379 41075 29385 41109
rect 29419 41075 29425 41109
rect 29379 41037 29425 41075
rect 29379 41003 29385 41037
rect 29419 41003 29425 41037
rect 29379 40965 29425 41003
rect 29379 40931 29385 40965
rect 29419 40931 29425 40965
rect 29379 40893 29425 40931
rect 29379 40859 29385 40893
rect 29419 40859 29425 40893
rect 29379 40821 29425 40859
rect 29379 40787 29385 40821
rect 29419 40787 29425 40821
rect 29379 40749 29425 40787
rect 29379 40715 29385 40749
rect 29419 40715 29425 40749
rect 29379 40677 29425 40715
rect 29379 40643 29385 40677
rect 29419 40643 29425 40677
rect 29379 40605 29425 40643
rect 29379 40571 29385 40605
rect 29419 40571 29425 40605
rect 29379 40533 29425 40571
rect 29379 40499 29385 40533
rect 29419 40499 29425 40533
rect 29379 40461 29425 40499
rect 29379 40427 29385 40461
rect 29419 40427 29425 40461
rect 29379 40389 29425 40427
rect 29379 40355 29385 40389
rect 29419 40355 29425 40389
rect 29379 40317 29425 40355
rect 29379 40283 29385 40317
rect 29419 40283 29425 40317
rect 29379 40245 29425 40283
rect 29379 40211 29385 40245
rect 29419 40211 29425 40245
rect 29379 40173 29425 40211
rect 29379 40139 29385 40173
rect 29419 40139 29425 40173
rect 29379 40101 29425 40139
rect 29379 40067 29385 40101
rect 29419 40067 29425 40101
rect 29379 40029 29425 40067
rect 29379 39995 29385 40029
rect 29419 39995 29425 40029
rect 28211 39923 28217 39957
rect 28251 39923 28257 39957
rect 28350 39924 28356 39976
rect 28408 39964 28414 39976
rect 29379 39964 29425 39995
rect 29837 41181 29883 41197
rect 29837 41147 29843 41181
rect 29877 41147 29883 41181
rect 29837 41109 29883 41147
rect 29837 41075 29843 41109
rect 29877 41075 29883 41109
rect 29837 41037 29883 41075
rect 29837 41003 29843 41037
rect 29877 41003 29883 41037
rect 29837 40965 29883 41003
rect 29837 40931 29843 40965
rect 29877 40931 29883 40965
rect 29837 40893 29883 40931
rect 29837 40859 29843 40893
rect 29877 40859 29883 40893
rect 29837 40821 29883 40859
rect 29837 40787 29843 40821
rect 29877 40787 29883 40821
rect 29837 40749 29883 40787
rect 29837 40715 29843 40749
rect 29877 40715 29883 40749
rect 29837 40677 29883 40715
rect 29837 40643 29843 40677
rect 29877 40643 29883 40677
rect 29837 40605 29883 40643
rect 29837 40571 29843 40605
rect 29877 40571 29883 40605
rect 29837 40533 29883 40571
rect 29837 40499 29843 40533
rect 29877 40499 29883 40533
rect 29837 40461 29883 40499
rect 29837 40427 29843 40461
rect 29877 40427 29883 40461
rect 29837 40389 29883 40427
rect 29837 40355 29843 40389
rect 29877 40355 29883 40389
rect 29837 40317 29883 40355
rect 29837 40283 29843 40317
rect 29877 40283 29883 40317
rect 29837 40245 29883 40283
rect 29837 40211 29843 40245
rect 29877 40211 29883 40245
rect 29837 40173 29883 40211
rect 29837 40139 29843 40173
rect 29877 40139 29883 40173
rect 29837 40101 29883 40139
rect 29837 40067 29843 40101
rect 29877 40067 29883 40101
rect 29837 40029 29883 40067
rect 29837 39995 29843 40029
rect 29877 39995 29883 40029
rect 29837 39964 29883 39995
rect 28408 39957 29425 39964
rect 28408 39936 29385 39957
rect 28408 39924 28414 39936
rect 28211 39907 28257 39923
rect 29379 39923 29385 39936
rect 29419 39923 29425 39957
rect 29379 39907 29425 39923
rect 29472 39957 29883 39964
rect 29472 39936 29843 39957
rect 22186 39788 22192 39840
rect 22244 39828 22250 39840
rect 22741 39831 22799 39837
rect 22741 39828 22753 39831
rect 22244 39800 22753 39828
rect 22244 39788 22250 39800
rect 22741 39797 22753 39800
rect 22787 39797 22799 39831
rect 22741 39791 22799 39797
rect 23750 39788 23756 39840
rect 23808 39828 23814 39840
rect 28074 39828 28080 39840
rect 23808 39800 27936 39828
rect 28019 39800 28080 39828
rect 23808 39788 23814 39800
rect 27908 39760 27936 39800
rect 28074 39788 28080 39800
rect 28132 39788 28138 39840
rect 28166 39760 28172 39772
rect 27908 39732 28172 39760
rect 28166 39720 28172 39732
rect 28224 39720 28230 39772
rect 29472 39760 29500 39936
rect 29837 39923 29843 39936
rect 29877 39923 29883 39957
rect 29837 39907 29883 39923
rect 30295 41181 30341 41197
rect 30295 41147 30301 41181
rect 30335 41147 30341 41181
rect 30295 41109 30341 41147
rect 30295 41075 30301 41109
rect 30335 41075 30341 41109
rect 30295 41037 30341 41075
rect 30295 41003 30301 41037
rect 30335 41003 30341 41037
rect 30295 40965 30341 41003
rect 30295 40931 30301 40965
rect 30335 40931 30341 40965
rect 30295 40893 30341 40931
rect 30295 40859 30301 40893
rect 30335 40859 30341 40893
rect 30295 40821 30341 40859
rect 30295 40787 30301 40821
rect 30335 40787 30341 40821
rect 30295 40749 30341 40787
rect 30295 40715 30301 40749
rect 30335 40715 30341 40749
rect 30295 40677 30341 40715
rect 30295 40643 30301 40677
rect 30335 40643 30341 40677
rect 30295 40605 30341 40643
rect 30295 40571 30301 40605
rect 30335 40571 30341 40605
rect 30295 40533 30341 40571
rect 30295 40499 30301 40533
rect 30335 40499 30341 40533
rect 30295 40461 30341 40499
rect 30295 40427 30301 40461
rect 30335 40427 30341 40461
rect 30295 40389 30341 40427
rect 30295 40355 30301 40389
rect 30335 40355 30341 40389
rect 30295 40317 30341 40355
rect 30295 40283 30301 40317
rect 30335 40283 30341 40317
rect 30295 40245 30341 40283
rect 30295 40211 30301 40245
rect 30335 40211 30341 40245
rect 30295 40173 30341 40211
rect 30295 40139 30301 40173
rect 30335 40139 30341 40173
rect 30295 40101 30341 40139
rect 30295 40067 30301 40101
rect 30335 40067 30341 40101
rect 30295 40029 30341 40067
rect 30295 39995 30301 40029
rect 30335 39995 30341 40029
rect 30295 39957 30341 39995
rect 30295 39923 30301 39957
rect 30335 39923 30341 39957
rect 30295 39907 30341 39923
rect 30753 41181 30799 41197
rect 30753 41147 30759 41181
rect 30793 41147 30799 41181
rect 30753 41109 30799 41147
rect 30753 41075 30759 41109
rect 30793 41075 30799 41109
rect 30753 41037 30799 41075
rect 30753 41003 30759 41037
rect 30793 41003 30799 41037
rect 30753 40965 30799 41003
rect 30753 40931 30759 40965
rect 30793 40931 30799 40965
rect 30753 40893 30799 40931
rect 30753 40859 30759 40893
rect 30793 40859 30799 40893
rect 30753 40821 30799 40859
rect 30753 40787 30759 40821
rect 30793 40787 30799 40821
rect 30753 40749 30799 40787
rect 30753 40715 30759 40749
rect 30793 40715 30799 40749
rect 30753 40677 30799 40715
rect 30753 40643 30759 40677
rect 30793 40643 30799 40677
rect 30753 40605 30799 40643
rect 30753 40571 30759 40605
rect 30793 40571 30799 40605
rect 30753 40533 30799 40571
rect 30753 40499 30759 40533
rect 30793 40499 30799 40533
rect 30753 40461 30799 40499
rect 30753 40427 30759 40461
rect 30793 40427 30799 40461
rect 30753 40389 30799 40427
rect 30753 40355 30759 40389
rect 30793 40355 30799 40389
rect 30753 40317 30799 40355
rect 30753 40283 30759 40317
rect 30793 40283 30799 40317
rect 30753 40245 30799 40283
rect 30753 40211 30759 40245
rect 30793 40211 30799 40245
rect 30753 40173 30799 40211
rect 30753 40139 30759 40173
rect 30793 40139 30799 40173
rect 30753 40101 30799 40139
rect 30753 40067 30759 40101
rect 30793 40067 30799 40101
rect 30753 40029 30799 40067
rect 30753 39995 30759 40029
rect 30793 39995 30799 40029
rect 30753 39957 30799 39995
rect 30753 39923 30759 39957
rect 30793 39923 30799 39957
rect 30753 39907 30799 39923
rect 31211 41181 31257 41197
rect 31211 41147 31217 41181
rect 31251 41147 31257 41181
rect 31211 41109 31257 41147
rect 31211 41075 31217 41109
rect 31251 41075 31257 41109
rect 31211 41037 31257 41075
rect 31211 41003 31217 41037
rect 31251 41003 31257 41037
rect 31211 40965 31257 41003
rect 31211 40931 31217 40965
rect 31251 40931 31257 40965
rect 31211 40893 31257 40931
rect 31211 40859 31217 40893
rect 31251 40859 31257 40893
rect 31211 40821 31257 40859
rect 31211 40787 31217 40821
rect 31251 40787 31257 40821
rect 31211 40749 31257 40787
rect 31211 40715 31217 40749
rect 31251 40715 31257 40749
rect 31211 40677 31257 40715
rect 31211 40643 31217 40677
rect 31251 40643 31257 40677
rect 31211 40605 31257 40643
rect 31211 40571 31217 40605
rect 31251 40571 31257 40605
rect 31211 40533 31257 40571
rect 31211 40499 31217 40533
rect 31251 40499 31257 40533
rect 31211 40461 31257 40499
rect 31211 40427 31217 40461
rect 31251 40427 31257 40461
rect 31211 40389 31257 40427
rect 31211 40355 31217 40389
rect 31251 40355 31257 40389
rect 31211 40317 31257 40355
rect 31211 40283 31217 40317
rect 31251 40283 31257 40317
rect 31211 40245 31257 40283
rect 31211 40211 31217 40245
rect 31251 40211 31257 40245
rect 31211 40173 31257 40211
rect 31211 40139 31217 40173
rect 31251 40139 31257 40173
rect 31211 40101 31257 40139
rect 31211 40067 31217 40101
rect 31251 40067 31257 40101
rect 31211 40029 31257 40067
rect 31211 39995 31217 40029
rect 31251 39995 31257 40029
rect 31211 39957 31257 39995
rect 31211 39923 31217 39957
rect 31251 39923 31257 39957
rect 31211 39907 31257 39923
rect 31669 41181 31715 41197
rect 31669 41147 31675 41181
rect 31709 41147 31715 41181
rect 31669 41109 31715 41147
rect 31669 41075 31675 41109
rect 31709 41075 31715 41109
rect 31669 41037 31715 41075
rect 31669 41003 31675 41037
rect 31709 41003 31715 41037
rect 31669 40965 31715 41003
rect 31669 40931 31675 40965
rect 31709 40931 31715 40965
rect 31669 40893 31715 40931
rect 31669 40859 31675 40893
rect 31709 40859 31715 40893
rect 31669 40821 31715 40859
rect 31669 40787 31675 40821
rect 31709 40787 31715 40821
rect 31669 40749 31715 40787
rect 31669 40715 31675 40749
rect 31709 40715 31715 40749
rect 31669 40677 31715 40715
rect 31669 40643 31675 40677
rect 31709 40643 31715 40677
rect 31669 40605 31715 40643
rect 31669 40571 31675 40605
rect 31709 40571 31715 40605
rect 31669 40533 31715 40571
rect 31669 40499 31675 40533
rect 31709 40499 31715 40533
rect 31669 40461 31715 40499
rect 31669 40427 31675 40461
rect 31709 40427 31715 40461
rect 31669 40389 31715 40427
rect 31669 40355 31675 40389
rect 31709 40355 31715 40389
rect 31669 40317 31715 40355
rect 31669 40283 31675 40317
rect 31709 40283 31715 40317
rect 31669 40245 31715 40283
rect 31669 40211 31675 40245
rect 31709 40211 31715 40245
rect 31669 40173 31715 40211
rect 31669 40139 31675 40173
rect 31709 40139 31715 40173
rect 31669 40101 31715 40139
rect 31669 40067 31675 40101
rect 31709 40067 31715 40101
rect 31669 40029 31715 40067
rect 31669 39995 31675 40029
rect 31709 39995 31715 40029
rect 31669 39957 31715 39995
rect 31669 39923 31675 39957
rect 31709 39923 31715 39957
rect 31669 39907 31715 39923
rect 32127 41181 32173 41197
rect 32127 41147 32133 41181
rect 32167 41147 32173 41181
rect 32127 41109 32173 41147
rect 32127 41075 32133 41109
rect 32167 41075 32173 41109
rect 32127 41037 32173 41075
rect 32127 41003 32133 41037
rect 32167 41003 32173 41037
rect 32127 40965 32173 41003
rect 32127 40931 32133 40965
rect 32167 40931 32173 40965
rect 32127 40893 32173 40931
rect 32127 40859 32133 40893
rect 32167 40859 32173 40893
rect 32127 40821 32173 40859
rect 32127 40787 32133 40821
rect 32167 40787 32173 40821
rect 32127 40749 32173 40787
rect 32127 40715 32133 40749
rect 32167 40715 32173 40749
rect 32127 40677 32173 40715
rect 32127 40643 32133 40677
rect 32167 40643 32173 40677
rect 32127 40605 32173 40643
rect 32127 40571 32133 40605
rect 32167 40571 32173 40605
rect 32127 40533 32173 40571
rect 32127 40499 32133 40533
rect 32167 40499 32173 40533
rect 32127 40461 32173 40499
rect 32127 40427 32133 40461
rect 32167 40427 32173 40461
rect 32127 40389 32173 40427
rect 32127 40355 32133 40389
rect 32167 40355 32173 40389
rect 32127 40317 32173 40355
rect 32127 40283 32133 40317
rect 32167 40283 32173 40317
rect 32127 40245 32173 40283
rect 32127 40211 32133 40245
rect 32167 40211 32173 40245
rect 32127 40173 32173 40211
rect 32127 40139 32133 40173
rect 32167 40139 32173 40173
rect 32127 40101 32173 40139
rect 32127 40067 32133 40101
rect 32167 40067 32173 40101
rect 32127 40029 32173 40067
rect 32127 39995 32133 40029
rect 32167 39995 32173 40029
rect 32127 39957 32173 39995
rect 32127 39923 32133 39957
rect 32167 39923 32173 39957
rect 32127 39907 32173 39923
rect 32585 41181 32631 41197
rect 32585 41147 32591 41181
rect 32625 41147 32631 41181
rect 32585 41109 32631 41147
rect 32585 41075 32591 41109
rect 32625 41075 32631 41109
rect 32585 41037 32631 41075
rect 32585 41003 32591 41037
rect 32625 41003 32631 41037
rect 32585 40965 32631 41003
rect 32585 40931 32591 40965
rect 32625 40931 32631 40965
rect 32585 40893 32631 40931
rect 32585 40859 32591 40893
rect 32625 40859 32631 40893
rect 32585 40821 32631 40859
rect 32585 40787 32591 40821
rect 32625 40787 32631 40821
rect 32585 40749 32631 40787
rect 32585 40715 32591 40749
rect 32625 40715 32631 40749
rect 32585 40677 32631 40715
rect 32585 40643 32591 40677
rect 32625 40643 32631 40677
rect 32585 40605 32631 40643
rect 32585 40571 32591 40605
rect 32625 40571 32631 40605
rect 32585 40533 32631 40571
rect 32585 40499 32591 40533
rect 32625 40499 32631 40533
rect 32585 40461 32631 40499
rect 32585 40427 32591 40461
rect 32625 40427 32631 40461
rect 32585 40389 32631 40427
rect 32585 40355 32591 40389
rect 32625 40355 32631 40389
rect 32585 40317 32631 40355
rect 32585 40283 32591 40317
rect 32625 40283 32631 40317
rect 32585 40245 32631 40283
rect 32585 40211 32591 40245
rect 32625 40211 32631 40245
rect 32585 40173 32631 40211
rect 32585 40139 32591 40173
rect 32625 40139 32631 40173
rect 32585 40101 32631 40139
rect 32585 40067 32591 40101
rect 32625 40067 32631 40101
rect 32585 40029 32631 40067
rect 32585 39995 32591 40029
rect 32625 39995 32631 40029
rect 32585 39957 32631 39995
rect 32585 39923 32591 39957
rect 32625 39923 32631 39957
rect 32585 39907 32631 39923
rect 33043 41181 33089 41197
rect 33043 41147 33049 41181
rect 33083 41147 33089 41181
rect 33043 41109 33089 41147
rect 33043 41075 33049 41109
rect 33083 41075 33089 41109
rect 33043 41037 33089 41075
rect 33043 41003 33049 41037
rect 33083 41003 33089 41037
rect 33043 40965 33089 41003
rect 33043 40931 33049 40965
rect 33083 40931 33089 40965
rect 33043 40893 33089 40931
rect 33043 40859 33049 40893
rect 33083 40859 33089 40893
rect 33043 40821 33089 40859
rect 33043 40787 33049 40821
rect 33083 40787 33089 40821
rect 33043 40749 33089 40787
rect 33043 40715 33049 40749
rect 33083 40715 33089 40749
rect 33043 40677 33089 40715
rect 33043 40643 33049 40677
rect 33083 40643 33089 40677
rect 33043 40605 33089 40643
rect 33043 40571 33049 40605
rect 33083 40571 33089 40605
rect 33043 40533 33089 40571
rect 33043 40499 33049 40533
rect 33083 40499 33089 40533
rect 33043 40461 33089 40499
rect 33043 40427 33049 40461
rect 33083 40427 33089 40461
rect 33043 40389 33089 40427
rect 33043 40355 33049 40389
rect 33083 40355 33089 40389
rect 33043 40317 33089 40355
rect 33043 40283 33049 40317
rect 33083 40283 33089 40317
rect 33043 40245 33089 40283
rect 33043 40211 33049 40245
rect 33083 40211 33089 40245
rect 33043 40173 33089 40211
rect 33043 40139 33049 40173
rect 33083 40139 33089 40173
rect 33043 40101 33089 40139
rect 33043 40067 33049 40101
rect 33083 40067 33089 40101
rect 33043 40029 33089 40067
rect 33043 39995 33049 40029
rect 33083 39995 33089 40029
rect 33043 39957 33089 39995
rect 33043 39923 33049 39957
rect 33083 39923 33089 39957
rect 33043 39907 33089 39923
rect 33501 41181 33547 41197
rect 33501 41147 33507 41181
rect 33541 41147 33547 41181
rect 33501 41109 33547 41147
rect 33501 41075 33507 41109
rect 33541 41075 33547 41109
rect 33501 41037 33547 41075
rect 33501 41003 33507 41037
rect 33541 41003 33547 41037
rect 33501 40965 33547 41003
rect 33501 40931 33507 40965
rect 33541 40931 33547 40965
rect 33501 40893 33547 40931
rect 33501 40859 33507 40893
rect 33541 40859 33547 40893
rect 33501 40821 33547 40859
rect 33501 40787 33507 40821
rect 33541 40787 33547 40821
rect 33501 40749 33547 40787
rect 33501 40715 33507 40749
rect 33541 40715 33547 40749
rect 33501 40677 33547 40715
rect 33501 40643 33507 40677
rect 33541 40643 33547 40677
rect 33501 40605 33547 40643
rect 33501 40571 33507 40605
rect 33541 40571 33547 40605
rect 33501 40533 33547 40571
rect 33501 40499 33507 40533
rect 33541 40499 33547 40533
rect 33501 40461 33547 40499
rect 33501 40427 33507 40461
rect 33541 40427 33547 40461
rect 33501 40389 33547 40427
rect 33501 40355 33507 40389
rect 33541 40355 33547 40389
rect 33501 40317 33547 40355
rect 33501 40283 33507 40317
rect 33541 40283 33547 40317
rect 33501 40245 33547 40283
rect 33501 40211 33507 40245
rect 33541 40211 33547 40245
rect 33501 40173 33547 40211
rect 33501 40139 33507 40173
rect 33541 40139 33547 40173
rect 33501 40101 33547 40139
rect 33501 40067 33507 40101
rect 33541 40067 33547 40101
rect 33501 40029 33547 40067
rect 33501 39995 33507 40029
rect 33541 39995 33547 40029
rect 33501 39957 33547 39995
rect 33501 39923 33507 39957
rect 33541 39923 33547 39957
rect 33501 39907 33547 39923
rect 33959 41181 34005 41197
rect 33959 41147 33965 41181
rect 33999 41147 34005 41181
rect 33959 41109 34005 41147
rect 33959 41075 33965 41109
rect 33999 41075 34005 41109
rect 33959 41037 34005 41075
rect 33959 41003 33965 41037
rect 33999 41003 34005 41037
rect 33959 40965 34005 41003
rect 33959 40931 33965 40965
rect 33999 40931 34005 40965
rect 33959 40893 34005 40931
rect 33959 40859 33965 40893
rect 33999 40859 34005 40893
rect 33959 40821 34005 40859
rect 33959 40787 33965 40821
rect 33999 40787 34005 40821
rect 33959 40749 34005 40787
rect 33959 40715 33965 40749
rect 33999 40715 34005 40749
rect 33959 40677 34005 40715
rect 33959 40643 33965 40677
rect 33999 40643 34005 40677
rect 33959 40605 34005 40643
rect 33959 40571 33965 40605
rect 33999 40571 34005 40605
rect 33959 40533 34005 40571
rect 33959 40499 33965 40533
rect 33999 40499 34005 40533
rect 33959 40461 34005 40499
rect 33959 40427 33965 40461
rect 33999 40427 34005 40461
rect 33959 40389 34005 40427
rect 33959 40355 33965 40389
rect 33999 40355 34005 40389
rect 33959 40317 34005 40355
rect 33959 40283 33965 40317
rect 33999 40283 34005 40317
rect 33959 40245 34005 40283
rect 33959 40211 33965 40245
rect 33999 40211 34005 40245
rect 33959 40173 34005 40211
rect 33959 40139 33965 40173
rect 33999 40139 34005 40173
rect 33959 40101 34005 40139
rect 33959 40067 33965 40101
rect 33999 40067 34005 40101
rect 33959 40029 34005 40067
rect 33959 39995 33965 40029
rect 33999 39995 34005 40029
rect 33959 39957 34005 39995
rect 33959 39923 33965 39957
rect 33999 39923 34005 39957
rect 33959 39907 34005 39923
rect 34417 41181 34463 41197
rect 34417 41147 34423 41181
rect 34457 41147 34463 41181
rect 34417 41109 34463 41147
rect 34417 41075 34423 41109
rect 34457 41075 34463 41109
rect 34417 41037 34463 41075
rect 34417 41003 34423 41037
rect 34457 41003 34463 41037
rect 34417 40965 34463 41003
rect 34417 40931 34423 40965
rect 34457 40931 34463 40965
rect 34417 40893 34463 40931
rect 34417 40859 34423 40893
rect 34457 40859 34463 40893
rect 34417 40821 34463 40859
rect 34417 40787 34423 40821
rect 34457 40787 34463 40821
rect 34417 40749 34463 40787
rect 34417 40715 34423 40749
rect 34457 40715 34463 40749
rect 34417 40677 34463 40715
rect 34417 40643 34423 40677
rect 34457 40643 34463 40677
rect 34417 40605 34463 40643
rect 34417 40571 34423 40605
rect 34457 40571 34463 40605
rect 34417 40533 34463 40571
rect 34417 40499 34423 40533
rect 34457 40499 34463 40533
rect 34417 40461 34463 40499
rect 34417 40427 34423 40461
rect 34457 40427 34463 40461
rect 34417 40389 34463 40427
rect 34417 40355 34423 40389
rect 34457 40355 34463 40389
rect 34417 40317 34463 40355
rect 34417 40283 34423 40317
rect 34457 40283 34463 40317
rect 34417 40245 34463 40283
rect 34417 40211 34423 40245
rect 34457 40211 34463 40245
rect 34417 40173 34463 40211
rect 34417 40139 34423 40173
rect 34457 40139 34463 40173
rect 34417 40101 34463 40139
rect 34417 40067 34423 40101
rect 34457 40067 34463 40101
rect 34417 40029 34463 40067
rect 34417 39995 34423 40029
rect 34457 39995 34463 40029
rect 34417 39957 34463 39995
rect 34417 39923 34423 39957
rect 34457 39923 34463 39957
rect 34417 39907 34463 39923
rect 34875 41181 34921 41197
rect 34875 41147 34881 41181
rect 34915 41147 34921 41181
rect 34875 41109 34921 41147
rect 41966 41122 41972 41132
rect 34875 41075 34881 41109
rect 34915 41075 34921 41109
rect 34875 41037 34921 41075
rect 41810 41116 41972 41122
rect 42024 41122 42030 41132
rect 42024 41116 52478 41122
rect 41810 41082 41830 41116
rect 41864 41082 41920 41116
rect 41954 41082 41972 41116
rect 42044 41082 42100 41116
rect 42134 41082 42190 41116
rect 42224 41082 42280 41116
rect 42314 41082 42370 41116
rect 42404 41082 42460 41116
rect 42494 41082 42550 41116
rect 42584 41082 42640 41116
rect 42674 41082 42730 41116
rect 42764 41082 42820 41116
rect 42854 41082 42910 41116
rect 42944 41082 43000 41116
rect 43034 41082 43170 41116
rect 43204 41082 43260 41116
rect 43294 41082 43350 41116
rect 43384 41082 43440 41116
rect 43474 41082 43530 41116
rect 43564 41082 43620 41116
rect 43654 41082 43710 41116
rect 43744 41082 43800 41116
rect 43834 41082 43890 41116
rect 43924 41082 43980 41116
rect 44014 41082 44070 41116
rect 44104 41082 44160 41116
rect 44194 41082 44250 41116
rect 44284 41082 44340 41116
rect 44374 41082 44510 41116
rect 44544 41082 44600 41116
rect 44634 41082 44690 41116
rect 44724 41082 44780 41116
rect 44814 41082 44870 41116
rect 44904 41082 44960 41116
rect 44994 41082 45050 41116
rect 45084 41082 45140 41116
rect 45174 41082 45230 41116
rect 45264 41082 45320 41116
rect 45354 41082 45410 41116
rect 45444 41082 45500 41116
rect 45534 41082 45590 41116
rect 45624 41082 45680 41116
rect 45714 41082 45850 41116
rect 45884 41082 45940 41116
rect 45974 41082 46030 41116
rect 46064 41082 46120 41116
rect 46154 41082 46210 41116
rect 46244 41082 46300 41116
rect 46334 41082 46390 41116
rect 46424 41082 46480 41116
rect 46514 41082 46570 41116
rect 46604 41082 46660 41116
rect 46694 41082 46750 41116
rect 46784 41082 46840 41116
rect 46874 41082 46930 41116
rect 46964 41082 47020 41116
rect 47054 41082 47190 41116
rect 47224 41082 47280 41116
rect 47314 41082 47370 41116
rect 47404 41082 47460 41116
rect 47494 41082 47550 41116
rect 47584 41082 47640 41116
rect 47674 41082 47730 41116
rect 47764 41082 47820 41116
rect 47854 41082 47910 41116
rect 47944 41082 48000 41116
rect 48034 41082 48090 41116
rect 48124 41082 48180 41116
rect 48214 41082 48270 41116
rect 48304 41082 48360 41116
rect 48394 41082 48530 41116
rect 48564 41082 48620 41116
rect 48654 41082 48710 41116
rect 48744 41082 48800 41116
rect 48834 41082 48890 41116
rect 48924 41082 48980 41116
rect 49014 41082 49070 41116
rect 49104 41082 49160 41116
rect 49194 41082 49250 41116
rect 49284 41082 49340 41116
rect 49374 41082 49430 41116
rect 49464 41082 49520 41116
rect 49554 41082 49610 41116
rect 49644 41082 49700 41116
rect 49734 41082 49870 41116
rect 49904 41082 49960 41116
rect 49994 41082 50050 41116
rect 50084 41082 50140 41116
rect 50174 41082 50230 41116
rect 50264 41082 50320 41116
rect 50354 41082 50410 41116
rect 50444 41082 50500 41116
rect 50534 41082 50590 41116
rect 50624 41082 50680 41116
rect 50714 41082 50770 41116
rect 50804 41082 50860 41116
rect 50894 41082 50950 41116
rect 50984 41082 51040 41116
rect 51074 41082 51210 41116
rect 51244 41082 51300 41116
rect 51334 41082 51390 41116
rect 51424 41082 51480 41116
rect 51514 41082 51570 41116
rect 51604 41082 51660 41116
rect 51694 41082 51750 41116
rect 51784 41082 51840 41116
rect 51874 41082 51930 41116
rect 51964 41082 52020 41116
rect 52054 41082 52110 41116
rect 52144 41082 52200 41116
rect 52234 41082 52290 41116
rect 52324 41082 52380 41116
rect 52414 41082 52478 41116
rect 41810 41080 41972 41082
rect 42024 41080 52478 41082
rect 41810 41052 52478 41080
rect 34875 41003 34881 41037
rect 34915 41003 34921 41037
rect 34875 40965 34921 41003
rect 34875 40931 34881 40965
rect 34915 40931 34921 40965
rect 41974 40956 52314 40972
rect 34875 40893 34921 40931
rect 34875 40859 34881 40893
rect 34915 40859 34921 40893
rect 34875 40821 34921 40859
rect 34875 40787 34881 40821
rect 34915 40787 34921 40821
rect 34875 40749 34921 40787
rect 34875 40715 34881 40749
rect 34915 40715 34921 40749
rect 34875 40677 34921 40715
rect 34875 40643 34881 40677
rect 34915 40643 34921 40677
rect 34875 40605 34921 40643
rect 34875 40571 34881 40605
rect 34915 40571 34921 40605
rect 34875 40533 34921 40571
rect 34875 40499 34881 40533
rect 34915 40499 34921 40533
rect 34875 40461 34921 40499
rect 34875 40427 34881 40461
rect 34915 40427 34921 40461
rect 34875 40389 34921 40427
rect 34875 40355 34881 40389
rect 34915 40355 34921 40389
rect 34875 40317 34921 40355
rect 34875 40283 34881 40317
rect 34915 40283 34921 40317
rect 34875 40245 34921 40283
rect 34875 40211 34881 40245
rect 34915 40211 34921 40245
rect 34875 40173 34921 40211
rect 34875 40139 34881 40173
rect 34915 40139 34921 40173
rect 37282 40929 37328 40952
rect 37282 40895 37288 40929
rect 37322 40895 37328 40929
rect 37282 40857 37328 40895
rect 37282 40823 37288 40857
rect 37322 40823 37328 40857
rect 37282 40785 37328 40823
rect 37282 40751 37288 40785
rect 37322 40751 37328 40785
rect 37282 40713 37328 40751
rect 37282 40679 37288 40713
rect 37322 40679 37328 40713
rect 37282 40641 37328 40679
rect 37282 40607 37288 40641
rect 37322 40607 37328 40641
rect 37282 40569 37328 40607
rect 37282 40535 37288 40569
rect 37322 40535 37328 40569
rect 37282 40497 37328 40535
rect 37282 40463 37288 40497
rect 37322 40463 37328 40497
rect 37282 40425 37328 40463
rect 37282 40391 37288 40425
rect 37322 40391 37328 40425
rect 37282 40353 37328 40391
rect 37282 40319 37288 40353
rect 37322 40319 37328 40353
rect 37282 40281 37328 40319
rect 37282 40247 37288 40281
rect 37322 40247 37328 40281
rect 37282 40209 37328 40247
rect 37282 40175 37288 40209
rect 37322 40175 37328 40209
rect 37282 40152 37328 40175
rect 37740 40929 37786 40952
rect 37740 40895 37746 40929
rect 37780 40895 37786 40929
rect 37740 40857 37786 40895
rect 37740 40823 37746 40857
rect 37780 40823 37786 40857
rect 37740 40785 37786 40823
rect 37740 40751 37746 40785
rect 37780 40751 37786 40785
rect 37740 40713 37786 40751
rect 37740 40679 37746 40713
rect 37780 40679 37786 40713
rect 37740 40641 37786 40679
rect 37740 40607 37746 40641
rect 37780 40607 37786 40641
rect 37740 40569 37786 40607
rect 37740 40535 37746 40569
rect 37780 40535 37786 40569
rect 37740 40497 37786 40535
rect 37740 40463 37746 40497
rect 37780 40463 37786 40497
rect 37740 40425 37786 40463
rect 37740 40391 37746 40425
rect 37780 40391 37786 40425
rect 37740 40353 37786 40391
rect 37740 40319 37746 40353
rect 37780 40319 37786 40353
rect 37740 40281 37786 40319
rect 37740 40247 37746 40281
rect 37780 40247 37786 40281
rect 37740 40209 37786 40247
rect 37740 40175 37746 40209
rect 37780 40175 37786 40209
rect 37740 40152 37786 40175
rect 38198 40929 38244 40952
rect 38198 40895 38204 40929
rect 38238 40895 38244 40929
rect 38198 40857 38244 40895
rect 38198 40823 38204 40857
rect 38238 40823 38244 40857
rect 38198 40785 38244 40823
rect 38198 40751 38204 40785
rect 38238 40751 38244 40785
rect 38198 40713 38244 40751
rect 38198 40679 38204 40713
rect 38238 40679 38244 40713
rect 38198 40641 38244 40679
rect 38198 40607 38204 40641
rect 38238 40607 38244 40641
rect 38198 40569 38244 40607
rect 38198 40535 38204 40569
rect 38238 40535 38244 40569
rect 38198 40497 38244 40535
rect 38198 40463 38204 40497
rect 38238 40463 38244 40497
rect 38198 40425 38244 40463
rect 38198 40391 38204 40425
rect 38238 40391 38244 40425
rect 38198 40353 38244 40391
rect 38198 40319 38204 40353
rect 38238 40319 38244 40353
rect 38198 40281 38244 40319
rect 38198 40247 38204 40281
rect 38238 40247 38244 40281
rect 38656 40929 38702 40952
rect 38656 40895 38662 40929
rect 38696 40895 38702 40929
rect 38656 40857 38702 40895
rect 38656 40823 38662 40857
rect 38696 40823 38702 40857
rect 38656 40785 38702 40823
rect 38656 40751 38662 40785
rect 38696 40751 38702 40785
rect 38656 40713 38702 40751
rect 38656 40679 38662 40713
rect 38696 40679 38702 40713
rect 38656 40641 38702 40679
rect 38656 40607 38662 40641
rect 38696 40607 38702 40641
rect 38656 40569 38702 40607
rect 38656 40535 38662 40569
rect 38696 40535 38702 40569
rect 38656 40497 38702 40535
rect 38656 40463 38662 40497
rect 38696 40463 38702 40497
rect 38656 40425 38702 40463
rect 38656 40391 38662 40425
rect 38696 40391 38702 40425
rect 38656 40353 38702 40391
rect 38656 40319 38662 40353
rect 38696 40319 38702 40353
rect 38656 40281 38702 40319
rect 38198 40236 38244 40247
rect 38562 40236 38568 40248
rect 38198 40209 38568 40236
rect 38198 40175 38204 40209
rect 38238 40208 38568 40209
rect 38238 40175 38244 40208
rect 38562 40196 38568 40208
rect 38620 40196 38626 40248
rect 38656 40247 38662 40281
rect 38696 40247 38702 40281
rect 38656 40209 38702 40247
rect 38198 40152 38244 40175
rect 38656 40175 38662 40209
rect 38696 40175 38702 40209
rect 38656 40152 38702 40175
rect 39114 40929 39160 40952
rect 39114 40895 39120 40929
rect 39154 40895 39160 40929
rect 39114 40857 39160 40895
rect 39114 40823 39120 40857
rect 39154 40823 39160 40857
rect 39114 40785 39160 40823
rect 39114 40751 39120 40785
rect 39154 40751 39160 40785
rect 39114 40713 39160 40751
rect 39114 40679 39120 40713
rect 39154 40679 39160 40713
rect 39114 40641 39160 40679
rect 39114 40607 39120 40641
rect 39154 40607 39160 40641
rect 39114 40569 39160 40607
rect 39114 40535 39120 40569
rect 39154 40535 39160 40569
rect 39114 40497 39160 40535
rect 39114 40463 39120 40497
rect 39154 40463 39160 40497
rect 39114 40425 39160 40463
rect 39114 40391 39120 40425
rect 39154 40391 39160 40425
rect 39114 40353 39160 40391
rect 39114 40319 39120 40353
rect 39154 40319 39160 40353
rect 39114 40281 39160 40319
rect 39114 40247 39120 40281
rect 39154 40247 39160 40281
rect 39114 40209 39160 40247
rect 39114 40175 39120 40209
rect 39154 40175 39160 40209
rect 39114 40152 39160 40175
rect 39572 40929 39618 40952
rect 39572 40895 39578 40929
rect 39612 40895 39618 40929
rect 39572 40857 39618 40895
rect 39572 40823 39578 40857
rect 39612 40823 39618 40857
rect 39572 40785 39618 40823
rect 39572 40751 39578 40785
rect 39612 40751 39618 40785
rect 39572 40713 39618 40751
rect 39572 40679 39578 40713
rect 39612 40679 39618 40713
rect 39572 40641 39618 40679
rect 39572 40607 39578 40641
rect 39612 40607 39618 40641
rect 39572 40569 39618 40607
rect 39572 40535 39578 40569
rect 39612 40535 39618 40569
rect 39572 40497 39618 40535
rect 39572 40463 39578 40497
rect 39612 40463 39618 40497
rect 39572 40425 39618 40463
rect 39572 40391 39578 40425
rect 39612 40391 39618 40425
rect 39572 40353 39618 40391
rect 39572 40319 39578 40353
rect 39612 40319 39618 40353
rect 39572 40281 39618 40319
rect 39572 40247 39578 40281
rect 39612 40247 39618 40281
rect 39572 40209 39618 40247
rect 39572 40175 39578 40209
rect 39612 40175 39618 40209
rect 39572 40152 39618 40175
rect 40030 40929 40076 40952
rect 40030 40895 40036 40929
rect 40070 40895 40076 40929
rect 40030 40857 40076 40895
rect 40030 40823 40036 40857
rect 40070 40823 40076 40857
rect 40030 40785 40076 40823
rect 40030 40751 40036 40785
rect 40070 40751 40076 40785
rect 40030 40713 40076 40751
rect 40030 40679 40036 40713
rect 40070 40679 40076 40713
rect 40030 40641 40076 40679
rect 40030 40607 40036 40641
rect 40070 40607 40076 40641
rect 40030 40569 40076 40607
rect 40030 40535 40036 40569
rect 40070 40535 40076 40569
rect 40030 40497 40076 40535
rect 40030 40463 40036 40497
rect 40070 40463 40076 40497
rect 40030 40425 40076 40463
rect 40030 40391 40036 40425
rect 40070 40391 40076 40425
rect 40030 40353 40076 40391
rect 40030 40319 40036 40353
rect 40070 40319 40076 40353
rect 40030 40281 40076 40319
rect 40030 40247 40036 40281
rect 40070 40247 40076 40281
rect 40030 40209 40076 40247
rect 40030 40175 40036 40209
rect 40070 40175 40076 40209
rect 40030 40152 40076 40175
rect 40488 40929 40534 40952
rect 40488 40895 40494 40929
rect 40528 40895 40534 40929
rect 40488 40857 40534 40895
rect 40488 40823 40494 40857
rect 40528 40823 40534 40857
rect 40488 40785 40534 40823
rect 40488 40751 40494 40785
rect 40528 40751 40534 40785
rect 40488 40713 40534 40751
rect 40488 40679 40494 40713
rect 40528 40679 40534 40713
rect 40488 40641 40534 40679
rect 40488 40607 40494 40641
rect 40528 40607 40534 40641
rect 40488 40569 40534 40607
rect 40488 40535 40494 40569
rect 40528 40535 40534 40569
rect 40488 40497 40534 40535
rect 40488 40463 40494 40497
rect 40528 40463 40534 40497
rect 40488 40425 40534 40463
rect 40488 40391 40494 40425
rect 40528 40391 40534 40425
rect 40488 40353 40534 40391
rect 40488 40319 40494 40353
rect 40528 40319 40534 40353
rect 40488 40281 40534 40319
rect 40488 40247 40494 40281
rect 40528 40247 40534 40281
rect 40488 40209 40534 40247
rect 40488 40175 40494 40209
rect 40528 40175 40534 40209
rect 40488 40152 40534 40175
rect 40946 40929 40992 40952
rect 40946 40895 40952 40929
rect 40986 40895 40992 40929
rect 40946 40857 40992 40895
rect 40946 40823 40952 40857
rect 40986 40823 40992 40857
rect 40946 40785 40992 40823
rect 40946 40751 40952 40785
rect 40986 40751 40992 40785
rect 40946 40713 40992 40751
rect 40946 40679 40952 40713
rect 40986 40679 40992 40713
rect 40946 40641 40992 40679
rect 40946 40607 40952 40641
rect 40986 40607 40992 40641
rect 40946 40569 40992 40607
rect 40946 40535 40952 40569
rect 40986 40535 40992 40569
rect 40946 40497 40992 40535
rect 40946 40463 40952 40497
rect 40986 40463 40992 40497
rect 40946 40425 40992 40463
rect 40946 40391 40952 40425
rect 40986 40391 40992 40425
rect 40946 40353 40992 40391
rect 40946 40319 40952 40353
rect 40986 40319 40992 40353
rect 40946 40281 40992 40319
rect 40946 40247 40952 40281
rect 40986 40247 40992 40281
rect 40946 40209 40992 40247
rect 40946 40175 40952 40209
rect 40986 40175 40992 40209
rect 40946 40152 40992 40175
rect 41404 40929 41450 40952
rect 41404 40895 41410 40929
rect 41444 40895 41450 40929
rect 41974 40928 41994 40956
rect 41404 40857 41450 40895
rect 41966 40876 41972 40928
rect 42028 40922 42084 40956
rect 42118 40922 42174 40956
rect 42208 40922 42264 40956
rect 42298 40922 42354 40956
rect 42388 40922 42444 40956
rect 42478 40922 42534 40956
rect 42568 40922 42624 40956
rect 42658 40922 42714 40956
rect 42748 40922 42804 40956
rect 42838 40922 42894 40956
rect 42928 40922 43334 40956
rect 43368 40922 43424 40956
rect 43458 40922 43514 40956
rect 43548 40922 43604 40956
rect 43638 40922 43694 40956
rect 43728 40922 43784 40956
rect 43818 40922 43874 40956
rect 43908 40922 43964 40956
rect 43998 40922 44054 40956
rect 44088 40922 44144 40956
rect 44178 40922 44234 40956
rect 44268 40922 44674 40956
rect 44708 40922 44764 40956
rect 44798 40922 44854 40956
rect 44888 40922 44944 40956
rect 44978 40922 45034 40956
rect 45068 40922 45124 40956
rect 45158 40922 45214 40956
rect 45248 40922 45304 40956
rect 45338 40922 45394 40956
rect 45428 40922 45484 40956
rect 45518 40922 45574 40956
rect 45608 40922 46014 40956
rect 46048 40922 46104 40956
rect 46138 40922 46194 40956
rect 46228 40922 46284 40956
rect 46318 40922 46374 40956
rect 46408 40922 46464 40956
rect 46498 40922 46554 40956
rect 46588 40922 46644 40956
rect 46678 40922 46734 40956
rect 46768 40922 46824 40956
rect 46858 40922 46914 40956
rect 46948 40922 47354 40956
rect 47388 40922 47444 40956
rect 47478 40922 47534 40956
rect 47568 40922 47624 40956
rect 47658 40922 47714 40956
rect 47748 40922 47804 40956
rect 47838 40922 47894 40956
rect 47928 40922 47984 40956
rect 48018 40922 48074 40956
rect 48108 40922 48164 40956
rect 48198 40922 48254 40956
rect 48288 40922 48694 40956
rect 48728 40922 48784 40956
rect 48818 40922 48874 40956
rect 48908 40922 48964 40956
rect 48998 40922 49054 40956
rect 49088 40922 49144 40956
rect 49178 40922 49234 40956
rect 49268 40922 49324 40956
rect 49358 40922 49414 40956
rect 49448 40922 49504 40956
rect 49538 40922 49594 40956
rect 49628 40922 50034 40956
rect 50068 40922 50124 40956
rect 50158 40922 50214 40956
rect 50248 40922 50304 40956
rect 50338 40922 50394 40956
rect 50428 40922 50484 40956
rect 50518 40922 50574 40956
rect 50608 40922 50664 40956
rect 50698 40922 50754 40956
rect 50788 40922 50844 40956
rect 50878 40922 50934 40956
rect 50968 40922 51374 40956
rect 51408 40922 51464 40956
rect 51498 40922 51554 40956
rect 51588 40922 51644 40956
rect 51678 40922 51734 40956
rect 51768 40922 51824 40956
rect 51858 40922 51914 40956
rect 51948 40922 52004 40956
rect 52038 40922 52094 40956
rect 52128 40922 52184 40956
rect 52218 40922 52274 40956
rect 52308 40922 52314 40956
rect 42024 40902 52314 40922
rect 42024 40876 42030 40902
rect 41404 40823 41410 40857
rect 41444 40823 41450 40857
rect 41404 40785 41450 40823
rect 41404 40751 41410 40785
rect 41444 40751 41450 40785
rect 41404 40713 41450 40751
rect 41404 40679 41410 40713
rect 41444 40679 41450 40713
rect 41404 40641 41450 40679
rect 41404 40607 41410 40641
rect 41444 40607 41450 40641
rect 41404 40569 41450 40607
rect 41404 40535 41410 40569
rect 41444 40535 41450 40569
rect 41404 40497 41450 40535
rect 41404 40463 41410 40497
rect 41444 40463 41450 40497
rect 41404 40425 41450 40463
rect 41404 40391 41410 40425
rect 41444 40391 41450 40425
rect 41404 40353 41450 40391
rect 41404 40319 41410 40353
rect 41444 40319 41450 40353
rect 41404 40281 41450 40319
rect 41404 40247 41410 40281
rect 41444 40247 41450 40281
rect 41404 40209 41450 40247
rect 41404 40175 41410 40209
rect 41444 40175 41450 40209
rect 42148 40792 52140 40798
rect 42148 40752 44088 40792
rect 42148 40718 42180 40752
rect 42214 40718 42280 40752
rect 42314 40718 42380 40752
rect 42414 40718 42480 40752
rect 42514 40718 42580 40752
rect 42614 40718 42680 40752
rect 42714 40718 43520 40752
rect 43554 40718 43620 40752
rect 43654 40718 43720 40752
rect 43754 40718 43820 40752
rect 43854 40718 43920 40752
rect 43954 40718 44020 40752
rect 44054 40740 44088 40752
rect 44140 40752 52140 40792
rect 44140 40740 44860 40752
rect 44054 40718 44860 40740
rect 44894 40718 44960 40752
rect 44994 40718 45060 40752
rect 45094 40718 45160 40752
rect 45194 40718 45260 40752
rect 45294 40718 45360 40752
rect 45394 40718 46200 40752
rect 46234 40718 46300 40752
rect 46334 40718 46400 40752
rect 46434 40718 46500 40752
rect 46534 40718 46600 40752
rect 46634 40718 46700 40752
rect 46734 40718 47540 40752
rect 47574 40718 47640 40752
rect 47674 40718 47740 40752
rect 47774 40718 47840 40752
rect 47874 40718 47940 40752
rect 47974 40718 48040 40752
rect 48074 40718 48880 40752
rect 48914 40718 48980 40752
rect 49014 40718 49080 40752
rect 49114 40718 49180 40752
rect 49214 40718 49280 40752
rect 49314 40718 49380 40752
rect 49414 40718 50220 40752
rect 50254 40718 50320 40752
rect 50354 40718 50420 40752
rect 50454 40718 50520 40752
rect 50554 40718 50620 40752
rect 50654 40718 50720 40752
rect 50754 40718 51560 40752
rect 51594 40718 51660 40752
rect 51694 40718 51760 40752
rect 51794 40718 51860 40752
rect 51894 40718 51960 40752
rect 51994 40718 52060 40752
rect 52094 40718 52140 40752
rect 42148 40652 52140 40718
rect 42148 40618 42180 40652
rect 42214 40618 42280 40652
rect 42314 40618 42380 40652
rect 42414 40618 42480 40652
rect 42514 40618 42580 40652
rect 42614 40618 42680 40652
rect 42714 40618 43520 40652
rect 43554 40618 43620 40652
rect 43654 40618 43720 40652
rect 43754 40618 43820 40652
rect 43854 40618 43920 40652
rect 43954 40618 44020 40652
rect 44054 40618 44860 40652
rect 44894 40618 44960 40652
rect 44994 40618 45060 40652
rect 45094 40618 45160 40652
rect 45194 40618 45260 40652
rect 45294 40618 45360 40652
rect 45394 40618 46200 40652
rect 46234 40618 46300 40652
rect 46334 40618 46400 40652
rect 46434 40618 46500 40652
rect 46534 40618 46600 40652
rect 46634 40618 46700 40652
rect 46734 40618 47540 40652
rect 47574 40618 47640 40652
rect 47674 40618 47740 40652
rect 47774 40618 47840 40652
rect 47874 40618 47940 40652
rect 47974 40618 48040 40652
rect 48074 40618 48880 40652
rect 48914 40618 48980 40652
rect 49014 40618 49080 40652
rect 49114 40618 49180 40652
rect 49214 40618 49280 40652
rect 49314 40618 49380 40652
rect 49414 40618 50220 40652
rect 50254 40618 50320 40652
rect 50354 40618 50420 40652
rect 50454 40618 50520 40652
rect 50554 40618 50620 40652
rect 50654 40618 50720 40652
rect 50754 40618 51560 40652
rect 51594 40618 51660 40652
rect 51694 40618 51760 40652
rect 51794 40618 51860 40652
rect 51894 40618 51960 40652
rect 51994 40618 52060 40652
rect 52094 40618 52140 40652
rect 42148 40552 52140 40618
rect 42148 40518 42180 40552
rect 42214 40518 42280 40552
rect 42314 40518 42380 40552
rect 42414 40518 42480 40552
rect 42514 40518 42580 40552
rect 42614 40518 42680 40552
rect 42714 40518 43520 40552
rect 43554 40518 43620 40552
rect 43654 40518 43720 40552
rect 43754 40518 43820 40552
rect 43854 40518 43920 40552
rect 43954 40518 44020 40552
rect 44054 40518 44860 40552
rect 44894 40518 44960 40552
rect 44994 40518 45060 40552
rect 45094 40518 45160 40552
rect 45194 40518 45260 40552
rect 45294 40518 45360 40552
rect 45394 40518 46200 40552
rect 46234 40518 46300 40552
rect 46334 40518 46400 40552
rect 46434 40518 46500 40552
rect 46534 40518 46600 40552
rect 46634 40518 46700 40552
rect 46734 40518 47540 40552
rect 47574 40518 47640 40552
rect 47674 40518 47740 40552
rect 47774 40518 47840 40552
rect 47874 40518 47940 40552
rect 47974 40518 48040 40552
rect 48074 40518 48880 40552
rect 48914 40518 48980 40552
rect 49014 40518 49080 40552
rect 49114 40518 49180 40552
rect 49214 40518 49280 40552
rect 49314 40518 49380 40552
rect 49414 40518 50220 40552
rect 50254 40518 50320 40552
rect 50354 40518 50420 40552
rect 50454 40518 50520 40552
rect 50554 40518 50620 40552
rect 50654 40518 50720 40552
rect 50754 40518 51560 40552
rect 51594 40518 51660 40552
rect 51694 40518 51760 40552
rect 51794 40518 51860 40552
rect 51894 40518 51960 40552
rect 51994 40518 52060 40552
rect 52094 40518 52140 40552
rect 42148 40452 52140 40518
rect 42148 40418 42180 40452
rect 42214 40418 42280 40452
rect 42314 40418 42380 40452
rect 42414 40418 42480 40452
rect 42514 40418 42580 40452
rect 42614 40418 42680 40452
rect 42714 40418 43520 40452
rect 43554 40418 43620 40452
rect 43654 40418 43720 40452
rect 43754 40418 43820 40452
rect 43854 40418 43920 40452
rect 43954 40418 44020 40452
rect 44054 40418 44860 40452
rect 44894 40418 44960 40452
rect 44994 40418 45060 40452
rect 45094 40418 45160 40452
rect 45194 40418 45260 40452
rect 45294 40418 45360 40452
rect 45394 40418 46200 40452
rect 46234 40418 46300 40452
rect 46334 40418 46400 40452
rect 46434 40418 46500 40452
rect 46534 40418 46600 40452
rect 46634 40418 46700 40452
rect 46734 40418 47540 40452
rect 47574 40418 47640 40452
rect 47674 40418 47740 40452
rect 47774 40418 47840 40452
rect 47874 40418 47940 40452
rect 47974 40418 48040 40452
rect 48074 40418 48880 40452
rect 48914 40418 48980 40452
rect 49014 40418 49080 40452
rect 49114 40418 49180 40452
rect 49214 40418 49280 40452
rect 49314 40418 49380 40452
rect 49414 40418 50220 40452
rect 50254 40418 50320 40452
rect 50354 40418 50420 40452
rect 50454 40418 50520 40452
rect 50554 40418 50620 40452
rect 50654 40418 50720 40452
rect 50754 40418 51560 40452
rect 51594 40418 51660 40452
rect 51694 40418 51760 40452
rect 51794 40418 51860 40452
rect 51894 40418 51960 40452
rect 51994 40418 52060 40452
rect 52094 40418 52140 40452
rect 42148 40352 52140 40418
rect 42148 40318 42180 40352
rect 42214 40318 42280 40352
rect 42314 40318 42380 40352
rect 42414 40318 42480 40352
rect 42514 40318 42580 40352
rect 42614 40318 42680 40352
rect 42714 40318 43520 40352
rect 43554 40318 43620 40352
rect 43654 40318 43720 40352
rect 43754 40318 43820 40352
rect 43854 40318 43920 40352
rect 43954 40318 44020 40352
rect 44054 40318 44860 40352
rect 44894 40318 44960 40352
rect 44994 40318 45060 40352
rect 45094 40318 45160 40352
rect 45194 40318 45260 40352
rect 45294 40318 45360 40352
rect 45394 40318 46200 40352
rect 46234 40318 46300 40352
rect 46334 40318 46400 40352
rect 46434 40318 46500 40352
rect 46534 40318 46600 40352
rect 46634 40318 46700 40352
rect 46734 40318 47540 40352
rect 47574 40318 47640 40352
rect 47674 40318 47740 40352
rect 47774 40318 47840 40352
rect 47874 40318 47940 40352
rect 47974 40318 48040 40352
rect 48074 40318 48880 40352
rect 48914 40318 48980 40352
rect 49014 40318 49080 40352
rect 49114 40318 49180 40352
rect 49214 40318 49280 40352
rect 49314 40318 49380 40352
rect 49414 40318 50220 40352
rect 50254 40318 50320 40352
rect 50354 40318 50420 40352
rect 50454 40318 50520 40352
rect 50554 40318 50620 40352
rect 50654 40318 50720 40352
rect 50754 40318 51560 40352
rect 51594 40318 51660 40352
rect 51694 40318 51760 40352
rect 51794 40318 51860 40352
rect 51894 40318 51960 40352
rect 51994 40318 52060 40352
rect 52094 40318 52140 40352
rect 42148 40252 52140 40318
rect 42148 40248 42180 40252
rect 42148 40196 42156 40248
rect 42214 40218 42280 40252
rect 42314 40218 42380 40252
rect 42414 40218 42480 40252
rect 42514 40218 42580 40252
rect 42614 40218 42680 40252
rect 42714 40218 43520 40252
rect 43554 40218 43620 40252
rect 43654 40218 43720 40252
rect 43754 40218 43820 40252
rect 43854 40218 43920 40252
rect 43954 40218 44020 40252
rect 44054 40218 44860 40252
rect 44894 40218 44960 40252
rect 44994 40218 45060 40252
rect 45094 40218 45160 40252
rect 45194 40218 45260 40252
rect 45294 40218 45360 40252
rect 45394 40218 46200 40252
rect 46234 40218 46300 40252
rect 46334 40218 46400 40252
rect 46434 40218 46500 40252
rect 46534 40218 46600 40252
rect 46634 40218 46700 40252
rect 46734 40218 47540 40252
rect 47574 40218 47640 40252
rect 47674 40218 47740 40252
rect 47774 40218 47840 40252
rect 47874 40218 47940 40252
rect 47974 40218 48040 40252
rect 48074 40218 48880 40252
rect 48914 40218 48980 40252
rect 49014 40218 49080 40252
rect 49114 40218 49180 40252
rect 49214 40218 49280 40252
rect 49314 40218 49380 40252
rect 49414 40218 50220 40252
rect 50254 40218 50320 40252
rect 50354 40218 50420 40252
rect 50454 40218 50520 40252
rect 50554 40218 50620 40252
rect 50654 40218 50720 40252
rect 50754 40218 51560 40252
rect 51594 40218 51660 40252
rect 51694 40218 51760 40252
rect 51794 40218 51860 40252
rect 51894 40218 51960 40252
rect 51994 40218 52060 40252
rect 52094 40218 52140 40252
rect 42208 40196 52140 40218
rect 42148 40186 52140 40196
rect 41404 40152 41450 40175
rect 34875 40101 34921 40139
rect 34875 40067 34881 40101
rect 34915 40067 34921 40101
rect 34875 40029 34921 40067
rect 35802 40060 35808 40112
rect 35860 40100 35866 40112
rect 37752 40100 37780 40152
rect 35860 40072 37780 40100
rect 35860 40060 35866 40072
rect 34875 39995 34881 40029
rect 34915 39995 34921 40029
rect 34875 39957 34921 39995
rect 34875 39923 34881 39957
rect 34915 39923 34921 39957
rect 34875 39907 34921 39923
rect 41417 39899 41475 39905
rect 41417 39865 41429 39899
rect 41463 39896 41475 39899
rect 48314 39896 48320 39908
rect 41463 39868 48320 39896
rect 41463 39865 41475 39868
rect 41417 39859 41475 39865
rect 48314 39856 48320 39868
rect 48372 39856 48378 39908
rect 28276 39732 29500 39760
rect 28276 39701 28304 39732
rect 28261 39695 28319 39701
rect 28261 39661 28273 39695
rect 28307 39661 28319 39695
rect 29454 39692 29460 39704
rect 29399 39664 29460 39692
rect 28261 39655 28319 39661
rect 29454 39652 29460 39664
rect 29512 39652 29518 39704
rect 900 39610 57536 39612
rect 900 39494 922 39610
rect 2510 39569 55926 39610
rect 2510 39535 6493 39569
rect 6527 39535 6893 39569
rect 6927 39535 7293 39569
rect 7327 39535 7693 39569
rect 7727 39535 8093 39569
rect 8127 39535 8493 39569
rect 8527 39535 8893 39569
rect 8927 39535 9293 39569
rect 9327 39535 9693 39569
rect 9727 39535 10093 39569
rect 10127 39535 10493 39569
rect 10527 39535 10893 39569
rect 10927 39535 11293 39569
rect 11327 39535 11693 39569
rect 11727 39535 12093 39569
rect 12127 39535 12493 39569
rect 12527 39535 12893 39569
rect 12927 39535 13293 39569
rect 13327 39535 15313 39569
rect 15347 39568 15713 39569
rect 15347 39535 15476 39568
rect 2510 39516 15476 39535
rect 15528 39535 15713 39568
rect 15747 39535 16113 39569
rect 16147 39535 16513 39569
rect 16547 39535 16913 39569
rect 16947 39535 17313 39569
rect 17347 39535 17713 39569
rect 17747 39535 18113 39569
rect 18147 39535 18513 39569
rect 18547 39535 18913 39569
rect 18947 39535 19313 39569
rect 19347 39535 19713 39569
rect 19747 39535 20113 39569
rect 20147 39535 20513 39569
rect 20547 39535 20913 39569
rect 20947 39535 21313 39569
rect 21347 39535 21713 39569
rect 21747 39535 22113 39569
rect 22147 39535 22857 39569
rect 22891 39535 23257 39569
rect 23291 39535 23657 39569
rect 23691 39535 24057 39569
rect 24091 39535 24457 39569
rect 24491 39535 24857 39569
rect 24891 39535 25257 39569
rect 25291 39535 25657 39569
rect 25691 39535 26057 39569
rect 26091 39535 26457 39569
rect 26491 39535 26857 39569
rect 26891 39535 27257 39569
rect 27291 39535 27657 39569
rect 27691 39535 28057 39569
rect 28091 39535 29521 39569
rect 29555 39535 29921 39569
rect 29955 39535 30321 39569
rect 30355 39535 30721 39569
rect 30755 39535 31121 39569
rect 31155 39535 31521 39569
rect 31555 39535 31921 39569
rect 31955 39535 32321 39569
rect 32355 39535 32721 39569
rect 32755 39535 33121 39569
rect 33155 39535 33521 39569
rect 33555 39535 33921 39569
rect 33955 39535 34321 39569
rect 34355 39535 34721 39569
rect 34755 39535 37459 39569
rect 37493 39535 37859 39569
rect 37893 39535 38259 39569
rect 38293 39535 38659 39569
rect 38693 39535 39059 39569
rect 39093 39535 39459 39569
rect 39493 39535 39859 39569
rect 39893 39535 40259 39569
rect 40293 39535 40659 39569
rect 40693 39535 41059 39569
rect 41093 39535 41967 39569
rect 42001 39568 42167 39569
rect 42024 39535 42167 39568
rect 42201 39535 42367 39569
rect 42401 39535 42567 39569
rect 42601 39535 42767 39569
rect 42801 39535 42967 39569
rect 43001 39535 43167 39569
rect 43201 39535 43367 39569
rect 43401 39535 43567 39569
rect 43601 39535 43767 39569
rect 43801 39535 43967 39569
rect 44001 39535 44167 39569
rect 44201 39535 44367 39569
rect 44401 39535 44567 39569
rect 44601 39535 44767 39569
rect 44801 39535 44967 39569
rect 45001 39535 45167 39569
rect 45201 39535 45367 39569
rect 45401 39535 45567 39569
rect 45601 39535 45767 39569
rect 45801 39535 45967 39569
rect 46001 39535 46167 39569
rect 46201 39535 46367 39569
rect 46401 39535 46567 39569
rect 46601 39535 46767 39569
rect 46801 39535 46967 39569
rect 47001 39535 47167 39569
rect 47201 39535 47367 39569
rect 47401 39535 47567 39569
rect 47601 39535 47767 39569
rect 47801 39535 47967 39569
rect 48001 39535 48167 39569
rect 48201 39535 48367 39569
rect 48401 39535 48567 39569
rect 48601 39535 48767 39569
rect 48801 39535 48967 39569
rect 49001 39535 49167 39569
rect 49201 39535 49367 39569
rect 49401 39535 49567 39569
rect 49601 39535 49767 39569
rect 49801 39535 49967 39569
rect 50001 39535 50167 39569
rect 50201 39535 50367 39569
rect 50401 39535 50567 39569
rect 50601 39535 50767 39569
rect 50801 39535 50967 39569
rect 51001 39535 51167 39569
rect 51201 39535 51367 39569
rect 51401 39535 51567 39569
rect 51601 39535 51767 39569
rect 51801 39535 51967 39569
rect 52001 39535 52167 39569
rect 52201 39535 52367 39569
rect 52401 39535 55926 39569
rect 15528 39516 41972 39535
rect 42024 39516 55926 39535
rect 2510 39494 55926 39516
rect 57514 39494 57536 39610
rect 900 39492 57536 39494
rect 14366 38088 14372 38140
rect 14424 38088 14430 38140
rect 14384 38060 14412 38088
rect 25774 38060 25780 38072
rect 14384 38032 25780 38060
rect 25774 38020 25780 38032
rect 25832 38020 25838 38072
rect 34422 37952 34428 38004
rect 34480 37992 34486 38004
rect 35802 37992 35808 38004
rect 34480 37964 35808 37992
rect 34480 37952 34486 37964
rect 35802 37952 35808 37964
rect 35860 37952 35866 38004
rect 3348 37730 55088 37732
rect 3348 37614 3370 37730
rect 4958 37689 53478 37730
rect 4958 37655 12175 37689
rect 12209 37655 12375 37689
rect 12409 37655 12575 37689
rect 12609 37655 12775 37689
rect 12809 37655 12975 37689
rect 13009 37655 13175 37689
rect 13209 37655 13861 37689
rect 13895 37655 14061 37689
rect 14095 37655 14261 37689
rect 14295 37655 14461 37689
rect 14495 37655 14661 37689
rect 14695 37655 14861 37689
rect 14895 37655 15061 37689
rect 15095 37655 15261 37689
rect 15295 37655 15461 37689
rect 15495 37655 15661 37689
rect 15695 37655 15861 37689
rect 15895 37655 16605 37689
rect 16639 37655 16805 37689
rect 16839 37655 17005 37689
rect 17039 37655 17205 37689
rect 17239 37655 17405 37689
rect 17439 37655 17605 37689
rect 17639 37655 17805 37689
rect 17839 37655 18005 37689
rect 18039 37655 18205 37689
rect 18239 37655 18405 37689
rect 18439 37655 18605 37689
rect 18639 37655 19351 37689
rect 19385 37655 19551 37689
rect 19585 37655 19751 37689
rect 19785 37655 19951 37689
rect 19985 37655 20151 37689
rect 20185 37655 20351 37689
rect 20385 37655 20551 37689
rect 20585 37655 20751 37689
rect 20785 37655 20951 37689
rect 20985 37655 21151 37689
rect 21185 37655 21351 37689
rect 21385 37655 21551 37689
rect 21585 37655 21751 37689
rect 21785 37655 21951 37689
rect 21985 37655 22681 37689
rect 22715 37655 22881 37689
rect 22915 37655 23081 37689
rect 23115 37655 23281 37689
rect 23315 37655 23481 37689
rect 23515 37655 23681 37689
rect 23715 37655 23881 37689
rect 23915 37655 24081 37689
rect 24115 37655 24281 37689
rect 24315 37655 24481 37689
rect 24515 37655 24681 37689
rect 24715 37655 25601 37689
rect 25635 37655 26001 37689
rect 26035 37655 26401 37689
rect 26435 37655 26801 37689
rect 26835 37655 27201 37689
rect 27235 37655 27601 37689
rect 27635 37655 28001 37689
rect 28035 37655 28401 37689
rect 28435 37655 28801 37689
rect 28835 37655 29201 37689
rect 29235 37655 30111 37689
rect 30145 37655 30511 37689
rect 30545 37655 30911 37689
rect 30945 37655 31311 37689
rect 31345 37655 31711 37689
rect 31745 37655 32111 37689
rect 32145 37655 32511 37689
rect 32545 37655 32911 37689
rect 32945 37655 33311 37689
rect 33345 37664 33711 37689
rect 33345 37655 33416 37664
rect 4958 37614 33416 37655
rect 3348 37612 33416 37614
rect 33468 37655 33711 37664
rect 33745 37655 34111 37689
rect 34145 37655 34511 37689
rect 34545 37655 34911 37689
rect 34945 37655 35311 37689
rect 35345 37655 35711 37689
rect 35745 37655 36111 37689
rect 36145 37655 36511 37689
rect 36545 37655 36911 37689
rect 36945 37655 37655 37689
rect 37689 37655 38055 37689
rect 38089 37655 38455 37689
rect 38489 37655 38855 37689
rect 38889 37655 39255 37689
rect 39289 37655 39655 37689
rect 39689 37655 40055 37689
rect 40089 37655 41967 37689
rect 42001 37655 42167 37689
rect 42201 37655 42367 37689
rect 42401 37655 42567 37689
rect 42601 37655 42767 37689
rect 42801 37655 42967 37689
rect 43001 37655 43167 37689
rect 43201 37655 43367 37689
rect 43401 37655 43567 37689
rect 43601 37655 43767 37689
rect 43801 37655 43967 37689
rect 44001 37655 44167 37689
rect 44201 37655 44367 37689
rect 44401 37655 44567 37689
rect 44601 37655 44767 37689
rect 44801 37655 44967 37689
rect 45001 37655 45167 37689
rect 45201 37655 45367 37689
rect 45401 37655 45567 37689
rect 45601 37655 45767 37689
rect 45801 37655 45967 37689
rect 46001 37655 46167 37689
rect 46201 37655 46367 37689
rect 46401 37655 46567 37689
rect 46601 37655 46767 37689
rect 46801 37655 46967 37689
rect 47001 37655 47167 37689
rect 47201 37655 47367 37689
rect 47401 37655 47567 37689
rect 47601 37655 47767 37689
rect 47801 37655 47967 37689
rect 48001 37655 48167 37689
rect 48201 37655 48367 37689
rect 48401 37655 48567 37689
rect 48601 37655 48767 37689
rect 48801 37655 48967 37689
rect 49001 37655 49167 37689
rect 49201 37655 49367 37689
rect 49401 37655 49567 37689
rect 49601 37655 49767 37689
rect 49801 37655 49967 37689
rect 50001 37655 50167 37689
rect 50201 37655 50367 37689
rect 50401 37655 50567 37689
rect 50601 37655 50767 37689
rect 50801 37655 50967 37689
rect 51001 37655 51167 37689
rect 51201 37655 51367 37689
rect 51401 37655 51567 37689
rect 51601 37655 51767 37689
rect 51801 37655 51967 37689
rect 52001 37655 52167 37689
rect 52201 37655 52367 37689
rect 52401 37655 53478 37689
rect 33468 37614 53478 37655
rect 55066 37614 55088 37730
rect 33468 37612 55088 37614
rect 22278 37516 22284 37528
rect 21652 37488 22284 37516
rect 13689 37421 14099 37433
rect 12894 37136 12900 37188
rect 12952 37136 12958 37188
rect 12912 37037 12940 37136
rect 12357 36992 12967 37037
rect 12357 36958 12388 36992
rect 12422 36958 12488 36992
rect 12522 36958 12588 36992
rect 12622 36958 12688 36992
rect 12722 36958 12788 36992
rect 12822 36958 12888 36992
rect 12922 36958 12967 36992
rect 12357 36892 12967 36958
rect 12357 36858 12388 36892
rect 12422 36858 12488 36892
rect 12522 36858 12588 36892
rect 12622 36858 12688 36892
rect 12722 36858 12788 36892
rect 12822 36858 12888 36892
rect 12922 36858 12967 36892
rect 13689 36883 13697 37421
rect 14091 36904 14099 37421
rect 15697 37421 16107 37433
rect 15562 36904 15568 36916
rect 14091 36883 15568 36904
rect 13689 36876 15568 36883
rect 13689 36871 14099 36876
rect 15562 36864 15568 36876
rect 15620 36864 15626 36916
rect 15697 36883 15704 37421
rect 16098 36883 16107 37421
rect 15697 36871 16107 36883
rect 16433 37421 16843 37433
rect 16433 36883 16441 37421
rect 16835 36883 16843 37421
rect 16433 36871 16580 36883
rect 12357 36792 12967 36858
rect 12357 36758 12388 36792
rect 12422 36758 12488 36792
rect 12522 36758 12588 36792
rect 12622 36758 12688 36792
rect 12722 36758 12788 36792
rect 12822 36758 12888 36792
rect 12922 36758 12967 36792
rect 12357 36692 12967 36758
rect 12357 36658 12388 36692
rect 12422 36658 12488 36692
rect 12522 36658 12588 36692
rect 12622 36658 12688 36692
rect 12722 36658 12788 36692
rect 12822 36658 12888 36692
rect 12922 36658 12967 36692
rect 12357 36592 12967 36658
rect 12357 36558 12388 36592
rect 12422 36558 12488 36592
rect 12522 36558 12588 36592
rect 12622 36558 12688 36592
rect 12722 36558 12788 36592
rect 12822 36558 12888 36592
rect 12922 36558 12967 36592
rect 12357 36492 12967 36558
rect 12357 36458 12388 36492
rect 12422 36458 12488 36492
rect 12522 36458 12588 36492
rect 12622 36458 12688 36492
rect 12722 36458 12788 36492
rect 12822 36458 12888 36492
rect 12922 36458 12967 36492
rect 12357 36427 12967 36458
rect 13689 36461 14099 36473
rect 13081 36295 13139 36301
rect 13081 36261 13093 36295
rect 13127 36261 13139 36295
rect 13081 36255 13139 36261
rect 13096 36156 13124 36255
rect 13265 36159 13323 36165
rect 13265 36156 13277 36159
rect 13096 36128 13277 36156
rect 13265 36125 13277 36128
rect 13311 36125 13323 36159
rect 13265 36119 13323 36125
rect 13280 35852 13308 36119
rect 13689 35923 13697 36461
rect 14091 35923 14099 36461
rect 13689 35912 13912 35923
rect 13964 35912 14099 35923
rect 13689 35911 14099 35912
rect 15686 36461 16118 36871
rect 16574 36864 16580 36871
rect 16632 36871 16843 36883
rect 18441 37421 18851 37433
rect 18441 36883 18448 37421
rect 18842 36883 18851 37421
rect 18441 36871 18851 36883
rect 19178 37421 19588 37433
rect 19178 36883 19186 37421
rect 19580 37380 19588 37421
rect 21652 37380 21680 37488
rect 22278 37476 22284 37488
rect 22336 37476 22342 37528
rect 37568 37525 37596 37612
rect 37553 37519 37611 37525
rect 37553 37485 37565 37519
rect 37599 37485 37611 37519
rect 37553 37479 37611 37485
rect 19580 37352 21680 37380
rect 21760 37421 22170 37433
rect 19580 36883 19588 37352
rect 19178 36871 19588 36883
rect 21760 36883 21767 37421
rect 22161 36883 22170 37421
rect 22509 37421 22919 37433
rect 21760 36871 22170 36883
rect 16632 36864 16638 36871
rect 15686 35923 15704 36461
rect 16098 35923 16118 36461
rect 16433 36461 16843 36473
rect 16206 36388 16212 36440
rect 16264 36428 16270 36440
rect 16433 36428 16441 36461
rect 16264 36400 16441 36428
rect 16264 36388 16270 36400
rect 15686 35907 16118 35923
rect 16433 35923 16441 36400
rect 16835 35923 16843 36461
rect 16433 35911 16843 35923
rect 18430 36461 18862 36871
rect 18430 35923 18448 36461
rect 18842 35923 18862 36461
rect 18430 35907 18862 35923
rect 19178 36461 19588 36473
rect 19178 35923 19186 36461
rect 19580 35923 19588 36461
rect 19178 35911 19588 35923
rect 21749 36461 22181 36871
rect 22370 36864 22376 36916
rect 22428 36904 22434 36916
rect 22509 36904 22517 37421
rect 22428 36883 22517 36904
rect 22911 36883 22919 37421
rect 22428 36876 22919 36883
rect 22428 36864 22434 36876
rect 22509 36871 22919 36876
rect 24517 37421 24927 37433
rect 24517 36883 24524 37421
rect 24918 36883 24927 37421
rect 37513 37421 37559 37437
rect 37513 37387 37519 37421
rect 37553 37387 37559 37421
rect 37513 37349 37559 37387
rect 37513 37315 37519 37349
rect 37553 37315 37559 37349
rect 37513 37277 37559 37315
rect 37513 37243 37519 37277
rect 37553 37243 37559 37277
rect 37513 37205 37559 37243
rect 24517 36871 24927 36883
rect 25424 37169 25470 37192
rect 25424 37135 25430 37169
rect 25464 37135 25470 37169
rect 25774 37136 25780 37188
rect 25832 37176 25838 37188
rect 25882 37176 25928 37192
rect 25832 37169 25928 37176
rect 25832 37148 25888 37169
rect 25832 37136 25838 37148
rect 25424 37097 25470 37135
rect 25424 37063 25430 37097
rect 25464 37063 25470 37097
rect 25424 37025 25470 37063
rect 25424 36991 25430 37025
rect 25464 36991 25470 37025
rect 25424 36953 25470 36991
rect 25424 36919 25430 36953
rect 25464 36919 25470 36953
rect 25424 36881 25470 36919
rect 21749 35923 21767 36461
rect 22161 35923 22181 36461
rect 22509 36461 22919 36473
rect 22278 36388 22284 36440
rect 22336 36428 22342 36440
rect 22509 36428 22517 36461
rect 22336 36400 22517 36428
rect 22336 36388 22342 36400
rect 19260 35852 19288 35911
rect 21749 35907 22181 35923
rect 22509 35923 22517 36400
rect 22911 35923 22919 36461
rect 22509 35911 22919 35923
rect 24506 36461 24938 36871
rect 24506 35923 24524 36461
rect 24918 35923 24938 36461
rect 25424 36847 25430 36881
rect 25464 36847 25470 36881
rect 25424 36809 25470 36847
rect 25424 36775 25430 36809
rect 25464 36775 25470 36809
rect 25424 36737 25470 36775
rect 25424 36703 25430 36737
rect 25464 36703 25470 36737
rect 25424 36665 25470 36703
rect 25424 36631 25430 36665
rect 25464 36631 25470 36665
rect 25424 36593 25470 36631
rect 25424 36559 25430 36593
rect 25464 36559 25470 36593
rect 25424 36521 25470 36559
rect 25424 36487 25430 36521
rect 25464 36487 25470 36521
rect 25424 36449 25470 36487
rect 25424 36415 25430 36449
rect 25464 36415 25470 36449
rect 25424 36392 25470 36415
rect 25882 37135 25888 37148
rect 25922 37135 25928 37169
rect 25882 37097 25928 37135
rect 25882 37063 25888 37097
rect 25922 37063 25928 37097
rect 25882 37025 25928 37063
rect 25882 36991 25888 37025
rect 25922 36991 25928 37025
rect 25882 36953 25928 36991
rect 25882 36919 25888 36953
rect 25922 36919 25928 36953
rect 25882 36881 25928 36919
rect 25882 36847 25888 36881
rect 25922 36847 25928 36881
rect 25882 36809 25928 36847
rect 25882 36775 25888 36809
rect 25922 36775 25928 36809
rect 25882 36737 25928 36775
rect 25882 36703 25888 36737
rect 25922 36703 25928 36737
rect 25882 36665 25928 36703
rect 25882 36631 25888 36665
rect 25922 36631 25928 36665
rect 25882 36593 25928 36631
rect 25882 36559 25888 36593
rect 25922 36559 25928 36593
rect 25882 36521 25928 36559
rect 25882 36487 25888 36521
rect 25922 36487 25928 36521
rect 25882 36449 25928 36487
rect 25882 36415 25888 36449
rect 25922 36415 25928 36449
rect 25882 36392 25928 36415
rect 26340 37169 26386 37192
rect 26340 37135 26346 37169
rect 26380 37135 26386 37169
rect 26340 37097 26386 37135
rect 26340 37063 26346 37097
rect 26380 37063 26386 37097
rect 26340 37025 26386 37063
rect 26340 36991 26346 37025
rect 26380 36991 26386 37025
rect 26340 36953 26386 36991
rect 26340 36919 26346 36953
rect 26380 36919 26386 36953
rect 26340 36881 26386 36919
rect 26340 36847 26346 36881
rect 26380 36847 26386 36881
rect 26340 36809 26386 36847
rect 26340 36775 26346 36809
rect 26380 36775 26386 36809
rect 26340 36737 26386 36775
rect 26340 36703 26346 36737
rect 26380 36703 26386 36737
rect 26340 36665 26386 36703
rect 26340 36631 26346 36665
rect 26380 36631 26386 36665
rect 26340 36593 26386 36631
rect 26340 36559 26346 36593
rect 26380 36559 26386 36593
rect 26340 36521 26386 36559
rect 26340 36487 26346 36521
rect 26380 36487 26386 36521
rect 26340 36449 26386 36487
rect 26340 36415 26346 36449
rect 26380 36415 26386 36449
rect 26340 36392 26386 36415
rect 26798 37169 26844 37192
rect 26798 37135 26804 37169
rect 26838 37135 26844 37169
rect 26798 37097 26844 37135
rect 26798 37063 26804 37097
rect 26838 37063 26844 37097
rect 26798 37025 26844 37063
rect 26798 36991 26804 37025
rect 26838 36991 26844 37025
rect 26798 36953 26844 36991
rect 26798 36919 26804 36953
rect 26838 36919 26844 36953
rect 26798 36881 26844 36919
rect 26798 36847 26804 36881
rect 26838 36847 26844 36881
rect 26798 36809 26844 36847
rect 26798 36775 26804 36809
rect 26838 36775 26844 36809
rect 26798 36737 26844 36775
rect 26798 36703 26804 36737
rect 26838 36703 26844 36737
rect 26798 36665 26844 36703
rect 26798 36631 26804 36665
rect 26838 36631 26844 36665
rect 26798 36593 26844 36631
rect 26798 36559 26804 36593
rect 26838 36559 26844 36593
rect 26798 36521 26844 36559
rect 26798 36487 26804 36521
rect 26838 36487 26844 36521
rect 26798 36449 26844 36487
rect 26798 36415 26804 36449
rect 26838 36415 26844 36449
rect 26798 36392 26844 36415
rect 27256 37169 27302 37192
rect 27256 37135 27262 37169
rect 27296 37135 27302 37169
rect 27256 37097 27302 37135
rect 27256 37063 27262 37097
rect 27296 37063 27302 37097
rect 27256 37025 27302 37063
rect 27256 36991 27262 37025
rect 27296 36991 27302 37025
rect 27256 36953 27302 36991
rect 27256 36919 27262 36953
rect 27296 36919 27302 36953
rect 27256 36881 27302 36919
rect 27256 36847 27262 36881
rect 27296 36847 27302 36881
rect 27256 36809 27302 36847
rect 27256 36775 27262 36809
rect 27296 36775 27302 36809
rect 27256 36737 27302 36775
rect 27256 36703 27262 36737
rect 27296 36703 27302 36737
rect 27256 36665 27302 36703
rect 27256 36631 27262 36665
rect 27296 36631 27302 36665
rect 27256 36593 27302 36631
rect 27256 36559 27262 36593
rect 27296 36559 27302 36593
rect 27256 36521 27302 36559
rect 27256 36487 27262 36521
rect 27296 36487 27302 36521
rect 27256 36449 27302 36487
rect 27256 36415 27262 36449
rect 27296 36415 27302 36449
rect 27256 36392 27302 36415
rect 27714 37169 27760 37192
rect 27714 37135 27720 37169
rect 27754 37135 27760 37169
rect 27714 37097 27760 37135
rect 27714 37063 27720 37097
rect 27754 37063 27760 37097
rect 27714 37025 27760 37063
rect 27714 36991 27720 37025
rect 27754 36991 27760 37025
rect 27714 36953 27760 36991
rect 27714 36919 27720 36953
rect 27754 36919 27760 36953
rect 27714 36881 27760 36919
rect 27714 36847 27720 36881
rect 27754 36847 27760 36881
rect 27714 36809 27760 36847
rect 27714 36775 27720 36809
rect 27754 36775 27760 36809
rect 27714 36737 27760 36775
rect 27714 36703 27720 36737
rect 27754 36703 27760 36737
rect 27714 36665 27760 36703
rect 27714 36631 27720 36665
rect 27754 36631 27760 36665
rect 27714 36593 27760 36631
rect 27714 36559 27720 36593
rect 27754 36559 27760 36593
rect 27714 36521 27760 36559
rect 27714 36487 27720 36521
rect 27754 36487 27760 36521
rect 27714 36449 27760 36487
rect 27714 36415 27720 36449
rect 27754 36415 27760 36449
rect 27714 36392 27760 36415
rect 28172 37169 28218 37192
rect 28172 37135 28178 37169
rect 28212 37135 28218 37169
rect 28172 37097 28218 37135
rect 28172 37063 28178 37097
rect 28212 37063 28218 37097
rect 28172 37025 28218 37063
rect 28172 36991 28178 37025
rect 28212 36991 28218 37025
rect 28172 36953 28218 36991
rect 28172 36919 28178 36953
rect 28212 36919 28218 36953
rect 28172 36881 28218 36919
rect 28172 36847 28178 36881
rect 28212 36847 28218 36881
rect 28172 36809 28218 36847
rect 28172 36775 28178 36809
rect 28212 36775 28218 36809
rect 28172 36737 28218 36775
rect 28172 36703 28178 36737
rect 28212 36703 28218 36737
rect 28172 36665 28218 36703
rect 28172 36631 28178 36665
rect 28212 36631 28218 36665
rect 28172 36593 28218 36631
rect 28172 36559 28178 36593
rect 28212 36559 28218 36593
rect 28172 36521 28218 36559
rect 28172 36487 28178 36521
rect 28212 36487 28218 36521
rect 28172 36449 28218 36487
rect 28172 36415 28178 36449
rect 28212 36415 28218 36449
rect 28172 36392 28218 36415
rect 28630 37169 28676 37192
rect 28630 37135 28636 37169
rect 28670 37135 28676 37169
rect 28630 37097 28676 37135
rect 28630 37063 28636 37097
rect 28670 37063 28676 37097
rect 28630 37025 28676 37063
rect 28630 36991 28636 37025
rect 28670 36991 28676 37025
rect 28630 36953 28676 36991
rect 28630 36919 28636 36953
rect 28670 36919 28676 36953
rect 28630 36881 28676 36919
rect 28630 36847 28636 36881
rect 28670 36847 28676 36881
rect 28630 36809 28676 36847
rect 28630 36775 28636 36809
rect 28670 36775 28676 36809
rect 28630 36737 28676 36775
rect 28630 36703 28636 36737
rect 28670 36703 28676 36737
rect 28630 36665 28676 36703
rect 28630 36631 28636 36665
rect 28670 36631 28676 36665
rect 28630 36593 28676 36631
rect 28630 36559 28636 36593
rect 28670 36559 28676 36593
rect 28630 36521 28676 36559
rect 28630 36487 28636 36521
rect 28670 36487 28676 36521
rect 28630 36449 28676 36487
rect 28630 36415 28636 36449
rect 28670 36415 28676 36449
rect 28630 36392 28676 36415
rect 29088 37169 29134 37192
rect 29088 37135 29094 37169
rect 29128 37135 29134 37169
rect 29088 37097 29134 37135
rect 29088 37063 29094 37097
rect 29128 37063 29134 37097
rect 29088 37025 29134 37063
rect 29088 36991 29094 37025
rect 29128 36991 29134 37025
rect 29088 36972 29134 36991
rect 29546 37176 29592 37192
rect 34422 37176 34428 37188
rect 29546 37169 34428 37176
rect 29546 37135 29552 37169
rect 29586 37148 34428 37169
rect 29586 37135 29592 37148
rect 34422 37136 34428 37148
rect 34480 37136 34486 37188
rect 37513 37171 37519 37205
rect 37553 37171 37559 37205
rect 29546 37097 29592 37135
rect 29546 37063 29552 37097
rect 29586 37063 29592 37097
rect 29546 37025 29592 37063
rect 29546 36991 29552 37025
rect 29586 36991 29592 37025
rect 29454 36972 29460 36984
rect 29088 36953 29460 36972
rect 29088 36919 29094 36953
rect 29128 36944 29460 36953
rect 29128 36919 29134 36944
rect 29454 36932 29460 36944
rect 29512 36932 29518 36984
rect 29546 36953 29592 36991
rect 29088 36881 29134 36919
rect 29088 36847 29094 36881
rect 29128 36847 29134 36881
rect 29088 36809 29134 36847
rect 29088 36775 29094 36809
rect 29128 36775 29134 36809
rect 29088 36737 29134 36775
rect 29088 36703 29094 36737
rect 29128 36703 29134 36737
rect 29088 36665 29134 36703
rect 29088 36631 29094 36665
rect 29128 36631 29134 36665
rect 29088 36593 29134 36631
rect 29088 36559 29094 36593
rect 29128 36559 29134 36593
rect 29088 36521 29134 36559
rect 29088 36487 29094 36521
rect 29128 36487 29134 36521
rect 29088 36449 29134 36487
rect 29088 36415 29094 36449
rect 29128 36415 29134 36449
rect 29088 36392 29134 36415
rect 29546 36919 29552 36953
rect 29586 36919 29592 36953
rect 29546 36881 29592 36919
rect 29546 36847 29552 36881
rect 29586 36847 29592 36881
rect 29546 36809 29592 36847
rect 29546 36775 29552 36809
rect 29586 36775 29592 36809
rect 29546 36737 29592 36775
rect 29546 36703 29552 36737
rect 29586 36703 29592 36737
rect 29546 36665 29592 36703
rect 29546 36631 29552 36665
rect 29586 36631 29592 36665
rect 29546 36593 29592 36631
rect 29546 36559 29552 36593
rect 29586 36559 29592 36593
rect 29546 36521 29592 36559
rect 29546 36487 29552 36521
rect 29586 36487 29592 36521
rect 29546 36449 29592 36487
rect 29546 36415 29552 36449
rect 29586 36415 29592 36449
rect 29546 36392 29592 36415
rect 37513 37133 37559 37171
rect 37513 37099 37519 37133
rect 37553 37099 37559 37133
rect 37513 37061 37559 37099
rect 37513 37027 37519 37061
rect 37553 37027 37559 37061
rect 37513 36989 37559 37027
rect 37513 36955 37519 36989
rect 37553 36955 37559 36989
rect 37513 36917 37559 36955
rect 37513 36883 37519 36917
rect 37553 36883 37559 36917
rect 37513 36845 37559 36883
rect 37513 36811 37519 36845
rect 37553 36811 37559 36845
rect 37513 36773 37559 36811
rect 37513 36739 37519 36773
rect 37553 36739 37559 36773
rect 37513 36701 37559 36739
rect 37513 36667 37519 36701
rect 37553 36667 37559 36701
rect 37513 36629 37559 36667
rect 37513 36595 37519 36629
rect 37553 36595 37559 36629
rect 37513 36557 37559 36595
rect 37513 36523 37519 36557
rect 37553 36523 37559 36557
rect 37513 36485 37559 36523
rect 37513 36451 37519 36485
rect 37553 36451 37559 36485
rect 37513 36413 37559 36451
rect 37513 36379 37519 36413
rect 37553 36379 37559 36413
rect 37513 36341 37559 36379
rect 37513 36307 37519 36341
rect 37553 36307 37559 36341
rect 37513 36269 37559 36307
rect 37513 36235 37519 36269
rect 37553 36235 37559 36269
rect 37513 36197 37559 36235
rect 28074 36156 28080 36168
rect 28019 36128 28080 36156
rect 28074 36116 28080 36128
rect 28132 36116 28138 36168
rect 37513 36163 37519 36197
rect 37553 36163 37559 36197
rect 37513 36147 37559 36163
rect 37971 37421 38017 37437
rect 37971 37387 37977 37421
rect 38011 37387 38017 37421
rect 37971 37349 38017 37387
rect 37971 37315 37977 37349
rect 38011 37315 38017 37349
rect 37971 37277 38017 37315
rect 37971 37243 37977 37277
rect 38011 37243 38017 37277
rect 37971 37205 38017 37243
rect 37971 37171 37977 37205
rect 38011 37171 38017 37205
rect 37971 37133 38017 37171
rect 37971 37099 37977 37133
rect 38011 37099 38017 37133
rect 37971 37061 38017 37099
rect 37971 37027 37977 37061
rect 38011 37027 38017 37061
rect 37971 36989 38017 37027
rect 37971 36955 37977 36989
rect 38011 36955 38017 36989
rect 37971 36917 38017 36955
rect 37971 36883 37977 36917
rect 38011 36883 38017 36917
rect 37971 36845 38017 36883
rect 37971 36811 37977 36845
rect 38011 36811 38017 36845
rect 37971 36773 38017 36811
rect 37971 36739 37977 36773
rect 38011 36739 38017 36773
rect 37971 36701 38017 36739
rect 37971 36667 37977 36701
rect 38011 36667 38017 36701
rect 37971 36629 38017 36667
rect 37971 36595 37977 36629
rect 38011 36595 38017 36629
rect 37971 36557 38017 36595
rect 37971 36523 37977 36557
rect 38011 36523 38017 36557
rect 37971 36485 38017 36523
rect 37971 36451 37977 36485
rect 38011 36451 38017 36485
rect 37971 36413 38017 36451
rect 37971 36379 37977 36413
rect 38011 36379 38017 36413
rect 37971 36341 38017 36379
rect 37971 36307 37977 36341
rect 38011 36307 38017 36341
rect 37971 36269 38017 36307
rect 37971 36235 37977 36269
rect 38011 36235 38017 36269
rect 37971 36197 38017 36235
rect 37971 36163 37977 36197
rect 38011 36163 38017 36197
rect 37971 36147 38017 36163
rect 38429 37421 38475 37437
rect 38429 37387 38435 37421
rect 38469 37387 38475 37421
rect 38429 37349 38475 37387
rect 38429 37315 38435 37349
rect 38469 37315 38475 37349
rect 38429 37277 38475 37315
rect 38429 37243 38435 37277
rect 38469 37243 38475 37277
rect 38429 37205 38475 37243
rect 38429 37171 38435 37205
rect 38469 37171 38475 37205
rect 38429 37133 38475 37171
rect 38429 37099 38435 37133
rect 38469 37099 38475 37133
rect 38429 37061 38475 37099
rect 38429 37027 38435 37061
rect 38469 37027 38475 37061
rect 38429 36989 38475 37027
rect 38429 36955 38435 36989
rect 38469 36955 38475 36989
rect 38429 36917 38475 36955
rect 38429 36883 38435 36917
rect 38469 36883 38475 36917
rect 38429 36845 38475 36883
rect 38429 36811 38435 36845
rect 38469 36811 38475 36845
rect 38429 36773 38475 36811
rect 38429 36739 38435 36773
rect 38469 36739 38475 36773
rect 38429 36701 38475 36739
rect 38429 36667 38435 36701
rect 38469 36667 38475 36701
rect 38429 36629 38475 36667
rect 38429 36595 38435 36629
rect 38469 36595 38475 36629
rect 38429 36557 38475 36595
rect 38429 36523 38435 36557
rect 38469 36523 38475 36557
rect 38429 36485 38475 36523
rect 38429 36451 38435 36485
rect 38469 36451 38475 36485
rect 38429 36413 38475 36451
rect 38429 36379 38435 36413
rect 38469 36379 38475 36413
rect 38429 36341 38475 36379
rect 38429 36307 38435 36341
rect 38469 36307 38475 36341
rect 38429 36269 38475 36307
rect 38429 36235 38435 36269
rect 38469 36235 38475 36269
rect 38429 36197 38475 36235
rect 38429 36163 38435 36197
rect 38469 36163 38475 36197
rect 38429 36147 38475 36163
rect 38887 37421 38933 37437
rect 38887 37387 38893 37421
rect 38927 37387 38933 37421
rect 38887 37349 38933 37387
rect 38887 37315 38893 37349
rect 38927 37315 38933 37349
rect 38887 37277 38933 37315
rect 38887 37243 38893 37277
rect 38927 37243 38933 37277
rect 38887 37205 38933 37243
rect 38887 37171 38893 37205
rect 38927 37171 38933 37205
rect 38887 37133 38933 37171
rect 38887 37099 38893 37133
rect 38927 37099 38933 37133
rect 38887 37061 38933 37099
rect 38887 37027 38893 37061
rect 38927 37027 38933 37061
rect 38887 36989 38933 37027
rect 38887 36955 38893 36989
rect 38927 36955 38933 36989
rect 38887 36917 38933 36955
rect 38887 36883 38893 36917
rect 38927 36883 38933 36917
rect 38887 36845 38933 36883
rect 38887 36811 38893 36845
rect 38927 36811 38933 36845
rect 38887 36773 38933 36811
rect 38887 36739 38893 36773
rect 38927 36739 38933 36773
rect 38887 36701 38933 36739
rect 38887 36667 38893 36701
rect 38927 36667 38933 36701
rect 38887 36629 38933 36667
rect 38887 36595 38893 36629
rect 38927 36595 38933 36629
rect 38887 36557 38933 36595
rect 38887 36523 38893 36557
rect 38927 36523 38933 36557
rect 38887 36485 38933 36523
rect 38887 36451 38893 36485
rect 38927 36451 38933 36485
rect 38887 36413 38933 36451
rect 38887 36379 38893 36413
rect 38927 36379 38933 36413
rect 38887 36341 38933 36379
rect 38887 36307 38893 36341
rect 38927 36307 38933 36341
rect 38887 36269 38933 36307
rect 38887 36235 38893 36269
rect 38927 36235 38933 36269
rect 38887 36197 38933 36235
rect 38887 36163 38893 36197
rect 38927 36163 38933 36197
rect 38887 36147 38933 36163
rect 39345 37421 39391 37437
rect 39345 37387 39351 37421
rect 39385 37387 39391 37421
rect 39345 37349 39391 37387
rect 39345 37315 39351 37349
rect 39385 37315 39391 37349
rect 39345 37277 39391 37315
rect 39345 37243 39351 37277
rect 39385 37243 39391 37277
rect 39345 37205 39391 37243
rect 39345 37171 39351 37205
rect 39385 37171 39391 37205
rect 39345 37133 39391 37171
rect 39345 37099 39351 37133
rect 39385 37099 39391 37133
rect 39345 37061 39391 37099
rect 39345 37027 39351 37061
rect 39385 37027 39391 37061
rect 39345 36989 39391 37027
rect 39345 36955 39351 36989
rect 39385 36955 39391 36989
rect 39345 36917 39391 36955
rect 39345 36883 39351 36917
rect 39385 36883 39391 36917
rect 39345 36845 39391 36883
rect 39345 36811 39351 36845
rect 39385 36811 39391 36845
rect 39345 36773 39391 36811
rect 39345 36739 39351 36773
rect 39385 36739 39391 36773
rect 39345 36701 39391 36739
rect 39345 36667 39351 36701
rect 39385 36667 39391 36701
rect 39345 36629 39391 36667
rect 39345 36595 39351 36629
rect 39385 36595 39391 36629
rect 39345 36557 39391 36595
rect 39345 36523 39351 36557
rect 39385 36523 39391 36557
rect 39345 36485 39391 36523
rect 39345 36451 39351 36485
rect 39385 36451 39391 36485
rect 39345 36413 39391 36451
rect 39345 36379 39351 36413
rect 39385 36379 39391 36413
rect 39345 36341 39391 36379
rect 39345 36307 39351 36341
rect 39385 36307 39391 36341
rect 39345 36269 39391 36307
rect 39345 36235 39351 36269
rect 39385 36235 39391 36269
rect 39345 36197 39391 36235
rect 39345 36163 39351 36197
rect 39385 36163 39391 36197
rect 39345 36147 39391 36163
rect 39803 37421 39849 37437
rect 39803 37387 39809 37421
rect 39843 37387 39849 37421
rect 39803 37349 39849 37387
rect 39803 37315 39809 37349
rect 39843 37315 39849 37349
rect 39803 37277 39849 37315
rect 39803 37243 39809 37277
rect 39843 37243 39849 37277
rect 39803 37205 39849 37243
rect 39803 37171 39809 37205
rect 39843 37171 39849 37205
rect 39803 37133 39849 37171
rect 39803 37099 39809 37133
rect 39843 37099 39849 37133
rect 39803 37061 39849 37099
rect 39803 37027 39809 37061
rect 39843 37027 39849 37061
rect 39803 36989 39849 37027
rect 39803 36955 39809 36989
rect 39843 36955 39849 36989
rect 39803 36917 39849 36955
rect 39803 36883 39809 36917
rect 39843 36883 39849 36917
rect 39803 36845 39849 36883
rect 39803 36811 39809 36845
rect 39843 36811 39849 36845
rect 39803 36773 39849 36811
rect 39803 36739 39809 36773
rect 39843 36739 39849 36773
rect 39803 36701 39849 36739
rect 39803 36667 39809 36701
rect 39843 36667 39849 36701
rect 39803 36629 39849 36667
rect 39803 36595 39809 36629
rect 39843 36595 39849 36629
rect 39803 36557 39849 36595
rect 39803 36523 39809 36557
rect 39843 36523 39849 36557
rect 39803 36485 39849 36523
rect 39803 36451 39809 36485
rect 39843 36451 39849 36485
rect 39803 36413 39849 36451
rect 39803 36379 39809 36413
rect 39843 36379 39849 36413
rect 39803 36341 39849 36379
rect 39803 36307 39809 36341
rect 39843 36307 39849 36341
rect 39803 36269 39849 36307
rect 39803 36235 39809 36269
rect 39843 36235 39849 36269
rect 39803 36197 39849 36235
rect 39803 36163 39809 36197
rect 39843 36163 39849 36197
rect 39803 36147 39849 36163
rect 40261 37421 40307 37437
rect 40261 37387 40267 37421
rect 40301 37387 40307 37421
rect 40261 37349 40307 37387
rect 40261 37315 40267 37349
rect 40301 37315 40307 37349
rect 40261 37277 40307 37315
rect 41810 37356 52478 37362
rect 41810 37322 41830 37356
rect 41864 37322 41920 37356
rect 41954 37322 42010 37356
rect 42044 37322 42100 37356
rect 42134 37322 42190 37356
rect 42224 37322 42280 37356
rect 42314 37322 42370 37356
rect 42404 37322 42460 37356
rect 42494 37322 42550 37356
rect 42584 37322 42640 37356
rect 42674 37322 42730 37356
rect 42764 37322 42820 37356
rect 42854 37322 42910 37356
rect 42944 37322 43000 37356
rect 43034 37322 43170 37356
rect 43204 37322 43260 37356
rect 43294 37322 43350 37356
rect 43384 37322 43440 37356
rect 43474 37322 43530 37356
rect 43564 37322 43620 37356
rect 43654 37322 43710 37356
rect 43744 37322 43800 37356
rect 43834 37322 43890 37356
rect 43924 37322 43980 37356
rect 44014 37322 44070 37356
rect 44104 37322 44160 37356
rect 44194 37322 44250 37356
rect 44284 37322 44340 37356
rect 44374 37322 44510 37356
rect 44544 37322 44600 37356
rect 44634 37322 44690 37356
rect 44724 37322 44780 37356
rect 44814 37322 44870 37356
rect 44904 37322 44960 37356
rect 44994 37322 45050 37356
rect 45084 37322 45140 37356
rect 45174 37322 45230 37356
rect 45264 37322 45320 37356
rect 45354 37322 45410 37356
rect 45444 37322 45500 37356
rect 45534 37322 45590 37356
rect 45624 37322 45680 37356
rect 45714 37322 45850 37356
rect 45884 37322 45940 37356
rect 45974 37322 46030 37356
rect 46064 37322 46120 37356
rect 46154 37322 46210 37356
rect 46244 37322 46300 37356
rect 46334 37322 46390 37356
rect 46424 37322 46480 37356
rect 46514 37322 46570 37356
rect 46604 37322 46660 37356
rect 46694 37322 46750 37356
rect 46784 37322 46840 37356
rect 46874 37322 46930 37356
rect 46964 37322 47020 37356
rect 47054 37322 47190 37356
rect 47224 37322 47280 37356
rect 47314 37322 47370 37356
rect 47404 37322 47460 37356
rect 47494 37322 47550 37356
rect 47584 37322 47640 37356
rect 47674 37322 47730 37356
rect 47764 37322 47820 37356
rect 47854 37322 47910 37356
rect 47944 37322 48000 37356
rect 48034 37322 48090 37356
rect 48124 37322 48180 37356
rect 48214 37322 48270 37356
rect 48304 37322 48360 37356
rect 48394 37322 48530 37356
rect 48564 37322 48620 37356
rect 48654 37322 48710 37356
rect 48744 37322 48800 37356
rect 48834 37322 48890 37356
rect 48924 37322 48980 37356
rect 49014 37322 49070 37356
rect 49104 37322 49160 37356
rect 49194 37322 49250 37356
rect 49284 37322 49340 37356
rect 49374 37322 49430 37356
rect 49464 37322 49520 37356
rect 49554 37322 49610 37356
rect 49644 37322 49700 37356
rect 49734 37322 49870 37356
rect 49904 37322 49960 37356
rect 49994 37322 50050 37356
rect 50084 37322 50140 37356
rect 50174 37322 50230 37356
rect 50264 37322 50320 37356
rect 50354 37322 50410 37356
rect 50444 37322 50500 37356
rect 50534 37322 50590 37356
rect 50624 37322 50680 37356
rect 50714 37322 50770 37356
rect 50804 37322 50860 37356
rect 50894 37322 50950 37356
rect 50984 37322 51040 37356
rect 51074 37322 51210 37356
rect 51244 37322 51300 37356
rect 51334 37322 51390 37356
rect 51424 37322 51480 37356
rect 51514 37322 51570 37356
rect 51604 37322 51660 37356
rect 51694 37322 51750 37356
rect 51784 37322 51840 37356
rect 51874 37322 51930 37356
rect 51964 37322 52020 37356
rect 52054 37322 52110 37356
rect 52144 37322 52200 37356
rect 52234 37322 52290 37356
rect 52324 37322 52380 37356
rect 52414 37322 52478 37356
rect 41810 37292 52478 37322
rect 40261 37243 40267 37277
rect 40301 37243 40307 37277
rect 40261 37205 40307 37243
rect 41984 37212 42012 37292
rect 40261 37171 40267 37205
rect 40301 37171 40307 37205
rect 41974 37196 52314 37212
rect 41974 37188 41994 37196
rect 40261 37133 40307 37171
rect 41966 37136 41972 37188
rect 42028 37162 42084 37196
rect 42118 37162 42174 37196
rect 42208 37162 42264 37196
rect 42298 37162 42354 37196
rect 42388 37162 42444 37196
rect 42478 37162 42534 37196
rect 42568 37162 42624 37196
rect 42658 37162 42714 37196
rect 42748 37162 42804 37196
rect 42838 37162 42894 37196
rect 42928 37162 43334 37196
rect 43368 37162 43424 37196
rect 43458 37162 43514 37196
rect 43548 37162 43604 37196
rect 43638 37162 43694 37196
rect 43728 37162 43784 37196
rect 43818 37162 43874 37196
rect 43908 37162 43964 37196
rect 43998 37162 44054 37196
rect 44088 37162 44144 37196
rect 44178 37162 44234 37196
rect 44268 37162 44674 37196
rect 44708 37162 44764 37196
rect 44798 37162 44854 37196
rect 44888 37162 44944 37196
rect 44978 37162 45034 37196
rect 45068 37162 45124 37196
rect 45158 37162 45214 37196
rect 45248 37162 45304 37196
rect 45338 37162 45394 37196
rect 45428 37162 45484 37196
rect 45518 37162 45574 37196
rect 45608 37162 46014 37196
rect 46048 37162 46104 37196
rect 46138 37162 46194 37196
rect 46228 37162 46284 37196
rect 46318 37162 46374 37196
rect 46408 37162 46464 37196
rect 46498 37162 46554 37196
rect 46588 37162 46644 37196
rect 46678 37162 46734 37196
rect 46768 37162 46824 37196
rect 46858 37162 46914 37196
rect 46948 37162 47354 37196
rect 47388 37162 47444 37196
rect 47478 37162 47534 37196
rect 47568 37162 47624 37196
rect 47658 37162 47714 37196
rect 47748 37162 47804 37196
rect 47838 37162 47894 37196
rect 47928 37162 47984 37196
rect 48018 37162 48074 37196
rect 48108 37162 48164 37196
rect 48198 37162 48254 37196
rect 48288 37162 48694 37196
rect 48728 37162 48784 37196
rect 48818 37162 48874 37196
rect 48908 37162 48964 37196
rect 48998 37162 49054 37196
rect 49088 37162 49144 37196
rect 49178 37162 49234 37196
rect 49268 37162 49324 37196
rect 49358 37162 49414 37196
rect 49448 37162 49504 37196
rect 49538 37162 49594 37196
rect 49628 37162 50034 37196
rect 50068 37162 50124 37196
rect 50158 37162 50214 37196
rect 50248 37162 50304 37196
rect 50338 37162 50394 37196
rect 50428 37162 50484 37196
rect 50518 37162 50574 37196
rect 50608 37162 50664 37196
rect 50698 37162 50754 37196
rect 50788 37162 50844 37196
rect 50878 37162 50934 37196
rect 50968 37162 51374 37196
rect 51408 37162 51464 37196
rect 51498 37162 51554 37196
rect 51588 37162 51644 37196
rect 51678 37162 51734 37196
rect 51768 37162 51824 37196
rect 51858 37162 51914 37196
rect 51948 37162 52004 37196
rect 52038 37162 52094 37196
rect 52128 37162 52184 37196
rect 52218 37162 52274 37196
rect 52308 37162 52314 37196
rect 42024 37142 52314 37162
rect 42024 37136 42030 37142
rect 40261 37099 40267 37133
rect 40301 37099 40307 37133
rect 40261 37061 40307 37099
rect 40261 37027 40267 37061
rect 40301 37027 40307 37061
rect 40261 36989 40307 37027
rect 40261 36955 40267 36989
rect 40301 36955 40307 36989
rect 40261 36917 40307 36955
rect 40261 36883 40267 36917
rect 40301 36883 40307 36917
rect 40261 36845 40307 36883
rect 40261 36811 40267 36845
rect 40301 36811 40307 36845
rect 40261 36773 40307 36811
rect 40261 36739 40267 36773
rect 40301 36739 40307 36773
rect 40261 36701 40307 36739
rect 40261 36667 40267 36701
rect 40301 36667 40307 36701
rect 40261 36629 40307 36667
rect 40261 36595 40267 36629
rect 40301 36595 40307 36629
rect 40261 36557 40307 36595
rect 40261 36523 40267 36557
rect 40301 36523 40307 36557
rect 40261 36485 40307 36523
rect 40261 36451 40267 36485
rect 40301 36451 40307 36485
rect 40261 36413 40307 36451
rect 42148 36992 52140 37038
rect 42148 36958 42180 36992
rect 42214 36958 42280 36992
rect 42314 36958 42380 36992
rect 42414 36958 42480 36992
rect 42514 36958 42580 36992
rect 42614 36958 42680 36992
rect 42714 36958 43520 36992
rect 43554 36958 43620 36992
rect 43654 36958 43720 36992
rect 43754 36958 43820 36992
rect 43854 36958 43920 36992
rect 43954 36958 44020 36992
rect 44054 36958 44860 36992
rect 44894 36958 44960 36992
rect 44994 36958 45060 36992
rect 45094 36958 45160 36992
rect 45194 36958 45260 36992
rect 45294 36958 45360 36992
rect 45394 36958 46200 36992
rect 46234 36958 46300 36992
rect 46334 36958 46400 36992
rect 46434 36958 46500 36992
rect 46534 36958 46600 36992
rect 46634 36958 46700 36992
rect 46734 36958 47540 36992
rect 47574 36958 47640 36992
rect 47674 36958 47740 36992
rect 47774 36958 47840 36992
rect 47874 36958 47940 36992
rect 47974 36958 48040 36992
rect 48074 36958 48880 36992
rect 48914 36958 48980 36992
rect 49014 36958 49080 36992
rect 49114 36958 49180 36992
rect 49214 36958 49280 36992
rect 49314 36958 49380 36992
rect 49414 36958 50220 36992
rect 50254 36958 50320 36992
rect 50354 36958 50420 36992
rect 50454 36958 50520 36992
rect 50554 36958 50620 36992
rect 50654 36958 50720 36992
rect 50754 36958 51560 36992
rect 51594 36958 51660 36992
rect 51694 36958 51760 36992
rect 51794 36958 51860 36992
rect 51894 36958 51960 36992
rect 51994 36958 52060 36992
rect 52094 36958 52140 36992
rect 42148 36892 52140 36958
rect 42148 36858 42180 36892
rect 42214 36858 42280 36892
rect 42314 36858 42380 36892
rect 42414 36858 42480 36892
rect 42514 36858 42580 36892
rect 42614 36858 42680 36892
rect 42714 36858 43520 36892
rect 43554 36858 43620 36892
rect 43654 36858 43720 36892
rect 43754 36858 43820 36892
rect 43854 36858 43920 36892
rect 43954 36858 44020 36892
rect 44054 36858 44860 36892
rect 44894 36858 44960 36892
rect 44994 36858 45060 36892
rect 45094 36858 45160 36892
rect 45194 36858 45260 36892
rect 45294 36858 45360 36892
rect 45394 36858 46200 36892
rect 46234 36858 46300 36892
rect 46334 36858 46400 36892
rect 46434 36858 46500 36892
rect 46534 36858 46600 36892
rect 46634 36858 46700 36892
rect 46734 36858 47540 36892
rect 47574 36858 47640 36892
rect 47674 36858 47740 36892
rect 47774 36858 47840 36892
rect 47874 36858 47940 36892
rect 47974 36858 48040 36892
rect 48074 36858 48880 36892
rect 48914 36858 48980 36892
rect 49014 36858 49080 36892
rect 49114 36858 49180 36892
rect 49214 36858 49280 36892
rect 49314 36858 49380 36892
rect 49414 36858 50220 36892
rect 50254 36858 50320 36892
rect 50354 36858 50420 36892
rect 50454 36858 50520 36892
rect 50554 36858 50620 36892
rect 50654 36858 50720 36892
rect 50754 36858 51560 36892
rect 51594 36858 51660 36892
rect 51694 36858 51760 36892
rect 51794 36858 51860 36892
rect 51894 36858 51960 36892
rect 51994 36858 52060 36892
rect 52094 36858 52140 36892
rect 42148 36792 52140 36858
rect 42148 36758 42180 36792
rect 42214 36758 42280 36792
rect 42314 36758 42380 36792
rect 42414 36758 42480 36792
rect 42514 36758 42580 36792
rect 42614 36758 42680 36792
rect 42714 36758 43520 36792
rect 43554 36758 43620 36792
rect 43654 36758 43720 36792
rect 43754 36758 43820 36792
rect 43854 36758 43920 36792
rect 43954 36758 44020 36792
rect 44054 36758 44860 36792
rect 44894 36758 44960 36792
rect 44994 36758 45060 36792
rect 45094 36758 45160 36792
rect 45194 36758 45260 36792
rect 45294 36758 45360 36792
rect 45394 36758 46200 36792
rect 46234 36758 46300 36792
rect 46334 36758 46400 36792
rect 46434 36758 46500 36792
rect 46534 36758 46600 36792
rect 46634 36758 46700 36792
rect 46734 36758 47540 36792
rect 47574 36758 47640 36792
rect 47674 36758 47740 36792
rect 47774 36758 47840 36792
rect 47874 36758 47940 36792
rect 47974 36758 48040 36792
rect 48074 36758 48880 36792
rect 48914 36758 48980 36792
rect 49014 36758 49080 36792
rect 49114 36758 49180 36792
rect 49214 36758 49280 36792
rect 49314 36758 49380 36792
rect 49414 36758 50220 36792
rect 50254 36758 50320 36792
rect 50354 36758 50420 36792
rect 50454 36758 50520 36792
rect 50554 36758 50620 36792
rect 50654 36758 50720 36792
rect 50754 36758 51560 36792
rect 51594 36758 51660 36792
rect 51694 36758 51760 36792
rect 51794 36758 51860 36792
rect 51894 36758 51960 36792
rect 51994 36758 52060 36792
rect 52094 36758 52140 36792
rect 42148 36692 52140 36758
rect 42148 36658 42180 36692
rect 42214 36658 42280 36692
rect 42314 36658 42380 36692
rect 42414 36658 42480 36692
rect 42514 36658 42580 36692
rect 42614 36658 42680 36692
rect 42714 36658 43520 36692
rect 43554 36658 43620 36692
rect 43654 36658 43720 36692
rect 43754 36658 43820 36692
rect 43854 36658 43920 36692
rect 43954 36658 44020 36692
rect 44054 36658 44860 36692
rect 44894 36658 44960 36692
rect 44994 36658 45060 36692
rect 45094 36658 45160 36692
rect 45194 36658 45260 36692
rect 45294 36658 45360 36692
rect 45394 36658 46200 36692
rect 46234 36658 46300 36692
rect 46334 36658 46400 36692
rect 46434 36658 46500 36692
rect 46534 36658 46600 36692
rect 46634 36658 46700 36692
rect 46734 36658 47540 36692
rect 47574 36658 47640 36692
rect 47674 36658 47740 36692
rect 47774 36658 47840 36692
rect 47874 36658 47940 36692
rect 47974 36658 48040 36692
rect 48074 36658 48880 36692
rect 48914 36658 48980 36692
rect 49014 36658 49080 36692
rect 49114 36658 49180 36692
rect 49214 36658 49280 36692
rect 49314 36658 49380 36692
rect 49414 36658 50220 36692
rect 50254 36658 50320 36692
rect 50354 36658 50420 36692
rect 50454 36658 50520 36692
rect 50554 36658 50620 36692
rect 50654 36658 50720 36692
rect 50754 36658 51560 36692
rect 51594 36658 51660 36692
rect 51694 36658 51760 36692
rect 51794 36658 51860 36692
rect 51894 36658 51960 36692
rect 51994 36658 52060 36692
rect 52094 36658 52140 36692
rect 42148 36592 52140 36658
rect 42148 36558 42180 36592
rect 42214 36558 42280 36592
rect 42314 36558 42380 36592
rect 42414 36558 42480 36592
rect 42514 36558 42580 36592
rect 42614 36558 42680 36592
rect 42714 36558 43520 36592
rect 43554 36558 43620 36592
rect 43654 36558 43720 36592
rect 43754 36558 43820 36592
rect 43854 36558 43920 36592
rect 43954 36558 44020 36592
rect 44054 36558 44860 36592
rect 44894 36558 44960 36592
rect 44994 36558 45060 36592
rect 45094 36558 45160 36592
rect 45194 36558 45260 36592
rect 45294 36558 45360 36592
rect 45394 36558 46200 36592
rect 46234 36558 46300 36592
rect 46334 36558 46400 36592
rect 46434 36558 46500 36592
rect 46534 36558 46600 36592
rect 46634 36558 46700 36592
rect 46734 36558 47540 36592
rect 47574 36558 47640 36592
rect 47674 36558 47740 36592
rect 47774 36558 47840 36592
rect 47874 36558 47940 36592
rect 47974 36558 48040 36592
rect 48074 36558 48880 36592
rect 48914 36558 48980 36592
rect 49014 36558 49080 36592
rect 49114 36558 49180 36592
rect 49214 36558 49280 36592
rect 49314 36558 49380 36592
rect 49414 36558 50220 36592
rect 50254 36558 50320 36592
rect 50354 36558 50420 36592
rect 50454 36558 50520 36592
rect 50554 36558 50620 36592
rect 50654 36558 50720 36592
rect 50754 36558 51560 36592
rect 51594 36558 51660 36592
rect 51694 36558 51760 36592
rect 51794 36558 51860 36592
rect 51894 36558 51960 36592
rect 51994 36558 52060 36592
rect 52094 36558 52140 36592
rect 42148 36508 52140 36558
rect 42148 36456 42156 36508
rect 42208 36492 52140 36508
rect 42214 36458 42280 36492
rect 42314 36458 42380 36492
rect 42414 36458 42480 36492
rect 42514 36458 42580 36492
rect 42614 36458 42680 36492
rect 42714 36458 43520 36492
rect 43554 36458 43620 36492
rect 43654 36458 43720 36492
rect 43754 36458 43820 36492
rect 43854 36458 43920 36492
rect 43954 36458 44020 36492
rect 44054 36458 44860 36492
rect 44894 36458 44960 36492
rect 44994 36458 45060 36492
rect 45094 36458 45160 36492
rect 45194 36458 45260 36492
rect 45294 36458 45360 36492
rect 45394 36458 46200 36492
rect 46234 36458 46300 36492
rect 46334 36458 46400 36492
rect 46434 36458 46500 36492
rect 46534 36458 46600 36492
rect 46634 36458 46700 36492
rect 46734 36458 47540 36492
rect 47574 36458 47640 36492
rect 47674 36458 47740 36492
rect 47774 36458 47840 36492
rect 47874 36458 47940 36492
rect 47974 36458 48040 36492
rect 48074 36458 48880 36492
rect 48914 36458 48980 36492
rect 49014 36458 49080 36492
rect 49114 36458 49180 36492
rect 49214 36458 49280 36492
rect 49314 36458 49380 36492
rect 49414 36458 50220 36492
rect 50254 36458 50320 36492
rect 50354 36458 50420 36492
rect 50454 36458 50520 36492
rect 50554 36458 50620 36492
rect 50654 36458 50720 36492
rect 50754 36458 51560 36492
rect 51594 36458 51660 36492
rect 51694 36458 51760 36492
rect 51794 36458 51860 36492
rect 51894 36458 51960 36492
rect 51994 36458 52060 36492
rect 52094 36458 52140 36492
rect 42208 36456 52140 36458
rect 42148 36426 52140 36456
rect 40261 36379 40267 36413
rect 40301 36379 40307 36413
rect 40261 36341 40307 36379
rect 40261 36307 40267 36341
rect 40301 36307 40307 36341
rect 40261 36269 40307 36307
rect 40261 36235 40267 36269
rect 40301 36235 40307 36269
rect 40261 36197 40307 36235
rect 40261 36163 40267 36197
rect 40301 36163 40307 36197
rect 40261 36147 40307 36163
rect 37553 36057 37611 36063
rect 37553 36032 37565 36057
rect 37599 36032 37611 36057
rect 37550 35980 37556 36032
rect 37608 35980 37614 36032
rect 38562 35952 38568 35964
rect 38507 35924 38568 35952
rect 24506 35907 24938 35923
rect 38562 35912 38568 35924
rect 38620 35912 38626 35964
rect 900 35850 57536 35852
rect 900 35734 922 35850
rect 2510 35828 55926 35850
rect 2510 35809 41972 35828
rect 42024 35809 55926 35828
rect 2510 35775 12175 35809
rect 12209 35775 12375 35809
rect 12409 35775 12575 35809
rect 12609 35775 12775 35809
rect 12809 35775 12975 35809
rect 13009 35775 13175 35809
rect 13209 35775 13861 35809
rect 13895 35775 14061 35809
rect 14095 35775 14261 35809
rect 14295 35775 14461 35809
rect 14495 35775 14661 35809
rect 14695 35775 14861 35809
rect 14895 35775 15061 35809
rect 15095 35775 15261 35809
rect 15295 35775 15461 35809
rect 15495 35775 15661 35809
rect 15695 35775 15861 35809
rect 15895 35775 16605 35809
rect 16639 35775 16805 35809
rect 16839 35775 17005 35809
rect 17039 35775 17205 35809
rect 17239 35775 17405 35809
rect 17439 35775 17605 35809
rect 17639 35775 17805 35809
rect 17839 35775 18005 35809
rect 18039 35775 18205 35809
rect 18239 35775 18405 35809
rect 18439 35775 18605 35809
rect 18639 35775 19351 35809
rect 19385 35775 19551 35809
rect 19585 35775 19751 35809
rect 19785 35775 19951 35809
rect 19985 35775 20151 35809
rect 20185 35775 20351 35809
rect 20385 35775 20551 35809
rect 20585 35775 20751 35809
rect 20785 35775 20951 35809
rect 20985 35775 21151 35809
rect 21185 35775 21351 35809
rect 21385 35775 21551 35809
rect 21585 35775 21751 35809
rect 21785 35775 21951 35809
rect 21985 35775 22681 35809
rect 22715 35775 22881 35809
rect 22915 35775 23081 35809
rect 23115 35775 23281 35809
rect 23315 35775 23481 35809
rect 23515 35775 23681 35809
rect 23715 35775 23881 35809
rect 23915 35775 24081 35809
rect 24115 35775 24281 35809
rect 24315 35775 24481 35809
rect 24515 35775 24681 35809
rect 24715 35775 25601 35809
rect 25635 35775 26001 35809
rect 26035 35775 26401 35809
rect 26435 35775 26801 35809
rect 26835 35775 27201 35809
rect 27235 35775 27601 35809
rect 27635 35775 28001 35809
rect 28035 35775 28401 35809
rect 28435 35775 28801 35809
rect 28835 35775 29201 35809
rect 29235 35775 30111 35809
rect 30145 35775 30511 35809
rect 30545 35775 30911 35809
rect 30945 35775 31311 35809
rect 31345 35775 31711 35809
rect 31745 35775 32111 35809
rect 32145 35775 32511 35809
rect 32545 35775 32911 35809
rect 32945 35775 33311 35809
rect 33345 35775 33711 35809
rect 33745 35775 34111 35809
rect 34145 35775 34511 35809
rect 34545 35775 34911 35809
rect 34945 35775 35311 35809
rect 35345 35775 35711 35809
rect 35745 35775 36111 35809
rect 36145 35775 36511 35809
rect 36545 35775 36911 35809
rect 36945 35775 37655 35809
rect 37689 35775 38055 35809
rect 38089 35775 38455 35809
rect 38489 35775 38855 35809
rect 38889 35775 39255 35809
rect 39289 35775 39655 35809
rect 39689 35775 40055 35809
rect 40089 35775 41967 35809
rect 42024 35776 42167 35809
rect 42001 35775 42167 35776
rect 42201 35775 42367 35809
rect 42401 35775 42567 35809
rect 42601 35775 42767 35809
rect 42801 35775 42967 35809
rect 43001 35775 43167 35809
rect 43201 35775 43367 35809
rect 43401 35775 43567 35809
rect 43601 35775 43767 35809
rect 43801 35775 43967 35809
rect 44001 35775 44167 35809
rect 44201 35775 44367 35809
rect 44401 35775 44567 35809
rect 44601 35775 44767 35809
rect 44801 35775 44967 35809
rect 45001 35775 45167 35809
rect 45201 35775 45367 35809
rect 45401 35775 45567 35809
rect 45601 35775 45767 35809
rect 45801 35775 45967 35809
rect 46001 35775 46167 35809
rect 46201 35775 46367 35809
rect 46401 35775 46567 35809
rect 46601 35775 46767 35809
rect 46801 35775 46967 35809
rect 47001 35775 47167 35809
rect 47201 35775 47367 35809
rect 47401 35775 47567 35809
rect 47601 35775 47767 35809
rect 47801 35775 47967 35809
rect 48001 35775 48167 35809
rect 48201 35775 48367 35809
rect 48401 35775 48567 35809
rect 48601 35775 48767 35809
rect 48801 35775 48967 35809
rect 49001 35775 49167 35809
rect 49201 35775 49367 35809
rect 49401 35775 49567 35809
rect 49601 35775 49767 35809
rect 49801 35775 49967 35809
rect 50001 35775 50167 35809
rect 50201 35775 50367 35809
rect 50401 35775 50567 35809
rect 50601 35775 50767 35809
rect 50801 35775 50967 35809
rect 51001 35775 51167 35809
rect 51201 35775 51367 35809
rect 51401 35775 51567 35809
rect 51601 35775 51767 35809
rect 51801 35775 51967 35809
rect 52001 35775 52167 35809
rect 52201 35775 52367 35809
rect 52401 35775 55926 35809
rect 2510 35734 55926 35775
rect 57514 35734 57536 35850
rect 900 35732 57536 35734
rect 3348 33970 55088 33972
rect 3348 33854 3370 33970
rect 4958 33929 53478 33970
rect 4958 33895 19447 33929
rect 19481 33895 19647 33929
rect 19681 33895 19847 33929
rect 19881 33895 20047 33929
rect 20081 33895 20247 33929
rect 20281 33895 20447 33929
rect 20481 33895 20647 33929
rect 20681 33895 20847 33929
rect 20881 33895 21047 33929
rect 21081 33895 21247 33929
rect 21281 33895 21447 33929
rect 21481 33895 22193 33929
rect 22227 33895 22393 33929
rect 22427 33895 22593 33929
rect 22627 33895 22793 33929
rect 22827 33895 22993 33929
rect 23027 33895 23193 33929
rect 23227 33895 23393 33929
rect 23427 33895 23593 33929
rect 23627 33895 23793 33929
rect 23827 33895 23993 33929
rect 24027 33895 24193 33929
rect 24227 33895 24393 33929
rect 24427 33895 24593 33929
rect 24627 33895 24793 33929
rect 24827 33895 26387 33929
rect 26421 33895 26787 33929
rect 26821 33895 27187 33929
rect 27221 33895 27587 33929
rect 27621 33895 27987 33929
rect 28021 33895 28387 33929
rect 28421 33895 28787 33929
rect 28821 33895 29187 33929
rect 29221 33895 29587 33929
rect 29621 33895 29987 33929
rect 30021 33895 30387 33929
rect 30421 33895 30787 33929
rect 30821 33895 31187 33929
rect 31221 33895 31587 33929
rect 31621 33895 31987 33929
rect 32021 33895 32387 33929
rect 32421 33895 32787 33929
rect 32821 33895 33187 33929
rect 33221 33924 33835 33929
rect 33221 33895 33416 33924
rect 4958 33872 33416 33895
rect 33468 33895 33835 33924
rect 33869 33895 34235 33929
rect 34269 33895 34635 33929
rect 34669 33895 35035 33929
rect 35069 33895 35435 33929
rect 35469 33895 35835 33929
rect 35869 33895 36235 33929
rect 36269 33895 36635 33929
rect 36669 33895 37035 33929
rect 37069 33895 37435 33929
rect 37469 33895 37835 33929
rect 37869 33895 38235 33929
rect 38269 33895 38635 33929
rect 38669 33895 39035 33929
rect 39069 33895 39435 33929
rect 39469 33895 39835 33929
rect 39869 33895 40235 33929
rect 40269 33895 40635 33929
rect 40669 33895 41967 33929
rect 42001 33895 42167 33929
rect 42201 33895 42367 33929
rect 42401 33895 42567 33929
rect 42601 33895 42767 33929
rect 42801 33895 42967 33929
rect 43001 33895 43167 33929
rect 43201 33895 43367 33929
rect 43401 33895 43567 33929
rect 43601 33895 43767 33929
rect 43801 33895 43967 33929
rect 44001 33895 44167 33929
rect 44201 33895 44367 33929
rect 44401 33895 44567 33929
rect 44601 33895 44767 33929
rect 44801 33895 44967 33929
rect 45001 33895 45167 33929
rect 45201 33895 45367 33929
rect 45401 33895 45567 33929
rect 45601 33895 45767 33929
rect 45801 33895 45967 33929
rect 46001 33895 46167 33929
rect 46201 33895 46367 33929
rect 46401 33895 46567 33929
rect 46601 33895 46767 33929
rect 46801 33895 46967 33929
rect 47001 33895 47167 33929
rect 47201 33895 47367 33929
rect 47401 33895 47567 33929
rect 47601 33895 47767 33929
rect 47801 33895 47967 33929
rect 48001 33895 48167 33929
rect 48201 33895 48367 33929
rect 48401 33895 48567 33929
rect 48601 33895 48767 33929
rect 48801 33895 48967 33929
rect 49001 33895 49167 33929
rect 49201 33895 49367 33929
rect 49401 33895 49567 33929
rect 49601 33895 49767 33929
rect 49801 33895 49967 33929
rect 50001 33895 50167 33929
rect 50201 33895 50367 33929
rect 50401 33895 50567 33929
rect 50601 33895 50767 33929
rect 50801 33895 50967 33929
rect 51001 33895 51167 33929
rect 51201 33895 51367 33929
rect 51401 33895 51567 33929
rect 51601 33895 51767 33929
rect 51801 33895 51967 33929
rect 52001 33895 52167 33929
rect 52201 33895 52367 33929
rect 52401 33895 53478 33929
rect 33468 33872 53478 33895
rect 4958 33854 53478 33872
rect 55066 33854 55088 33970
rect 3348 33852 55088 33854
rect 48682 33736 48688 33788
rect 48740 33736 48746 33788
rect 48700 33708 48728 33736
rect 48700 33680 58466 33708
rect 19275 33661 19685 33673
rect 19275 33123 19283 33661
rect 19677 33123 19685 33661
rect 19275 33111 19685 33123
rect 21283 33661 21693 33673
rect 21283 33123 21290 33661
rect 21684 33123 21693 33661
rect 21283 33111 21693 33123
rect 22020 33661 22430 33673
rect 22020 33123 22028 33661
rect 22422 33164 22430 33661
rect 24602 33661 25012 33673
rect 24486 33164 24492 33176
rect 22422 33136 24492 33164
rect 22422 33123 22430 33136
rect 24486 33124 24492 33136
rect 24544 33124 24550 33176
rect 22020 33111 22430 33123
rect 24602 33123 24609 33661
rect 25003 33123 25012 33661
rect 41810 33596 52478 33602
rect 41810 33562 41830 33596
rect 41864 33584 41920 33596
rect 41864 33562 41880 33584
rect 41954 33562 42010 33596
rect 42044 33562 42100 33596
rect 42134 33562 42190 33596
rect 42224 33562 42280 33596
rect 42314 33562 42370 33596
rect 42404 33562 42460 33596
rect 42494 33562 42550 33596
rect 42584 33562 42640 33596
rect 42674 33562 42730 33596
rect 42764 33562 42820 33596
rect 42854 33562 42910 33596
rect 42944 33562 43000 33596
rect 43034 33562 43170 33596
rect 43204 33562 43260 33596
rect 43294 33562 43350 33596
rect 43384 33562 43440 33596
rect 43474 33562 43530 33596
rect 43564 33562 43620 33596
rect 43654 33562 43710 33596
rect 43744 33562 43800 33596
rect 43834 33562 43890 33596
rect 43924 33562 43980 33596
rect 44014 33562 44070 33596
rect 44104 33562 44160 33596
rect 44194 33562 44250 33596
rect 44284 33562 44340 33596
rect 44374 33562 44510 33596
rect 44544 33562 44600 33596
rect 44634 33562 44690 33596
rect 44724 33562 44780 33596
rect 44814 33562 44870 33596
rect 44904 33562 44960 33596
rect 44994 33562 45050 33596
rect 45084 33562 45140 33596
rect 45174 33562 45230 33596
rect 45264 33562 45320 33596
rect 45354 33562 45410 33596
rect 45444 33562 45500 33596
rect 45534 33562 45590 33596
rect 45624 33562 45680 33596
rect 45714 33562 45850 33596
rect 45884 33562 45940 33596
rect 45974 33562 46030 33596
rect 46064 33562 46120 33596
rect 46154 33562 46210 33596
rect 46244 33562 46300 33596
rect 46334 33562 46390 33596
rect 46424 33562 46480 33596
rect 46514 33562 46570 33596
rect 46604 33562 46660 33596
rect 46694 33562 46750 33596
rect 46784 33562 46840 33596
rect 46874 33562 46930 33596
rect 46964 33562 47020 33596
rect 47054 33562 47190 33596
rect 47224 33562 47280 33596
rect 47314 33562 47370 33596
rect 47404 33562 47460 33596
rect 47494 33562 47550 33596
rect 47584 33562 47640 33596
rect 47674 33562 47730 33596
rect 47764 33562 47820 33596
rect 47854 33562 47910 33596
rect 47944 33562 48000 33596
rect 48034 33562 48090 33596
rect 48124 33562 48180 33596
rect 48214 33562 48270 33596
rect 48304 33562 48360 33596
rect 48394 33562 48530 33596
rect 48564 33562 48620 33596
rect 48654 33562 48710 33596
rect 48744 33562 48800 33596
rect 48834 33562 48890 33596
rect 48924 33562 48980 33596
rect 49014 33562 49070 33596
rect 49104 33562 49160 33596
rect 49194 33562 49250 33596
rect 49284 33562 49340 33596
rect 49374 33562 49430 33596
rect 49464 33562 49520 33596
rect 49554 33562 49610 33596
rect 49644 33562 49700 33596
rect 49734 33562 49870 33596
rect 49904 33562 49960 33596
rect 49994 33562 50050 33596
rect 50084 33562 50140 33596
rect 50174 33562 50230 33596
rect 50264 33562 50320 33596
rect 50354 33562 50410 33596
rect 50444 33562 50500 33596
rect 50534 33562 50590 33596
rect 50624 33562 50680 33596
rect 50714 33562 50770 33596
rect 50804 33562 50860 33596
rect 50894 33562 50950 33596
rect 50984 33562 51040 33596
rect 51074 33562 51210 33596
rect 51244 33562 51300 33596
rect 51334 33562 51390 33596
rect 51424 33562 51480 33596
rect 51514 33562 51570 33596
rect 51604 33562 51660 33596
rect 51694 33562 51750 33596
rect 51784 33562 51840 33596
rect 51874 33562 51930 33596
rect 51964 33562 52020 33596
rect 52054 33562 52110 33596
rect 52144 33562 52200 33596
rect 52234 33562 52290 33596
rect 52324 33562 52380 33596
rect 52414 33562 52478 33596
rect 41810 33532 41880 33562
rect 41932 33532 52478 33562
rect 42720 33452 42748 33532
rect 41974 33436 52314 33452
rect 58438 33436 58466 33680
rect 41974 33402 41994 33436
rect 42028 33402 42084 33436
rect 42118 33402 42174 33436
rect 42208 33402 42264 33436
rect 42298 33402 42354 33436
rect 42388 33402 42444 33436
rect 42478 33402 42534 33436
rect 42568 33402 42624 33436
rect 42658 33402 42714 33436
rect 42748 33402 42804 33436
rect 42838 33402 42894 33436
rect 42928 33402 43334 33436
rect 43368 33402 43424 33436
rect 43458 33402 43514 33436
rect 43548 33402 43604 33436
rect 43638 33402 43694 33436
rect 43728 33402 43784 33436
rect 43818 33402 43874 33436
rect 43908 33402 43964 33436
rect 43998 33402 44054 33436
rect 44088 33402 44144 33436
rect 44178 33402 44234 33436
rect 44268 33402 44674 33436
rect 44708 33402 44764 33436
rect 44798 33402 44854 33436
rect 44888 33402 44944 33436
rect 44978 33402 45034 33436
rect 45068 33402 45124 33436
rect 45158 33402 45214 33436
rect 45248 33402 45304 33436
rect 45338 33402 45394 33436
rect 45428 33402 45484 33436
rect 45518 33402 45574 33436
rect 45608 33402 46014 33436
rect 46048 33402 46104 33436
rect 46138 33402 46194 33436
rect 46228 33402 46284 33436
rect 46318 33402 46374 33436
rect 46408 33402 46464 33436
rect 46498 33402 46554 33436
rect 46588 33402 46644 33436
rect 46678 33402 46734 33436
rect 46768 33402 46824 33436
rect 46858 33402 46914 33436
rect 46948 33402 47354 33436
rect 47388 33402 47444 33436
rect 47478 33402 47534 33436
rect 47568 33402 47624 33436
rect 47658 33402 47714 33436
rect 47748 33402 47804 33436
rect 47838 33402 47894 33436
rect 47928 33402 47984 33436
rect 48018 33402 48074 33436
rect 48108 33402 48164 33436
rect 48198 33402 48254 33436
rect 48288 33402 48694 33436
rect 48728 33402 48784 33436
rect 48818 33402 48874 33436
rect 48908 33402 48964 33436
rect 48998 33402 49054 33436
rect 49088 33402 49144 33436
rect 49178 33402 49234 33436
rect 49268 33402 49324 33436
rect 49358 33402 49414 33436
rect 49448 33402 49504 33436
rect 49538 33402 49594 33436
rect 49628 33402 50034 33436
rect 50068 33402 50124 33436
rect 50158 33402 50214 33436
rect 50248 33402 50304 33436
rect 50338 33402 50394 33436
rect 50428 33402 50484 33436
rect 50518 33402 50574 33436
rect 50608 33402 50664 33436
rect 50698 33402 50754 33436
rect 50788 33402 50844 33436
rect 50878 33402 50934 33436
rect 50968 33402 51374 33436
rect 51408 33402 51464 33436
rect 51498 33402 51554 33436
rect 51588 33402 51644 33436
rect 51678 33402 51734 33436
rect 51768 33402 51824 33436
rect 51858 33402 51914 33436
rect 51948 33402 52004 33436
rect 52038 33402 52094 33436
rect 52128 33402 52184 33436
rect 52218 33402 52274 33436
rect 52308 33402 52314 33436
rect 58393 33408 58512 33436
rect 41974 33382 52314 33402
rect 24602 33111 25012 33123
rect 42148 33244 52140 33278
rect 42148 33192 42156 33244
rect 42208 33232 52140 33244
rect 42214 33198 42280 33232
rect 42314 33198 42380 33232
rect 42414 33198 42480 33232
rect 42514 33198 42580 33232
rect 42614 33198 42680 33232
rect 42714 33198 43520 33232
rect 43554 33198 43620 33232
rect 43654 33198 43720 33232
rect 43754 33198 43820 33232
rect 43854 33198 43920 33232
rect 43954 33198 44020 33232
rect 44054 33198 44860 33232
rect 44894 33198 44960 33232
rect 44994 33198 45060 33232
rect 45094 33198 45160 33232
rect 45194 33198 45260 33232
rect 45294 33198 45360 33232
rect 45394 33198 46200 33232
rect 46234 33198 46300 33232
rect 46334 33198 46400 33232
rect 46434 33198 46500 33232
rect 46534 33198 46600 33232
rect 46634 33198 46700 33232
rect 46734 33198 47540 33232
rect 47574 33198 47640 33232
rect 47674 33198 47740 33232
rect 47774 33198 47840 33232
rect 47874 33198 47940 33232
rect 47974 33198 48040 33232
rect 48074 33198 48880 33232
rect 48914 33198 48980 33232
rect 49014 33198 49080 33232
rect 49114 33198 49180 33232
rect 49214 33198 49280 33232
rect 49314 33198 49380 33232
rect 49414 33198 50220 33232
rect 50254 33198 50320 33232
rect 50354 33198 50420 33232
rect 50454 33198 50520 33232
rect 50554 33198 50620 33232
rect 50654 33198 50720 33232
rect 50754 33198 51560 33232
rect 51594 33198 51660 33232
rect 51694 33198 51760 33232
rect 51794 33198 51860 33232
rect 51894 33198 51960 33232
rect 51994 33198 52060 33232
rect 52094 33198 52140 33232
rect 42208 33192 52140 33198
rect 42148 33132 52140 33192
rect 19275 32701 19685 32713
rect 16574 32648 16580 32700
rect 16632 32688 16638 32700
rect 19275 32688 19283 32701
rect 16632 32660 19283 32688
rect 16632 32648 16638 32660
rect 19275 32163 19283 32660
rect 19677 32163 19685 32701
rect 19275 32151 19685 32163
rect 21272 32701 21704 33111
rect 21272 32163 21290 32701
rect 21684 32163 21704 32701
rect 21272 32147 21704 32163
rect 22020 32701 22430 32713
rect 22020 32163 22028 32701
rect 22422 32163 22430 32701
rect 22020 32151 22430 32163
rect 24591 32701 25023 33111
rect 24591 32163 24609 32701
rect 25003 32163 25023 32701
rect 42148 33098 42180 33132
rect 42214 33098 42280 33132
rect 42314 33098 42380 33132
rect 42414 33098 42480 33132
rect 42514 33098 42580 33132
rect 42614 33098 42680 33132
rect 42714 33098 43520 33132
rect 43554 33098 43620 33132
rect 43654 33098 43720 33132
rect 43754 33098 43820 33132
rect 43854 33098 43920 33132
rect 43954 33098 44020 33132
rect 44054 33098 44860 33132
rect 44894 33098 44960 33132
rect 44994 33098 45060 33132
rect 45094 33098 45160 33132
rect 45194 33098 45260 33132
rect 45294 33098 45360 33132
rect 45394 33098 46200 33132
rect 46234 33098 46300 33132
rect 46334 33098 46400 33132
rect 46434 33098 46500 33132
rect 46534 33098 46600 33132
rect 46634 33098 46700 33132
rect 46734 33098 47540 33132
rect 47574 33098 47640 33132
rect 47674 33098 47740 33132
rect 47774 33098 47840 33132
rect 47874 33098 47940 33132
rect 47974 33098 48040 33132
rect 48074 33098 48880 33132
rect 48914 33098 48980 33132
rect 49014 33098 49080 33132
rect 49114 33098 49180 33132
rect 49214 33098 49280 33132
rect 49314 33098 49380 33132
rect 49414 33098 50220 33132
rect 50254 33098 50320 33132
rect 50354 33098 50420 33132
rect 50454 33098 50520 33132
rect 50554 33098 50620 33132
rect 50654 33098 50720 33132
rect 50754 33098 51560 33132
rect 51594 33098 51660 33132
rect 51694 33098 51760 33132
rect 51794 33098 51860 33132
rect 51894 33098 51960 33132
rect 51994 33098 52060 33132
rect 52094 33098 52140 33132
rect 42148 33032 52140 33098
rect 42148 32998 42180 33032
rect 42214 32998 42280 33032
rect 42314 32998 42380 33032
rect 42414 32998 42480 33032
rect 42514 32998 42580 33032
rect 42614 32998 42680 33032
rect 42714 32998 43520 33032
rect 43554 32998 43620 33032
rect 43654 32998 43720 33032
rect 43754 32998 43820 33032
rect 43854 32998 43920 33032
rect 43954 32998 44020 33032
rect 44054 32998 44860 33032
rect 44894 32998 44960 33032
rect 44994 32998 45060 33032
rect 45094 32998 45160 33032
rect 45194 32998 45260 33032
rect 45294 32998 45360 33032
rect 45394 32998 46200 33032
rect 46234 32998 46300 33032
rect 46334 32998 46400 33032
rect 46434 32998 46500 33032
rect 46534 32998 46600 33032
rect 46634 32998 46700 33032
rect 46734 32998 47540 33032
rect 47574 32998 47640 33032
rect 47674 32998 47740 33032
rect 47774 32998 47840 33032
rect 47874 32998 47940 33032
rect 47974 32998 48040 33032
rect 48074 32998 48880 33032
rect 48914 32998 48980 33032
rect 49014 32998 49080 33032
rect 49114 32998 49180 33032
rect 49214 32998 49280 33032
rect 49314 32998 49380 33032
rect 49414 32998 50220 33032
rect 50254 32998 50320 33032
rect 50354 32998 50420 33032
rect 50454 32998 50520 33032
rect 50554 32998 50620 33032
rect 50654 32998 50720 33032
rect 50754 32998 51560 33032
rect 51594 32998 51660 33032
rect 51694 32998 51760 33032
rect 51794 32998 51860 33032
rect 51894 32998 51960 33032
rect 51994 32998 52060 33032
rect 52094 32998 52140 33032
rect 42148 32932 52140 32998
rect 42148 32898 42180 32932
rect 42214 32898 42280 32932
rect 42314 32898 42380 32932
rect 42414 32898 42480 32932
rect 42514 32898 42580 32932
rect 42614 32898 42680 32932
rect 42714 32898 43520 32932
rect 43554 32898 43620 32932
rect 43654 32898 43720 32932
rect 43754 32898 43820 32932
rect 43854 32898 43920 32932
rect 43954 32898 44020 32932
rect 44054 32898 44860 32932
rect 44894 32898 44960 32932
rect 44994 32898 45060 32932
rect 45094 32898 45160 32932
rect 45194 32898 45260 32932
rect 45294 32898 45360 32932
rect 45394 32898 46200 32932
rect 46234 32898 46300 32932
rect 46334 32898 46400 32932
rect 46434 32898 46500 32932
rect 46534 32898 46600 32932
rect 46634 32898 46700 32932
rect 46734 32898 47540 32932
rect 47574 32898 47640 32932
rect 47674 32898 47740 32932
rect 47774 32898 47840 32932
rect 47874 32898 47940 32932
rect 47974 32898 48040 32932
rect 48074 32898 48880 32932
rect 48914 32898 48980 32932
rect 49014 32898 49080 32932
rect 49114 32898 49180 32932
rect 49214 32898 49280 32932
rect 49314 32898 49380 32932
rect 49414 32898 50220 32932
rect 50254 32898 50320 32932
rect 50354 32898 50420 32932
rect 50454 32898 50520 32932
rect 50554 32898 50620 32932
rect 50654 32898 50720 32932
rect 50754 32898 51560 32932
rect 51594 32898 51660 32932
rect 51694 32898 51760 32932
rect 51794 32898 51860 32932
rect 51894 32898 51960 32932
rect 51994 32898 52060 32932
rect 52094 32898 52140 32932
rect 42148 32832 52140 32898
rect 42148 32798 42180 32832
rect 42214 32798 42280 32832
rect 42314 32798 42380 32832
rect 42414 32798 42480 32832
rect 42514 32798 42580 32832
rect 42614 32798 42680 32832
rect 42714 32798 43520 32832
rect 43554 32798 43620 32832
rect 43654 32798 43720 32832
rect 43754 32798 43820 32832
rect 43854 32798 43920 32832
rect 43954 32798 44020 32832
rect 44054 32798 44860 32832
rect 44894 32798 44960 32832
rect 44994 32798 45060 32832
rect 45094 32798 45160 32832
rect 45194 32798 45260 32832
rect 45294 32798 45360 32832
rect 45394 32798 46200 32832
rect 46234 32798 46300 32832
rect 46334 32798 46400 32832
rect 46434 32798 46500 32832
rect 46534 32798 46600 32832
rect 46634 32798 46700 32832
rect 46734 32798 47540 32832
rect 47574 32798 47640 32832
rect 47674 32798 47740 32832
rect 47774 32798 47840 32832
rect 47874 32798 47940 32832
rect 47974 32798 48040 32832
rect 48074 32798 48880 32832
rect 48914 32798 48980 32832
rect 49014 32798 49080 32832
rect 49114 32798 49180 32832
rect 49214 32798 49280 32832
rect 49314 32798 49380 32832
rect 49414 32798 50220 32832
rect 50254 32798 50320 32832
rect 50354 32798 50420 32832
rect 50454 32798 50520 32832
rect 50554 32798 50620 32832
rect 50654 32798 50720 32832
rect 50754 32798 51560 32832
rect 51594 32798 51660 32832
rect 51694 32798 51760 32832
rect 51794 32798 51860 32832
rect 51894 32798 51960 32832
rect 51994 32798 52060 32832
rect 52094 32798 52140 32832
rect 42148 32732 52140 32798
rect 42148 32698 42180 32732
rect 42214 32700 42280 32732
rect 42214 32698 42248 32700
rect 42314 32698 42380 32732
rect 42414 32698 42480 32732
rect 42514 32698 42580 32732
rect 42614 32698 42680 32732
rect 42714 32698 43520 32732
rect 43554 32698 43620 32732
rect 43654 32698 43720 32732
rect 43754 32698 43820 32732
rect 43854 32698 43920 32732
rect 43954 32698 44020 32732
rect 44054 32698 44860 32732
rect 44894 32698 44960 32732
rect 44994 32698 45060 32732
rect 45094 32698 45160 32732
rect 45194 32698 45260 32732
rect 45294 32698 45360 32732
rect 45394 32698 46200 32732
rect 46234 32698 46300 32732
rect 46334 32698 46400 32732
rect 46434 32698 46500 32732
rect 46534 32698 46600 32732
rect 46634 32698 46700 32732
rect 46734 32698 47540 32732
rect 47574 32698 47640 32732
rect 47674 32698 47740 32732
rect 47774 32698 47840 32732
rect 47874 32698 47940 32732
rect 47974 32698 48040 32732
rect 48074 32698 48880 32732
rect 48914 32698 48980 32732
rect 49014 32698 49080 32732
rect 49114 32698 49180 32732
rect 49214 32698 49280 32732
rect 49314 32698 49380 32732
rect 49414 32698 50220 32732
rect 50254 32698 50320 32732
rect 50354 32698 50420 32732
rect 50454 32698 50520 32732
rect 50554 32698 50620 32732
rect 50654 32698 50720 32732
rect 50754 32698 51560 32732
rect 51594 32698 51660 32732
rect 51694 32698 51760 32732
rect 51794 32698 51860 32732
rect 51894 32698 51960 32732
rect 51994 32698 52060 32732
rect 52094 32698 52140 32732
rect 42148 32666 42248 32698
rect 42242 32648 42248 32666
rect 42300 32666 52140 32698
rect 42300 32648 42306 32666
rect 22388 32092 22416 32151
rect 24591 32147 25023 32163
rect 900 32090 57536 32092
rect 900 31974 922 32090
rect 2510 32049 55926 32090
rect 2510 32015 19447 32049
rect 19481 32015 19647 32049
rect 19681 32015 19847 32049
rect 19881 32015 20047 32049
rect 20081 32015 20247 32049
rect 20281 32015 20447 32049
rect 20481 32015 20647 32049
rect 20681 32015 20847 32049
rect 20881 32015 21047 32049
rect 21081 32015 21247 32049
rect 21281 32015 21447 32049
rect 21481 32015 22193 32049
rect 22227 32015 22393 32049
rect 22427 32015 22593 32049
rect 22627 32015 22793 32049
rect 22827 32015 22993 32049
rect 23027 32015 23193 32049
rect 23227 32015 23393 32049
rect 23427 32015 23593 32049
rect 23627 32015 23793 32049
rect 23827 32015 23993 32049
rect 24027 32015 24193 32049
rect 24227 32015 24393 32049
rect 24427 32015 24593 32049
rect 24627 32015 24793 32049
rect 24827 32015 26387 32049
rect 26421 32015 26787 32049
rect 26821 32015 27187 32049
rect 27221 32015 27587 32049
rect 27621 32015 27987 32049
rect 28021 32015 28387 32049
rect 28421 32015 28787 32049
rect 28821 32015 29187 32049
rect 29221 32015 29587 32049
rect 29621 32015 29987 32049
rect 30021 32015 30387 32049
rect 30421 32015 30787 32049
rect 30821 32015 31187 32049
rect 31221 32015 31587 32049
rect 31621 32015 31987 32049
rect 32021 32015 32387 32049
rect 32421 32015 32787 32049
rect 32821 32015 33187 32049
rect 33221 32015 33835 32049
rect 33869 32015 34235 32049
rect 34269 32015 34635 32049
rect 34669 32015 35035 32049
rect 35069 32015 35435 32049
rect 35469 32015 35835 32049
rect 35869 32015 36235 32049
rect 36269 32015 36635 32049
rect 36669 32015 37035 32049
rect 37069 32015 37435 32049
rect 37469 32015 37835 32049
rect 37869 32015 38235 32049
rect 38269 32015 38635 32049
rect 38669 32015 39035 32049
rect 39069 32015 39435 32049
rect 39469 32015 39835 32049
rect 39869 32015 40235 32049
rect 40269 32015 40635 32049
rect 40669 32015 41967 32049
rect 42001 32015 42167 32049
rect 42201 32015 42367 32049
rect 42401 32015 42567 32049
rect 42601 32015 42767 32049
rect 42801 32015 42967 32049
rect 43001 32015 43167 32049
rect 43201 32015 43367 32049
rect 43401 32015 43567 32049
rect 43601 32015 43767 32049
rect 43801 32015 43967 32049
rect 44001 32015 44167 32049
rect 44201 32015 44367 32049
rect 44401 32015 44567 32049
rect 44601 32015 44767 32049
rect 44801 32015 44967 32049
rect 45001 32015 45167 32049
rect 45201 32015 45367 32049
rect 45401 32015 45567 32049
rect 45601 32015 45767 32049
rect 45801 32015 45967 32049
rect 46001 32015 46167 32049
rect 46201 32015 46367 32049
rect 46401 32015 46567 32049
rect 46601 32015 46767 32049
rect 46801 32015 46967 32049
rect 47001 32015 47167 32049
rect 47201 32015 47367 32049
rect 47401 32015 47567 32049
rect 47601 32015 47767 32049
rect 47801 32015 47967 32049
rect 48001 32015 48167 32049
rect 48201 32015 48367 32049
rect 48401 32015 48567 32049
rect 48601 32015 48767 32049
rect 48801 32015 48967 32049
rect 49001 32015 49167 32049
rect 49201 32015 49367 32049
rect 49401 32015 49567 32049
rect 49601 32015 49767 32049
rect 49801 32015 49967 32049
rect 50001 32015 50167 32049
rect 50201 32015 50367 32049
rect 50401 32015 50567 32049
rect 50601 32015 50767 32049
rect 50801 32015 50967 32049
rect 51001 32015 51167 32049
rect 51201 32015 51367 32049
rect 51401 32015 51567 32049
rect 51601 32015 51767 32049
rect 51801 32015 51967 32049
rect 52001 32015 52167 32049
rect 52201 32015 52367 32049
rect 52401 32015 55926 32049
rect 2510 31974 55926 32015
rect 57514 31974 57536 32090
rect 900 31972 57536 31974
rect 3348 30210 55088 30212
rect 3348 30094 3370 30210
rect 4958 30184 53478 30210
rect 4958 30169 33416 30184
rect 4958 30135 16703 30169
rect 16737 30135 16903 30169
rect 16937 30135 17103 30169
rect 17137 30135 17303 30169
rect 17337 30135 17503 30169
rect 17537 30135 17703 30169
rect 17737 30135 17903 30169
rect 17937 30135 18103 30169
rect 18137 30135 18303 30169
rect 18337 30135 18503 30169
rect 18537 30135 18703 30169
rect 18737 30135 19447 30169
rect 19481 30135 19647 30169
rect 19681 30135 19847 30169
rect 19881 30135 20047 30169
rect 20081 30135 20247 30169
rect 20281 30135 20447 30169
rect 20481 30135 20647 30169
rect 20681 30135 20847 30169
rect 20881 30135 21047 30169
rect 21081 30135 21247 30169
rect 21281 30135 21447 30169
rect 21481 30135 22191 30169
rect 22225 30135 22391 30169
rect 22425 30135 22591 30169
rect 22625 30135 22791 30169
rect 22825 30135 22991 30169
rect 23025 30135 23191 30169
rect 23225 30135 23391 30169
rect 23425 30135 23591 30169
rect 23625 30135 23791 30169
rect 23825 30135 23991 30169
rect 24025 30135 24191 30169
rect 24225 30135 27385 30169
rect 27419 30135 27585 30169
rect 27619 30135 27785 30169
rect 27819 30135 27985 30169
rect 28019 30135 28185 30169
rect 28219 30135 28385 30169
rect 28419 30135 28585 30169
rect 28619 30135 28785 30169
rect 28819 30135 28985 30169
rect 29019 30135 29185 30169
rect 29219 30135 29385 30169
rect 29419 30135 30111 30169
rect 30145 30135 30511 30169
rect 30545 30135 30911 30169
rect 30945 30135 31311 30169
rect 31345 30135 31711 30169
rect 31745 30135 32111 30169
rect 32145 30135 32511 30169
rect 32545 30135 32911 30169
rect 32945 30135 33311 30169
rect 33345 30135 33416 30169
rect 4958 30132 33416 30135
rect 33468 30169 53478 30184
rect 33468 30135 33711 30169
rect 33745 30135 34111 30169
rect 34145 30135 34511 30169
rect 34545 30135 34911 30169
rect 34945 30135 35311 30169
rect 35345 30135 35711 30169
rect 35745 30135 36111 30169
rect 36145 30135 36511 30169
rect 36545 30135 36911 30169
rect 36945 30135 37655 30169
rect 37689 30135 38055 30169
rect 38089 30135 38455 30169
rect 38489 30135 38855 30169
rect 38889 30135 39255 30169
rect 39289 30135 39655 30169
rect 39689 30135 40055 30169
rect 40089 30135 41967 30169
rect 42001 30135 42167 30169
rect 42201 30135 42367 30169
rect 42401 30135 42567 30169
rect 42601 30135 42767 30169
rect 42801 30135 42967 30169
rect 43001 30135 43167 30169
rect 43201 30135 43367 30169
rect 43401 30135 43567 30169
rect 43601 30135 43767 30169
rect 43801 30135 43967 30169
rect 44001 30135 44167 30169
rect 44201 30135 44367 30169
rect 44401 30135 44567 30169
rect 44601 30135 44767 30169
rect 44801 30135 44967 30169
rect 45001 30135 45167 30169
rect 45201 30135 45367 30169
rect 45401 30135 45567 30169
rect 45601 30135 45767 30169
rect 45801 30135 45967 30169
rect 46001 30135 46167 30169
rect 46201 30135 46367 30169
rect 46401 30135 46567 30169
rect 46601 30135 46767 30169
rect 46801 30135 46967 30169
rect 47001 30135 47167 30169
rect 47201 30135 47367 30169
rect 47401 30135 47567 30169
rect 47601 30135 47767 30169
rect 47801 30135 47967 30169
rect 48001 30135 48167 30169
rect 48201 30135 48367 30169
rect 48401 30135 48567 30169
rect 48601 30135 48767 30169
rect 48801 30135 48967 30169
rect 49001 30135 49167 30169
rect 49201 30135 49367 30169
rect 49401 30135 49567 30169
rect 49601 30135 49767 30169
rect 49801 30135 49967 30169
rect 50001 30135 50167 30169
rect 50201 30135 50367 30169
rect 50401 30135 50567 30169
rect 50601 30135 50767 30169
rect 50801 30135 50967 30169
rect 51001 30135 51167 30169
rect 51201 30135 51367 30169
rect 51401 30135 51567 30169
rect 51601 30135 51767 30169
rect 51801 30135 51967 30169
rect 52001 30135 52167 30169
rect 52201 30135 52367 30169
rect 52401 30135 53478 30169
rect 33468 30132 53478 30135
rect 4958 30094 53478 30132
rect 55066 30094 55088 30210
rect 3348 30092 55088 30094
rect 20898 29996 20904 30048
rect 20956 30036 20962 30048
rect 22370 30036 22376 30048
rect 20956 30008 22376 30036
rect 20956 29996 20962 30008
rect 22370 29996 22376 30008
rect 22428 29996 22434 30048
rect 40328 30005 40356 30092
rect 40313 29999 40371 30005
rect 40313 29965 40325 29999
rect 40359 29965 40371 29999
rect 40313 29959 40371 29965
rect 16531 29901 16941 29913
rect 16531 29363 16539 29901
rect 16933 29363 16941 29901
rect 16531 29351 16941 29363
rect 18539 29901 18949 29913
rect 18539 29363 18546 29901
rect 18940 29363 18949 29901
rect 19275 29901 19685 29913
rect 19058 29384 19064 29436
rect 19116 29424 19122 29436
rect 19275 29424 19283 29901
rect 19116 29396 19283 29424
rect 19116 29384 19122 29396
rect 18539 29351 18949 29363
rect 19275 29363 19283 29396
rect 19677 29363 19685 29901
rect 19275 29351 19685 29363
rect 21283 29901 21693 29913
rect 21283 29363 21290 29901
rect 21684 29363 21693 29901
rect 21283 29351 21693 29363
rect 22019 29912 22429 29913
rect 22019 29901 22192 29912
rect 22244 29901 22429 29912
rect 22019 29363 22027 29901
rect 22421 29363 22429 29901
rect 22019 29351 22429 29363
rect 24027 29901 24437 29913
rect 24027 29363 24034 29901
rect 24428 29363 24437 29901
rect 24027 29351 24437 29363
rect 27213 29901 27623 29913
rect 27213 29363 27221 29901
rect 27615 29363 27623 29901
rect 27213 29351 27623 29363
rect 29221 29901 29631 29913
rect 29221 29363 29228 29901
rect 29622 29363 29631 29901
rect 29221 29351 29631 29363
rect 37513 29901 37559 29917
rect 37513 29867 37519 29901
rect 37553 29867 37559 29901
rect 37513 29829 37559 29867
rect 37513 29795 37519 29829
rect 37553 29795 37559 29829
rect 37513 29757 37559 29795
rect 37513 29723 37519 29757
rect 37553 29723 37559 29757
rect 37513 29685 37559 29723
rect 37513 29651 37519 29685
rect 37553 29651 37559 29685
rect 37513 29613 37559 29651
rect 37513 29579 37519 29613
rect 37553 29579 37559 29613
rect 37513 29541 37559 29579
rect 37513 29507 37519 29541
rect 37553 29507 37559 29541
rect 37513 29469 37559 29507
rect 37513 29435 37519 29469
rect 37553 29435 37559 29469
rect 37513 29397 37559 29435
rect 37513 29363 37519 29397
rect 37553 29363 37559 29397
rect 16531 28948 16941 28953
rect 18414 28948 18420 28960
rect 16531 28941 18420 28948
rect 16531 28403 16539 28941
rect 16933 28920 18420 28941
rect 16933 28403 16941 28920
rect 18414 28908 18420 28920
rect 18472 28908 18478 28960
rect 18528 28941 18960 29351
rect 16531 28391 16941 28403
rect 18528 28403 18546 28941
rect 18940 28403 18960 28941
rect 18528 28387 18960 28403
rect 19275 28948 19685 28953
rect 20898 28948 20904 28960
rect 19275 28941 20904 28948
rect 19275 28403 19283 28941
rect 19677 28920 20904 28941
rect 19677 28403 19685 28920
rect 20898 28908 20904 28920
rect 20956 28908 20962 28960
rect 21272 28941 21704 29351
rect 19275 28391 19685 28403
rect 21272 28403 21290 28941
rect 21684 28403 21704 28941
rect 21732 28960 21784 28966
rect 22019 28948 22429 28953
rect 21784 28941 22429 28948
rect 21784 28920 22027 28941
rect 21732 28902 21784 28908
rect 21272 28387 21704 28403
rect 22019 28403 22027 28920
rect 22421 28403 22429 28941
rect 22019 28391 22429 28403
rect 24016 28941 24448 29351
rect 24016 28403 24034 28941
rect 24428 28403 24448 28941
rect 24486 28908 24492 28960
rect 24544 28948 24550 28960
rect 27213 28948 27623 28953
rect 24544 28941 27623 28948
rect 24544 28920 27221 28941
rect 24544 28908 24550 28920
rect 24016 28387 24448 28403
rect 27213 28403 27221 28920
rect 27615 28403 27623 28941
rect 27213 28391 27623 28403
rect 29210 28941 29642 29351
rect 29210 28403 29228 28941
rect 29622 28403 29642 28941
rect 37513 29325 37559 29363
rect 37513 29291 37519 29325
rect 37553 29291 37559 29325
rect 37513 29253 37559 29291
rect 37513 29219 37519 29253
rect 37553 29219 37559 29253
rect 37513 29181 37559 29219
rect 37513 29147 37519 29181
rect 37553 29147 37559 29181
rect 37513 29109 37559 29147
rect 37513 29075 37519 29109
rect 37553 29075 37559 29109
rect 37513 29037 37559 29075
rect 37513 29003 37519 29037
rect 37553 29003 37559 29037
rect 37513 28965 37559 29003
rect 37513 28931 37519 28965
rect 37553 28931 37559 28965
rect 37513 28893 37559 28931
rect 37513 28859 37519 28893
rect 37553 28859 37559 28893
rect 37513 28821 37559 28859
rect 37513 28787 37519 28821
rect 37553 28787 37559 28821
rect 37513 28749 37559 28787
rect 37513 28715 37519 28749
rect 37553 28715 37559 28749
rect 37513 28677 37559 28715
rect 37513 28643 37519 28677
rect 37553 28643 37559 28677
rect 37513 28627 37559 28643
rect 37971 29901 38017 29917
rect 37971 29867 37977 29901
rect 38011 29867 38017 29901
rect 37971 29829 38017 29867
rect 37971 29795 37977 29829
rect 38011 29795 38017 29829
rect 37971 29757 38017 29795
rect 37971 29723 37977 29757
rect 38011 29723 38017 29757
rect 37971 29685 38017 29723
rect 37971 29651 37977 29685
rect 38011 29651 38017 29685
rect 37971 29613 38017 29651
rect 37971 29579 37977 29613
rect 38011 29579 38017 29613
rect 37971 29541 38017 29579
rect 37971 29507 37977 29541
rect 38011 29507 38017 29541
rect 37971 29469 38017 29507
rect 37971 29435 37977 29469
rect 38011 29435 38017 29469
rect 37971 29397 38017 29435
rect 37971 29363 37977 29397
rect 38011 29363 38017 29397
rect 37971 29325 38017 29363
rect 37971 29291 37977 29325
rect 38011 29291 38017 29325
rect 37971 29253 38017 29291
rect 37971 29219 37977 29253
rect 38011 29219 38017 29253
rect 37971 29181 38017 29219
rect 37971 29147 37977 29181
rect 38011 29147 38017 29181
rect 37971 29109 38017 29147
rect 37971 29075 37977 29109
rect 38011 29075 38017 29109
rect 37971 29037 38017 29075
rect 37971 29003 37977 29037
rect 38011 29003 38017 29037
rect 37971 28965 38017 29003
rect 37971 28931 37977 28965
rect 38011 28931 38017 28965
rect 37971 28893 38017 28931
rect 37971 28859 37977 28893
rect 38011 28859 38017 28893
rect 37971 28821 38017 28859
rect 37971 28787 37977 28821
rect 38011 28787 38017 28821
rect 37971 28749 38017 28787
rect 37971 28715 37977 28749
rect 38011 28715 38017 28749
rect 37971 28677 38017 28715
rect 37971 28643 37977 28677
rect 38011 28643 38017 28677
rect 37971 28627 38017 28643
rect 38429 29901 38475 29917
rect 38429 29867 38435 29901
rect 38469 29867 38475 29901
rect 38429 29829 38475 29867
rect 38429 29795 38435 29829
rect 38469 29795 38475 29829
rect 38429 29757 38475 29795
rect 38429 29723 38435 29757
rect 38469 29723 38475 29757
rect 38429 29685 38475 29723
rect 38429 29651 38435 29685
rect 38469 29651 38475 29685
rect 38429 29613 38475 29651
rect 38429 29579 38435 29613
rect 38469 29579 38475 29613
rect 38429 29541 38475 29579
rect 38429 29507 38435 29541
rect 38469 29507 38475 29541
rect 38429 29469 38475 29507
rect 38429 29435 38435 29469
rect 38469 29435 38475 29469
rect 38429 29397 38475 29435
rect 38429 29363 38435 29397
rect 38469 29363 38475 29397
rect 38429 29325 38475 29363
rect 38429 29291 38435 29325
rect 38469 29291 38475 29325
rect 38429 29253 38475 29291
rect 38429 29219 38435 29253
rect 38469 29219 38475 29253
rect 38429 29181 38475 29219
rect 38429 29147 38435 29181
rect 38469 29147 38475 29181
rect 38429 29109 38475 29147
rect 38429 29075 38435 29109
rect 38469 29075 38475 29109
rect 38429 29037 38475 29075
rect 38429 29003 38435 29037
rect 38469 29003 38475 29037
rect 38429 28965 38475 29003
rect 38429 28931 38435 28965
rect 38469 28931 38475 28965
rect 38429 28893 38475 28931
rect 38429 28859 38435 28893
rect 38469 28859 38475 28893
rect 38429 28821 38475 28859
rect 38429 28787 38435 28821
rect 38469 28787 38475 28821
rect 38429 28749 38475 28787
rect 38429 28715 38435 28749
rect 38469 28715 38475 28749
rect 38429 28677 38475 28715
rect 38429 28643 38435 28677
rect 38469 28643 38475 28677
rect 38429 28627 38475 28643
rect 38887 29901 38933 29917
rect 38887 29867 38893 29901
rect 38927 29867 38933 29901
rect 38887 29829 38933 29867
rect 38887 29795 38893 29829
rect 38927 29795 38933 29829
rect 38887 29757 38933 29795
rect 38887 29723 38893 29757
rect 38927 29723 38933 29757
rect 38887 29685 38933 29723
rect 38887 29651 38893 29685
rect 38927 29651 38933 29685
rect 38887 29613 38933 29651
rect 38887 29579 38893 29613
rect 38927 29579 38933 29613
rect 38887 29541 38933 29579
rect 38887 29507 38893 29541
rect 38927 29507 38933 29541
rect 38887 29469 38933 29507
rect 38887 29435 38893 29469
rect 38927 29435 38933 29469
rect 38887 29397 38933 29435
rect 38887 29363 38893 29397
rect 38927 29363 38933 29397
rect 38887 29325 38933 29363
rect 38887 29291 38893 29325
rect 38927 29291 38933 29325
rect 38887 29253 38933 29291
rect 38887 29219 38893 29253
rect 38927 29219 38933 29253
rect 38887 29181 38933 29219
rect 38887 29147 38893 29181
rect 38927 29147 38933 29181
rect 38887 29109 38933 29147
rect 38887 29075 38893 29109
rect 38927 29075 38933 29109
rect 38887 29037 38933 29075
rect 38887 29003 38893 29037
rect 38927 29003 38933 29037
rect 38887 28965 38933 29003
rect 38887 28931 38893 28965
rect 38927 28931 38933 28965
rect 38887 28893 38933 28931
rect 38887 28859 38893 28893
rect 38927 28859 38933 28893
rect 38887 28821 38933 28859
rect 38887 28787 38893 28821
rect 38927 28787 38933 28821
rect 38887 28749 38933 28787
rect 38887 28715 38893 28749
rect 38927 28715 38933 28749
rect 38887 28677 38933 28715
rect 38887 28643 38893 28677
rect 38927 28643 38933 28677
rect 38887 28627 38933 28643
rect 39345 29901 39391 29917
rect 39345 29867 39351 29901
rect 39385 29867 39391 29901
rect 39345 29829 39391 29867
rect 39345 29795 39351 29829
rect 39385 29795 39391 29829
rect 39345 29757 39391 29795
rect 39345 29723 39351 29757
rect 39385 29723 39391 29757
rect 39345 29685 39391 29723
rect 39345 29651 39351 29685
rect 39385 29651 39391 29685
rect 39345 29613 39391 29651
rect 39345 29579 39351 29613
rect 39385 29579 39391 29613
rect 39345 29541 39391 29579
rect 39345 29507 39351 29541
rect 39385 29507 39391 29541
rect 39345 29469 39391 29507
rect 39345 29435 39351 29469
rect 39385 29435 39391 29469
rect 39345 29397 39391 29435
rect 39345 29363 39351 29397
rect 39385 29363 39391 29397
rect 39345 29325 39391 29363
rect 39345 29291 39351 29325
rect 39385 29291 39391 29325
rect 39345 29253 39391 29291
rect 39345 29219 39351 29253
rect 39385 29219 39391 29253
rect 39345 29181 39391 29219
rect 39345 29147 39351 29181
rect 39385 29147 39391 29181
rect 39345 29109 39391 29147
rect 39345 29075 39351 29109
rect 39385 29075 39391 29109
rect 39345 29037 39391 29075
rect 39345 29003 39351 29037
rect 39385 29003 39391 29037
rect 39345 28965 39391 29003
rect 39345 28931 39351 28965
rect 39385 28931 39391 28965
rect 39345 28893 39391 28931
rect 39345 28859 39351 28893
rect 39385 28859 39391 28893
rect 39345 28821 39391 28859
rect 39345 28787 39351 28821
rect 39385 28787 39391 28821
rect 39345 28749 39391 28787
rect 39345 28715 39351 28749
rect 39385 28715 39391 28749
rect 39345 28677 39391 28715
rect 39345 28643 39351 28677
rect 39385 28643 39391 28677
rect 39345 28627 39391 28643
rect 39803 29901 39849 29917
rect 39803 29867 39809 29901
rect 39843 29867 39849 29901
rect 39803 29829 39849 29867
rect 39803 29795 39809 29829
rect 39843 29795 39849 29829
rect 39803 29757 39849 29795
rect 39803 29723 39809 29757
rect 39843 29723 39849 29757
rect 39803 29685 39849 29723
rect 39803 29651 39809 29685
rect 39843 29651 39849 29685
rect 39803 29613 39849 29651
rect 39803 29579 39809 29613
rect 39843 29579 39849 29613
rect 39803 29541 39849 29579
rect 39803 29507 39809 29541
rect 39843 29507 39849 29541
rect 39803 29469 39849 29507
rect 39803 29435 39809 29469
rect 39843 29435 39849 29469
rect 39803 29397 39849 29435
rect 39803 29363 39809 29397
rect 39843 29363 39849 29397
rect 39803 29325 39849 29363
rect 39803 29291 39809 29325
rect 39843 29291 39849 29325
rect 39803 29253 39849 29291
rect 39803 29219 39809 29253
rect 39843 29219 39849 29253
rect 39803 29181 39849 29219
rect 39803 29147 39809 29181
rect 39843 29147 39849 29181
rect 39803 29109 39849 29147
rect 39803 29075 39809 29109
rect 39843 29075 39849 29109
rect 39803 29037 39849 29075
rect 39803 29003 39809 29037
rect 39843 29003 39849 29037
rect 39803 28965 39849 29003
rect 39803 28931 39809 28965
rect 39843 28931 39849 28965
rect 39803 28893 39849 28931
rect 39803 28859 39809 28893
rect 39843 28859 39849 28893
rect 39803 28821 39849 28859
rect 39803 28787 39809 28821
rect 39843 28787 39849 28821
rect 39803 28749 39849 28787
rect 39803 28715 39809 28749
rect 39843 28715 39849 28749
rect 39803 28677 39849 28715
rect 39803 28643 39809 28677
rect 39843 28643 39849 28677
rect 39803 28627 39849 28643
rect 40261 29901 40307 29917
rect 40261 29867 40267 29901
rect 40301 29867 40307 29901
rect 40261 29829 40307 29867
rect 40261 29795 40267 29829
rect 40301 29795 40307 29829
rect 40261 29757 40307 29795
rect 41810 29836 52478 29842
rect 41810 29802 41830 29836
rect 41864 29802 41920 29836
rect 41954 29802 42010 29836
rect 42044 29802 42100 29836
rect 42134 29802 42190 29836
rect 42224 29802 42280 29836
rect 42314 29802 42370 29836
rect 42404 29802 42460 29836
rect 42494 29802 42550 29836
rect 42584 29802 42640 29836
rect 42674 29802 42730 29836
rect 42764 29802 42820 29836
rect 42854 29802 42910 29836
rect 42944 29802 43000 29836
rect 43034 29802 43170 29836
rect 43204 29802 43260 29836
rect 43294 29802 43350 29836
rect 43384 29802 43440 29836
rect 43474 29802 43530 29836
rect 43564 29802 43620 29836
rect 43654 29802 43710 29836
rect 43744 29802 43800 29836
rect 43834 29802 43890 29836
rect 43924 29802 43980 29836
rect 44014 29802 44070 29836
rect 44104 29802 44160 29836
rect 44194 29802 44250 29836
rect 44284 29802 44340 29836
rect 44374 29802 44510 29836
rect 44544 29802 44600 29836
rect 44634 29802 44690 29836
rect 44724 29802 44780 29836
rect 44814 29802 44870 29836
rect 44904 29802 44960 29836
rect 44994 29802 45050 29836
rect 45084 29802 45140 29836
rect 45174 29802 45230 29836
rect 45264 29802 45320 29836
rect 45354 29802 45410 29836
rect 45444 29802 45500 29836
rect 45534 29802 45590 29836
rect 45624 29802 45680 29836
rect 45714 29802 45850 29836
rect 45884 29802 45940 29836
rect 45974 29802 46030 29836
rect 46064 29802 46120 29836
rect 46154 29802 46210 29836
rect 46244 29802 46300 29836
rect 46334 29802 46390 29836
rect 46424 29802 46480 29836
rect 46514 29802 46570 29836
rect 46604 29802 46660 29836
rect 46694 29802 46750 29836
rect 46784 29802 46840 29836
rect 46874 29802 46930 29836
rect 46964 29802 47020 29836
rect 47054 29802 47190 29836
rect 47224 29802 47280 29836
rect 47314 29802 47370 29836
rect 47404 29802 47460 29836
rect 47494 29802 47550 29836
rect 47584 29802 47640 29836
rect 47674 29802 47730 29836
rect 47764 29802 47820 29836
rect 47854 29802 47910 29836
rect 47944 29802 48000 29836
rect 48034 29802 48090 29836
rect 48124 29802 48180 29836
rect 48214 29802 48270 29836
rect 48304 29802 48360 29836
rect 48394 29802 48530 29836
rect 48564 29802 48620 29836
rect 48654 29802 48710 29836
rect 48744 29802 48800 29836
rect 48834 29802 48890 29836
rect 48924 29802 48980 29836
rect 49014 29802 49070 29836
rect 49104 29802 49160 29836
rect 49194 29802 49250 29836
rect 49284 29802 49340 29836
rect 49374 29802 49430 29836
rect 49464 29802 49520 29836
rect 49554 29802 49610 29836
rect 49644 29802 49700 29836
rect 49734 29802 49870 29836
rect 49904 29802 49960 29836
rect 49994 29802 50050 29836
rect 50084 29802 50140 29836
rect 50174 29802 50230 29836
rect 50264 29802 50320 29836
rect 50354 29802 50410 29836
rect 50444 29802 50500 29836
rect 50534 29802 50590 29836
rect 50624 29802 50680 29836
rect 50714 29802 50770 29836
rect 50804 29802 50860 29836
rect 50894 29802 50950 29836
rect 50984 29802 51040 29836
rect 51074 29802 51210 29836
rect 51244 29802 51300 29836
rect 51334 29802 51390 29836
rect 51424 29802 51480 29836
rect 51514 29802 51570 29836
rect 51604 29802 51660 29836
rect 51694 29802 51750 29836
rect 51784 29802 51840 29836
rect 51874 29802 51930 29836
rect 51964 29802 52020 29836
rect 52054 29802 52110 29836
rect 52144 29802 52200 29836
rect 52234 29802 52290 29836
rect 52324 29802 52380 29836
rect 52414 29802 52478 29836
rect 41810 29772 52478 29802
rect 40261 29723 40267 29757
rect 40301 29723 40307 29757
rect 40261 29685 40307 29723
rect 42168 29708 42196 29772
rect 42150 29692 42156 29708
rect 40261 29651 40267 29685
rect 40301 29651 40307 29685
rect 40261 29613 40307 29651
rect 41974 29676 42156 29692
rect 42208 29692 42214 29708
rect 42208 29676 52314 29692
rect 41974 29642 41994 29676
rect 42028 29642 42084 29676
rect 42118 29656 42156 29676
rect 42118 29642 42174 29656
rect 42208 29642 42264 29676
rect 42298 29642 42354 29676
rect 42388 29642 42444 29676
rect 42478 29642 42534 29676
rect 42568 29642 42624 29676
rect 42658 29642 42714 29676
rect 42748 29642 42804 29676
rect 42838 29642 42894 29676
rect 42928 29642 43334 29676
rect 43368 29642 43424 29676
rect 43458 29642 43514 29676
rect 43548 29642 43604 29676
rect 43638 29642 43694 29676
rect 43728 29642 43784 29676
rect 43818 29642 43874 29676
rect 43908 29642 43964 29676
rect 43998 29642 44054 29676
rect 44088 29642 44144 29676
rect 44178 29642 44234 29676
rect 44268 29642 44674 29676
rect 44708 29642 44764 29676
rect 44798 29642 44854 29676
rect 44888 29642 44944 29676
rect 44978 29642 45034 29676
rect 45068 29642 45124 29676
rect 45158 29642 45214 29676
rect 45248 29642 45304 29676
rect 45338 29642 45394 29676
rect 45428 29642 45484 29676
rect 45518 29642 45574 29676
rect 45608 29642 46014 29676
rect 46048 29642 46104 29676
rect 46138 29642 46194 29676
rect 46228 29642 46284 29676
rect 46318 29642 46374 29676
rect 46408 29642 46464 29676
rect 46498 29642 46554 29676
rect 46588 29642 46644 29676
rect 46678 29642 46734 29676
rect 46768 29642 46824 29676
rect 46858 29642 46914 29676
rect 46948 29642 47354 29676
rect 47388 29642 47444 29676
rect 47478 29642 47534 29676
rect 47568 29642 47624 29676
rect 47658 29642 47714 29676
rect 47748 29642 47804 29676
rect 47838 29642 47894 29676
rect 47928 29642 47984 29676
rect 48018 29642 48074 29676
rect 48108 29642 48164 29676
rect 48198 29642 48254 29676
rect 48288 29642 48694 29676
rect 48728 29642 48784 29676
rect 48818 29642 48874 29676
rect 48908 29642 48964 29676
rect 48998 29642 49054 29676
rect 49088 29642 49144 29676
rect 49178 29642 49234 29676
rect 49268 29642 49324 29676
rect 49358 29642 49414 29676
rect 49448 29642 49504 29676
rect 49538 29642 49594 29676
rect 49628 29642 50034 29676
rect 50068 29642 50124 29676
rect 50158 29642 50214 29676
rect 50248 29642 50304 29676
rect 50338 29642 50394 29676
rect 50428 29642 50484 29676
rect 50518 29642 50574 29676
rect 50608 29642 50664 29676
rect 50698 29642 50754 29676
rect 50788 29642 50844 29676
rect 50878 29642 50934 29676
rect 50968 29642 51374 29676
rect 51408 29642 51464 29676
rect 51498 29642 51554 29676
rect 51588 29642 51644 29676
rect 51678 29642 51734 29676
rect 51768 29642 51824 29676
rect 51858 29642 51914 29676
rect 51948 29642 52004 29676
rect 52038 29642 52094 29676
rect 52128 29642 52184 29676
rect 52218 29642 52274 29676
rect 52308 29642 52314 29676
rect 41974 29622 52314 29642
rect 40261 29579 40267 29613
rect 40301 29579 40307 29613
rect 40261 29541 40307 29579
rect 40261 29507 40267 29541
rect 40301 29507 40307 29541
rect 40261 29469 40307 29507
rect 40261 29435 40267 29469
rect 40301 29435 40307 29469
rect 40261 29397 40307 29435
rect 40261 29363 40267 29397
rect 40301 29363 40307 29397
rect 40261 29325 40307 29363
rect 40261 29291 40267 29325
rect 40301 29291 40307 29325
rect 40261 29253 40307 29291
rect 40261 29219 40267 29253
rect 40301 29219 40307 29253
rect 40261 29181 40307 29219
rect 40261 29147 40267 29181
rect 40301 29147 40307 29181
rect 40261 29109 40307 29147
rect 40261 29075 40267 29109
rect 40301 29075 40307 29109
rect 40261 29037 40307 29075
rect 40261 29003 40267 29037
rect 40301 29003 40307 29037
rect 40261 28965 40307 29003
rect 40261 28931 40267 28965
rect 40301 28931 40307 28965
rect 40261 28893 40307 28931
rect 42148 29504 52140 29518
rect 42148 29472 42248 29504
rect 42300 29472 52140 29504
rect 42148 29438 42180 29472
rect 42214 29452 42248 29472
rect 42214 29438 42280 29452
rect 42314 29438 42380 29472
rect 42414 29438 42480 29472
rect 42514 29438 42580 29472
rect 42614 29438 42680 29472
rect 42714 29438 43520 29472
rect 43554 29438 43620 29472
rect 43654 29438 43720 29472
rect 43754 29438 43820 29472
rect 43854 29438 43920 29472
rect 43954 29438 44020 29472
rect 44054 29438 44860 29472
rect 44894 29438 44960 29472
rect 44994 29438 45060 29472
rect 45094 29438 45160 29472
rect 45194 29438 45260 29472
rect 45294 29438 45360 29472
rect 45394 29438 46200 29472
rect 46234 29438 46300 29472
rect 46334 29438 46400 29472
rect 46434 29438 46500 29472
rect 46534 29438 46600 29472
rect 46634 29438 46700 29472
rect 46734 29438 47540 29472
rect 47574 29438 47640 29472
rect 47674 29438 47740 29472
rect 47774 29438 47840 29472
rect 47874 29438 47940 29472
rect 47974 29438 48040 29472
rect 48074 29438 48880 29472
rect 48914 29438 48980 29472
rect 49014 29438 49080 29472
rect 49114 29438 49180 29472
rect 49214 29438 49280 29472
rect 49314 29438 49380 29472
rect 49414 29438 50220 29472
rect 50254 29438 50320 29472
rect 50354 29438 50420 29472
rect 50454 29438 50520 29472
rect 50554 29438 50620 29472
rect 50654 29438 50720 29472
rect 50754 29438 51560 29472
rect 51594 29438 51660 29472
rect 51694 29438 51760 29472
rect 51794 29438 51860 29472
rect 51894 29438 51960 29472
rect 51994 29438 52060 29472
rect 52094 29438 52140 29472
rect 42148 29372 52140 29438
rect 42148 29338 42180 29372
rect 42214 29338 42280 29372
rect 42314 29338 42380 29372
rect 42414 29338 42480 29372
rect 42514 29338 42580 29372
rect 42614 29338 42680 29372
rect 42714 29338 43520 29372
rect 43554 29338 43620 29372
rect 43654 29338 43720 29372
rect 43754 29338 43820 29372
rect 43854 29338 43920 29372
rect 43954 29338 44020 29372
rect 44054 29338 44860 29372
rect 44894 29338 44960 29372
rect 44994 29338 45060 29372
rect 45094 29338 45160 29372
rect 45194 29338 45260 29372
rect 45294 29338 45360 29372
rect 45394 29338 46200 29372
rect 46234 29338 46300 29372
rect 46334 29338 46400 29372
rect 46434 29338 46500 29372
rect 46534 29338 46600 29372
rect 46634 29338 46700 29372
rect 46734 29338 47540 29372
rect 47574 29338 47640 29372
rect 47674 29338 47740 29372
rect 47774 29338 47840 29372
rect 47874 29338 47940 29372
rect 47974 29338 48040 29372
rect 48074 29338 48880 29372
rect 48914 29338 48980 29372
rect 49014 29338 49080 29372
rect 49114 29338 49180 29372
rect 49214 29338 49280 29372
rect 49314 29338 49380 29372
rect 49414 29338 50220 29372
rect 50254 29338 50320 29372
rect 50354 29338 50420 29372
rect 50454 29338 50520 29372
rect 50554 29338 50620 29372
rect 50654 29338 50720 29372
rect 50754 29338 51560 29372
rect 51594 29338 51660 29372
rect 51694 29338 51760 29372
rect 51794 29338 51860 29372
rect 51894 29338 51960 29372
rect 51994 29338 52060 29372
rect 52094 29338 52140 29372
rect 42148 29272 52140 29338
rect 42148 29238 42180 29272
rect 42214 29238 42280 29272
rect 42314 29238 42380 29272
rect 42414 29238 42480 29272
rect 42514 29238 42580 29272
rect 42614 29238 42680 29272
rect 42714 29238 43520 29272
rect 43554 29238 43620 29272
rect 43654 29238 43720 29272
rect 43754 29238 43820 29272
rect 43854 29238 43920 29272
rect 43954 29238 44020 29272
rect 44054 29238 44860 29272
rect 44894 29238 44960 29272
rect 44994 29238 45060 29272
rect 45094 29238 45160 29272
rect 45194 29238 45260 29272
rect 45294 29238 45360 29272
rect 45394 29238 46200 29272
rect 46234 29238 46300 29272
rect 46334 29238 46400 29272
rect 46434 29238 46500 29272
rect 46534 29238 46600 29272
rect 46634 29238 46700 29272
rect 46734 29238 47540 29272
rect 47574 29238 47640 29272
rect 47674 29238 47740 29272
rect 47774 29238 47840 29272
rect 47874 29238 47940 29272
rect 47974 29238 48040 29272
rect 48074 29238 48880 29272
rect 48914 29238 48980 29272
rect 49014 29238 49080 29272
rect 49114 29238 49180 29272
rect 49214 29238 49280 29272
rect 49314 29238 49380 29272
rect 49414 29238 50220 29272
rect 50254 29238 50320 29272
rect 50354 29238 50420 29272
rect 50454 29238 50520 29272
rect 50554 29238 50620 29272
rect 50654 29238 50720 29272
rect 50754 29238 51560 29272
rect 51594 29238 51660 29272
rect 51694 29238 51760 29272
rect 51794 29238 51860 29272
rect 51894 29238 51960 29272
rect 51994 29238 52060 29272
rect 52094 29238 52140 29272
rect 42148 29172 52140 29238
rect 42148 29138 42180 29172
rect 42214 29138 42280 29172
rect 42314 29138 42380 29172
rect 42414 29138 42480 29172
rect 42514 29138 42580 29172
rect 42614 29138 42680 29172
rect 42714 29138 43520 29172
rect 43554 29138 43620 29172
rect 43654 29138 43720 29172
rect 43754 29138 43820 29172
rect 43854 29138 43920 29172
rect 43954 29138 44020 29172
rect 44054 29138 44860 29172
rect 44894 29138 44960 29172
rect 44994 29138 45060 29172
rect 45094 29138 45160 29172
rect 45194 29138 45260 29172
rect 45294 29138 45360 29172
rect 45394 29138 46200 29172
rect 46234 29138 46300 29172
rect 46334 29138 46400 29172
rect 46434 29138 46500 29172
rect 46534 29138 46600 29172
rect 46634 29138 46700 29172
rect 46734 29138 47540 29172
rect 47574 29138 47640 29172
rect 47674 29138 47740 29172
rect 47774 29138 47840 29172
rect 47874 29138 47940 29172
rect 47974 29138 48040 29172
rect 48074 29138 48880 29172
rect 48914 29138 48980 29172
rect 49014 29138 49080 29172
rect 49114 29138 49180 29172
rect 49214 29138 49280 29172
rect 49314 29138 49380 29172
rect 49414 29138 50220 29172
rect 50254 29138 50320 29172
rect 50354 29138 50420 29172
rect 50454 29138 50520 29172
rect 50554 29138 50620 29172
rect 50654 29138 50720 29172
rect 50754 29138 51560 29172
rect 51594 29138 51660 29172
rect 51694 29138 51760 29172
rect 51794 29138 51860 29172
rect 51894 29138 51960 29172
rect 51994 29138 52060 29172
rect 52094 29138 52140 29172
rect 42148 29072 52140 29138
rect 42148 29038 42180 29072
rect 42214 29038 42280 29072
rect 42314 29038 42380 29072
rect 42414 29038 42480 29072
rect 42514 29038 42580 29072
rect 42614 29038 42680 29072
rect 42714 29038 43520 29072
rect 43554 29038 43620 29072
rect 43654 29038 43720 29072
rect 43754 29038 43820 29072
rect 43854 29038 43920 29072
rect 43954 29038 44020 29072
rect 44054 29038 44860 29072
rect 44894 29038 44960 29072
rect 44994 29038 45060 29072
rect 45094 29038 45160 29072
rect 45194 29038 45260 29072
rect 45294 29038 45360 29072
rect 45394 29038 46200 29072
rect 46234 29038 46300 29072
rect 46334 29038 46400 29072
rect 46434 29038 46500 29072
rect 46534 29038 46600 29072
rect 46634 29038 46700 29072
rect 46734 29038 47540 29072
rect 47574 29038 47640 29072
rect 47674 29038 47740 29072
rect 47774 29038 47840 29072
rect 47874 29038 47940 29072
rect 47974 29038 48040 29072
rect 48074 29038 48880 29072
rect 48914 29038 48980 29072
rect 49014 29038 49080 29072
rect 49114 29038 49180 29072
rect 49214 29038 49280 29072
rect 49314 29038 49380 29072
rect 49414 29038 50220 29072
rect 50254 29038 50320 29072
rect 50354 29038 50420 29072
rect 50454 29038 50520 29072
rect 50554 29038 50620 29072
rect 50654 29038 50720 29072
rect 50754 29038 51560 29072
rect 51594 29038 51660 29072
rect 51694 29038 51760 29072
rect 51794 29038 51860 29072
rect 51894 29038 51960 29072
rect 51994 29038 52060 29072
rect 52094 29038 52140 29072
rect 42148 28972 52140 29038
rect 42148 28938 42180 28972
rect 42214 28938 42280 28972
rect 42314 28938 42380 28972
rect 42414 28938 42480 28972
rect 42514 28938 42580 28972
rect 42614 28938 42680 28972
rect 42714 28938 43520 28972
rect 43554 28938 43620 28972
rect 43654 28938 43720 28972
rect 43754 28938 43820 28972
rect 43854 28938 43920 28972
rect 43954 28938 44020 28972
rect 44054 28938 44860 28972
rect 44894 28938 44960 28972
rect 44994 28938 45060 28972
rect 45094 28938 45160 28972
rect 45194 28938 45260 28972
rect 45294 28938 45360 28972
rect 45394 28938 46200 28972
rect 46234 28938 46300 28972
rect 46334 28938 46400 28972
rect 46434 28938 46500 28972
rect 46534 28938 46600 28972
rect 46634 28938 46700 28972
rect 46734 28938 47540 28972
rect 47574 28938 47640 28972
rect 47674 28938 47740 28972
rect 47774 28938 47840 28972
rect 47874 28938 47940 28972
rect 47974 28938 48040 28972
rect 48074 28960 48880 28972
rect 48074 28938 48412 28960
rect 42148 28908 48412 28938
rect 48464 28938 48880 28960
rect 48914 28938 48980 28972
rect 49014 28938 49080 28972
rect 49114 28938 49180 28972
rect 49214 28938 49280 28972
rect 49314 28938 49380 28972
rect 49414 28938 50220 28972
rect 50254 28938 50320 28972
rect 50354 28938 50420 28972
rect 50454 28938 50520 28972
rect 50554 28938 50620 28972
rect 50654 28938 50720 28972
rect 50754 28938 51560 28972
rect 51594 28938 51660 28972
rect 51694 28938 51760 28972
rect 51794 28938 51860 28972
rect 51894 28938 51960 28972
rect 51994 28938 52060 28972
rect 52094 28938 52140 28972
rect 48464 28908 52140 28938
rect 42148 28906 52140 28908
rect 40261 28859 40267 28893
rect 40301 28859 40307 28893
rect 40261 28821 40307 28859
rect 40261 28787 40267 28821
rect 40301 28787 40307 28821
rect 40261 28749 40307 28787
rect 40261 28715 40267 28749
rect 40301 28715 40307 28749
rect 40261 28677 40307 28715
rect 40261 28643 40267 28677
rect 40301 28643 40307 28677
rect 40261 28627 40307 28643
rect 38565 28543 38623 28549
rect 38565 28509 38577 28543
rect 38611 28509 38623 28543
rect 38565 28503 38623 28509
rect 38580 28416 38608 28503
rect 38562 28404 38568 28416
rect 29210 28387 29642 28403
rect 38507 28376 38568 28404
rect 38562 28364 38568 28376
rect 38620 28364 38626 28416
rect 900 28330 57536 28332
rect 900 28214 922 28330
rect 2510 28289 55926 28330
rect 2510 28255 16703 28289
rect 16737 28255 16903 28289
rect 16937 28255 17103 28289
rect 17137 28255 17303 28289
rect 17337 28255 17503 28289
rect 17537 28255 17703 28289
rect 17737 28255 17903 28289
rect 17937 28255 18103 28289
rect 18137 28255 18303 28289
rect 18337 28255 18503 28289
rect 18537 28255 18703 28289
rect 18737 28255 19447 28289
rect 19481 28255 19647 28289
rect 19681 28255 19847 28289
rect 19881 28255 20047 28289
rect 20081 28255 20247 28289
rect 20281 28255 20447 28289
rect 20481 28255 20647 28289
rect 20681 28255 20847 28289
rect 20881 28255 21047 28289
rect 21081 28255 21247 28289
rect 21281 28255 21447 28289
rect 21481 28255 22191 28289
rect 22225 28255 22391 28289
rect 22425 28255 22591 28289
rect 22625 28255 22791 28289
rect 22825 28255 22991 28289
rect 23025 28255 23191 28289
rect 23225 28255 23391 28289
rect 23425 28255 23591 28289
rect 23625 28255 23791 28289
rect 23825 28255 23991 28289
rect 24025 28255 24191 28289
rect 24225 28255 27385 28289
rect 27419 28255 27585 28289
rect 27619 28255 27785 28289
rect 27819 28255 27985 28289
rect 28019 28255 28185 28289
rect 28219 28255 28385 28289
rect 28419 28255 28585 28289
rect 28619 28255 28785 28289
rect 28819 28255 28985 28289
rect 29019 28255 29185 28289
rect 29219 28255 29385 28289
rect 29419 28255 30111 28289
rect 30145 28255 30511 28289
rect 30545 28255 30911 28289
rect 30945 28255 31311 28289
rect 31345 28255 31711 28289
rect 31745 28255 32111 28289
rect 32145 28255 32511 28289
rect 32545 28255 32911 28289
rect 32945 28255 33311 28289
rect 33345 28255 33711 28289
rect 33745 28255 34111 28289
rect 34145 28255 34511 28289
rect 34545 28255 34911 28289
rect 34945 28255 35311 28289
rect 35345 28255 35711 28289
rect 35745 28255 36111 28289
rect 36145 28255 36511 28289
rect 36545 28255 36911 28289
rect 36945 28255 37655 28289
rect 37689 28255 38055 28289
rect 38089 28255 38455 28289
rect 38489 28255 38855 28289
rect 38889 28255 39255 28289
rect 39289 28255 39655 28289
rect 39689 28255 40055 28289
rect 40089 28255 41967 28289
rect 42001 28280 42167 28289
rect 42201 28280 42367 28289
rect 42001 28255 42156 28280
rect 42208 28255 42367 28280
rect 42401 28255 42567 28289
rect 42601 28255 42767 28289
rect 42801 28255 42967 28289
rect 43001 28255 43167 28289
rect 43201 28255 43367 28289
rect 43401 28255 43567 28289
rect 43601 28255 43767 28289
rect 43801 28255 43967 28289
rect 44001 28255 44167 28289
rect 44201 28255 44367 28289
rect 44401 28255 44567 28289
rect 44601 28255 44767 28289
rect 44801 28255 44967 28289
rect 45001 28255 45167 28289
rect 45201 28255 45367 28289
rect 45401 28255 45567 28289
rect 45601 28255 45767 28289
rect 45801 28255 45967 28289
rect 46001 28255 46167 28289
rect 46201 28255 46367 28289
rect 46401 28255 46567 28289
rect 46601 28255 46767 28289
rect 46801 28255 46967 28289
rect 47001 28255 47167 28289
rect 47201 28255 47367 28289
rect 47401 28255 47567 28289
rect 47601 28255 47767 28289
rect 47801 28255 47967 28289
rect 48001 28255 48167 28289
rect 48201 28255 48367 28289
rect 48401 28255 48567 28289
rect 48601 28255 48767 28289
rect 48801 28255 48967 28289
rect 49001 28255 49167 28289
rect 49201 28255 49367 28289
rect 49401 28255 49567 28289
rect 49601 28255 49767 28289
rect 49801 28255 49967 28289
rect 50001 28255 50167 28289
rect 50201 28255 50367 28289
rect 50401 28255 50567 28289
rect 50601 28255 50767 28289
rect 50801 28255 50967 28289
rect 51001 28255 51167 28289
rect 51201 28255 51367 28289
rect 51401 28255 51567 28289
rect 51601 28255 51767 28289
rect 51801 28255 51967 28289
rect 52001 28255 52167 28289
rect 52201 28255 52367 28289
rect 52401 28255 55926 28289
rect 2510 28228 42156 28255
rect 42208 28228 55926 28255
rect 2510 28214 55926 28228
rect 57514 28214 57536 28330
rect 900 28212 57536 28214
rect 3348 26450 55088 26452
rect 3348 26334 3370 26450
rect 4958 26444 53478 26450
rect 4958 26409 33416 26444
rect 4958 26375 22583 26409
rect 22617 26375 22783 26409
rect 22817 26375 22983 26409
rect 23017 26375 23183 26409
rect 23217 26375 23383 26409
rect 23417 26375 23583 26409
rect 23617 26375 23783 26409
rect 23817 26375 23983 26409
rect 24017 26375 24183 26409
rect 24217 26375 24383 26409
rect 24417 26375 24583 26409
rect 24617 26375 25601 26409
rect 25635 26375 26001 26409
rect 26035 26375 26401 26409
rect 26435 26375 26801 26409
rect 26835 26375 27201 26409
rect 27235 26375 27601 26409
rect 27635 26375 28001 26409
rect 28035 26375 28401 26409
rect 28435 26375 28801 26409
rect 28835 26375 29201 26409
rect 29235 26375 30111 26409
rect 30145 26375 30511 26409
rect 30545 26375 30911 26409
rect 30945 26375 31311 26409
rect 31345 26375 31711 26409
rect 31745 26375 32111 26409
rect 32145 26375 32511 26409
rect 32545 26375 32911 26409
rect 32945 26375 33311 26409
rect 33345 26392 33416 26409
rect 33468 26409 53478 26444
rect 33468 26392 33711 26409
rect 33345 26375 33711 26392
rect 33745 26375 34111 26409
rect 34145 26375 34511 26409
rect 34545 26375 34911 26409
rect 34945 26375 35311 26409
rect 35345 26375 35711 26409
rect 35745 26375 36111 26409
rect 36145 26375 36511 26409
rect 36545 26375 36911 26409
rect 36945 26375 37577 26409
rect 37611 26375 37777 26409
rect 37811 26375 37977 26409
rect 38011 26375 38177 26409
rect 38211 26375 38377 26409
rect 38411 26375 38577 26409
rect 38611 26375 38777 26409
rect 38811 26375 38977 26409
rect 39011 26375 39177 26409
rect 39211 26375 39377 26409
rect 39411 26375 39577 26409
rect 39611 26375 40321 26409
rect 40355 26375 40521 26409
rect 40555 26375 40721 26409
rect 40755 26375 40921 26409
rect 40955 26375 41121 26409
rect 41155 26375 41321 26409
rect 41355 26375 41521 26409
rect 41555 26375 41721 26409
rect 41755 26375 41921 26409
rect 41955 26375 42121 26409
rect 42155 26375 42321 26409
rect 42355 26375 43065 26409
rect 43099 26375 43265 26409
rect 43299 26375 43465 26409
rect 43499 26375 43665 26409
rect 43699 26375 43865 26409
rect 43899 26375 44065 26409
rect 44099 26375 44265 26409
rect 44299 26375 44465 26409
rect 44499 26375 44665 26409
rect 44699 26375 44865 26409
rect 44899 26375 45065 26409
rect 45099 26375 45809 26409
rect 45843 26375 46009 26409
rect 46043 26375 46209 26409
rect 46243 26375 46409 26409
rect 46443 26375 46609 26409
rect 46643 26375 46809 26409
rect 46843 26375 47009 26409
rect 47043 26375 47209 26409
rect 47243 26375 47409 26409
rect 47443 26375 47609 26409
rect 47643 26375 47809 26409
rect 47843 26375 48553 26409
rect 48587 26375 48753 26409
rect 48787 26375 48953 26409
rect 48987 26375 49153 26409
rect 49187 26375 49353 26409
rect 49387 26375 49553 26409
rect 49587 26375 49753 26409
rect 49787 26375 49953 26409
rect 49987 26375 50153 26409
rect 50187 26375 50353 26409
rect 50387 26375 50553 26409
rect 50587 26375 53478 26409
rect 4958 26334 53478 26375
rect 55066 26334 55088 26450
rect 3348 26332 55088 26334
rect 39942 26228 39948 26240
rect 37752 26200 39948 26228
rect 37752 26153 37780 26200
rect 39942 26188 39948 26200
rect 40000 26188 40006 26240
rect 41432 26200 45692 26228
rect 41432 26172 41460 26200
rect 22411 26141 22821 26153
rect 13906 25848 13912 25900
rect 13964 25888 13970 25900
rect 22411 25888 22419 26141
rect 13964 25860 22419 25888
rect 13964 25848 13970 25860
rect 22411 25603 22419 25860
rect 22813 25603 22821 26141
rect 22411 25591 22821 25603
rect 24419 26141 24829 26153
rect 24419 25603 24426 26141
rect 24820 25603 24829 26141
rect 37405 26141 37815 26153
rect 24419 25591 24829 25603
rect 25424 25889 25470 25912
rect 25424 25855 25430 25889
rect 25464 25855 25470 25889
rect 25424 25817 25470 25855
rect 25424 25783 25430 25817
rect 25464 25783 25470 25817
rect 25424 25745 25470 25783
rect 25424 25711 25430 25745
rect 25464 25711 25470 25745
rect 25424 25673 25470 25711
rect 25424 25639 25430 25673
rect 25464 25639 25470 25673
rect 25424 25601 25470 25639
rect 22411 25181 22821 25193
rect 22411 24643 22419 25181
rect 22813 24664 22821 25181
rect 24408 25181 24840 25591
rect 22922 24664 22928 24676
rect 22813 24643 22928 24664
rect 22411 24636 22928 24643
rect 22411 24631 22821 24636
rect 22922 24624 22928 24636
rect 22980 24624 22986 24676
rect 24408 24643 24426 25181
rect 24820 24643 24840 25181
rect 25424 25567 25430 25601
rect 25464 25567 25470 25601
rect 25424 25529 25470 25567
rect 25424 25495 25430 25529
rect 25464 25495 25470 25529
rect 25424 25457 25470 25495
rect 25424 25423 25430 25457
rect 25464 25423 25470 25457
rect 25424 25385 25470 25423
rect 25424 25351 25430 25385
rect 25464 25351 25470 25385
rect 25424 25313 25470 25351
rect 25424 25279 25430 25313
rect 25464 25279 25470 25313
rect 25424 25241 25470 25279
rect 25424 25207 25430 25241
rect 25464 25207 25470 25241
rect 25424 25169 25470 25207
rect 25424 25152 25430 25169
rect 25406 25100 25412 25152
rect 25464 25100 25470 25169
rect 25882 25889 25928 25912
rect 25882 25855 25888 25889
rect 25922 25855 25928 25889
rect 25882 25817 25928 25855
rect 25882 25783 25888 25817
rect 25922 25783 25928 25817
rect 25882 25745 25928 25783
rect 25882 25711 25888 25745
rect 25922 25711 25928 25745
rect 25882 25673 25928 25711
rect 25882 25639 25888 25673
rect 25922 25639 25928 25673
rect 25882 25601 25928 25639
rect 25882 25567 25888 25601
rect 25922 25567 25928 25601
rect 25882 25529 25928 25567
rect 25882 25495 25888 25529
rect 25922 25495 25928 25529
rect 25882 25457 25928 25495
rect 25882 25423 25888 25457
rect 25922 25423 25928 25457
rect 25882 25385 25928 25423
rect 25882 25351 25888 25385
rect 25922 25351 25928 25385
rect 25882 25313 25928 25351
rect 25882 25279 25888 25313
rect 25922 25279 25928 25313
rect 25882 25241 25928 25279
rect 25882 25207 25888 25241
rect 25922 25207 25928 25241
rect 25882 25169 25928 25207
rect 25882 25135 25888 25169
rect 25922 25135 25928 25169
rect 25882 25112 25928 25135
rect 26340 25889 26386 25912
rect 26340 25855 26346 25889
rect 26380 25855 26386 25889
rect 26340 25817 26386 25855
rect 26340 25783 26346 25817
rect 26380 25783 26386 25817
rect 26340 25745 26386 25783
rect 26340 25711 26346 25745
rect 26380 25711 26386 25745
rect 26340 25673 26386 25711
rect 26340 25639 26346 25673
rect 26380 25639 26386 25673
rect 26340 25601 26386 25639
rect 26340 25567 26346 25601
rect 26380 25567 26386 25601
rect 26340 25529 26386 25567
rect 26340 25495 26346 25529
rect 26380 25495 26386 25529
rect 26340 25457 26386 25495
rect 26340 25423 26346 25457
rect 26380 25423 26386 25457
rect 26340 25385 26386 25423
rect 26340 25351 26346 25385
rect 26380 25351 26386 25385
rect 26340 25313 26386 25351
rect 26340 25279 26346 25313
rect 26380 25279 26386 25313
rect 26340 25241 26386 25279
rect 26340 25207 26346 25241
rect 26380 25207 26386 25241
rect 26340 25169 26386 25207
rect 26340 25135 26346 25169
rect 26380 25135 26386 25169
rect 26340 25112 26386 25135
rect 26798 25889 26844 25912
rect 26798 25855 26804 25889
rect 26838 25855 26844 25889
rect 26798 25817 26844 25855
rect 26798 25783 26804 25817
rect 26838 25783 26844 25817
rect 26798 25745 26844 25783
rect 26798 25711 26804 25745
rect 26838 25711 26844 25745
rect 26798 25673 26844 25711
rect 26798 25639 26804 25673
rect 26838 25639 26844 25673
rect 26798 25601 26844 25639
rect 26798 25567 26804 25601
rect 26838 25567 26844 25601
rect 26798 25529 26844 25567
rect 26798 25495 26804 25529
rect 26838 25495 26844 25529
rect 26798 25457 26844 25495
rect 26798 25423 26804 25457
rect 26838 25423 26844 25457
rect 26798 25385 26844 25423
rect 26798 25351 26804 25385
rect 26838 25351 26844 25385
rect 26798 25313 26844 25351
rect 26798 25279 26804 25313
rect 26838 25279 26844 25313
rect 26798 25241 26844 25279
rect 26798 25207 26804 25241
rect 26838 25207 26844 25241
rect 26798 25169 26844 25207
rect 26798 25135 26804 25169
rect 26838 25135 26844 25169
rect 26798 25112 26844 25135
rect 27256 25889 27302 25912
rect 27256 25855 27262 25889
rect 27296 25855 27302 25889
rect 27256 25817 27302 25855
rect 27256 25783 27262 25817
rect 27296 25783 27302 25817
rect 27256 25745 27302 25783
rect 27256 25711 27262 25745
rect 27296 25711 27302 25745
rect 27256 25673 27302 25711
rect 27256 25639 27262 25673
rect 27296 25639 27302 25673
rect 27256 25601 27302 25639
rect 27256 25567 27262 25601
rect 27296 25567 27302 25601
rect 27256 25529 27302 25567
rect 27256 25495 27262 25529
rect 27296 25495 27302 25529
rect 27256 25457 27302 25495
rect 27256 25423 27262 25457
rect 27296 25423 27302 25457
rect 27256 25385 27302 25423
rect 27256 25351 27262 25385
rect 27296 25351 27302 25385
rect 27256 25313 27302 25351
rect 27256 25279 27262 25313
rect 27296 25279 27302 25313
rect 27256 25241 27302 25279
rect 27256 25207 27262 25241
rect 27296 25207 27302 25241
rect 27256 25169 27302 25207
rect 27256 25135 27262 25169
rect 27296 25135 27302 25169
rect 27256 25112 27302 25135
rect 27714 25889 27760 25912
rect 27714 25855 27720 25889
rect 27754 25855 27760 25889
rect 27714 25817 27760 25855
rect 27714 25783 27720 25817
rect 27754 25783 27760 25817
rect 27714 25745 27760 25783
rect 27714 25711 27720 25745
rect 27754 25711 27760 25745
rect 27714 25673 27760 25711
rect 27714 25639 27720 25673
rect 27754 25639 27760 25673
rect 27714 25601 27760 25639
rect 27714 25567 27720 25601
rect 27754 25567 27760 25601
rect 27714 25529 27760 25567
rect 27714 25495 27720 25529
rect 27754 25495 27760 25529
rect 27714 25457 27760 25495
rect 27714 25423 27720 25457
rect 27754 25423 27760 25457
rect 27714 25385 27760 25423
rect 27714 25351 27720 25385
rect 27754 25351 27760 25385
rect 27714 25313 27760 25351
rect 27714 25279 27720 25313
rect 27754 25279 27760 25313
rect 27714 25241 27760 25279
rect 27714 25207 27720 25241
rect 27754 25207 27760 25241
rect 27714 25169 27760 25207
rect 27714 25135 27720 25169
rect 27754 25135 27760 25169
rect 27714 25112 27760 25135
rect 28172 25889 28218 25912
rect 28172 25855 28178 25889
rect 28212 25855 28218 25889
rect 28172 25817 28218 25855
rect 28172 25783 28178 25817
rect 28212 25783 28218 25817
rect 28172 25745 28218 25783
rect 28172 25711 28178 25745
rect 28212 25711 28218 25745
rect 28172 25673 28218 25711
rect 28172 25639 28178 25673
rect 28212 25639 28218 25673
rect 28172 25601 28218 25639
rect 28172 25567 28178 25601
rect 28212 25567 28218 25601
rect 28172 25529 28218 25567
rect 28172 25495 28178 25529
rect 28212 25495 28218 25529
rect 28172 25457 28218 25495
rect 28172 25423 28178 25457
rect 28212 25423 28218 25457
rect 28172 25385 28218 25423
rect 28172 25351 28178 25385
rect 28212 25351 28218 25385
rect 28172 25313 28218 25351
rect 28172 25279 28178 25313
rect 28212 25279 28218 25313
rect 28172 25241 28218 25279
rect 28172 25207 28178 25241
rect 28212 25207 28218 25241
rect 28172 25169 28218 25207
rect 28172 25135 28178 25169
rect 28212 25135 28218 25169
rect 28172 25112 28218 25135
rect 28630 25889 28676 25912
rect 28630 25855 28636 25889
rect 28670 25855 28676 25889
rect 28630 25817 28676 25855
rect 28630 25783 28636 25817
rect 28670 25783 28676 25817
rect 28630 25745 28676 25783
rect 28630 25711 28636 25745
rect 28670 25711 28676 25745
rect 28630 25673 28676 25711
rect 28630 25639 28636 25673
rect 28670 25639 28676 25673
rect 28630 25601 28676 25639
rect 28630 25567 28636 25601
rect 28670 25567 28676 25601
rect 28630 25529 28676 25567
rect 28630 25495 28636 25529
rect 28670 25495 28676 25529
rect 28630 25457 28676 25495
rect 28630 25423 28636 25457
rect 28670 25423 28676 25457
rect 28630 25385 28676 25423
rect 28630 25351 28636 25385
rect 28670 25351 28676 25385
rect 28630 25313 28676 25351
rect 28630 25279 28636 25313
rect 28670 25279 28676 25313
rect 28630 25241 28676 25279
rect 28630 25207 28636 25241
rect 28670 25207 28676 25241
rect 28630 25169 28676 25207
rect 28630 25135 28636 25169
rect 28670 25135 28676 25169
rect 28630 25112 28676 25135
rect 29088 25889 29134 25912
rect 29088 25855 29094 25889
rect 29128 25855 29134 25889
rect 29088 25817 29134 25855
rect 29088 25783 29094 25817
rect 29128 25783 29134 25817
rect 29088 25752 29134 25783
rect 29546 25889 29592 25912
rect 29546 25855 29552 25889
rect 29586 25855 29592 25889
rect 29546 25817 29592 25855
rect 29546 25783 29552 25817
rect 29586 25783 29592 25817
rect 29454 25752 29460 25764
rect 29088 25745 29460 25752
rect 29088 25711 29094 25745
rect 29128 25724 29460 25745
rect 29128 25711 29134 25724
rect 29454 25712 29460 25724
rect 29512 25712 29518 25764
rect 29546 25745 29592 25783
rect 29088 25673 29134 25711
rect 29088 25639 29094 25673
rect 29128 25639 29134 25673
rect 29088 25601 29134 25639
rect 29088 25567 29094 25601
rect 29128 25567 29134 25601
rect 29088 25529 29134 25567
rect 29088 25495 29094 25529
rect 29128 25495 29134 25529
rect 29088 25457 29134 25495
rect 29088 25423 29094 25457
rect 29128 25423 29134 25457
rect 29088 25385 29134 25423
rect 29088 25351 29094 25385
rect 29128 25351 29134 25385
rect 29088 25313 29134 25351
rect 29088 25279 29094 25313
rect 29128 25279 29134 25313
rect 29088 25241 29134 25279
rect 29088 25207 29094 25241
rect 29128 25207 29134 25241
rect 29088 25169 29134 25207
rect 29088 25135 29094 25169
rect 29128 25135 29134 25169
rect 29088 25112 29134 25135
rect 29546 25711 29552 25745
rect 29586 25711 29592 25745
rect 29546 25673 29592 25711
rect 29546 25639 29552 25673
rect 29586 25639 29592 25673
rect 29546 25601 29592 25639
rect 29546 25567 29552 25601
rect 29586 25567 29592 25601
rect 37405 25603 37413 26141
rect 37807 25603 37815 26141
rect 37405 25591 37815 25603
rect 39413 26141 39823 26153
rect 39413 25603 39420 26141
rect 39814 25603 39823 26141
rect 40149 26141 40559 26153
rect 40149 25628 40157 26141
rect 39413 25591 39823 25603
rect 29546 25529 29592 25567
rect 29546 25495 29552 25529
rect 29586 25495 29592 25529
rect 29546 25457 29592 25495
rect 29546 25423 29552 25457
rect 29586 25423 29592 25457
rect 29546 25385 29592 25423
rect 29546 25351 29552 25385
rect 29586 25351 29592 25385
rect 29546 25313 29592 25351
rect 29546 25279 29552 25313
rect 29586 25279 29592 25313
rect 29546 25241 29592 25279
rect 29546 25207 29552 25241
rect 29586 25207 29592 25241
rect 29546 25169 29592 25207
rect 29546 25135 29552 25169
rect 29586 25135 29592 25169
rect 29546 25112 29592 25135
rect 37405 25181 37815 25193
rect 24408 24627 24840 24643
rect 25884 24572 25912 25112
rect 27522 24868 27528 24880
rect 27467 24840 27528 24868
rect 27522 24828 27528 24840
rect 27580 24828 27586 24880
rect 37405 24676 37413 25181
rect 37366 24624 37372 24676
rect 37807 24643 37815 25181
rect 37424 24631 37815 24643
rect 39402 25181 39834 25591
rect 40126 25576 40132 25628
rect 40551 25603 40559 26141
rect 41414 26120 41420 26172
rect 41472 26120 41478 26172
rect 45664 26153 45692 26200
rect 46014 26188 46020 26240
rect 46072 26228 46078 26240
rect 48498 26228 48504 26240
rect 46072 26200 48504 26228
rect 46072 26188 46078 26200
rect 48498 26188 48504 26200
rect 48556 26188 48562 26240
rect 42157 26141 42567 26153
rect 40184 25591 40559 25603
rect 42157 25603 42164 26141
rect 42558 25603 42567 26141
rect 42893 26141 43303 26153
rect 42702 25644 42708 25696
rect 42760 25684 42766 25696
rect 42893 25684 42901 26141
rect 42760 25656 42901 25684
rect 42760 25644 42766 25656
rect 42157 25591 42567 25603
rect 42893 25603 42901 25656
rect 43295 25603 43303 26141
rect 42893 25591 43303 25603
rect 44901 26141 45311 26153
rect 44901 25603 44908 26141
rect 45302 25603 45311 26141
rect 44901 25591 45311 25603
rect 45637 26141 46047 26153
rect 45637 25603 45645 26141
rect 46039 25603 46047 26141
rect 45637 25591 46047 25603
rect 47645 26141 48055 26153
rect 47645 25603 47652 26141
rect 48046 25603 48055 26141
rect 47645 25591 48055 25603
rect 48381 26141 48791 26153
rect 48381 25603 48389 26141
rect 48783 25603 48791 26141
rect 48381 25591 48596 25603
rect 40184 25576 40190 25591
rect 39402 24643 39420 25181
rect 39814 24643 39834 25181
rect 40149 25181 40559 25193
rect 39942 25100 39948 25152
rect 40000 25140 40006 25152
rect 40149 25140 40157 25181
rect 40000 25112 40157 25140
rect 40000 25100 40006 25112
rect 37424 24624 37430 24631
rect 39402 24627 39834 24643
rect 40149 24643 40157 25112
rect 40551 24643 40559 25181
rect 40149 24631 40559 24643
rect 42146 25181 42578 25591
rect 42146 24643 42164 25181
rect 42558 24643 42578 25181
rect 42893 25181 43303 25193
rect 42893 24676 42901 25181
rect 42146 24627 42578 24643
rect 42886 24624 42892 24676
rect 43295 24643 43303 25181
rect 42944 24631 43303 24643
rect 44890 25181 45322 25591
rect 44890 24643 44908 25181
rect 45302 24643 45322 25181
rect 42944 24624 42950 24631
rect 44890 24627 45322 24643
rect 45637 25181 46047 25193
rect 45637 24643 45645 25181
rect 46039 25152 46047 25181
rect 47634 25181 48066 25591
rect 48590 25576 48596 25591
rect 48648 25591 48791 25603
rect 50389 26141 50799 26153
rect 50389 25603 50396 26141
rect 50790 25603 50799 26141
rect 50389 25591 50799 25603
rect 48648 25576 48654 25591
rect 46072 25100 46078 25152
rect 46039 24643 46047 25100
rect 45637 24631 46047 24643
rect 47634 24643 47652 25181
rect 48046 24643 48066 25181
rect 47634 24627 48066 24643
rect 48381 25181 48791 25193
rect 48381 24643 48389 25181
rect 48783 24643 48791 25181
rect 48381 24631 48791 24643
rect 50378 25181 50810 25591
rect 50378 24643 50396 25181
rect 50790 24643 50810 25181
rect 50378 24627 50810 24643
rect 900 24570 57536 24572
rect 900 24454 922 24570
rect 2510 24529 55926 24570
rect 2510 24495 22583 24529
rect 22617 24495 22783 24529
rect 22817 24495 22983 24529
rect 23017 24495 23183 24529
rect 23217 24495 23383 24529
rect 23417 24495 23583 24529
rect 23617 24495 23783 24529
rect 23817 24495 23983 24529
rect 24017 24495 24183 24529
rect 24217 24495 24383 24529
rect 24417 24495 24583 24529
rect 24617 24495 25601 24529
rect 25635 24495 26001 24529
rect 26035 24495 26401 24529
rect 26435 24495 26801 24529
rect 26835 24495 27201 24529
rect 27235 24495 27601 24529
rect 27635 24495 28001 24529
rect 28035 24495 28401 24529
rect 28435 24495 28801 24529
rect 28835 24495 29201 24529
rect 29235 24495 30111 24529
rect 30145 24495 30511 24529
rect 30545 24495 30911 24529
rect 30945 24495 31311 24529
rect 31345 24495 31711 24529
rect 31745 24495 32111 24529
rect 32145 24495 32511 24529
rect 32545 24495 32911 24529
rect 32945 24495 33311 24529
rect 33345 24495 33711 24529
rect 33745 24495 34111 24529
rect 34145 24495 34511 24529
rect 34545 24495 34911 24529
rect 34945 24495 35311 24529
rect 35345 24495 35711 24529
rect 35745 24495 36111 24529
rect 36145 24495 36511 24529
rect 36545 24495 36911 24529
rect 36945 24495 37577 24529
rect 37611 24495 37777 24529
rect 37811 24495 37977 24529
rect 38011 24495 38177 24529
rect 38211 24495 38377 24529
rect 38411 24495 38577 24529
rect 38611 24495 38777 24529
rect 38811 24495 38977 24529
rect 39011 24495 39177 24529
rect 39211 24495 39377 24529
rect 39411 24495 39577 24529
rect 39611 24495 40321 24529
rect 40355 24495 40521 24529
rect 40555 24495 40721 24529
rect 40755 24495 40921 24529
rect 40955 24495 41121 24529
rect 41155 24495 41321 24529
rect 41355 24495 41521 24529
rect 41555 24495 41721 24529
rect 41755 24495 41921 24529
rect 41955 24495 42121 24529
rect 42155 24495 42321 24529
rect 42355 24495 43065 24529
rect 43099 24495 43265 24529
rect 43299 24495 43465 24529
rect 43499 24495 43665 24529
rect 43699 24495 43865 24529
rect 43899 24495 44065 24529
rect 44099 24495 44265 24529
rect 44299 24495 44465 24529
rect 44499 24495 44665 24529
rect 44699 24495 44865 24529
rect 44899 24495 45065 24529
rect 45099 24495 45809 24529
rect 45843 24495 46009 24529
rect 46043 24495 46209 24529
rect 46243 24495 46409 24529
rect 46443 24495 46609 24529
rect 46643 24495 46809 24529
rect 46843 24495 47009 24529
rect 47043 24495 47209 24529
rect 47243 24495 47409 24529
rect 47443 24495 47609 24529
rect 47643 24495 47809 24529
rect 47843 24495 48553 24529
rect 48587 24495 48753 24529
rect 48787 24495 48953 24529
rect 48987 24495 49153 24529
rect 49187 24495 49353 24529
rect 49387 24495 49553 24529
rect 49587 24495 49753 24529
rect 49787 24495 49953 24529
rect 49987 24495 50153 24529
rect 50187 24495 50353 24529
rect 50387 24495 50553 24529
rect 50587 24495 55926 24529
rect 2510 24454 55926 24495
rect 57514 24454 57536 24570
rect 900 24452 57536 24454
rect 38286 24148 38292 24200
rect 38344 24188 38350 24200
rect 42886 24188 42892 24200
rect 38344 24160 42892 24188
rect 38344 24148 38350 24160
rect 42886 24148 42892 24160
rect 42944 24148 42950 24200
rect 30926 23400 30932 23452
rect 30984 23440 30990 23452
rect 37366 23440 37372 23452
rect 30984 23412 37372 23440
rect 30984 23400 30990 23412
rect 37366 23400 37372 23412
rect 37424 23400 37430 23452
rect 3348 22690 55088 22692
rect 3348 22574 3370 22690
rect 4958 22649 53478 22690
rect 4958 22615 24053 22649
rect 24087 22615 24253 22649
rect 24287 22615 24453 22649
rect 24487 22615 24653 22649
rect 24687 22615 24853 22649
rect 24887 22615 25053 22649
rect 25087 22615 25253 22649
rect 25287 22615 25453 22649
rect 25487 22615 25653 22649
rect 25687 22615 25853 22649
rect 25887 22615 26053 22649
rect 26087 22615 27385 22649
rect 27419 22615 27585 22649
rect 27619 22615 27785 22649
rect 27819 22615 27985 22649
rect 28019 22615 28185 22649
rect 28219 22615 28385 22649
rect 28419 22615 28585 22649
rect 28619 22615 28785 22649
rect 28819 22615 28985 22649
rect 29019 22615 29185 22649
rect 29219 22615 29385 22649
rect 29419 22615 30129 22649
rect 30163 22615 30329 22649
rect 30363 22615 30529 22649
rect 30563 22615 30729 22649
rect 30763 22615 30929 22649
rect 30963 22615 31129 22649
rect 31163 22615 31329 22649
rect 31363 22615 31529 22649
rect 31563 22615 31729 22649
rect 31763 22615 31929 22649
rect 31963 22615 32129 22649
rect 32163 22615 33363 22649
rect 33397 22615 33563 22649
rect 33597 22615 33763 22649
rect 33797 22615 33963 22649
rect 33997 22615 34163 22649
rect 34197 22615 34363 22649
rect 34397 22615 34563 22649
rect 34597 22615 34763 22649
rect 34797 22615 34963 22649
rect 34997 22615 35163 22649
rect 35197 22615 35363 22649
rect 35397 22615 37577 22649
rect 37611 22615 37777 22649
rect 37811 22615 37977 22649
rect 38011 22615 38177 22649
rect 38211 22615 38377 22649
rect 38411 22615 38577 22649
rect 38611 22615 38777 22649
rect 38811 22615 38977 22649
rect 39011 22615 39177 22649
rect 39211 22615 39377 22649
rect 39411 22615 39577 22649
rect 39611 22615 40321 22649
rect 40355 22615 40521 22649
rect 40555 22615 40721 22649
rect 40755 22615 40921 22649
rect 40955 22615 41121 22649
rect 41155 22615 41321 22649
rect 41355 22615 41521 22649
rect 41555 22615 41721 22649
rect 41755 22615 41921 22649
rect 41955 22615 42121 22649
rect 42155 22615 42321 22649
rect 42355 22615 48553 22649
rect 48587 22615 48753 22649
rect 48787 22615 48953 22649
rect 48987 22615 49153 22649
rect 49187 22615 49353 22649
rect 49387 22615 49553 22649
rect 49587 22615 49753 22649
rect 49787 22615 49953 22649
rect 49987 22615 50153 22649
rect 50187 22615 50353 22649
rect 50387 22615 50553 22649
rect 50587 22615 53478 22649
rect 4958 22574 53478 22615
rect 55066 22574 55088 22690
rect 3348 22572 55088 22574
rect 34974 22448 34980 22500
rect 35032 22488 35038 22500
rect 40126 22488 40132 22500
rect 35032 22460 40132 22488
rect 35032 22448 35038 22460
rect 40126 22448 40132 22460
rect 40184 22448 40190 22500
rect 42702 22488 42708 22500
rect 40512 22460 42708 22488
rect 40512 22393 40540 22460
rect 42702 22448 42708 22460
rect 42760 22448 42766 22500
rect 48498 22448 48504 22500
rect 48556 22448 48562 22500
rect 48516 22393 48544 22448
rect 23881 22381 24291 22393
rect 22922 22312 22928 22364
rect 22980 22352 22986 22364
rect 23881 22352 23889 22381
rect 22980 22324 23889 22352
rect 22980 22312 22986 22324
rect 23881 21843 23889 22324
rect 24283 21843 24291 22381
rect 23881 21831 24291 21843
rect 25889 22381 26299 22393
rect 25889 21843 25896 22381
rect 26290 21843 26299 22381
rect 25889 21831 26299 21843
rect 27213 22381 27623 22393
rect 27213 21843 27221 22381
rect 27615 21876 27623 22381
rect 29221 22381 29631 22393
rect 29086 21876 29092 21888
rect 27615 21848 29092 21876
rect 27615 21843 27623 21848
rect 27213 21831 27623 21843
rect 29086 21836 29092 21848
rect 29144 21836 29150 21888
rect 29221 21843 29228 22381
rect 29622 21843 29631 22381
rect 29221 21831 29631 21843
rect 29957 22381 30367 22393
rect 29957 21843 29965 22381
rect 30359 22352 30367 22381
rect 31965 22381 32375 22393
rect 30926 22352 30932 22364
rect 30359 22324 30932 22352
rect 30359 21843 30367 22324
rect 30926 22312 30932 22324
rect 30984 22312 30990 22364
rect 29957 21831 30367 21843
rect 31965 21843 31972 22381
rect 32366 21843 32375 22381
rect 31965 21831 32375 21843
rect 33191 22381 33601 22393
rect 33191 21843 33199 22381
rect 33593 21876 33601 22381
rect 35199 22381 35609 22393
rect 35066 21876 35072 21888
rect 33593 21848 35072 21876
rect 33593 21843 33601 21848
rect 33191 21831 33601 21843
rect 35066 21836 35072 21848
rect 35124 21836 35130 21888
rect 35199 21843 35206 22381
rect 35600 21843 35609 22381
rect 35199 21831 35609 21843
rect 37405 22381 37815 22393
rect 37405 21843 37413 22381
rect 37807 22352 37815 22381
rect 39413 22381 39823 22393
rect 38286 22352 38292 22364
rect 37807 22324 38292 22352
rect 37807 21843 37815 22324
rect 38286 22312 38292 22324
rect 38344 22312 38350 22364
rect 37405 21831 37815 21843
rect 39413 21843 39420 22381
rect 39814 21843 39823 22381
rect 39413 21831 39823 21843
rect 40149 22381 40559 22393
rect 40149 21843 40157 22381
rect 40551 21843 40559 22381
rect 40149 21831 40559 21843
rect 42157 22381 42567 22393
rect 42157 21843 42164 22381
rect 42558 21843 42567 22381
rect 42157 21831 42567 21843
rect 48381 22381 48791 22393
rect 48381 21843 48389 22381
rect 48783 21843 48791 22381
rect 48381 21831 48791 21843
rect 50389 22381 50799 22393
rect 50389 21843 50396 22381
rect 50790 21843 50799 22381
rect 50389 21831 50799 21843
rect 23881 21421 24291 21433
rect 16666 21360 16672 21412
rect 16724 21400 16730 21412
rect 23881 21400 23889 21421
rect 16724 21372 23889 21400
rect 16724 21360 16730 21372
rect 23881 20883 23889 21372
rect 24283 20883 24291 21421
rect 23881 20871 24291 20883
rect 25878 21421 26310 21831
rect 25878 20883 25896 21421
rect 26290 20883 26310 21421
rect 25878 20867 26310 20883
rect 27213 21421 27623 21433
rect 27213 20883 27221 21421
rect 27615 20883 27623 21421
rect 27213 20871 27623 20883
rect 29210 21421 29642 21831
rect 29210 20883 29228 21421
rect 29622 20883 29642 21421
rect 29957 21421 30367 21433
rect 29730 21360 29736 21412
rect 29788 21400 29794 21412
rect 29957 21400 29965 21421
rect 29788 21372 29965 21400
rect 29788 21360 29794 21372
rect 29210 20867 29642 20883
rect 29957 20883 29965 21372
rect 30359 20883 30367 21421
rect 29957 20871 30367 20883
rect 31954 21421 32386 21831
rect 31954 20883 31972 21421
rect 32366 20883 32386 21421
rect 31954 20867 32386 20883
rect 33191 21421 33601 21433
rect 33191 20883 33199 21421
rect 33593 21400 33601 21421
rect 35188 21421 35620 21831
rect 34974 21400 34980 21412
rect 33593 21372 34980 21400
rect 33593 20883 33601 21372
rect 34974 21360 34980 21372
rect 35032 21360 35038 21412
rect 33191 20871 33601 20883
rect 35188 20883 35206 21421
rect 35600 20883 35620 21421
rect 37405 21421 37815 21433
rect 35710 21360 35716 21412
rect 35768 21400 35774 21412
rect 37405 21400 37413 21421
rect 35768 21372 37413 21400
rect 35768 21360 35774 21372
rect 35188 20867 35620 20883
rect 37405 20883 37413 21372
rect 37807 20883 37815 21421
rect 37405 20871 37815 20883
rect 39402 21421 39834 21831
rect 39402 20883 39420 21421
rect 39814 20883 39834 21421
rect 39402 20867 39834 20883
rect 40149 21421 40559 21433
rect 40149 20883 40157 21421
rect 40551 21400 40559 21421
rect 42146 21421 42578 21831
rect 41414 21400 41420 21412
rect 40551 21372 41420 21400
rect 40551 20883 40559 21372
rect 41414 21360 41420 21372
rect 41472 21360 41478 21412
rect 40149 20871 40559 20883
rect 42146 20883 42164 21421
rect 42558 20883 42578 21421
rect 42146 20867 42578 20883
rect 48381 21421 48791 21433
rect 48381 20883 48389 21421
rect 48783 20883 48791 21421
rect 48381 20871 48791 20883
rect 50378 21421 50810 21831
rect 50378 20883 50396 21421
rect 50790 20883 50810 21421
rect 50378 20867 50810 20883
rect 900 20810 57536 20812
rect 900 20694 922 20810
rect 2510 20769 55926 20810
rect 2510 20735 24053 20769
rect 24087 20735 24253 20769
rect 24287 20735 24453 20769
rect 24487 20735 24653 20769
rect 24687 20735 24853 20769
rect 24887 20735 25053 20769
rect 25087 20735 25253 20769
rect 25287 20735 25453 20769
rect 25487 20735 25653 20769
rect 25687 20735 25853 20769
rect 25887 20735 26053 20769
rect 26087 20735 27385 20769
rect 27419 20735 27585 20769
rect 27619 20735 27785 20769
rect 27819 20735 27985 20769
rect 28019 20735 28185 20769
rect 28219 20735 28385 20769
rect 28419 20735 28585 20769
rect 28619 20735 28785 20769
rect 28819 20735 28985 20769
rect 29019 20735 29185 20769
rect 29219 20735 29385 20769
rect 29419 20735 30129 20769
rect 30163 20735 30329 20769
rect 30363 20735 30529 20769
rect 30563 20735 30729 20769
rect 30763 20735 30929 20769
rect 30963 20735 31129 20769
rect 31163 20735 31329 20769
rect 31363 20735 31529 20769
rect 31563 20735 31729 20769
rect 31763 20735 31929 20769
rect 31963 20735 32129 20769
rect 32163 20735 33363 20769
rect 33397 20735 33563 20769
rect 33597 20735 33763 20769
rect 33797 20735 33963 20769
rect 33997 20735 34163 20769
rect 34197 20735 34363 20769
rect 34397 20735 34563 20769
rect 34597 20735 34763 20769
rect 34797 20735 34963 20769
rect 34997 20735 35163 20769
rect 35197 20735 35363 20769
rect 35397 20735 37577 20769
rect 37611 20735 37777 20769
rect 37811 20735 37977 20769
rect 38011 20735 38177 20769
rect 38211 20735 38377 20769
rect 38411 20735 38577 20769
rect 38611 20735 38777 20769
rect 38811 20735 38977 20769
rect 39011 20735 39177 20769
rect 39211 20735 39377 20769
rect 39411 20735 39577 20769
rect 39611 20735 40321 20769
rect 40355 20735 40521 20769
rect 40555 20735 40721 20769
rect 40755 20735 40921 20769
rect 40955 20735 41121 20769
rect 41155 20735 41321 20769
rect 41355 20735 41521 20769
rect 41555 20735 41721 20769
rect 41755 20735 41921 20769
rect 41955 20735 42121 20769
rect 42155 20735 42321 20769
rect 42355 20735 48553 20769
rect 48587 20735 48753 20769
rect 48787 20735 48953 20769
rect 48987 20735 49153 20769
rect 49187 20735 49353 20769
rect 49387 20735 49553 20769
rect 49587 20735 49753 20769
rect 49787 20735 49953 20769
rect 49987 20735 50153 20769
rect 50187 20735 50353 20769
rect 50387 20735 50553 20769
rect 50587 20735 55926 20769
rect 2510 20694 55926 20735
rect 57514 20694 57536 20810
rect 900 20692 57536 20694
rect 3348 18930 55088 18932
rect 3348 18814 3370 18930
rect 4958 18889 53478 18930
rect 4958 18855 25013 18889
rect 25047 18855 25413 18889
rect 25447 18855 25813 18889
rect 25847 18855 26213 18889
rect 26247 18855 26613 18889
rect 26647 18855 27013 18889
rect 27047 18855 27413 18889
rect 27447 18855 27813 18889
rect 27847 18855 28213 18889
rect 28247 18855 28613 18889
rect 28647 18855 29013 18889
rect 29047 18855 29413 18889
rect 29447 18855 29813 18889
rect 29847 18855 30213 18889
rect 30247 18855 30613 18889
rect 30647 18855 31013 18889
rect 31047 18855 31413 18889
rect 31447 18855 31813 18889
rect 31847 18855 32213 18889
rect 32247 18855 32613 18889
rect 32647 18855 33013 18889
rect 33047 18855 33413 18889
rect 33447 18855 33813 18889
rect 33847 18855 34213 18889
rect 34247 18855 34613 18889
rect 34647 18855 35013 18889
rect 35047 18855 35413 18889
rect 35447 18855 35813 18889
rect 35847 18855 36213 18889
rect 36247 18855 36613 18889
rect 36647 18855 37013 18889
rect 37047 18855 37413 18889
rect 37447 18855 37813 18889
rect 37847 18855 38213 18889
rect 38247 18855 38613 18889
rect 38647 18855 39013 18889
rect 39047 18855 39413 18889
rect 39447 18855 39813 18889
rect 39847 18855 40213 18889
rect 40247 18855 40613 18889
rect 40647 18855 41013 18889
rect 41047 18855 41413 18889
rect 41447 18855 41813 18889
rect 41847 18855 42213 18889
rect 42247 18855 42613 18889
rect 42647 18855 43013 18889
rect 43047 18855 43413 18889
rect 43447 18855 43813 18889
rect 43847 18855 44213 18889
rect 44247 18855 44613 18889
rect 44647 18855 45013 18889
rect 45047 18855 45413 18889
rect 45447 18855 45813 18889
rect 45847 18855 46213 18889
rect 46247 18855 46613 18889
rect 46647 18855 47013 18889
rect 47047 18855 47413 18889
rect 47447 18855 47813 18889
rect 47847 18855 48213 18889
rect 48247 18855 48613 18889
rect 48647 18855 49013 18889
rect 49047 18855 49413 18889
rect 49447 18855 49813 18889
rect 49847 18855 50213 18889
rect 50247 18855 50613 18889
rect 50647 18855 51013 18889
rect 51047 18855 51413 18889
rect 51447 18855 51813 18889
rect 51847 18855 52213 18889
rect 52247 18855 53478 18889
rect 4958 18814 53478 18855
rect 55066 18814 55088 18930
rect 3348 18812 55088 18814
rect 25332 18637 25360 18812
rect 24871 18621 24917 18637
rect 24871 18587 24877 18621
rect 24911 18587 24917 18621
rect 24871 18549 24917 18587
rect 24871 18515 24877 18549
rect 24911 18515 24917 18549
rect 24871 18477 24917 18515
rect 24871 18443 24877 18477
rect 24911 18443 24917 18477
rect 24871 18405 24917 18443
rect 24871 18371 24877 18405
rect 24911 18371 24917 18405
rect 24871 18333 24917 18371
rect 24871 18299 24877 18333
rect 24911 18299 24917 18333
rect 24871 18261 24917 18299
rect 24871 18227 24877 18261
rect 24911 18227 24917 18261
rect 24871 18189 24917 18227
rect 24871 18155 24877 18189
rect 24911 18155 24917 18189
rect 24871 18117 24917 18155
rect 24871 18083 24877 18117
rect 24911 18083 24917 18117
rect 24871 18045 24917 18083
rect 24871 18011 24877 18045
rect 24911 18011 24917 18045
rect 24871 17973 24917 18011
rect 24871 17939 24877 17973
rect 24911 17939 24917 17973
rect 24871 17901 24917 17939
rect 24871 17867 24877 17901
rect 24911 17867 24917 17901
rect 24871 17829 24917 17867
rect 24871 17795 24877 17829
rect 24911 17795 24917 17829
rect 24871 17757 24917 17795
rect 24871 17723 24877 17757
rect 24911 17723 24917 17757
rect 24871 17685 24917 17723
rect 24871 17651 24877 17685
rect 24911 17651 24917 17685
rect 24871 17613 24917 17651
rect 24871 17579 24877 17613
rect 24911 17579 24917 17613
rect 24871 17541 24917 17579
rect 24871 17507 24877 17541
rect 24911 17507 24917 17541
rect 24871 17469 24917 17507
rect 24871 17435 24877 17469
rect 24911 17435 24917 17469
rect 24871 17397 24917 17435
rect 24871 17363 24877 17397
rect 24911 17363 24917 17397
rect 24871 17347 24917 17363
rect 25329 18621 25375 18637
rect 25329 18587 25335 18621
rect 25369 18587 25375 18621
rect 25329 18549 25375 18587
rect 25329 18515 25335 18549
rect 25369 18515 25375 18549
rect 25329 18477 25375 18515
rect 25329 18443 25335 18477
rect 25369 18443 25375 18477
rect 25329 18405 25375 18443
rect 25329 18371 25335 18405
rect 25369 18371 25375 18405
rect 25329 18333 25375 18371
rect 25329 18299 25335 18333
rect 25369 18299 25375 18333
rect 25329 18261 25375 18299
rect 25329 18227 25335 18261
rect 25369 18227 25375 18261
rect 25329 18189 25375 18227
rect 25329 18155 25335 18189
rect 25369 18155 25375 18189
rect 25329 18117 25375 18155
rect 25329 18083 25335 18117
rect 25369 18083 25375 18117
rect 25329 18045 25375 18083
rect 25329 18011 25335 18045
rect 25369 18011 25375 18045
rect 25329 17973 25375 18011
rect 25329 17939 25335 17973
rect 25369 17939 25375 17973
rect 25329 17901 25375 17939
rect 25329 17867 25335 17901
rect 25369 17867 25375 17901
rect 25329 17829 25375 17867
rect 25329 17795 25335 17829
rect 25369 17795 25375 17829
rect 25329 17757 25375 17795
rect 25329 17723 25335 17757
rect 25369 17723 25375 17757
rect 25329 17685 25375 17723
rect 25329 17651 25335 17685
rect 25369 17651 25375 17685
rect 25329 17613 25375 17651
rect 25329 17579 25335 17613
rect 25369 17579 25375 17613
rect 25329 17541 25375 17579
rect 25329 17507 25335 17541
rect 25369 17507 25375 17541
rect 25329 17469 25375 17507
rect 25329 17435 25335 17469
rect 25369 17435 25375 17469
rect 25329 17397 25375 17435
rect 25329 17363 25335 17397
rect 25369 17363 25375 17397
rect 25329 17347 25375 17363
rect 25787 18621 25833 18637
rect 25787 18587 25793 18621
rect 25827 18587 25833 18621
rect 25787 18549 25833 18587
rect 25787 18515 25793 18549
rect 25827 18515 25833 18549
rect 25787 18477 25833 18515
rect 25787 18443 25793 18477
rect 25827 18443 25833 18477
rect 25787 18405 25833 18443
rect 25787 18371 25793 18405
rect 25827 18371 25833 18405
rect 25787 18333 25833 18371
rect 25787 18299 25793 18333
rect 25827 18299 25833 18333
rect 25787 18261 25833 18299
rect 25787 18227 25793 18261
rect 25827 18227 25833 18261
rect 25787 18189 25833 18227
rect 25787 18155 25793 18189
rect 25827 18155 25833 18189
rect 25787 18117 25833 18155
rect 25787 18083 25793 18117
rect 25827 18083 25833 18117
rect 25787 18045 25833 18083
rect 25787 18011 25793 18045
rect 25827 18011 25833 18045
rect 25787 17973 25833 18011
rect 25787 17939 25793 17973
rect 25827 17939 25833 17973
rect 25787 17901 25833 17939
rect 25787 17867 25793 17901
rect 25827 17867 25833 17901
rect 25787 17829 25833 17867
rect 25787 17795 25793 17829
rect 25827 17795 25833 17829
rect 25787 17757 25833 17795
rect 25787 17723 25793 17757
rect 25827 17723 25833 17757
rect 25787 17685 25833 17723
rect 25787 17651 25793 17685
rect 25827 17651 25833 17685
rect 25787 17613 25833 17651
rect 25787 17579 25793 17613
rect 25827 17579 25833 17613
rect 25787 17541 25833 17579
rect 25787 17507 25793 17541
rect 25827 17507 25833 17541
rect 25787 17469 25833 17507
rect 25787 17435 25793 17469
rect 25827 17435 25833 17469
rect 25787 17397 25833 17435
rect 25787 17363 25793 17397
rect 25827 17363 25833 17397
rect 25787 17347 25833 17363
rect 26245 18621 26291 18637
rect 26245 18587 26251 18621
rect 26285 18587 26291 18621
rect 26245 18549 26291 18587
rect 26245 18515 26251 18549
rect 26285 18515 26291 18549
rect 26245 18477 26291 18515
rect 26245 18443 26251 18477
rect 26285 18443 26291 18477
rect 26245 18405 26291 18443
rect 26245 18371 26251 18405
rect 26285 18371 26291 18405
rect 26245 18333 26291 18371
rect 26245 18299 26251 18333
rect 26285 18299 26291 18333
rect 26245 18261 26291 18299
rect 26245 18227 26251 18261
rect 26285 18227 26291 18261
rect 26245 18189 26291 18227
rect 26245 18155 26251 18189
rect 26285 18155 26291 18189
rect 26245 18117 26291 18155
rect 26245 18083 26251 18117
rect 26285 18083 26291 18117
rect 26245 18045 26291 18083
rect 26245 18011 26251 18045
rect 26285 18011 26291 18045
rect 26245 17973 26291 18011
rect 26245 17939 26251 17973
rect 26285 17939 26291 17973
rect 26245 17901 26291 17939
rect 26245 17867 26251 17901
rect 26285 17867 26291 17901
rect 26245 17829 26291 17867
rect 26245 17795 26251 17829
rect 26285 17795 26291 17829
rect 26245 17757 26291 17795
rect 26245 17723 26251 17757
rect 26285 17723 26291 17757
rect 26245 17685 26291 17723
rect 26245 17651 26251 17685
rect 26285 17651 26291 17685
rect 26245 17613 26291 17651
rect 26245 17579 26251 17613
rect 26285 17579 26291 17613
rect 26245 17541 26291 17579
rect 26245 17507 26251 17541
rect 26285 17507 26291 17541
rect 26245 17469 26291 17507
rect 26245 17435 26251 17469
rect 26285 17435 26291 17469
rect 26245 17397 26291 17435
rect 26245 17363 26251 17397
rect 26285 17363 26291 17397
rect 26245 17347 26291 17363
rect 26703 18621 26749 18637
rect 26703 18587 26709 18621
rect 26743 18587 26749 18621
rect 26703 18549 26749 18587
rect 26703 18515 26709 18549
rect 26743 18515 26749 18549
rect 26703 18477 26749 18515
rect 26703 18443 26709 18477
rect 26743 18443 26749 18477
rect 26703 18405 26749 18443
rect 26703 18371 26709 18405
rect 26743 18371 26749 18405
rect 26703 18333 26749 18371
rect 26703 18299 26709 18333
rect 26743 18299 26749 18333
rect 26703 18261 26749 18299
rect 26703 18227 26709 18261
rect 26743 18227 26749 18261
rect 26703 18189 26749 18227
rect 26703 18155 26709 18189
rect 26743 18155 26749 18189
rect 26703 18117 26749 18155
rect 26703 18083 26709 18117
rect 26743 18083 26749 18117
rect 26703 18045 26749 18083
rect 26703 18011 26709 18045
rect 26743 18011 26749 18045
rect 26703 17973 26749 18011
rect 26703 17939 26709 17973
rect 26743 17939 26749 17973
rect 26703 17901 26749 17939
rect 26703 17867 26709 17901
rect 26743 17867 26749 17901
rect 26703 17829 26749 17867
rect 26703 17795 26709 17829
rect 26743 17795 26749 17829
rect 26703 17757 26749 17795
rect 26703 17723 26709 17757
rect 26743 17723 26749 17757
rect 26703 17685 26749 17723
rect 26703 17651 26709 17685
rect 26743 17651 26749 17685
rect 26703 17613 26749 17651
rect 26703 17579 26709 17613
rect 26743 17579 26749 17613
rect 26703 17541 26749 17579
rect 26703 17507 26709 17541
rect 26743 17507 26749 17541
rect 26703 17469 26749 17507
rect 26703 17435 26709 17469
rect 26743 17435 26749 17469
rect 26703 17397 26749 17435
rect 26703 17363 26709 17397
rect 26743 17363 26749 17397
rect 26703 17347 26749 17363
rect 27161 18621 27207 18637
rect 27161 18587 27167 18621
rect 27201 18587 27207 18621
rect 27161 18549 27207 18587
rect 27161 18515 27167 18549
rect 27201 18515 27207 18549
rect 27161 18477 27207 18515
rect 27161 18443 27167 18477
rect 27201 18443 27207 18477
rect 27161 18405 27207 18443
rect 27161 18371 27167 18405
rect 27201 18371 27207 18405
rect 27161 18333 27207 18371
rect 27161 18299 27167 18333
rect 27201 18299 27207 18333
rect 27161 18261 27207 18299
rect 27161 18227 27167 18261
rect 27201 18227 27207 18261
rect 27161 18189 27207 18227
rect 27161 18155 27167 18189
rect 27201 18155 27207 18189
rect 27161 18117 27207 18155
rect 27161 18083 27167 18117
rect 27201 18083 27207 18117
rect 27161 18045 27207 18083
rect 27161 18011 27167 18045
rect 27201 18011 27207 18045
rect 27161 17973 27207 18011
rect 27161 17939 27167 17973
rect 27201 17939 27207 17973
rect 27161 17901 27207 17939
rect 27161 17867 27167 17901
rect 27201 17867 27207 17901
rect 27161 17829 27207 17867
rect 27161 17795 27167 17829
rect 27201 17795 27207 17829
rect 27161 17757 27207 17795
rect 27161 17723 27167 17757
rect 27201 17723 27207 17757
rect 27161 17685 27207 17723
rect 27161 17651 27167 17685
rect 27201 17651 27207 17685
rect 27161 17613 27207 17651
rect 27161 17579 27167 17613
rect 27201 17579 27207 17613
rect 27161 17541 27207 17579
rect 27161 17507 27167 17541
rect 27201 17507 27207 17541
rect 27161 17469 27207 17507
rect 27161 17435 27167 17469
rect 27201 17435 27207 17469
rect 27161 17397 27207 17435
rect 27161 17363 27167 17397
rect 27201 17363 27207 17397
rect 27161 17347 27207 17363
rect 27619 18621 27665 18637
rect 27619 18587 27625 18621
rect 27659 18587 27665 18621
rect 27619 18549 27665 18587
rect 27619 18515 27625 18549
rect 27659 18515 27665 18549
rect 27619 18477 27665 18515
rect 27619 18443 27625 18477
rect 27659 18443 27665 18477
rect 27619 18405 27665 18443
rect 27619 18371 27625 18405
rect 27659 18371 27665 18405
rect 27619 18333 27665 18371
rect 27619 18299 27625 18333
rect 27659 18299 27665 18333
rect 27619 18261 27665 18299
rect 27619 18227 27625 18261
rect 27659 18227 27665 18261
rect 27619 18189 27665 18227
rect 27619 18155 27625 18189
rect 27659 18155 27665 18189
rect 27619 18117 27665 18155
rect 27619 18083 27625 18117
rect 27659 18083 27665 18117
rect 27619 18045 27665 18083
rect 27619 18011 27625 18045
rect 27659 18011 27665 18045
rect 27619 17973 27665 18011
rect 27619 17939 27625 17973
rect 27659 17939 27665 17973
rect 27619 17901 27665 17939
rect 27619 17867 27625 17901
rect 27659 17867 27665 17901
rect 27619 17829 27665 17867
rect 27619 17795 27625 17829
rect 27659 17795 27665 17829
rect 27619 17757 27665 17795
rect 27619 17723 27625 17757
rect 27659 17723 27665 17757
rect 27619 17685 27665 17723
rect 27619 17651 27625 17685
rect 27659 17651 27665 17685
rect 27619 17613 27665 17651
rect 27619 17579 27625 17613
rect 27659 17579 27665 17613
rect 27619 17541 27665 17579
rect 27619 17507 27625 17541
rect 27659 17507 27665 17541
rect 27619 17469 27665 17507
rect 27619 17435 27625 17469
rect 27659 17435 27665 17469
rect 27619 17397 27665 17435
rect 27619 17363 27625 17397
rect 27659 17363 27665 17397
rect 27619 17347 27665 17363
rect 28077 18621 28123 18637
rect 28077 18587 28083 18621
rect 28117 18587 28123 18621
rect 28077 18549 28123 18587
rect 28077 18515 28083 18549
rect 28117 18515 28123 18549
rect 28077 18477 28123 18515
rect 28077 18443 28083 18477
rect 28117 18443 28123 18477
rect 28077 18405 28123 18443
rect 28077 18371 28083 18405
rect 28117 18371 28123 18405
rect 28077 18333 28123 18371
rect 28077 18299 28083 18333
rect 28117 18299 28123 18333
rect 28077 18261 28123 18299
rect 28077 18227 28083 18261
rect 28117 18227 28123 18261
rect 28077 18189 28123 18227
rect 28077 18155 28083 18189
rect 28117 18155 28123 18189
rect 28077 18117 28123 18155
rect 28077 18083 28083 18117
rect 28117 18083 28123 18117
rect 28077 18045 28123 18083
rect 28077 18011 28083 18045
rect 28117 18011 28123 18045
rect 28077 17973 28123 18011
rect 28077 17939 28083 17973
rect 28117 17939 28123 17973
rect 28077 17901 28123 17939
rect 28077 17867 28083 17901
rect 28117 17867 28123 17901
rect 28077 17829 28123 17867
rect 28077 17795 28083 17829
rect 28117 17795 28123 17829
rect 28077 17757 28123 17795
rect 28077 17723 28083 17757
rect 28117 17723 28123 17757
rect 28077 17685 28123 17723
rect 28077 17651 28083 17685
rect 28117 17651 28123 17685
rect 28077 17613 28123 17651
rect 28077 17579 28083 17613
rect 28117 17579 28123 17613
rect 28077 17541 28123 17579
rect 28077 17507 28083 17541
rect 28117 17507 28123 17541
rect 28077 17469 28123 17507
rect 28077 17435 28083 17469
rect 28117 17435 28123 17469
rect 28077 17397 28123 17435
rect 28077 17363 28083 17397
rect 28117 17363 28123 17397
rect 28077 17347 28123 17363
rect 28535 18621 28581 18637
rect 28535 18587 28541 18621
rect 28575 18587 28581 18621
rect 28535 18549 28581 18587
rect 28535 18515 28541 18549
rect 28575 18515 28581 18549
rect 28535 18477 28581 18515
rect 28535 18443 28541 18477
rect 28575 18443 28581 18477
rect 28535 18405 28581 18443
rect 28535 18371 28541 18405
rect 28575 18371 28581 18405
rect 28535 18333 28581 18371
rect 28535 18299 28541 18333
rect 28575 18299 28581 18333
rect 28535 18261 28581 18299
rect 28535 18227 28541 18261
rect 28575 18227 28581 18261
rect 28535 18189 28581 18227
rect 28535 18155 28541 18189
rect 28575 18155 28581 18189
rect 28535 18117 28581 18155
rect 28535 18083 28541 18117
rect 28575 18083 28581 18117
rect 28535 18045 28581 18083
rect 28535 18011 28541 18045
rect 28575 18011 28581 18045
rect 28535 17973 28581 18011
rect 28535 17939 28541 17973
rect 28575 17939 28581 17973
rect 28535 17901 28581 17939
rect 28535 17867 28541 17901
rect 28575 17867 28581 17901
rect 28535 17829 28581 17867
rect 28535 17795 28541 17829
rect 28575 17795 28581 17829
rect 28535 17757 28581 17795
rect 28535 17723 28541 17757
rect 28575 17723 28581 17757
rect 28535 17685 28581 17723
rect 28535 17651 28541 17685
rect 28575 17651 28581 17685
rect 28535 17613 28581 17651
rect 28535 17579 28541 17613
rect 28575 17579 28581 17613
rect 28535 17541 28581 17579
rect 28535 17507 28541 17541
rect 28575 17507 28581 17541
rect 28535 17469 28581 17507
rect 28535 17435 28541 17469
rect 28575 17435 28581 17469
rect 28535 17397 28581 17435
rect 28535 17363 28541 17397
rect 28575 17363 28581 17397
rect 28535 17347 28581 17363
rect 28993 18621 29039 18637
rect 28993 18587 28999 18621
rect 29033 18587 29039 18621
rect 28993 18549 29039 18587
rect 28993 18515 28999 18549
rect 29033 18515 29039 18549
rect 28993 18477 29039 18515
rect 28993 18443 28999 18477
rect 29033 18443 29039 18477
rect 28993 18405 29039 18443
rect 28993 18371 28999 18405
rect 29033 18371 29039 18405
rect 28993 18333 29039 18371
rect 28993 18299 28999 18333
rect 29033 18299 29039 18333
rect 28993 18261 29039 18299
rect 28993 18227 28999 18261
rect 29033 18227 29039 18261
rect 28993 18189 29039 18227
rect 28993 18155 28999 18189
rect 29033 18155 29039 18189
rect 28993 18117 29039 18155
rect 28993 18083 28999 18117
rect 29033 18083 29039 18117
rect 28993 18045 29039 18083
rect 28993 18011 28999 18045
rect 29033 18011 29039 18045
rect 28993 17973 29039 18011
rect 28993 17939 28999 17973
rect 29033 17939 29039 17973
rect 28993 17901 29039 17939
rect 28993 17867 28999 17901
rect 29033 17867 29039 17901
rect 28993 17829 29039 17867
rect 28993 17795 28999 17829
rect 29033 17795 29039 17829
rect 28993 17757 29039 17795
rect 28993 17723 28999 17757
rect 29033 17723 29039 17757
rect 28993 17685 29039 17723
rect 28993 17651 28999 17685
rect 29033 17651 29039 17685
rect 28993 17613 29039 17651
rect 28993 17579 28999 17613
rect 29033 17579 29039 17613
rect 28993 17541 29039 17579
rect 28993 17507 28999 17541
rect 29033 17507 29039 17541
rect 28993 17469 29039 17507
rect 28993 17435 28999 17469
rect 29033 17435 29039 17469
rect 28993 17397 29039 17435
rect 28993 17363 28999 17397
rect 29033 17363 29039 17397
rect 28993 17347 29039 17363
rect 29451 18621 29497 18637
rect 29451 18587 29457 18621
rect 29491 18587 29497 18621
rect 29451 18549 29497 18587
rect 29451 18515 29457 18549
rect 29491 18515 29497 18549
rect 29451 18477 29497 18515
rect 29451 18443 29457 18477
rect 29491 18443 29497 18477
rect 29451 18405 29497 18443
rect 29451 18371 29457 18405
rect 29491 18371 29497 18405
rect 29451 18333 29497 18371
rect 29451 18299 29457 18333
rect 29491 18299 29497 18333
rect 29451 18261 29497 18299
rect 29451 18227 29457 18261
rect 29491 18227 29497 18261
rect 29451 18189 29497 18227
rect 29451 18155 29457 18189
rect 29491 18155 29497 18189
rect 29451 18117 29497 18155
rect 29451 18083 29457 18117
rect 29491 18083 29497 18117
rect 29451 18045 29497 18083
rect 29451 18011 29457 18045
rect 29491 18011 29497 18045
rect 29451 17973 29497 18011
rect 29451 17939 29457 17973
rect 29491 17939 29497 17973
rect 29451 17901 29497 17939
rect 29451 17867 29457 17901
rect 29491 17867 29497 17901
rect 29451 17829 29497 17867
rect 29451 17795 29457 17829
rect 29491 17795 29497 17829
rect 29451 17757 29497 17795
rect 29451 17723 29457 17757
rect 29491 17723 29497 17757
rect 29451 17685 29497 17723
rect 29451 17651 29457 17685
rect 29491 17651 29497 17685
rect 29451 17613 29497 17651
rect 29451 17579 29457 17613
rect 29491 17579 29497 17613
rect 29451 17541 29497 17579
rect 29451 17507 29457 17541
rect 29491 17507 29497 17541
rect 29451 17469 29497 17507
rect 29451 17435 29457 17469
rect 29491 17435 29497 17469
rect 29451 17397 29497 17435
rect 29451 17363 29457 17397
rect 29491 17363 29497 17397
rect 29451 17347 29497 17363
rect 29909 18621 29955 18637
rect 29909 18587 29915 18621
rect 29949 18587 29955 18621
rect 29909 18549 29955 18587
rect 29909 18515 29915 18549
rect 29949 18515 29955 18549
rect 29909 18477 29955 18515
rect 29909 18443 29915 18477
rect 29949 18443 29955 18477
rect 29909 18405 29955 18443
rect 29909 18371 29915 18405
rect 29949 18371 29955 18405
rect 29909 18333 29955 18371
rect 29909 18299 29915 18333
rect 29949 18299 29955 18333
rect 29909 18261 29955 18299
rect 29909 18227 29915 18261
rect 29949 18227 29955 18261
rect 29909 18189 29955 18227
rect 29909 18155 29915 18189
rect 29949 18155 29955 18189
rect 29909 18117 29955 18155
rect 29909 18083 29915 18117
rect 29949 18083 29955 18117
rect 29909 18045 29955 18083
rect 29909 18011 29915 18045
rect 29949 18011 29955 18045
rect 29909 17973 29955 18011
rect 29909 17939 29915 17973
rect 29949 17939 29955 17973
rect 29909 17901 29955 17939
rect 29909 17867 29915 17901
rect 29949 17867 29955 17901
rect 29909 17829 29955 17867
rect 29909 17795 29915 17829
rect 29949 17795 29955 17829
rect 29909 17757 29955 17795
rect 29909 17723 29915 17757
rect 29949 17723 29955 17757
rect 29909 17685 29955 17723
rect 29909 17651 29915 17685
rect 29949 17651 29955 17685
rect 29909 17613 29955 17651
rect 29909 17579 29915 17613
rect 29949 17579 29955 17613
rect 29909 17541 29955 17579
rect 29909 17507 29915 17541
rect 29949 17507 29955 17541
rect 29909 17469 29955 17507
rect 29909 17435 29915 17469
rect 29949 17435 29955 17469
rect 29909 17397 29955 17435
rect 29909 17363 29915 17397
rect 29949 17363 29955 17397
rect 29909 17347 29955 17363
rect 30367 18621 30413 18637
rect 30367 18587 30373 18621
rect 30407 18587 30413 18621
rect 30367 18549 30413 18587
rect 30367 18515 30373 18549
rect 30407 18515 30413 18549
rect 30367 18477 30413 18515
rect 30367 18443 30373 18477
rect 30407 18443 30413 18477
rect 30367 18405 30413 18443
rect 30367 18371 30373 18405
rect 30407 18371 30413 18405
rect 30367 18333 30413 18371
rect 30367 18299 30373 18333
rect 30407 18299 30413 18333
rect 30367 18261 30413 18299
rect 30367 18227 30373 18261
rect 30407 18227 30413 18261
rect 30367 18189 30413 18227
rect 30367 18155 30373 18189
rect 30407 18155 30413 18189
rect 30367 18117 30413 18155
rect 30367 18083 30373 18117
rect 30407 18083 30413 18117
rect 30367 18045 30413 18083
rect 30367 18011 30373 18045
rect 30407 18011 30413 18045
rect 30367 17973 30413 18011
rect 30367 17939 30373 17973
rect 30407 17939 30413 17973
rect 30367 17901 30413 17939
rect 30367 17867 30373 17901
rect 30407 17867 30413 17901
rect 30367 17829 30413 17867
rect 30367 17795 30373 17829
rect 30407 17795 30413 17829
rect 30367 17757 30413 17795
rect 30367 17723 30373 17757
rect 30407 17723 30413 17757
rect 30367 17685 30413 17723
rect 30367 17651 30373 17685
rect 30407 17651 30413 17685
rect 30367 17613 30413 17651
rect 30367 17579 30373 17613
rect 30407 17579 30413 17613
rect 30367 17541 30413 17579
rect 30367 17507 30373 17541
rect 30407 17507 30413 17541
rect 30367 17469 30413 17507
rect 30367 17435 30373 17469
rect 30407 17435 30413 17469
rect 30367 17397 30413 17435
rect 30367 17363 30373 17397
rect 30407 17363 30413 17397
rect 30367 17347 30413 17363
rect 30825 18621 30871 18637
rect 30825 18587 30831 18621
rect 30865 18587 30871 18621
rect 30825 18549 30871 18587
rect 30825 18515 30831 18549
rect 30865 18515 30871 18549
rect 30825 18477 30871 18515
rect 30825 18443 30831 18477
rect 30865 18443 30871 18477
rect 30825 18405 30871 18443
rect 30825 18371 30831 18405
rect 30865 18371 30871 18405
rect 30825 18333 30871 18371
rect 30825 18299 30831 18333
rect 30865 18299 30871 18333
rect 30825 18261 30871 18299
rect 30825 18227 30831 18261
rect 30865 18227 30871 18261
rect 30825 18189 30871 18227
rect 30825 18155 30831 18189
rect 30865 18155 30871 18189
rect 30825 18117 30871 18155
rect 30825 18083 30831 18117
rect 30865 18083 30871 18117
rect 30825 18045 30871 18083
rect 30825 18011 30831 18045
rect 30865 18011 30871 18045
rect 30825 17973 30871 18011
rect 30825 17939 30831 17973
rect 30865 17939 30871 17973
rect 30825 17901 30871 17939
rect 30825 17867 30831 17901
rect 30865 17867 30871 17901
rect 30825 17829 30871 17867
rect 30825 17795 30831 17829
rect 30865 17795 30871 17829
rect 30825 17757 30871 17795
rect 30825 17723 30831 17757
rect 30865 17723 30871 17757
rect 30825 17685 30871 17723
rect 30825 17651 30831 17685
rect 30865 17651 30871 17685
rect 30825 17613 30871 17651
rect 30825 17579 30831 17613
rect 30865 17579 30871 17613
rect 30825 17541 30871 17579
rect 30825 17507 30831 17541
rect 30865 17507 30871 17541
rect 30825 17469 30871 17507
rect 30825 17435 30831 17469
rect 30865 17435 30871 17469
rect 30825 17397 30871 17435
rect 30825 17363 30831 17397
rect 30865 17363 30871 17397
rect 30825 17347 30871 17363
rect 31283 18621 31329 18637
rect 31283 18587 31289 18621
rect 31323 18587 31329 18621
rect 31283 18549 31329 18587
rect 31283 18515 31289 18549
rect 31323 18515 31329 18549
rect 31283 18477 31329 18515
rect 31283 18443 31289 18477
rect 31323 18443 31329 18477
rect 31283 18405 31329 18443
rect 31283 18371 31289 18405
rect 31323 18371 31329 18405
rect 31283 18333 31329 18371
rect 31283 18299 31289 18333
rect 31323 18299 31329 18333
rect 31283 18261 31329 18299
rect 31283 18227 31289 18261
rect 31323 18227 31329 18261
rect 31283 18189 31329 18227
rect 31283 18155 31289 18189
rect 31323 18155 31329 18189
rect 31283 18117 31329 18155
rect 31283 18083 31289 18117
rect 31323 18083 31329 18117
rect 31283 18045 31329 18083
rect 31283 18011 31289 18045
rect 31323 18011 31329 18045
rect 31283 17973 31329 18011
rect 31283 17939 31289 17973
rect 31323 17939 31329 17973
rect 31283 17901 31329 17939
rect 31283 17867 31289 17901
rect 31323 17867 31329 17901
rect 31283 17829 31329 17867
rect 31283 17795 31289 17829
rect 31323 17795 31329 17829
rect 31283 17757 31329 17795
rect 31283 17723 31289 17757
rect 31323 17723 31329 17757
rect 31283 17685 31329 17723
rect 31283 17651 31289 17685
rect 31323 17651 31329 17685
rect 31283 17613 31329 17651
rect 31283 17579 31289 17613
rect 31323 17579 31329 17613
rect 31283 17541 31329 17579
rect 31283 17507 31289 17541
rect 31323 17507 31329 17541
rect 31283 17469 31329 17507
rect 31283 17435 31289 17469
rect 31323 17435 31329 17469
rect 31283 17397 31329 17435
rect 31283 17363 31289 17397
rect 31323 17363 31329 17397
rect 31283 17347 31329 17363
rect 31741 18621 31787 18637
rect 31741 18587 31747 18621
rect 31781 18587 31787 18621
rect 31741 18549 31787 18587
rect 31741 18515 31747 18549
rect 31781 18515 31787 18549
rect 31741 18477 31787 18515
rect 31741 18443 31747 18477
rect 31781 18443 31787 18477
rect 31741 18405 31787 18443
rect 31741 18371 31747 18405
rect 31781 18371 31787 18405
rect 31741 18333 31787 18371
rect 31741 18299 31747 18333
rect 31781 18299 31787 18333
rect 31741 18261 31787 18299
rect 31741 18227 31747 18261
rect 31781 18227 31787 18261
rect 31741 18189 31787 18227
rect 31741 18155 31747 18189
rect 31781 18155 31787 18189
rect 31741 18117 31787 18155
rect 31741 18083 31747 18117
rect 31781 18083 31787 18117
rect 31741 18045 31787 18083
rect 31741 18011 31747 18045
rect 31781 18011 31787 18045
rect 31741 17973 31787 18011
rect 31741 17939 31747 17973
rect 31781 17939 31787 17973
rect 31741 17901 31787 17939
rect 31741 17867 31747 17901
rect 31781 17867 31787 17901
rect 31741 17829 31787 17867
rect 31741 17795 31747 17829
rect 31781 17795 31787 17829
rect 31741 17757 31787 17795
rect 31741 17723 31747 17757
rect 31781 17723 31787 17757
rect 31741 17685 31787 17723
rect 31741 17651 31747 17685
rect 31781 17651 31787 17685
rect 31741 17613 31787 17651
rect 31741 17579 31747 17613
rect 31781 17579 31787 17613
rect 31741 17541 31787 17579
rect 31741 17507 31747 17541
rect 31781 17507 31787 17541
rect 31741 17469 31787 17507
rect 31741 17435 31747 17469
rect 31781 17435 31787 17469
rect 31741 17397 31787 17435
rect 31741 17363 31747 17397
rect 31781 17363 31787 17397
rect 31741 17347 31787 17363
rect 32199 18621 32245 18637
rect 32199 18587 32205 18621
rect 32239 18587 32245 18621
rect 32199 18549 32245 18587
rect 32199 18515 32205 18549
rect 32239 18515 32245 18549
rect 32199 18477 32245 18515
rect 32199 18443 32205 18477
rect 32239 18443 32245 18477
rect 32199 18405 32245 18443
rect 32199 18371 32205 18405
rect 32239 18371 32245 18405
rect 32199 18333 32245 18371
rect 32199 18299 32205 18333
rect 32239 18299 32245 18333
rect 32199 18261 32245 18299
rect 32199 18227 32205 18261
rect 32239 18227 32245 18261
rect 32199 18189 32245 18227
rect 32199 18155 32205 18189
rect 32239 18155 32245 18189
rect 32199 18117 32245 18155
rect 32199 18083 32205 18117
rect 32239 18083 32245 18117
rect 32199 18045 32245 18083
rect 32199 18011 32205 18045
rect 32239 18011 32245 18045
rect 32199 17973 32245 18011
rect 32199 17939 32205 17973
rect 32239 17939 32245 17973
rect 32199 17901 32245 17939
rect 32199 17867 32205 17901
rect 32239 17867 32245 17901
rect 32199 17829 32245 17867
rect 32199 17795 32205 17829
rect 32239 17795 32245 17829
rect 32199 17757 32245 17795
rect 32199 17723 32205 17757
rect 32239 17723 32245 17757
rect 32199 17685 32245 17723
rect 32199 17651 32205 17685
rect 32239 17651 32245 17685
rect 32199 17613 32245 17651
rect 32199 17579 32205 17613
rect 32239 17579 32245 17613
rect 32199 17541 32245 17579
rect 32199 17507 32205 17541
rect 32239 17507 32245 17541
rect 32199 17469 32245 17507
rect 32199 17435 32205 17469
rect 32239 17435 32245 17469
rect 32199 17397 32245 17435
rect 32199 17363 32205 17397
rect 32239 17363 32245 17397
rect 32199 17347 32245 17363
rect 32657 18621 32703 18637
rect 32657 18587 32663 18621
rect 32697 18587 32703 18621
rect 32657 18549 32703 18587
rect 32657 18515 32663 18549
rect 32697 18515 32703 18549
rect 32657 18477 32703 18515
rect 32657 18443 32663 18477
rect 32697 18443 32703 18477
rect 32657 18405 32703 18443
rect 32657 18371 32663 18405
rect 32697 18371 32703 18405
rect 32657 18333 32703 18371
rect 32657 18299 32663 18333
rect 32697 18299 32703 18333
rect 32657 18261 32703 18299
rect 32657 18227 32663 18261
rect 32697 18227 32703 18261
rect 32657 18189 32703 18227
rect 32657 18155 32663 18189
rect 32697 18155 32703 18189
rect 32657 18117 32703 18155
rect 32657 18083 32663 18117
rect 32697 18083 32703 18117
rect 32657 18045 32703 18083
rect 32657 18011 32663 18045
rect 32697 18011 32703 18045
rect 32657 17973 32703 18011
rect 32657 17939 32663 17973
rect 32697 17939 32703 17973
rect 32657 17901 32703 17939
rect 32657 17867 32663 17901
rect 32697 17867 32703 17901
rect 32657 17829 32703 17867
rect 32657 17795 32663 17829
rect 32697 17795 32703 17829
rect 32657 17757 32703 17795
rect 32657 17723 32663 17757
rect 32697 17723 32703 17757
rect 32657 17685 32703 17723
rect 32657 17651 32663 17685
rect 32697 17651 32703 17685
rect 32657 17613 32703 17651
rect 32657 17579 32663 17613
rect 32697 17579 32703 17613
rect 32657 17541 32703 17579
rect 32657 17507 32663 17541
rect 32697 17507 32703 17541
rect 32657 17469 32703 17507
rect 32657 17435 32663 17469
rect 32697 17435 32703 17469
rect 32657 17397 32703 17435
rect 32657 17363 32663 17397
rect 32697 17363 32703 17397
rect 32657 17347 32703 17363
rect 33115 18621 33161 18637
rect 33115 18587 33121 18621
rect 33155 18587 33161 18621
rect 33115 18549 33161 18587
rect 33115 18515 33121 18549
rect 33155 18515 33161 18549
rect 33115 18477 33161 18515
rect 33115 18443 33121 18477
rect 33155 18443 33161 18477
rect 33115 18405 33161 18443
rect 33115 18371 33121 18405
rect 33155 18371 33161 18405
rect 33115 18333 33161 18371
rect 33115 18299 33121 18333
rect 33155 18299 33161 18333
rect 33115 18261 33161 18299
rect 33115 18227 33121 18261
rect 33155 18227 33161 18261
rect 33115 18189 33161 18227
rect 33115 18155 33121 18189
rect 33155 18155 33161 18189
rect 33115 18117 33161 18155
rect 33115 18083 33121 18117
rect 33155 18083 33161 18117
rect 33115 18045 33161 18083
rect 33115 18011 33121 18045
rect 33155 18011 33161 18045
rect 33115 17973 33161 18011
rect 33115 17939 33121 17973
rect 33155 17939 33161 17973
rect 33115 17901 33161 17939
rect 33115 17867 33121 17901
rect 33155 17867 33161 17901
rect 33115 17829 33161 17867
rect 33115 17795 33121 17829
rect 33155 17795 33161 17829
rect 33115 17757 33161 17795
rect 33115 17723 33121 17757
rect 33155 17723 33161 17757
rect 33115 17685 33161 17723
rect 33115 17651 33121 17685
rect 33155 17651 33161 17685
rect 33115 17613 33161 17651
rect 33115 17579 33121 17613
rect 33155 17579 33161 17613
rect 33115 17541 33161 17579
rect 33115 17507 33121 17541
rect 33155 17507 33161 17541
rect 33115 17469 33161 17507
rect 33115 17435 33121 17469
rect 33155 17435 33161 17469
rect 33115 17397 33161 17435
rect 33115 17363 33121 17397
rect 33155 17363 33161 17397
rect 33115 17347 33161 17363
rect 33573 18621 33619 18637
rect 33573 18587 33579 18621
rect 33613 18587 33619 18621
rect 33573 18549 33619 18587
rect 33573 18515 33579 18549
rect 33613 18515 33619 18549
rect 33573 18477 33619 18515
rect 33573 18443 33579 18477
rect 33613 18443 33619 18477
rect 33573 18405 33619 18443
rect 33573 18371 33579 18405
rect 33613 18371 33619 18405
rect 33573 18333 33619 18371
rect 33573 18299 33579 18333
rect 33613 18299 33619 18333
rect 33573 18261 33619 18299
rect 33573 18227 33579 18261
rect 33613 18227 33619 18261
rect 33573 18189 33619 18227
rect 33573 18155 33579 18189
rect 33613 18155 33619 18189
rect 33573 18117 33619 18155
rect 33573 18083 33579 18117
rect 33613 18083 33619 18117
rect 33573 18045 33619 18083
rect 33573 18011 33579 18045
rect 33613 18011 33619 18045
rect 33573 17973 33619 18011
rect 33573 17939 33579 17973
rect 33613 17939 33619 17973
rect 33573 17901 33619 17939
rect 33573 17867 33579 17901
rect 33613 17867 33619 17901
rect 33573 17829 33619 17867
rect 33573 17795 33579 17829
rect 33613 17795 33619 17829
rect 33573 17757 33619 17795
rect 33573 17723 33579 17757
rect 33613 17723 33619 17757
rect 33573 17685 33619 17723
rect 33573 17651 33579 17685
rect 33613 17651 33619 17685
rect 33573 17613 33619 17651
rect 33573 17579 33579 17613
rect 33613 17579 33619 17613
rect 33573 17541 33619 17579
rect 33573 17507 33579 17541
rect 33613 17507 33619 17541
rect 33573 17469 33619 17507
rect 33573 17435 33579 17469
rect 33613 17435 33619 17469
rect 33573 17397 33619 17435
rect 33573 17363 33579 17397
rect 33613 17363 33619 17397
rect 33573 17347 33619 17363
rect 34031 18621 34077 18637
rect 34031 18587 34037 18621
rect 34071 18587 34077 18621
rect 34031 18549 34077 18587
rect 34031 18515 34037 18549
rect 34071 18515 34077 18549
rect 34031 18477 34077 18515
rect 34031 18443 34037 18477
rect 34071 18443 34077 18477
rect 34031 18405 34077 18443
rect 34031 18371 34037 18405
rect 34071 18371 34077 18405
rect 34031 18333 34077 18371
rect 34031 18299 34037 18333
rect 34071 18299 34077 18333
rect 34031 18261 34077 18299
rect 34031 18227 34037 18261
rect 34071 18227 34077 18261
rect 34031 18189 34077 18227
rect 34031 18155 34037 18189
rect 34071 18155 34077 18189
rect 34031 18117 34077 18155
rect 34031 18083 34037 18117
rect 34071 18083 34077 18117
rect 34031 18045 34077 18083
rect 34031 18011 34037 18045
rect 34071 18011 34077 18045
rect 34031 17973 34077 18011
rect 34031 17939 34037 17973
rect 34071 17939 34077 17973
rect 34031 17901 34077 17939
rect 34031 17867 34037 17901
rect 34071 17867 34077 17901
rect 34031 17829 34077 17867
rect 34031 17795 34037 17829
rect 34071 17795 34077 17829
rect 34031 17757 34077 17795
rect 34031 17723 34037 17757
rect 34071 17723 34077 17757
rect 34031 17685 34077 17723
rect 34031 17651 34037 17685
rect 34071 17651 34077 17685
rect 34031 17613 34077 17651
rect 34031 17579 34037 17613
rect 34071 17579 34077 17613
rect 34031 17541 34077 17579
rect 34031 17507 34037 17541
rect 34071 17507 34077 17541
rect 34031 17469 34077 17507
rect 34031 17435 34037 17469
rect 34071 17435 34077 17469
rect 34031 17397 34077 17435
rect 34031 17363 34037 17397
rect 34071 17363 34077 17397
rect 34031 17347 34077 17363
rect 34489 18621 34535 18637
rect 34489 18587 34495 18621
rect 34529 18587 34535 18621
rect 34489 18549 34535 18587
rect 34489 18515 34495 18549
rect 34529 18515 34535 18549
rect 34489 18477 34535 18515
rect 34489 18443 34495 18477
rect 34529 18443 34535 18477
rect 34489 18405 34535 18443
rect 34489 18371 34495 18405
rect 34529 18371 34535 18405
rect 34489 18333 34535 18371
rect 34489 18299 34495 18333
rect 34529 18299 34535 18333
rect 34489 18261 34535 18299
rect 34489 18227 34495 18261
rect 34529 18227 34535 18261
rect 34489 18189 34535 18227
rect 34489 18155 34495 18189
rect 34529 18155 34535 18189
rect 34489 18117 34535 18155
rect 34489 18083 34495 18117
rect 34529 18083 34535 18117
rect 34489 18045 34535 18083
rect 34489 18011 34495 18045
rect 34529 18011 34535 18045
rect 34489 17973 34535 18011
rect 34489 17939 34495 17973
rect 34529 17939 34535 17973
rect 34489 17901 34535 17939
rect 34489 17867 34495 17901
rect 34529 17867 34535 17901
rect 34489 17829 34535 17867
rect 34489 17795 34495 17829
rect 34529 17795 34535 17829
rect 34489 17757 34535 17795
rect 34489 17723 34495 17757
rect 34529 17723 34535 17757
rect 34489 17685 34535 17723
rect 34489 17651 34495 17685
rect 34529 17651 34535 17685
rect 34489 17613 34535 17651
rect 34489 17579 34495 17613
rect 34529 17579 34535 17613
rect 34489 17541 34535 17579
rect 34489 17507 34495 17541
rect 34529 17507 34535 17541
rect 34489 17469 34535 17507
rect 34489 17435 34495 17469
rect 34529 17435 34535 17469
rect 34489 17397 34535 17435
rect 34489 17363 34495 17397
rect 34529 17363 34535 17397
rect 34489 17347 34535 17363
rect 34947 18621 34993 18637
rect 34947 18587 34953 18621
rect 34987 18587 34993 18621
rect 34947 18549 34993 18587
rect 34947 18515 34953 18549
rect 34987 18515 34993 18549
rect 34947 18477 34993 18515
rect 34947 18443 34953 18477
rect 34987 18443 34993 18477
rect 34947 18405 34993 18443
rect 34947 18371 34953 18405
rect 34987 18371 34993 18405
rect 34947 18333 34993 18371
rect 34947 18299 34953 18333
rect 34987 18299 34993 18333
rect 34947 18261 34993 18299
rect 34947 18227 34953 18261
rect 34987 18227 34993 18261
rect 34947 18189 34993 18227
rect 34947 18155 34953 18189
rect 34987 18155 34993 18189
rect 34947 18117 34993 18155
rect 34947 18083 34953 18117
rect 34987 18083 34993 18117
rect 34947 18045 34993 18083
rect 34947 18011 34953 18045
rect 34987 18011 34993 18045
rect 34947 17973 34993 18011
rect 34947 17939 34953 17973
rect 34987 17939 34993 17973
rect 34947 17901 34993 17939
rect 34947 17867 34953 17901
rect 34987 17867 34993 17901
rect 34947 17829 34993 17867
rect 34947 17795 34953 17829
rect 34987 17795 34993 17829
rect 34947 17757 34993 17795
rect 34947 17723 34953 17757
rect 34987 17723 34993 17757
rect 34947 17685 34993 17723
rect 34947 17651 34953 17685
rect 34987 17651 34993 17685
rect 34947 17613 34993 17651
rect 34947 17579 34953 17613
rect 34987 17579 34993 17613
rect 34947 17541 34993 17579
rect 34947 17507 34953 17541
rect 34987 17507 34993 17541
rect 34947 17469 34993 17507
rect 34947 17435 34953 17469
rect 34987 17435 34993 17469
rect 34947 17397 34993 17435
rect 34947 17363 34953 17397
rect 34987 17363 34993 17397
rect 34947 17347 34993 17363
rect 35405 18621 35451 18637
rect 35405 18587 35411 18621
rect 35445 18587 35451 18621
rect 35405 18549 35451 18587
rect 35405 18515 35411 18549
rect 35445 18515 35451 18549
rect 35405 18477 35451 18515
rect 35405 18443 35411 18477
rect 35445 18443 35451 18477
rect 35405 18405 35451 18443
rect 35405 18371 35411 18405
rect 35445 18371 35451 18405
rect 35405 18333 35451 18371
rect 35405 18299 35411 18333
rect 35445 18299 35451 18333
rect 35405 18261 35451 18299
rect 35405 18227 35411 18261
rect 35445 18227 35451 18261
rect 35405 18189 35451 18227
rect 35405 18155 35411 18189
rect 35445 18155 35451 18189
rect 35405 18117 35451 18155
rect 35405 18083 35411 18117
rect 35445 18083 35451 18117
rect 35405 18045 35451 18083
rect 35405 18011 35411 18045
rect 35445 18011 35451 18045
rect 35405 17973 35451 18011
rect 35405 17939 35411 17973
rect 35445 17939 35451 17973
rect 35405 17901 35451 17939
rect 35405 17867 35411 17901
rect 35445 17867 35451 17901
rect 35405 17829 35451 17867
rect 35405 17795 35411 17829
rect 35445 17795 35451 17829
rect 35405 17757 35451 17795
rect 35405 17723 35411 17757
rect 35445 17723 35451 17757
rect 35405 17685 35451 17723
rect 35405 17651 35411 17685
rect 35445 17651 35451 17685
rect 35405 17613 35451 17651
rect 35405 17579 35411 17613
rect 35445 17579 35451 17613
rect 35405 17541 35451 17579
rect 35405 17507 35411 17541
rect 35445 17507 35451 17541
rect 35405 17469 35451 17507
rect 35405 17435 35411 17469
rect 35445 17435 35451 17469
rect 35405 17397 35451 17435
rect 35405 17363 35411 17397
rect 35445 17363 35451 17397
rect 35405 17347 35451 17363
rect 35863 18621 35909 18637
rect 35863 18587 35869 18621
rect 35903 18587 35909 18621
rect 35863 18549 35909 18587
rect 35863 18515 35869 18549
rect 35903 18515 35909 18549
rect 35863 18477 35909 18515
rect 35863 18443 35869 18477
rect 35903 18443 35909 18477
rect 35863 18405 35909 18443
rect 35863 18371 35869 18405
rect 35903 18371 35909 18405
rect 35863 18333 35909 18371
rect 35863 18299 35869 18333
rect 35903 18299 35909 18333
rect 35863 18261 35909 18299
rect 35863 18227 35869 18261
rect 35903 18227 35909 18261
rect 35863 18189 35909 18227
rect 35863 18155 35869 18189
rect 35903 18155 35909 18189
rect 35863 18117 35909 18155
rect 35863 18083 35869 18117
rect 35903 18083 35909 18117
rect 35863 18045 35909 18083
rect 35863 18011 35869 18045
rect 35903 18011 35909 18045
rect 35863 17973 35909 18011
rect 35863 17939 35869 17973
rect 35903 17939 35909 17973
rect 35863 17901 35909 17939
rect 35863 17867 35869 17901
rect 35903 17867 35909 17901
rect 35863 17829 35909 17867
rect 35863 17795 35869 17829
rect 35903 17795 35909 17829
rect 35863 17757 35909 17795
rect 35863 17723 35869 17757
rect 35903 17723 35909 17757
rect 35863 17685 35909 17723
rect 35863 17651 35869 17685
rect 35903 17651 35909 17685
rect 35863 17613 35909 17651
rect 35863 17579 35869 17613
rect 35903 17579 35909 17613
rect 35863 17541 35909 17579
rect 35863 17507 35869 17541
rect 35903 17507 35909 17541
rect 35863 17469 35909 17507
rect 35863 17435 35869 17469
rect 35903 17435 35909 17469
rect 35863 17397 35909 17435
rect 35863 17363 35869 17397
rect 35903 17363 35909 17397
rect 35863 17347 35909 17363
rect 36321 18621 36367 18637
rect 36321 18587 36327 18621
rect 36361 18587 36367 18621
rect 36321 18549 36367 18587
rect 36321 18515 36327 18549
rect 36361 18515 36367 18549
rect 36321 18477 36367 18515
rect 36321 18443 36327 18477
rect 36361 18443 36367 18477
rect 36321 18405 36367 18443
rect 36321 18371 36327 18405
rect 36361 18371 36367 18405
rect 36321 18333 36367 18371
rect 36321 18299 36327 18333
rect 36361 18299 36367 18333
rect 36321 18261 36367 18299
rect 36321 18227 36327 18261
rect 36361 18227 36367 18261
rect 36321 18189 36367 18227
rect 36321 18155 36327 18189
rect 36361 18155 36367 18189
rect 36321 18117 36367 18155
rect 36321 18083 36327 18117
rect 36361 18083 36367 18117
rect 36321 18045 36367 18083
rect 36321 18011 36327 18045
rect 36361 18011 36367 18045
rect 36321 17973 36367 18011
rect 36321 17939 36327 17973
rect 36361 17939 36367 17973
rect 36321 17901 36367 17939
rect 36321 17867 36327 17901
rect 36361 17867 36367 17901
rect 36321 17829 36367 17867
rect 36321 17795 36327 17829
rect 36361 17795 36367 17829
rect 36321 17757 36367 17795
rect 36321 17723 36327 17757
rect 36361 17723 36367 17757
rect 36321 17685 36367 17723
rect 36321 17651 36327 17685
rect 36361 17651 36367 17685
rect 36321 17613 36367 17651
rect 36321 17579 36327 17613
rect 36361 17579 36367 17613
rect 36321 17541 36367 17579
rect 36321 17507 36327 17541
rect 36361 17507 36367 17541
rect 36321 17469 36367 17507
rect 36321 17435 36327 17469
rect 36361 17435 36367 17469
rect 36321 17397 36367 17435
rect 36321 17363 36327 17397
rect 36361 17363 36367 17397
rect 36321 17347 36367 17363
rect 36779 18621 36825 18637
rect 36779 18587 36785 18621
rect 36819 18587 36825 18621
rect 36779 18549 36825 18587
rect 36779 18515 36785 18549
rect 36819 18515 36825 18549
rect 36779 18477 36825 18515
rect 36779 18443 36785 18477
rect 36819 18443 36825 18477
rect 36779 18405 36825 18443
rect 36779 18371 36785 18405
rect 36819 18371 36825 18405
rect 36779 18333 36825 18371
rect 36779 18299 36785 18333
rect 36819 18299 36825 18333
rect 36779 18261 36825 18299
rect 36779 18227 36785 18261
rect 36819 18227 36825 18261
rect 36779 18189 36825 18227
rect 36779 18155 36785 18189
rect 36819 18155 36825 18189
rect 36779 18117 36825 18155
rect 36779 18083 36785 18117
rect 36819 18083 36825 18117
rect 36779 18045 36825 18083
rect 36779 18011 36785 18045
rect 36819 18011 36825 18045
rect 36779 17973 36825 18011
rect 36779 17939 36785 17973
rect 36819 17939 36825 17973
rect 36779 17901 36825 17939
rect 36779 17867 36785 17901
rect 36819 17867 36825 17901
rect 36779 17829 36825 17867
rect 36779 17795 36785 17829
rect 36819 17795 36825 17829
rect 36779 17757 36825 17795
rect 36779 17723 36785 17757
rect 36819 17723 36825 17757
rect 36779 17685 36825 17723
rect 36779 17651 36785 17685
rect 36819 17651 36825 17685
rect 36779 17613 36825 17651
rect 36779 17579 36785 17613
rect 36819 17579 36825 17613
rect 36779 17541 36825 17579
rect 36779 17507 36785 17541
rect 36819 17507 36825 17541
rect 36779 17469 36825 17507
rect 36779 17435 36785 17469
rect 36819 17435 36825 17469
rect 36779 17397 36825 17435
rect 36779 17363 36785 17397
rect 36819 17363 36825 17397
rect 36779 17347 36825 17363
rect 37237 18621 37283 18637
rect 37237 18587 37243 18621
rect 37277 18587 37283 18621
rect 37237 18549 37283 18587
rect 37237 18515 37243 18549
rect 37277 18515 37283 18549
rect 37237 18477 37283 18515
rect 37237 18443 37243 18477
rect 37277 18443 37283 18477
rect 37237 18405 37283 18443
rect 37237 18371 37243 18405
rect 37277 18371 37283 18405
rect 37237 18333 37283 18371
rect 37237 18299 37243 18333
rect 37277 18299 37283 18333
rect 37237 18261 37283 18299
rect 37237 18227 37243 18261
rect 37277 18227 37283 18261
rect 37237 18189 37283 18227
rect 37237 18155 37243 18189
rect 37277 18155 37283 18189
rect 37237 18117 37283 18155
rect 37237 18083 37243 18117
rect 37277 18083 37283 18117
rect 37237 18045 37283 18083
rect 37237 18011 37243 18045
rect 37277 18011 37283 18045
rect 37237 17973 37283 18011
rect 37237 17939 37243 17973
rect 37277 17939 37283 17973
rect 37237 17901 37283 17939
rect 37237 17867 37243 17901
rect 37277 17867 37283 17901
rect 37237 17829 37283 17867
rect 37237 17795 37243 17829
rect 37277 17795 37283 17829
rect 37237 17757 37283 17795
rect 37237 17723 37243 17757
rect 37277 17723 37283 17757
rect 37237 17685 37283 17723
rect 37237 17651 37243 17685
rect 37277 17651 37283 17685
rect 37237 17613 37283 17651
rect 37237 17579 37243 17613
rect 37277 17579 37283 17613
rect 37237 17541 37283 17579
rect 37237 17507 37243 17541
rect 37277 17507 37283 17541
rect 37237 17469 37283 17507
rect 37237 17435 37243 17469
rect 37277 17435 37283 17469
rect 37237 17397 37283 17435
rect 37237 17363 37243 17397
rect 37277 17363 37283 17397
rect 37237 17347 37283 17363
rect 37695 18621 37741 18637
rect 37695 18587 37701 18621
rect 37735 18587 37741 18621
rect 37695 18549 37741 18587
rect 37695 18515 37701 18549
rect 37735 18515 37741 18549
rect 37695 18477 37741 18515
rect 37695 18443 37701 18477
rect 37735 18443 37741 18477
rect 37695 18405 37741 18443
rect 37695 18371 37701 18405
rect 37735 18371 37741 18405
rect 37695 18333 37741 18371
rect 37695 18299 37701 18333
rect 37735 18299 37741 18333
rect 37695 18261 37741 18299
rect 37695 18227 37701 18261
rect 37735 18227 37741 18261
rect 37695 18189 37741 18227
rect 37695 18155 37701 18189
rect 37735 18155 37741 18189
rect 37695 18117 37741 18155
rect 37695 18083 37701 18117
rect 37735 18083 37741 18117
rect 37695 18045 37741 18083
rect 37695 18011 37701 18045
rect 37735 18011 37741 18045
rect 37695 17973 37741 18011
rect 37695 17939 37701 17973
rect 37735 17939 37741 17973
rect 37695 17901 37741 17939
rect 37695 17867 37701 17901
rect 37735 17867 37741 17901
rect 37695 17829 37741 17867
rect 37695 17795 37701 17829
rect 37735 17795 37741 17829
rect 37695 17757 37741 17795
rect 37695 17723 37701 17757
rect 37735 17723 37741 17757
rect 37695 17685 37741 17723
rect 37695 17651 37701 17685
rect 37735 17651 37741 17685
rect 37695 17613 37741 17651
rect 37695 17579 37701 17613
rect 37735 17579 37741 17613
rect 37695 17541 37741 17579
rect 37695 17507 37701 17541
rect 37735 17507 37741 17541
rect 37695 17469 37741 17507
rect 37695 17435 37701 17469
rect 37735 17435 37741 17469
rect 37695 17397 37741 17435
rect 37695 17363 37701 17397
rect 37735 17363 37741 17397
rect 37695 17347 37741 17363
rect 38153 18621 38199 18637
rect 38153 18587 38159 18621
rect 38193 18587 38199 18621
rect 38153 18549 38199 18587
rect 38153 18515 38159 18549
rect 38193 18515 38199 18549
rect 38153 18477 38199 18515
rect 38153 18443 38159 18477
rect 38193 18443 38199 18477
rect 38153 18405 38199 18443
rect 38153 18371 38159 18405
rect 38193 18371 38199 18405
rect 38153 18333 38199 18371
rect 38153 18299 38159 18333
rect 38193 18299 38199 18333
rect 38153 18261 38199 18299
rect 38153 18227 38159 18261
rect 38193 18227 38199 18261
rect 38153 18189 38199 18227
rect 38153 18155 38159 18189
rect 38193 18155 38199 18189
rect 38153 18117 38199 18155
rect 38153 18083 38159 18117
rect 38193 18083 38199 18117
rect 38153 18045 38199 18083
rect 38153 18011 38159 18045
rect 38193 18011 38199 18045
rect 38153 17973 38199 18011
rect 38153 17939 38159 17973
rect 38193 17939 38199 17973
rect 38153 17901 38199 17939
rect 38153 17867 38159 17901
rect 38193 17867 38199 17901
rect 38153 17829 38199 17867
rect 38153 17795 38159 17829
rect 38193 17795 38199 17829
rect 38153 17757 38199 17795
rect 38153 17723 38159 17757
rect 38193 17723 38199 17757
rect 38153 17685 38199 17723
rect 38153 17651 38159 17685
rect 38193 17651 38199 17685
rect 38153 17613 38199 17651
rect 38153 17579 38159 17613
rect 38193 17579 38199 17613
rect 38153 17541 38199 17579
rect 38153 17507 38159 17541
rect 38193 17507 38199 17541
rect 38153 17469 38199 17507
rect 38153 17435 38159 17469
rect 38193 17435 38199 17469
rect 38153 17397 38199 17435
rect 38153 17363 38159 17397
rect 38193 17363 38199 17397
rect 38153 17347 38199 17363
rect 38611 18621 38657 18637
rect 38611 18587 38617 18621
rect 38651 18587 38657 18621
rect 38611 18549 38657 18587
rect 38611 18515 38617 18549
rect 38651 18515 38657 18549
rect 38611 18477 38657 18515
rect 38611 18443 38617 18477
rect 38651 18443 38657 18477
rect 38611 18405 38657 18443
rect 38611 18371 38617 18405
rect 38651 18371 38657 18405
rect 38611 18333 38657 18371
rect 38611 18299 38617 18333
rect 38651 18299 38657 18333
rect 38611 18261 38657 18299
rect 38611 18227 38617 18261
rect 38651 18227 38657 18261
rect 38611 18189 38657 18227
rect 38611 18155 38617 18189
rect 38651 18155 38657 18189
rect 38611 18117 38657 18155
rect 38611 18083 38617 18117
rect 38651 18083 38657 18117
rect 38611 18045 38657 18083
rect 38611 18011 38617 18045
rect 38651 18011 38657 18045
rect 38611 17973 38657 18011
rect 38611 17939 38617 17973
rect 38651 17939 38657 17973
rect 38611 17901 38657 17939
rect 38611 17867 38617 17901
rect 38651 17867 38657 17901
rect 38611 17829 38657 17867
rect 38611 17795 38617 17829
rect 38651 17795 38657 17829
rect 38611 17757 38657 17795
rect 38611 17723 38617 17757
rect 38651 17723 38657 17757
rect 38611 17685 38657 17723
rect 38611 17651 38617 17685
rect 38651 17651 38657 17685
rect 38611 17613 38657 17651
rect 38611 17579 38617 17613
rect 38651 17579 38657 17613
rect 38611 17541 38657 17579
rect 38611 17507 38617 17541
rect 38651 17507 38657 17541
rect 38611 17469 38657 17507
rect 38611 17435 38617 17469
rect 38651 17435 38657 17469
rect 38611 17397 38657 17435
rect 38611 17363 38617 17397
rect 38651 17363 38657 17397
rect 38611 17347 38657 17363
rect 39069 18621 39115 18637
rect 39069 18587 39075 18621
rect 39109 18587 39115 18621
rect 39069 18549 39115 18587
rect 39069 18515 39075 18549
rect 39109 18515 39115 18549
rect 39069 18477 39115 18515
rect 39069 18443 39075 18477
rect 39109 18443 39115 18477
rect 39069 18405 39115 18443
rect 39069 18371 39075 18405
rect 39109 18371 39115 18405
rect 39069 18333 39115 18371
rect 39069 18299 39075 18333
rect 39109 18299 39115 18333
rect 39069 18261 39115 18299
rect 39069 18227 39075 18261
rect 39109 18227 39115 18261
rect 39069 18189 39115 18227
rect 39069 18155 39075 18189
rect 39109 18155 39115 18189
rect 39069 18117 39115 18155
rect 39069 18083 39075 18117
rect 39109 18083 39115 18117
rect 39069 18045 39115 18083
rect 39069 18011 39075 18045
rect 39109 18011 39115 18045
rect 39069 17973 39115 18011
rect 39069 17939 39075 17973
rect 39109 17939 39115 17973
rect 39069 17901 39115 17939
rect 39069 17867 39075 17901
rect 39109 17867 39115 17901
rect 39069 17829 39115 17867
rect 39069 17795 39075 17829
rect 39109 17795 39115 17829
rect 39069 17757 39115 17795
rect 39069 17723 39075 17757
rect 39109 17723 39115 17757
rect 39069 17685 39115 17723
rect 39069 17651 39075 17685
rect 39109 17651 39115 17685
rect 39069 17613 39115 17651
rect 39069 17579 39075 17613
rect 39109 17579 39115 17613
rect 39069 17541 39115 17579
rect 39069 17507 39075 17541
rect 39109 17507 39115 17541
rect 39069 17469 39115 17507
rect 39069 17435 39075 17469
rect 39109 17435 39115 17469
rect 39069 17397 39115 17435
rect 39069 17363 39075 17397
rect 39109 17363 39115 17397
rect 39069 17347 39115 17363
rect 39527 18621 39573 18637
rect 39527 18587 39533 18621
rect 39567 18587 39573 18621
rect 39527 18549 39573 18587
rect 39527 18515 39533 18549
rect 39567 18515 39573 18549
rect 39527 18477 39573 18515
rect 39527 18443 39533 18477
rect 39567 18443 39573 18477
rect 39527 18405 39573 18443
rect 39527 18371 39533 18405
rect 39567 18371 39573 18405
rect 39527 18333 39573 18371
rect 39527 18299 39533 18333
rect 39567 18299 39573 18333
rect 39527 18261 39573 18299
rect 39527 18227 39533 18261
rect 39567 18227 39573 18261
rect 39527 18189 39573 18227
rect 39527 18155 39533 18189
rect 39567 18155 39573 18189
rect 39527 18117 39573 18155
rect 39527 18083 39533 18117
rect 39567 18083 39573 18117
rect 39527 18045 39573 18083
rect 39527 18011 39533 18045
rect 39567 18011 39573 18045
rect 39527 17973 39573 18011
rect 39527 17939 39533 17973
rect 39567 17939 39573 17973
rect 39527 17901 39573 17939
rect 39527 17867 39533 17901
rect 39567 17867 39573 17901
rect 39527 17829 39573 17867
rect 39527 17795 39533 17829
rect 39567 17795 39573 17829
rect 39527 17757 39573 17795
rect 39527 17723 39533 17757
rect 39567 17723 39573 17757
rect 39527 17685 39573 17723
rect 39527 17651 39533 17685
rect 39567 17651 39573 17685
rect 39527 17613 39573 17651
rect 39527 17579 39533 17613
rect 39567 17579 39573 17613
rect 39527 17541 39573 17579
rect 39527 17507 39533 17541
rect 39567 17507 39573 17541
rect 39527 17469 39573 17507
rect 39527 17435 39533 17469
rect 39567 17435 39573 17469
rect 39527 17397 39573 17435
rect 39527 17363 39533 17397
rect 39567 17363 39573 17397
rect 39527 17347 39573 17363
rect 39985 18621 40031 18637
rect 39985 18587 39991 18621
rect 40025 18587 40031 18621
rect 39985 18549 40031 18587
rect 39985 18515 39991 18549
rect 40025 18515 40031 18549
rect 39985 18477 40031 18515
rect 39985 18443 39991 18477
rect 40025 18443 40031 18477
rect 39985 18405 40031 18443
rect 39985 18371 39991 18405
rect 40025 18371 40031 18405
rect 39985 18333 40031 18371
rect 39985 18299 39991 18333
rect 40025 18299 40031 18333
rect 39985 18261 40031 18299
rect 39985 18227 39991 18261
rect 40025 18227 40031 18261
rect 39985 18189 40031 18227
rect 39985 18155 39991 18189
rect 40025 18155 40031 18189
rect 39985 18117 40031 18155
rect 39985 18083 39991 18117
rect 40025 18083 40031 18117
rect 39985 18045 40031 18083
rect 39985 18011 39991 18045
rect 40025 18011 40031 18045
rect 39985 17973 40031 18011
rect 39985 17939 39991 17973
rect 40025 17939 40031 17973
rect 39985 17901 40031 17939
rect 39985 17867 39991 17901
rect 40025 17867 40031 17901
rect 39985 17829 40031 17867
rect 39985 17795 39991 17829
rect 40025 17795 40031 17829
rect 39985 17757 40031 17795
rect 39985 17723 39991 17757
rect 40025 17723 40031 17757
rect 39985 17685 40031 17723
rect 39985 17651 39991 17685
rect 40025 17651 40031 17685
rect 39985 17613 40031 17651
rect 39985 17579 39991 17613
rect 40025 17579 40031 17613
rect 39985 17541 40031 17579
rect 39985 17507 39991 17541
rect 40025 17507 40031 17541
rect 39985 17469 40031 17507
rect 39985 17435 39991 17469
rect 40025 17435 40031 17469
rect 39985 17397 40031 17435
rect 39985 17363 39991 17397
rect 40025 17363 40031 17397
rect 39985 17347 40031 17363
rect 40443 18621 40489 18637
rect 40443 18587 40449 18621
rect 40483 18587 40489 18621
rect 40443 18549 40489 18587
rect 40443 18515 40449 18549
rect 40483 18515 40489 18549
rect 40443 18477 40489 18515
rect 40443 18443 40449 18477
rect 40483 18443 40489 18477
rect 40443 18405 40489 18443
rect 40443 18371 40449 18405
rect 40483 18371 40489 18405
rect 40443 18333 40489 18371
rect 40443 18299 40449 18333
rect 40483 18299 40489 18333
rect 40443 18261 40489 18299
rect 40443 18227 40449 18261
rect 40483 18227 40489 18261
rect 40443 18189 40489 18227
rect 40443 18155 40449 18189
rect 40483 18155 40489 18189
rect 40443 18117 40489 18155
rect 40443 18083 40449 18117
rect 40483 18083 40489 18117
rect 40443 18045 40489 18083
rect 40443 18011 40449 18045
rect 40483 18011 40489 18045
rect 40443 17973 40489 18011
rect 40443 17939 40449 17973
rect 40483 17939 40489 17973
rect 40443 17901 40489 17939
rect 40443 17867 40449 17901
rect 40483 17867 40489 17901
rect 40443 17829 40489 17867
rect 40443 17795 40449 17829
rect 40483 17795 40489 17829
rect 40443 17757 40489 17795
rect 40443 17723 40449 17757
rect 40483 17723 40489 17757
rect 40443 17685 40489 17723
rect 40443 17651 40449 17685
rect 40483 17651 40489 17685
rect 40443 17613 40489 17651
rect 40443 17579 40449 17613
rect 40483 17579 40489 17613
rect 40443 17541 40489 17579
rect 40443 17507 40449 17541
rect 40483 17507 40489 17541
rect 40443 17469 40489 17507
rect 40443 17435 40449 17469
rect 40483 17435 40489 17469
rect 40443 17397 40489 17435
rect 40443 17363 40449 17397
rect 40483 17363 40489 17397
rect 40443 17347 40489 17363
rect 40901 18621 40947 18637
rect 40901 18587 40907 18621
rect 40941 18587 40947 18621
rect 40901 18549 40947 18587
rect 40901 18515 40907 18549
rect 40941 18515 40947 18549
rect 40901 18477 40947 18515
rect 40901 18443 40907 18477
rect 40941 18443 40947 18477
rect 40901 18405 40947 18443
rect 40901 18371 40907 18405
rect 40941 18371 40947 18405
rect 40901 18333 40947 18371
rect 40901 18299 40907 18333
rect 40941 18299 40947 18333
rect 40901 18261 40947 18299
rect 40901 18227 40907 18261
rect 40941 18227 40947 18261
rect 40901 18189 40947 18227
rect 40901 18155 40907 18189
rect 40941 18155 40947 18189
rect 40901 18117 40947 18155
rect 40901 18083 40907 18117
rect 40941 18083 40947 18117
rect 40901 18045 40947 18083
rect 40901 18011 40907 18045
rect 40941 18011 40947 18045
rect 40901 17973 40947 18011
rect 40901 17939 40907 17973
rect 40941 17939 40947 17973
rect 40901 17901 40947 17939
rect 40901 17867 40907 17901
rect 40941 17867 40947 17901
rect 40901 17829 40947 17867
rect 40901 17795 40907 17829
rect 40941 17795 40947 17829
rect 40901 17757 40947 17795
rect 40901 17723 40907 17757
rect 40941 17723 40947 17757
rect 40901 17685 40947 17723
rect 40901 17651 40907 17685
rect 40941 17651 40947 17685
rect 40901 17613 40947 17651
rect 40901 17579 40907 17613
rect 40941 17579 40947 17613
rect 40901 17541 40947 17579
rect 40901 17507 40907 17541
rect 40941 17507 40947 17541
rect 40901 17469 40947 17507
rect 40901 17435 40907 17469
rect 40941 17435 40947 17469
rect 40901 17397 40947 17435
rect 40901 17363 40907 17397
rect 40941 17363 40947 17397
rect 40901 17347 40947 17363
rect 41359 18621 41405 18637
rect 41359 18587 41365 18621
rect 41399 18587 41405 18621
rect 41359 18549 41405 18587
rect 41359 18515 41365 18549
rect 41399 18515 41405 18549
rect 41359 18477 41405 18515
rect 41359 18443 41365 18477
rect 41399 18443 41405 18477
rect 41359 18405 41405 18443
rect 41359 18371 41365 18405
rect 41399 18371 41405 18405
rect 41359 18333 41405 18371
rect 41359 18299 41365 18333
rect 41399 18299 41405 18333
rect 41359 18261 41405 18299
rect 41359 18227 41365 18261
rect 41399 18227 41405 18261
rect 41359 18189 41405 18227
rect 41359 18155 41365 18189
rect 41399 18155 41405 18189
rect 41359 18117 41405 18155
rect 41359 18083 41365 18117
rect 41399 18083 41405 18117
rect 41359 18045 41405 18083
rect 41359 18011 41365 18045
rect 41399 18011 41405 18045
rect 41359 17973 41405 18011
rect 41359 17939 41365 17973
rect 41399 17939 41405 17973
rect 41359 17901 41405 17939
rect 41359 17867 41365 17901
rect 41399 17867 41405 17901
rect 41359 17829 41405 17867
rect 41359 17795 41365 17829
rect 41399 17795 41405 17829
rect 41359 17757 41405 17795
rect 41359 17723 41365 17757
rect 41399 17723 41405 17757
rect 41359 17685 41405 17723
rect 41359 17651 41365 17685
rect 41399 17651 41405 17685
rect 41359 17613 41405 17651
rect 41359 17579 41365 17613
rect 41399 17579 41405 17613
rect 41359 17541 41405 17579
rect 41359 17507 41365 17541
rect 41399 17507 41405 17541
rect 41359 17469 41405 17507
rect 41359 17435 41365 17469
rect 41399 17435 41405 17469
rect 41359 17397 41405 17435
rect 41359 17363 41365 17397
rect 41399 17363 41405 17397
rect 41359 17347 41405 17363
rect 41817 18621 41863 18637
rect 41817 18587 41823 18621
rect 41857 18587 41863 18621
rect 41817 18549 41863 18587
rect 41817 18515 41823 18549
rect 41857 18515 41863 18549
rect 41817 18477 41863 18515
rect 41817 18443 41823 18477
rect 41857 18443 41863 18477
rect 41817 18405 41863 18443
rect 41817 18371 41823 18405
rect 41857 18371 41863 18405
rect 41817 18333 41863 18371
rect 41817 18299 41823 18333
rect 41857 18299 41863 18333
rect 41817 18261 41863 18299
rect 41817 18227 41823 18261
rect 41857 18227 41863 18261
rect 41817 18189 41863 18227
rect 41817 18155 41823 18189
rect 41857 18155 41863 18189
rect 41817 18117 41863 18155
rect 41817 18083 41823 18117
rect 41857 18083 41863 18117
rect 41817 18045 41863 18083
rect 41817 18011 41823 18045
rect 41857 18011 41863 18045
rect 41817 17973 41863 18011
rect 41817 17939 41823 17973
rect 41857 17939 41863 17973
rect 41817 17901 41863 17939
rect 41817 17867 41823 17901
rect 41857 17867 41863 17901
rect 41817 17829 41863 17867
rect 41817 17795 41823 17829
rect 41857 17795 41863 17829
rect 41817 17757 41863 17795
rect 41817 17723 41823 17757
rect 41857 17723 41863 17757
rect 41817 17685 41863 17723
rect 41817 17651 41823 17685
rect 41857 17651 41863 17685
rect 41817 17613 41863 17651
rect 41817 17579 41823 17613
rect 41857 17579 41863 17613
rect 41817 17541 41863 17579
rect 41817 17507 41823 17541
rect 41857 17507 41863 17541
rect 41817 17469 41863 17507
rect 41817 17435 41823 17469
rect 41857 17435 41863 17469
rect 41817 17397 41863 17435
rect 41817 17363 41823 17397
rect 41857 17363 41863 17397
rect 41817 17347 41863 17363
rect 42275 18621 42321 18637
rect 42275 18587 42281 18621
rect 42315 18587 42321 18621
rect 42275 18549 42321 18587
rect 42275 18515 42281 18549
rect 42315 18515 42321 18549
rect 42275 18477 42321 18515
rect 42275 18443 42281 18477
rect 42315 18443 42321 18477
rect 42275 18405 42321 18443
rect 42275 18371 42281 18405
rect 42315 18371 42321 18405
rect 42275 18333 42321 18371
rect 42275 18299 42281 18333
rect 42315 18299 42321 18333
rect 42275 18261 42321 18299
rect 42275 18227 42281 18261
rect 42315 18227 42321 18261
rect 42275 18189 42321 18227
rect 42275 18155 42281 18189
rect 42315 18155 42321 18189
rect 42275 18117 42321 18155
rect 42275 18083 42281 18117
rect 42315 18083 42321 18117
rect 42275 18045 42321 18083
rect 42275 18011 42281 18045
rect 42315 18011 42321 18045
rect 42275 17973 42321 18011
rect 42275 17939 42281 17973
rect 42315 17939 42321 17973
rect 42275 17901 42321 17939
rect 42275 17867 42281 17901
rect 42315 17867 42321 17901
rect 42275 17829 42321 17867
rect 42275 17795 42281 17829
rect 42315 17795 42321 17829
rect 42275 17757 42321 17795
rect 42275 17723 42281 17757
rect 42315 17723 42321 17757
rect 42275 17685 42321 17723
rect 42275 17651 42281 17685
rect 42315 17651 42321 17685
rect 42275 17613 42321 17651
rect 42275 17579 42281 17613
rect 42315 17579 42321 17613
rect 42275 17541 42321 17579
rect 42275 17507 42281 17541
rect 42315 17507 42321 17541
rect 42275 17469 42321 17507
rect 42275 17435 42281 17469
rect 42315 17435 42321 17469
rect 42275 17397 42321 17435
rect 42275 17363 42281 17397
rect 42315 17363 42321 17397
rect 42275 17347 42321 17363
rect 42733 18621 42779 18637
rect 42733 18587 42739 18621
rect 42773 18587 42779 18621
rect 42733 18549 42779 18587
rect 42733 18515 42739 18549
rect 42773 18515 42779 18549
rect 42733 18477 42779 18515
rect 42733 18443 42739 18477
rect 42773 18443 42779 18477
rect 42733 18405 42779 18443
rect 42733 18371 42739 18405
rect 42773 18371 42779 18405
rect 42733 18333 42779 18371
rect 42733 18299 42739 18333
rect 42773 18299 42779 18333
rect 42733 18261 42779 18299
rect 42733 18227 42739 18261
rect 42773 18227 42779 18261
rect 42733 18189 42779 18227
rect 42733 18155 42739 18189
rect 42773 18155 42779 18189
rect 42733 18117 42779 18155
rect 42733 18083 42739 18117
rect 42773 18083 42779 18117
rect 42733 18045 42779 18083
rect 42733 18011 42739 18045
rect 42773 18011 42779 18045
rect 42733 17973 42779 18011
rect 42733 17939 42739 17973
rect 42773 17939 42779 17973
rect 42733 17901 42779 17939
rect 42733 17867 42739 17901
rect 42773 17867 42779 17901
rect 42733 17829 42779 17867
rect 42733 17795 42739 17829
rect 42773 17795 42779 17829
rect 42733 17757 42779 17795
rect 42733 17723 42739 17757
rect 42773 17723 42779 17757
rect 42733 17685 42779 17723
rect 42733 17651 42739 17685
rect 42773 17651 42779 17685
rect 42733 17613 42779 17651
rect 42733 17579 42739 17613
rect 42773 17579 42779 17613
rect 42733 17541 42779 17579
rect 42733 17507 42739 17541
rect 42773 17507 42779 17541
rect 42733 17469 42779 17507
rect 42733 17435 42739 17469
rect 42773 17435 42779 17469
rect 42733 17397 42779 17435
rect 42733 17363 42739 17397
rect 42773 17363 42779 17397
rect 42733 17347 42779 17363
rect 43191 18621 43237 18637
rect 43191 18587 43197 18621
rect 43231 18587 43237 18621
rect 43191 18549 43237 18587
rect 43191 18515 43197 18549
rect 43231 18515 43237 18549
rect 43191 18477 43237 18515
rect 43191 18443 43197 18477
rect 43231 18443 43237 18477
rect 43191 18405 43237 18443
rect 43191 18371 43197 18405
rect 43231 18371 43237 18405
rect 43191 18333 43237 18371
rect 43191 18299 43197 18333
rect 43231 18299 43237 18333
rect 43191 18261 43237 18299
rect 43191 18227 43197 18261
rect 43231 18227 43237 18261
rect 43191 18189 43237 18227
rect 43191 18155 43197 18189
rect 43231 18155 43237 18189
rect 43191 18117 43237 18155
rect 43191 18083 43197 18117
rect 43231 18083 43237 18117
rect 43191 18045 43237 18083
rect 43191 18011 43197 18045
rect 43231 18011 43237 18045
rect 43191 17973 43237 18011
rect 43191 17939 43197 17973
rect 43231 17939 43237 17973
rect 43191 17901 43237 17939
rect 43191 17867 43197 17901
rect 43231 17867 43237 17901
rect 43191 17829 43237 17867
rect 43191 17795 43197 17829
rect 43231 17795 43237 17829
rect 43191 17757 43237 17795
rect 43191 17723 43197 17757
rect 43231 17723 43237 17757
rect 43191 17685 43237 17723
rect 43191 17651 43197 17685
rect 43231 17651 43237 17685
rect 43191 17613 43237 17651
rect 43191 17579 43197 17613
rect 43231 17579 43237 17613
rect 43191 17541 43237 17579
rect 43191 17507 43197 17541
rect 43231 17507 43237 17541
rect 43191 17469 43237 17507
rect 43191 17435 43197 17469
rect 43231 17435 43237 17469
rect 43191 17397 43237 17435
rect 43191 17363 43197 17397
rect 43231 17363 43237 17397
rect 43191 17347 43237 17363
rect 43649 18621 43695 18637
rect 43649 18587 43655 18621
rect 43689 18587 43695 18621
rect 43649 18549 43695 18587
rect 43649 18515 43655 18549
rect 43689 18515 43695 18549
rect 43649 18477 43695 18515
rect 43649 18443 43655 18477
rect 43689 18443 43695 18477
rect 43649 18405 43695 18443
rect 43649 18371 43655 18405
rect 43689 18371 43695 18405
rect 43649 18333 43695 18371
rect 43649 18299 43655 18333
rect 43689 18299 43695 18333
rect 43649 18261 43695 18299
rect 43649 18227 43655 18261
rect 43689 18227 43695 18261
rect 43649 18189 43695 18227
rect 43649 18155 43655 18189
rect 43689 18155 43695 18189
rect 43649 18117 43695 18155
rect 43649 18083 43655 18117
rect 43689 18083 43695 18117
rect 43649 18045 43695 18083
rect 43649 18011 43655 18045
rect 43689 18011 43695 18045
rect 43649 17973 43695 18011
rect 43649 17939 43655 17973
rect 43689 17939 43695 17973
rect 43649 17901 43695 17939
rect 43649 17867 43655 17901
rect 43689 17867 43695 17901
rect 43649 17829 43695 17867
rect 43649 17795 43655 17829
rect 43689 17795 43695 17829
rect 43649 17757 43695 17795
rect 43649 17723 43655 17757
rect 43689 17723 43695 17757
rect 43649 17685 43695 17723
rect 43649 17651 43655 17685
rect 43689 17651 43695 17685
rect 43649 17613 43695 17651
rect 43649 17579 43655 17613
rect 43689 17579 43695 17613
rect 43649 17541 43695 17579
rect 43649 17507 43655 17541
rect 43689 17507 43695 17541
rect 43649 17469 43695 17507
rect 43649 17435 43655 17469
rect 43689 17435 43695 17469
rect 43649 17397 43695 17435
rect 44107 18621 44153 18637
rect 44107 18587 44113 18621
rect 44147 18587 44153 18621
rect 44107 18549 44153 18587
rect 44107 18515 44113 18549
rect 44147 18515 44153 18549
rect 44107 18477 44153 18515
rect 44107 18443 44113 18477
rect 44147 18443 44153 18477
rect 44107 18405 44153 18443
rect 44107 18371 44113 18405
rect 44147 18371 44153 18405
rect 44107 18333 44153 18371
rect 44107 18299 44113 18333
rect 44147 18299 44153 18333
rect 44107 18261 44153 18299
rect 44107 18227 44113 18261
rect 44147 18227 44153 18261
rect 44107 18189 44153 18227
rect 44107 18155 44113 18189
rect 44147 18155 44153 18189
rect 44107 18117 44153 18155
rect 44107 18083 44113 18117
rect 44147 18083 44153 18117
rect 44107 18045 44153 18083
rect 44107 18011 44113 18045
rect 44147 18011 44153 18045
rect 44107 17973 44153 18011
rect 44107 17939 44113 17973
rect 44147 17939 44153 17973
rect 44107 17901 44153 17939
rect 44107 17867 44113 17901
rect 44147 17867 44153 17901
rect 44107 17829 44153 17867
rect 44107 17795 44113 17829
rect 44147 17795 44153 17829
rect 44107 17757 44153 17795
rect 44107 17723 44113 17757
rect 44147 17723 44153 17757
rect 44107 17685 44153 17723
rect 44107 17651 44113 17685
rect 44147 17651 44153 17685
rect 44107 17613 44153 17651
rect 44107 17579 44113 17613
rect 44147 17579 44153 17613
rect 44107 17541 44153 17579
rect 44107 17507 44113 17541
rect 44147 17507 44153 17541
rect 44107 17469 44153 17507
rect 44107 17435 44113 17469
rect 44147 17435 44153 17469
rect 43649 17363 43655 17397
rect 43689 17363 43695 17397
rect 43649 17347 43695 17363
rect 43990 17348 43996 17400
rect 44048 17388 44054 17400
rect 44107 17397 44153 17435
rect 44107 17388 44113 17397
rect 44048 17363 44113 17388
rect 44147 17363 44153 17397
rect 44048 17360 44153 17363
rect 44048 17348 44054 17360
rect 44107 17347 44153 17360
rect 44565 18621 44611 18637
rect 44565 18587 44571 18621
rect 44605 18587 44611 18621
rect 44565 18549 44611 18587
rect 44565 18515 44571 18549
rect 44605 18515 44611 18549
rect 44565 18477 44611 18515
rect 44565 18443 44571 18477
rect 44605 18443 44611 18477
rect 44565 18405 44611 18443
rect 44565 18371 44571 18405
rect 44605 18371 44611 18405
rect 44565 18333 44611 18371
rect 44565 18299 44571 18333
rect 44605 18299 44611 18333
rect 44565 18261 44611 18299
rect 44565 18227 44571 18261
rect 44605 18227 44611 18261
rect 44565 18189 44611 18227
rect 44565 18155 44571 18189
rect 44605 18155 44611 18189
rect 44565 18117 44611 18155
rect 44565 18083 44571 18117
rect 44605 18083 44611 18117
rect 44565 18045 44611 18083
rect 44565 18011 44571 18045
rect 44605 18011 44611 18045
rect 44565 17973 44611 18011
rect 44565 17939 44571 17973
rect 44605 17939 44611 17973
rect 44565 17901 44611 17939
rect 44565 17867 44571 17901
rect 44605 17867 44611 17901
rect 44565 17829 44611 17867
rect 44565 17795 44571 17829
rect 44605 17795 44611 17829
rect 44565 17757 44611 17795
rect 44565 17723 44571 17757
rect 44605 17723 44611 17757
rect 44565 17685 44611 17723
rect 44565 17651 44571 17685
rect 44605 17651 44611 17685
rect 44565 17613 44611 17651
rect 44565 17579 44571 17613
rect 44605 17579 44611 17613
rect 44565 17541 44611 17579
rect 44565 17507 44571 17541
rect 44605 17507 44611 17541
rect 44565 17469 44611 17507
rect 44565 17435 44571 17469
rect 44605 17435 44611 17469
rect 44565 17397 44611 17435
rect 44565 17363 44571 17397
rect 44605 17363 44611 17397
rect 44565 17347 44611 17363
rect 45023 18621 45069 18637
rect 45023 18587 45029 18621
rect 45063 18587 45069 18621
rect 45023 18549 45069 18587
rect 45023 18515 45029 18549
rect 45063 18515 45069 18549
rect 45023 18477 45069 18515
rect 45023 18443 45029 18477
rect 45063 18443 45069 18477
rect 45023 18405 45069 18443
rect 45023 18371 45029 18405
rect 45063 18371 45069 18405
rect 45023 18333 45069 18371
rect 45023 18299 45029 18333
rect 45063 18299 45069 18333
rect 45023 18261 45069 18299
rect 45023 18227 45029 18261
rect 45063 18227 45069 18261
rect 45023 18189 45069 18227
rect 45023 18155 45029 18189
rect 45063 18155 45069 18189
rect 45023 18117 45069 18155
rect 45023 18083 45029 18117
rect 45063 18083 45069 18117
rect 45023 18045 45069 18083
rect 45023 18011 45029 18045
rect 45063 18011 45069 18045
rect 45023 17973 45069 18011
rect 45023 17939 45029 17973
rect 45063 17939 45069 17973
rect 45023 17901 45069 17939
rect 45023 17867 45029 17901
rect 45063 17867 45069 17901
rect 45023 17829 45069 17867
rect 45023 17795 45029 17829
rect 45063 17795 45069 17829
rect 45023 17757 45069 17795
rect 45023 17723 45029 17757
rect 45063 17723 45069 17757
rect 45023 17685 45069 17723
rect 45023 17651 45029 17685
rect 45063 17651 45069 17685
rect 45023 17613 45069 17651
rect 45023 17579 45029 17613
rect 45063 17579 45069 17613
rect 45023 17541 45069 17579
rect 45023 17507 45029 17541
rect 45063 17507 45069 17541
rect 45023 17469 45069 17507
rect 45023 17435 45029 17469
rect 45063 17435 45069 17469
rect 45023 17397 45069 17435
rect 45023 17363 45029 17397
rect 45063 17363 45069 17397
rect 45023 17347 45069 17363
rect 45481 18621 45527 18637
rect 45481 18587 45487 18621
rect 45521 18587 45527 18621
rect 45481 18549 45527 18587
rect 45481 18515 45487 18549
rect 45521 18515 45527 18549
rect 45481 18477 45527 18515
rect 45481 18443 45487 18477
rect 45521 18443 45527 18477
rect 45481 18405 45527 18443
rect 45481 18371 45487 18405
rect 45521 18371 45527 18405
rect 45481 18333 45527 18371
rect 45481 18299 45487 18333
rect 45521 18299 45527 18333
rect 45481 18261 45527 18299
rect 45481 18227 45487 18261
rect 45521 18227 45527 18261
rect 45481 18189 45527 18227
rect 45481 18155 45487 18189
rect 45521 18155 45527 18189
rect 45481 18117 45527 18155
rect 45481 18083 45487 18117
rect 45521 18083 45527 18117
rect 45481 18045 45527 18083
rect 45481 18011 45487 18045
rect 45521 18011 45527 18045
rect 45481 17973 45527 18011
rect 45481 17939 45487 17973
rect 45521 17939 45527 17973
rect 45481 17901 45527 17939
rect 45481 17867 45487 17901
rect 45521 17867 45527 17901
rect 45481 17829 45527 17867
rect 45481 17795 45487 17829
rect 45521 17795 45527 17829
rect 45481 17757 45527 17795
rect 45481 17723 45487 17757
rect 45521 17723 45527 17757
rect 45481 17685 45527 17723
rect 45481 17651 45487 17685
rect 45521 17651 45527 17685
rect 45481 17613 45527 17651
rect 45481 17579 45487 17613
rect 45521 17579 45527 17613
rect 45481 17541 45527 17579
rect 45481 17507 45487 17541
rect 45521 17507 45527 17541
rect 45481 17469 45527 17507
rect 45481 17435 45487 17469
rect 45521 17435 45527 17469
rect 45481 17397 45527 17435
rect 45481 17363 45487 17397
rect 45521 17363 45527 17397
rect 45481 17347 45527 17363
rect 45939 18621 45985 18637
rect 45939 18587 45945 18621
rect 45979 18587 45985 18621
rect 45939 18549 45985 18587
rect 45939 18515 45945 18549
rect 45979 18515 45985 18549
rect 45939 18477 45985 18515
rect 45939 18443 45945 18477
rect 45979 18443 45985 18477
rect 45939 18405 45985 18443
rect 45939 18371 45945 18405
rect 45979 18371 45985 18405
rect 45939 18333 45985 18371
rect 45939 18299 45945 18333
rect 45979 18299 45985 18333
rect 45939 18261 45985 18299
rect 45939 18227 45945 18261
rect 45979 18227 45985 18261
rect 45939 18189 45985 18227
rect 45939 18155 45945 18189
rect 45979 18155 45985 18189
rect 45939 18117 45985 18155
rect 45939 18083 45945 18117
rect 45979 18083 45985 18117
rect 45939 18045 45985 18083
rect 45939 18011 45945 18045
rect 45979 18011 45985 18045
rect 45939 17973 45985 18011
rect 45939 17939 45945 17973
rect 45979 17939 45985 17973
rect 45939 17901 45985 17939
rect 45939 17867 45945 17901
rect 45979 17867 45985 17901
rect 45939 17829 45985 17867
rect 45939 17795 45945 17829
rect 45979 17795 45985 17829
rect 45939 17757 45985 17795
rect 45939 17723 45945 17757
rect 45979 17723 45985 17757
rect 45939 17685 45985 17723
rect 45939 17651 45945 17685
rect 45979 17651 45985 17685
rect 45939 17613 45985 17651
rect 45939 17579 45945 17613
rect 45979 17579 45985 17613
rect 45939 17541 45985 17579
rect 45939 17507 45945 17541
rect 45979 17507 45985 17541
rect 45939 17469 45985 17507
rect 45939 17435 45945 17469
rect 45979 17435 45985 17469
rect 45939 17397 45985 17435
rect 45939 17363 45945 17397
rect 45979 17363 45985 17397
rect 45939 17347 45985 17363
rect 46397 18621 46443 18637
rect 46397 18587 46403 18621
rect 46437 18587 46443 18621
rect 46397 18549 46443 18587
rect 46397 18515 46403 18549
rect 46437 18515 46443 18549
rect 46397 18477 46443 18515
rect 46397 18443 46403 18477
rect 46437 18443 46443 18477
rect 46397 18405 46443 18443
rect 46397 18371 46403 18405
rect 46437 18371 46443 18405
rect 46397 18333 46443 18371
rect 46397 18299 46403 18333
rect 46437 18299 46443 18333
rect 46397 18261 46443 18299
rect 46397 18227 46403 18261
rect 46437 18227 46443 18261
rect 46397 18189 46443 18227
rect 46397 18155 46403 18189
rect 46437 18155 46443 18189
rect 46397 18117 46443 18155
rect 46397 18083 46403 18117
rect 46437 18083 46443 18117
rect 46397 18045 46443 18083
rect 46397 18011 46403 18045
rect 46437 18011 46443 18045
rect 46397 17973 46443 18011
rect 46397 17939 46403 17973
rect 46437 17939 46443 17973
rect 46397 17901 46443 17939
rect 46397 17867 46403 17901
rect 46437 17867 46443 17901
rect 46397 17829 46443 17867
rect 46397 17795 46403 17829
rect 46437 17795 46443 17829
rect 46397 17757 46443 17795
rect 46397 17723 46403 17757
rect 46437 17723 46443 17757
rect 46397 17685 46443 17723
rect 46397 17651 46403 17685
rect 46437 17651 46443 17685
rect 46397 17613 46443 17651
rect 46397 17579 46403 17613
rect 46437 17579 46443 17613
rect 46397 17541 46443 17579
rect 46397 17507 46403 17541
rect 46437 17507 46443 17541
rect 46397 17469 46443 17507
rect 46397 17435 46403 17469
rect 46437 17435 46443 17469
rect 46397 17397 46443 17435
rect 46397 17363 46403 17397
rect 46437 17363 46443 17397
rect 46397 17347 46443 17363
rect 46855 18621 46901 18637
rect 46855 18587 46861 18621
rect 46895 18587 46901 18621
rect 46855 18549 46901 18587
rect 46855 18515 46861 18549
rect 46895 18515 46901 18549
rect 46855 18477 46901 18515
rect 46855 18443 46861 18477
rect 46895 18443 46901 18477
rect 46855 18405 46901 18443
rect 46855 18371 46861 18405
rect 46895 18371 46901 18405
rect 46855 18333 46901 18371
rect 46855 18299 46861 18333
rect 46895 18299 46901 18333
rect 46855 18261 46901 18299
rect 46855 18227 46861 18261
rect 46895 18227 46901 18261
rect 46855 18189 46901 18227
rect 46855 18155 46861 18189
rect 46895 18155 46901 18189
rect 46855 18117 46901 18155
rect 46855 18083 46861 18117
rect 46895 18083 46901 18117
rect 46855 18045 46901 18083
rect 46855 18011 46861 18045
rect 46895 18011 46901 18045
rect 46855 17973 46901 18011
rect 46855 17939 46861 17973
rect 46895 17939 46901 17973
rect 46855 17901 46901 17939
rect 46855 17867 46861 17901
rect 46895 17867 46901 17901
rect 46855 17829 46901 17867
rect 46855 17795 46861 17829
rect 46895 17795 46901 17829
rect 46855 17757 46901 17795
rect 46855 17723 46861 17757
rect 46895 17723 46901 17757
rect 46855 17685 46901 17723
rect 46855 17651 46861 17685
rect 46895 17651 46901 17685
rect 46855 17613 46901 17651
rect 46855 17579 46861 17613
rect 46895 17579 46901 17613
rect 46855 17541 46901 17579
rect 46855 17507 46861 17541
rect 46895 17507 46901 17541
rect 46855 17469 46901 17507
rect 46855 17435 46861 17469
rect 46895 17435 46901 17469
rect 46855 17397 46901 17435
rect 46855 17363 46861 17397
rect 46895 17363 46901 17397
rect 46855 17347 46901 17363
rect 47313 18621 47359 18637
rect 47313 18587 47319 18621
rect 47353 18587 47359 18621
rect 47313 18549 47359 18587
rect 47313 18515 47319 18549
rect 47353 18515 47359 18549
rect 47313 18477 47359 18515
rect 47313 18443 47319 18477
rect 47353 18443 47359 18477
rect 47313 18405 47359 18443
rect 47313 18371 47319 18405
rect 47353 18371 47359 18405
rect 47313 18333 47359 18371
rect 47313 18299 47319 18333
rect 47353 18299 47359 18333
rect 47313 18261 47359 18299
rect 47313 18227 47319 18261
rect 47353 18227 47359 18261
rect 47313 18189 47359 18227
rect 47313 18155 47319 18189
rect 47353 18155 47359 18189
rect 47313 18117 47359 18155
rect 47313 18083 47319 18117
rect 47353 18083 47359 18117
rect 47313 18045 47359 18083
rect 47313 18011 47319 18045
rect 47353 18011 47359 18045
rect 47313 17973 47359 18011
rect 47313 17939 47319 17973
rect 47353 17939 47359 17973
rect 47313 17901 47359 17939
rect 47313 17867 47319 17901
rect 47353 17867 47359 17901
rect 47313 17829 47359 17867
rect 47313 17795 47319 17829
rect 47353 17795 47359 17829
rect 47313 17757 47359 17795
rect 47313 17723 47319 17757
rect 47353 17723 47359 17757
rect 47313 17685 47359 17723
rect 47313 17651 47319 17685
rect 47353 17651 47359 17685
rect 47313 17613 47359 17651
rect 47313 17579 47319 17613
rect 47353 17579 47359 17613
rect 47313 17541 47359 17579
rect 47313 17507 47319 17541
rect 47353 17507 47359 17541
rect 47313 17469 47359 17507
rect 47313 17435 47319 17469
rect 47353 17435 47359 17469
rect 47313 17397 47359 17435
rect 47313 17363 47319 17397
rect 47353 17363 47359 17397
rect 47313 17347 47359 17363
rect 47771 18621 47817 18637
rect 47771 18587 47777 18621
rect 47811 18587 47817 18621
rect 47771 18549 47817 18587
rect 47771 18515 47777 18549
rect 47811 18515 47817 18549
rect 47771 18477 47817 18515
rect 47771 18443 47777 18477
rect 47811 18443 47817 18477
rect 47771 18405 47817 18443
rect 47771 18371 47777 18405
rect 47811 18371 47817 18405
rect 47771 18333 47817 18371
rect 47771 18299 47777 18333
rect 47811 18299 47817 18333
rect 47771 18261 47817 18299
rect 47771 18227 47777 18261
rect 47811 18227 47817 18261
rect 47771 18189 47817 18227
rect 47771 18155 47777 18189
rect 47811 18155 47817 18189
rect 47771 18117 47817 18155
rect 47771 18083 47777 18117
rect 47811 18083 47817 18117
rect 47771 18045 47817 18083
rect 47771 18011 47777 18045
rect 47811 18011 47817 18045
rect 47771 17973 47817 18011
rect 47771 17939 47777 17973
rect 47811 17939 47817 17973
rect 47771 17901 47817 17939
rect 47771 17867 47777 17901
rect 47811 17867 47817 17901
rect 47771 17829 47817 17867
rect 47771 17795 47777 17829
rect 47811 17795 47817 17829
rect 47771 17757 47817 17795
rect 47771 17723 47777 17757
rect 47811 17723 47817 17757
rect 47771 17685 47817 17723
rect 47771 17651 47777 17685
rect 47811 17651 47817 17685
rect 47771 17613 47817 17651
rect 47771 17579 47777 17613
rect 47811 17579 47817 17613
rect 47771 17541 47817 17579
rect 47771 17507 47777 17541
rect 47811 17507 47817 17541
rect 47771 17469 47817 17507
rect 47771 17435 47777 17469
rect 47811 17435 47817 17469
rect 47771 17397 47817 17435
rect 47771 17363 47777 17397
rect 47811 17363 47817 17397
rect 47771 17347 47817 17363
rect 48229 18621 48275 18637
rect 48229 18587 48235 18621
rect 48269 18587 48275 18621
rect 48229 18549 48275 18587
rect 48229 18515 48235 18549
rect 48269 18515 48275 18549
rect 48229 18477 48275 18515
rect 48229 18443 48235 18477
rect 48269 18443 48275 18477
rect 48229 18405 48275 18443
rect 48229 18371 48235 18405
rect 48269 18371 48275 18405
rect 48229 18333 48275 18371
rect 48229 18299 48235 18333
rect 48269 18299 48275 18333
rect 48229 18261 48275 18299
rect 48229 18227 48235 18261
rect 48269 18227 48275 18261
rect 48229 18189 48275 18227
rect 48229 18155 48235 18189
rect 48269 18155 48275 18189
rect 48229 18117 48275 18155
rect 48229 18083 48235 18117
rect 48269 18083 48275 18117
rect 48229 18045 48275 18083
rect 48229 18011 48235 18045
rect 48269 18011 48275 18045
rect 48229 17973 48275 18011
rect 48229 17939 48235 17973
rect 48269 17939 48275 17973
rect 48229 17901 48275 17939
rect 48229 17867 48235 17901
rect 48269 17867 48275 17901
rect 48229 17829 48275 17867
rect 48229 17795 48235 17829
rect 48269 17795 48275 17829
rect 48229 17757 48275 17795
rect 48229 17723 48235 17757
rect 48269 17723 48275 17757
rect 48229 17685 48275 17723
rect 48229 17651 48235 17685
rect 48269 17651 48275 17685
rect 48229 17613 48275 17651
rect 48229 17579 48235 17613
rect 48269 17579 48275 17613
rect 48229 17541 48275 17579
rect 48229 17507 48235 17541
rect 48269 17507 48275 17541
rect 48229 17469 48275 17507
rect 48229 17435 48235 17469
rect 48269 17435 48275 17469
rect 48229 17397 48275 17435
rect 48229 17363 48235 17397
rect 48269 17363 48275 17397
rect 48229 17347 48275 17363
rect 48687 18621 48733 18637
rect 48687 18587 48693 18621
rect 48727 18587 48733 18621
rect 48687 18549 48733 18587
rect 48687 18515 48693 18549
rect 48727 18515 48733 18549
rect 48687 18477 48733 18515
rect 48687 18443 48693 18477
rect 48727 18443 48733 18477
rect 48687 18405 48733 18443
rect 48687 18371 48693 18405
rect 48727 18371 48733 18405
rect 48687 18333 48733 18371
rect 48687 18299 48693 18333
rect 48727 18299 48733 18333
rect 48687 18261 48733 18299
rect 48687 18227 48693 18261
rect 48727 18227 48733 18261
rect 48687 18189 48733 18227
rect 48687 18155 48693 18189
rect 48727 18155 48733 18189
rect 48687 18117 48733 18155
rect 48687 18083 48693 18117
rect 48727 18083 48733 18117
rect 48687 18045 48733 18083
rect 48687 18011 48693 18045
rect 48727 18011 48733 18045
rect 48687 17973 48733 18011
rect 48687 17939 48693 17973
rect 48727 17939 48733 17973
rect 48687 17901 48733 17939
rect 48687 17867 48693 17901
rect 48727 17867 48733 17901
rect 48687 17829 48733 17867
rect 48687 17795 48693 17829
rect 48727 17795 48733 17829
rect 48687 17757 48733 17795
rect 48687 17723 48693 17757
rect 48727 17723 48733 17757
rect 48687 17685 48733 17723
rect 48687 17651 48693 17685
rect 48727 17651 48733 17685
rect 48687 17613 48733 17651
rect 48687 17579 48693 17613
rect 48727 17579 48733 17613
rect 48687 17541 48733 17579
rect 48687 17507 48693 17541
rect 48727 17507 48733 17541
rect 48687 17469 48733 17507
rect 48687 17435 48693 17469
rect 48727 17435 48733 17469
rect 48687 17397 48733 17435
rect 48687 17363 48693 17397
rect 48727 17363 48733 17397
rect 48687 17347 48733 17363
rect 49145 18621 49191 18637
rect 49145 18587 49151 18621
rect 49185 18587 49191 18621
rect 49145 18549 49191 18587
rect 49145 18515 49151 18549
rect 49185 18515 49191 18549
rect 49145 18477 49191 18515
rect 49145 18443 49151 18477
rect 49185 18443 49191 18477
rect 49145 18405 49191 18443
rect 49145 18371 49151 18405
rect 49185 18371 49191 18405
rect 49145 18333 49191 18371
rect 49145 18299 49151 18333
rect 49185 18299 49191 18333
rect 49145 18261 49191 18299
rect 49145 18227 49151 18261
rect 49185 18227 49191 18261
rect 49145 18189 49191 18227
rect 49145 18155 49151 18189
rect 49185 18155 49191 18189
rect 49145 18117 49191 18155
rect 49145 18083 49151 18117
rect 49185 18083 49191 18117
rect 49145 18045 49191 18083
rect 49145 18011 49151 18045
rect 49185 18011 49191 18045
rect 49145 17973 49191 18011
rect 49145 17939 49151 17973
rect 49185 17939 49191 17973
rect 49145 17901 49191 17939
rect 49145 17867 49151 17901
rect 49185 17867 49191 17901
rect 49145 17829 49191 17867
rect 49145 17795 49151 17829
rect 49185 17795 49191 17829
rect 49145 17757 49191 17795
rect 49145 17723 49151 17757
rect 49185 17723 49191 17757
rect 49145 17685 49191 17723
rect 49145 17651 49151 17685
rect 49185 17651 49191 17685
rect 49145 17613 49191 17651
rect 49145 17579 49151 17613
rect 49185 17579 49191 17613
rect 49145 17541 49191 17579
rect 49145 17507 49151 17541
rect 49185 17507 49191 17541
rect 49145 17469 49191 17507
rect 49145 17435 49151 17469
rect 49185 17435 49191 17469
rect 49145 17397 49191 17435
rect 49145 17363 49151 17397
rect 49185 17363 49191 17397
rect 49145 17347 49191 17363
rect 49603 18621 49649 18637
rect 49603 18587 49609 18621
rect 49643 18587 49649 18621
rect 49603 18549 49649 18587
rect 49603 18515 49609 18549
rect 49643 18515 49649 18549
rect 49603 18477 49649 18515
rect 49603 18443 49609 18477
rect 49643 18443 49649 18477
rect 49603 18405 49649 18443
rect 49603 18371 49609 18405
rect 49643 18371 49649 18405
rect 49603 18333 49649 18371
rect 49603 18299 49609 18333
rect 49643 18299 49649 18333
rect 49603 18261 49649 18299
rect 49603 18227 49609 18261
rect 49643 18227 49649 18261
rect 49603 18189 49649 18227
rect 49603 18155 49609 18189
rect 49643 18155 49649 18189
rect 49603 18117 49649 18155
rect 49603 18083 49609 18117
rect 49643 18083 49649 18117
rect 49603 18045 49649 18083
rect 49603 18011 49609 18045
rect 49643 18011 49649 18045
rect 49603 17973 49649 18011
rect 49603 17939 49609 17973
rect 49643 17939 49649 17973
rect 49603 17901 49649 17939
rect 49603 17867 49609 17901
rect 49643 17867 49649 17901
rect 49603 17829 49649 17867
rect 49603 17795 49609 17829
rect 49643 17795 49649 17829
rect 49603 17757 49649 17795
rect 49603 17723 49609 17757
rect 49643 17723 49649 17757
rect 49603 17685 49649 17723
rect 49603 17651 49609 17685
rect 49643 17651 49649 17685
rect 49603 17613 49649 17651
rect 49603 17579 49609 17613
rect 49643 17579 49649 17613
rect 49603 17541 49649 17579
rect 49603 17507 49609 17541
rect 49643 17507 49649 17541
rect 49603 17469 49649 17507
rect 49603 17435 49609 17469
rect 49643 17435 49649 17469
rect 49603 17397 49649 17435
rect 49603 17363 49609 17397
rect 49643 17363 49649 17397
rect 49603 17347 49649 17363
rect 50061 18621 50107 18637
rect 50061 18587 50067 18621
rect 50101 18587 50107 18621
rect 50061 18549 50107 18587
rect 50061 18515 50067 18549
rect 50101 18515 50107 18549
rect 50061 18477 50107 18515
rect 50061 18443 50067 18477
rect 50101 18443 50107 18477
rect 50061 18405 50107 18443
rect 50061 18371 50067 18405
rect 50101 18371 50107 18405
rect 50061 18333 50107 18371
rect 50061 18299 50067 18333
rect 50101 18299 50107 18333
rect 50061 18261 50107 18299
rect 50061 18227 50067 18261
rect 50101 18227 50107 18261
rect 50061 18189 50107 18227
rect 50061 18155 50067 18189
rect 50101 18155 50107 18189
rect 50061 18117 50107 18155
rect 50061 18083 50067 18117
rect 50101 18083 50107 18117
rect 50061 18045 50107 18083
rect 50061 18011 50067 18045
rect 50101 18011 50107 18045
rect 50061 17973 50107 18011
rect 50061 17939 50067 17973
rect 50101 17939 50107 17973
rect 50061 17901 50107 17939
rect 50061 17867 50067 17901
rect 50101 17867 50107 17901
rect 50061 17829 50107 17867
rect 50061 17795 50067 17829
rect 50101 17795 50107 17829
rect 50061 17757 50107 17795
rect 50061 17723 50067 17757
rect 50101 17723 50107 17757
rect 50061 17685 50107 17723
rect 50061 17651 50067 17685
rect 50101 17651 50107 17685
rect 50061 17613 50107 17651
rect 50061 17579 50067 17613
rect 50101 17579 50107 17613
rect 50061 17541 50107 17579
rect 50061 17507 50067 17541
rect 50101 17507 50107 17541
rect 50061 17469 50107 17507
rect 50061 17435 50067 17469
rect 50101 17435 50107 17469
rect 50061 17397 50107 17435
rect 50061 17363 50067 17397
rect 50101 17363 50107 17397
rect 50061 17347 50107 17363
rect 50519 18621 50565 18637
rect 50519 18587 50525 18621
rect 50559 18587 50565 18621
rect 50519 18549 50565 18587
rect 50519 18515 50525 18549
rect 50559 18515 50565 18549
rect 50519 18477 50565 18515
rect 50519 18443 50525 18477
rect 50559 18443 50565 18477
rect 50519 18405 50565 18443
rect 50519 18371 50525 18405
rect 50559 18371 50565 18405
rect 50519 18333 50565 18371
rect 50519 18299 50525 18333
rect 50559 18299 50565 18333
rect 50519 18261 50565 18299
rect 50519 18227 50525 18261
rect 50559 18227 50565 18261
rect 50519 18189 50565 18227
rect 50519 18155 50525 18189
rect 50559 18155 50565 18189
rect 50519 18117 50565 18155
rect 50519 18083 50525 18117
rect 50559 18083 50565 18117
rect 50519 18045 50565 18083
rect 50519 18011 50525 18045
rect 50559 18011 50565 18045
rect 50519 17973 50565 18011
rect 50519 17939 50525 17973
rect 50559 17939 50565 17973
rect 50519 17901 50565 17939
rect 50519 17867 50525 17901
rect 50559 17867 50565 17901
rect 50519 17829 50565 17867
rect 50519 17795 50525 17829
rect 50559 17795 50565 17829
rect 50519 17757 50565 17795
rect 50519 17723 50525 17757
rect 50559 17723 50565 17757
rect 50519 17685 50565 17723
rect 50519 17651 50525 17685
rect 50559 17651 50565 17685
rect 50519 17613 50565 17651
rect 50519 17579 50525 17613
rect 50559 17579 50565 17613
rect 50519 17541 50565 17579
rect 50519 17507 50525 17541
rect 50559 17507 50565 17541
rect 50519 17469 50565 17507
rect 50519 17435 50525 17469
rect 50559 17435 50565 17469
rect 50519 17397 50565 17435
rect 50519 17363 50525 17397
rect 50559 17363 50565 17397
rect 50519 17347 50565 17363
rect 50977 18621 51023 18637
rect 50977 18587 50983 18621
rect 51017 18587 51023 18621
rect 50977 18549 51023 18587
rect 50977 18515 50983 18549
rect 51017 18515 51023 18549
rect 50977 18477 51023 18515
rect 50977 18443 50983 18477
rect 51017 18443 51023 18477
rect 50977 18405 51023 18443
rect 50977 18371 50983 18405
rect 51017 18371 51023 18405
rect 50977 18333 51023 18371
rect 50977 18299 50983 18333
rect 51017 18299 51023 18333
rect 50977 18261 51023 18299
rect 50977 18227 50983 18261
rect 51017 18227 51023 18261
rect 50977 18189 51023 18227
rect 50977 18155 50983 18189
rect 51017 18155 51023 18189
rect 50977 18117 51023 18155
rect 50977 18083 50983 18117
rect 51017 18083 51023 18117
rect 50977 18045 51023 18083
rect 50977 18011 50983 18045
rect 51017 18011 51023 18045
rect 50977 17973 51023 18011
rect 50977 17939 50983 17973
rect 51017 17939 51023 17973
rect 50977 17901 51023 17939
rect 50977 17867 50983 17901
rect 51017 17867 51023 17901
rect 50977 17829 51023 17867
rect 50977 17795 50983 17829
rect 51017 17795 51023 17829
rect 50977 17757 51023 17795
rect 50977 17723 50983 17757
rect 51017 17723 51023 17757
rect 50977 17685 51023 17723
rect 50977 17651 50983 17685
rect 51017 17651 51023 17685
rect 50977 17613 51023 17651
rect 50977 17579 50983 17613
rect 51017 17579 51023 17613
rect 50977 17541 51023 17579
rect 50977 17507 50983 17541
rect 51017 17507 51023 17541
rect 50977 17469 51023 17507
rect 50977 17435 50983 17469
rect 51017 17435 51023 17469
rect 50977 17397 51023 17435
rect 50977 17363 50983 17397
rect 51017 17363 51023 17397
rect 50977 17347 51023 17363
rect 51435 18621 51481 18637
rect 51435 18587 51441 18621
rect 51475 18587 51481 18621
rect 51435 18549 51481 18587
rect 51435 18515 51441 18549
rect 51475 18515 51481 18549
rect 51435 18477 51481 18515
rect 51435 18443 51441 18477
rect 51475 18443 51481 18477
rect 51435 18405 51481 18443
rect 51435 18371 51441 18405
rect 51475 18371 51481 18405
rect 51435 18333 51481 18371
rect 51435 18299 51441 18333
rect 51475 18299 51481 18333
rect 51435 18261 51481 18299
rect 51435 18227 51441 18261
rect 51475 18227 51481 18261
rect 51435 18189 51481 18227
rect 51435 18155 51441 18189
rect 51475 18155 51481 18189
rect 51435 18117 51481 18155
rect 51435 18083 51441 18117
rect 51475 18083 51481 18117
rect 51435 18045 51481 18083
rect 51435 18011 51441 18045
rect 51475 18011 51481 18045
rect 51435 17973 51481 18011
rect 51435 17939 51441 17973
rect 51475 17939 51481 17973
rect 51435 17901 51481 17939
rect 51435 17867 51441 17901
rect 51475 17867 51481 17901
rect 51435 17829 51481 17867
rect 51435 17795 51441 17829
rect 51475 17795 51481 17829
rect 51435 17757 51481 17795
rect 51435 17723 51441 17757
rect 51475 17723 51481 17757
rect 51435 17685 51481 17723
rect 51435 17651 51441 17685
rect 51475 17651 51481 17685
rect 51435 17613 51481 17651
rect 51435 17579 51441 17613
rect 51475 17579 51481 17613
rect 51435 17541 51481 17579
rect 51435 17507 51441 17541
rect 51475 17507 51481 17541
rect 51435 17469 51481 17507
rect 51435 17435 51441 17469
rect 51475 17435 51481 17469
rect 51435 17397 51481 17435
rect 51435 17363 51441 17397
rect 51475 17363 51481 17397
rect 51435 17347 51481 17363
rect 51893 18621 51939 18637
rect 51893 18587 51899 18621
rect 51933 18587 51939 18621
rect 51893 18549 51939 18587
rect 51893 18515 51899 18549
rect 51933 18515 51939 18549
rect 51893 18477 51939 18515
rect 51893 18443 51899 18477
rect 51933 18443 51939 18477
rect 51893 18405 51939 18443
rect 51893 18371 51899 18405
rect 51933 18371 51939 18405
rect 51893 18333 51939 18371
rect 51893 18299 51899 18333
rect 51933 18299 51939 18333
rect 51893 18261 51939 18299
rect 51893 18227 51899 18261
rect 51933 18227 51939 18261
rect 51893 18189 51939 18227
rect 51893 18155 51899 18189
rect 51933 18155 51939 18189
rect 51893 18117 51939 18155
rect 51893 18083 51899 18117
rect 51933 18083 51939 18117
rect 51893 18045 51939 18083
rect 51893 18011 51899 18045
rect 51933 18011 51939 18045
rect 51893 17973 51939 18011
rect 51893 17939 51899 17973
rect 51933 17939 51939 17973
rect 51893 17901 51939 17939
rect 51893 17867 51899 17901
rect 51933 17867 51939 17901
rect 51893 17829 51939 17867
rect 51893 17795 51899 17829
rect 51933 17795 51939 17829
rect 51893 17757 51939 17795
rect 51893 17723 51899 17757
rect 51933 17723 51939 17757
rect 51893 17685 51939 17723
rect 51893 17651 51899 17685
rect 51933 17651 51939 17685
rect 51893 17613 51939 17651
rect 51893 17579 51899 17613
rect 51933 17579 51939 17613
rect 51893 17541 51939 17579
rect 51893 17507 51899 17541
rect 51933 17507 51939 17541
rect 51893 17469 51939 17507
rect 51893 17435 51899 17469
rect 51933 17435 51939 17469
rect 51893 17397 51939 17435
rect 51893 17363 51899 17397
rect 51933 17363 51939 17397
rect 51893 17347 51939 17363
rect 52351 18621 52397 18637
rect 52351 18587 52357 18621
rect 52391 18587 52397 18621
rect 52351 18549 52397 18587
rect 52351 18515 52357 18549
rect 52391 18515 52397 18549
rect 52351 18477 52397 18515
rect 52351 18443 52357 18477
rect 52391 18443 52397 18477
rect 52351 18405 52397 18443
rect 52351 18371 52357 18405
rect 52391 18371 52397 18405
rect 52351 18333 52397 18371
rect 52351 18299 52357 18333
rect 52391 18299 52397 18333
rect 52351 18261 52397 18299
rect 52351 18227 52357 18261
rect 52391 18227 52397 18261
rect 52351 18189 52397 18227
rect 52351 18155 52357 18189
rect 52391 18155 52397 18189
rect 52351 18117 52397 18155
rect 52351 18083 52357 18117
rect 52391 18083 52397 18117
rect 52351 18045 52397 18083
rect 52351 18011 52357 18045
rect 52391 18011 52397 18045
rect 52351 17973 52397 18011
rect 52351 17939 52357 17973
rect 52391 17939 52397 17973
rect 52351 17901 52397 17939
rect 52351 17867 52357 17901
rect 52391 17867 52397 17901
rect 52351 17829 52397 17867
rect 52351 17795 52357 17829
rect 52391 17795 52397 17829
rect 52351 17757 52397 17795
rect 52351 17723 52357 17757
rect 52391 17723 52397 17757
rect 52351 17685 52397 17723
rect 52351 17651 52357 17685
rect 52391 17651 52397 17685
rect 52351 17613 52397 17651
rect 52351 17579 52357 17613
rect 52391 17579 52397 17613
rect 52351 17541 52397 17579
rect 52351 17507 52357 17541
rect 52391 17507 52397 17541
rect 52351 17469 52397 17507
rect 52351 17435 52357 17469
rect 52391 17435 52397 17469
rect 52351 17397 52397 17435
rect 52351 17363 52357 17397
rect 52391 17363 52397 17397
rect 52351 17347 52397 17363
rect 34330 17252 34336 17264
rect 34275 17224 34336 17252
rect 34330 17212 34336 17224
rect 34388 17212 34394 17264
rect 25406 17144 25412 17196
rect 25464 17144 25470 17196
rect 25409 17119 25421 17144
rect 25455 17119 25467 17144
rect 25409 17113 25467 17119
rect 900 17050 57536 17052
rect 900 16934 922 17050
rect 2510 17009 55926 17050
rect 2510 16975 25013 17009
rect 25047 16975 25413 17009
rect 25447 16975 25813 17009
rect 25847 16975 26213 17009
rect 26247 16975 26613 17009
rect 26647 16975 27013 17009
rect 27047 16975 27413 17009
rect 27447 16975 27813 17009
rect 27847 16975 28213 17009
rect 28247 16975 28613 17009
rect 28647 16975 29013 17009
rect 29047 16975 29413 17009
rect 29447 16975 29813 17009
rect 29847 16975 30213 17009
rect 30247 16975 30613 17009
rect 30647 16975 31013 17009
rect 31047 16975 31413 17009
rect 31447 16975 31813 17009
rect 31847 16975 32213 17009
rect 32247 16975 32613 17009
rect 32647 16975 33013 17009
rect 33047 16975 33413 17009
rect 33447 16975 33813 17009
rect 33847 16975 34213 17009
rect 34247 16975 34613 17009
rect 34647 16975 35013 17009
rect 35047 16975 35413 17009
rect 35447 16975 35813 17009
rect 35847 16975 36213 17009
rect 36247 16975 36613 17009
rect 36647 16975 37013 17009
rect 37047 16975 37413 17009
rect 37447 16975 37813 17009
rect 37847 16975 38213 17009
rect 38247 16975 38613 17009
rect 38647 16975 39013 17009
rect 39047 16975 39413 17009
rect 39447 16975 39813 17009
rect 39847 16975 40213 17009
rect 40247 16975 40613 17009
rect 40647 16975 41013 17009
rect 41047 16975 41413 17009
rect 41447 16975 41813 17009
rect 41847 16975 42213 17009
rect 42247 16975 42613 17009
rect 42647 16975 43013 17009
rect 43047 16975 43413 17009
rect 43447 16975 43813 17009
rect 43847 16975 44213 17009
rect 44247 16975 44613 17009
rect 44647 16975 45013 17009
rect 45047 16975 45413 17009
rect 45447 16975 45813 17009
rect 45847 16975 46213 17009
rect 46247 16975 46613 17009
rect 46647 16975 47013 17009
rect 47047 16975 47413 17009
rect 47447 16975 47813 17009
rect 47847 16975 48213 17009
rect 48247 16975 48613 17009
rect 48647 16975 49013 17009
rect 49047 16975 49413 17009
rect 49447 16975 49813 17009
rect 49847 16975 50213 17009
rect 50247 16975 50613 17009
rect 50647 16975 51013 17009
rect 51047 16975 51413 17009
rect 51447 16975 51813 17009
rect 51847 16975 52213 17009
rect 52247 16975 55926 17009
rect 2510 16934 55926 16975
rect 57514 16934 57536 17050
rect 900 16932 57536 16934
rect 3348 15170 55088 15172
rect 3348 15054 3370 15170
rect 4958 15129 53478 15170
rect 4958 15095 44045 15129
rect 44079 15095 44245 15129
rect 44279 15095 44445 15129
rect 44479 15095 44645 15129
rect 44679 15095 44845 15129
rect 44879 15095 45045 15129
rect 45079 15095 45245 15129
rect 45279 15095 45445 15129
rect 45479 15095 45645 15129
rect 45679 15095 45845 15129
rect 45879 15095 46045 15129
rect 46079 15095 46789 15129
rect 46823 15095 46989 15129
rect 47023 15095 47189 15129
rect 47223 15095 47389 15129
rect 47423 15095 47589 15129
rect 47623 15095 47789 15129
rect 47823 15095 47989 15129
rect 48023 15095 48189 15129
rect 48223 15095 48389 15129
rect 48423 15095 48589 15129
rect 48623 15095 48789 15129
rect 48823 15095 49533 15129
rect 49567 15095 49733 15129
rect 49767 15095 49933 15129
rect 49967 15095 50133 15129
rect 50167 15095 50333 15129
rect 50367 15095 50533 15129
rect 50567 15095 50733 15129
rect 50767 15095 50933 15129
rect 50967 15095 51133 15129
rect 51167 15095 51333 15129
rect 51367 15095 51533 15129
rect 51567 15095 53478 15129
rect 4958 15054 53478 15095
rect 55066 15054 55088 15170
rect 3348 15052 55088 15054
rect 49050 15008 49056 15020
rect 44192 14980 49056 15008
rect 44192 14873 44220 14980
rect 49050 14968 49056 14980
rect 49108 14968 49114 15020
rect 44376 14912 49096 14940
rect 44376 14884 44404 14912
rect 43873 14861 44283 14873
rect 43873 14323 43881 14861
rect 44275 14323 44283 14861
rect 44358 14832 44364 14884
rect 44416 14832 44422 14884
rect 45881 14861 46291 14873
rect 43873 14311 44283 14323
rect 45881 14323 45888 14861
rect 46282 14323 46291 14861
rect 45881 14311 46291 14323
rect 46617 14861 47027 14873
rect 46617 14323 46625 14861
rect 47019 14323 47027 14861
rect 46617 14311 46664 14323
rect 43873 13901 44283 13913
rect 43873 13363 43881 13901
rect 44275 13864 44283 13901
rect 45870 13901 46302 14311
rect 46658 14288 46664 14311
rect 46716 14311 47027 14323
rect 48625 14861 49035 14873
rect 48625 14323 48632 14861
rect 49026 14323 49035 14861
rect 49068 14872 49096 14912
rect 49361 14872 49771 14873
rect 49068 14861 49771 14872
rect 49068 14844 49369 14861
rect 48625 14311 49035 14323
rect 49361 14323 49369 14844
rect 49763 14323 49771 14861
rect 49361 14311 49771 14323
rect 51369 14861 51779 14873
rect 51369 14323 51376 14861
rect 51770 14323 51779 14861
rect 51369 14311 51779 14323
rect 46716 14288 46722 14311
rect 44324 13812 44330 13864
rect 44275 13363 44283 13812
rect 43873 13351 44283 13363
rect 45870 13363 45888 13901
rect 46282 13363 46302 13901
rect 45870 13347 46302 13363
rect 46617 13901 47027 13913
rect 46617 13363 46625 13901
rect 47019 13363 47027 13901
rect 46617 13351 46940 13363
rect 46934 13336 46940 13351
rect 46992 13351 47027 13363
rect 48614 13901 49046 14311
rect 48614 13363 48632 13901
rect 49026 13363 49046 13901
rect 46992 13336 46998 13351
rect 48614 13347 49046 13363
rect 49361 13901 49771 13913
rect 49361 13363 49369 13901
rect 49763 13363 49771 13901
rect 49361 13351 49516 13363
rect 49510 13336 49516 13351
rect 49568 13351 49771 13363
rect 51358 13901 51790 14311
rect 51358 13363 51376 13901
rect 51770 13363 51790 13901
rect 49568 13336 49574 13351
rect 51358 13347 51790 13363
rect 900 13290 57536 13292
rect 900 13174 922 13290
rect 2510 13249 55926 13290
rect 2510 13215 44045 13249
rect 44079 13215 44245 13249
rect 44279 13215 44445 13249
rect 44479 13215 44645 13249
rect 44679 13215 44845 13249
rect 44879 13215 45045 13249
rect 45079 13215 45245 13249
rect 45279 13215 45445 13249
rect 45479 13215 45645 13249
rect 45679 13215 45845 13249
rect 45879 13215 46045 13249
rect 46079 13215 46789 13249
rect 46823 13215 46989 13249
rect 47023 13215 47189 13249
rect 47223 13215 47389 13249
rect 47423 13215 47589 13249
rect 47623 13215 47789 13249
rect 47823 13215 47989 13249
rect 48023 13215 48189 13249
rect 48223 13215 48389 13249
rect 48423 13215 48589 13249
rect 48623 13215 48789 13249
rect 48823 13215 49533 13249
rect 49567 13215 49733 13249
rect 49767 13215 49933 13249
rect 49967 13215 50133 13249
rect 50167 13215 50333 13249
rect 50367 13215 50533 13249
rect 50567 13215 50733 13249
rect 50767 13215 50933 13249
rect 50967 13215 51133 13249
rect 51167 13215 51333 13249
rect 51367 13215 51533 13249
rect 51567 13215 55926 13249
rect 2510 13174 55926 13215
rect 57514 13174 57536 13290
rect 900 13172 57536 13174
rect 3348 11410 55088 11412
rect 3348 11294 3370 11410
rect 4958 11369 53478 11410
rect 4958 11335 43947 11369
rect 43981 11335 44147 11369
rect 44181 11335 44347 11369
rect 44381 11335 44547 11369
rect 44581 11335 44747 11369
rect 44781 11335 44947 11369
rect 44981 11335 45147 11369
rect 45181 11335 45347 11369
rect 45381 11335 45547 11369
rect 45581 11335 45747 11369
rect 45781 11335 45947 11369
rect 45981 11335 46691 11369
rect 46725 11335 46891 11369
rect 46925 11335 47091 11369
rect 47125 11335 47291 11369
rect 47325 11335 47491 11369
rect 47525 11335 47691 11369
rect 47725 11335 47891 11369
rect 47925 11335 48091 11369
rect 48125 11335 48291 11369
rect 48325 11335 48491 11369
rect 48525 11335 48691 11369
rect 48725 11335 49435 11369
rect 49469 11335 49635 11369
rect 49669 11335 49835 11369
rect 49869 11335 50035 11369
rect 50069 11335 50235 11369
rect 50269 11335 50435 11369
rect 50469 11335 50635 11369
rect 50669 11335 50835 11369
rect 50869 11335 51035 11369
rect 51069 11335 51235 11369
rect 51269 11335 51435 11369
rect 51469 11335 53478 11369
rect 4958 11294 53478 11335
rect 55066 11294 55088 11410
rect 3348 11292 55088 11294
rect 44726 11160 44732 11212
rect 44784 11200 44790 11212
rect 44784 11172 46336 11200
rect 44784 11160 44790 11172
rect 43775 11101 44185 11113
rect 43775 10563 43783 11101
rect 44177 10563 44185 11101
rect 43775 10551 44185 10563
rect 45783 11101 46193 11113
rect 45783 10563 45790 11101
rect 46184 10563 46193 11101
rect 46308 11064 46336 11172
rect 46934 11160 46940 11212
rect 46992 11200 46998 11212
rect 46992 11172 49004 11200
rect 46992 11160 46998 11172
rect 46519 11101 46929 11113
rect 46519 11064 46527 11101
rect 46308 11036 46527 11064
rect 45783 10551 46193 10563
rect 46519 10563 46527 11036
rect 46921 10563 46929 11101
rect 46519 10551 46929 10563
rect 48527 11101 48937 11113
rect 48527 10563 48534 11101
rect 48928 10563 48937 11101
rect 48976 11064 49004 11172
rect 49263 11101 49673 11113
rect 49263 11064 49271 11101
rect 48976 11036 49271 11064
rect 48527 10551 48937 10563
rect 49263 10563 49271 11036
rect 49665 10563 49673 11101
rect 49263 10551 49673 10563
rect 51271 11101 51681 11113
rect 51271 10563 51278 11101
rect 51672 10563 51681 11101
rect 51271 10551 51681 10563
rect 43775 10141 44185 10153
rect 43775 9603 43783 10141
rect 44177 9636 44185 10141
rect 45772 10141 46204 10551
rect 45646 9636 45652 9648
rect 44177 9608 45652 9636
rect 44177 9603 44185 9608
rect 43775 9591 44185 9603
rect 45646 9596 45652 9608
rect 45704 9596 45710 9648
rect 45772 9603 45790 10141
rect 46184 9603 46204 10141
rect 45772 9587 46204 9603
rect 46519 10141 46929 10153
rect 46519 9603 46527 10141
rect 46921 9603 46929 10141
rect 46519 9591 46929 9603
rect 48516 10141 48948 10551
rect 48516 9603 48534 10141
rect 48928 9603 48948 10141
rect 49263 10141 49673 10153
rect 49050 10072 49056 10124
rect 49108 10112 49114 10124
rect 49263 10112 49271 10141
rect 49108 10084 49271 10112
rect 49108 10072 49114 10084
rect 48516 9587 48948 9603
rect 49263 9603 49271 10084
rect 49665 9603 49673 10141
rect 49263 9591 49673 9603
rect 51260 10141 51692 10551
rect 51260 9603 51278 10141
rect 51672 9603 51692 10141
rect 51260 9587 51692 9603
rect 900 9530 57536 9532
rect 900 9414 922 9530
rect 2510 9489 55926 9530
rect 2510 9455 43947 9489
rect 43981 9455 44147 9489
rect 44181 9455 44347 9489
rect 44381 9455 44547 9489
rect 44581 9455 44747 9489
rect 44781 9455 44947 9489
rect 44981 9455 45147 9489
rect 45181 9455 45347 9489
rect 45381 9455 45547 9489
rect 45581 9455 45747 9489
rect 45781 9455 45947 9489
rect 45981 9455 46691 9489
rect 46725 9455 46891 9489
rect 46925 9455 47091 9489
rect 47125 9455 47291 9489
rect 47325 9455 47491 9489
rect 47525 9455 47691 9489
rect 47725 9455 47891 9489
rect 47925 9455 48091 9489
rect 48125 9455 48291 9489
rect 48325 9455 48491 9489
rect 48525 9455 48691 9489
rect 48725 9455 49435 9489
rect 49469 9455 49635 9489
rect 49669 9455 49835 9489
rect 49869 9455 50035 9489
rect 50069 9455 50235 9489
rect 50269 9455 50435 9489
rect 50469 9455 50635 9489
rect 50669 9455 50835 9489
rect 50869 9455 51035 9489
rect 51069 9455 51235 9489
rect 51269 9455 51435 9489
rect 51469 9455 55926 9489
rect 2510 9414 55926 9455
rect 57514 9414 57536 9530
rect 900 9412 57536 9414
rect 45646 9324 45652 9376
rect 45704 9364 45710 9376
rect 49878 9364 49884 9376
rect 45704 9336 49884 9364
rect 45704 9324 45710 9336
rect 49878 9324 49884 9336
rect 49936 9324 49942 9376
rect 3348 7650 55088 7652
rect 3348 7534 3370 7650
rect 4958 7609 53478 7650
rect 4958 7575 44731 7609
rect 44765 7575 44931 7609
rect 44965 7575 45131 7609
rect 45165 7575 45331 7609
rect 45365 7575 45531 7609
rect 45565 7575 45731 7609
rect 45765 7575 45931 7609
rect 45965 7575 46131 7609
rect 46165 7575 46331 7609
rect 46365 7575 46531 7609
rect 46565 7575 46731 7609
rect 46765 7575 47475 7609
rect 47509 7575 47675 7609
rect 47709 7575 47875 7609
rect 47909 7575 48075 7609
rect 48109 7575 48275 7609
rect 48309 7575 48475 7609
rect 48509 7575 48675 7609
rect 48709 7575 48875 7609
rect 48909 7575 49075 7609
rect 49109 7575 49275 7609
rect 49309 7575 49475 7609
rect 49509 7575 50219 7609
rect 50253 7575 50419 7609
rect 50453 7575 50619 7609
rect 50653 7575 50819 7609
rect 50853 7575 51019 7609
rect 51053 7575 51219 7609
rect 51253 7575 51419 7609
rect 51453 7575 51619 7609
rect 51653 7575 51819 7609
rect 51853 7575 52019 7609
rect 52053 7575 52219 7609
rect 52253 7575 53478 7609
rect 4958 7534 53478 7575
rect 55066 7534 55088 7650
rect 3348 7532 55088 7534
rect 49786 7460 49792 7472
rect 46492 7432 49792 7460
rect 44559 7341 44969 7353
rect 44559 6803 44567 7341
rect 44961 7324 44969 7341
rect 46492 7324 46520 7432
rect 49786 7420 49792 7432
rect 49844 7420 49850 7472
rect 44961 7296 46520 7324
rect 46567 7341 46977 7353
rect 44961 6803 44969 7296
rect 44559 6791 44969 6803
rect 46567 6803 46574 7341
rect 46968 6803 46977 7341
rect 46567 6791 46977 6803
rect 47303 7341 47713 7353
rect 47303 6803 47311 7341
rect 47705 7324 47713 7341
rect 49311 7341 49721 7353
rect 49142 7324 49148 7336
rect 47705 7296 49148 7324
rect 47705 6803 47713 7296
rect 49142 7284 49148 7296
rect 49200 7284 49206 7336
rect 47303 6791 47713 6803
rect 49311 6803 49318 7341
rect 49712 6803 49721 7341
rect 50047 7341 50457 7353
rect 49878 7284 49884 7336
rect 49936 7324 49942 7336
rect 50047 7324 50055 7341
rect 49936 7296 50055 7324
rect 49936 7284 49942 7296
rect 49311 6791 49721 6803
rect 50047 6803 50055 7296
rect 50449 6803 50457 7341
rect 50047 6791 50457 6803
rect 52055 7341 52465 7353
rect 52055 6803 52062 7341
rect 52456 6803 52465 7341
rect 52055 6791 52465 6803
rect 44559 6384 44969 6393
rect 44559 6381 44732 6384
rect 44784 6381 44969 6384
rect 44559 5843 44567 6381
rect 44961 5843 44969 6381
rect 44559 5831 44969 5843
rect 46556 6381 46988 6791
rect 46556 5843 46574 6381
rect 46968 5843 46988 6381
rect 46556 5827 46988 5843
rect 47303 6381 47713 6393
rect 47303 5843 47311 6381
rect 47705 5843 47713 6381
rect 47303 5831 47713 5843
rect 49300 6381 49732 6791
rect 49300 5843 49318 6381
rect 49712 5843 49732 6381
rect 49786 6332 49792 6384
rect 49844 6372 49850 6384
rect 50047 6381 50457 6393
rect 50047 6372 50055 6381
rect 49844 6344 50055 6372
rect 49844 6332 49850 6344
rect 47320 5772 47348 5831
rect 49300 5827 49732 5843
rect 50047 5843 50055 6344
rect 50449 5843 50457 6381
rect 50047 5831 50457 5843
rect 52044 6381 52476 6791
rect 52044 5843 52062 6381
rect 52456 5843 52476 6381
rect 52044 5827 52476 5843
rect 900 5770 57536 5772
rect 900 5654 922 5770
rect 2510 5729 55926 5770
rect 2510 5695 44731 5729
rect 44765 5695 44931 5729
rect 44965 5695 45131 5729
rect 45165 5695 45331 5729
rect 45365 5695 45531 5729
rect 45565 5695 45731 5729
rect 45765 5695 45931 5729
rect 45965 5695 46131 5729
rect 46165 5695 46331 5729
rect 46365 5695 46531 5729
rect 46565 5695 46731 5729
rect 46765 5695 47475 5729
rect 47509 5695 47675 5729
rect 47709 5695 47875 5729
rect 47909 5695 48075 5729
rect 48109 5695 48275 5729
rect 48309 5695 48475 5729
rect 48509 5695 48675 5729
rect 48709 5695 48875 5729
rect 48909 5695 49075 5729
rect 49109 5695 49275 5729
rect 49309 5695 49475 5729
rect 49509 5695 50219 5729
rect 50253 5695 50419 5729
rect 50453 5695 50619 5729
rect 50653 5695 50819 5729
rect 50853 5695 51019 5729
rect 51053 5695 51219 5729
rect 51253 5695 51419 5729
rect 51453 5695 51619 5729
rect 51653 5695 51819 5729
rect 51853 5695 52019 5729
rect 52053 5695 52219 5729
rect 52253 5695 55926 5729
rect 2510 5654 55926 5695
rect 57514 5654 57536 5770
rect 900 5652 57536 5654
rect 25498 4496 25504 4548
rect 25556 4536 25562 4548
rect 27522 4536 27528 4548
rect 25556 4508 27528 4536
rect 25556 4496 25562 4508
rect 27522 4496 27528 4508
rect 27580 4496 27586 4548
<< via1 >>
rect 922 50774 2510 50890
rect 55926 50774 57514 50890
rect 3370 48894 4958 49010
rect 53478 48894 55066 49010
rect 20996 48016 21048 48068
rect 19432 47268 19484 47320
rect 23756 47200 23808 47252
rect 48320 47472 48372 47524
rect 29460 47243 29512 47252
rect 29460 47209 29469 47243
rect 29469 47209 29503 47243
rect 29503 47209 29512 47243
rect 29460 47200 29512 47209
rect 922 47014 2510 47130
rect 17684 47064 17736 47116
rect 55926 47014 57514 47130
rect 3370 45134 4958 45250
rect 53478 45134 55066 45250
rect 14372 43707 14424 43716
rect 14372 43673 14381 43707
rect 14381 43673 14415 43707
rect 14415 43673 14424 43707
rect 14372 43664 14424 43673
rect 14556 43503 14608 43512
rect 14556 43469 14565 43503
rect 14565 43469 14599 43503
rect 14599 43469 14608 43503
rect 14556 43460 14608 43469
rect 22192 43664 22244 43716
rect 43260 44716 43312 44736
rect 43260 44684 43294 44716
rect 43294 44684 43312 44716
rect 44088 43800 44140 43852
rect 15016 43571 15068 43580
rect 15016 43537 15025 43571
rect 15025 43537 15059 43571
rect 15059 43537 15068 43571
rect 15016 43528 15068 43537
rect 29460 43469 29512 43478
rect 29460 43435 29469 43469
rect 29469 43435 29503 43469
rect 29503 43435 29512 43469
rect 29460 43426 29512 43435
rect 922 43254 2510 43370
rect 8300 43256 8352 43308
rect 43260 43256 43312 43308
rect 55926 43254 57514 43370
rect 3370 41374 4958 41490
rect 53478 41374 55066 41490
rect 28356 39924 28408 39976
rect 22192 39788 22244 39840
rect 23756 39788 23808 39840
rect 28080 39831 28132 39840
rect 28080 39797 28089 39831
rect 28089 39797 28123 39831
rect 28123 39797 28132 39831
rect 28080 39788 28132 39797
rect 28172 39720 28224 39772
rect 41972 41116 42024 41132
rect 41972 41082 42010 41116
rect 42010 41082 42024 41116
rect 41972 41080 42024 41082
rect 38568 40196 38620 40248
rect 41972 40922 41994 40928
rect 41994 40922 42024 40928
rect 41972 40876 42024 40922
rect 44088 40740 44140 40792
rect 42156 40218 42180 40248
rect 42180 40218 42208 40248
rect 42156 40196 42208 40218
rect 35808 40060 35860 40112
rect 48320 39856 48372 39908
rect 29460 39695 29512 39704
rect 29460 39661 29469 39695
rect 29469 39661 29503 39695
rect 29503 39661 29512 39695
rect 29460 39652 29512 39661
rect 922 39494 2510 39610
rect 15476 39516 15528 39568
rect 41972 39535 42001 39568
rect 42001 39535 42024 39568
rect 41972 39516 42024 39535
rect 55926 39494 57514 39610
rect 14372 38088 14424 38140
rect 25780 38020 25832 38072
rect 34428 37952 34480 38004
rect 35808 37952 35860 38004
rect 3370 37614 4958 37730
rect 33416 37612 33468 37664
rect 53478 37614 55066 37730
rect 12900 37136 12952 37188
rect 15568 36864 15620 36916
rect 16580 36883 16632 36916
rect 13912 35923 13964 35964
rect 13912 35912 13964 35923
rect 16580 36864 16632 36883
rect 22284 37476 22336 37528
rect 16212 36388 16264 36440
rect 22376 36864 22428 36916
rect 25780 37136 25832 37188
rect 22284 36388 22336 36440
rect 34428 37136 34480 37188
rect 29460 36932 29512 36984
rect 28080 36159 28132 36168
rect 28080 36125 28089 36159
rect 28089 36125 28123 36159
rect 28123 36125 28132 36159
rect 28080 36116 28132 36125
rect 41972 37162 41994 37188
rect 41994 37162 42024 37188
rect 41972 37136 42024 37162
rect 42156 36492 42208 36508
rect 42156 36458 42180 36492
rect 42180 36458 42208 36492
rect 42156 36456 42208 36458
rect 37556 36023 37565 36032
rect 37565 36023 37599 36032
rect 37599 36023 37608 36032
rect 37556 35980 37608 36023
rect 38568 35955 38620 35964
rect 38568 35921 38577 35955
rect 38577 35921 38611 35955
rect 38611 35921 38620 35955
rect 38568 35912 38620 35921
rect 922 35734 2510 35850
rect 41972 35809 42024 35828
rect 41972 35776 42001 35809
rect 42001 35776 42024 35809
rect 55926 35734 57514 35850
rect 3370 33854 4958 33970
rect 33416 33872 33468 33924
rect 53478 33854 55066 33970
rect 48688 33736 48740 33788
rect 19432 33600 19484 33652
rect 24492 33124 24544 33176
rect 41880 33562 41920 33584
rect 41920 33562 41932 33584
rect 41880 33532 41932 33562
rect 42156 33232 42208 33244
rect 42156 33198 42180 33232
rect 42180 33198 42208 33232
rect 42156 33192 42208 33198
rect 16580 32648 16632 32700
rect 42248 32698 42280 32700
rect 42280 32698 42300 32700
rect 42248 32648 42300 32698
rect 922 31974 2510 32090
rect 55926 31974 57514 32090
rect 3370 30094 4958 30210
rect 33416 30132 33468 30184
rect 53478 30094 55066 30210
rect 20904 29996 20956 30048
rect 22376 29996 22428 30048
rect 16672 29384 16724 29436
rect 19064 29384 19116 29436
rect 22192 29901 22244 29912
rect 22192 29860 22244 29901
rect 27436 29384 27488 29436
rect 18420 28908 18472 28960
rect 20904 28908 20956 28960
rect 21732 28908 21784 28960
rect 24492 28908 24544 28960
rect 42156 29676 42208 29708
rect 42156 29656 42174 29676
rect 42174 29656 42208 29676
rect 42248 29472 42300 29504
rect 42248 29452 42280 29472
rect 42280 29452 42300 29472
rect 48412 28908 48464 28960
rect 38568 28407 38620 28416
rect 38568 28373 38577 28407
rect 38577 28373 38611 28407
rect 38611 28373 38620 28407
rect 38568 28364 38620 28373
rect 922 28214 2510 28330
rect 42156 28255 42167 28280
rect 42167 28255 42201 28280
rect 42201 28255 42208 28280
rect 42156 28228 42208 28255
rect 55926 28214 57514 28330
rect 3370 26334 4958 26450
rect 33416 26392 33468 26444
rect 53478 26334 55066 26450
rect 39948 26188 40000 26240
rect 13912 25848 13964 25900
rect 22928 24624 22980 24676
rect 25412 25135 25430 25152
rect 25430 25135 25464 25152
rect 25412 25100 25464 25135
rect 29460 25712 29512 25764
rect 27528 24871 27580 24880
rect 27528 24837 27537 24871
rect 27537 24837 27571 24871
rect 27571 24837 27580 24871
rect 27528 24828 27580 24837
rect 37372 24643 37413 24676
rect 37413 24643 37424 24676
rect 37372 24624 37424 24643
rect 40132 25603 40157 25628
rect 40157 25603 40184 25628
rect 41420 26120 41472 26172
rect 46020 26188 46072 26240
rect 48504 26188 48556 26240
rect 40132 25576 40184 25603
rect 42708 25644 42760 25696
rect 48596 25603 48648 25628
rect 39948 25100 40000 25152
rect 42892 24643 42901 24676
rect 42901 24643 42944 24676
rect 42892 24624 42944 24643
rect 48596 25576 48648 25603
rect 46020 25100 46039 25152
rect 46039 25100 46072 25152
rect 48412 25100 48464 25152
rect 922 24454 2510 24570
rect 55926 24454 57514 24570
rect 38292 24148 38344 24200
rect 42892 24148 42944 24200
rect 30932 23400 30984 23452
rect 37372 23400 37424 23452
rect 3370 22574 4958 22690
rect 53478 22574 55066 22690
rect 34980 22448 35032 22500
rect 40132 22448 40184 22500
rect 42708 22448 42760 22500
rect 48504 22448 48556 22500
rect 22928 22312 22980 22364
rect 29092 21836 29144 21888
rect 30932 22312 30984 22364
rect 35072 21836 35124 21888
rect 38292 22312 38344 22364
rect 16672 21360 16724 21412
rect 27436 21360 27488 21412
rect 29736 21360 29788 21412
rect 34980 21360 35032 21412
rect 35716 21360 35768 21412
rect 41420 21360 41472 21412
rect 48596 21360 48648 21412
rect 922 20694 2510 20810
rect 55926 20694 57514 20810
rect 3370 18814 4958 18930
rect 53478 18814 55066 18930
rect 43996 17348 44048 17400
rect 34336 17255 34388 17264
rect 34336 17221 34345 17255
rect 34345 17221 34379 17255
rect 34379 17221 34388 17255
rect 34336 17212 34388 17221
rect 25412 17153 25464 17196
rect 25412 17144 25421 17153
rect 25421 17144 25455 17153
rect 25455 17144 25464 17153
rect 922 16934 2510 17050
rect 55926 16934 57514 17050
rect 3370 15054 4958 15170
rect 53478 15054 55066 15170
rect 49056 14968 49108 15020
rect 44364 14832 44416 14884
rect 46664 14323 46716 14340
rect 46664 14288 46716 14323
rect 44272 13812 44275 13864
rect 44275 13812 44324 13864
rect 46940 13363 46992 13388
rect 46940 13336 46992 13363
rect 49516 13363 49568 13388
rect 49516 13336 49568 13363
rect 922 13174 2510 13290
rect 55926 13174 57514 13290
rect 3370 11294 4958 11410
rect 53478 11294 55066 11410
rect 44732 11160 44784 11212
rect 43996 11024 44048 11076
rect 46940 11160 46992 11212
rect 45652 9596 45704 9648
rect 46664 10072 46716 10124
rect 49056 10072 49108 10124
rect 922 9414 2510 9530
rect 55926 9414 57514 9530
rect 45652 9324 45704 9376
rect 49884 9324 49936 9376
rect 3370 7534 4958 7650
rect 53478 7534 55066 7650
rect 49792 7420 49844 7472
rect 49148 7284 49200 7336
rect 49884 7284 49936 7336
rect 44732 6381 44784 6384
rect 44732 6332 44784 6381
rect 49792 6332 49844 6384
rect 922 5654 2510 5770
rect 55926 5654 57514 5770
rect 25504 4496 25556 4548
rect 27528 4496 27580 4548
<< metal2 >>
rect 900 50890 2532 50892
rect 900 50774 922 50890
rect 2510 50774 2532 50890
rect 900 50772 2532 50774
rect 55904 50890 57536 50892
rect 55904 50774 55926 50890
rect 57514 50774 57536 50890
rect 55904 50772 57536 50774
rect 3348 49010 4980 49012
rect 3348 48894 3370 49010
rect 4958 48894 4980 49010
rect 3348 48892 4980 48894
rect 53456 49010 55088 49012
rect 53456 48894 53478 49010
rect 55066 48894 55088 49010
rect 53456 48892 55088 48894
rect 5916 48710 6116 48722
rect 5916 48654 5948 48710
rect 6004 48654 6028 48710
rect 6084 48654 6116 48710
rect 5916 48642 6116 48654
rect 13364 48710 13564 48722
rect 13364 48654 13396 48710
rect 13452 48654 13476 48710
rect 13532 48654 13564 48710
rect 13364 48642 13564 48654
rect 20996 48068 21048 48074
rect 20996 48010 21048 48016
rect 19432 47320 19484 47326
rect 5938 47290 6098 47312
rect 5938 47234 5990 47290
rect 6046 47234 6098 47290
rect 5938 47212 6098 47234
rect 13386 47290 13546 47312
rect 13386 47234 13438 47290
rect 13494 47234 13546 47290
rect 19432 47262 19484 47268
rect 13386 47212 13546 47234
rect 17682 47132 17738 47141
rect 900 47130 2532 47132
rect 900 47014 922 47130
rect 2510 47014 2532 47130
rect 17682 47067 17684 47076
rect 17736 47067 17738 47076
rect 17684 47058 17736 47064
rect 17696 47044 17724 47058
rect 900 47012 2532 47014
rect 3348 45250 4980 45252
rect 3348 45134 3370 45250
rect 4958 45134 4980 45250
rect 3348 45132 4980 45134
rect 5916 44950 6116 44962
rect 5916 44894 5948 44950
rect 6004 44894 6028 44950
rect 6084 44894 6116 44950
rect 5916 44882 6116 44894
rect 15014 43838 15070 43847
rect 15014 43773 15070 43782
rect 14372 43716 14424 43722
rect 14372 43658 14424 43664
rect 5938 43530 6098 43552
rect 5938 43474 5990 43530
rect 6046 43474 6098 43530
rect 5938 43452 6098 43474
rect 900 43370 2532 43372
rect 900 43254 922 43370
rect 2510 43254 2532 43370
rect 8298 43350 8354 43359
rect 8298 43285 8300 43294
rect 900 43252 2532 43254
rect 8352 43285 8354 43294
rect 8300 43250 8352 43256
rect 3348 41490 4980 41492
rect 3348 41374 3370 41490
rect 4958 41374 4980 41490
rect 3348 41372 4980 41374
rect 6308 41190 6508 41202
rect 6308 41134 6340 41190
rect 6396 41134 6420 41190
rect 6476 41134 6508 41190
rect 6308 41122 6508 41134
rect 6330 39770 6490 39792
rect 6330 39714 6382 39770
rect 6438 39714 6490 39770
rect 6330 39692 6490 39714
rect 900 39610 2532 39612
rect 900 39494 922 39610
rect 2510 39494 2532 39610
rect 900 39492 2532 39494
rect 14384 38146 14412 43658
rect 15028 43586 15056 43773
rect 15016 43580 15068 43586
rect 15016 43522 15068 43528
rect 14556 43512 14608 43518
rect 14554 43472 14556 43481
rect 14608 43472 14610 43481
rect 14554 43407 14610 43416
rect 15128 41190 15328 41202
rect 15128 41134 15160 41190
rect 15216 41134 15240 41190
rect 15296 41134 15328 41190
rect 15128 41122 15328 41134
rect 15150 39770 15310 39792
rect 15150 39714 15202 39770
rect 15258 39714 15310 39770
rect 15150 39692 15310 39714
rect 15474 39690 15530 39699
rect 15474 39625 15530 39634
rect 15488 39574 15516 39625
rect 15476 39568 15528 39574
rect 15476 39510 15528 39516
rect 14372 38140 14424 38146
rect 14372 38082 14424 38088
rect 3348 37730 4980 37732
rect 3348 37614 3370 37730
rect 4958 37614 4980 37730
rect 3348 37612 4980 37614
rect 12898 37250 12954 37259
rect 12898 37188 12954 37194
rect 12898 37185 12900 37188
rect 12952 37185 12954 37188
rect 12900 37130 12952 37136
rect 15568 36916 15620 36922
rect 16580 36916 16632 36922
rect 15620 36876 16252 36904
rect 15568 36858 15620 36864
rect 16224 36446 16252 36876
rect 16580 36858 16632 36864
rect 16212 36440 16264 36446
rect 16212 36382 16264 36388
rect 13912 35964 13964 35970
rect 13912 35906 13964 35912
rect 900 35850 2532 35852
rect 900 35734 922 35850
rect 2510 35734 2532 35850
rect 900 35732 2532 35734
rect 3348 33970 4980 33972
rect 3348 33854 3370 33970
rect 4958 33854 4980 33970
rect 3348 33852 4980 33854
rect 900 32090 2532 32092
rect 900 31974 922 32090
rect 2510 31974 2532 32090
rect 900 31972 2532 31974
rect 3348 30210 4980 30212
rect 3348 30094 3370 30210
rect 4958 30094 4980 30210
rect 3348 30092 4980 30094
rect 900 28330 2532 28332
rect 900 28214 922 28330
rect 2510 28214 2532 28330
rect 900 28212 2532 28214
rect 3348 26450 4980 26452
rect 3348 26334 3370 26450
rect 4958 26334 4980 26450
rect 3348 26332 4980 26334
rect 13924 25906 13952 35906
rect 16592 32706 16620 36858
rect 19444 33658 19472 47262
rect 19432 33652 19484 33658
rect 19432 33594 19484 33600
rect 16580 32700 16632 32706
rect 16580 32642 16632 32648
rect 20904 30048 20956 30054
rect 20904 29990 20956 29996
rect 16672 29436 16724 29442
rect 19064 29436 19116 29442
rect 16672 29378 16724 29384
rect 18432 29396 19064 29424
rect 13912 25900 13964 25906
rect 13912 25842 13964 25848
rect 900 24570 2532 24572
rect 900 24454 922 24570
rect 2510 24454 2532 24570
rect 900 24452 2532 24454
rect 3348 22690 4980 22692
rect 3348 22574 3370 22690
rect 4958 22574 4980 22690
rect 3348 22572 4980 22574
rect 16684 21418 16712 29378
rect 18432 28966 18460 29396
rect 19064 29378 19116 29384
rect 20916 28966 20944 29990
rect 21008 29152 21036 48010
rect 48320 47524 48372 47530
rect 48320 47466 48372 47472
rect 23756 47252 23808 47258
rect 23756 47194 23808 47200
rect 29460 47252 29512 47258
rect 29460 47194 29512 47200
rect 22192 43716 22244 43722
rect 22192 43658 22244 43664
rect 22204 41407 22232 43658
rect 23768 43481 23796 47194
rect 29472 43484 29500 47194
rect 43260 44736 43312 44742
rect 43260 44678 43312 44684
rect 23754 43472 23810 43481
rect 29460 43478 29512 43484
rect 29460 43420 29512 43426
rect 23754 43407 23810 43416
rect 22190 41398 22246 41407
rect 22190 41333 22246 41342
rect 22204 39846 22232 41333
rect 23768 39846 23796 43407
rect 28356 39976 28408 39982
rect 28356 39918 28408 39924
rect 22192 39840 22244 39846
rect 22192 39782 22244 39788
rect 23756 39840 23808 39846
rect 23756 39782 23808 39788
rect 28080 39840 28132 39846
rect 28080 39782 28132 39788
rect 22204 29918 22232 39782
rect 25780 38072 25832 38078
rect 25780 38014 25832 38020
rect 22284 37528 22336 37534
rect 22284 37470 22336 37476
rect 22296 36446 22324 37470
rect 25792 37194 25820 38014
rect 25780 37188 25832 37194
rect 25780 37130 25832 37136
rect 22376 36916 22428 36922
rect 22376 36858 22428 36864
rect 22284 36440 22336 36446
rect 22284 36382 22336 36388
rect 22388 30054 22416 36858
rect 28092 36174 28120 39782
rect 28172 39772 28224 39778
rect 28368 39760 28396 39918
rect 28224 39732 28396 39760
rect 28172 39714 28224 39720
rect 29472 39710 29500 43420
rect 43272 43314 43300 44678
rect 44088 43852 44140 43858
rect 44088 43794 44140 43800
rect 43260 43308 43312 43314
rect 43260 43250 43312 43256
rect 41972 41132 42024 41138
rect 41972 41074 42024 41080
rect 41984 40934 42012 41074
rect 41972 40928 42024 40934
rect 41972 40870 42024 40876
rect 38568 40248 38620 40254
rect 38568 40190 38620 40196
rect 35808 40112 35860 40118
rect 35808 40054 35860 40060
rect 29460 39704 29512 39710
rect 29460 39646 29512 39652
rect 29472 37015 29500 39646
rect 35820 38010 35848 40054
rect 34428 38004 34480 38010
rect 34428 37946 34480 37952
rect 35808 38004 35860 38010
rect 35808 37946 35860 37952
rect 33416 37664 33468 37670
rect 33414 37616 33416 37625
rect 33468 37616 33470 37625
rect 33414 37551 33470 37560
rect 29926 37430 30126 37442
rect 29926 37374 29958 37430
rect 30014 37374 30038 37430
rect 30094 37374 30126 37430
rect 29926 37362 30126 37374
rect 34440 37194 34468 37946
rect 34428 37188 34480 37194
rect 34428 37130 34480 37136
rect 29458 37006 29514 37015
rect 29458 36941 29460 36950
rect 29512 36941 29514 36950
rect 29460 36926 29512 36932
rect 29472 36918 29500 36926
rect 28080 36168 28132 36174
rect 28080 36110 28132 36116
rect 37554 36032 37610 36039
rect 29948 36010 30108 36032
rect 29948 35954 30000 36010
rect 30056 35954 30108 36010
rect 37554 36030 37556 36032
rect 37608 36030 37610 36032
rect 37554 35965 37610 35974
rect 38580 35970 38608 40190
rect 41984 39574 42012 40870
rect 44100 40798 44128 43794
rect 44088 40792 44140 40798
rect 44088 40734 44140 40740
rect 42156 40248 42208 40254
rect 42156 40190 42208 40196
rect 41972 39568 42024 39574
rect 41972 39510 42024 39516
rect 41972 37188 42024 37194
rect 41972 37130 42024 37136
rect 29948 35932 30108 35954
rect 37568 35942 37596 35965
rect 38568 35964 38620 35970
rect 38568 35906 38620 35912
rect 33414 33924 33470 33930
rect 33414 33872 33416 33924
rect 33468 33872 33470 33924
rect 33414 33834 33470 33872
rect 33414 33769 33470 33778
rect 26202 33670 26402 33682
rect 26202 33614 26234 33670
rect 26290 33614 26314 33670
rect 26370 33614 26402 33670
rect 26202 33602 26402 33614
rect 33650 33670 33850 33682
rect 33650 33614 33682 33670
rect 33738 33614 33762 33670
rect 33818 33614 33850 33670
rect 33650 33602 33850 33614
rect 24492 33176 24544 33182
rect 24492 33118 24544 33124
rect 22376 30048 22428 30054
rect 22376 29990 22428 29996
rect 22192 29912 22244 29918
rect 22192 29854 22244 29860
rect 21008 29124 21772 29152
rect 21744 28966 21772 29124
rect 24504 28966 24532 33118
rect 26224 32250 26384 32272
rect 26224 32194 26276 32250
rect 26332 32194 26384 32250
rect 26224 32172 26384 32194
rect 33672 32250 33832 32272
rect 33672 32194 33724 32250
rect 33780 32194 33832 32250
rect 33672 32172 33832 32194
rect 33416 30184 33468 30190
rect 33414 30174 33416 30183
rect 33468 30174 33470 30183
rect 33414 30109 33470 30118
rect 33428 30093 33456 30109
rect 29926 29910 30126 29922
rect 29926 29854 29958 29910
rect 30014 29854 30038 29910
rect 30094 29854 30126 29910
rect 29926 29842 30126 29854
rect 27436 29436 27488 29442
rect 27436 29378 27488 29384
rect 18420 28960 18472 28966
rect 18420 28902 18472 28908
rect 20904 28960 20956 28966
rect 20904 28902 20956 28908
rect 21732 28960 21784 28966
rect 21732 28902 21784 28908
rect 24492 28960 24544 28966
rect 24492 28902 24544 28908
rect 25412 25152 25464 25158
rect 25412 25094 25464 25100
rect 22928 24676 22980 24682
rect 22928 24618 22980 24624
rect 22940 22370 22968 24618
rect 22928 22364 22980 22370
rect 22928 22306 22980 22312
rect 16672 21412 16724 21418
rect 16672 21354 16724 21360
rect 900 20810 2532 20812
rect 900 20694 922 20810
rect 2510 20694 2532 20810
rect 900 20692 2532 20694
rect 3348 18930 4980 18932
rect 3348 18814 3370 18930
rect 4958 18814 4980 18930
rect 3348 18812 4980 18814
rect 25424 17202 25452 25094
rect 27448 21418 27476 29378
rect 29948 28490 30108 28512
rect 29948 28434 30000 28490
rect 30056 28434 30108 28490
rect 29948 28412 30108 28434
rect 38580 28422 38608 35906
rect 41984 35834 42012 37130
rect 42168 36514 42196 40190
rect 48332 39914 48360 47466
rect 55904 47130 57536 47132
rect 55904 47014 55926 47130
rect 57514 47014 57536 47130
rect 55904 47012 57536 47014
rect 53456 45250 55088 45252
rect 53456 45134 53478 45250
rect 55066 45134 55088 45250
rect 53456 45132 55088 45134
rect 55904 43370 57536 43372
rect 55904 43254 55926 43370
rect 57514 43254 57536 43370
rect 55904 43252 57536 43254
rect 53456 41490 55088 41492
rect 53456 41374 53478 41490
rect 55066 41374 55088 41490
rect 53456 41372 55088 41374
rect 48320 39908 48372 39914
rect 48320 39850 48372 39856
rect 48332 37176 48360 39850
rect 55904 39610 57536 39612
rect 55904 39494 55926 39610
rect 57514 39494 57536 39610
rect 55904 39492 57536 39494
rect 53456 37730 55088 37732
rect 53456 37614 53478 37730
rect 55066 37614 55088 37730
rect 53456 37612 55088 37614
rect 48332 37148 48544 37176
rect 42156 36508 42208 36514
rect 42156 36450 42208 36456
rect 41972 35828 42024 35834
rect 41972 35770 42024 35776
rect 41984 33776 42012 35770
rect 41892 33748 42012 33776
rect 41892 33590 41920 33748
rect 41880 33584 41932 33590
rect 41880 33526 41932 33532
rect 42168 33250 42196 36450
rect 48516 33776 48544 37148
rect 55904 35850 57536 35852
rect 55904 35734 55926 35850
rect 57514 35734 57536 35850
rect 55904 35732 57536 35734
rect 53456 33970 55088 33972
rect 53456 33854 53478 33970
rect 55066 33854 55088 33970
rect 53456 33852 55088 33854
rect 48688 33788 48740 33794
rect 48516 33748 48688 33776
rect 42156 33244 42208 33250
rect 42156 33186 42208 33192
rect 42248 32700 42300 32706
rect 42248 32642 42300 32648
rect 42156 29708 42208 29714
rect 42156 29650 42208 29656
rect 38568 28416 38620 28422
rect 38568 28358 38620 28364
rect 42168 28286 42196 29650
rect 42260 29510 42288 32642
rect 42248 29504 42300 29510
rect 42248 29446 42300 29452
rect 48412 28960 48464 28966
rect 48412 28902 48464 28908
rect 42156 28280 42208 28286
rect 42156 28222 42208 28228
rect 33416 26444 33468 26450
rect 33414 26392 33416 26401
rect 33468 26392 33470 26401
rect 33414 26327 33470 26336
rect 39948 26240 40000 26246
rect 39948 26182 40000 26188
rect 46020 26240 46072 26246
rect 46020 26182 46072 26188
rect 29926 26150 30126 26162
rect 29926 26094 29958 26150
rect 30014 26094 30038 26150
rect 30094 26094 30126 26150
rect 29926 26082 30126 26094
rect 29458 25782 29514 25791
rect 29458 25717 29460 25726
rect 29512 25717 29514 25726
rect 29460 25706 29512 25712
rect 29472 25694 29500 25706
rect 39960 25158 39988 26182
rect 41420 26172 41472 26178
rect 41420 26114 41472 26120
rect 40132 25628 40184 25634
rect 40132 25570 40184 25576
rect 39948 25152 40000 25158
rect 39948 25094 40000 25100
rect 27528 24880 27580 24886
rect 27528 24822 27580 24828
rect 27436 21412 27488 21418
rect 27436 21354 27488 21360
rect 25412 17196 25464 17202
rect 25412 17138 25464 17144
rect 900 17050 2532 17052
rect 900 16934 922 17050
rect 2510 16934 2532 17050
rect 900 16932 2532 16934
rect 3348 15170 4980 15172
rect 3348 15054 3370 15170
rect 4958 15054 4980 15170
rect 3348 15052 4980 15054
rect 900 13290 2532 13292
rect 900 13174 922 13290
rect 2510 13174 2532 13290
rect 900 13172 2532 13174
rect 3348 11410 4980 11412
rect 3348 11294 3370 11410
rect 4958 11294 4980 11410
rect 3348 11292 4980 11294
rect 900 9530 2532 9532
rect 900 9414 922 9530
rect 2510 9414 2532 9530
rect 900 9412 2532 9414
rect 3348 7650 4980 7652
rect 3348 7534 3370 7650
rect 4958 7534 4980 7650
rect 3348 7532 4980 7534
rect 900 5770 2532 5772
rect 900 5654 922 5770
rect 2510 5654 2532 5770
rect 900 5652 2532 5654
rect 27540 4554 27568 24822
rect 29948 24730 30108 24752
rect 29948 24674 30000 24730
rect 30056 24674 30108 24730
rect 29948 24652 30108 24674
rect 37372 24676 37424 24682
rect 37372 24618 37424 24624
rect 37384 23458 37412 24618
rect 38292 24200 38344 24206
rect 38292 24142 38344 24148
rect 30932 23452 30984 23458
rect 30932 23394 30984 23400
rect 37372 23452 37424 23458
rect 37372 23394 37424 23400
rect 30944 22370 30972 23394
rect 34980 22500 35032 22506
rect 34980 22442 35032 22448
rect 30932 22364 30984 22370
rect 30932 22306 30984 22312
rect 29092 21888 29144 21894
rect 29092 21830 29144 21836
rect 29104 21400 29132 21830
rect 34992 21418 35020 22442
rect 38304 22370 38332 24142
rect 40144 22506 40172 25570
rect 40132 22500 40184 22506
rect 40132 22442 40184 22448
rect 38292 22364 38344 22370
rect 38292 22306 38344 22312
rect 35072 21888 35124 21894
rect 35072 21830 35124 21836
rect 29736 21412 29788 21418
rect 29104 21372 29736 21400
rect 29736 21354 29788 21360
rect 34980 21412 35032 21418
rect 35084 21400 35112 21830
rect 41432 21418 41460 26114
rect 42708 25696 42760 25702
rect 42708 25638 42760 25644
rect 42720 22506 42748 25638
rect 46032 25158 46060 26182
rect 48424 25158 48452 28902
rect 48516 26246 48544 33748
rect 48688 33730 48740 33736
rect 55904 32090 57536 32092
rect 55904 31974 55926 32090
rect 57514 31974 57536 32090
rect 55904 31972 57536 31974
rect 53456 30210 55088 30212
rect 53456 30094 53478 30210
rect 55066 30094 55088 30210
rect 53456 30092 55088 30094
rect 55904 28330 57536 28332
rect 55904 28214 55926 28330
rect 57514 28214 57536 28330
rect 55904 28212 57536 28214
rect 53456 26450 55088 26452
rect 53456 26334 53478 26450
rect 55066 26334 55088 26450
rect 53456 26332 55088 26334
rect 48504 26240 48556 26246
rect 48504 26182 48556 26188
rect 46020 25152 46072 25158
rect 46020 25094 46072 25100
rect 48412 25152 48464 25158
rect 48412 25094 48464 25100
rect 42892 24676 42944 24682
rect 42892 24618 42944 24624
rect 42904 24206 42932 24618
rect 42892 24200 42944 24206
rect 42892 24142 42944 24148
rect 48516 22506 48544 26182
rect 48596 25628 48648 25634
rect 48596 25570 48648 25576
rect 42708 22500 42760 22506
rect 42708 22442 42760 22448
rect 48504 22500 48556 22506
rect 48504 22442 48556 22448
rect 48608 21418 48636 25570
rect 55904 24570 57536 24572
rect 55904 24454 55926 24570
rect 57514 24454 57536 24570
rect 55904 24452 57536 24454
rect 53456 22690 55088 22692
rect 53456 22574 53478 22690
rect 55066 22574 55088 22690
rect 53456 22572 55088 22574
rect 35716 21412 35768 21418
rect 35084 21372 35716 21400
rect 34980 21354 35032 21360
rect 35716 21354 35768 21360
rect 41420 21412 41472 21418
rect 41420 21354 41472 21360
rect 48596 21412 48648 21418
rect 48596 21354 48648 21360
rect 55904 20810 57536 20812
rect 55904 20694 55926 20810
rect 57514 20694 57536 20810
rect 55904 20692 57536 20694
rect 53456 18930 55088 18932
rect 53456 18814 53478 18930
rect 55066 18814 55088 18930
rect 53456 18812 55088 18814
rect 43996 17400 44048 17406
rect 43996 17342 44048 17348
rect 34336 17264 34388 17270
rect 34336 17206 34388 17212
rect 25504 4548 25556 4554
rect 25504 4490 25556 4496
rect 27528 4548 27580 4554
rect 27528 4490 27580 4496
rect 25516 0 25544 4490
rect 34348 0 34376 17206
rect 44008 11082 44036 17342
rect 55904 17050 57536 17052
rect 55904 16934 55926 17050
rect 57514 16934 57536 17050
rect 55904 16932 57536 16934
rect 53456 15170 55088 15172
rect 53456 15054 53478 15170
rect 55066 15054 55088 15170
rect 53456 15052 55088 15054
rect 49056 15020 49108 15026
rect 49056 14962 49108 14968
rect 44364 14884 44416 14890
rect 44284 14844 44364 14872
rect 44284 13870 44312 14844
rect 44364 14826 44416 14832
rect 46664 14340 46716 14346
rect 46664 14282 46716 14288
rect 44272 13864 44324 13870
rect 44272 13806 44324 13812
rect 44732 11212 44784 11218
rect 44732 11154 44784 11160
rect 43996 11076 44048 11082
rect 43996 11018 44048 11024
rect 44744 6390 44772 11154
rect 46676 10130 46704 14282
rect 46940 13388 46992 13394
rect 46940 13330 46992 13336
rect 46952 11218 46980 13330
rect 46940 11212 46992 11218
rect 46940 11154 46992 11160
rect 49068 10130 49096 14962
rect 49516 13388 49568 13394
rect 49516 13330 49568 13336
rect 46664 10124 46716 10130
rect 46664 10066 46716 10072
rect 49056 10124 49108 10130
rect 49056 10066 49108 10072
rect 45652 9648 45704 9654
rect 45652 9590 45704 9596
rect 45664 9382 45692 9590
rect 45652 9376 45704 9382
rect 45652 9318 45704 9324
rect 49528 7528 49556 13330
rect 55904 13290 57536 13292
rect 55904 13174 55926 13290
rect 57514 13174 57536 13290
rect 55904 13172 57536 13174
rect 53456 11410 55088 11412
rect 53456 11294 53478 11410
rect 55066 11294 55088 11410
rect 53456 11292 55088 11294
rect 55904 9530 57536 9532
rect 55904 9414 55926 9530
rect 57514 9414 57536 9530
rect 55904 9412 57536 9414
rect 49884 9376 49936 9382
rect 49884 9318 49936 9324
rect 49160 7500 49556 7528
rect 49160 7342 49188 7500
rect 49792 7472 49844 7478
rect 49792 7414 49844 7420
rect 49148 7336 49200 7342
rect 49148 7278 49200 7284
rect 49804 6390 49832 7414
rect 49896 7342 49924 9318
rect 53456 7650 55088 7652
rect 53456 7534 53478 7650
rect 55066 7534 55088 7650
rect 53456 7532 55088 7534
rect 49884 7336 49936 7342
rect 49884 7278 49936 7284
rect 44732 6384 44784 6390
rect 44732 6326 44784 6332
rect 49792 6384 49844 6390
rect 49792 6326 49844 6332
rect 55904 5770 57536 5772
rect 55904 5654 55926 5770
rect 57514 5654 57536 5770
rect 55904 5652 57536 5654
<< via2 >>
rect 928 50804 984 50860
rect 1008 50804 1064 50860
rect 1088 50804 1144 50860
rect 1168 50804 1224 50860
rect 1248 50804 1304 50860
rect 1328 50804 1384 50860
rect 1408 50804 1464 50860
rect 1488 50804 1544 50860
rect 1568 50804 1624 50860
rect 1648 50804 1704 50860
rect 1728 50804 1784 50860
rect 1808 50804 1864 50860
rect 1888 50804 1944 50860
rect 1968 50804 2024 50860
rect 2048 50804 2104 50860
rect 2128 50804 2184 50860
rect 2208 50804 2264 50860
rect 2288 50804 2344 50860
rect 2368 50804 2424 50860
rect 2448 50804 2504 50860
rect 55932 50804 55988 50860
rect 56012 50804 56068 50860
rect 56092 50804 56148 50860
rect 56172 50804 56228 50860
rect 56252 50804 56308 50860
rect 56332 50804 56388 50860
rect 56412 50804 56468 50860
rect 56492 50804 56548 50860
rect 56572 50804 56628 50860
rect 56652 50804 56708 50860
rect 56732 50804 56788 50860
rect 56812 50804 56868 50860
rect 56892 50804 56948 50860
rect 56972 50804 57028 50860
rect 57052 50804 57108 50860
rect 57132 50804 57188 50860
rect 57212 50804 57268 50860
rect 57292 50804 57348 50860
rect 57372 50804 57428 50860
rect 57452 50804 57508 50860
rect 3376 48924 3432 48980
rect 3456 48924 3512 48980
rect 3536 48924 3592 48980
rect 3616 48924 3672 48980
rect 3696 48924 3752 48980
rect 3776 48924 3832 48980
rect 3856 48924 3912 48980
rect 3936 48924 3992 48980
rect 4016 48924 4072 48980
rect 4096 48924 4152 48980
rect 4176 48924 4232 48980
rect 4256 48924 4312 48980
rect 4336 48924 4392 48980
rect 4416 48924 4472 48980
rect 4496 48924 4552 48980
rect 4576 48924 4632 48980
rect 4656 48924 4712 48980
rect 4736 48924 4792 48980
rect 4816 48924 4872 48980
rect 4896 48924 4952 48980
rect 53484 48924 53540 48980
rect 53564 48924 53620 48980
rect 53644 48924 53700 48980
rect 53724 48924 53780 48980
rect 53804 48924 53860 48980
rect 53884 48924 53940 48980
rect 53964 48924 54020 48980
rect 54044 48924 54100 48980
rect 54124 48924 54180 48980
rect 54204 48924 54260 48980
rect 54284 48924 54340 48980
rect 54364 48924 54420 48980
rect 54444 48924 54500 48980
rect 54524 48924 54580 48980
rect 54604 48924 54660 48980
rect 54684 48924 54740 48980
rect 54764 48924 54820 48980
rect 54844 48924 54900 48980
rect 54924 48924 54980 48980
rect 55004 48924 55060 48980
rect 5948 48654 6004 48710
rect 6028 48654 6084 48710
rect 13396 48654 13452 48710
rect 13476 48654 13532 48710
rect 5990 47234 6046 47290
rect 13438 47234 13494 47290
rect 928 47044 984 47100
rect 1008 47044 1064 47100
rect 1088 47044 1144 47100
rect 1168 47044 1224 47100
rect 1248 47044 1304 47100
rect 1328 47044 1384 47100
rect 1408 47044 1464 47100
rect 1488 47044 1544 47100
rect 1568 47044 1624 47100
rect 1648 47044 1704 47100
rect 1728 47044 1784 47100
rect 1808 47044 1864 47100
rect 1888 47044 1944 47100
rect 1968 47044 2024 47100
rect 2048 47044 2104 47100
rect 2128 47044 2184 47100
rect 2208 47044 2264 47100
rect 2288 47044 2344 47100
rect 2368 47044 2424 47100
rect 2448 47044 2504 47100
rect 17682 47116 17738 47132
rect 17682 47076 17684 47116
rect 17684 47076 17736 47116
rect 17736 47076 17738 47116
rect 3376 45164 3432 45220
rect 3456 45164 3512 45220
rect 3536 45164 3592 45220
rect 3616 45164 3672 45220
rect 3696 45164 3752 45220
rect 3776 45164 3832 45220
rect 3856 45164 3912 45220
rect 3936 45164 3992 45220
rect 4016 45164 4072 45220
rect 4096 45164 4152 45220
rect 4176 45164 4232 45220
rect 4256 45164 4312 45220
rect 4336 45164 4392 45220
rect 4416 45164 4472 45220
rect 4496 45164 4552 45220
rect 4576 45164 4632 45220
rect 4656 45164 4712 45220
rect 4736 45164 4792 45220
rect 4816 45164 4872 45220
rect 4896 45164 4952 45220
rect 5948 44894 6004 44950
rect 6028 44894 6084 44950
rect 15014 43782 15070 43838
rect 5990 43474 6046 43530
rect 928 43284 984 43340
rect 1008 43284 1064 43340
rect 1088 43284 1144 43340
rect 1168 43284 1224 43340
rect 1248 43284 1304 43340
rect 1328 43284 1384 43340
rect 1408 43284 1464 43340
rect 1488 43284 1544 43340
rect 1568 43284 1624 43340
rect 1648 43284 1704 43340
rect 1728 43284 1784 43340
rect 1808 43284 1864 43340
rect 1888 43284 1944 43340
rect 1968 43284 2024 43340
rect 2048 43284 2104 43340
rect 2128 43284 2184 43340
rect 2208 43284 2264 43340
rect 2288 43284 2344 43340
rect 2368 43284 2424 43340
rect 2448 43284 2504 43340
rect 8298 43308 8354 43350
rect 8298 43294 8300 43308
rect 8300 43294 8352 43308
rect 8352 43294 8354 43308
rect 3376 41404 3432 41460
rect 3456 41404 3512 41460
rect 3536 41404 3592 41460
rect 3616 41404 3672 41460
rect 3696 41404 3752 41460
rect 3776 41404 3832 41460
rect 3856 41404 3912 41460
rect 3936 41404 3992 41460
rect 4016 41404 4072 41460
rect 4096 41404 4152 41460
rect 4176 41404 4232 41460
rect 4256 41404 4312 41460
rect 4336 41404 4392 41460
rect 4416 41404 4472 41460
rect 4496 41404 4552 41460
rect 4576 41404 4632 41460
rect 4656 41404 4712 41460
rect 4736 41404 4792 41460
rect 4816 41404 4872 41460
rect 4896 41404 4952 41460
rect 6340 41134 6396 41190
rect 6420 41134 6476 41190
rect 6382 39714 6438 39770
rect 928 39524 984 39580
rect 1008 39524 1064 39580
rect 1088 39524 1144 39580
rect 1168 39524 1224 39580
rect 1248 39524 1304 39580
rect 1328 39524 1384 39580
rect 1408 39524 1464 39580
rect 1488 39524 1544 39580
rect 1568 39524 1624 39580
rect 1648 39524 1704 39580
rect 1728 39524 1784 39580
rect 1808 39524 1864 39580
rect 1888 39524 1944 39580
rect 1968 39524 2024 39580
rect 2048 39524 2104 39580
rect 2128 39524 2184 39580
rect 2208 39524 2264 39580
rect 2288 39524 2344 39580
rect 2368 39524 2424 39580
rect 2448 39524 2504 39580
rect 14554 43460 14556 43472
rect 14556 43460 14608 43472
rect 14608 43460 14610 43472
rect 14554 43416 14610 43460
rect 15160 41134 15216 41190
rect 15240 41134 15296 41190
rect 15202 39714 15258 39770
rect 15474 39634 15530 39690
rect 3376 37644 3432 37700
rect 3456 37644 3512 37700
rect 3536 37644 3592 37700
rect 3616 37644 3672 37700
rect 3696 37644 3752 37700
rect 3776 37644 3832 37700
rect 3856 37644 3912 37700
rect 3936 37644 3992 37700
rect 4016 37644 4072 37700
rect 4096 37644 4152 37700
rect 4176 37644 4232 37700
rect 4256 37644 4312 37700
rect 4336 37644 4392 37700
rect 4416 37644 4472 37700
rect 4496 37644 4552 37700
rect 4576 37644 4632 37700
rect 4656 37644 4712 37700
rect 4736 37644 4792 37700
rect 4816 37644 4872 37700
rect 4896 37644 4952 37700
rect 12898 37194 12954 37250
rect 928 35764 984 35820
rect 1008 35764 1064 35820
rect 1088 35764 1144 35820
rect 1168 35764 1224 35820
rect 1248 35764 1304 35820
rect 1328 35764 1384 35820
rect 1408 35764 1464 35820
rect 1488 35764 1544 35820
rect 1568 35764 1624 35820
rect 1648 35764 1704 35820
rect 1728 35764 1784 35820
rect 1808 35764 1864 35820
rect 1888 35764 1944 35820
rect 1968 35764 2024 35820
rect 2048 35764 2104 35820
rect 2128 35764 2184 35820
rect 2208 35764 2264 35820
rect 2288 35764 2344 35820
rect 2368 35764 2424 35820
rect 2448 35764 2504 35820
rect 3376 33884 3432 33940
rect 3456 33884 3512 33940
rect 3536 33884 3592 33940
rect 3616 33884 3672 33940
rect 3696 33884 3752 33940
rect 3776 33884 3832 33940
rect 3856 33884 3912 33940
rect 3936 33884 3992 33940
rect 4016 33884 4072 33940
rect 4096 33884 4152 33940
rect 4176 33884 4232 33940
rect 4256 33884 4312 33940
rect 4336 33884 4392 33940
rect 4416 33884 4472 33940
rect 4496 33884 4552 33940
rect 4576 33884 4632 33940
rect 4656 33884 4712 33940
rect 4736 33884 4792 33940
rect 4816 33884 4872 33940
rect 4896 33884 4952 33940
rect 928 32004 984 32060
rect 1008 32004 1064 32060
rect 1088 32004 1144 32060
rect 1168 32004 1224 32060
rect 1248 32004 1304 32060
rect 1328 32004 1384 32060
rect 1408 32004 1464 32060
rect 1488 32004 1544 32060
rect 1568 32004 1624 32060
rect 1648 32004 1704 32060
rect 1728 32004 1784 32060
rect 1808 32004 1864 32060
rect 1888 32004 1944 32060
rect 1968 32004 2024 32060
rect 2048 32004 2104 32060
rect 2128 32004 2184 32060
rect 2208 32004 2264 32060
rect 2288 32004 2344 32060
rect 2368 32004 2424 32060
rect 2448 32004 2504 32060
rect 3376 30124 3432 30180
rect 3456 30124 3512 30180
rect 3536 30124 3592 30180
rect 3616 30124 3672 30180
rect 3696 30124 3752 30180
rect 3776 30124 3832 30180
rect 3856 30124 3912 30180
rect 3936 30124 3992 30180
rect 4016 30124 4072 30180
rect 4096 30124 4152 30180
rect 4176 30124 4232 30180
rect 4256 30124 4312 30180
rect 4336 30124 4392 30180
rect 4416 30124 4472 30180
rect 4496 30124 4552 30180
rect 4576 30124 4632 30180
rect 4656 30124 4712 30180
rect 4736 30124 4792 30180
rect 4816 30124 4872 30180
rect 4896 30124 4952 30180
rect 928 28244 984 28300
rect 1008 28244 1064 28300
rect 1088 28244 1144 28300
rect 1168 28244 1224 28300
rect 1248 28244 1304 28300
rect 1328 28244 1384 28300
rect 1408 28244 1464 28300
rect 1488 28244 1544 28300
rect 1568 28244 1624 28300
rect 1648 28244 1704 28300
rect 1728 28244 1784 28300
rect 1808 28244 1864 28300
rect 1888 28244 1944 28300
rect 1968 28244 2024 28300
rect 2048 28244 2104 28300
rect 2128 28244 2184 28300
rect 2208 28244 2264 28300
rect 2288 28244 2344 28300
rect 2368 28244 2424 28300
rect 2448 28244 2504 28300
rect 3376 26364 3432 26420
rect 3456 26364 3512 26420
rect 3536 26364 3592 26420
rect 3616 26364 3672 26420
rect 3696 26364 3752 26420
rect 3776 26364 3832 26420
rect 3856 26364 3912 26420
rect 3936 26364 3992 26420
rect 4016 26364 4072 26420
rect 4096 26364 4152 26420
rect 4176 26364 4232 26420
rect 4256 26364 4312 26420
rect 4336 26364 4392 26420
rect 4416 26364 4472 26420
rect 4496 26364 4552 26420
rect 4576 26364 4632 26420
rect 4656 26364 4712 26420
rect 4736 26364 4792 26420
rect 4816 26364 4872 26420
rect 4896 26364 4952 26420
rect 928 24484 984 24540
rect 1008 24484 1064 24540
rect 1088 24484 1144 24540
rect 1168 24484 1224 24540
rect 1248 24484 1304 24540
rect 1328 24484 1384 24540
rect 1408 24484 1464 24540
rect 1488 24484 1544 24540
rect 1568 24484 1624 24540
rect 1648 24484 1704 24540
rect 1728 24484 1784 24540
rect 1808 24484 1864 24540
rect 1888 24484 1944 24540
rect 1968 24484 2024 24540
rect 2048 24484 2104 24540
rect 2128 24484 2184 24540
rect 2208 24484 2264 24540
rect 2288 24484 2344 24540
rect 2368 24484 2424 24540
rect 2448 24484 2504 24540
rect 3376 22604 3432 22660
rect 3456 22604 3512 22660
rect 3536 22604 3592 22660
rect 3616 22604 3672 22660
rect 3696 22604 3752 22660
rect 3776 22604 3832 22660
rect 3856 22604 3912 22660
rect 3936 22604 3992 22660
rect 4016 22604 4072 22660
rect 4096 22604 4152 22660
rect 4176 22604 4232 22660
rect 4256 22604 4312 22660
rect 4336 22604 4392 22660
rect 4416 22604 4472 22660
rect 4496 22604 4552 22660
rect 4576 22604 4632 22660
rect 4656 22604 4712 22660
rect 4736 22604 4792 22660
rect 4816 22604 4872 22660
rect 4896 22604 4952 22660
rect 23754 43416 23810 43472
rect 22190 41342 22246 41398
rect 33414 37612 33416 37616
rect 33416 37612 33468 37616
rect 33468 37612 33470 37616
rect 33414 37560 33470 37612
rect 29958 37374 30014 37430
rect 30038 37374 30094 37430
rect 29458 36984 29514 37006
rect 29458 36950 29460 36984
rect 29460 36950 29512 36984
rect 29512 36950 29514 36984
rect 30000 35954 30056 36010
rect 37554 35980 37556 36030
rect 37556 35980 37608 36030
rect 37608 35980 37610 36030
rect 37554 35974 37610 35980
rect 33414 33778 33470 33834
rect 26234 33614 26290 33670
rect 26314 33614 26370 33670
rect 33682 33614 33738 33670
rect 33762 33614 33818 33670
rect 26276 32194 26332 32250
rect 33724 32194 33780 32250
rect 33414 30132 33416 30174
rect 33416 30132 33468 30174
rect 33468 30132 33470 30174
rect 33414 30118 33470 30132
rect 29958 29854 30014 29910
rect 30038 29854 30094 29910
rect 928 20724 984 20780
rect 1008 20724 1064 20780
rect 1088 20724 1144 20780
rect 1168 20724 1224 20780
rect 1248 20724 1304 20780
rect 1328 20724 1384 20780
rect 1408 20724 1464 20780
rect 1488 20724 1544 20780
rect 1568 20724 1624 20780
rect 1648 20724 1704 20780
rect 1728 20724 1784 20780
rect 1808 20724 1864 20780
rect 1888 20724 1944 20780
rect 1968 20724 2024 20780
rect 2048 20724 2104 20780
rect 2128 20724 2184 20780
rect 2208 20724 2264 20780
rect 2288 20724 2344 20780
rect 2368 20724 2424 20780
rect 2448 20724 2504 20780
rect 3376 18844 3432 18900
rect 3456 18844 3512 18900
rect 3536 18844 3592 18900
rect 3616 18844 3672 18900
rect 3696 18844 3752 18900
rect 3776 18844 3832 18900
rect 3856 18844 3912 18900
rect 3936 18844 3992 18900
rect 4016 18844 4072 18900
rect 4096 18844 4152 18900
rect 4176 18844 4232 18900
rect 4256 18844 4312 18900
rect 4336 18844 4392 18900
rect 4416 18844 4472 18900
rect 4496 18844 4552 18900
rect 4576 18844 4632 18900
rect 4656 18844 4712 18900
rect 4736 18844 4792 18900
rect 4816 18844 4872 18900
rect 4896 18844 4952 18900
rect 30000 28434 30056 28490
rect 55932 47044 55988 47100
rect 56012 47044 56068 47100
rect 56092 47044 56148 47100
rect 56172 47044 56228 47100
rect 56252 47044 56308 47100
rect 56332 47044 56388 47100
rect 56412 47044 56468 47100
rect 56492 47044 56548 47100
rect 56572 47044 56628 47100
rect 56652 47044 56708 47100
rect 56732 47044 56788 47100
rect 56812 47044 56868 47100
rect 56892 47044 56948 47100
rect 56972 47044 57028 47100
rect 57052 47044 57108 47100
rect 57132 47044 57188 47100
rect 57212 47044 57268 47100
rect 57292 47044 57348 47100
rect 57372 47044 57428 47100
rect 57452 47044 57508 47100
rect 53484 45164 53540 45220
rect 53564 45164 53620 45220
rect 53644 45164 53700 45220
rect 53724 45164 53780 45220
rect 53804 45164 53860 45220
rect 53884 45164 53940 45220
rect 53964 45164 54020 45220
rect 54044 45164 54100 45220
rect 54124 45164 54180 45220
rect 54204 45164 54260 45220
rect 54284 45164 54340 45220
rect 54364 45164 54420 45220
rect 54444 45164 54500 45220
rect 54524 45164 54580 45220
rect 54604 45164 54660 45220
rect 54684 45164 54740 45220
rect 54764 45164 54820 45220
rect 54844 45164 54900 45220
rect 54924 45164 54980 45220
rect 55004 45164 55060 45220
rect 55932 43284 55988 43340
rect 56012 43284 56068 43340
rect 56092 43284 56148 43340
rect 56172 43284 56228 43340
rect 56252 43284 56308 43340
rect 56332 43284 56388 43340
rect 56412 43284 56468 43340
rect 56492 43284 56548 43340
rect 56572 43284 56628 43340
rect 56652 43284 56708 43340
rect 56732 43284 56788 43340
rect 56812 43284 56868 43340
rect 56892 43284 56948 43340
rect 56972 43284 57028 43340
rect 57052 43284 57108 43340
rect 57132 43284 57188 43340
rect 57212 43284 57268 43340
rect 57292 43284 57348 43340
rect 57372 43284 57428 43340
rect 57452 43284 57508 43340
rect 53484 41404 53540 41460
rect 53564 41404 53620 41460
rect 53644 41404 53700 41460
rect 53724 41404 53780 41460
rect 53804 41404 53860 41460
rect 53884 41404 53940 41460
rect 53964 41404 54020 41460
rect 54044 41404 54100 41460
rect 54124 41404 54180 41460
rect 54204 41404 54260 41460
rect 54284 41404 54340 41460
rect 54364 41404 54420 41460
rect 54444 41404 54500 41460
rect 54524 41404 54580 41460
rect 54604 41404 54660 41460
rect 54684 41404 54740 41460
rect 54764 41404 54820 41460
rect 54844 41404 54900 41460
rect 54924 41404 54980 41460
rect 55004 41404 55060 41460
rect 55932 39524 55988 39580
rect 56012 39524 56068 39580
rect 56092 39524 56148 39580
rect 56172 39524 56228 39580
rect 56252 39524 56308 39580
rect 56332 39524 56388 39580
rect 56412 39524 56468 39580
rect 56492 39524 56548 39580
rect 56572 39524 56628 39580
rect 56652 39524 56708 39580
rect 56732 39524 56788 39580
rect 56812 39524 56868 39580
rect 56892 39524 56948 39580
rect 56972 39524 57028 39580
rect 57052 39524 57108 39580
rect 57132 39524 57188 39580
rect 57212 39524 57268 39580
rect 57292 39524 57348 39580
rect 57372 39524 57428 39580
rect 57452 39524 57508 39580
rect 53484 37644 53540 37700
rect 53564 37644 53620 37700
rect 53644 37644 53700 37700
rect 53724 37644 53780 37700
rect 53804 37644 53860 37700
rect 53884 37644 53940 37700
rect 53964 37644 54020 37700
rect 54044 37644 54100 37700
rect 54124 37644 54180 37700
rect 54204 37644 54260 37700
rect 54284 37644 54340 37700
rect 54364 37644 54420 37700
rect 54444 37644 54500 37700
rect 54524 37644 54580 37700
rect 54604 37644 54660 37700
rect 54684 37644 54740 37700
rect 54764 37644 54820 37700
rect 54844 37644 54900 37700
rect 54924 37644 54980 37700
rect 55004 37644 55060 37700
rect 55932 35764 55988 35820
rect 56012 35764 56068 35820
rect 56092 35764 56148 35820
rect 56172 35764 56228 35820
rect 56252 35764 56308 35820
rect 56332 35764 56388 35820
rect 56412 35764 56468 35820
rect 56492 35764 56548 35820
rect 56572 35764 56628 35820
rect 56652 35764 56708 35820
rect 56732 35764 56788 35820
rect 56812 35764 56868 35820
rect 56892 35764 56948 35820
rect 56972 35764 57028 35820
rect 57052 35764 57108 35820
rect 57132 35764 57188 35820
rect 57212 35764 57268 35820
rect 57292 35764 57348 35820
rect 57372 35764 57428 35820
rect 57452 35764 57508 35820
rect 53484 33884 53540 33940
rect 53564 33884 53620 33940
rect 53644 33884 53700 33940
rect 53724 33884 53780 33940
rect 53804 33884 53860 33940
rect 53884 33884 53940 33940
rect 53964 33884 54020 33940
rect 54044 33884 54100 33940
rect 54124 33884 54180 33940
rect 54204 33884 54260 33940
rect 54284 33884 54340 33940
rect 54364 33884 54420 33940
rect 54444 33884 54500 33940
rect 54524 33884 54580 33940
rect 54604 33884 54660 33940
rect 54684 33884 54740 33940
rect 54764 33884 54820 33940
rect 54844 33884 54900 33940
rect 54924 33884 54980 33940
rect 55004 33884 55060 33940
rect 33414 26336 33470 26392
rect 29958 26094 30014 26150
rect 30038 26094 30094 26150
rect 29458 25764 29514 25782
rect 29458 25726 29460 25764
rect 29460 25726 29512 25764
rect 29512 25726 29514 25764
rect 928 16964 984 17020
rect 1008 16964 1064 17020
rect 1088 16964 1144 17020
rect 1168 16964 1224 17020
rect 1248 16964 1304 17020
rect 1328 16964 1384 17020
rect 1408 16964 1464 17020
rect 1488 16964 1544 17020
rect 1568 16964 1624 17020
rect 1648 16964 1704 17020
rect 1728 16964 1784 17020
rect 1808 16964 1864 17020
rect 1888 16964 1944 17020
rect 1968 16964 2024 17020
rect 2048 16964 2104 17020
rect 2128 16964 2184 17020
rect 2208 16964 2264 17020
rect 2288 16964 2344 17020
rect 2368 16964 2424 17020
rect 2448 16964 2504 17020
rect 3376 15084 3432 15140
rect 3456 15084 3512 15140
rect 3536 15084 3592 15140
rect 3616 15084 3672 15140
rect 3696 15084 3752 15140
rect 3776 15084 3832 15140
rect 3856 15084 3912 15140
rect 3936 15084 3992 15140
rect 4016 15084 4072 15140
rect 4096 15084 4152 15140
rect 4176 15084 4232 15140
rect 4256 15084 4312 15140
rect 4336 15084 4392 15140
rect 4416 15084 4472 15140
rect 4496 15084 4552 15140
rect 4576 15084 4632 15140
rect 4656 15084 4712 15140
rect 4736 15084 4792 15140
rect 4816 15084 4872 15140
rect 4896 15084 4952 15140
rect 928 13204 984 13260
rect 1008 13204 1064 13260
rect 1088 13204 1144 13260
rect 1168 13204 1224 13260
rect 1248 13204 1304 13260
rect 1328 13204 1384 13260
rect 1408 13204 1464 13260
rect 1488 13204 1544 13260
rect 1568 13204 1624 13260
rect 1648 13204 1704 13260
rect 1728 13204 1784 13260
rect 1808 13204 1864 13260
rect 1888 13204 1944 13260
rect 1968 13204 2024 13260
rect 2048 13204 2104 13260
rect 2128 13204 2184 13260
rect 2208 13204 2264 13260
rect 2288 13204 2344 13260
rect 2368 13204 2424 13260
rect 2448 13204 2504 13260
rect 3376 11324 3432 11380
rect 3456 11324 3512 11380
rect 3536 11324 3592 11380
rect 3616 11324 3672 11380
rect 3696 11324 3752 11380
rect 3776 11324 3832 11380
rect 3856 11324 3912 11380
rect 3936 11324 3992 11380
rect 4016 11324 4072 11380
rect 4096 11324 4152 11380
rect 4176 11324 4232 11380
rect 4256 11324 4312 11380
rect 4336 11324 4392 11380
rect 4416 11324 4472 11380
rect 4496 11324 4552 11380
rect 4576 11324 4632 11380
rect 4656 11324 4712 11380
rect 4736 11324 4792 11380
rect 4816 11324 4872 11380
rect 4896 11324 4952 11380
rect 928 9444 984 9500
rect 1008 9444 1064 9500
rect 1088 9444 1144 9500
rect 1168 9444 1224 9500
rect 1248 9444 1304 9500
rect 1328 9444 1384 9500
rect 1408 9444 1464 9500
rect 1488 9444 1544 9500
rect 1568 9444 1624 9500
rect 1648 9444 1704 9500
rect 1728 9444 1784 9500
rect 1808 9444 1864 9500
rect 1888 9444 1944 9500
rect 1968 9444 2024 9500
rect 2048 9444 2104 9500
rect 2128 9444 2184 9500
rect 2208 9444 2264 9500
rect 2288 9444 2344 9500
rect 2368 9444 2424 9500
rect 2448 9444 2504 9500
rect 3376 7564 3432 7620
rect 3456 7564 3512 7620
rect 3536 7564 3592 7620
rect 3616 7564 3672 7620
rect 3696 7564 3752 7620
rect 3776 7564 3832 7620
rect 3856 7564 3912 7620
rect 3936 7564 3992 7620
rect 4016 7564 4072 7620
rect 4096 7564 4152 7620
rect 4176 7564 4232 7620
rect 4256 7564 4312 7620
rect 4336 7564 4392 7620
rect 4416 7564 4472 7620
rect 4496 7564 4552 7620
rect 4576 7564 4632 7620
rect 4656 7564 4712 7620
rect 4736 7564 4792 7620
rect 4816 7564 4872 7620
rect 4896 7564 4952 7620
rect 928 5684 984 5740
rect 1008 5684 1064 5740
rect 1088 5684 1144 5740
rect 1168 5684 1224 5740
rect 1248 5684 1304 5740
rect 1328 5684 1384 5740
rect 1408 5684 1464 5740
rect 1488 5684 1544 5740
rect 1568 5684 1624 5740
rect 1648 5684 1704 5740
rect 1728 5684 1784 5740
rect 1808 5684 1864 5740
rect 1888 5684 1944 5740
rect 1968 5684 2024 5740
rect 2048 5684 2104 5740
rect 2128 5684 2184 5740
rect 2208 5684 2264 5740
rect 2288 5684 2344 5740
rect 2368 5684 2424 5740
rect 2448 5684 2504 5740
rect 30000 24674 30056 24730
rect 55932 32004 55988 32060
rect 56012 32004 56068 32060
rect 56092 32004 56148 32060
rect 56172 32004 56228 32060
rect 56252 32004 56308 32060
rect 56332 32004 56388 32060
rect 56412 32004 56468 32060
rect 56492 32004 56548 32060
rect 56572 32004 56628 32060
rect 56652 32004 56708 32060
rect 56732 32004 56788 32060
rect 56812 32004 56868 32060
rect 56892 32004 56948 32060
rect 56972 32004 57028 32060
rect 57052 32004 57108 32060
rect 57132 32004 57188 32060
rect 57212 32004 57268 32060
rect 57292 32004 57348 32060
rect 57372 32004 57428 32060
rect 57452 32004 57508 32060
rect 53484 30124 53540 30180
rect 53564 30124 53620 30180
rect 53644 30124 53700 30180
rect 53724 30124 53780 30180
rect 53804 30124 53860 30180
rect 53884 30124 53940 30180
rect 53964 30124 54020 30180
rect 54044 30124 54100 30180
rect 54124 30124 54180 30180
rect 54204 30124 54260 30180
rect 54284 30124 54340 30180
rect 54364 30124 54420 30180
rect 54444 30124 54500 30180
rect 54524 30124 54580 30180
rect 54604 30124 54660 30180
rect 54684 30124 54740 30180
rect 54764 30124 54820 30180
rect 54844 30124 54900 30180
rect 54924 30124 54980 30180
rect 55004 30124 55060 30180
rect 55932 28244 55988 28300
rect 56012 28244 56068 28300
rect 56092 28244 56148 28300
rect 56172 28244 56228 28300
rect 56252 28244 56308 28300
rect 56332 28244 56388 28300
rect 56412 28244 56468 28300
rect 56492 28244 56548 28300
rect 56572 28244 56628 28300
rect 56652 28244 56708 28300
rect 56732 28244 56788 28300
rect 56812 28244 56868 28300
rect 56892 28244 56948 28300
rect 56972 28244 57028 28300
rect 57052 28244 57108 28300
rect 57132 28244 57188 28300
rect 57212 28244 57268 28300
rect 57292 28244 57348 28300
rect 57372 28244 57428 28300
rect 57452 28244 57508 28300
rect 53484 26364 53540 26420
rect 53564 26364 53620 26420
rect 53644 26364 53700 26420
rect 53724 26364 53780 26420
rect 53804 26364 53860 26420
rect 53884 26364 53940 26420
rect 53964 26364 54020 26420
rect 54044 26364 54100 26420
rect 54124 26364 54180 26420
rect 54204 26364 54260 26420
rect 54284 26364 54340 26420
rect 54364 26364 54420 26420
rect 54444 26364 54500 26420
rect 54524 26364 54580 26420
rect 54604 26364 54660 26420
rect 54684 26364 54740 26420
rect 54764 26364 54820 26420
rect 54844 26364 54900 26420
rect 54924 26364 54980 26420
rect 55004 26364 55060 26420
rect 55932 24484 55988 24540
rect 56012 24484 56068 24540
rect 56092 24484 56148 24540
rect 56172 24484 56228 24540
rect 56252 24484 56308 24540
rect 56332 24484 56388 24540
rect 56412 24484 56468 24540
rect 56492 24484 56548 24540
rect 56572 24484 56628 24540
rect 56652 24484 56708 24540
rect 56732 24484 56788 24540
rect 56812 24484 56868 24540
rect 56892 24484 56948 24540
rect 56972 24484 57028 24540
rect 57052 24484 57108 24540
rect 57132 24484 57188 24540
rect 57212 24484 57268 24540
rect 57292 24484 57348 24540
rect 57372 24484 57428 24540
rect 57452 24484 57508 24540
rect 53484 22604 53540 22660
rect 53564 22604 53620 22660
rect 53644 22604 53700 22660
rect 53724 22604 53780 22660
rect 53804 22604 53860 22660
rect 53884 22604 53940 22660
rect 53964 22604 54020 22660
rect 54044 22604 54100 22660
rect 54124 22604 54180 22660
rect 54204 22604 54260 22660
rect 54284 22604 54340 22660
rect 54364 22604 54420 22660
rect 54444 22604 54500 22660
rect 54524 22604 54580 22660
rect 54604 22604 54660 22660
rect 54684 22604 54740 22660
rect 54764 22604 54820 22660
rect 54844 22604 54900 22660
rect 54924 22604 54980 22660
rect 55004 22604 55060 22660
rect 55932 20724 55988 20780
rect 56012 20724 56068 20780
rect 56092 20724 56148 20780
rect 56172 20724 56228 20780
rect 56252 20724 56308 20780
rect 56332 20724 56388 20780
rect 56412 20724 56468 20780
rect 56492 20724 56548 20780
rect 56572 20724 56628 20780
rect 56652 20724 56708 20780
rect 56732 20724 56788 20780
rect 56812 20724 56868 20780
rect 56892 20724 56948 20780
rect 56972 20724 57028 20780
rect 57052 20724 57108 20780
rect 57132 20724 57188 20780
rect 57212 20724 57268 20780
rect 57292 20724 57348 20780
rect 57372 20724 57428 20780
rect 57452 20724 57508 20780
rect 53484 18844 53540 18900
rect 53564 18844 53620 18900
rect 53644 18844 53700 18900
rect 53724 18844 53780 18900
rect 53804 18844 53860 18900
rect 53884 18844 53940 18900
rect 53964 18844 54020 18900
rect 54044 18844 54100 18900
rect 54124 18844 54180 18900
rect 54204 18844 54260 18900
rect 54284 18844 54340 18900
rect 54364 18844 54420 18900
rect 54444 18844 54500 18900
rect 54524 18844 54580 18900
rect 54604 18844 54660 18900
rect 54684 18844 54740 18900
rect 54764 18844 54820 18900
rect 54844 18844 54900 18900
rect 54924 18844 54980 18900
rect 55004 18844 55060 18900
rect 55932 16964 55988 17020
rect 56012 16964 56068 17020
rect 56092 16964 56148 17020
rect 56172 16964 56228 17020
rect 56252 16964 56308 17020
rect 56332 16964 56388 17020
rect 56412 16964 56468 17020
rect 56492 16964 56548 17020
rect 56572 16964 56628 17020
rect 56652 16964 56708 17020
rect 56732 16964 56788 17020
rect 56812 16964 56868 17020
rect 56892 16964 56948 17020
rect 56972 16964 57028 17020
rect 57052 16964 57108 17020
rect 57132 16964 57188 17020
rect 57212 16964 57268 17020
rect 57292 16964 57348 17020
rect 57372 16964 57428 17020
rect 57452 16964 57508 17020
rect 53484 15084 53540 15140
rect 53564 15084 53620 15140
rect 53644 15084 53700 15140
rect 53724 15084 53780 15140
rect 53804 15084 53860 15140
rect 53884 15084 53940 15140
rect 53964 15084 54020 15140
rect 54044 15084 54100 15140
rect 54124 15084 54180 15140
rect 54204 15084 54260 15140
rect 54284 15084 54340 15140
rect 54364 15084 54420 15140
rect 54444 15084 54500 15140
rect 54524 15084 54580 15140
rect 54604 15084 54660 15140
rect 54684 15084 54740 15140
rect 54764 15084 54820 15140
rect 54844 15084 54900 15140
rect 54924 15084 54980 15140
rect 55004 15084 55060 15140
rect 55932 13204 55988 13260
rect 56012 13204 56068 13260
rect 56092 13204 56148 13260
rect 56172 13204 56228 13260
rect 56252 13204 56308 13260
rect 56332 13204 56388 13260
rect 56412 13204 56468 13260
rect 56492 13204 56548 13260
rect 56572 13204 56628 13260
rect 56652 13204 56708 13260
rect 56732 13204 56788 13260
rect 56812 13204 56868 13260
rect 56892 13204 56948 13260
rect 56972 13204 57028 13260
rect 57052 13204 57108 13260
rect 57132 13204 57188 13260
rect 57212 13204 57268 13260
rect 57292 13204 57348 13260
rect 57372 13204 57428 13260
rect 57452 13204 57508 13260
rect 53484 11324 53540 11380
rect 53564 11324 53620 11380
rect 53644 11324 53700 11380
rect 53724 11324 53780 11380
rect 53804 11324 53860 11380
rect 53884 11324 53940 11380
rect 53964 11324 54020 11380
rect 54044 11324 54100 11380
rect 54124 11324 54180 11380
rect 54204 11324 54260 11380
rect 54284 11324 54340 11380
rect 54364 11324 54420 11380
rect 54444 11324 54500 11380
rect 54524 11324 54580 11380
rect 54604 11324 54660 11380
rect 54684 11324 54740 11380
rect 54764 11324 54820 11380
rect 54844 11324 54900 11380
rect 54924 11324 54980 11380
rect 55004 11324 55060 11380
rect 55932 9444 55988 9500
rect 56012 9444 56068 9500
rect 56092 9444 56148 9500
rect 56172 9444 56228 9500
rect 56252 9444 56308 9500
rect 56332 9444 56388 9500
rect 56412 9444 56468 9500
rect 56492 9444 56548 9500
rect 56572 9444 56628 9500
rect 56652 9444 56708 9500
rect 56732 9444 56788 9500
rect 56812 9444 56868 9500
rect 56892 9444 56948 9500
rect 56972 9444 57028 9500
rect 57052 9444 57108 9500
rect 57132 9444 57188 9500
rect 57212 9444 57268 9500
rect 57292 9444 57348 9500
rect 57372 9444 57428 9500
rect 57452 9444 57508 9500
rect 53484 7564 53540 7620
rect 53564 7564 53620 7620
rect 53644 7564 53700 7620
rect 53724 7564 53780 7620
rect 53804 7564 53860 7620
rect 53884 7564 53940 7620
rect 53964 7564 54020 7620
rect 54044 7564 54100 7620
rect 54124 7564 54180 7620
rect 54204 7564 54260 7620
rect 54284 7564 54340 7620
rect 54364 7564 54420 7620
rect 54444 7564 54500 7620
rect 54524 7564 54580 7620
rect 54604 7564 54660 7620
rect 54684 7564 54740 7620
rect 54764 7564 54820 7620
rect 54844 7564 54900 7620
rect 54924 7564 54980 7620
rect 55004 7564 55060 7620
rect 55932 5684 55988 5740
rect 56012 5684 56068 5740
rect 56092 5684 56148 5740
rect 56172 5684 56228 5740
rect 56252 5684 56308 5740
rect 56332 5684 56388 5740
rect 56412 5684 56468 5740
rect 56492 5684 56548 5740
rect 56572 5684 56628 5740
rect 56652 5684 56708 5740
rect 56732 5684 56788 5740
rect 56812 5684 56868 5740
rect 56892 5684 56948 5740
rect 56972 5684 57028 5740
rect 57052 5684 57108 5740
rect 57132 5684 57188 5740
rect 57212 5684 57268 5740
rect 57292 5684 57348 5740
rect 57372 5684 57428 5740
rect 57452 5684 57508 5740
<< metal3 >>
rect 900 50864 2532 50892
rect 900 50800 924 50864
rect 988 50800 1004 50864
rect 1068 50800 1084 50864
rect 1148 50800 1164 50864
rect 1228 50800 1244 50864
rect 1308 50800 1324 50864
rect 1388 50800 1404 50864
rect 1468 50800 1484 50864
rect 1548 50800 1564 50864
rect 1628 50800 1644 50864
rect 1708 50800 1724 50864
rect 1788 50800 1804 50864
rect 1868 50800 1884 50864
rect 1948 50800 1964 50864
rect 2028 50800 2044 50864
rect 2108 50800 2124 50864
rect 2188 50800 2204 50864
rect 2268 50800 2284 50864
rect 2348 50800 2364 50864
rect 2428 50800 2444 50864
rect 2508 50800 2532 50864
rect 900 50772 2532 50800
rect 55904 50864 57536 50892
rect 55904 50800 55928 50864
rect 55992 50800 56008 50864
rect 56072 50800 56088 50864
rect 56152 50800 56168 50864
rect 56232 50800 56248 50864
rect 56312 50800 56328 50864
rect 56392 50800 56408 50864
rect 56472 50800 56488 50864
rect 56552 50800 56568 50864
rect 56632 50800 56648 50864
rect 56712 50800 56728 50864
rect 56792 50800 56808 50864
rect 56872 50800 56888 50864
rect 56952 50800 56968 50864
rect 57032 50800 57048 50864
rect 57112 50800 57128 50864
rect 57192 50800 57208 50864
rect 57272 50800 57288 50864
rect 57352 50800 57368 50864
rect 57432 50800 57448 50864
rect 57512 50800 57536 50864
rect 55904 50772 57536 50800
rect 3348 48984 4980 49012
rect 3348 48920 3372 48984
rect 3436 48920 3452 48984
rect 3516 48920 3532 48984
rect 3596 48920 3612 48984
rect 3676 48920 3692 48984
rect 3756 48920 3772 48984
rect 3836 48920 3852 48984
rect 3916 48920 3932 48984
rect 3996 48920 4012 48984
rect 4076 48920 4092 48984
rect 4156 48920 4172 48984
rect 4236 48920 4252 48984
rect 4316 48920 4332 48984
rect 4396 48920 4412 48984
rect 4476 48920 4492 48984
rect 4556 48920 4572 48984
rect 4636 48920 4652 48984
rect 4716 48920 4732 48984
rect 4796 48920 4812 48984
rect 4876 48920 4892 48984
rect 4956 48920 4980 48984
rect 3348 48892 4980 48920
rect 53456 48984 55088 49012
rect 53456 48920 53480 48984
rect 53544 48920 53560 48984
rect 53624 48920 53640 48984
rect 53704 48920 53720 48984
rect 53784 48920 53800 48984
rect 53864 48920 53880 48984
rect 53944 48920 53960 48984
rect 54024 48920 54040 48984
rect 54104 48920 54120 48984
rect 54184 48920 54200 48984
rect 54264 48920 54280 48984
rect 54344 48920 54360 48984
rect 54424 48920 54440 48984
rect 54504 48920 54520 48984
rect 54584 48920 54600 48984
rect 54664 48920 54680 48984
rect 54744 48920 54760 48984
rect 54824 48920 54840 48984
rect 54904 48920 54920 48984
rect 54984 48920 55000 48984
rect 55064 48920 55088 48984
rect 53456 48892 55088 48920
rect 5916 48710 13088 48722
rect 5916 48654 5948 48710
rect 6004 48654 6028 48710
rect 6084 48694 13088 48710
rect 6084 48654 6532 48694
rect 5916 48630 6532 48654
rect 6596 48630 7251 48694
rect 7315 48630 7970 48694
rect 8034 48630 8689 48694
rect 8753 48630 9408 48694
rect 9472 48630 10127 48694
rect 10191 48630 10846 48694
rect 10910 48630 11565 48694
rect 11629 48630 12284 48694
rect 12348 48630 13003 48694
rect 13067 48630 13088 48694
rect 5916 48614 13088 48630
rect 5916 48550 6532 48614
rect 6596 48550 7251 48614
rect 7315 48550 7970 48614
rect 8034 48550 8689 48614
rect 8753 48550 9408 48614
rect 9472 48550 10127 48614
rect 10191 48550 10846 48614
rect 10910 48550 11565 48614
rect 11629 48550 12284 48614
rect 12348 48550 13003 48614
rect 13067 48550 13088 48614
rect 5916 48534 13088 48550
rect 5916 48470 6532 48534
rect 6596 48470 7251 48534
rect 7315 48470 7970 48534
rect 8034 48470 8689 48534
rect 8753 48470 9408 48534
rect 9472 48470 10127 48534
rect 10191 48470 10846 48534
rect 10910 48470 11565 48534
rect 11629 48470 12284 48534
rect 12348 48470 13003 48534
rect 13067 48470 13088 48534
rect 5916 48454 13088 48470
rect 5916 48390 6532 48454
rect 6596 48390 7251 48454
rect 7315 48390 7970 48454
rect 8034 48390 8689 48454
rect 8753 48390 9408 48454
rect 9472 48390 10127 48454
rect 10191 48390 10846 48454
rect 10910 48390 11565 48454
rect 11629 48390 12284 48454
rect 12348 48390 13003 48454
rect 13067 48390 13088 48454
rect 5916 48374 13088 48390
rect 5916 48310 6532 48374
rect 6596 48310 7251 48374
rect 7315 48310 7970 48374
rect 8034 48310 8689 48374
rect 8753 48310 9408 48374
rect 9472 48310 10127 48374
rect 10191 48310 10846 48374
rect 10910 48310 11565 48374
rect 11629 48310 12284 48374
rect 12348 48310 13003 48374
rect 13067 48310 13088 48374
rect 5916 48294 13088 48310
rect 5916 48230 6532 48294
rect 6596 48230 7251 48294
rect 7315 48230 7970 48294
rect 8034 48230 8689 48294
rect 8753 48230 9408 48294
rect 9472 48230 10127 48294
rect 10191 48230 10846 48294
rect 10910 48230 11565 48294
rect 11629 48230 12284 48294
rect 12348 48230 13003 48294
rect 13067 48230 13088 48294
rect 5916 48214 13088 48230
rect 5916 48150 6532 48214
rect 6596 48150 7251 48214
rect 7315 48150 7970 48214
rect 8034 48150 8689 48214
rect 8753 48150 9408 48214
rect 9472 48150 10127 48214
rect 10191 48150 10846 48214
rect 10910 48150 11565 48214
rect 11629 48150 12284 48214
rect 12348 48150 13003 48214
rect 13067 48150 13088 48214
rect 5916 47994 13088 48150
rect 5916 47930 6532 47994
rect 6596 47930 7251 47994
rect 7315 47930 7970 47994
rect 8034 47930 8689 47994
rect 8753 47930 9408 47994
rect 9472 47930 10127 47994
rect 10191 47930 10846 47994
rect 10910 47930 11565 47994
rect 11629 47930 12284 47994
rect 12348 47930 13003 47994
rect 13067 47930 13088 47994
rect 5916 47914 13088 47930
rect 5916 47850 6532 47914
rect 6596 47850 7251 47914
rect 7315 47850 7970 47914
rect 8034 47850 8689 47914
rect 8753 47850 9408 47914
rect 9472 47850 10127 47914
rect 10191 47850 10846 47914
rect 10910 47850 11565 47914
rect 11629 47850 12284 47914
rect 12348 47850 13003 47914
rect 13067 47850 13088 47914
rect 5916 47834 13088 47850
rect 5916 47770 6532 47834
rect 6596 47770 7251 47834
rect 7315 47770 7970 47834
rect 8034 47770 8689 47834
rect 8753 47770 9408 47834
rect 9472 47770 10127 47834
rect 10191 47770 10846 47834
rect 10910 47770 11565 47834
rect 11629 47770 12284 47834
rect 12348 47770 13003 47834
rect 13067 47770 13088 47834
rect 5916 47754 13088 47770
rect 5916 47690 6532 47754
rect 6596 47690 7251 47754
rect 7315 47690 7970 47754
rect 8034 47690 8689 47754
rect 8753 47690 9408 47754
rect 9472 47690 10127 47754
rect 10191 47690 10846 47754
rect 10910 47690 11565 47754
rect 11629 47690 12284 47754
rect 12348 47690 13003 47754
rect 13067 47690 13088 47754
rect 5916 47674 13088 47690
rect 5916 47610 6532 47674
rect 6596 47610 7251 47674
rect 7315 47610 7970 47674
rect 8034 47610 8689 47674
rect 8753 47610 9408 47674
rect 9472 47610 10127 47674
rect 10191 47610 10846 47674
rect 10910 47610 11565 47674
rect 11629 47610 12284 47674
rect 12348 47610 13003 47674
rect 13067 47610 13088 47674
rect 5916 47594 13088 47610
rect 5916 47530 6532 47594
rect 6596 47530 7251 47594
rect 7315 47530 7970 47594
rect 8034 47530 8689 47594
rect 8753 47530 9408 47594
rect 9472 47530 10127 47594
rect 10191 47530 10846 47594
rect 10910 47530 11565 47594
rect 11629 47530 12284 47594
rect 12348 47530 13003 47594
rect 13067 47530 13088 47594
rect 5916 47514 13088 47530
rect 5916 47450 6532 47514
rect 6596 47450 7251 47514
rect 7315 47450 7970 47514
rect 8034 47450 8689 47514
rect 8753 47450 9408 47514
rect 9472 47450 10127 47514
rect 10191 47450 10846 47514
rect 10910 47450 11565 47514
rect 11629 47450 12284 47514
rect 12348 47450 13003 47514
rect 13067 47450 13088 47514
rect 5916 47422 13088 47450
rect 13364 48710 20536 48722
rect 13364 48654 13396 48710
rect 13452 48654 13476 48710
rect 13532 48694 20536 48710
rect 13532 48654 13980 48694
rect 13364 48630 13980 48654
rect 14044 48630 14699 48694
rect 14763 48630 15418 48694
rect 15482 48630 16137 48694
rect 16201 48630 16856 48694
rect 16920 48630 17575 48694
rect 17639 48630 18294 48694
rect 18358 48630 19013 48694
rect 19077 48630 19732 48694
rect 19796 48630 20451 48694
rect 20515 48630 20536 48694
rect 13364 48614 20536 48630
rect 13364 48550 13980 48614
rect 14044 48550 14699 48614
rect 14763 48550 15418 48614
rect 15482 48550 16137 48614
rect 16201 48550 16856 48614
rect 16920 48550 17575 48614
rect 17639 48550 18294 48614
rect 18358 48550 19013 48614
rect 19077 48550 19732 48614
rect 19796 48550 20451 48614
rect 20515 48550 20536 48614
rect 13364 48534 20536 48550
rect 13364 48470 13980 48534
rect 14044 48470 14699 48534
rect 14763 48470 15418 48534
rect 15482 48470 16137 48534
rect 16201 48470 16856 48534
rect 16920 48470 17575 48534
rect 17639 48470 18294 48534
rect 18358 48470 19013 48534
rect 19077 48470 19732 48534
rect 19796 48470 20451 48534
rect 20515 48470 20536 48534
rect 13364 48454 20536 48470
rect 13364 48390 13980 48454
rect 14044 48390 14699 48454
rect 14763 48390 15418 48454
rect 15482 48390 16137 48454
rect 16201 48390 16856 48454
rect 16920 48390 17575 48454
rect 17639 48390 18294 48454
rect 18358 48390 19013 48454
rect 19077 48390 19732 48454
rect 19796 48390 20451 48454
rect 20515 48390 20536 48454
rect 13364 48374 20536 48390
rect 13364 48310 13980 48374
rect 14044 48310 14699 48374
rect 14763 48310 15418 48374
rect 15482 48310 16137 48374
rect 16201 48310 16856 48374
rect 16920 48310 17575 48374
rect 17639 48310 18294 48374
rect 18358 48310 19013 48374
rect 19077 48310 19732 48374
rect 19796 48310 20451 48374
rect 20515 48310 20536 48374
rect 13364 48294 20536 48310
rect 13364 48230 13980 48294
rect 14044 48230 14699 48294
rect 14763 48230 15418 48294
rect 15482 48230 16137 48294
rect 16201 48230 16856 48294
rect 16920 48230 17575 48294
rect 17639 48230 18294 48294
rect 18358 48230 19013 48294
rect 19077 48230 19732 48294
rect 19796 48230 20451 48294
rect 20515 48230 20536 48294
rect 13364 48214 20536 48230
rect 13364 48150 13980 48214
rect 14044 48150 14699 48214
rect 14763 48150 15418 48214
rect 15482 48150 16137 48214
rect 16201 48150 16856 48214
rect 16920 48150 17575 48214
rect 17639 48150 18294 48214
rect 18358 48150 19013 48214
rect 19077 48150 19732 48214
rect 19796 48150 20451 48214
rect 20515 48150 20536 48214
rect 13364 47994 20536 48150
rect 13364 47930 13980 47994
rect 14044 47930 14699 47994
rect 14763 47930 15418 47994
rect 15482 47930 16137 47994
rect 16201 47930 16856 47994
rect 16920 47930 17575 47994
rect 17639 47930 18294 47994
rect 18358 47930 19013 47994
rect 19077 47930 19732 47994
rect 19796 47930 20451 47994
rect 20515 47930 20536 47994
rect 13364 47914 20536 47930
rect 13364 47850 13980 47914
rect 14044 47850 14699 47914
rect 14763 47850 15418 47914
rect 15482 47850 16137 47914
rect 16201 47850 16856 47914
rect 16920 47850 17575 47914
rect 17639 47850 18294 47914
rect 18358 47850 19013 47914
rect 19077 47850 19732 47914
rect 19796 47850 20451 47914
rect 20515 47850 20536 47914
rect 13364 47834 20536 47850
rect 13364 47770 13980 47834
rect 14044 47770 14699 47834
rect 14763 47770 15418 47834
rect 15482 47770 16137 47834
rect 16201 47770 16856 47834
rect 16920 47770 17575 47834
rect 17639 47770 18294 47834
rect 18358 47770 19013 47834
rect 19077 47770 19732 47834
rect 19796 47770 20451 47834
rect 20515 47770 20536 47834
rect 13364 47754 20536 47770
rect 13364 47690 13980 47754
rect 14044 47690 14699 47754
rect 14763 47690 15418 47754
rect 15482 47690 16137 47754
rect 16201 47690 16856 47754
rect 16920 47690 17575 47754
rect 17639 47690 18294 47754
rect 18358 47690 19013 47754
rect 19077 47690 19732 47754
rect 19796 47690 20451 47754
rect 20515 47690 20536 47754
rect 13364 47674 20536 47690
rect 13364 47610 13980 47674
rect 14044 47610 14699 47674
rect 14763 47610 15418 47674
rect 15482 47610 16137 47674
rect 16201 47610 16856 47674
rect 16920 47610 17575 47674
rect 17639 47610 18294 47674
rect 18358 47610 19013 47674
rect 19077 47610 19732 47674
rect 19796 47610 20451 47674
rect 20515 47610 20536 47674
rect 13364 47594 20536 47610
rect 13364 47530 13980 47594
rect 14044 47530 14699 47594
rect 14763 47530 15418 47594
rect 15482 47530 16137 47594
rect 16201 47530 16856 47594
rect 16920 47530 17575 47594
rect 17639 47530 18294 47594
rect 18358 47530 19013 47594
rect 19077 47530 19732 47594
rect 19796 47530 20451 47594
rect 20515 47530 20536 47594
rect 13364 47514 20536 47530
rect 13364 47450 13980 47514
rect 14044 47450 14699 47514
rect 14763 47450 15418 47514
rect 15482 47450 16137 47514
rect 16201 47450 16856 47514
rect 16920 47450 17575 47514
rect 17639 47450 18294 47514
rect 18358 47450 19013 47514
rect 19077 47450 19732 47514
rect 19796 47450 20451 47514
rect 20515 47450 20536 47514
rect 13364 47422 20536 47450
rect 5918 47294 6118 47322
rect 5918 47230 5946 47294
rect 6010 47290 6026 47294
rect 6010 47230 6026 47234
rect 6090 47230 6118 47294
rect 5918 47202 6118 47230
rect 13366 47294 13566 47322
rect 13366 47230 13394 47294
rect 13458 47290 13474 47294
rect 13458 47230 13474 47234
rect 13538 47230 13566 47294
rect 13366 47202 13566 47230
rect 17677 47136 17743 47137
rect 17672 47134 17678 47136
rect 900 47104 2532 47132
rect 900 47040 924 47104
rect 988 47040 1004 47104
rect 1068 47040 1084 47104
rect 1148 47040 1164 47104
rect 1228 47040 1244 47104
rect 1308 47040 1324 47104
rect 1388 47040 1404 47104
rect 1468 47040 1484 47104
rect 1548 47040 1564 47104
rect 1628 47040 1644 47104
rect 1708 47040 1724 47104
rect 1788 47040 1804 47104
rect 1868 47040 1884 47104
rect 1948 47040 1964 47104
rect 2028 47040 2044 47104
rect 2108 47040 2124 47104
rect 2188 47040 2204 47104
rect 2268 47040 2284 47104
rect 2348 47040 2364 47104
rect 2428 47040 2444 47104
rect 2508 47040 2532 47104
rect 17588 47074 17678 47134
rect 17672 47072 17678 47074
rect 17742 47072 17748 47136
rect 55904 47104 57536 47132
rect 17677 47071 17743 47072
rect 900 47012 2532 47040
rect 55904 47040 55928 47104
rect 55992 47040 56008 47104
rect 56072 47040 56088 47104
rect 56152 47040 56168 47104
rect 56232 47040 56248 47104
rect 56312 47040 56328 47104
rect 56392 47040 56408 47104
rect 56472 47040 56488 47104
rect 56552 47040 56568 47104
rect 56632 47040 56648 47104
rect 56712 47040 56728 47104
rect 56792 47040 56808 47104
rect 56872 47040 56888 47104
rect 56952 47040 56968 47104
rect 57032 47040 57048 47104
rect 57112 47040 57128 47104
rect 57192 47040 57208 47104
rect 57272 47040 57288 47104
rect 57352 47040 57368 47104
rect 57432 47040 57448 47104
rect 57512 47040 57536 47104
rect 55904 47012 57536 47040
rect 3348 45224 4980 45252
rect 3348 45160 3372 45224
rect 3436 45160 3452 45224
rect 3516 45160 3532 45224
rect 3596 45160 3612 45224
rect 3676 45160 3692 45224
rect 3756 45160 3772 45224
rect 3836 45160 3852 45224
rect 3916 45160 3932 45224
rect 3996 45160 4012 45224
rect 4076 45160 4092 45224
rect 4156 45160 4172 45224
rect 4236 45160 4252 45224
rect 4316 45160 4332 45224
rect 4396 45160 4412 45224
rect 4476 45160 4492 45224
rect 4556 45160 4572 45224
rect 4636 45160 4652 45224
rect 4716 45160 4732 45224
rect 4796 45160 4812 45224
rect 4876 45160 4892 45224
rect 4956 45160 4980 45224
rect 3348 45132 4980 45160
rect 53456 45224 55088 45252
rect 53456 45160 53480 45224
rect 53544 45160 53560 45224
rect 53624 45160 53640 45224
rect 53704 45160 53720 45224
rect 53784 45160 53800 45224
rect 53864 45160 53880 45224
rect 53944 45160 53960 45224
rect 54024 45160 54040 45224
rect 54104 45160 54120 45224
rect 54184 45160 54200 45224
rect 54264 45160 54280 45224
rect 54344 45160 54360 45224
rect 54424 45160 54440 45224
rect 54504 45160 54520 45224
rect 54584 45160 54600 45224
rect 54664 45160 54680 45224
rect 54744 45160 54760 45224
rect 54824 45160 54840 45224
rect 54904 45160 54920 45224
rect 54984 45160 55000 45224
rect 55064 45160 55088 45224
rect 53456 45132 55088 45160
rect 5916 44950 13088 44962
rect 5916 44894 5948 44950
rect 6004 44894 6028 44950
rect 6084 44934 13088 44950
rect 6084 44894 6532 44934
rect 5916 44870 6532 44894
rect 6596 44870 7251 44934
rect 7315 44870 7970 44934
rect 8034 44870 8689 44934
rect 8753 44870 9408 44934
rect 9472 44870 10127 44934
rect 10191 44870 10846 44934
rect 10910 44870 11565 44934
rect 11629 44870 12284 44934
rect 12348 44870 13003 44934
rect 13067 44870 13088 44934
rect 5916 44854 13088 44870
rect 5916 44790 6532 44854
rect 6596 44790 7251 44854
rect 7315 44790 7970 44854
rect 8034 44790 8689 44854
rect 8753 44790 9408 44854
rect 9472 44790 10127 44854
rect 10191 44790 10846 44854
rect 10910 44790 11565 44854
rect 11629 44790 12284 44854
rect 12348 44790 13003 44854
rect 13067 44790 13088 44854
rect 5916 44774 13088 44790
rect 5916 44710 6532 44774
rect 6596 44710 7251 44774
rect 7315 44710 7970 44774
rect 8034 44710 8689 44774
rect 8753 44710 9408 44774
rect 9472 44710 10127 44774
rect 10191 44710 10846 44774
rect 10910 44710 11565 44774
rect 11629 44710 12284 44774
rect 12348 44710 13003 44774
rect 13067 44710 13088 44774
rect 5916 44694 13088 44710
rect 5916 44630 6532 44694
rect 6596 44630 7251 44694
rect 7315 44630 7970 44694
rect 8034 44630 8689 44694
rect 8753 44630 9408 44694
rect 9472 44630 10127 44694
rect 10191 44630 10846 44694
rect 10910 44630 11565 44694
rect 11629 44630 12284 44694
rect 12348 44630 13003 44694
rect 13067 44630 13088 44694
rect 5916 44614 13088 44630
rect 5916 44550 6532 44614
rect 6596 44550 7251 44614
rect 7315 44550 7970 44614
rect 8034 44550 8689 44614
rect 8753 44550 9408 44614
rect 9472 44550 10127 44614
rect 10191 44550 10846 44614
rect 10910 44550 11565 44614
rect 11629 44550 12284 44614
rect 12348 44550 13003 44614
rect 13067 44550 13088 44614
rect 5916 44534 13088 44550
rect 5916 44470 6532 44534
rect 6596 44470 7251 44534
rect 7315 44470 7970 44534
rect 8034 44470 8689 44534
rect 8753 44470 9408 44534
rect 9472 44470 10127 44534
rect 10191 44470 10846 44534
rect 10910 44470 11565 44534
rect 11629 44470 12284 44534
rect 12348 44470 13003 44534
rect 13067 44470 13088 44534
rect 5916 44454 13088 44470
rect 5916 44390 6532 44454
rect 6596 44390 7251 44454
rect 7315 44390 7970 44454
rect 8034 44390 8689 44454
rect 8753 44390 9408 44454
rect 9472 44390 10127 44454
rect 10191 44390 10846 44454
rect 10910 44390 11565 44454
rect 11629 44390 12284 44454
rect 12348 44390 13003 44454
rect 13067 44390 13088 44454
rect 5916 44234 13088 44390
rect 5916 44170 6532 44234
rect 6596 44170 7251 44234
rect 7315 44170 7970 44234
rect 8034 44170 8689 44234
rect 8753 44170 9408 44234
rect 9472 44170 10127 44234
rect 10191 44170 10846 44234
rect 10910 44170 11565 44234
rect 11629 44170 12284 44234
rect 12348 44170 13003 44234
rect 13067 44170 13088 44234
rect 5916 44154 13088 44170
rect 5916 44090 6532 44154
rect 6596 44090 7251 44154
rect 7315 44090 7970 44154
rect 8034 44090 8689 44154
rect 8753 44090 9408 44154
rect 9472 44090 10127 44154
rect 10191 44090 10846 44154
rect 10910 44090 11565 44154
rect 11629 44090 12284 44154
rect 12348 44090 13003 44154
rect 13067 44090 13088 44154
rect 5916 44074 13088 44090
rect 5916 44010 6532 44074
rect 6596 44010 7251 44074
rect 7315 44010 7970 44074
rect 8034 44010 8689 44074
rect 8753 44010 9408 44074
rect 9472 44010 10127 44074
rect 10191 44010 10846 44074
rect 10910 44010 11565 44074
rect 11629 44010 12284 44074
rect 12348 44010 13003 44074
rect 13067 44010 13088 44074
rect 5916 43994 13088 44010
rect 5916 43930 6532 43994
rect 6596 43930 7251 43994
rect 7315 43930 7970 43994
rect 8034 43930 8689 43994
rect 8753 43930 9408 43994
rect 9472 43930 10127 43994
rect 10191 43930 10846 43994
rect 10910 43930 11565 43994
rect 11629 43930 12284 43994
rect 12348 43930 13003 43994
rect 13067 43930 13088 43994
rect 5916 43914 13088 43930
rect 5916 43850 6532 43914
rect 6596 43850 7251 43914
rect 7315 43850 7970 43914
rect 8034 43850 8689 43914
rect 8753 43850 9408 43914
rect 9472 43850 10127 43914
rect 10191 43850 10846 43914
rect 10910 43850 11565 43914
rect 11629 43850 12284 43914
rect 12348 43850 13003 43914
rect 13067 43850 13088 43914
rect 5916 43834 13088 43850
rect 5916 43770 6532 43834
rect 6596 43770 7251 43834
rect 7315 43770 7970 43834
rect 8034 43770 8689 43834
rect 8753 43770 9408 43834
rect 9472 43770 10127 43834
rect 10191 43770 10846 43834
rect 10910 43770 11565 43834
rect 11629 43770 12284 43834
rect 12348 43770 13003 43834
rect 13067 43770 13088 43834
rect 13394 43778 13400 43842
rect 13464 43840 13470 43842
rect 15009 43840 15075 43843
rect 13464 43838 15075 43840
rect 13464 43782 15014 43838
rect 15070 43782 15075 43838
rect 13464 43780 15075 43782
rect 13464 43778 13470 43780
rect 15009 43777 15075 43780
rect 5916 43754 13088 43770
rect 5916 43690 6532 43754
rect 6596 43690 7251 43754
rect 7315 43690 7970 43754
rect 8034 43690 8689 43754
rect 8753 43690 9408 43754
rect 9472 43690 10127 43754
rect 10191 43690 10846 43754
rect 10910 43690 11565 43754
rect 11629 43690 12284 43754
rect 12348 43690 13003 43754
rect 13067 43690 13088 43754
rect 5916 43662 13088 43690
rect 5918 43534 6118 43562
rect 5918 43470 5946 43534
rect 6010 43530 6026 43534
rect 6010 43470 6026 43474
rect 6090 43470 6118 43534
rect 5918 43442 6118 43470
rect 14549 43474 14615 43477
rect 23749 43474 23815 43477
rect 14549 43472 23815 43474
rect 14549 43416 14554 43472
rect 14610 43416 23754 43472
rect 23810 43416 23815 43472
rect 14549 43414 23815 43416
rect 14549 43411 14615 43414
rect 23749 43411 23815 43414
rect 900 43344 2532 43372
rect 8293 43354 8359 43355
rect 900 43280 924 43344
rect 988 43280 1004 43344
rect 1068 43280 1084 43344
rect 1148 43280 1164 43344
rect 1228 43280 1244 43344
rect 1308 43280 1324 43344
rect 1388 43280 1404 43344
rect 1468 43280 1484 43344
rect 1548 43280 1564 43344
rect 1628 43280 1644 43344
rect 1708 43280 1724 43344
rect 1788 43280 1804 43344
rect 1868 43280 1884 43344
rect 1948 43280 1964 43344
rect 2028 43280 2044 43344
rect 2108 43280 2124 43344
rect 2188 43280 2204 43344
rect 2268 43280 2284 43344
rect 2348 43280 2364 43344
rect 2428 43280 2444 43344
rect 2508 43280 2532 43344
rect 8288 43290 8294 43354
rect 8358 43352 8364 43354
rect 8358 43292 8448 43352
rect 55904 43344 57536 43372
rect 8358 43290 8364 43292
rect 8293 43289 8359 43290
rect 900 43252 2532 43280
rect 55904 43280 55928 43344
rect 55992 43280 56008 43344
rect 56072 43280 56088 43344
rect 56152 43280 56168 43344
rect 56232 43280 56248 43344
rect 56312 43280 56328 43344
rect 56392 43280 56408 43344
rect 56472 43280 56488 43344
rect 56552 43280 56568 43344
rect 56632 43280 56648 43344
rect 56712 43280 56728 43344
rect 56792 43280 56808 43344
rect 56872 43280 56888 43344
rect 56952 43280 56968 43344
rect 57032 43280 57048 43344
rect 57112 43280 57128 43344
rect 57192 43280 57208 43344
rect 57272 43280 57288 43344
rect 57352 43280 57368 43344
rect 57432 43280 57448 43344
rect 57512 43280 57536 43344
rect 55904 43252 57536 43280
rect 3348 41464 4980 41492
rect 3348 41400 3372 41464
rect 3436 41400 3452 41464
rect 3516 41400 3532 41464
rect 3596 41400 3612 41464
rect 3676 41400 3692 41464
rect 3756 41400 3772 41464
rect 3836 41400 3852 41464
rect 3916 41400 3932 41464
rect 3996 41400 4012 41464
rect 4076 41400 4092 41464
rect 4156 41400 4172 41464
rect 4236 41400 4252 41464
rect 4316 41400 4332 41464
rect 4396 41400 4412 41464
rect 4476 41400 4492 41464
rect 4556 41400 4572 41464
rect 4636 41400 4652 41464
rect 4716 41400 4732 41464
rect 4796 41400 4812 41464
rect 4876 41400 4892 41464
rect 4956 41400 4980 41464
rect 53456 41464 55088 41492
rect 22185 41402 22251 41403
rect 6908 41400 6914 41402
rect 3348 41372 4980 41400
rect 5168 41340 6914 41400
rect 5168 41034 5228 41340
rect 6908 41338 6914 41340
rect 6978 41338 6984 41402
rect 22185 41400 22232 41402
rect 22142 41398 22232 41400
rect 22142 41342 22190 41398
rect 22142 41340 22232 41342
rect 22185 41338 22232 41340
rect 22296 41338 22302 41402
rect 53456 41400 53480 41464
rect 53544 41400 53560 41464
rect 53624 41400 53640 41464
rect 53704 41400 53720 41464
rect 53784 41400 53800 41464
rect 53864 41400 53880 41464
rect 53944 41400 53960 41464
rect 54024 41400 54040 41464
rect 54104 41400 54120 41464
rect 54184 41400 54200 41464
rect 54264 41400 54280 41464
rect 54344 41400 54360 41464
rect 54424 41400 54440 41464
rect 54504 41400 54520 41464
rect 54584 41400 54600 41464
rect 54664 41400 54680 41464
rect 54744 41400 54760 41464
rect 54824 41400 54840 41464
rect 54904 41400 54920 41464
rect 54984 41400 55000 41464
rect 55064 41400 55088 41464
rect 53456 41372 55088 41400
rect 22185 41337 22251 41338
rect 0 40974 5228 41034
rect 6308 41190 13480 41202
rect 6308 41134 6340 41190
rect 6396 41134 6420 41190
rect 6476 41174 13480 41190
rect 6476 41134 6924 41174
rect 6308 41110 6924 41134
rect 6988 41110 7643 41174
rect 7707 41110 8362 41174
rect 8426 41110 9081 41174
rect 9145 41110 9800 41174
rect 9864 41110 10519 41174
rect 10583 41110 11238 41174
rect 11302 41110 11957 41174
rect 12021 41110 12676 41174
rect 12740 41110 13395 41174
rect 13459 41110 13480 41174
rect 6308 41094 13480 41110
rect 6308 41030 6924 41094
rect 6988 41030 7643 41094
rect 7707 41030 8362 41094
rect 8426 41030 9081 41094
rect 9145 41030 9800 41094
rect 9864 41030 10519 41094
rect 10583 41030 11238 41094
rect 11302 41030 11957 41094
rect 12021 41030 12676 41094
rect 12740 41030 13395 41094
rect 13459 41030 13480 41094
rect 6308 41014 13480 41030
rect 6308 40950 6924 41014
rect 6988 40950 7643 41014
rect 7707 40950 8362 41014
rect 8426 40950 9081 41014
rect 9145 40950 9800 41014
rect 9864 40950 10519 41014
rect 10583 40950 11238 41014
rect 11302 40950 11957 41014
rect 12021 40950 12676 41014
rect 12740 40950 13395 41014
rect 13459 40950 13480 41014
rect 6308 40934 13480 40950
rect 6308 40870 6924 40934
rect 6988 40870 7643 40934
rect 7707 40870 8362 40934
rect 8426 40870 9081 40934
rect 9145 40870 9800 40934
rect 9864 40870 10519 40934
rect 10583 40870 11238 40934
rect 11302 40870 11957 40934
rect 12021 40870 12676 40934
rect 12740 40870 13395 40934
rect 13459 40870 13480 40934
rect 6308 40854 13480 40870
rect 6308 40790 6924 40854
rect 6988 40790 7643 40854
rect 7707 40790 8362 40854
rect 8426 40790 9081 40854
rect 9145 40790 9800 40854
rect 9864 40790 10519 40854
rect 10583 40790 11238 40854
rect 11302 40790 11957 40854
rect 12021 40790 12676 40854
rect 12740 40790 13395 40854
rect 13459 40790 13480 40854
rect 6308 40774 13480 40790
rect 6308 40710 6924 40774
rect 6988 40710 7643 40774
rect 7707 40710 8362 40774
rect 8426 40710 9081 40774
rect 9145 40710 9800 40774
rect 9864 40710 10519 40774
rect 10583 40710 11238 40774
rect 11302 40710 11957 40774
rect 12021 40710 12676 40774
rect 12740 40710 13395 40774
rect 13459 40710 13480 40774
rect 6308 40694 13480 40710
rect 6308 40630 6924 40694
rect 6988 40630 7643 40694
rect 7707 40630 8362 40694
rect 8426 40630 9081 40694
rect 9145 40630 9800 40694
rect 9864 40630 10519 40694
rect 10583 40630 11238 40694
rect 11302 40630 11957 40694
rect 12021 40630 12676 40694
rect 12740 40630 13395 40694
rect 13459 40630 13480 40694
rect 6308 40474 13480 40630
rect 6308 40410 6924 40474
rect 6988 40410 7643 40474
rect 7707 40410 8362 40474
rect 8426 40410 9081 40474
rect 9145 40410 9800 40474
rect 9864 40410 10519 40474
rect 10583 40410 11238 40474
rect 11302 40410 11957 40474
rect 12021 40410 12676 40474
rect 12740 40410 13395 40474
rect 13459 40410 13480 40474
rect 6308 40394 13480 40410
rect 6308 40330 6924 40394
rect 6988 40330 7643 40394
rect 7707 40330 8362 40394
rect 8426 40330 9081 40394
rect 9145 40330 9800 40394
rect 9864 40330 10519 40394
rect 10583 40330 11238 40394
rect 11302 40330 11957 40394
rect 12021 40330 12676 40394
rect 12740 40330 13395 40394
rect 13459 40330 13480 40394
rect 6308 40314 13480 40330
rect 6308 40250 6924 40314
rect 6988 40250 7643 40314
rect 7707 40250 8362 40314
rect 8426 40250 9081 40314
rect 9145 40250 9800 40314
rect 9864 40250 10519 40314
rect 10583 40250 11238 40314
rect 11302 40250 11957 40314
rect 12021 40250 12676 40314
rect 12740 40250 13395 40314
rect 13459 40250 13480 40314
rect 6308 40234 13480 40250
rect 6308 40170 6924 40234
rect 6988 40170 7643 40234
rect 7707 40170 8362 40234
rect 8426 40170 9081 40234
rect 9145 40170 9800 40234
rect 9864 40170 10519 40234
rect 10583 40170 11238 40234
rect 11302 40170 11957 40234
rect 12021 40170 12676 40234
rect 12740 40170 13395 40234
rect 13459 40170 13480 40234
rect 6308 40154 13480 40170
rect 6308 40090 6924 40154
rect 6988 40090 7643 40154
rect 7707 40090 8362 40154
rect 8426 40090 9081 40154
rect 9145 40090 9800 40154
rect 9864 40090 10519 40154
rect 10583 40090 11238 40154
rect 11302 40090 11957 40154
rect 12021 40090 12676 40154
rect 12740 40090 13395 40154
rect 13459 40090 13480 40154
rect 6308 40074 13480 40090
rect 6308 40010 6924 40074
rect 6988 40010 7643 40074
rect 7707 40010 8362 40074
rect 8426 40010 9081 40074
rect 9145 40010 9800 40074
rect 9864 40010 10519 40074
rect 10583 40010 11238 40074
rect 11302 40010 11957 40074
rect 12021 40010 12676 40074
rect 12740 40010 13395 40074
rect 13459 40010 13480 40074
rect 6308 39994 13480 40010
rect 6308 39930 6924 39994
rect 6988 39930 7643 39994
rect 7707 39930 8362 39994
rect 8426 39930 9081 39994
rect 9145 39930 9800 39994
rect 9864 39930 10519 39994
rect 10583 39930 11238 39994
rect 11302 39930 11957 39994
rect 12021 39930 12676 39994
rect 12740 39930 13395 39994
rect 13459 39930 13480 39994
rect 6308 39902 13480 39930
rect 15128 41190 22300 41202
rect 15128 41134 15160 41190
rect 15216 41134 15240 41190
rect 15296 41174 22300 41190
rect 15296 41134 15744 41174
rect 15128 41110 15744 41134
rect 15808 41110 16463 41174
rect 16527 41110 17182 41174
rect 17246 41110 17901 41174
rect 17965 41110 18620 41174
rect 18684 41110 19339 41174
rect 19403 41110 20058 41174
rect 20122 41110 20777 41174
rect 20841 41110 21496 41174
rect 21560 41110 22215 41174
rect 22279 41110 22300 41174
rect 15128 41094 22300 41110
rect 15128 41030 15744 41094
rect 15808 41030 16463 41094
rect 16527 41030 17182 41094
rect 17246 41030 17901 41094
rect 17965 41030 18620 41094
rect 18684 41030 19339 41094
rect 19403 41030 20058 41094
rect 20122 41030 20777 41094
rect 20841 41030 21496 41094
rect 21560 41030 22215 41094
rect 22279 41030 22300 41094
rect 15128 41014 22300 41030
rect 15128 40950 15744 41014
rect 15808 40950 16463 41014
rect 16527 40950 17182 41014
rect 17246 40950 17901 41014
rect 17965 40950 18620 41014
rect 18684 40950 19339 41014
rect 19403 40950 20058 41014
rect 20122 40950 20777 41014
rect 20841 40950 21496 41014
rect 21560 40950 22215 41014
rect 22279 40950 22300 41014
rect 15128 40934 22300 40950
rect 15128 40870 15744 40934
rect 15808 40870 16463 40934
rect 16527 40870 17182 40934
rect 17246 40870 17901 40934
rect 17965 40870 18620 40934
rect 18684 40870 19339 40934
rect 19403 40870 20058 40934
rect 20122 40870 20777 40934
rect 20841 40870 21496 40934
rect 21560 40870 22215 40934
rect 22279 40870 22300 40934
rect 15128 40854 22300 40870
rect 15128 40790 15744 40854
rect 15808 40790 16463 40854
rect 16527 40790 17182 40854
rect 17246 40790 17901 40854
rect 17965 40790 18620 40854
rect 18684 40790 19339 40854
rect 19403 40790 20058 40854
rect 20122 40790 20777 40854
rect 20841 40790 21496 40854
rect 21560 40790 22215 40854
rect 22279 40790 22300 40854
rect 15128 40774 22300 40790
rect 15128 40710 15744 40774
rect 15808 40710 16463 40774
rect 16527 40710 17182 40774
rect 17246 40710 17901 40774
rect 17965 40710 18620 40774
rect 18684 40710 19339 40774
rect 19403 40710 20058 40774
rect 20122 40710 20777 40774
rect 20841 40710 21496 40774
rect 21560 40710 22215 40774
rect 22279 40710 22300 40774
rect 15128 40694 22300 40710
rect 15128 40630 15744 40694
rect 15808 40630 16463 40694
rect 16527 40630 17182 40694
rect 17246 40630 17901 40694
rect 17965 40630 18620 40694
rect 18684 40630 19339 40694
rect 19403 40630 20058 40694
rect 20122 40630 20777 40694
rect 20841 40630 21496 40694
rect 21560 40630 22215 40694
rect 22279 40630 22300 40694
rect 15128 40474 22300 40630
rect 15128 40410 15744 40474
rect 15808 40410 16463 40474
rect 16527 40410 17182 40474
rect 17246 40410 17901 40474
rect 17965 40410 18620 40474
rect 18684 40410 19339 40474
rect 19403 40410 20058 40474
rect 20122 40410 20777 40474
rect 20841 40410 21496 40474
rect 21560 40410 22215 40474
rect 22279 40410 22300 40474
rect 15128 40394 22300 40410
rect 15128 40330 15744 40394
rect 15808 40330 16463 40394
rect 16527 40330 17182 40394
rect 17246 40330 17901 40394
rect 17965 40330 18620 40394
rect 18684 40330 19339 40394
rect 19403 40330 20058 40394
rect 20122 40330 20777 40394
rect 20841 40330 21496 40394
rect 21560 40330 22215 40394
rect 22279 40330 22300 40394
rect 15128 40314 22300 40330
rect 15128 40250 15744 40314
rect 15808 40250 16463 40314
rect 16527 40250 17182 40314
rect 17246 40250 17901 40314
rect 17965 40250 18620 40314
rect 18684 40250 19339 40314
rect 19403 40250 20058 40314
rect 20122 40250 20777 40314
rect 20841 40250 21496 40314
rect 21560 40250 22215 40314
rect 22279 40250 22300 40314
rect 15128 40234 22300 40250
rect 15128 40170 15744 40234
rect 15808 40170 16463 40234
rect 16527 40170 17182 40234
rect 17246 40170 17901 40234
rect 17965 40170 18620 40234
rect 18684 40170 19339 40234
rect 19403 40170 20058 40234
rect 20122 40170 20777 40234
rect 20841 40170 21496 40234
rect 21560 40170 22215 40234
rect 22279 40170 22300 40234
rect 15128 40154 22300 40170
rect 15128 40090 15744 40154
rect 15808 40090 16463 40154
rect 16527 40090 17182 40154
rect 17246 40090 17901 40154
rect 17965 40090 18620 40154
rect 18684 40090 19339 40154
rect 19403 40090 20058 40154
rect 20122 40090 20777 40154
rect 20841 40090 21496 40154
rect 21560 40090 22215 40154
rect 22279 40090 22300 40154
rect 15128 40074 22300 40090
rect 15128 40010 15744 40074
rect 15808 40010 16463 40074
rect 16527 40010 17182 40074
rect 17246 40010 17901 40074
rect 17965 40010 18620 40074
rect 18684 40010 19339 40074
rect 19403 40010 20058 40074
rect 20122 40010 20777 40074
rect 20841 40010 21496 40074
rect 21560 40010 22215 40074
rect 22279 40010 22300 40074
rect 15128 39994 22300 40010
rect 15128 39930 15744 39994
rect 15808 39930 16463 39994
rect 16527 39930 17182 39994
rect 17246 39930 17901 39994
rect 17965 39930 18620 39994
rect 18684 39930 19339 39994
rect 19403 39930 20058 39994
rect 20122 39930 20777 39994
rect 20841 39930 21496 39994
rect 21560 39930 22215 39994
rect 22279 39930 22300 39994
rect 15128 39902 22300 39930
rect 6310 39774 6510 39802
rect 6310 39710 6338 39774
rect 6402 39770 6418 39774
rect 6402 39710 6418 39714
rect 6482 39710 6510 39774
rect 6310 39682 6510 39710
rect 15130 39774 15330 39802
rect 15130 39710 15158 39774
rect 15222 39770 15238 39774
rect 15222 39710 15238 39714
rect 15302 39710 15330 39774
rect 15130 39682 15330 39710
rect 15469 39694 15535 39695
rect 15464 39630 15470 39694
rect 15534 39692 15540 39694
rect 15534 39632 15624 39692
rect 15534 39630 15540 39632
rect 15469 39629 15535 39630
rect 900 39584 2532 39612
rect 900 39520 924 39584
rect 988 39520 1004 39584
rect 1068 39520 1084 39584
rect 1148 39520 1164 39584
rect 1228 39520 1244 39584
rect 1308 39520 1324 39584
rect 1388 39520 1404 39584
rect 1468 39520 1484 39584
rect 1548 39520 1564 39584
rect 1628 39520 1644 39584
rect 1708 39520 1724 39584
rect 1788 39520 1804 39584
rect 1868 39520 1884 39584
rect 1948 39520 1964 39584
rect 2028 39520 2044 39584
rect 2108 39520 2124 39584
rect 2188 39520 2204 39584
rect 2268 39520 2284 39584
rect 2348 39520 2364 39584
rect 2428 39520 2444 39584
rect 2508 39520 2532 39584
rect 900 39492 2532 39520
rect 55904 39584 57536 39612
rect 55904 39520 55928 39584
rect 55992 39520 56008 39584
rect 56072 39520 56088 39584
rect 56152 39520 56168 39584
rect 56232 39520 56248 39584
rect 56312 39520 56328 39584
rect 56392 39520 56408 39584
rect 56472 39520 56488 39584
rect 56552 39520 56568 39584
rect 56632 39520 56648 39584
rect 56712 39520 56728 39584
rect 56792 39520 56808 39584
rect 56872 39520 56888 39584
rect 56952 39520 56968 39584
rect 57032 39520 57048 39584
rect 57112 39520 57128 39584
rect 57192 39520 57208 39584
rect 57272 39520 57288 39584
rect 57352 39520 57368 39584
rect 57432 39520 57448 39584
rect 57512 39520 57536 39584
rect 55904 39492 57536 39520
rect 3348 37704 4980 37732
rect 3348 37640 3372 37704
rect 3436 37640 3452 37704
rect 3516 37640 3532 37704
rect 3596 37640 3612 37704
rect 3676 37640 3692 37704
rect 3756 37640 3772 37704
rect 3836 37640 3852 37704
rect 3916 37640 3932 37704
rect 3996 37640 4012 37704
rect 4076 37640 4092 37704
rect 4156 37640 4172 37704
rect 4236 37640 4252 37704
rect 4316 37640 4332 37704
rect 4396 37640 4412 37704
rect 4476 37640 4492 37704
rect 4556 37640 4572 37704
rect 4636 37640 4652 37704
rect 4716 37640 4732 37704
rect 4796 37640 4812 37704
rect 4876 37640 4892 37704
rect 4956 37640 4980 37704
rect 3348 37612 4980 37640
rect 53456 37704 55088 37732
rect 53456 37640 53480 37704
rect 53544 37640 53560 37704
rect 53624 37640 53640 37704
rect 53704 37640 53720 37704
rect 53784 37640 53800 37704
rect 53864 37640 53880 37704
rect 53944 37640 53960 37704
rect 54024 37640 54040 37704
rect 54104 37640 54120 37704
rect 54184 37640 54200 37704
rect 54264 37640 54280 37704
rect 54344 37640 54360 37704
rect 54424 37640 54440 37704
rect 54504 37640 54520 37704
rect 54584 37640 54600 37704
rect 54664 37640 54680 37704
rect 54744 37640 54760 37704
rect 54824 37640 54840 37704
rect 54904 37640 54920 37704
rect 54984 37640 55000 37704
rect 55064 37640 55088 37704
rect 33409 37620 33475 37621
rect 33404 37618 33410 37620
rect 33320 37558 33410 37618
rect 33404 37556 33410 37558
rect 33474 37556 33480 37620
rect 53456 37612 55088 37640
rect 33409 37555 33475 37556
rect 29926 37430 37098 37442
rect 29926 37374 29958 37430
rect 30014 37374 30038 37430
rect 30094 37414 37098 37430
rect 30094 37374 30542 37414
rect 29926 37350 30542 37374
rect 30606 37350 31261 37414
rect 31325 37350 31980 37414
rect 32044 37350 32699 37414
rect 32763 37350 33418 37414
rect 33482 37350 34137 37414
rect 34201 37350 34856 37414
rect 34920 37350 35575 37414
rect 35639 37350 36294 37414
rect 36358 37350 37013 37414
rect 37077 37350 37098 37414
rect 29926 37334 37098 37350
rect 29926 37270 30542 37334
rect 30606 37270 31261 37334
rect 31325 37270 31980 37334
rect 32044 37270 32699 37334
rect 32763 37270 33418 37334
rect 33482 37270 34137 37334
rect 34201 37270 34856 37334
rect 34920 37270 35575 37334
rect 35639 37270 36294 37334
rect 36358 37270 37013 37334
rect 37077 37270 37098 37334
rect 12893 37252 12959 37255
rect 29926 37254 37098 37270
rect 13532 37252 13538 37254
rect 12893 37250 13538 37252
rect 12893 37194 12898 37250
rect 12954 37194 13538 37250
rect 12893 37192 13538 37194
rect 12893 37189 12959 37192
rect 13532 37190 13538 37192
rect 13602 37190 13608 37254
rect 29926 37190 30542 37254
rect 30606 37190 31261 37254
rect 31325 37190 31980 37254
rect 32044 37190 32699 37254
rect 32763 37190 33418 37254
rect 33482 37190 34137 37254
rect 34201 37190 34856 37254
rect 34920 37190 35575 37254
rect 35639 37190 36294 37254
rect 36358 37190 37013 37254
rect 37077 37190 37098 37254
rect 29926 37174 37098 37190
rect 29926 37110 30542 37174
rect 30606 37110 31261 37174
rect 31325 37110 31980 37174
rect 32044 37110 32699 37174
rect 32763 37110 33418 37174
rect 33482 37110 34137 37174
rect 34201 37110 34856 37174
rect 34920 37110 35575 37174
rect 35639 37110 36294 37174
rect 36358 37110 37013 37174
rect 37077 37110 37098 37174
rect 29926 37094 37098 37110
rect 29926 37030 30542 37094
rect 30606 37030 31261 37094
rect 31325 37030 31980 37094
rect 32044 37030 32699 37094
rect 32763 37030 33418 37094
rect 33482 37030 34137 37094
rect 34201 37030 34856 37094
rect 34920 37030 35575 37094
rect 35639 37030 36294 37094
rect 36358 37030 37013 37094
rect 37077 37030 37098 37094
rect 29926 37014 37098 37030
rect 29453 37008 29519 37011
rect 29678 37008 29684 37010
rect 29453 37006 29684 37008
rect 29453 36950 29458 37006
rect 29514 36950 29684 37006
rect 29453 36948 29684 36950
rect 29453 36945 29519 36948
rect 29678 36946 29684 36948
rect 29748 36946 29754 37010
rect 29926 36950 30542 37014
rect 30606 36950 31261 37014
rect 31325 36950 31980 37014
rect 32044 36950 32699 37014
rect 32763 36950 33418 37014
rect 33482 36950 34137 37014
rect 34201 36950 34856 37014
rect 34920 36950 35575 37014
rect 35639 36950 36294 37014
rect 36358 36950 37013 37014
rect 37077 36950 37098 37014
rect 29926 36934 37098 36950
rect 29926 36870 30542 36934
rect 30606 36870 31261 36934
rect 31325 36870 31980 36934
rect 32044 36870 32699 36934
rect 32763 36870 33418 36934
rect 33482 36870 34137 36934
rect 34201 36870 34856 36934
rect 34920 36870 35575 36934
rect 35639 36870 36294 36934
rect 36358 36870 37013 36934
rect 37077 36870 37098 36934
rect 29926 36714 37098 36870
rect 29926 36650 30542 36714
rect 30606 36650 31261 36714
rect 31325 36650 31980 36714
rect 32044 36650 32699 36714
rect 32763 36650 33418 36714
rect 33482 36650 34137 36714
rect 34201 36650 34856 36714
rect 34920 36650 35575 36714
rect 35639 36650 36294 36714
rect 36358 36650 37013 36714
rect 37077 36650 37098 36714
rect 29926 36634 37098 36650
rect 29926 36570 30542 36634
rect 30606 36570 31261 36634
rect 31325 36570 31980 36634
rect 32044 36570 32699 36634
rect 32763 36570 33418 36634
rect 33482 36570 34137 36634
rect 34201 36570 34856 36634
rect 34920 36570 35575 36634
rect 35639 36570 36294 36634
rect 36358 36570 37013 36634
rect 37077 36570 37098 36634
rect 29926 36554 37098 36570
rect 29926 36490 30542 36554
rect 30606 36490 31261 36554
rect 31325 36490 31980 36554
rect 32044 36490 32699 36554
rect 32763 36490 33418 36554
rect 33482 36490 34137 36554
rect 34201 36490 34856 36554
rect 34920 36490 35575 36554
rect 35639 36490 36294 36554
rect 36358 36490 37013 36554
rect 37077 36490 37098 36554
rect 29926 36474 37098 36490
rect 29926 36410 30542 36474
rect 30606 36410 31261 36474
rect 31325 36410 31980 36474
rect 32044 36410 32699 36474
rect 32763 36410 33418 36474
rect 33482 36410 34137 36474
rect 34201 36410 34856 36474
rect 34920 36410 35575 36474
rect 35639 36410 36294 36474
rect 36358 36410 37013 36474
rect 37077 36410 37098 36474
rect 29926 36394 37098 36410
rect 29926 36330 30542 36394
rect 30606 36330 31261 36394
rect 31325 36330 31980 36394
rect 32044 36330 32699 36394
rect 32763 36330 33418 36394
rect 33482 36330 34137 36394
rect 34201 36330 34856 36394
rect 34920 36330 35575 36394
rect 35639 36330 36294 36394
rect 36358 36330 37013 36394
rect 37077 36330 37098 36394
rect 29926 36314 37098 36330
rect 29926 36250 30542 36314
rect 30606 36250 31261 36314
rect 31325 36250 31980 36314
rect 32044 36250 32699 36314
rect 32763 36250 33418 36314
rect 33482 36250 34137 36314
rect 34201 36250 34856 36314
rect 34920 36250 35575 36314
rect 35639 36250 36294 36314
rect 36358 36250 37013 36314
rect 37077 36250 37098 36314
rect 29926 36234 37098 36250
rect 29926 36170 30542 36234
rect 30606 36170 31261 36234
rect 31325 36170 31980 36234
rect 32044 36170 32699 36234
rect 32763 36170 33418 36234
rect 33482 36170 34137 36234
rect 34201 36170 34856 36234
rect 34920 36170 35575 36234
rect 35639 36170 36294 36234
rect 36358 36170 37013 36234
rect 37077 36170 37098 36234
rect 29926 36142 37098 36170
rect 29928 36014 30128 36042
rect 37549 36034 37615 36035
rect 37544 36032 37550 36034
rect 29928 35950 29956 36014
rect 30020 36010 30036 36014
rect 30020 35950 30036 35954
rect 30100 35950 30128 36014
rect 37460 35972 37550 36032
rect 37544 35970 37550 35972
rect 37614 35970 37620 36034
rect 37549 35969 37615 35970
rect 29928 35922 30128 35950
rect 900 35824 2532 35852
rect 900 35760 924 35824
rect 988 35760 1004 35824
rect 1068 35760 1084 35824
rect 1148 35760 1164 35824
rect 1228 35760 1244 35824
rect 1308 35760 1324 35824
rect 1388 35760 1404 35824
rect 1468 35760 1484 35824
rect 1548 35760 1564 35824
rect 1628 35760 1644 35824
rect 1708 35760 1724 35824
rect 1788 35760 1804 35824
rect 1868 35760 1884 35824
rect 1948 35760 1964 35824
rect 2028 35760 2044 35824
rect 2108 35760 2124 35824
rect 2188 35760 2204 35824
rect 2268 35760 2284 35824
rect 2348 35760 2364 35824
rect 2428 35760 2444 35824
rect 2508 35760 2532 35824
rect 900 35732 2532 35760
rect 55904 35824 57536 35852
rect 55904 35760 55928 35824
rect 55992 35760 56008 35824
rect 56072 35760 56088 35824
rect 56152 35760 56168 35824
rect 56232 35760 56248 35824
rect 56312 35760 56328 35824
rect 56392 35760 56408 35824
rect 56472 35760 56488 35824
rect 56552 35760 56568 35824
rect 56632 35760 56648 35824
rect 56712 35760 56728 35824
rect 56792 35760 56808 35824
rect 56872 35760 56888 35824
rect 56952 35760 56968 35824
rect 57032 35760 57048 35824
rect 57112 35760 57128 35824
rect 57192 35760 57208 35824
rect 57272 35760 57288 35824
rect 57352 35760 57368 35824
rect 57432 35760 57448 35824
rect 57512 35760 57536 35824
rect 55904 35732 57536 35760
rect 3348 33944 4980 33972
rect 3348 33880 3372 33944
rect 3436 33880 3452 33944
rect 3516 33880 3532 33944
rect 3596 33880 3612 33944
rect 3676 33880 3692 33944
rect 3756 33880 3772 33944
rect 3836 33880 3852 33944
rect 3916 33880 3932 33944
rect 3996 33880 4012 33944
rect 4076 33880 4092 33944
rect 4156 33880 4172 33944
rect 4236 33880 4252 33944
rect 4316 33880 4332 33944
rect 4396 33880 4412 33944
rect 4476 33880 4492 33944
rect 4556 33880 4572 33944
rect 4636 33880 4652 33944
rect 4716 33880 4732 33944
rect 4796 33880 4812 33944
rect 4876 33880 4892 33944
rect 4956 33880 4980 33944
rect 3348 33852 4980 33880
rect 53456 33944 55088 33972
rect 53456 33880 53480 33944
rect 53544 33880 53560 33944
rect 53624 33880 53640 33944
rect 53704 33880 53720 33944
rect 53784 33880 53800 33944
rect 53864 33880 53880 33944
rect 53944 33880 53960 33944
rect 54024 33880 54040 33944
rect 54104 33880 54120 33944
rect 54184 33880 54200 33944
rect 54264 33880 54280 33944
rect 54344 33880 54360 33944
rect 54424 33880 54440 33944
rect 54504 33880 54520 33944
rect 54584 33880 54600 33944
rect 54664 33880 54680 33944
rect 54744 33880 54760 33944
rect 54824 33880 54840 33944
rect 54904 33880 54920 33944
rect 54984 33880 55000 33944
rect 55064 33880 55088 33944
rect 53456 33852 55088 33880
rect 33266 33774 33272 33838
rect 33336 33836 33342 33838
rect 33409 33836 33475 33839
rect 34094 33836 34100 33838
rect 33336 33834 34100 33836
rect 33336 33778 33414 33834
rect 33470 33778 34100 33834
rect 33336 33776 34100 33778
rect 33336 33774 33342 33776
rect 33409 33773 33475 33776
rect 34094 33774 34100 33776
rect 34164 33774 34170 33838
rect 26202 33670 33374 33682
rect 26202 33614 26234 33670
rect 26290 33614 26314 33670
rect 26370 33654 33374 33670
rect 26370 33614 26818 33654
rect 26202 33590 26818 33614
rect 26882 33590 27537 33654
rect 27601 33590 28256 33654
rect 28320 33590 28975 33654
rect 29039 33590 29694 33654
rect 29758 33590 30413 33654
rect 30477 33590 31132 33654
rect 31196 33590 31851 33654
rect 31915 33590 32570 33654
rect 32634 33590 33289 33654
rect 33353 33590 33374 33654
rect 26202 33574 33374 33590
rect 26202 33510 26818 33574
rect 26882 33510 27537 33574
rect 27601 33510 28256 33574
rect 28320 33510 28975 33574
rect 29039 33510 29694 33574
rect 29758 33510 30413 33574
rect 30477 33510 31132 33574
rect 31196 33510 31851 33574
rect 31915 33510 32570 33574
rect 32634 33510 33289 33574
rect 33353 33510 33374 33574
rect 26202 33494 33374 33510
rect 26202 33430 26818 33494
rect 26882 33430 27537 33494
rect 27601 33430 28256 33494
rect 28320 33430 28975 33494
rect 29039 33430 29694 33494
rect 29758 33430 30413 33494
rect 30477 33430 31132 33494
rect 31196 33430 31851 33494
rect 31915 33430 32570 33494
rect 32634 33430 33289 33494
rect 33353 33430 33374 33494
rect 26202 33414 33374 33430
rect 26202 33350 26818 33414
rect 26882 33350 27537 33414
rect 27601 33350 28256 33414
rect 28320 33350 28975 33414
rect 29039 33350 29694 33414
rect 29758 33350 30413 33414
rect 30477 33350 31132 33414
rect 31196 33350 31851 33414
rect 31915 33350 32570 33414
rect 32634 33350 33289 33414
rect 33353 33350 33374 33414
rect 26202 33334 33374 33350
rect 26202 33270 26818 33334
rect 26882 33270 27537 33334
rect 27601 33270 28256 33334
rect 28320 33270 28975 33334
rect 29039 33270 29694 33334
rect 29758 33270 30413 33334
rect 30477 33270 31132 33334
rect 31196 33270 31851 33334
rect 31915 33270 32570 33334
rect 32634 33270 33289 33334
rect 33353 33270 33374 33334
rect 26202 33254 33374 33270
rect 26202 33190 26818 33254
rect 26882 33190 27537 33254
rect 27601 33190 28256 33254
rect 28320 33190 28975 33254
rect 29039 33190 29694 33254
rect 29758 33190 30413 33254
rect 30477 33190 31132 33254
rect 31196 33190 31851 33254
rect 31915 33190 32570 33254
rect 32634 33190 33289 33254
rect 33353 33190 33374 33254
rect 26202 33174 33374 33190
rect 26202 33110 26818 33174
rect 26882 33110 27537 33174
rect 27601 33110 28256 33174
rect 28320 33110 28975 33174
rect 29039 33110 29694 33174
rect 29758 33110 30413 33174
rect 30477 33110 31132 33174
rect 31196 33110 31851 33174
rect 31915 33110 32570 33174
rect 32634 33110 33289 33174
rect 33353 33110 33374 33174
rect 26202 32954 33374 33110
rect 26202 32890 26818 32954
rect 26882 32890 27537 32954
rect 27601 32890 28256 32954
rect 28320 32890 28975 32954
rect 29039 32890 29694 32954
rect 29758 32890 30413 32954
rect 30477 32890 31132 32954
rect 31196 32890 31851 32954
rect 31915 32890 32570 32954
rect 32634 32890 33289 32954
rect 33353 32890 33374 32954
rect 26202 32874 33374 32890
rect 26202 32810 26818 32874
rect 26882 32810 27537 32874
rect 27601 32810 28256 32874
rect 28320 32810 28975 32874
rect 29039 32810 29694 32874
rect 29758 32810 30413 32874
rect 30477 32810 31132 32874
rect 31196 32810 31851 32874
rect 31915 32810 32570 32874
rect 32634 32810 33289 32874
rect 33353 32810 33374 32874
rect 26202 32794 33374 32810
rect 26202 32730 26818 32794
rect 26882 32730 27537 32794
rect 27601 32730 28256 32794
rect 28320 32730 28975 32794
rect 29039 32730 29694 32794
rect 29758 32730 30413 32794
rect 30477 32730 31132 32794
rect 31196 32730 31851 32794
rect 31915 32730 32570 32794
rect 32634 32730 33289 32794
rect 33353 32730 33374 32794
rect 26202 32714 33374 32730
rect 26202 32650 26818 32714
rect 26882 32650 27537 32714
rect 27601 32650 28256 32714
rect 28320 32650 28975 32714
rect 29039 32650 29694 32714
rect 29758 32650 30413 32714
rect 30477 32650 31132 32714
rect 31196 32650 31851 32714
rect 31915 32650 32570 32714
rect 32634 32650 33289 32714
rect 33353 32650 33374 32714
rect 26202 32634 33374 32650
rect 26202 32570 26818 32634
rect 26882 32570 27537 32634
rect 27601 32570 28256 32634
rect 28320 32570 28975 32634
rect 29039 32570 29694 32634
rect 29758 32570 30413 32634
rect 30477 32570 31132 32634
rect 31196 32570 31851 32634
rect 31915 32570 32570 32634
rect 32634 32570 33289 32634
rect 33353 32570 33374 32634
rect 26202 32554 33374 32570
rect 26202 32490 26818 32554
rect 26882 32490 27537 32554
rect 27601 32490 28256 32554
rect 28320 32490 28975 32554
rect 29039 32490 29694 32554
rect 29758 32490 30413 32554
rect 30477 32490 31132 32554
rect 31196 32490 31851 32554
rect 31915 32490 32570 32554
rect 32634 32490 33289 32554
rect 33353 32490 33374 32554
rect 26202 32474 33374 32490
rect 26202 32410 26818 32474
rect 26882 32410 27537 32474
rect 27601 32410 28256 32474
rect 28320 32410 28975 32474
rect 29039 32410 29694 32474
rect 29758 32410 30413 32474
rect 30477 32410 31132 32474
rect 31196 32410 31851 32474
rect 31915 32410 32570 32474
rect 32634 32410 33289 32474
rect 33353 32410 33374 32474
rect 26202 32382 33374 32410
rect 33650 33670 40822 33682
rect 33650 33614 33682 33670
rect 33738 33614 33762 33670
rect 33818 33654 40822 33670
rect 33818 33614 34266 33654
rect 33650 33590 34266 33614
rect 34330 33590 34985 33654
rect 35049 33590 35704 33654
rect 35768 33590 36423 33654
rect 36487 33590 37142 33654
rect 37206 33590 37861 33654
rect 37925 33590 38580 33654
rect 38644 33590 39299 33654
rect 39363 33590 40018 33654
rect 40082 33590 40737 33654
rect 40801 33590 40822 33654
rect 33650 33574 40822 33590
rect 33650 33510 34266 33574
rect 34330 33510 34985 33574
rect 35049 33510 35704 33574
rect 35768 33510 36423 33574
rect 36487 33510 37142 33574
rect 37206 33510 37861 33574
rect 37925 33510 38580 33574
rect 38644 33510 39299 33574
rect 39363 33510 40018 33574
rect 40082 33510 40737 33574
rect 40801 33510 40822 33574
rect 33650 33494 40822 33510
rect 33650 33430 34266 33494
rect 34330 33430 34985 33494
rect 35049 33430 35704 33494
rect 35768 33430 36423 33494
rect 36487 33430 37142 33494
rect 37206 33430 37861 33494
rect 37925 33430 38580 33494
rect 38644 33430 39299 33494
rect 39363 33430 40018 33494
rect 40082 33430 40737 33494
rect 40801 33430 40822 33494
rect 33650 33414 40822 33430
rect 33650 33350 34266 33414
rect 34330 33350 34985 33414
rect 35049 33350 35704 33414
rect 35768 33350 36423 33414
rect 36487 33350 37142 33414
rect 37206 33350 37861 33414
rect 37925 33350 38580 33414
rect 38644 33350 39299 33414
rect 39363 33350 40018 33414
rect 40082 33350 40737 33414
rect 40801 33350 40822 33414
rect 33650 33334 40822 33350
rect 33650 33270 34266 33334
rect 34330 33270 34985 33334
rect 35049 33270 35704 33334
rect 35768 33270 36423 33334
rect 36487 33270 37142 33334
rect 37206 33270 37861 33334
rect 37925 33270 38580 33334
rect 38644 33270 39299 33334
rect 39363 33270 40018 33334
rect 40082 33270 40737 33334
rect 40801 33270 40822 33334
rect 33650 33254 40822 33270
rect 33650 33190 34266 33254
rect 34330 33190 34985 33254
rect 35049 33190 35704 33254
rect 35768 33190 36423 33254
rect 36487 33190 37142 33254
rect 37206 33190 37861 33254
rect 37925 33190 38580 33254
rect 38644 33190 39299 33254
rect 39363 33190 40018 33254
rect 40082 33190 40737 33254
rect 40801 33190 40822 33254
rect 33650 33174 40822 33190
rect 33650 33110 34266 33174
rect 34330 33110 34985 33174
rect 35049 33110 35704 33174
rect 35768 33110 36423 33174
rect 36487 33110 37142 33174
rect 37206 33110 37861 33174
rect 37925 33110 38580 33174
rect 38644 33110 39299 33174
rect 39363 33110 40018 33174
rect 40082 33110 40737 33174
rect 40801 33110 40822 33174
rect 33650 32954 40822 33110
rect 33650 32890 34266 32954
rect 34330 32890 34985 32954
rect 35049 32890 35704 32954
rect 35768 32890 36423 32954
rect 36487 32890 37142 32954
rect 37206 32890 37861 32954
rect 37925 32890 38580 32954
rect 38644 32890 39299 32954
rect 39363 32890 40018 32954
rect 40082 32890 40737 32954
rect 40801 32890 40822 32954
rect 33650 32874 40822 32890
rect 33650 32810 34266 32874
rect 34330 32810 34985 32874
rect 35049 32810 35704 32874
rect 35768 32810 36423 32874
rect 36487 32810 37142 32874
rect 37206 32810 37861 32874
rect 37925 32810 38580 32874
rect 38644 32810 39299 32874
rect 39363 32810 40018 32874
rect 40082 32810 40737 32874
rect 40801 32810 40822 32874
rect 33650 32794 40822 32810
rect 33650 32730 34266 32794
rect 34330 32730 34985 32794
rect 35049 32730 35704 32794
rect 35768 32730 36423 32794
rect 36487 32730 37142 32794
rect 37206 32730 37861 32794
rect 37925 32730 38580 32794
rect 38644 32730 39299 32794
rect 39363 32730 40018 32794
rect 40082 32730 40737 32794
rect 40801 32730 40822 32794
rect 33650 32714 40822 32730
rect 33650 32650 34266 32714
rect 34330 32650 34985 32714
rect 35049 32650 35704 32714
rect 35768 32650 36423 32714
rect 36487 32650 37142 32714
rect 37206 32650 37861 32714
rect 37925 32650 38580 32714
rect 38644 32650 39299 32714
rect 39363 32650 40018 32714
rect 40082 32650 40737 32714
rect 40801 32650 40822 32714
rect 33650 32634 40822 32650
rect 33650 32570 34266 32634
rect 34330 32570 34985 32634
rect 35049 32570 35704 32634
rect 35768 32570 36423 32634
rect 36487 32570 37142 32634
rect 37206 32570 37861 32634
rect 37925 32570 38580 32634
rect 38644 32570 39299 32634
rect 39363 32570 40018 32634
rect 40082 32570 40737 32634
rect 40801 32570 40822 32634
rect 33650 32554 40822 32570
rect 33650 32490 34266 32554
rect 34330 32490 34985 32554
rect 35049 32490 35704 32554
rect 35768 32490 36423 32554
rect 36487 32490 37142 32554
rect 37206 32490 37861 32554
rect 37925 32490 38580 32554
rect 38644 32490 39299 32554
rect 39363 32490 40018 32554
rect 40082 32490 40737 32554
rect 40801 32490 40822 32554
rect 33650 32474 40822 32490
rect 33650 32410 34266 32474
rect 34330 32410 34985 32474
rect 35049 32410 35704 32474
rect 35768 32410 36423 32474
rect 36487 32410 37142 32474
rect 37206 32410 37861 32474
rect 37925 32410 38580 32474
rect 38644 32410 39299 32474
rect 39363 32410 40018 32474
rect 40082 32410 40737 32474
rect 40801 32410 40822 32474
rect 33650 32382 40822 32410
rect 26204 32254 26404 32282
rect 26204 32190 26232 32254
rect 26296 32250 26312 32254
rect 26296 32190 26312 32194
rect 26376 32190 26404 32254
rect 26204 32162 26404 32190
rect 33652 32254 33852 32282
rect 33652 32190 33680 32254
rect 33744 32250 33760 32254
rect 33744 32190 33760 32194
rect 33824 32190 33852 32254
rect 33652 32162 33852 32190
rect 900 32064 2532 32092
rect 900 32000 924 32064
rect 988 32000 1004 32064
rect 1068 32000 1084 32064
rect 1148 32000 1164 32064
rect 1228 32000 1244 32064
rect 1308 32000 1324 32064
rect 1388 32000 1404 32064
rect 1468 32000 1484 32064
rect 1548 32000 1564 32064
rect 1628 32000 1644 32064
rect 1708 32000 1724 32064
rect 1788 32000 1804 32064
rect 1868 32000 1884 32064
rect 1948 32000 1964 32064
rect 2028 32000 2044 32064
rect 2108 32000 2124 32064
rect 2188 32000 2204 32064
rect 2268 32000 2284 32064
rect 2348 32000 2364 32064
rect 2428 32000 2444 32064
rect 2508 32000 2532 32064
rect 900 31972 2532 32000
rect 55904 32064 57536 32092
rect 55904 32000 55928 32064
rect 55992 32000 56008 32064
rect 56072 32000 56088 32064
rect 56152 32000 56168 32064
rect 56232 32000 56248 32064
rect 56312 32000 56328 32064
rect 56392 32000 56408 32064
rect 56472 32000 56488 32064
rect 56552 32000 56568 32064
rect 56632 32000 56648 32064
rect 56712 32000 56728 32064
rect 56792 32000 56808 32064
rect 56872 32000 56888 32064
rect 56952 32000 56968 32064
rect 57032 32000 57048 32064
rect 57112 32000 57128 32064
rect 57192 32000 57208 32064
rect 57272 32000 57288 32064
rect 57352 32000 57368 32064
rect 57432 32000 57448 32064
rect 57512 32000 57536 32064
rect 55904 31972 57536 32000
rect 3348 30184 4980 30212
rect 3348 30120 3372 30184
rect 3436 30120 3452 30184
rect 3516 30120 3532 30184
rect 3596 30120 3612 30184
rect 3676 30120 3692 30184
rect 3756 30120 3772 30184
rect 3836 30120 3852 30184
rect 3916 30120 3932 30184
rect 3996 30120 4012 30184
rect 4076 30120 4092 30184
rect 4156 30120 4172 30184
rect 4236 30120 4252 30184
rect 4316 30120 4332 30184
rect 4396 30120 4412 30184
rect 4476 30120 4492 30184
rect 4556 30120 4572 30184
rect 4636 30120 4652 30184
rect 4716 30120 4732 30184
rect 4796 30120 4812 30184
rect 4876 30120 4892 30184
rect 4956 30120 4980 30184
rect 53456 30184 55088 30212
rect 33409 30178 33475 30179
rect 33404 30176 33410 30178
rect 3348 30092 4980 30120
rect 33320 30116 33410 30176
rect 33404 30114 33410 30116
rect 33474 30114 33480 30178
rect 53456 30120 53480 30184
rect 53544 30120 53560 30184
rect 53624 30120 53640 30184
rect 53704 30120 53720 30184
rect 53784 30120 53800 30184
rect 53864 30120 53880 30184
rect 53944 30120 53960 30184
rect 54024 30120 54040 30184
rect 54104 30120 54120 30184
rect 54184 30120 54200 30184
rect 54264 30120 54280 30184
rect 54344 30120 54360 30184
rect 54424 30120 54440 30184
rect 54504 30120 54520 30184
rect 54584 30120 54600 30184
rect 54664 30120 54680 30184
rect 54744 30120 54760 30184
rect 54824 30120 54840 30184
rect 54904 30120 54920 30184
rect 54984 30120 55000 30184
rect 55064 30120 55088 30184
rect 33409 30113 33475 30114
rect 53456 30092 55088 30120
rect 29926 29910 37098 29922
rect 29926 29854 29958 29910
rect 30014 29854 30038 29910
rect 30094 29894 37098 29910
rect 30094 29854 30542 29894
rect 29926 29830 30542 29854
rect 30606 29830 31261 29894
rect 31325 29830 31980 29894
rect 32044 29830 32699 29894
rect 32763 29830 33418 29894
rect 33482 29830 34137 29894
rect 34201 29830 34856 29894
rect 34920 29830 35575 29894
rect 35639 29830 36294 29894
rect 36358 29830 37013 29894
rect 37077 29830 37098 29894
rect 29926 29814 37098 29830
rect 29926 29750 30542 29814
rect 30606 29750 31261 29814
rect 31325 29750 31980 29814
rect 32044 29750 32699 29814
rect 32763 29750 33418 29814
rect 33482 29750 34137 29814
rect 34201 29750 34856 29814
rect 34920 29750 35575 29814
rect 35639 29750 36294 29814
rect 36358 29750 37013 29814
rect 37077 29750 37098 29814
rect 29926 29734 37098 29750
rect 29926 29670 30542 29734
rect 30606 29670 31261 29734
rect 31325 29670 31980 29734
rect 32044 29670 32699 29734
rect 32763 29670 33418 29734
rect 33482 29670 34137 29734
rect 34201 29670 34856 29734
rect 34920 29670 35575 29734
rect 35639 29670 36294 29734
rect 36358 29670 37013 29734
rect 37077 29670 37098 29734
rect 29926 29654 37098 29670
rect 29926 29590 30542 29654
rect 30606 29590 31261 29654
rect 31325 29590 31980 29654
rect 32044 29590 32699 29654
rect 32763 29590 33418 29654
rect 33482 29590 34137 29654
rect 34201 29590 34856 29654
rect 34920 29590 35575 29654
rect 35639 29590 36294 29654
rect 36358 29590 37013 29654
rect 37077 29590 37098 29654
rect 29926 29574 37098 29590
rect 29926 29510 30542 29574
rect 30606 29510 31261 29574
rect 31325 29510 31980 29574
rect 32044 29510 32699 29574
rect 32763 29510 33418 29574
rect 33482 29510 34137 29574
rect 34201 29510 34856 29574
rect 34920 29510 35575 29574
rect 35639 29510 36294 29574
rect 36358 29510 37013 29574
rect 37077 29510 37098 29574
rect 29926 29494 37098 29510
rect 29926 29430 30542 29494
rect 30606 29430 31261 29494
rect 31325 29430 31980 29494
rect 32044 29430 32699 29494
rect 32763 29430 33418 29494
rect 33482 29430 34137 29494
rect 34201 29430 34856 29494
rect 34920 29430 35575 29494
rect 35639 29430 36294 29494
rect 36358 29430 37013 29494
rect 37077 29430 37098 29494
rect 29926 29414 37098 29430
rect 29926 29350 30542 29414
rect 30606 29350 31261 29414
rect 31325 29350 31980 29414
rect 32044 29350 32699 29414
rect 32763 29350 33418 29414
rect 33482 29350 34137 29414
rect 34201 29350 34856 29414
rect 34920 29350 35575 29414
rect 35639 29350 36294 29414
rect 36358 29350 37013 29414
rect 37077 29350 37098 29414
rect 29926 29194 37098 29350
rect 29926 29130 30542 29194
rect 30606 29130 31261 29194
rect 31325 29130 31980 29194
rect 32044 29130 32699 29194
rect 32763 29130 33418 29194
rect 33482 29130 34137 29194
rect 34201 29130 34856 29194
rect 34920 29130 35575 29194
rect 35639 29130 36294 29194
rect 36358 29130 37013 29194
rect 37077 29130 37098 29194
rect 29926 29114 37098 29130
rect 29926 29050 30542 29114
rect 30606 29050 31261 29114
rect 31325 29050 31980 29114
rect 32044 29050 32699 29114
rect 32763 29050 33418 29114
rect 33482 29050 34137 29114
rect 34201 29050 34856 29114
rect 34920 29050 35575 29114
rect 35639 29050 36294 29114
rect 36358 29050 37013 29114
rect 37077 29050 37098 29114
rect 29926 29034 37098 29050
rect 29926 28970 30542 29034
rect 30606 28970 31261 29034
rect 31325 28970 31980 29034
rect 32044 28970 32699 29034
rect 32763 28970 33418 29034
rect 33482 28970 34137 29034
rect 34201 28970 34856 29034
rect 34920 28970 35575 29034
rect 35639 28970 36294 29034
rect 36358 28970 37013 29034
rect 37077 28970 37098 29034
rect 29926 28954 37098 28970
rect 29926 28890 30542 28954
rect 30606 28890 31261 28954
rect 31325 28890 31980 28954
rect 32044 28890 32699 28954
rect 32763 28890 33418 28954
rect 33482 28890 34137 28954
rect 34201 28890 34856 28954
rect 34920 28890 35575 28954
rect 35639 28890 36294 28954
rect 36358 28890 37013 28954
rect 37077 28890 37098 28954
rect 29926 28874 37098 28890
rect 29926 28810 30542 28874
rect 30606 28810 31261 28874
rect 31325 28810 31980 28874
rect 32044 28810 32699 28874
rect 32763 28810 33418 28874
rect 33482 28810 34137 28874
rect 34201 28810 34856 28874
rect 34920 28810 35575 28874
rect 35639 28810 36294 28874
rect 36358 28810 37013 28874
rect 37077 28810 37098 28874
rect 29926 28794 37098 28810
rect 29926 28730 30542 28794
rect 30606 28730 31261 28794
rect 31325 28730 31980 28794
rect 32044 28730 32699 28794
rect 32763 28730 33418 28794
rect 33482 28730 34137 28794
rect 34201 28730 34856 28794
rect 34920 28730 35575 28794
rect 35639 28730 36294 28794
rect 36358 28730 37013 28794
rect 37077 28730 37098 28794
rect 29926 28714 37098 28730
rect 29926 28650 30542 28714
rect 30606 28650 31261 28714
rect 31325 28650 31980 28714
rect 32044 28650 32699 28714
rect 32763 28650 33418 28714
rect 33482 28650 34137 28714
rect 34201 28650 34856 28714
rect 34920 28650 35575 28714
rect 35639 28650 36294 28714
rect 36358 28650 37013 28714
rect 37077 28650 37098 28714
rect 29926 28622 37098 28650
rect 29928 28494 30128 28522
rect 29928 28430 29956 28494
rect 30020 28490 30036 28494
rect 30020 28430 30036 28434
rect 30100 28430 30128 28494
rect 29928 28402 30128 28430
rect 900 28304 2532 28332
rect 900 28240 924 28304
rect 988 28240 1004 28304
rect 1068 28240 1084 28304
rect 1148 28240 1164 28304
rect 1228 28240 1244 28304
rect 1308 28240 1324 28304
rect 1388 28240 1404 28304
rect 1468 28240 1484 28304
rect 1548 28240 1564 28304
rect 1628 28240 1644 28304
rect 1708 28240 1724 28304
rect 1788 28240 1804 28304
rect 1868 28240 1884 28304
rect 1948 28240 1964 28304
rect 2028 28240 2044 28304
rect 2108 28240 2124 28304
rect 2188 28240 2204 28304
rect 2268 28240 2284 28304
rect 2348 28240 2364 28304
rect 2428 28240 2444 28304
rect 2508 28240 2532 28304
rect 900 28212 2532 28240
rect 55904 28304 57536 28332
rect 55904 28240 55928 28304
rect 55992 28240 56008 28304
rect 56072 28240 56088 28304
rect 56152 28240 56168 28304
rect 56232 28240 56248 28304
rect 56312 28240 56328 28304
rect 56392 28240 56408 28304
rect 56472 28240 56488 28304
rect 56552 28240 56568 28304
rect 56632 28240 56648 28304
rect 56712 28240 56728 28304
rect 56792 28240 56808 28304
rect 56872 28240 56888 28304
rect 56952 28240 56968 28304
rect 57032 28240 57048 28304
rect 57112 28240 57128 28304
rect 57192 28240 57208 28304
rect 57272 28240 57288 28304
rect 57352 28240 57368 28304
rect 57432 28240 57448 28304
rect 57512 28240 57536 28304
rect 55904 28212 57536 28240
rect 3348 26424 4980 26452
rect 3348 26360 3372 26424
rect 3436 26360 3452 26424
rect 3516 26360 3532 26424
rect 3596 26360 3612 26424
rect 3676 26360 3692 26424
rect 3756 26360 3772 26424
rect 3836 26360 3852 26424
rect 3916 26360 3932 26424
rect 3996 26360 4012 26424
rect 4076 26360 4092 26424
rect 4156 26360 4172 26424
rect 4236 26360 4252 26424
rect 4316 26360 4332 26424
rect 4396 26360 4412 26424
rect 4476 26360 4492 26424
rect 4556 26360 4572 26424
rect 4636 26360 4652 26424
rect 4716 26360 4732 26424
rect 4796 26360 4812 26424
rect 4876 26360 4892 26424
rect 4956 26360 4980 26424
rect 53456 26424 55088 26452
rect 33409 26396 33475 26397
rect 33404 26394 33410 26396
rect 3348 26332 4980 26360
rect 33320 26334 33410 26394
rect 33404 26332 33410 26334
rect 33474 26332 33480 26396
rect 53456 26360 53480 26424
rect 53544 26360 53560 26424
rect 53624 26360 53640 26424
rect 53704 26360 53720 26424
rect 53784 26360 53800 26424
rect 53864 26360 53880 26424
rect 53944 26360 53960 26424
rect 54024 26360 54040 26424
rect 54104 26360 54120 26424
rect 54184 26360 54200 26424
rect 54264 26360 54280 26424
rect 54344 26360 54360 26424
rect 54424 26360 54440 26424
rect 54504 26360 54520 26424
rect 54584 26360 54600 26424
rect 54664 26360 54680 26424
rect 54744 26360 54760 26424
rect 54824 26360 54840 26424
rect 54904 26360 54920 26424
rect 54984 26360 55000 26424
rect 55064 26360 55088 26424
rect 53456 26332 55088 26360
rect 33409 26331 33475 26332
rect 29926 26150 37098 26162
rect 29926 26094 29958 26150
rect 30014 26094 30038 26150
rect 30094 26134 37098 26150
rect 30094 26094 30542 26134
rect 29926 26070 30542 26094
rect 30606 26070 31261 26134
rect 31325 26070 31980 26134
rect 32044 26070 32699 26134
rect 32763 26070 33418 26134
rect 33482 26070 34137 26134
rect 34201 26070 34856 26134
rect 34920 26070 35575 26134
rect 35639 26070 36294 26134
rect 36358 26070 37013 26134
rect 37077 26070 37098 26134
rect 29926 26054 37098 26070
rect 29926 25990 30542 26054
rect 30606 25990 31261 26054
rect 31325 25990 31980 26054
rect 32044 25990 32699 26054
rect 32763 25990 33418 26054
rect 33482 25990 34137 26054
rect 34201 25990 34856 26054
rect 34920 25990 35575 26054
rect 35639 25990 36294 26054
rect 36358 25990 37013 26054
rect 37077 25990 37098 26054
rect 29926 25974 37098 25990
rect 29926 25910 30542 25974
rect 30606 25910 31261 25974
rect 31325 25910 31980 25974
rect 32044 25910 32699 25974
rect 32763 25910 33418 25974
rect 33482 25910 34137 25974
rect 34201 25910 34856 25974
rect 34920 25910 35575 25974
rect 35639 25910 36294 25974
rect 36358 25910 37013 25974
rect 37077 25910 37098 25974
rect 29926 25894 37098 25910
rect 29926 25830 30542 25894
rect 30606 25830 31261 25894
rect 31325 25830 31980 25894
rect 32044 25830 32699 25894
rect 32763 25830 33418 25894
rect 33482 25830 34137 25894
rect 34201 25830 34856 25894
rect 34920 25830 35575 25894
rect 35639 25830 36294 25894
rect 36358 25830 37013 25894
rect 37077 25830 37098 25894
rect 29926 25814 37098 25830
rect 29453 25784 29519 25787
rect 29678 25784 29684 25786
rect 29453 25782 29684 25784
rect 29453 25726 29458 25782
rect 29514 25726 29684 25782
rect 29453 25724 29684 25726
rect 29453 25721 29519 25724
rect 29678 25722 29684 25724
rect 29748 25722 29754 25786
rect 29926 25750 30542 25814
rect 30606 25750 31261 25814
rect 31325 25750 31980 25814
rect 32044 25750 32699 25814
rect 32763 25750 33418 25814
rect 33482 25750 34137 25814
rect 34201 25750 34856 25814
rect 34920 25750 35575 25814
rect 35639 25750 36294 25814
rect 36358 25750 37013 25814
rect 37077 25750 37098 25814
rect 29926 25734 37098 25750
rect 29926 25670 30542 25734
rect 30606 25670 31261 25734
rect 31325 25670 31980 25734
rect 32044 25670 32699 25734
rect 32763 25670 33418 25734
rect 33482 25670 34137 25734
rect 34201 25670 34856 25734
rect 34920 25670 35575 25734
rect 35639 25670 36294 25734
rect 36358 25670 37013 25734
rect 37077 25670 37098 25734
rect 29926 25654 37098 25670
rect 29926 25590 30542 25654
rect 30606 25590 31261 25654
rect 31325 25590 31980 25654
rect 32044 25590 32699 25654
rect 32763 25590 33418 25654
rect 33482 25590 34137 25654
rect 34201 25590 34856 25654
rect 34920 25590 35575 25654
rect 35639 25590 36294 25654
rect 36358 25590 37013 25654
rect 37077 25590 37098 25654
rect 29926 25434 37098 25590
rect 29926 25370 30542 25434
rect 30606 25370 31261 25434
rect 31325 25370 31980 25434
rect 32044 25370 32699 25434
rect 32763 25370 33418 25434
rect 33482 25370 34137 25434
rect 34201 25370 34856 25434
rect 34920 25370 35575 25434
rect 35639 25370 36294 25434
rect 36358 25370 37013 25434
rect 37077 25370 37098 25434
rect 29926 25354 37098 25370
rect 29926 25290 30542 25354
rect 30606 25290 31261 25354
rect 31325 25290 31980 25354
rect 32044 25290 32699 25354
rect 32763 25290 33418 25354
rect 33482 25290 34137 25354
rect 34201 25290 34856 25354
rect 34920 25290 35575 25354
rect 35639 25290 36294 25354
rect 36358 25290 37013 25354
rect 37077 25290 37098 25354
rect 29926 25274 37098 25290
rect 29926 25210 30542 25274
rect 30606 25210 31261 25274
rect 31325 25210 31980 25274
rect 32044 25210 32699 25274
rect 32763 25210 33418 25274
rect 33482 25210 34137 25274
rect 34201 25210 34856 25274
rect 34920 25210 35575 25274
rect 35639 25210 36294 25274
rect 36358 25210 37013 25274
rect 37077 25210 37098 25274
rect 29926 25194 37098 25210
rect 29926 25130 30542 25194
rect 30606 25130 31261 25194
rect 31325 25130 31980 25194
rect 32044 25130 32699 25194
rect 32763 25130 33418 25194
rect 33482 25130 34137 25194
rect 34201 25130 34856 25194
rect 34920 25130 35575 25194
rect 35639 25130 36294 25194
rect 36358 25130 37013 25194
rect 37077 25130 37098 25194
rect 29926 25114 37098 25130
rect 29926 25050 30542 25114
rect 30606 25050 31261 25114
rect 31325 25050 31980 25114
rect 32044 25050 32699 25114
rect 32763 25050 33418 25114
rect 33482 25050 34137 25114
rect 34201 25050 34856 25114
rect 34920 25050 35575 25114
rect 35639 25050 36294 25114
rect 36358 25050 37013 25114
rect 37077 25050 37098 25114
rect 29926 25034 37098 25050
rect 29926 24970 30542 25034
rect 30606 24970 31261 25034
rect 31325 24970 31980 25034
rect 32044 24970 32699 25034
rect 32763 24970 33418 25034
rect 33482 24970 34137 25034
rect 34201 24970 34856 25034
rect 34920 24970 35575 25034
rect 35639 24970 36294 25034
rect 36358 24970 37013 25034
rect 37077 24970 37098 25034
rect 29926 24954 37098 24970
rect 29926 24890 30542 24954
rect 30606 24890 31261 24954
rect 31325 24890 31980 24954
rect 32044 24890 32699 24954
rect 32763 24890 33418 24954
rect 33482 24890 34137 24954
rect 34201 24890 34856 24954
rect 34920 24890 35575 24954
rect 35639 24890 36294 24954
rect 36358 24890 37013 24954
rect 37077 24890 37098 24954
rect 29926 24862 37098 24890
rect 29928 24734 30128 24762
rect 29928 24670 29956 24734
rect 30020 24730 30036 24734
rect 30020 24670 30036 24674
rect 30100 24670 30128 24734
rect 29928 24642 30128 24670
rect 900 24544 2532 24572
rect 900 24480 924 24544
rect 988 24480 1004 24544
rect 1068 24480 1084 24544
rect 1148 24480 1164 24544
rect 1228 24480 1244 24544
rect 1308 24480 1324 24544
rect 1388 24480 1404 24544
rect 1468 24480 1484 24544
rect 1548 24480 1564 24544
rect 1628 24480 1644 24544
rect 1708 24480 1724 24544
rect 1788 24480 1804 24544
rect 1868 24480 1884 24544
rect 1948 24480 1964 24544
rect 2028 24480 2044 24544
rect 2108 24480 2124 24544
rect 2188 24480 2204 24544
rect 2268 24480 2284 24544
rect 2348 24480 2364 24544
rect 2428 24480 2444 24544
rect 2508 24480 2532 24544
rect 900 24452 2532 24480
rect 55904 24544 57536 24572
rect 55904 24480 55928 24544
rect 55992 24480 56008 24544
rect 56072 24480 56088 24544
rect 56152 24480 56168 24544
rect 56232 24480 56248 24544
rect 56312 24480 56328 24544
rect 56392 24480 56408 24544
rect 56472 24480 56488 24544
rect 56552 24480 56568 24544
rect 56632 24480 56648 24544
rect 56712 24480 56728 24544
rect 56792 24480 56808 24544
rect 56872 24480 56888 24544
rect 56952 24480 56968 24544
rect 57032 24480 57048 24544
rect 57112 24480 57128 24544
rect 57192 24480 57208 24544
rect 57272 24480 57288 24544
rect 57352 24480 57368 24544
rect 57432 24480 57448 24544
rect 57512 24480 57536 24544
rect 55904 24452 57536 24480
rect 3348 22664 4980 22692
rect 3348 22600 3372 22664
rect 3436 22600 3452 22664
rect 3516 22600 3532 22664
rect 3596 22600 3612 22664
rect 3676 22600 3692 22664
rect 3756 22600 3772 22664
rect 3836 22600 3852 22664
rect 3916 22600 3932 22664
rect 3996 22600 4012 22664
rect 4076 22600 4092 22664
rect 4156 22600 4172 22664
rect 4236 22600 4252 22664
rect 4316 22600 4332 22664
rect 4396 22600 4412 22664
rect 4476 22600 4492 22664
rect 4556 22600 4572 22664
rect 4636 22600 4652 22664
rect 4716 22600 4732 22664
rect 4796 22600 4812 22664
rect 4876 22600 4892 22664
rect 4956 22600 4980 22664
rect 3348 22572 4980 22600
rect 53456 22664 55088 22692
rect 53456 22600 53480 22664
rect 53544 22600 53560 22664
rect 53624 22600 53640 22664
rect 53704 22600 53720 22664
rect 53784 22600 53800 22664
rect 53864 22600 53880 22664
rect 53944 22600 53960 22664
rect 54024 22600 54040 22664
rect 54104 22600 54120 22664
rect 54184 22600 54200 22664
rect 54264 22600 54280 22664
rect 54344 22600 54360 22664
rect 54424 22600 54440 22664
rect 54504 22600 54520 22664
rect 54584 22600 54600 22664
rect 54664 22600 54680 22664
rect 54744 22600 54760 22664
rect 54824 22600 54840 22664
rect 54904 22600 54920 22664
rect 54984 22600 55000 22664
rect 55064 22600 55088 22664
rect 53456 22572 55088 22600
rect 900 20784 2532 20812
rect 900 20720 924 20784
rect 988 20720 1004 20784
rect 1068 20720 1084 20784
rect 1148 20720 1164 20784
rect 1228 20720 1244 20784
rect 1308 20720 1324 20784
rect 1388 20720 1404 20784
rect 1468 20720 1484 20784
rect 1548 20720 1564 20784
rect 1628 20720 1644 20784
rect 1708 20720 1724 20784
rect 1788 20720 1804 20784
rect 1868 20720 1884 20784
rect 1948 20720 1964 20784
rect 2028 20720 2044 20784
rect 2108 20720 2124 20784
rect 2188 20720 2204 20784
rect 2268 20720 2284 20784
rect 2348 20720 2364 20784
rect 2428 20720 2444 20784
rect 2508 20720 2532 20784
rect 900 20692 2532 20720
rect 55904 20784 57536 20812
rect 55904 20720 55928 20784
rect 55992 20720 56008 20784
rect 56072 20720 56088 20784
rect 56152 20720 56168 20784
rect 56232 20720 56248 20784
rect 56312 20720 56328 20784
rect 56392 20720 56408 20784
rect 56472 20720 56488 20784
rect 56552 20720 56568 20784
rect 56632 20720 56648 20784
rect 56712 20720 56728 20784
rect 56792 20720 56808 20784
rect 56872 20720 56888 20784
rect 56952 20720 56968 20784
rect 57032 20720 57048 20784
rect 57112 20720 57128 20784
rect 57192 20720 57208 20784
rect 57272 20720 57288 20784
rect 57352 20720 57368 20784
rect 57432 20720 57448 20784
rect 57512 20720 57536 20784
rect 55904 20692 57536 20720
rect 3348 18904 4980 18932
rect 3348 18840 3372 18904
rect 3436 18840 3452 18904
rect 3516 18840 3532 18904
rect 3596 18840 3612 18904
rect 3676 18840 3692 18904
rect 3756 18840 3772 18904
rect 3836 18840 3852 18904
rect 3916 18840 3932 18904
rect 3996 18840 4012 18904
rect 4076 18840 4092 18904
rect 4156 18840 4172 18904
rect 4236 18840 4252 18904
rect 4316 18840 4332 18904
rect 4396 18840 4412 18904
rect 4476 18840 4492 18904
rect 4556 18840 4572 18904
rect 4636 18840 4652 18904
rect 4716 18840 4732 18904
rect 4796 18840 4812 18904
rect 4876 18840 4892 18904
rect 4956 18840 4980 18904
rect 3348 18812 4980 18840
rect 53456 18904 55088 18932
rect 53456 18840 53480 18904
rect 53544 18840 53560 18904
rect 53624 18840 53640 18904
rect 53704 18840 53720 18904
rect 53784 18840 53800 18904
rect 53864 18840 53880 18904
rect 53944 18840 53960 18904
rect 54024 18840 54040 18904
rect 54104 18840 54120 18904
rect 54184 18840 54200 18904
rect 54264 18840 54280 18904
rect 54344 18840 54360 18904
rect 54424 18840 54440 18904
rect 54504 18840 54520 18904
rect 54584 18840 54600 18904
rect 54664 18840 54680 18904
rect 54744 18840 54760 18904
rect 54824 18840 54840 18904
rect 54904 18840 54920 18904
rect 54984 18840 55000 18904
rect 55064 18840 55088 18904
rect 53456 18812 55088 18840
rect 900 17024 2532 17052
rect 900 16960 924 17024
rect 988 16960 1004 17024
rect 1068 16960 1084 17024
rect 1148 16960 1164 17024
rect 1228 16960 1244 17024
rect 1308 16960 1324 17024
rect 1388 16960 1404 17024
rect 1468 16960 1484 17024
rect 1548 16960 1564 17024
rect 1628 16960 1644 17024
rect 1708 16960 1724 17024
rect 1788 16960 1804 17024
rect 1868 16960 1884 17024
rect 1948 16960 1964 17024
rect 2028 16960 2044 17024
rect 2108 16960 2124 17024
rect 2188 16960 2204 17024
rect 2268 16960 2284 17024
rect 2348 16960 2364 17024
rect 2428 16960 2444 17024
rect 2508 16960 2532 17024
rect 900 16932 2532 16960
rect 55904 17024 57536 17052
rect 55904 16960 55928 17024
rect 55992 16960 56008 17024
rect 56072 16960 56088 17024
rect 56152 16960 56168 17024
rect 56232 16960 56248 17024
rect 56312 16960 56328 17024
rect 56392 16960 56408 17024
rect 56472 16960 56488 17024
rect 56552 16960 56568 17024
rect 56632 16960 56648 17024
rect 56712 16960 56728 17024
rect 56792 16960 56808 17024
rect 56872 16960 56888 17024
rect 56952 16960 56968 17024
rect 57032 16960 57048 17024
rect 57112 16960 57128 17024
rect 57192 16960 57208 17024
rect 57272 16960 57288 17024
rect 57352 16960 57368 17024
rect 57432 16960 57448 17024
rect 57512 16960 57536 17024
rect 55904 16932 57536 16960
rect 3348 15144 4980 15172
rect 3348 15080 3372 15144
rect 3436 15080 3452 15144
rect 3516 15080 3532 15144
rect 3596 15080 3612 15144
rect 3676 15080 3692 15144
rect 3756 15080 3772 15144
rect 3836 15080 3852 15144
rect 3916 15080 3932 15144
rect 3996 15080 4012 15144
rect 4076 15080 4092 15144
rect 4156 15080 4172 15144
rect 4236 15080 4252 15144
rect 4316 15080 4332 15144
rect 4396 15080 4412 15144
rect 4476 15080 4492 15144
rect 4556 15080 4572 15144
rect 4636 15080 4652 15144
rect 4716 15080 4732 15144
rect 4796 15080 4812 15144
rect 4876 15080 4892 15144
rect 4956 15080 4980 15144
rect 3348 15052 4980 15080
rect 53456 15144 55088 15172
rect 53456 15080 53480 15144
rect 53544 15080 53560 15144
rect 53624 15080 53640 15144
rect 53704 15080 53720 15144
rect 53784 15080 53800 15144
rect 53864 15080 53880 15144
rect 53944 15080 53960 15144
rect 54024 15080 54040 15144
rect 54104 15080 54120 15144
rect 54184 15080 54200 15144
rect 54264 15080 54280 15144
rect 54344 15080 54360 15144
rect 54424 15080 54440 15144
rect 54504 15080 54520 15144
rect 54584 15080 54600 15144
rect 54664 15080 54680 15144
rect 54744 15080 54760 15144
rect 54824 15080 54840 15144
rect 54904 15080 54920 15144
rect 54984 15080 55000 15144
rect 55064 15080 55088 15144
rect 53456 15052 55088 15080
rect 900 13264 2532 13292
rect 900 13200 924 13264
rect 988 13200 1004 13264
rect 1068 13200 1084 13264
rect 1148 13200 1164 13264
rect 1228 13200 1244 13264
rect 1308 13200 1324 13264
rect 1388 13200 1404 13264
rect 1468 13200 1484 13264
rect 1548 13200 1564 13264
rect 1628 13200 1644 13264
rect 1708 13200 1724 13264
rect 1788 13200 1804 13264
rect 1868 13200 1884 13264
rect 1948 13200 1964 13264
rect 2028 13200 2044 13264
rect 2108 13200 2124 13264
rect 2188 13200 2204 13264
rect 2268 13200 2284 13264
rect 2348 13200 2364 13264
rect 2428 13200 2444 13264
rect 2508 13200 2532 13264
rect 900 13172 2532 13200
rect 55904 13264 57536 13292
rect 55904 13200 55928 13264
rect 55992 13200 56008 13264
rect 56072 13200 56088 13264
rect 56152 13200 56168 13264
rect 56232 13200 56248 13264
rect 56312 13200 56328 13264
rect 56392 13200 56408 13264
rect 56472 13200 56488 13264
rect 56552 13200 56568 13264
rect 56632 13200 56648 13264
rect 56712 13200 56728 13264
rect 56792 13200 56808 13264
rect 56872 13200 56888 13264
rect 56952 13200 56968 13264
rect 57032 13200 57048 13264
rect 57112 13200 57128 13264
rect 57192 13200 57208 13264
rect 57272 13200 57288 13264
rect 57352 13200 57368 13264
rect 57432 13200 57448 13264
rect 57512 13200 57536 13264
rect 55904 13172 57536 13200
rect 3348 11384 4980 11412
rect 3348 11320 3372 11384
rect 3436 11320 3452 11384
rect 3516 11320 3532 11384
rect 3596 11320 3612 11384
rect 3676 11320 3692 11384
rect 3756 11320 3772 11384
rect 3836 11320 3852 11384
rect 3916 11320 3932 11384
rect 3996 11320 4012 11384
rect 4076 11320 4092 11384
rect 4156 11320 4172 11384
rect 4236 11320 4252 11384
rect 4316 11320 4332 11384
rect 4396 11320 4412 11384
rect 4476 11320 4492 11384
rect 4556 11320 4572 11384
rect 4636 11320 4652 11384
rect 4716 11320 4732 11384
rect 4796 11320 4812 11384
rect 4876 11320 4892 11384
rect 4956 11320 4980 11384
rect 3348 11292 4980 11320
rect 53456 11384 55088 11412
rect 53456 11320 53480 11384
rect 53544 11320 53560 11384
rect 53624 11320 53640 11384
rect 53704 11320 53720 11384
rect 53784 11320 53800 11384
rect 53864 11320 53880 11384
rect 53944 11320 53960 11384
rect 54024 11320 54040 11384
rect 54104 11320 54120 11384
rect 54184 11320 54200 11384
rect 54264 11320 54280 11384
rect 54344 11320 54360 11384
rect 54424 11320 54440 11384
rect 54504 11320 54520 11384
rect 54584 11320 54600 11384
rect 54664 11320 54680 11384
rect 54744 11320 54760 11384
rect 54824 11320 54840 11384
rect 54904 11320 54920 11384
rect 54984 11320 55000 11384
rect 55064 11320 55088 11384
rect 53456 11292 55088 11320
rect 900 9504 2532 9532
rect 900 9440 924 9504
rect 988 9440 1004 9504
rect 1068 9440 1084 9504
rect 1148 9440 1164 9504
rect 1228 9440 1244 9504
rect 1308 9440 1324 9504
rect 1388 9440 1404 9504
rect 1468 9440 1484 9504
rect 1548 9440 1564 9504
rect 1628 9440 1644 9504
rect 1708 9440 1724 9504
rect 1788 9440 1804 9504
rect 1868 9440 1884 9504
rect 1948 9440 1964 9504
rect 2028 9440 2044 9504
rect 2108 9440 2124 9504
rect 2188 9440 2204 9504
rect 2268 9440 2284 9504
rect 2348 9440 2364 9504
rect 2428 9440 2444 9504
rect 2508 9440 2532 9504
rect 900 9412 2532 9440
rect 55904 9504 57536 9532
rect 55904 9440 55928 9504
rect 55992 9440 56008 9504
rect 56072 9440 56088 9504
rect 56152 9440 56168 9504
rect 56232 9440 56248 9504
rect 56312 9440 56328 9504
rect 56392 9440 56408 9504
rect 56472 9440 56488 9504
rect 56552 9440 56568 9504
rect 56632 9440 56648 9504
rect 56712 9440 56728 9504
rect 56792 9440 56808 9504
rect 56872 9440 56888 9504
rect 56952 9440 56968 9504
rect 57032 9440 57048 9504
rect 57112 9440 57128 9504
rect 57192 9440 57208 9504
rect 57272 9440 57288 9504
rect 57352 9440 57368 9504
rect 57432 9440 57448 9504
rect 57512 9440 57536 9504
rect 55904 9412 57536 9440
rect 3348 7624 4980 7652
rect 3348 7560 3372 7624
rect 3436 7560 3452 7624
rect 3516 7560 3532 7624
rect 3596 7560 3612 7624
rect 3676 7560 3692 7624
rect 3756 7560 3772 7624
rect 3836 7560 3852 7624
rect 3916 7560 3932 7624
rect 3996 7560 4012 7624
rect 4076 7560 4092 7624
rect 4156 7560 4172 7624
rect 4236 7560 4252 7624
rect 4316 7560 4332 7624
rect 4396 7560 4412 7624
rect 4476 7560 4492 7624
rect 4556 7560 4572 7624
rect 4636 7560 4652 7624
rect 4716 7560 4732 7624
rect 4796 7560 4812 7624
rect 4876 7560 4892 7624
rect 4956 7560 4980 7624
rect 3348 7532 4980 7560
rect 53456 7624 55088 7652
rect 53456 7560 53480 7624
rect 53544 7560 53560 7624
rect 53624 7560 53640 7624
rect 53704 7560 53720 7624
rect 53784 7560 53800 7624
rect 53864 7560 53880 7624
rect 53944 7560 53960 7624
rect 54024 7560 54040 7624
rect 54104 7560 54120 7624
rect 54184 7560 54200 7624
rect 54264 7560 54280 7624
rect 54344 7560 54360 7624
rect 54424 7560 54440 7624
rect 54504 7560 54520 7624
rect 54584 7560 54600 7624
rect 54664 7560 54680 7624
rect 54744 7560 54760 7624
rect 54824 7560 54840 7624
rect 54904 7560 54920 7624
rect 54984 7560 55000 7624
rect 55064 7560 55088 7624
rect 53456 7532 55088 7560
rect 900 5744 2532 5772
rect 900 5680 924 5744
rect 988 5680 1004 5744
rect 1068 5680 1084 5744
rect 1148 5680 1164 5744
rect 1228 5680 1244 5744
rect 1308 5680 1324 5744
rect 1388 5680 1404 5744
rect 1468 5680 1484 5744
rect 1548 5680 1564 5744
rect 1628 5680 1644 5744
rect 1708 5680 1724 5744
rect 1788 5680 1804 5744
rect 1868 5680 1884 5744
rect 1948 5680 1964 5744
rect 2028 5680 2044 5744
rect 2108 5680 2124 5744
rect 2188 5680 2204 5744
rect 2268 5680 2284 5744
rect 2348 5680 2364 5744
rect 2428 5680 2444 5744
rect 2508 5680 2532 5744
rect 900 5652 2532 5680
rect 55904 5744 57536 5772
rect 55904 5680 55928 5744
rect 55992 5680 56008 5744
rect 56072 5680 56088 5744
rect 56152 5680 56168 5744
rect 56232 5680 56248 5744
rect 56312 5680 56328 5744
rect 56392 5680 56408 5744
rect 56472 5680 56488 5744
rect 56552 5680 56568 5744
rect 56632 5680 56648 5744
rect 56712 5680 56728 5744
rect 56792 5680 56808 5744
rect 56872 5680 56888 5744
rect 56952 5680 56968 5744
rect 57032 5680 57048 5744
rect 57112 5680 57128 5744
rect 57192 5680 57208 5744
rect 57272 5680 57288 5744
rect 57352 5680 57368 5744
rect 57432 5680 57448 5744
rect 57512 5680 57536 5744
rect 55904 5652 57536 5680
<< via3 >>
rect 924 50860 988 50864
rect 924 50804 928 50860
rect 928 50804 984 50860
rect 984 50804 988 50860
rect 924 50800 988 50804
rect 1004 50860 1068 50864
rect 1004 50804 1008 50860
rect 1008 50804 1064 50860
rect 1064 50804 1068 50860
rect 1004 50800 1068 50804
rect 1084 50860 1148 50864
rect 1084 50804 1088 50860
rect 1088 50804 1144 50860
rect 1144 50804 1148 50860
rect 1084 50800 1148 50804
rect 1164 50860 1228 50864
rect 1164 50804 1168 50860
rect 1168 50804 1224 50860
rect 1224 50804 1228 50860
rect 1164 50800 1228 50804
rect 1244 50860 1308 50864
rect 1244 50804 1248 50860
rect 1248 50804 1304 50860
rect 1304 50804 1308 50860
rect 1244 50800 1308 50804
rect 1324 50860 1388 50864
rect 1324 50804 1328 50860
rect 1328 50804 1384 50860
rect 1384 50804 1388 50860
rect 1324 50800 1388 50804
rect 1404 50860 1468 50864
rect 1404 50804 1408 50860
rect 1408 50804 1464 50860
rect 1464 50804 1468 50860
rect 1404 50800 1468 50804
rect 1484 50860 1548 50864
rect 1484 50804 1488 50860
rect 1488 50804 1544 50860
rect 1544 50804 1548 50860
rect 1484 50800 1548 50804
rect 1564 50860 1628 50864
rect 1564 50804 1568 50860
rect 1568 50804 1624 50860
rect 1624 50804 1628 50860
rect 1564 50800 1628 50804
rect 1644 50860 1708 50864
rect 1644 50804 1648 50860
rect 1648 50804 1704 50860
rect 1704 50804 1708 50860
rect 1644 50800 1708 50804
rect 1724 50860 1788 50864
rect 1724 50804 1728 50860
rect 1728 50804 1784 50860
rect 1784 50804 1788 50860
rect 1724 50800 1788 50804
rect 1804 50860 1868 50864
rect 1804 50804 1808 50860
rect 1808 50804 1864 50860
rect 1864 50804 1868 50860
rect 1804 50800 1868 50804
rect 1884 50860 1948 50864
rect 1884 50804 1888 50860
rect 1888 50804 1944 50860
rect 1944 50804 1948 50860
rect 1884 50800 1948 50804
rect 1964 50860 2028 50864
rect 1964 50804 1968 50860
rect 1968 50804 2024 50860
rect 2024 50804 2028 50860
rect 1964 50800 2028 50804
rect 2044 50860 2108 50864
rect 2044 50804 2048 50860
rect 2048 50804 2104 50860
rect 2104 50804 2108 50860
rect 2044 50800 2108 50804
rect 2124 50860 2188 50864
rect 2124 50804 2128 50860
rect 2128 50804 2184 50860
rect 2184 50804 2188 50860
rect 2124 50800 2188 50804
rect 2204 50860 2268 50864
rect 2204 50804 2208 50860
rect 2208 50804 2264 50860
rect 2264 50804 2268 50860
rect 2204 50800 2268 50804
rect 2284 50860 2348 50864
rect 2284 50804 2288 50860
rect 2288 50804 2344 50860
rect 2344 50804 2348 50860
rect 2284 50800 2348 50804
rect 2364 50860 2428 50864
rect 2364 50804 2368 50860
rect 2368 50804 2424 50860
rect 2424 50804 2428 50860
rect 2364 50800 2428 50804
rect 2444 50860 2508 50864
rect 2444 50804 2448 50860
rect 2448 50804 2504 50860
rect 2504 50804 2508 50860
rect 2444 50800 2508 50804
rect 55928 50860 55992 50864
rect 55928 50804 55932 50860
rect 55932 50804 55988 50860
rect 55988 50804 55992 50860
rect 55928 50800 55992 50804
rect 56008 50860 56072 50864
rect 56008 50804 56012 50860
rect 56012 50804 56068 50860
rect 56068 50804 56072 50860
rect 56008 50800 56072 50804
rect 56088 50860 56152 50864
rect 56088 50804 56092 50860
rect 56092 50804 56148 50860
rect 56148 50804 56152 50860
rect 56088 50800 56152 50804
rect 56168 50860 56232 50864
rect 56168 50804 56172 50860
rect 56172 50804 56228 50860
rect 56228 50804 56232 50860
rect 56168 50800 56232 50804
rect 56248 50860 56312 50864
rect 56248 50804 56252 50860
rect 56252 50804 56308 50860
rect 56308 50804 56312 50860
rect 56248 50800 56312 50804
rect 56328 50860 56392 50864
rect 56328 50804 56332 50860
rect 56332 50804 56388 50860
rect 56388 50804 56392 50860
rect 56328 50800 56392 50804
rect 56408 50860 56472 50864
rect 56408 50804 56412 50860
rect 56412 50804 56468 50860
rect 56468 50804 56472 50860
rect 56408 50800 56472 50804
rect 56488 50860 56552 50864
rect 56488 50804 56492 50860
rect 56492 50804 56548 50860
rect 56548 50804 56552 50860
rect 56488 50800 56552 50804
rect 56568 50860 56632 50864
rect 56568 50804 56572 50860
rect 56572 50804 56628 50860
rect 56628 50804 56632 50860
rect 56568 50800 56632 50804
rect 56648 50860 56712 50864
rect 56648 50804 56652 50860
rect 56652 50804 56708 50860
rect 56708 50804 56712 50860
rect 56648 50800 56712 50804
rect 56728 50860 56792 50864
rect 56728 50804 56732 50860
rect 56732 50804 56788 50860
rect 56788 50804 56792 50860
rect 56728 50800 56792 50804
rect 56808 50860 56872 50864
rect 56808 50804 56812 50860
rect 56812 50804 56868 50860
rect 56868 50804 56872 50860
rect 56808 50800 56872 50804
rect 56888 50860 56952 50864
rect 56888 50804 56892 50860
rect 56892 50804 56948 50860
rect 56948 50804 56952 50860
rect 56888 50800 56952 50804
rect 56968 50860 57032 50864
rect 56968 50804 56972 50860
rect 56972 50804 57028 50860
rect 57028 50804 57032 50860
rect 56968 50800 57032 50804
rect 57048 50860 57112 50864
rect 57048 50804 57052 50860
rect 57052 50804 57108 50860
rect 57108 50804 57112 50860
rect 57048 50800 57112 50804
rect 57128 50860 57192 50864
rect 57128 50804 57132 50860
rect 57132 50804 57188 50860
rect 57188 50804 57192 50860
rect 57128 50800 57192 50804
rect 57208 50860 57272 50864
rect 57208 50804 57212 50860
rect 57212 50804 57268 50860
rect 57268 50804 57272 50860
rect 57208 50800 57272 50804
rect 57288 50860 57352 50864
rect 57288 50804 57292 50860
rect 57292 50804 57348 50860
rect 57348 50804 57352 50860
rect 57288 50800 57352 50804
rect 57368 50860 57432 50864
rect 57368 50804 57372 50860
rect 57372 50804 57428 50860
rect 57428 50804 57432 50860
rect 57368 50800 57432 50804
rect 57448 50860 57512 50864
rect 57448 50804 57452 50860
rect 57452 50804 57508 50860
rect 57508 50804 57512 50860
rect 57448 50800 57512 50804
rect 3372 48980 3436 48984
rect 3372 48924 3376 48980
rect 3376 48924 3432 48980
rect 3432 48924 3436 48980
rect 3372 48920 3436 48924
rect 3452 48980 3516 48984
rect 3452 48924 3456 48980
rect 3456 48924 3512 48980
rect 3512 48924 3516 48980
rect 3452 48920 3516 48924
rect 3532 48980 3596 48984
rect 3532 48924 3536 48980
rect 3536 48924 3592 48980
rect 3592 48924 3596 48980
rect 3532 48920 3596 48924
rect 3612 48980 3676 48984
rect 3612 48924 3616 48980
rect 3616 48924 3672 48980
rect 3672 48924 3676 48980
rect 3612 48920 3676 48924
rect 3692 48980 3756 48984
rect 3692 48924 3696 48980
rect 3696 48924 3752 48980
rect 3752 48924 3756 48980
rect 3692 48920 3756 48924
rect 3772 48980 3836 48984
rect 3772 48924 3776 48980
rect 3776 48924 3832 48980
rect 3832 48924 3836 48980
rect 3772 48920 3836 48924
rect 3852 48980 3916 48984
rect 3852 48924 3856 48980
rect 3856 48924 3912 48980
rect 3912 48924 3916 48980
rect 3852 48920 3916 48924
rect 3932 48980 3996 48984
rect 3932 48924 3936 48980
rect 3936 48924 3992 48980
rect 3992 48924 3996 48980
rect 3932 48920 3996 48924
rect 4012 48980 4076 48984
rect 4012 48924 4016 48980
rect 4016 48924 4072 48980
rect 4072 48924 4076 48980
rect 4012 48920 4076 48924
rect 4092 48980 4156 48984
rect 4092 48924 4096 48980
rect 4096 48924 4152 48980
rect 4152 48924 4156 48980
rect 4092 48920 4156 48924
rect 4172 48980 4236 48984
rect 4172 48924 4176 48980
rect 4176 48924 4232 48980
rect 4232 48924 4236 48980
rect 4172 48920 4236 48924
rect 4252 48980 4316 48984
rect 4252 48924 4256 48980
rect 4256 48924 4312 48980
rect 4312 48924 4316 48980
rect 4252 48920 4316 48924
rect 4332 48980 4396 48984
rect 4332 48924 4336 48980
rect 4336 48924 4392 48980
rect 4392 48924 4396 48980
rect 4332 48920 4396 48924
rect 4412 48980 4476 48984
rect 4412 48924 4416 48980
rect 4416 48924 4472 48980
rect 4472 48924 4476 48980
rect 4412 48920 4476 48924
rect 4492 48980 4556 48984
rect 4492 48924 4496 48980
rect 4496 48924 4552 48980
rect 4552 48924 4556 48980
rect 4492 48920 4556 48924
rect 4572 48980 4636 48984
rect 4572 48924 4576 48980
rect 4576 48924 4632 48980
rect 4632 48924 4636 48980
rect 4572 48920 4636 48924
rect 4652 48980 4716 48984
rect 4652 48924 4656 48980
rect 4656 48924 4712 48980
rect 4712 48924 4716 48980
rect 4652 48920 4716 48924
rect 4732 48980 4796 48984
rect 4732 48924 4736 48980
rect 4736 48924 4792 48980
rect 4792 48924 4796 48980
rect 4732 48920 4796 48924
rect 4812 48980 4876 48984
rect 4812 48924 4816 48980
rect 4816 48924 4872 48980
rect 4872 48924 4876 48980
rect 4812 48920 4876 48924
rect 4892 48980 4956 48984
rect 4892 48924 4896 48980
rect 4896 48924 4952 48980
rect 4952 48924 4956 48980
rect 4892 48920 4956 48924
rect 53480 48980 53544 48984
rect 53480 48924 53484 48980
rect 53484 48924 53540 48980
rect 53540 48924 53544 48980
rect 53480 48920 53544 48924
rect 53560 48980 53624 48984
rect 53560 48924 53564 48980
rect 53564 48924 53620 48980
rect 53620 48924 53624 48980
rect 53560 48920 53624 48924
rect 53640 48980 53704 48984
rect 53640 48924 53644 48980
rect 53644 48924 53700 48980
rect 53700 48924 53704 48980
rect 53640 48920 53704 48924
rect 53720 48980 53784 48984
rect 53720 48924 53724 48980
rect 53724 48924 53780 48980
rect 53780 48924 53784 48980
rect 53720 48920 53784 48924
rect 53800 48980 53864 48984
rect 53800 48924 53804 48980
rect 53804 48924 53860 48980
rect 53860 48924 53864 48980
rect 53800 48920 53864 48924
rect 53880 48980 53944 48984
rect 53880 48924 53884 48980
rect 53884 48924 53940 48980
rect 53940 48924 53944 48980
rect 53880 48920 53944 48924
rect 53960 48980 54024 48984
rect 53960 48924 53964 48980
rect 53964 48924 54020 48980
rect 54020 48924 54024 48980
rect 53960 48920 54024 48924
rect 54040 48980 54104 48984
rect 54040 48924 54044 48980
rect 54044 48924 54100 48980
rect 54100 48924 54104 48980
rect 54040 48920 54104 48924
rect 54120 48980 54184 48984
rect 54120 48924 54124 48980
rect 54124 48924 54180 48980
rect 54180 48924 54184 48980
rect 54120 48920 54184 48924
rect 54200 48980 54264 48984
rect 54200 48924 54204 48980
rect 54204 48924 54260 48980
rect 54260 48924 54264 48980
rect 54200 48920 54264 48924
rect 54280 48980 54344 48984
rect 54280 48924 54284 48980
rect 54284 48924 54340 48980
rect 54340 48924 54344 48980
rect 54280 48920 54344 48924
rect 54360 48980 54424 48984
rect 54360 48924 54364 48980
rect 54364 48924 54420 48980
rect 54420 48924 54424 48980
rect 54360 48920 54424 48924
rect 54440 48980 54504 48984
rect 54440 48924 54444 48980
rect 54444 48924 54500 48980
rect 54500 48924 54504 48980
rect 54440 48920 54504 48924
rect 54520 48980 54584 48984
rect 54520 48924 54524 48980
rect 54524 48924 54580 48980
rect 54580 48924 54584 48980
rect 54520 48920 54584 48924
rect 54600 48980 54664 48984
rect 54600 48924 54604 48980
rect 54604 48924 54660 48980
rect 54660 48924 54664 48980
rect 54600 48920 54664 48924
rect 54680 48980 54744 48984
rect 54680 48924 54684 48980
rect 54684 48924 54740 48980
rect 54740 48924 54744 48980
rect 54680 48920 54744 48924
rect 54760 48980 54824 48984
rect 54760 48924 54764 48980
rect 54764 48924 54820 48980
rect 54820 48924 54824 48980
rect 54760 48920 54824 48924
rect 54840 48980 54904 48984
rect 54840 48924 54844 48980
rect 54844 48924 54900 48980
rect 54900 48924 54904 48980
rect 54840 48920 54904 48924
rect 54920 48980 54984 48984
rect 54920 48924 54924 48980
rect 54924 48924 54980 48980
rect 54980 48924 54984 48980
rect 54920 48920 54984 48924
rect 55000 48980 55064 48984
rect 55000 48924 55004 48980
rect 55004 48924 55060 48980
rect 55060 48924 55064 48980
rect 55000 48920 55064 48924
rect 6532 48630 6596 48694
rect 7251 48630 7315 48694
rect 7970 48630 8034 48694
rect 8689 48630 8753 48694
rect 9408 48630 9472 48694
rect 10127 48630 10191 48694
rect 10846 48630 10910 48694
rect 11565 48630 11629 48694
rect 12284 48630 12348 48694
rect 13003 48630 13067 48694
rect 6532 48550 6596 48614
rect 7251 48550 7315 48614
rect 7970 48550 8034 48614
rect 8689 48550 8753 48614
rect 9408 48550 9472 48614
rect 10127 48550 10191 48614
rect 10846 48550 10910 48614
rect 11565 48550 11629 48614
rect 12284 48550 12348 48614
rect 13003 48550 13067 48614
rect 6532 48470 6596 48534
rect 7251 48470 7315 48534
rect 7970 48470 8034 48534
rect 8689 48470 8753 48534
rect 9408 48470 9472 48534
rect 10127 48470 10191 48534
rect 10846 48470 10910 48534
rect 11565 48470 11629 48534
rect 12284 48470 12348 48534
rect 13003 48470 13067 48534
rect 6532 48390 6596 48454
rect 7251 48390 7315 48454
rect 7970 48390 8034 48454
rect 8689 48390 8753 48454
rect 9408 48390 9472 48454
rect 10127 48390 10191 48454
rect 10846 48390 10910 48454
rect 11565 48390 11629 48454
rect 12284 48390 12348 48454
rect 13003 48390 13067 48454
rect 6532 48310 6596 48374
rect 7251 48310 7315 48374
rect 7970 48310 8034 48374
rect 8689 48310 8753 48374
rect 9408 48310 9472 48374
rect 10127 48310 10191 48374
rect 10846 48310 10910 48374
rect 11565 48310 11629 48374
rect 12284 48310 12348 48374
rect 13003 48310 13067 48374
rect 6532 48230 6596 48294
rect 7251 48230 7315 48294
rect 7970 48230 8034 48294
rect 8689 48230 8753 48294
rect 9408 48230 9472 48294
rect 10127 48230 10191 48294
rect 10846 48230 10910 48294
rect 11565 48230 11629 48294
rect 12284 48230 12348 48294
rect 13003 48230 13067 48294
rect 6532 48150 6596 48214
rect 7251 48150 7315 48214
rect 7970 48150 8034 48214
rect 8689 48150 8753 48214
rect 9408 48150 9472 48214
rect 10127 48150 10191 48214
rect 10846 48150 10910 48214
rect 11565 48150 11629 48214
rect 12284 48150 12348 48214
rect 13003 48150 13067 48214
rect 6532 47930 6596 47994
rect 7251 47930 7315 47994
rect 7970 47930 8034 47994
rect 8689 47930 8753 47994
rect 9408 47930 9472 47994
rect 10127 47930 10191 47994
rect 10846 47930 10910 47994
rect 11565 47930 11629 47994
rect 12284 47930 12348 47994
rect 13003 47930 13067 47994
rect 6532 47850 6596 47914
rect 7251 47850 7315 47914
rect 7970 47850 8034 47914
rect 8689 47850 8753 47914
rect 9408 47850 9472 47914
rect 10127 47850 10191 47914
rect 10846 47850 10910 47914
rect 11565 47850 11629 47914
rect 12284 47850 12348 47914
rect 13003 47850 13067 47914
rect 6532 47770 6596 47834
rect 7251 47770 7315 47834
rect 7970 47770 8034 47834
rect 8689 47770 8753 47834
rect 9408 47770 9472 47834
rect 10127 47770 10191 47834
rect 10846 47770 10910 47834
rect 11565 47770 11629 47834
rect 12284 47770 12348 47834
rect 13003 47770 13067 47834
rect 6532 47690 6596 47754
rect 7251 47690 7315 47754
rect 7970 47690 8034 47754
rect 8689 47690 8753 47754
rect 9408 47690 9472 47754
rect 10127 47690 10191 47754
rect 10846 47690 10910 47754
rect 11565 47690 11629 47754
rect 12284 47690 12348 47754
rect 13003 47690 13067 47754
rect 6532 47610 6596 47674
rect 7251 47610 7315 47674
rect 7970 47610 8034 47674
rect 8689 47610 8753 47674
rect 9408 47610 9472 47674
rect 10127 47610 10191 47674
rect 10846 47610 10910 47674
rect 11565 47610 11629 47674
rect 12284 47610 12348 47674
rect 13003 47610 13067 47674
rect 6532 47530 6596 47594
rect 7251 47530 7315 47594
rect 7970 47530 8034 47594
rect 8689 47530 8753 47594
rect 9408 47530 9472 47594
rect 10127 47530 10191 47594
rect 10846 47530 10910 47594
rect 11565 47530 11629 47594
rect 12284 47530 12348 47594
rect 13003 47530 13067 47594
rect 6532 47450 6596 47514
rect 7251 47450 7315 47514
rect 7970 47450 8034 47514
rect 8689 47450 8753 47514
rect 9408 47450 9472 47514
rect 10127 47450 10191 47514
rect 10846 47450 10910 47514
rect 11565 47450 11629 47514
rect 12284 47450 12348 47514
rect 13003 47450 13067 47514
rect 13980 48630 14044 48694
rect 14699 48630 14763 48694
rect 15418 48630 15482 48694
rect 16137 48630 16201 48694
rect 16856 48630 16920 48694
rect 17575 48630 17639 48694
rect 18294 48630 18358 48694
rect 19013 48630 19077 48694
rect 19732 48630 19796 48694
rect 20451 48630 20515 48694
rect 13980 48550 14044 48614
rect 14699 48550 14763 48614
rect 15418 48550 15482 48614
rect 16137 48550 16201 48614
rect 16856 48550 16920 48614
rect 17575 48550 17639 48614
rect 18294 48550 18358 48614
rect 19013 48550 19077 48614
rect 19732 48550 19796 48614
rect 20451 48550 20515 48614
rect 13980 48470 14044 48534
rect 14699 48470 14763 48534
rect 15418 48470 15482 48534
rect 16137 48470 16201 48534
rect 16856 48470 16920 48534
rect 17575 48470 17639 48534
rect 18294 48470 18358 48534
rect 19013 48470 19077 48534
rect 19732 48470 19796 48534
rect 20451 48470 20515 48534
rect 13980 48390 14044 48454
rect 14699 48390 14763 48454
rect 15418 48390 15482 48454
rect 16137 48390 16201 48454
rect 16856 48390 16920 48454
rect 17575 48390 17639 48454
rect 18294 48390 18358 48454
rect 19013 48390 19077 48454
rect 19732 48390 19796 48454
rect 20451 48390 20515 48454
rect 13980 48310 14044 48374
rect 14699 48310 14763 48374
rect 15418 48310 15482 48374
rect 16137 48310 16201 48374
rect 16856 48310 16920 48374
rect 17575 48310 17639 48374
rect 18294 48310 18358 48374
rect 19013 48310 19077 48374
rect 19732 48310 19796 48374
rect 20451 48310 20515 48374
rect 13980 48230 14044 48294
rect 14699 48230 14763 48294
rect 15418 48230 15482 48294
rect 16137 48230 16201 48294
rect 16856 48230 16920 48294
rect 17575 48230 17639 48294
rect 18294 48230 18358 48294
rect 19013 48230 19077 48294
rect 19732 48230 19796 48294
rect 20451 48230 20515 48294
rect 13980 48150 14044 48214
rect 14699 48150 14763 48214
rect 15418 48150 15482 48214
rect 16137 48150 16201 48214
rect 16856 48150 16920 48214
rect 17575 48150 17639 48214
rect 18294 48150 18358 48214
rect 19013 48150 19077 48214
rect 19732 48150 19796 48214
rect 20451 48150 20515 48214
rect 13980 47930 14044 47994
rect 14699 47930 14763 47994
rect 15418 47930 15482 47994
rect 16137 47930 16201 47994
rect 16856 47930 16920 47994
rect 17575 47930 17639 47994
rect 18294 47930 18358 47994
rect 19013 47930 19077 47994
rect 19732 47930 19796 47994
rect 20451 47930 20515 47994
rect 13980 47850 14044 47914
rect 14699 47850 14763 47914
rect 15418 47850 15482 47914
rect 16137 47850 16201 47914
rect 16856 47850 16920 47914
rect 17575 47850 17639 47914
rect 18294 47850 18358 47914
rect 19013 47850 19077 47914
rect 19732 47850 19796 47914
rect 20451 47850 20515 47914
rect 13980 47770 14044 47834
rect 14699 47770 14763 47834
rect 15418 47770 15482 47834
rect 16137 47770 16201 47834
rect 16856 47770 16920 47834
rect 17575 47770 17639 47834
rect 18294 47770 18358 47834
rect 19013 47770 19077 47834
rect 19732 47770 19796 47834
rect 20451 47770 20515 47834
rect 13980 47690 14044 47754
rect 14699 47690 14763 47754
rect 15418 47690 15482 47754
rect 16137 47690 16201 47754
rect 16856 47690 16920 47754
rect 17575 47690 17639 47754
rect 18294 47690 18358 47754
rect 19013 47690 19077 47754
rect 19732 47690 19796 47754
rect 20451 47690 20515 47754
rect 13980 47610 14044 47674
rect 14699 47610 14763 47674
rect 15418 47610 15482 47674
rect 16137 47610 16201 47674
rect 16856 47610 16920 47674
rect 17575 47610 17639 47674
rect 18294 47610 18358 47674
rect 19013 47610 19077 47674
rect 19732 47610 19796 47674
rect 20451 47610 20515 47674
rect 13980 47530 14044 47594
rect 14699 47530 14763 47594
rect 15418 47530 15482 47594
rect 16137 47530 16201 47594
rect 16856 47530 16920 47594
rect 17575 47530 17639 47594
rect 18294 47530 18358 47594
rect 19013 47530 19077 47594
rect 19732 47530 19796 47594
rect 20451 47530 20515 47594
rect 13980 47450 14044 47514
rect 14699 47450 14763 47514
rect 15418 47450 15482 47514
rect 16137 47450 16201 47514
rect 16856 47450 16920 47514
rect 17575 47450 17639 47514
rect 18294 47450 18358 47514
rect 19013 47450 19077 47514
rect 19732 47450 19796 47514
rect 20451 47450 20515 47514
rect 5946 47290 6010 47294
rect 6026 47290 6090 47294
rect 5946 47234 5990 47290
rect 5990 47234 6010 47290
rect 6026 47234 6046 47290
rect 6046 47234 6090 47290
rect 5946 47230 6010 47234
rect 6026 47230 6090 47234
rect 13394 47290 13458 47294
rect 13474 47290 13538 47294
rect 13394 47234 13438 47290
rect 13438 47234 13458 47290
rect 13474 47234 13494 47290
rect 13494 47234 13538 47290
rect 13394 47230 13458 47234
rect 13474 47230 13538 47234
rect 924 47100 988 47104
rect 924 47044 928 47100
rect 928 47044 984 47100
rect 984 47044 988 47100
rect 924 47040 988 47044
rect 1004 47100 1068 47104
rect 1004 47044 1008 47100
rect 1008 47044 1064 47100
rect 1064 47044 1068 47100
rect 1004 47040 1068 47044
rect 1084 47100 1148 47104
rect 1084 47044 1088 47100
rect 1088 47044 1144 47100
rect 1144 47044 1148 47100
rect 1084 47040 1148 47044
rect 1164 47100 1228 47104
rect 1164 47044 1168 47100
rect 1168 47044 1224 47100
rect 1224 47044 1228 47100
rect 1164 47040 1228 47044
rect 1244 47100 1308 47104
rect 1244 47044 1248 47100
rect 1248 47044 1304 47100
rect 1304 47044 1308 47100
rect 1244 47040 1308 47044
rect 1324 47100 1388 47104
rect 1324 47044 1328 47100
rect 1328 47044 1384 47100
rect 1384 47044 1388 47100
rect 1324 47040 1388 47044
rect 1404 47100 1468 47104
rect 1404 47044 1408 47100
rect 1408 47044 1464 47100
rect 1464 47044 1468 47100
rect 1404 47040 1468 47044
rect 1484 47100 1548 47104
rect 1484 47044 1488 47100
rect 1488 47044 1544 47100
rect 1544 47044 1548 47100
rect 1484 47040 1548 47044
rect 1564 47100 1628 47104
rect 1564 47044 1568 47100
rect 1568 47044 1624 47100
rect 1624 47044 1628 47100
rect 1564 47040 1628 47044
rect 1644 47100 1708 47104
rect 1644 47044 1648 47100
rect 1648 47044 1704 47100
rect 1704 47044 1708 47100
rect 1644 47040 1708 47044
rect 1724 47100 1788 47104
rect 1724 47044 1728 47100
rect 1728 47044 1784 47100
rect 1784 47044 1788 47100
rect 1724 47040 1788 47044
rect 1804 47100 1868 47104
rect 1804 47044 1808 47100
rect 1808 47044 1864 47100
rect 1864 47044 1868 47100
rect 1804 47040 1868 47044
rect 1884 47100 1948 47104
rect 1884 47044 1888 47100
rect 1888 47044 1944 47100
rect 1944 47044 1948 47100
rect 1884 47040 1948 47044
rect 1964 47100 2028 47104
rect 1964 47044 1968 47100
rect 1968 47044 2024 47100
rect 2024 47044 2028 47100
rect 1964 47040 2028 47044
rect 2044 47100 2108 47104
rect 2044 47044 2048 47100
rect 2048 47044 2104 47100
rect 2104 47044 2108 47100
rect 2044 47040 2108 47044
rect 2124 47100 2188 47104
rect 2124 47044 2128 47100
rect 2128 47044 2184 47100
rect 2184 47044 2188 47100
rect 2124 47040 2188 47044
rect 2204 47100 2268 47104
rect 2204 47044 2208 47100
rect 2208 47044 2264 47100
rect 2264 47044 2268 47100
rect 2204 47040 2268 47044
rect 2284 47100 2348 47104
rect 2284 47044 2288 47100
rect 2288 47044 2344 47100
rect 2344 47044 2348 47100
rect 2284 47040 2348 47044
rect 2364 47100 2428 47104
rect 2364 47044 2368 47100
rect 2368 47044 2424 47100
rect 2424 47044 2428 47100
rect 2364 47040 2428 47044
rect 2444 47100 2508 47104
rect 2444 47044 2448 47100
rect 2448 47044 2504 47100
rect 2504 47044 2508 47100
rect 2444 47040 2508 47044
rect 17678 47132 17742 47136
rect 17678 47076 17682 47132
rect 17682 47076 17738 47132
rect 17738 47076 17742 47132
rect 17678 47072 17742 47076
rect 55928 47100 55992 47104
rect 55928 47044 55932 47100
rect 55932 47044 55988 47100
rect 55988 47044 55992 47100
rect 55928 47040 55992 47044
rect 56008 47100 56072 47104
rect 56008 47044 56012 47100
rect 56012 47044 56068 47100
rect 56068 47044 56072 47100
rect 56008 47040 56072 47044
rect 56088 47100 56152 47104
rect 56088 47044 56092 47100
rect 56092 47044 56148 47100
rect 56148 47044 56152 47100
rect 56088 47040 56152 47044
rect 56168 47100 56232 47104
rect 56168 47044 56172 47100
rect 56172 47044 56228 47100
rect 56228 47044 56232 47100
rect 56168 47040 56232 47044
rect 56248 47100 56312 47104
rect 56248 47044 56252 47100
rect 56252 47044 56308 47100
rect 56308 47044 56312 47100
rect 56248 47040 56312 47044
rect 56328 47100 56392 47104
rect 56328 47044 56332 47100
rect 56332 47044 56388 47100
rect 56388 47044 56392 47100
rect 56328 47040 56392 47044
rect 56408 47100 56472 47104
rect 56408 47044 56412 47100
rect 56412 47044 56468 47100
rect 56468 47044 56472 47100
rect 56408 47040 56472 47044
rect 56488 47100 56552 47104
rect 56488 47044 56492 47100
rect 56492 47044 56548 47100
rect 56548 47044 56552 47100
rect 56488 47040 56552 47044
rect 56568 47100 56632 47104
rect 56568 47044 56572 47100
rect 56572 47044 56628 47100
rect 56628 47044 56632 47100
rect 56568 47040 56632 47044
rect 56648 47100 56712 47104
rect 56648 47044 56652 47100
rect 56652 47044 56708 47100
rect 56708 47044 56712 47100
rect 56648 47040 56712 47044
rect 56728 47100 56792 47104
rect 56728 47044 56732 47100
rect 56732 47044 56788 47100
rect 56788 47044 56792 47100
rect 56728 47040 56792 47044
rect 56808 47100 56872 47104
rect 56808 47044 56812 47100
rect 56812 47044 56868 47100
rect 56868 47044 56872 47100
rect 56808 47040 56872 47044
rect 56888 47100 56952 47104
rect 56888 47044 56892 47100
rect 56892 47044 56948 47100
rect 56948 47044 56952 47100
rect 56888 47040 56952 47044
rect 56968 47100 57032 47104
rect 56968 47044 56972 47100
rect 56972 47044 57028 47100
rect 57028 47044 57032 47100
rect 56968 47040 57032 47044
rect 57048 47100 57112 47104
rect 57048 47044 57052 47100
rect 57052 47044 57108 47100
rect 57108 47044 57112 47100
rect 57048 47040 57112 47044
rect 57128 47100 57192 47104
rect 57128 47044 57132 47100
rect 57132 47044 57188 47100
rect 57188 47044 57192 47100
rect 57128 47040 57192 47044
rect 57208 47100 57272 47104
rect 57208 47044 57212 47100
rect 57212 47044 57268 47100
rect 57268 47044 57272 47100
rect 57208 47040 57272 47044
rect 57288 47100 57352 47104
rect 57288 47044 57292 47100
rect 57292 47044 57348 47100
rect 57348 47044 57352 47100
rect 57288 47040 57352 47044
rect 57368 47100 57432 47104
rect 57368 47044 57372 47100
rect 57372 47044 57428 47100
rect 57428 47044 57432 47100
rect 57368 47040 57432 47044
rect 57448 47100 57512 47104
rect 57448 47044 57452 47100
rect 57452 47044 57508 47100
rect 57508 47044 57512 47100
rect 57448 47040 57512 47044
rect 3372 45220 3436 45224
rect 3372 45164 3376 45220
rect 3376 45164 3432 45220
rect 3432 45164 3436 45220
rect 3372 45160 3436 45164
rect 3452 45220 3516 45224
rect 3452 45164 3456 45220
rect 3456 45164 3512 45220
rect 3512 45164 3516 45220
rect 3452 45160 3516 45164
rect 3532 45220 3596 45224
rect 3532 45164 3536 45220
rect 3536 45164 3592 45220
rect 3592 45164 3596 45220
rect 3532 45160 3596 45164
rect 3612 45220 3676 45224
rect 3612 45164 3616 45220
rect 3616 45164 3672 45220
rect 3672 45164 3676 45220
rect 3612 45160 3676 45164
rect 3692 45220 3756 45224
rect 3692 45164 3696 45220
rect 3696 45164 3752 45220
rect 3752 45164 3756 45220
rect 3692 45160 3756 45164
rect 3772 45220 3836 45224
rect 3772 45164 3776 45220
rect 3776 45164 3832 45220
rect 3832 45164 3836 45220
rect 3772 45160 3836 45164
rect 3852 45220 3916 45224
rect 3852 45164 3856 45220
rect 3856 45164 3912 45220
rect 3912 45164 3916 45220
rect 3852 45160 3916 45164
rect 3932 45220 3996 45224
rect 3932 45164 3936 45220
rect 3936 45164 3992 45220
rect 3992 45164 3996 45220
rect 3932 45160 3996 45164
rect 4012 45220 4076 45224
rect 4012 45164 4016 45220
rect 4016 45164 4072 45220
rect 4072 45164 4076 45220
rect 4012 45160 4076 45164
rect 4092 45220 4156 45224
rect 4092 45164 4096 45220
rect 4096 45164 4152 45220
rect 4152 45164 4156 45220
rect 4092 45160 4156 45164
rect 4172 45220 4236 45224
rect 4172 45164 4176 45220
rect 4176 45164 4232 45220
rect 4232 45164 4236 45220
rect 4172 45160 4236 45164
rect 4252 45220 4316 45224
rect 4252 45164 4256 45220
rect 4256 45164 4312 45220
rect 4312 45164 4316 45220
rect 4252 45160 4316 45164
rect 4332 45220 4396 45224
rect 4332 45164 4336 45220
rect 4336 45164 4392 45220
rect 4392 45164 4396 45220
rect 4332 45160 4396 45164
rect 4412 45220 4476 45224
rect 4412 45164 4416 45220
rect 4416 45164 4472 45220
rect 4472 45164 4476 45220
rect 4412 45160 4476 45164
rect 4492 45220 4556 45224
rect 4492 45164 4496 45220
rect 4496 45164 4552 45220
rect 4552 45164 4556 45220
rect 4492 45160 4556 45164
rect 4572 45220 4636 45224
rect 4572 45164 4576 45220
rect 4576 45164 4632 45220
rect 4632 45164 4636 45220
rect 4572 45160 4636 45164
rect 4652 45220 4716 45224
rect 4652 45164 4656 45220
rect 4656 45164 4712 45220
rect 4712 45164 4716 45220
rect 4652 45160 4716 45164
rect 4732 45220 4796 45224
rect 4732 45164 4736 45220
rect 4736 45164 4792 45220
rect 4792 45164 4796 45220
rect 4732 45160 4796 45164
rect 4812 45220 4876 45224
rect 4812 45164 4816 45220
rect 4816 45164 4872 45220
rect 4872 45164 4876 45220
rect 4812 45160 4876 45164
rect 4892 45220 4956 45224
rect 4892 45164 4896 45220
rect 4896 45164 4952 45220
rect 4952 45164 4956 45220
rect 4892 45160 4956 45164
rect 53480 45220 53544 45224
rect 53480 45164 53484 45220
rect 53484 45164 53540 45220
rect 53540 45164 53544 45220
rect 53480 45160 53544 45164
rect 53560 45220 53624 45224
rect 53560 45164 53564 45220
rect 53564 45164 53620 45220
rect 53620 45164 53624 45220
rect 53560 45160 53624 45164
rect 53640 45220 53704 45224
rect 53640 45164 53644 45220
rect 53644 45164 53700 45220
rect 53700 45164 53704 45220
rect 53640 45160 53704 45164
rect 53720 45220 53784 45224
rect 53720 45164 53724 45220
rect 53724 45164 53780 45220
rect 53780 45164 53784 45220
rect 53720 45160 53784 45164
rect 53800 45220 53864 45224
rect 53800 45164 53804 45220
rect 53804 45164 53860 45220
rect 53860 45164 53864 45220
rect 53800 45160 53864 45164
rect 53880 45220 53944 45224
rect 53880 45164 53884 45220
rect 53884 45164 53940 45220
rect 53940 45164 53944 45220
rect 53880 45160 53944 45164
rect 53960 45220 54024 45224
rect 53960 45164 53964 45220
rect 53964 45164 54020 45220
rect 54020 45164 54024 45220
rect 53960 45160 54024 45164
rect 54040 45220 54104 45224
rect 54040 45164 54044 45220
rect 54044 45164 54100 45220
rect 54100 45164 54104 45220
rect 54040 45160 54104 45164
rect 54120 45220 54184 45224
rect 54120 45164 54124 45220
rect 54124 45164 54180 45220
rect 54180 45164 54184 45220
rect 54120 45160 54184 45164
rect 54200 45220 54264 45224
rect 54200 45164 54204 45220
rect 54204 45164 54260 45220
rect 54260 45164 54264 45220
rect 54200 45160 54264 45164
rect 54280 45220 54344 45224
rect 54280 45164 54284 45220
rect 54284 45164 54340 45220
rect 54340 45164 54344 45220
rect 54280 45160 54344 45164
rect 54360 45220 54424 45224
rect 54360 45164 54364 45220
rect 54364 45164 54420 45220
rect 54420 45164 54424 45220
rect 54360 45160 54424 45164
rect 54440 45220 54504 45224
rect 54440 45164 54444 45220
rect 54444 45164 54500 45220
rect 54500 45164 54504 45220
rect 54440 45160 54504 45164
rect 54520 45220 54584 45224
rect 54520 45164 54524 45220
rect 54524 45164 54580 45220
rect 54580 45164 54584 45220
rect 54520 45160 54584 45164
rect 54600 45220 54664 45224
rect 54600 45164 54604 45220
rect 54604 45164 54660 45220
rect 54660 45164 54664 45220
rect 54600 45160 54664 45164
rect 54680 45220 54744 45224
rect 54680 45164 54684 45220
rect 54684 45164 54740 45220
rect 54740 45164 54744 45220
rect 54680 45160 54744 45164
rect 54760 45220 54824 45224
rect 54760 45164 54764 45220
rect 54764 45164 54820 45220
rect 54820 45164 54824 45220
rect 54760 45160 54824 45164
rect 54840 45220 54904 45224
rect 54840 45164 54844 45220
rect 54844 45164 54900 45220
rect 54900 45164 54904 45220
rect 54840 45160 54904 45164
rect 54920 45220 54984 45224
rect 54920 45164 54924 45220
rect 54924 45164 54980 45220
rect 54980 45164 54984 45220
rect 54920 45160 54984 45164
rect 55000 45220 55064 45224
rect 55000 45164 55004 45220
rect 55004 45164 55060 45220
rect 55060 45164 55064 45220
rect 55000 45160 55064 45164
rect 6532 44870 6596 44934
rect 7251 44870 7315 44934
rect 7970 44870 8034 44934
rect 8689 44870 8753 44934
rect 9408 44870 9472 44934
rect 10127 44870 10191 44934
rect 10846 44870 10910 44934
rect 11565 44870 11629 44934
rect 12284 44870 12348 44934
rect 13003 44870 13067 44934
rect 6532 44790 6596 44854
rect 7251 44790 7315 44854
rect 7970 44790 8034 44854
rect 8689 44790 8753 44854
rect 9408 44790 9472 44854
rect 10127 44790 10191 44854
rect 10846 44790 10910 44854
rect 11565 44790 11629 44854
rect 12284 44790 12348 44854
rect 13003 44790 13067 44854
rect 6532 44710 6596 44774
rect 7251 44710 7315 44774
rect 7970 44710 8034 44774
rect 8689 44710 8753 44774
rect 9408 44710 9472 44774
rect 10127 44710 10191 44774
rect 10846 44710 10910 44774
rect 11565 44710 11629 44774
rect 12284 44710 12348 44774
rect 13003 44710 13067 44774
rect 6532 44630 6596 44694
rect 7251 44630 7315 44694
rect 7970 44630 8034 44694
rect 8689 44630 8753 44694
rect 9408 44630 9472 44694
rect 10127 44630 10191 44694
rect 10846 44630 10910 44694
rect 11565 44630 11629 44694
rect 12284 44630 12348 44694
rect 13003 44630 13067 44694
rect 6532 44550 6596 44614
rect 7251 44550 7315 44614
rect 7970 44550 8034 44614
rect 8689 44550 8753 44614
rect 9408 44550 9472 44614
rect 10127 44550 10191 44614
rect 10846 44550 10910 44614
rect 11565 44550 11629 44614
rect 12284 44550 12348 44614
rect 13003 44550 13067 44614
rect 6532 44470 6596 44534
rect 7251 44470 7315 44534
rect 7970 44470 8034 44534
rect 8689 44470 8753 44534
rect 9408 44470 9472 44534
rect 10127 44470 10191 44534
rect 10846 44470 10910 44534
rect 11565 44470 11629 44534
rect 12284 44470 12348 44534
rect 13003 44470 13067 44534
rect 6532 44390 6596 44454
rect 7251 44390 7315 44454
rect 7970 44390 8034 44454
rect 8689 44390 8753 44454
rect 9408 44390 9472 44454
rect 10127 44390 10191 44454
rect 10846 44390 10910 44454
rect 11565 44390 11629 44454
rect 12284 44390 12348 44454
rect 13003 44390 13067 44454
rect 6532 44170 6596 44234
rect 7251 44170 7315 44234
rect 7970 44170 8034 44234
rect 8689 44170 8753 44234
rect 9408 44170 9472 44234
rect 10127 44170 10191 44234
rect 10846 44170 10910 44234
rect 11565 44170 11629 44234
rect 12284 44170 12348 44234
rect 13003 44170 13067 44234
rect 6532 44090 6596 44154
rect 7251 44090 7315 44154
rect 7970 44090 8034 44154
rect 8689 44090 8753 44154
rect 9408 44090 9472 44154
rect 10127 44090 10191 44154
rect 10846 44090 10910 44154
rect 11565 44090 11629 44154
rect 12284 44090 12348 44154
rect 13003 44090 13067 44154
rect 6532 44010 6596 44074
rect 7251 44010 7315 44074
rect 7970 44010 8034 44074
rect 8689 44010 8753 44074
rect 9408 44010 9472 44074
rect 10127 44010 10191 44074
rect 10846 44010 10910 44074
rect 11565 44010 11629 44074
rect 12284 44010 12348 44074
rect 13003 44010 13067 44074
rect 6532 43930 6596 43994
rect 7251 43930 7315 43994
rect 7970 43930 8034 43994
rect 8689 43930 8753 43994
rect 9408 43930 9472 43994
rect 10127 43930 10191 43994
rect 10846 43930 10910 43994
rect 11565 43930 11629 43994
rect 12284 43930 12348 43994
rect 13003 43930 13067 43994
rect 6532 43850 6596 43914
rect 7251 43850 7315 43914
rect 7970 43850 8034 43914
rect 8689 43850 8753 43914
rect 9408 43850 9472 43914
rect 10127 43850 10191 43914
rect 10846 43850 10910 43914
rect 11565 43850 11629 43914
rect 12284 43850 12348 43914
rect 13003 43850 13067 43914
rect 6532 43770 6596 43834
rect 7251 43770 7315 43834
rect 7970 43770 8034 43834
rect 8689 43770 8753 43834
rect 9408 43770 9472 43834
rect 10127 43770 10191 43834
rect 10846 43770 10910 43834
rect 11565 43770 11629 43834
rect 12284 43770 12348 43834
rect 13003 43770 13067 43834
rect 13400 43778 13464 43842
rect 6532 43690 6596 43754
rect 7251 43690 7315 43754
rect 7970 43690 8034 43754
rect 8689 43690 8753 43754
rect 9408 43690 9472 43754
rect 10127 43690 10191 43754
rect 10846 43690 10910 43754
rect 11565 43690 11629 43754
rect 12284 43690 12348 43754
rect 13003 43690 13067 43754
rect 5946 43530 6010 43534
rect 6026 43530 6090 43534
rect 5946 43474 5990 43530
rect 5990 43474 6010 43530
rect 6026 43474 6046 43530
rect 6046 43474 6090 43530
rect 5946 43470 6010 43474
rect 6026 43470 6090 43474
rect 924 43340 988 43344
rect 924 43284 928 43340
rect 928 43284 984 43340
rect 984 43284 988 43340
rect 924 43280 988 43284
rect 1004 43340 1068 43344
rect 1004 43284 1008 43340
rect 1008 43284 1064 43340
rect 1064 43284 1068 43340
rect 1004 43280 1068 43284
rect 1084 43340 1148 43344
rect 1084 43284 1088 43340
rect 1088 43284 1144 43340
rect 1144 43284 1148 43340
rect 1084 43280 1148 43284
rect 1164 43340 1228 43344
rect 1164 43284 1168 43340
rect 1168 43284 1224 43340
rect 1224 43284 1228 43340
rect 1164 43280 1228 43284
rect 1244 43340 1308 43344
rect 1244 43284 1248 43340
rect 1248 43284 1304 43340
rect 1304 43284 1308 43340
rect 1244 43280 1308 43284
rect 1324 43340 1388 43344
rect 1324 43284 1328 43340
rect 1328 43284 1384 43340
rect 1384 43284 1388 43340
rect 1324 43280 1388 43284
rect 1404 43340 1468 43344
rect 1404 43284 1408 43340
rect 1408 43284 1464 43340
rect 1464 43284 1468 43340
rect 1404 43280 1468 43284
rect 1484 43340 1548 43344
rect 1484 43284 1488 43340
rect 1488 43284 1544 43340
rect 1544 43284 1548 43340
rect 1484 43280 1548 43284
rect 1564 43340 1628 43344
rect 1564 43284 1568 43340
rect 1568 43284 1624 43340
rect 1624 43284 1628 43340
rect 1564 43280 1628 43284
rect 1644 43340 1708 43344
rect 1644 43284 1648 43340
rect 1648 43284 1704 43340
rect 1704 43284 1708 43340
rect 1644 43280 1708 43284
rect 1724 43340 1788 43344
rect 1724 43284 1728 43340
rect 1728 43284 1784 43340
rect 1784 43284 1788 43340
rect 1724 43280 1788 43284
rect 1804 43340 1868 43344
rect 1804 43284 1808 43340
rect 1808 43284 1864 43340
rect 1864 43284 1868 43340
rect 1804 43280 1868 43284
rect 1884 43340 1948 43344
rect 1884 43284 1888 43340
rect 1888 43284 1944 43340
rect 1944 43284 1948 43340
rect 1884 43280 1948 43284
rect 1964 43340 2028 43344
rect 1964 43284 1968 43340
rect 1968 43284 2024 43340
rect 2024 43284 2028 43340
rect 1964 43280 2028 43284
rect 2044 43340 2108 43344
rect 2044 43284 2048 43340
rect 2048 43284 2104 43340
rect 2104 43284 2108 43340
rect 2044 43280 2108 43284
rect 2124 43340 2188 43344
rect 2124 43284 2128 43340
rect 2128 43284 2184 43340
rect 2184 43284 2188 43340
rect 2124 43280 2188 43284
rect 2204 43340 2268 43344
rect 2204 43284 2208 43340
rect 2208 43284 2264 43340
rect 2264 43284 2268 43340
rect 2204 43280 2268 43284
rect 2284 43340 2348 43344
rect 2284 43284 2288 43340
rect 2288 43284 2344 43340
rect 2344 43284 2348 43340
rect 2284 43280 2348 43284
rect 2364 43340 2428 43344
rect 2364 43284 2368 43340
rect 2368 43284 2424 43340
rect 2424 43284 2428 43340
rect 2364 43280 2428 43284
rect 2444 43340 2508 43344
rect 2444 43284 2448 43340
rect 2448 43284 2504 43340
rect 2504 43284 2508 43340
rect 2444 43280 2508 43284
rect 8294 43350 8358 43354
rect 8294 43294 8298 43350
rect 8298 43294 8354 43350
rect 8354 43294 8358 43350
rect 8294 43290 8358 43294
rect 55928 43340 55992 43344
rect 55928 43284 55932 43340
rect 55932 43284 55988 43340
rect 55988 43284 55992 43340
rect 55928 43280 55992 43284
rect 56008 43340 56072 43344
rect 56008 43284 56012 43340
rect 56012 43284 56068 43340
rect 56068 43284 56072 43340
rect 56008 43280 56072 43284
rect 56088 43340 56152 43344
rect 56088 43284 56092 43340
rect 56092 43284 56148 43340
rect 56148 43284 56152 43340
rect 56088 43280 56152 43284
rect 56168 43340 56232 43344
rect 56168 43284 56172 43340
rect 56172 43284 56228 43340
rect 56228 43284 56232 43340
rect 56168 43280 56232 43284
rect 56248 43340 56312 43344
rect 56248 43284 56252 43340
rect 56252 43284 56308 43340
rect 56308 43284 56312 43340
rect 56248 43280 56312 43284
rect 56328 43340 56392 43344
rect 56328 43284 56332 43340
rect 56332 43284 56388 43340
rect 56388 43284 56392 43340
rect 56328 43280 56392 43284
rect 56408 43340 56472 43344
rect 56408 43284 56412 43340
rect 56412 43284 56468 43340
rect 56468 43284 56472 43340
rect 56408 43280 56472 43284
rect 56488 43340 56552 43344
rect 56488 43284 56492 43340
rect 56492 43284 56548 43340
rect 56548 43284 56552 43340
rect 56488 43280 56552 43284
rect 56568 43340 56632 43344
rect 56568 43284 56572 43340
rect 56572 43284 56628 43340
rect 56628 43284 56632 43340
rect 56568 43280 56632 43284
rect 56648 43340 56712 43344
rect 56648 43284 56652 43340
rect 56652 43284 56708 43340
rect 56708 43284 56712 43340
rect 56648 43280 56712 43284
rect 56728 43340 56792 43344
rect 56728 43284 56732 43340
rect 56732 43284 56788 43340
rect 56788 43284 56792 43340
rect 56728 43280 56792 43284
rect 56808 43340 56872 43344
rect 56808 43284 56812 43340
rect 56812 43284 56868 43340
rect 56868 43284 56872 43340
rect 56808 43280 56872 43284
rect 56888 43340 56952 43344
rect 56888 43284 56892 43340
rect 56892 43284 56948 43340
rect 56948 43284 56952 43340
rect 56888 43280 56952 43284
rect 56968 43340 57032 43344
rect 56968 43284 56972 43340
rect 56972 43284 57028 43340
rect 57028 43284 57032 43340
rect 56968 43280 57032 43284
rect 57048 43340 57112 43344
rect 57048 43284 57052 43340
rect 57052 43284 57108 43340
rect 57108 43284 57112 43340
rect 57048 43280 57112 43284
rect 57128 43340 57192 43344
rect 57128 43284 57132 43340
rect 57132 43284 57188 43340
rect 57188 43284 57192 43340
rect 57128 43280 57192 43284
rect 57208 43340 57272 43344
rect 57208 43284 57212 43340
rect 57212 43284 57268 43340
rect 57268 43284 57272 43340
rect 57208 43280 57272 43284
rect 57288 43340 57352 43344
rect 57288 43284 57292 43340
rect 57292 43284 57348 43340
rect 57348 43284 57352 43340
rect 57288 43280 57352 43284
rect 57368 43340 57432 43344
rect 57368 43284 57372 43340
rect 57372 43284 57428 43340
rect 57428 43284 57432 43340
rect 57368 43280 57432 43284
rect 57448 43340 57512 43344
rect 57448 43284 57452 43340
rect 57452 43284 57508 43340
rect 57508 43284 57512 43340
rect 57448 43280 57512 43284
rect 3372 41460 3436 41464
rect 3372 41404 3376 41460
rect 3376 41404 3432 41460
rect 3432 41404 3436 41460
rect 3372 41400 3436 41404
rect 3452 41460 3516 41464
rect 3452 41404 3456 41460
rect 3456 41404 3512 41460
rect 3512 41404 3516 41460
rect 3452 41400 3516 41404
rect 3532 41460 3596 41464
rect 3532 41404 3536 41460
rect 3536 41404 3592 41460
rect 3592 41404 3596 41460
rect 3532 41400 3596 41404
rect 3612 41460 3676 41464
rect 3612 41404 3616 41460
rect 3616 41404 3672 41460
rect 3672 41404 3676 41460
rect 3612 41400 3676 41404
rect 3692 41460 3756 41464
rect 3692 41404 3696 41460
rect 3696 41404 3752 41460
rect 3752 41404 3756 41460
rect 3692 41400 3756 41404
rect 3772 41460 3836 41464
rect 3772 41404 3776 41460
rect 3776 41404 3832 41460
rect 3832 41404 3836 41460
rect 3772 41400 3836 41404
rect 3852 41460 3916 41464
rect 3852 41404 3856 41460
rect 3856 41404 3912 41460
rect 3912 41404 3916 41460
rect 3852 41400 3916 41404
rect 3932 41460 3996 41464
rect 3932 41404 3936 41460
rect 3936 41404 3992 41460
rect 3992 41404 3996 41460
rect 3932 41400 3996 41404
rect 4012 41460 4076 41464
rect 4012 41404 4016 41460
rect 4016 41404 4072 41460
rect 4072 41404 4076 41460
rect 4012 41400 4076 41404
rect 4092 41460 4156 41464
rect 4092 41404 4096 41460
rect 4096 41404 4152 41460
rect 4152 41404 4156 41460
rect 4092 41400 4156 41404
rect 4172 41460 4236 41464
rect 4172 41404 4176 41460
rect 4176 41404 4232 41460
rect 4232 41404 4236 41460
rect 4172 41400 4236 41404
rect 4252 41460 4316 41464
rect 4252 41404 4256 41460
rect 4256 41404 4312 41460
rect 4312 41404 4316 41460
rect 4252 41400 4316 41404
rect 4332 41460 4396 41464
rect 4332 41404 4336 41460
rect 4336 41404 4392 41460
rect 4392 41404 4396 41460
rect 4332 41400 4396 41404
rect 4412 41460 4476 41464
rect 4412 41404 4416 41460
rect 4416 41404 4472 41460
rect 4472 41404 4476 41460
rect 4412 41400 4476 41404
rect 4492 41460 4556 41464
rect 4492 41404 4496 41460
rect 4496 41404 4552 41460
rect 4552 41404 4556 41460
rect 4492 41400 4556 41404
rect 4572 41460 4636 41464
rect 4572 41404 4576 41460
rect 4576 41404 4632 41460
rect 4632 41404 4636 41460
rect 4572 41400 4636 41404
rect 4652 41460 4716 41464
rect 4652 41404 4656 41460
rect 4656 41404 4712 41460
rect 4712 41404 4716 41460
rect 4652 41400 4716 41404
rect 4732 41460 4796 41464
rect 4732 41404 4736 41460
rect 4736 41404 4792 41460
rect 4792 41404 4796 41460
rect 4732 41400 4796 41404
rect 4812 41460 4876 41464
rect 4812 41404 4816 41460
rect 4816 41404 4872 41460
rect 4872 41404 4876 41460
rect 4812 41400 4876 41404
rect 4892 41460 4956 41464
rect 4892 41404 4896 41460
rect 4896 41404 4952 41460
rect 4952 41404 4956 41460
rect 4892 41400 4956 41404
rect 6914 41338 6978 41402
rect 22232 41398 22296 41402
rect 22232 41342 22246 41398
rect 22246 41342 22296 41398
rect 22232 41338 22296 41342
rect 53480 41460 53544 41464
rect 53480 41404 53484 41460
rect 53484 41404 53540 41460
rect 53540 41404 53544 41460
rect 53480 41400 53544 41404
rect 53560 41460 53624 41464
rect 53560 41404 53564 41460
rect 53564 41404 53620 41460
rect 53620 41404 53624 41460
rect 53560 41400 53624 41404
rect 53640 41460 53704 41464
rect 53640 41404 53644 41460
rect 53644 41404 53700 41460
rect 53700 41404 53704 41460
rect 53640 41400 53704 41404
rect 53720 41460 53784 41464
rect 53720 41404 53724 41460
rect 53724 41404 53780 41460
rect 53780 41404 53784 41460
rect 53720 41400 53784 41404
rect 53800 41460 53864 41464
rect 53800 41404 53804 41460
rect 53804 41404 53860 41460
rect 53860 41404 53864 41460
rect 53800 41400 53864 41404
rect 53880 41460 53944 41464
rect 53880 41404 53884 41460
rect 53884 41404 53940 41460
rect 53940 41404 53944 41460
rect 53880 41400 53944 41404
rect 53960 41460 54024 41464
rect 53960 41404 53964 41460
rect 53964 41404 54020 41460
rect 54020 41404 54024 41460
rect 53960 41400 54024 41404
rect 54040 41460 54104 41464
rect 54040 41404 54044 41460
rect 54044 41404 54100 41460
rect 54100 41404 54104 41460
rect 54040 41400 54104 41404
rect 54120 41460 54184 41464
rect 54120 41404 54124 41460
rect 54124 41404 54180 41460
rect 54180 41404 54184 41460
rect 54120 41400 54184 41404
rect 54200 41460 54264 41464
rect 54200 41404 54204 41460
rect 54204 41404 54260 41460
rect 54260 41404 54264 41460
rect 54200 41400 54264 41404
rect 54280 41460 54344 41464
rect 54280 41404 54284 41460
rect 54284 41404 54340 41460
rect 54340 41404 54344 41460
rect 54280 41400 54344 41404
rect 54360 41460 54424 41464
rect 54360 41404 54364 41460
rect 54364 41404 54420 41460
rect 54420 41404 54424 41460
rect 54360 41400 54424 41404
rect 54440 41460 54504 41464
rect 54440 41404 54444 41460
rect 54444 41404 54500 41460
rect 54500 41404 54504 41460
rect 54440 41400 54504 41404
rect 54520 41460 54584 41464
rect 54520 41404 54524 41460
rect 54524 41404 54580 41460
rect 54580 41404 54584 41460
rect 54520 41400 54584 41404
rect 54600 41460 54664 41464
rect 54600 41404 54604 41460
rect 54604 41404 54660 41460
rect 54660 41404 54664 41460
rect 54600 41400 54664 41404
rect 54680 41460 54744 41464
rect 54680 41404 54684 41460
rect 54684 41404 54740 41460
rect 54740 41404 54744 41460
rect 54680 41400 54744 41404
rect 54760 41460 54824 41464
rect 54760 41404 54764 41460
rect 54764 41404 54820 41460
rect 54820 41404 54824 41460
rect 54760 41400 54824 41404
rect 54840 41460 54904 41464
rect 54840 41404 54844 41460
rect 54844 41404 54900 41460
rect 54900 41404 54904 41460
rect 54840 41400 54904 41404
rect 54920 41460 54984 41464
rect 54920 41404 54924 41460
rect 54924 41404 54980 41460
rect 54980 41404 54984 41460
rect 54920 41400 54984 41404
rect 55000 41460 55064 41464
rect 55000 41404 55004 41460
rect 55004 41404 55060 41460
rect 55060 41404 55064 41460
rect 55000 41400 55064 41404
rect 6924 41110 6988 41174
rect 7643 41110 7707 41174
rect 8362 41110 8426 41174
rect 9081 41110 9145 41174
rect 9800 41110 9864 41174
rect 10519 41110 10583 41174
rect 11238 41110 11302 41174
rect 11957 41110 12021 41174
rect 12676 41110 12740 41174
rect 13395 41110 13459 41174
rect 6924 41030 6988 41094
rect 7643 41030 7707 41094
rect 8362 41030 8426 41094
rect 9081 41030 9145 41094
rect 9800 41030 9864 41094
rect 10519 41030 10583 41094
rect 11238 41030 11302 41094
rect 11957 41030 12021 41094
rect 12676 41030 12740 41094
rect 13395 41030 13459 41094
rect 6924 40950 6988 41014
rect 7643 40950 7707 41014
rect 8362 40950 8426 41014
rect 9081 40950 9145 41014
rect 9800 40950 9864 41014
rect 10519 40950 10583 41014
rect 11238 40950 11302 41014
rect 11957 40950 12021 41014
rect 12676 40950 12740 41014
rect 13395 40950 13459 41014
rect 6924 40870 6988 40934
rect 7643 40870 7707 40934
rect 8362 40870 8426 40934
rect 9081 40870 9145 40934
rect 9800 40870 9864 40934
rect 10519 40870 10583 40934
rect 11238 40870 11302 40934
rect 11957 40870 12021 40934
rect 12676 40870 12740 40934
rect 13395 40870 13459 40934
rect 6924 40790 6988 40854
rect 7643 40790 7707 40854
rect 8362 40790 8426 40854
rect 9081 40790 9145 40854
rect 9800 40790 9864 40854
rect 10519 40790 10583 40854
rect 11238 40790 11302 40854
rect 11957 40790 12021 40854
rect 12676 40790 12740 40854
rect 13395 40790 13459 40854
rect 6924 40710 6988 40774
rect 7643 40710 7707 40774
rect 8362 40710 8426 40774
rect 9081 40710 9145 40774
rect 9800 40710 9864 40774
rect 10519 40710 10583 40774
rect 11238 40710 11302 40774
rect 11957 40710 12021 40774
rect 12676 40710 12740 40774
rect 13395 40710 13459 40774
rect 6924 40630 6988 40694
rect 7643 40630 7707 40694
rect 8362 40630 8426 40694
rect 9081 40630 9145 40694
rect 9800 40630 9864 40694
rect 10519 40630 10583 40694
rect 11238 40630 11302 40694
rect 11957 40630 12021 40694
rect 12676 40630 12740 40694
rect 13395 40630 13459 40694
rect 6924 40410 6988 40474
rect 7643 40410 7707 40474
rect 8362 40410 8426 40474
rect 9081 40410 9145 40474
rect 9800 40410 9864 40474
rect 10519 40410 10583 40474
rect 11238 40410 11302 40474
rect 11957 40410 12021 40474
rect 12676 40410 12740 40474
rect 13395 40410 13459 40474
rect 6924 40330 6988 40394
rect 7643 40330 7707 40394
rect 8362 40330 8426 40394
rect 9081 40330 9145 40394
rect 9800 40330 9864 40394
rect 10519 40330 10583 40394
rect 11238 40330 11302 40394
rect 11957 40330 12021 40394
rect 12676 40330 12740 40394
rect 13395 40330 13459 40394
rect 6924 40250 6988 40314
rect 7643 40250 7707 40314
rect 8362 40250 8426 40314
rect 9081 40250 9145 40314
rect 9800 40250 9864 40314
rect 10519 40250 10583 40314
rect 11238 40250 11302 40314
rect 11957 40250 12021 40314
rect 12676 40250 12740 40314
rect 13395 40250 13459 40314
rect 6924 40170 6988 40234
rect 7643 40170 7707 40234
rect 8362 40170 8426 40234
rect 9081 40170 9145 40234
rect 9800 40170 9864 40234
rect 10519 40170 10583 40234
rect 11238 40170 11302 40234
rect 11957 40170 12021 40234
rect 12676 40170 12740 40234
rect 13395 40170 13459 40234
rect 6924 40090 6988 40154
rect 7643 40090 7707 40154
rect 8362 40090 8426 40154
rect 9081 40090 9145 40154
rect 9800 40090 9864 40154
rect 10519 40090 10583 40154
rect 11238 40090 11302 40154
rect 11957 40090 12021 40154
rect 12676 40090 12740 40154
rect 13395 40090 13459 40154
rect 6924 40010 6988 40074
rect 7643 40010 7707 40074
rect 8362 40010 8426 40074
rect 9081 40010 9145 40074
rect 9800 40010 9864 40074
rect 10519 40010 10583 40074
rect 11238 40010 11302 40074
rect 11957 40010 12021 40074
rect 12676 40010 12740 40074
rect 13395 40010 13459 40074
rect 6924 39930 6988 39994
rect 7643 39930 7707 39994
rect 8362 39930 8426 39994
rect 9081 39930 9145 39994
rect 9800 39930 9864 39994
rect 10519 39930 10583 39994
rect 11238 39930 11302 39994
rect 11957 39930 12021 39994
rect 12676 39930 12740 39994
rect 13395 39930 13459 39994
rect 15744 41110 15808 41174
rect 16463 41110 16527 41174
rect 17182 41110 17246 41174
rect 17901 41110 17965 41174
rect 18620 41110 18684 41174
rect 19339 41110 19403 41174
rect 20058 41110 20122 41174
rect 20777 41110 20841 41174
rect 21496 41110 21560 41174
rect 22215 41110 22279 41174
rect 15744 41030 15808 41094
rect 16463 41030 16527 41094
rect 17182 41030 17246 41094
rect 17901 41030 17965 41094
rect 18620 41030 18684 41094
rect 19339 41030 19403 41094
rect 20058 41030 20122 41094
rect 20777 41030 20841 41094
rect 21496 41030 21560 41094
rect 22215 41030 22279 41094
rect 15744 40950 15808 41014
rect 16463 40950 16527 41014
rect 17182 40950 17246 41014
rect 17901 40950 17965 41014
rect 18620 40950 18684 41014
rect 19339 40950 19403 41014
rect 20058 40950 20122 41014
rect 20777 40950 20841 41014
rect 21496 40950 21560 41014
rect 22215 40950 22279 41014
rect 15744 40870 15808 40934
rect 16463 40870 16527 40934
rect 17182 40870 17246 40934
rect 17901 40870 17965 40934
rect 18620 40870 18684 40934
rect 19339 40870 19403 40934
rect 20058 40870 20122 40934
rect 20777 40870 20841 40934
rect 21496 40870 21560 40934
rect 22215 40870 22279 40934
rect 15744 40790 15808 40854
rect 16463 40790 16527 40854
rect 17182 40790 17246 40854
rect 17901 40790 17965 40854
rect 18620 40790 18684 40854
rect 19339 40790 19403 40854
rect 20058 40790 20122 40854
rect 20777 40790 20841 40854
rect 21496 40790 21560 40854
rect 22215 40790 22279 40854
rect 15744 40710 15808 40774
rect 16463 40710 16527 40774
rect 17182 40710 17246 40774
rect 17901 40710 17965 40774
rect 18620 40710 18684 40774
rect 19339 40710 19403 40774
rect 20058 40710 20122 40774
rect 20777 40710 20841 40774
rect 21496 40710 21560 40774
rect 22215 40710 22279 40774
rect 15744 40630 15808 40694
rect 16463 40630 16527 40694
rect 17182 40630 17246 40694
rect 17901 40630 17965 40694
rect 18620 40630 18684 40694
rect 19339 40630 19403 40694
rect 20058 40630 20122 40694
rect 20777 40630 20841 40694
rect 21496 40630 21560 40694
rect 22215 40630 22279 40694
rect 15744 40410 15808 40474
rect 16463 40410 16527 40474
rect 17182 40410 17246 40474
rect 17901 40410 17965 40474
rect 18620 40410 18684 40474
rect 19339 40410 19403 40474
rect 20058 40410 20122 40474
rect 20777 40410 20841 40474
rect 21496 40410 21560 40474
rect 22215 40410 22279 40474
rect 15744 40330 15808 40394
rect 16463 40330 16527 40394
rect 17182 40330 17246 40394
rect 17901 40330 17965 40394
rect 18620 40330 18684 40394
rect 19339 40330 19403 40394
rect 20058 40330 20122 40394
rect 20777 40330 20841 40394
rect 21496 40330 21560 40394
rect 22215 40330 22279 40394
rect 15744 40250 15808 40314
rect 16463 40250 16527 40314
rect 17182 40250 17246 40314
rect 17901 40250 17965 40314
rect 18620 40250 18684 40314
rect 19339 40250 19403 40314
rect 20058 40250 20122 40314
rect 20777 40250 20841 40314
rect 21496 40250 21560 40314
rect 22215 40250 22279 40314
rect 15744 40170 15808 40234
rect 16463 40170 16527 40234
rect 17182 40170 17246 40234
rect 17901 40170 17965 40234
rect 18620 40170 18684 40234
rect 19339 40170 19403 40234
rect 20058 40170 20122 40234
rect 20777 40170 20841 40234
rect 21496 40170 21560 40234
rect 22215 40170 22279 40234
rect 15744 40090 15808 40154
rect 16463 40090 16527 40154
rect 17182 40090 17246 40154
rect 17901 40090 17965 40154
rect 18620 40090 18684 40154
rect 19339 40090 19403 40154
rect 20058 40090 20122 40154
rect 20777 40090 20841 40154
rect 21496 40090 21560 40154
rect 22215 40090 22279 40154
rect 15744 40010 15808 40074
rect 16463 40010 16527 40074
rect 17182 40010 17246 40074
rect 17901 40010 17965 40074
rect 18620 40010 18684 40074
rect 19339 40010 19403 40074
rect 20058 40010 20122 40074
rect 20777 40010 20841 40074
rect 21496 40010 21560 40074
rect 22215 40010 22279 40074
rect 15744 39930 15808 39994
rect 16463 39930 16527 39994
rect 17182 39930 17246 39994
rect 17901 39930 17965 39994
rect 18620 39930 18684 39994
rect 19339 39930 19403 39994
rect 20058 39930 20122 39994
rect 20777 39930 20841 39994
rect 21496 39930 21560 39994
rect 22215 39930 22279 39994
rect 6338 39770 6402 39774
rect 6418 39770 6482 39774
rect 6338 39714 6382 39770
rect 6382 39714 6402 39770
rect 6418 39714 6438 39770
rect 6438 39714 6482 39770
rect 6338 39710 6402 39714
rect 6418 39710 6482 39714
rect 15158 39770 15222 39774
rect 15238 39770 15302 39774
rect 15158 39714 15202 39770
rect 15202 39714 15222 39770
rect 15238 39714 15258 39770
rect 15258 39714 15302 39770
rect 15158 39710 15222 39714
rect 15238 39710 15302 39714
rect 15470 39690 15534 39694
rect 15470 39634 15474 39690
rect 15474 39634 15530 39690
rect 15530 39634 15534 39690
rect 15470 39630 15534 39634
rect 924 39580 988 39584
rect 924 39524 928 39580
rect 928 39524 984 39580
rect 984 39524 988 39580
rect 924 39520 988 39524
rect 1004 39580 1068 39584
rect 1004 39524 1008 39580
rect 1008 39524 1064 39580
rect 1064 39524 1068 39580
rect 1004 39520 1068 39524
rect 1084 39580 1148 39584
rect 1084 39524 1088 39580
rect 1088 39524 1144 39580
rect 1144 39524 1148 39580
rect 1084 39520 1148 39524
rect 1164 39580 1228 39584
rect 1164 39524 1168 39580
rect 1168 39524 1224 39580
rect 1224 39524 1228 39580
rect 1164 39520 1228 39524
rect 1244 39580 1308 39584
rect 1244 39524 1248 39580
rect 1248 39524 1304 39580
rect 1304 39524 1308 39580
rect 1244 39520 1308 39524
rect 1324 39580 1388 39584
rect 1324 39524 1328 39580
rect 1328 39524 1384 39580
rect 1384 39524 1388 39580
rect 1324 39520 1388 39524
rect 1404 39580 1468 39584
rect 1404 39524 1408 39580
rect 1408 39524 1464 39580
rect 1464 39524 1468 39580
rect 1404 39520 1468 39524
rect 1484 39580 1548 39584
rect 1484 39524 1488 39580
rect 1488 39524 1544 39580
rect 1544 39524 1548 39580
rect 1484 39520 1548 39524
rect 1564 39580 1628 39584
rect 1564 39524 1568 39580
rect 1568 39524 1624 39580
rect 1624 39524 1628 39580
rect 1564 39520 1628 39524
rect 1644 39580 1708 39584
rect 1644 39524 1648 39580
rect 1648 39524 1704 39580
rect 1704 39524 1708 39580
rect 1644 39520 1708 39524
rect 1724 39580 1788 39584
rect 1724 39524 1728 39580
rect 1728 39524 1784 39580
rect 1784 39524 1788 39580
rect 1724 39520 1788 39524
rect 1804 39580 1868 39584
rect 1804 39524 1808 39580
rect 1808 39524 1864 39580
rect 1864 39524 1868 39580
rect 1804 39520 1868 39524
rect 1884 39580 1948 39584
rect 1884 39524 1888 39580
rect 1888 39524 1944 39580
rect 1944 39524 1948 39580
rect 1884 39520 1948 39524
rect 1964 39580 2028 39584
rect 1964 39524 1968 39580
rect 1968 39524 2024 39580
rect 2024 39524 2028 39580
rect 1964 39520 2028 39524
rect 2044 39580 2108 39584
rect 2044 39524 2048 39580
rect 2048 39524 2104 39580
rect 2104 39524 2108 39580
rect 2044 39520 2108 39524
rect 2124 39580 2188 39584
rect 2124 39524 2128 39580
rect 2128 39524 2184 39580
rect 2184 39524 2188 39580
rect 2124 39520 2188 39524
rect 2204 39580 2268 39584
rect 2204 39524 2208 39580
rect 2208 39524 2264 39580
rect 2264 39524 2268 39580
rect 2204 39520 2268 39524
rect 2284 39580 2348 39584
rect 2284 39524 2288 39580
rect 2288 39524 2344 39580
rect 2344 39524 2348 39580
rect 2284 39520 2348 39524
rect 2364 39580 2428 39584
rect 2364 39524 2368 39580
rect 2368 39524 2424 39580
rect 2424 39524 2428 39580
rect 2364 39520 2428 39524
rect 2444 39580 2508 39584
rect 2444 39524 2448 39580
rect 2448 39524 2504 39580
rect 2504 39524 2508 39580
rect 2444 39520 2508 39524
rect 55928 39580 55992 39584
rect 55928 39524 55932 39580
rect 55932 39524 55988 39580
rect 55988 39524 55992 39580
rect 55928 39520 55992 39524
rect 56008 39580 56072 39584
rect 56008 39524 56012 39580
rect 56012 39524 56068 39580
rect 56068 39524 56072 39580
rect 56008 39520 56072 39524
rect 56088 39580 56152 39584
rect 56088 39524 56092 39580
rect 56092 39524 56148 39580
rect 56148 39524 56152 39580
rect 56088 39520 56152 39524
rect 56168 39580 56232 39584
rect 56168 39524 56172 39580
rect 56172 39524 56228 39580
rect 56228 39524 56232 39580
rect 56168 39520 56232 39524
rect 56248 39580 56312 39584
rect 56248 39524 56252 39580
rect 56252 39524 56308 39580
rect 56308 39524 56312 39580
rect 56248 39520 56312 39524
rect 56328 39580 56392 39584
rect 56328 39524 56332 39580
rect 56332 39524 56388 39580
rect 56388 39524 56392 39580
rect 56328 39520 56392 39524
rect 56408 39580 56472 39584
rect 56408 39524 56412 39580
rect 56412 39524 56468 39580
rect 56468 39524 56472 39580
rect 56408 39520 56472 39524
rect 56488 39580 56552 39584
rect 56488 39524 56492 39580
rect 56492 39524 56548 39580
rect 56548 39524 56552 39580
rect 56488 39520 56552 39524
rect 56568 39580 56632 39584
rect 56568 39524 56572 39580
rect 56572 39524 56628 39580
rect 56628 39524 56632 39580
rect 56568 39520 56632 39524
rect 56648 39580 56712 39584
rect 56648 39524 56652 39580
rect 56652 39524 56708 39580
rect 56708 39524 56712 39580
rect 56648 39520 56712 39524
rect 56728 39580 56792 39584
rect 56728 39524 56732 39580
rect 56732 39524 56788 39580
rect 56788 39524 56792 39580
rect 56728 39520 56792 39524
rect 56808 39580 56872 39584
rect 56808 39524 56812 39580
rect 56812 39524 56868 39580
rect 56868 39524 56872 39580
rect 56808 39520 56872 39524
rect 56888 39580 56952 39584
rect 56888 39524 56892 39580
rect 56892 39524 56948 39580
rect 56948 39524 56952 39580
rect 56888 39520 56952 39524
rect 56968 39580 57032 39584
rect 56968 39524 56972 39580
rect 56972 39524 57028 39580
rect 57028 39524 57032 39580
rect 56968 39520 57032 39524
rect 57048 39580 57112 39584
rect 57048 39524 57052 39580
rect 57052 39524 57108 39580
rect 57108 39524 57112 39580
rect 57048 39520 57112 39524
rect 57128 39580 57192 39584
rect 57128 39524 57132 39580
rect 57132 39524 57188 39580
rect 57188 39524 57192 39580
rect 57128 39520 57192 39524
rect 57208 39580 57272 39584
rect 57208 39524 57212 39580
rect 57212 39524 57268 39580
rect 57268 39524 57272 39580
rect 57208 39520 57272 39524
rect 57288 39580 57352 39584
rect 57288 39524 57292 39580
rect 57292 39524 57348 39580
rect 57348 39524 57352 39580
rect 57288 39520 57352 39524
rect 57368 39580 57432 39584
rect 57368 39524 57372 39580
rect 57372 39524 57428 39580
rect 57428 39524 57432 39580
rect 57368 39520 57432 39524
rect 57448 39580 57512 39584
rect 57448 39524 57452 39580
rect 57452 39524 57508 39580
rect 57508 39524 57512 39580
rect 57448 39520 57512 39524
rect 3372 37700 3436 37704
rect 3372 37644 3376 37700
rect 3376 37644 3432 37700
rect 3432 37644 3436 37700
rect 3372 37640 3436 37644
rect 3452 37700 3516 37704
rect 3452 37644 3456 37700
rect 3456 37644 3512 37700
rect 3512 37644 3516 37700
rect 3452 37640 3516 37644
rect 3532 37700 3596 37704
rect 3532 37644 3536 37700
rect 3536 37644 3592 37700
rect 3592 37644 3596 37700
rect 3532 37640 3596 37644
rect 3612 37700 3676 37704
rect 3612 37644 3616 37700
rect 3616 37644 3672 37700
rect 3672 37644 3676 37700
rect 3612 37640 3676 37644
rect 3692 37700 3756 37704
rect 3692 37644 3696 37700
rect 3696 37644 3752 37700
rect 3752 37644 3756 37700
rect 3692 37640 3756 37644
rect 3772 37700 3836 37704
rect 3772 37644 3776 37700
rect 3776 37644 3832 37700
rect 3832 37644 3836 37700
rect 3772 37640 3836 37644
rect 3852 37700 3916 37704
rect 3852 37644 3856 37700
rect 3856 37644 3912 37700
rect 3912 37644 3916 37700
rect 3852 37640 3916 37644
rect 3932 37700 3996 37704
rect 3932 37644 3936 37700
rect 3936 37644 3992 37700
rect 3992 37644 3996 37700
rect 3932 37640 3996 37644
rect 4012 37700 4076 37704
rect 4012 37644 4016 37700
rect 4016 37644 4072 37700
rect 4072 37644 4076 37700
rect 4012 37640 4076 37644
rect 4092 37700 4156 37704
rect 4092 37644 4096 37700
rect 4096 37644 4152 37700
rect 4152 37644 4156 37700
rect 4092 37640 4156 37644
rect 4172 37700 4236 37704
rect 4172 37644 4176 37700
rect 4176 37644 4232 37700
rect 4232 37644 4236 37700
rect 4172 37640 4236 37644
rect 4252 37700 4316 37704
rect 4252 37644 4256 37700
rect 4256 37644 4312 37700
rect 4312 37644 4316 37700
rect 4252 37640 4316 37644
rect 4332 37700 4396 37704
rect 4332 37644 4336 37700
rect 4336 37644 4392 37700
rect 4392 37644 4396 37700
rect 4332 37640 4396 37644
rect 4412 37700 4476 37704
rect 4412 37644 4416 37700
rect 4416 37644 4472 37700
rect 4472 37644 4476 37700
rect 4412 37640 4476 37644
rect 4492 37700 4556 37704
rect 4492 37644 4496 37700
rect 4496 37644 4552 37700
rect 4552 37644 4556 37700
rect 4492 37640 4556 37644
rect 4572 37700 4636 37704
rect 4572 37644 4576 37700
rect 4576 37644 4632 37700
rect 4632 37644 4636 37700
rect 4572 37640 4636 37644
rect 4652 37700 4716 37704
rect 4652 37644 4656 37700
rect 4656 37644 4712 37700
rect 4712 37644 4716 37700
rect 4652 37640 4716 37644
rect 4732 37700 4796 37704
rect 4732 37644 4736 37700
rect 4736 37644 4792 37700
rect 4792 37644 4796 37700
rect 4732 37640 4796 37644
rect 4812 37700 4876 37704
rect 4812 37644 4816 37700
rect 4816 37644 4872 37700
rect 4872 37644 4876 37700
rect 4812 37640 4876 37644
rect 4892 37700 4956 37704
rect 4892 37644 4896 37700
rect 4896 37644 4952 37700
rect 4952 37644 4956 37700
rect 4892 37640 4956 37644
rect 53480 37700 53544 37704
rect 53480 37644 53484 37700
rect 53484 37644 53540 37700
rect 53540 37644 53544 37700
rect 53480 37640 53544 37644
rect 53560 37700 53624 37704
rect 53560 37644 53564 37700
rect 53564 37644 53620 37700
rect 53620 37644 53624 37700
rect 53560 37640 53624 37644
rect 53640 37700 53704 37704
rect 53640 37644 53644 37700
rect 53644 37644 53700 37700
rect 53700 37644 53704 37700
rect 53640 37640 53704 37644
rect 53720 37700 53784 37704
rect 53720 37644 53724 37700
rect 53724 37644 53780 37700
rect 53780 37644 53784 37700
rect 53720 37640 53784 37644
rect 53800 37700 53864 37704
rect 53800 37644 53804 37700
rect 53804 37644 53860 37700
rect 53860 37644 53864 37700
rect 53800 37640 53864 37644
rect 53880 37700 53944 37704
rect 53880 37644 53884 37700
rect 53884 37644 53940 37700
rect 53940 37644 53944 37700
rect 53880 37640 53944 37644
rect 53960 37700 54024 37704
rect 53960 37644 53964 37700
rect 53964 37644 54020 37700
rect 54020 37644 54024 37700
rect 53960 37640 54024 37644
rect 54040 37700 54104 37704
rect 54040 37644 54044 37700
rect 54044 37644 54100 37700
rect 54100 37644 54104 37700
rect 54040 37640 54104 37644
rect 54120 37700 54184 37704
rect 54120 37644 54124 37700
rect 54124 37644 54180 37700
rect 54180 37644 54184 37700
rect 54120 37640 54184 37644
rect 54200 37700 54264 37704
rect 54200 37644 54204 37700
rect 54204 37644 54260 37700
rect 54260 37644 54264 37700
rect 54200 37640 54264 37644
rect 54280 37700 54344 37704
rect 54280 37644 54284 37700
rect 54284 37644 54340 37700
rect 54340 37644 54344 37700
rect 54280 37640 54344 37644
rect 54360 37700 54424 37704
rect 54360 37644 54364 37700
rect 54364 37644 54420 37700
rect 54420 37644 54424 37700
rect 54360 37640 54424 37644
rect 54440 37700 54504 37704
rect 54440 37644 54444 37700
rect 54444 37644 54500 37700
rect 54500 37644 54504 37700
rect 54440 37640 54504 37644
rect 54520 37700 54584 37704
rect 54520 37644 54524 37700
rect 54524 37644 54580 37700
rect 54580 37644 54584 37700
rect 54520 37640 54584 37644
rect 54600 37700 54664 37704
rect 54600 37644 54604 37700
rect 54604 37644 54660 37700
rect 54660 37644 54664 37700
rect 54600 37640 54664 37644
rect 54680 37700 54744 37704
rect 54680 37644 54684 37700
rect 54684 37644 54740 37700
rect 54740 37644 54744 37700
rect 54680 37640 54744 37644
rect 54760 37700 54824 37704
rect 54760 37644 54764 37700
rect 54764 37644 54820 37700
rect 54820 37644 54824 37700
rect 54760 37640 54824 37644
rect 54840 37700 54904 37704
rect 54840 37644 54844 37700
rect 54844 37644 54900 37700
rect 54900 37644 54904 37700
rect 54840 37640 54904 37644
rect 54920 37700 54984 37704
rect 54920 37644 54924 37700
rect 54924 37644 54980 37700
rect 54980 37644 54984 37700
rect 54920 37640 54984 37644
rect 55000 37700 55064 37704
rect 55000 37644 55004 37700
rect 55004 37644 55060 37700
rect 55060 37644 55064 37700
rect 55000 37640 55064 37644
rect 33410 37616 33474 37620
rect 33410 37560 33414 37616
rect 33414 37560 33470 37616
rect 33470 37560 33474 37616
rect 33410 37556 33474 37560
rect 30542 37350 30606 37414
rect 31261 37350 31325 37414
rect 31980 37350 32044 37414
rect 32699 37350 32763 37414
rect 33418 37350 33482 37414
rect 34137 37350 34201 37414
rect 34856 37350 34920 37414
rect 35575 37350 35639 37414
rect 36294 37350 36358 37414
rect 37013 37350 37077 37414
rect 30542 37270 30606 37334
rect 31261 37270 31325 37334
rect 31980 37270 32044 37334
rect 32699 37270 32763 37334
rect 33418 37270 33482 37334
rect 34137 37270 34201 37334
rect 34856 37270 34920 37334
rect 35575 37270 35639 37334
rect 36294 37270 36358 37334
rect 37013 37270 37077 37334
rect 13538 37190 13602 37254
rect 30542 37190 30606 37254
rect 31261 37190 31325 37254
rect 31980 37190 32044 37254
rect 32699 37190 32763 37254
rect 33418 37190 33482 37254
rect 34137 37190 34201 37254
rect 34856 37190 34920 37254
rect 35575 37190 35639 37254
rect 36294 37190 36358 37254
rect 37013 37190 37077 37254
rect 30542 37110 30606 37174
rect 31261 37110 31325 37174
rect 31980 37110 32044 37174
rect 32699 37110 32763 37174
rect 33418 37110 33482 37174
rect 34137 37110 34201 37174
rect 34856 37110 34920 37174
rect 35575 37110 35639 37174
rect 36294 37110 36358 37174
rect 37013 37110 37077 37174
rect 30542 37030 30606 37094
rect 31261 37030 31325 37094
rect 31980 37030 32044 37094
rect 32699 37030 32763 37094
rect 33418 37030 33482 37094
rect 34137 37030 34201 37094
rect 34856 37030 34920 37094
rect 35575 37030 35639 37094
rect 36294 37030 36358 37094
rect 37013 37030 37077 37094
rect 29684 36946 29748 37010
rect 30542 36950 30606 37014
rect 31261 36950 31325 37014
rect 31980 36950 32044 37014
rect 32699 36950 32763 37014
rect 33418 36950 33482 37014
rect 34137 36950 34201 37014
rect 34856 36950 34920 37014
rect 35575 36950 35639 37014
rect 36294 36950 36358 37014
rect 37013 36950 37077 37014
rect 30542 36870 30606 36934
rect 31261 36870 31325 36934
rect 31980 36870 32044 36934
rect 32699 36870 32763 36934
rect 33418 36870 33482 36934
rect 34137 36870 34201 36934
rect 34856 36870 34920 36934
rect 35575 36870 35639 36934
rect 36294 36870 36358 36934
rect 37013 36870 37077 36934
rect 30542 36650 30606 36714
rect 31261 36650 31325 36714
rect 31980 36650 32044 36714
rect 32699 36650 32763 36714
rect 33418 36650 33482 36714
rect 34137 36650 34201 36714
rect 34856 36650 34920 36714
rect 35575 36650 35639 36714
rect 36294 36650 36358 36714
rect 37013 36650 37077 36714
rect 30542 36570 30606 36634
rect 31261 36570 31325 36634
rect 31980 36570 32044 36634
rect 32699 36570 32763 36634
rect 33418 36570 33482 36634
rect 34137 36570 34201 36634
rect 34856 36570 34920 36634
rect 35575 36570 35639 36634
rect 36294 36570 36358 36634
rect 37013 36570 37077 36634
rect 30542 36490 30606 36554
rect 31261 36490 31325 36554
rect 31980 36490 32044 36554
rect 32699 36490 32763 36554
rect 33418 36490 33482 36554
rect 34137 36490 34201 36554
rect 34856 36490 34920 36554
rect 35575 36490 35639 36554
rect 36294 36490 36358 36554
rect 37013 36490 37077 36554
rect 30542 36410 30606 36474
rect 31261 36410 31325 36474
rect 31980 36410 32044 36474
rect 32699 36410 32763 36474
rect 33418 36410 33482 36474
rect 34137 36410 34201 36474
rect 34856 36410 34920 36474
rect 35575 36410 35639 36474
rect 36294 36410 36358 36474
rect 37013 36410 37077 36474
rect 30542 36330 30606 36394
rect 31261 36330 31325 36394
rect 31980 36330 32044 36394
rect 32699 36330 32763 36394
rect 33418 36330 33482 36394
rect 34137 36330 34201 36394
rect 34856 36330 34920 36394
rect 35575 36330 35639 36394
rect 36294 36330 36358 36394
rect 37013 36330 37077 36394
rect 30542 36250 30606 36314
rect 31261 36250 31325 36314
rect 31980 36250 32044 36314
rect 32699 36250 32763 36314
rect 33418 36250 33482 36314
rect 34137 36250 34201 36314
rect 34856 36250 34920 36314
rect 35575 36250 35639 36314
rect 36294 36250 36358 36314
rect 37013 36250 37077 36314
rect 30542 36170 30606 36234
rect 31261 36170 31325 36234
rect 31980 36170 32044 36234
rect 32699 36170 32763 36234
rect 33418 36170 33482 36234
rect 34137 36170 34201 36234
rect 34856 36170 34920 36234
rect 35575 36170 35639 36234
rect 36294 36170 36358 36234
rect 37013 36170 37077 36234
rect 29956 36010 30020 36014
rect 30036 36010 30100 36014
rect 29956 35954 30000 36010
rect 30000 35954 30020 36010
rect 30036 35954 30056 36010
rect 30056 35954 30100 36010
rect 29956 35950 30020 35954
rect 30036 35950 30100 35954
rect 37550 36030 37614 36034
rect 37550 35974 37554 36030
rect 37554 35974 37610 36030
rect 37610 35974 37614 36030
rect 37550 35970 37614 35974
rect 924 35820 988 35824
rect 924 35764 928 35820
rect 928 35764 984 35820
rect 984 35764 988 35820
rect 924 35760 988 35764
rect 1004 35820 1068 35824
rect 1004 35764 1008 35820
rect 1008 35764 1064 35820
rect 1064 35764 1068 35820
rect 1004 35760 1068 35764
rect 1084 35820 1148 35824
rect 1084 35764 1088 35820
rect 1088 35764 1144 35820
rect 1144 35764 1148 35820
rect 1084 35760 1148 35764
rect 1164 35820 1228 35824
rect 1164 35764 1168 35820
rect 1168 35764 1224 35820
rect 1224 35764 1228 35820
rect 1164 35760 1228 35764
rect 1244 35820 1308 35824
rect 1244 35764 1248 35820
rect 1248 35764 1304 35820
rect 1304 35764 1308 35820
rect 1244 35760 1308 35764
rect 1324 35820 1388 35824
rect 1324 35764 1328 35820
rect 1328 35764 1384 35820
rect 1384 35764 1388 35820
rect 1324 35760 1388 35764
rect 1404 35820 1468 35824
rect 1404 35764 1408 35820
rect 1408 35764 1464 35820
rect 1464 35764 1468 35820
rect 1404 35760 1468 35764
rect 1484 35820 1548 35824
rect 1484 35764 1488 35820
rect 1488 35764 1544 35820
rect 1544 35764 1548 35820
rect 1484 35760 1548 35764
rect 1564 35820 1628 35824
rect 1564 35764 1568 35820
rect 1568 35764 1624 35820
rect 1624 35764 1628 35820
rect 1564 35760 1628 35764
rect 1644 35820 1708 35824
rect 1644 35764 1648 35820
rect 1648 35764 1704 35820
rect 1704 35764 1708 35820
rect 1644 35760 1708 35764
rect 1724 35820 1788 35824
rect 1724 35764 1728 35820
rect 1728 35764 1784 35820
rect 1784 35764 1788 35820
rect 1724 35760 1788 35764
rect 1804 35820 1868 35824
rect 1804 35764 1808 35820
rect 1808 35764 1864 35820
rect 1864 35764 1868 35820
rect 1804 35760 1868 35764
rect 1884 35820 1948 35824
rect 1884 35764 1888 35820
rect 1888 35764 1944 35820
rect 1944 35764 1948 35820
rect 1884 35760 1948 35764
rect 1964 35820 2028 35824
rect 1964 35764 1968 35820
rect 1968 35764 2024 35820
rect 2024 35764 2028 35820
rect 1964 35760 2028 35764
rect 2044 35820 2108 35824
rect 2044 35764 2048 35820
rect 2048 35764 2104 35820
rect 2104 35764 2108 35820
rect 2044 35760 2108 35764
rect 2124 35820 2188 35824
rect 2124 35764 2128 35820
rect 2128 35764 2184 35820
rect 2184 35764 2188 35820
rect 2124 35760 2188 35764
rect 2204 35820 2268 35824
rect 2204 35764 2208 35820
rect 2208 35764 2264 35820
rect 2264 35764 2268 35820
rect 2204 35760 2268 35764
rect 2284 35820 2348 35824
rect 2284 35764 2288 35820
rect 2288 35764 2344 35820
rect 2344 35764 2348 35820
rect 2284 35760 2348 35764
rect 2364 35820 2428 35824
rect 2364 35764 2368 35820
rect 2368 35764 2424 35820
rect 2424 35764 2428 35820
rect 2364 35760 2428 35764
rect 2444 35820 2508 35824
rect 2444 35764 2448 35820
rect 2448 35764 2504 35820
rect 2504 35764 2508 35820
rect 2444 35760 2508 35764
rect 55928 35820 55992 35824
rect 55928 35764 55932 35820
rect 55932 35764 55988 35820
rect 55988 35764 55992 35820
rect 55928 35760 55992 35764
rect 56008 35820 56072 35824
rect 56008 35764 56012 35820
rect 56012 35764 56068 35820
rect 56068 35764 56072 35820
rect 56008 35760 56072 35764
rect 56088 35820 56152 35824
rect 56088 35764 56092 35820
rect 56092 35764 56148 35820
rect 56148 35764 56152 35820
rect 56088 35760 56152 35764
rect 56168 35820 56232 35824
rect 56168 35764 56172 35820
rect 56172 35764 56228 35820
rect 56228 35764 56232 35820
rect 56168 35760 56232 35764
rect 56248 35820 56312 35824
rect 56248 35764 56252 35820
rect 56252 35764 56308 35820
rect 56308 35764 56312 35820
rect 56248 35760 56312 35764
rect 56328 35820 56392 35824
rect 56328 35764 56332 35820
rect 56332 35764 56388 35820
rect 56388 35764 56392 35820
rect 56328 35760 56392 35764
rect 56408 35820 56472 35824
rect 56408 35764 56412 35820
rect 56412 35764 56468 35820
rect 56468 35764 56472 35820
rect 56408 35760 56472 35764
rect 56488 35820 56552 35824
rect 56488 35764 56492 35820
rect 56492 35764 56548 35820
rect 56548 35764 56552 35820
rect 56488 35760 56552 35764
rect 56568 35820 56632 35824
rect 56568 35764 56572 35820
rect 56572 35764 56628 35820
rect 56628 35764 56632 35820
rect 56568 35760 56632 35764
rect 56648 35820 56712 35824
rect 56648 35764 56652 35820
rect 56652 35764 56708 35820
rect 56708 35764 56712 35820
rect 56648 35760 56712 35764
rect 56728 35820 56792 35824
rect 56728 35764 56732 35820
rect 56732 35764 56788 35820
rect 56788 35764 56792 35820
rect 56728 35760 56792 35764
rect 56808 35820 56872 35824
rect 56808 35764 56812 35820
rect 56812 35764 56868 35820
rect 56868 35764 56872 35820
rect 56808 35760 56872 35764
rect 56888 35820 56952 35824
rect 56888 35764 56892 35820
rect 56892 35764 56948 35820
rect 56948 35764 56952 35820
rect 56888 35760 56952 35764
rect 56968 35820 57032 35824
rect 56968 35764 56972 35820
rect 56972 35764 57028 35820
rect 57028 35764 57032 35820
rect 56968 35760 57032 35764
rect 57048 35820 57112 35824
rect 57048 35764 57052 35820
rect 57052 35764 57108 35820
rect 57108 35764 57112 35820
rect 57048 35760 57112 35764
rect 57128 35820 57192 35824
rect 57128 35764 57132 35820
rect 57132 35764 57188 35820
rect 57188 35764 57192 35820
rect 57128 35760 57192 35764
rect 57208 35820 57272 35824
rect 57208 35764 57212 35820
rect 57212 35764 57268 35820
rect 57268 35764 57272 35820
rect 57208 35760 57272 35764
rect 57288 35820 57352 35824
rect 57288 35764 57292 35820
rect 57292 35764 57348 35820
rect 57348 35764 57352 35820
rect 57288 35760 57352 35764
rect 57368 35820 57432 35824
rect 57368 35764 57372 35820
rect 57372 35764 57428 35820
rect 57428 35764 57432 35820
rect 57368 35760 57432 35764
rect 57448 35820 57512 35824
rect 57448 35764 57452 35820
rect 57452 35764 57508 35820
rect 57508 35764 57512 35820
rect 57448 35760 57512 35764
rect 3372 33940 3436 33944
rect 3372 33884 3376 33940
rect 3376 33884 3432 33940
rect 3432 33884 3436 33940
rect 3372 33880 3436 33884
rect 3452 33940 3516 33944
rect 3452 33884 3456 33940
rect 3456 33884 3512 33940
rect 3512 33884 3516 33940
rect 3452 33880 3516 33884
rect 3532 33940 3596 33944
rect 3532 33884 3536 33940
rect 3536 33884 3592 33940
rect 3592 33884 3596 33940
rect 3532 33880 3596 33884
rect 3612 33940 3676 33944
rect 3612 33884 3616 33940
rect 3616 33884 3672 33940
rect 3672 33884 3676 33940
rect 3612 33880 3676 33884
rect 3692 33940 3756 33944
rect 3692 33884 3696 33940
rect 3696 33884 3752 33940
rect 3752 33884 3756 33940
rect 3692 33880 3756 33884
rect 3772 33940 3836 33944
rect 3772 33884 3776 33940
rect 3776 33884 3832 33940
rect 3832 33884 3836 33940
rect 3772 33880 3836 33884
rect 3852 33940 3916 33944
rect 3852 33884 3856 33940
rect 3856 33884 3912 33940
rect 3912 33884 3916 33940
rect 3852 33880 3916 33884
rect 3932 33940 3996 33944
rect 3932 33884 3936 33940
rect 3936 33884 3992 33940
rect 3992 33884 3996 33940
rect 3932 33880 3996 33884
rect 4012 33940 4076 33944
rect 4012 33884 4016 33940
rect 4016 33884 4072 33940
rect 4072 33884 4076 33940
rect 4012 33880 4076 33884
rect 4092 33940 4156 33944
rect 4092 33884 4096 33940
rect 4096 33884 4152 33940
rect 4152 33884 4156 33940
rect 4092 33880 4156 33884
rect 4172 33940 4236 33944
rect 4172 33884 4176 33940
rect 4176 33884 4232 33940
rect 4232 33884 4236 33940
rect 4172 33880 4236 33884
rect 4252 33940 4316 33944
rect 4252 33884 4256 33940
rect 4256 33884 4312 33940
rect 4312 33884 4316 33940
rect 4252 33880 4316 33884
rect 4332 33940 4396 33944
rect 4332 33884 4336 33940
rect 4336 33884 4392 33940
rect 4392 33884 4396 33940
rect 4332 33880 4396 33884
rect 4412 33940 4476 33944
rect 4412 33884 4416 33940
rect 4416 33884 4472 33940
rect 4472 33884 4476 33940
rect 4412 33880 4476 33884
rect 4492 33940 4556 33944
rect 4492 33884 4496 33940
rect 4496 33884 4552 33940
rect 4552 33884 4556 33940
rect 4492 33880 4556 33884
rect 4572 33940 4636 33944
rect 4572 33884 4576 33940
rect 4576 33884 4632 33940
rect 4632 33884 4636 33940
rect 4572 33880 4636 33884
rect 4652 33940 4716 33944
rect 4652 33884 4656 33940
rect 4656 33884 4712 33940
rect 4712 33884 4716 33940
rect 4652 33880 4716 33884
rect 4732 33940 4796 33944
rect 4732 33884 4736 33940
rect 4736 33884 4792 33940
rect 4792 33884 4796 33940
rect 4732 33880 4796 33884
rect 4812 33940 4876 33944
rect 4812 33884 4816 33940
rect 4816 33884 4872 33940
rect 4872 33884 4876 33940
rect 4812 33880 4876 33884
rect 4892 33940 4956 33944
rect 4892 33884 4896 33940
rect 4896 33884 4952 33940
rect 4952 33884 4956 33940
rect 4892 33880 4956 33884
rect 53480 33940 53544 33944
rect 53480 33884 53484 33940
rect 53484 33884 53540 33940
rect 53540 33884 53544 33940
rect 53480 33880 53544 33884
rect 53560 33940 53624 33944
rect 53560 33884 53564 33940
rect 53564 33884 53620 33940
rect 53620 33884 53624 33940
rect 53560 33880 53624 33884
rect 53640 33940 53704 33944
rect 53640 33884 53644 33940
rect 53644 33884 53700 33940
rect 53700 33884 53704 33940
rect 53640 33880 53704 33884
rect 53720 33940 53784 33944
rect 53720 33884 53724 33940
rect 53724 33884 53780 33940
rect 53780 33884 53784 33940
rect 53720 33880 53784 33884
rect 53800 33940 53864 33944
rect 53800 33884 53804 33940
rect 53804 33884 53860 33940
rect 53860 33884 53864 33940
rect 53800 33880 53864 33884
rect 53880 33940 53944 33944
rect 53880 33884 53884 33940
rect 53884 33884 53940 33940
rect 53940 33884 53944 33940
rect 53880 33880 53944 33884
rect 53960 33940 54024 33944
rect 53960 33884 53964 33940
rect 53964 33884 54020 33940
rect 54020 33884 54024 33940
rect 53960 33880 54024 33884
rect 54040 33940 54104 33944
rect 54040 33884 54044 33940
rect 54044 33884 54100 33940
rect 54100 33884 54104 33940
rect 54040 33880 54104 33884
rect 54120 33940 54184 33944
rect 54120 33884 54124 33940
rect 54124 33884 54180 33940
rect 54180 33884 54184 33940
rect 54120 33880 54184 33884
rect 54200 33940 54264 33944
rect 54200 33884 54204 33940
rect 54204 33884 54260 33940
rect 54260 33884 54264 33940
rect 54200 33880 54264 33884
rect 54280 33940 54344 33944
rect 54280 33884 54284 33940
rect 54284 33884 54340 33940
rect 54340 33884 54344 33940
rect 54280 33880 54344 33884
rect 54360 33940 54424 33944
rect 54360 33884 54364 33940
rect 54364 33884 54420 33940
rect 54420 33884 54424 33940
rect 54360 33880 54424 33884
rect 54440 33940 54504 33944
rect 54440 33884 54444 33940
rect 54444 33884 54500 33940
rect 54500 33884 54504 33940
rect 54440 33880 54504 33884
rect 54520 33940 54584 33944
rect 54520 33884 54524 33940
rect 54524 33884 54580 33940
rect 54580 33884 54584 33940
rect 54520 33880 54584 33884
rect 54600 33940 54664 33944
rect 54600 33884 54604 33940
rect 54604 33884 54660 33940
rect 54660 33884 54664 33940
rect 54600 33880 54664 33884
rect 54680 33940 54744 33944
rect 54680 33884 54684 33940
rect 54684 33884 54740 33940
rect 54740 33884 54744 33940
rect 54680 33880 54744 33884
rect 54760 33940 54824 33944
rect 54760 33884 54764 33940
rect 54764 33884 54820 33940
rect 54820 33884 54824 33940
rect 54760 33880 54824 33884
rect 54840 33940 54904 33944
rect 54840 33884 54844 33940
rect 54844 33884 54900 33940
rect 54900 33884 54904 33940
rect 54840 33880 54904 33884
rect 54920 33940 54984 33944
rect 54920 33884 54924 33940
rect 54924 33884 54980 33940
rect 54980 33884 54984 33940
rect 54920 33880 54984 33884
rect 55000 33940 55064 33944
rect 55000 33884 55004 33940
rect 55004 33884 55060 33940
rect 55060 33884 55064 33940
rect 55000 33880 55064 33884
rect 33272 33774 33336 33838
rect 34100 33774 34164 33838
rect 26818 33590 26882 33654
rect 27537 33590 27601 33654
rect 28256 33590 28320 33654
rect 28975 33590 29039 33654
rect 29694 33590 29758 33654
rect 30413 33590 30477 33654
rect 31132 33590 31196 33654
rect 31851 33590 31915 33654
rect 32570 33590 32634 33654
rect 33289 33590 33353 33654
rect 26818 33510 26882 33574
rect 27537 33510 27601 33574
rect 28256 33510 28320 33574
rect 28975 33510 29039 33574
rect 29694 33510 29758 33574
rect 30413 33510 30477 33574
rect 31132 33510 31196 33574
rect 31851 33510 31915 33574
rect 32570 33510 32634 33574
rect 33289 33510 33353 33574
rect 26818 33430 26882 33494
rect 27537 33430 27601 33494
rect 28256 33430 28320 33494
rect 28975 33430 29039 33494
rect 29694 33430 29758 33494
rect 30413 33430 30477 33494
rect 31132 33430 31196 33494
rect 31851 33430 31915 33494
rect 32570 33430 32634 33494
rect 33289 33430 33353 33494
rect 26818 33350 26882 33414
rect 27537 33350 27601 33414
rect 28256 33350 28320 33414
rect 28975 33350 29039 33414
rect 29694 33350 29758 33414
rect 30413 33350 30477 33414
rect 31132 33350 31196 33414
rect 31851 33350 31915 33414
rect 32570 33350 32634 33414
rect 33289 33350 33353 33414
rect 26818 33270 26882 33334
rect 27537 33270 27601 33334
rect 28256 33270 28320 33334
rect 28975 33270 29039 33334
rect 29694 33270 29758 33334
rect 30413 33270 30477 33334
rect 31132 33270 31196 33334
rect 31851 33270 31915 33334
rect 32570 33270 32634 33334
rect 33289 33270 33353 33334
rect 26818 33190 26882 33254
rect 27537 33190 27601 33254
rect 28256 33190 28320 33254
rect 28975 33190 29039 33254
rect 29694 33190 29758 33254
rect 30413 33190 30477 33254
rect 31132 33190 31196 33254
rect 31851 33190 31915 33254
rect 32570 33190 32634 33254
rect 33289 33190 33353 33254
rect 26818 33110 26882 33174
rect 27537 33110 27601 33174
rect 28256 33110 28320 33174
rect 28975 33110 29039 33174
rect 29694 33110 29758 33174
rect 30413 33110 30477 33174
rect 31132 33110 31196 33174
rect 31851 33110 31915 33174
rect 32570 33110 32634 33174
rect 33289 33110 33353 33174
rect 26818 32890 26882 32954
rect 27537 32890 27601 32954
rect 28256 32890 28320 32954
rect 28975 32890 29039 32954
rect 29694 32890 29758 32954
rect 30413 32890 30477 32954
rect 31132 32890 31196 32954
rect 31851 32890 31915 32954
rect 32570 32890 32634 32954
rect 33289 32890 33353 32954
rect 26818 32810 26882 32874
rect 27537 32810 27601 32874
rect 28256 32810 28320 32874
rect 28975 32810 29039 32874
rect 29694 32810 29758 32874
rect 30413 32810 30477 32874
rect 31132 32810 31196 32874
rect 31851 32810 31915 32874
rect 32570 32810 32634 32874
rect 33289 32810 33353 32874
rect 26818 32730 26882 32794
rect 27537 32730 27601 32794
rect 28256 32730 28320 32794
rect 28975 32730 29039 32794
rect 29694 32730 29758 32794
rect 30413 32730 30477 32794
rect 31132 32730 31196 32794
rect 31851 32730 31915 32794
rect 32570 32730 32634 32794
rect 33289 32730 33353 32794
rect 26818 32650 26882 32714
rect 27537 32650 27601 32714
rect 28256 32650 28320 32714
rect 28975 32650 29039 32714
rect 29694 32650 29758 32714
rect 30413 32650 30477 32714
rect 31132 32650 31196 32714
rect 31851 32650 31915 32714
rect 32570 32650 32634 32714
rect 33289 32650 33353 32714
rect 26818 32570 26882 32634
rect 27537 32570 27601 32634
rect 28256 32570 28320 32634
rect 28975 32570 29039 32634
rect 29694 32570 29758 32634
rect 30413 32570 30477 32634
rect 31132 32570 31196 32634
rect 31851 32570 31915 32634
rect 32570 32570 32634 32634
rect 33289 32570 33353 32634
rect 26818 32490 26882 32554
rect 27537 32490 27601 32554
rect 28256 32490 28320 32554
rect 28975 32490 29039 32554
rect 29694 32490 29758 32554
rect 30413 32490 30477 32554
rect 31132 32490 31196 32554
rect 31851 32490 31915 32554
rect 32570 32490 32634 32554
rect 33289 32490 33353 32554
rect 26818 32410 26882 32474
rect 27537 32410 27601 32474
rect 28256 32410 28320 32474
rect 28975 32410 29039 32474
rect 29694 32410 29758 32474
rect 30413 32410 30477 32474
rect 31132 32410 31196 32474
rect 31851 32410 31915 32474
rect 32570 32410 32634 32474
rect 33289 32410 33353 32474
rect 34266 33590 34330 33654
rect 34985 33590 35049 33654
rect 35704 33590 35768 33654
rect 36423 33590 36487 33654
rect 37142 33590 37206 33654
rect 37861 33590 37925 33654
rect 38580 33590 38644 33654
rect 39299 33590 39363 33654
rect 40018 33590 40082 33654
rect 40737 33590 40801 33654
rect 34266 33510 34330 33574
rect 34985 33510 35049 33574
rect 35704 33510 35768 33574
rect 36423 33510 36487 33574
rect 37142 33510 37206 33574
rect 37861 33510 37925 33574
rect 38580 33510 38644 33574
rect 39299 33510 39363 33574
rect 40018 33510 40082 33574
rect 40737 33510 40801 33574
rect 34266 33430 34330 33494
rect 34985 33430 35049 33494
rect 35704 33430 35768 33494
rect 36423 33430 36487 33494
rect 37142 33430 37206 33494
rect 37861 33430 37925 33494
rect 38580 33430 38644 33494
rect 39299 33430 39363 33494
rect 40018 33430 40082 33494
rect 40737 33430 40801 33494
rect 34266 33350 34330 33414
rect 34985 33350 35049 33414
rect 35704 33350 35768 33414
rect 36423 33350 36487 33414
rect 37142 33350 37206 33414
rect 37861 33350 37925 33414
rect 38580 33350 38644 33414
rect 39299 33350 39363 33414
rect 40018 33350 40082 33414
rect 40737 33350 40801 33414
rect 34266 33270 34330 33334
rect 34985 33270 35049 33334
rect 35704 33270 35768 33334
rect 36423 33270 36487 33334
rect 37142 33270 37206 33334
rect 37861 33270 37925 33334
rect 38580 33270 38644 33334
rect 39299 33270 39363 33334
rect 40018 33270 40082 33334
rect 40737 33270 40801 33334
rect 34266 33190 34330 33254
rect 34985 33190 35049 33254
rect 35704 33190 35768 33254
rect 36423 33190 36487 33254
rect 37142 33190 37206 33254
rect 37861 33190 37925 33254
rect 38580 33190 38644 33254
rect 39299 33190 39363 33254
rect 40018 33190 40082 33254
rect 40737 33190 40801 33254
rect 34266 33110 34330 33174
rect 34985 33110 35049 33174
rect 35704 33110 35768 33174
rect 36423 33110 36487 33174
rect 37142 33110 37206 33174
rect 37861 33110 37925 33174
rect 38580 33110 38644 33174
rect 39299 33110 39363 33174
rect 40018 33110 40082 33174
rect 40737 33110 40801 33174
rect 34266 32890 34330 32954
rect 34985 32890 35049 32954
rect 35704 32890 35768 32954
rect 36423 32890 36487 32954
rect 37142 32890 37206 32954
rect 37861 32890 37925 32954
rect 38580 32890 38644 32954
rect 39299 32890 39363 32954
rect 40018 32890 40082 32954
rect 40737 32890 40801 32954
rect 34266 32810 34330 32874
rect 34985 32810 35049 32874
rect 35704 32810 35768 32874
rect 36423 32810 36487 32874
rect 37142 32810 37206 32874
rect 37861 32810 37925 32874
rect 38580 32810 38644 32874
rect 39299 32810 39363 32874
rect 40018 32810 40082 32874
rect 40737 32810 40801 32874
rect 34266 32730 34330 32794
rect 34985 32730 35049 32794
rect 35704 32730 35768 32794
rect 36423 32730 36487 32794
rect 37142 32730 37206 32794
rect 37861 32730 37925 32794
rect 38580 32730 38644 32794
rect 39299 32730 39363 32794
rect 40018 32730 40082 32794
rect 40737 32730 40801 32794
rect 34266 32650 34330 32714
rect 34985 32650 35049 32714
rect 35704 32650 35768 32714
rect 36423 32650 36487 32714
rect 37142 32650 37206 32714
rect 37861 32650 37925 32714
rect 38580 32650 38644 32714
rect 39299 32650 39363 32714
rect 40018 32650 40082 32714
rect 40737 32650 40801 32714
rect 34266 32570 34330 32634
rect 34985 32570 35049 32634
rect 35704 32570 35768 32634
rect 36423 32570 36487 32634
rect 37142 32570 37206 32634
rect 37861 32570 37925 32634
rect 38580 32570 38644 32634
rect 39299 32570 39363 32634
rect 40018 32570 40082 32634
rect 40737 32570 40801 32634
rect 34266 32490 34330 32554
rect 34985 32490 35049 32554
rect 35704 32490 35768 32554
rect 36423 32490 36487 32554
rect 37142 32490 37206 32554
rect 37861 32490 37925 32554
rect 38580 32490 38644 32554
rect 39299 32490 39363 32554
rect 40018 32490 40082 32554
rect 40737 32490 40801 32554
rect 34266 32410 34330 32474
rect 34985 32410 35049 32474
rect 35704 32410 35768 32474
rect 36423 32410 36487 32474
rect 37142 32410 37206 32474
rect 37861 32410 37925 32474
rect 38580 32410 38644 32474
rect 39299 32410 39363 32474
rect 40018 32410 40082 32474
rect 40737 32410 40801 32474
rect 26232 32250 26296 32254
rect 26312 32250 26376 32254
rect 26232 32194 26276 32250
rect 26276 32194 26296 32250
rect 26312 32194 26332 32250
rect 26332 32194 26376 32250
rect 26232 32190 26296 32194
rect 26312 32190 26376 32194
rect 33680 32250 33744 32254
rect 33760 32250 33824 32254
rect 33680 32194 33724 32250
rect 33724 32194 33744 32250
rect 33760 32194 33780 32250
rect 33780 32194 33824 32250
rect 33680 32190 33744 32194
rect 33760 32190 33824 32194
rect 924 32060 988 32064
rect 924 32004 928 32060
rect 928 32004 984 32060
rect 984 32004 988 32060
rect 924 32000 988 32004
rect 1004 32060 1068 32064
rect 1004 32004 1008 32060
rect 1008 32004 1064 32060
rect 1064 32004 1068 32060
rect 1004 32000 1068 32004
rect 1084 32060 1148 32064
rect 1084 32004 1088 32060
rect 1088 32004 1144 32060
rect 1144 32004 1148 32060
rect 1084 32000 1148 32004
rect 1164 32060 1228 32064
rect 1164 32004 1168 32060
rect 1168 32004 1224 32060
rect 1224 32004 1228 32060
rect 1164 32000 1228 32004
rect 1244 32060 1308 32064
rect 1244 32004 1248 32060
rect 1248 32004 1304 32060
rect 1304 32004 1308 32060
rect 1244 32000 1308 32004
rect 1324 32060 1388 32064
rect 1324 32004 1328 32060
rect 1328 32004 1384 32060
rect 1384 32004 1388 32060
rect 1324 32000 1388 32004
rect 1404 32060 1468 32064
rect 1404 32004 1408 32060
rect 1408 32004 1464 32060
rect 1464 32004 1468 32060
rect 1404 32000 1468 32004
rect 1484 32060 1548 32064
rect 1484 32004 1488 32060
rect 1488 32004 1544 32060
rect 1544 32004 1548 32060
rect 1484 32000 1548 32004
rect 1564 32060 1628 32064
rect 1564 32004 1568 32060
rect 1568 32004 1624 32060
rect 1624 32004 1628 32060
rect 1564 32000 1628 32004
rect 1644 32060 1708 32064
rect 1644 32004 1648 32060
rect 1648 32004 1704 32060
rect 1704 32004 1708 32060
rect 1644 32000 1708 32004
rect 1724 32060 1788 32064
rect 1724 32004 1728 32060
rect 1728 32004 1784 32060
rect 1784 32004 1788 32060
rect 1724 32000 1788 32004
rect 1804 32060 1868 32064
rect 1804 32004 1808 32060
rect 1808 32004 1864 32060
rect 1864 32004 1868 32060
rect 1804 32000 1868 32004
rect 1884 32060 1948 32064
rect 1884 32004 1888 32060
rect 1888 32004 1944 32060
rect 1944 32004 1948 32060
rect 1884 32000 1948 32004
rect 1964 32060 2028 32064
rect 1964 32004 1968 32060
rect 1968 32004 2024 32060
rect 2024 32004 2028 32060
rect 1964 32000 2028 32004
rect 2044 32060 2108 32064
rect 2044 32004 2048 32060
rect 2048 32004 2104 32060
rect 2104 32004 2108 32060
rect 2044 32000 2108 32004
rect 2124 32060 2188 32064
rect 2124 32004 2128 32060
rect 2128 32004 2184 32060
rect 2184 32004 2188 32060
rect 2124 32000 2188 32004
rect 2204 32060 2268 32064
rect 2204 32004 2208 32060
rect 2208 32004 2264 32060
rect 2264 32004 2268 32060
rect 2204 32000 2268 32004
rect 2284 32060 2348 32064
rect 2284 32004 2288 32060
rect 2288 32004 2344 32060
rect 2344 32004 2348 32060
rect 2284 32000 2348 32004
rect 2364 32060 2428 32064
rect 2364 32004 2368 32060
rect 2368 32004 2424 32060
rect 2424 32004 2428 32060
rect 2364 32000 2428 32004
rect 2444 32060 2508 32064
rect 2444 32004 2448 32060
rect 2448 32004 2504 32060
rect 2504 32004 2508 32060
rect 2444 32000 2508 32004
rect 55928 32060 55992 32064
rect 55928 32004 55932 32060
rect 55932 32004 55988 32060
rect 55988 32004 55992 32060
rect 55928 32000 55992 32004
rect 56008 32060 56072 32064
rect 56008 32004 56012 32060
rect 56012 32004 56068 32060
rect 56068 32004 56072 32060
rect 56008 32000 56072 32004
rect 56088 32060 56152 32064
rect 56088 32004 56092 32060
rect 56092 32004 56148 32060
rect 56148 32004 56152 32060
rect 56088 32000 56152 32004
rect 56168 32060 56232 32064
rect 56168 32004 56172 32060
rect 56172 32004 56228 32060
rect 56228 32004 56232 32060
rect 56168 32000 56232 32004
rect 56248 32060 56312 32064
rect 56248 32004 56252 32060
rect 56252 32004 56308 32060
rect 56308 32004 56312 32060
rect 56248 32000 56312 32004
rect 56328 32060 56392 32064
rect 56328 32004 56332 32060
rect 56332 32004 56388 32060
rect 56388 32004 56392 32060
rect 56328 32000 56392 32004
rect 56408 32060 56472 32064
rect 56408 32004 56412 32060
rect 56412 32004 56468 32060
rect 56468 32004 56472 32060
rect 56408 32000 56472 32004
rect 56488 32060 56552 32064
rect 56488 32004 56492 32060
rect 56492 32004 56548 32060
rect 56548 32004 56552 32060
rect 56488 32000 56552 32004
rect 56568 32060 56632 32064
rect 56568 32004 56572 32060
rect 56572 32004 56628 32060
rect 56628 32004 56632 32060
rect 56568 32000 56632 32004
rect 56648 32060 56712 32064
rect 56648 32004 56652 32060
rect 56652 32004 56708 32060
rect 56708 32004 56712 32060
rect 56648 32000 56712 32004
rect 56728 32060 56792 32064
rect 56728 32004 56732 32060
rect 56732 32004 56788 32060
rect 56788 32004 56792 32060
rect 56728 32000 56792 32004
rect 56808 32060 56872 32064
rect 56808 32004 56812 32060
rect 56812 32004 56868 32060
rect 56868 32004 56872 32060
rect 56808 32000 56872 32004
rect 56888 32060 56952 32064
rect 56888 32004 56892 32060
rect 56892 32004 56948 32060
rect 56948 32004 56952 32060
rect 56888 32000 56952 32004
rect 56968 32060 57032 32064
rect 56968 32004 56972 32060
rect 56972 32004 57028 32060
rect 57028 32004 57032 32060
rect 56968 32000 57032 32004
rect 57048 32060 57112 32064
rect 57048 32004 57052 32060
rect 57052 32004 57108 32060
rect 57108 32004 57112 32060
rect 57048 32000 57112 32004
rect 57128 32060 57192 32064
rect 57128 32004 57132 32060
rect 57132 32004 57188 32060
rect 57188 32004 57192 32060
rect 57128 32000 57192 32004
rect 57208 32060 57272 32064
rect 57208 32004 57212 32060
rect 57212 32004 57268 32060
rect 57268 32004 57272 32060
rect 57208 32000 57272 32004
rect 57288 32060 57352 32064
rect 57288 32004 57292 32060
rect 57292 32004 57348 32060
rect 57348 32004 57352 32060
rect 57288 32000 57352 32004
rect 57368 32060 57432 32064
rect 57368 32004 57372 32060
rect 57372 32004 57428 32060
rect 57428 32004 57432 32060
rect 57368 32000 57432 32004
rect 57448 32060 57512 32064
rect 57448 32004 57452 32060
rect 57452 32004 57508 32060
rect 57508 32004 57512 32060
rect 57448 32000 57512 32004
rect 3372 30180 3436 30184
rect 3372 30124 3376 30180
rect 3376 30124 3432 30180
rect 3432 30124 3436 30180
rect 3372 30120 3436 30124
rect 3452 30180 3516 30184
rect 3452 30124 3456 30180
rect 3456 30124 3512 30180
rect 3512 30124 3516 30180
rect 3452 30120 3516 30124
rect 3532 30180 3596 30184
rect 3532 30124 3536 30180
rect 3536 30124 3592 30180
rect 3592 30124 3596 30180
rect 3532 30120 3596 30124
rect 3612 30180 3676 30184
rect 3612 30124 3616 30180
rect 3616 30124 3672 30180
rect 3672 30124 3676 30180
rect 3612 30120 3676 30124
rect 3692 30180 3756 30184
rect 3692 30124 3696 30180
rect 3696 30124 3752 30180
rect 3752 30124 3756 30180
rect 3692 30120 3756 30124
rect 3772 30180 3836 30184
rect 3772 30124 3776 30180
rect 3776 30124 3832 30180
rect 3832 30124 3836 30180
rect 3772 30120 3836 30124
rect 3852 30180 3916 30184
rect 3852 30124 3856 30180
rect 3856 30124 3912 30180
rect 3912 30124 3916 30180
rect 3852 30120 3916 30124
rect 3932 30180 3996 30184
rect 3932 30124 3936 30180
rect 3936 30124 3992 30180
rect 3992 30124 3996 30180
rect 3932 30120 3996 30124
rect 4012 30180 4076 30184
rect 4012 30124 4016 30180
rect 4016 30124 4072 30180
rect 4072 30124 4076 30180
rect 4012 30120 4076 30124
rect 4092 30180 4156 30184
rect 4092 30124 4096 30180
rect 4096 30124 4152 30180
rect 4152 30124 4156 30180
rect 4092 30120 4156 30124
rect 4172 30180 4236 30184
rect 4172 30124 4176 30180
rect 4176 30124 4232 30180
rect 4232 30124 4236 30180
rect 4172 30120 4236 30124
rect 4252 30180 4316 30184
rect 4252 30124 4256 30180
rect 4256 30124 4312 30180
rect 4312 30124 4316 30180
rect 4252 30120 4316 30124
rect 4332 30180 4396 30184
rect 4332 30124 4336 30180
rect 4336 30124 4392 30180
rect 4392 30124 4396 30180
rect 4332 30120 4396 30124
rect 4412 30180 4476 30184
rect 4412 30124 4416 30180
rect 4416 30124 4472 30180
rect 4472 30124 4476 30180
rect 4412 30120 4476 30124
rect 4492 30180 4556 30184
rect 4492 30124 4496 30180
rect 4496 30124 4552 30180
rect 4552 30124 4556 30180
rect 4492 30120 4556 30124
rect 4572 30180 4636 30184
rect 4572 30124 4576 30180
rect 4576 30124 4632 30180
rect 4632 30124 4636 30180
rect 4572 30120 4636 30124
rect 4652 30180 4716 30184
rect 4652 30124 4656 30180
rect 4656 30124 4712 30180
rect 4712 30124 4716 30180
rect 4652 30120 4716 30124
rect 4732 30180 4796 30184
rect 4732 30124 4736 30180
rect 4736 30124 4792 30180
rect 4792 30124 4796 30180
rect 4732 30120 4796 30124
rect 4812 30180 4876 30184
rect 4812 30124 4816 30180
rect 4816 30124 4872 30180
rect 4872 30124 4876 30180
rect 4812 30120 4876 30124
rect 4892 30180 4956 30184
rect 4892 30124 4896 30180
rect 4896 30124 4952 30180
rect 4952 30124 4956 30180
rect 4892 30120 4956 30124
rect 33410 30174 33474 30178
rect 33410 30118 33414 30174
rect 33414 30118 33470 30174
rect 33470 30118 33474 30174
rect 33410 30114 33474 30118
rect 53480 30180 53544 30184
rect 53480 30124 53484 30180
rect 53484 30124 53540 30180
rect 53540 30124 53544 30180
rect 53480 30120 53544 30124
rect 53560 30180 53624 30184
rect 53560 30124 53564 30180
rect 53564 30124 53620 30180
rect 53620 30124 53624 30180
rect 53560 30120 53624 30124
rect 53640 30180 53704 30184
rect 53640 30124 53644 30180
rect 53644 30124 53700 30180
rect 53700 30124 53704 30180
rect 53640 30120 53704 30124
rect 53720 30180 53784 30184
rect 53720 30124 53724 30180
rect 53724 30124 53780 30180
rect 53780 30124 53784 30180
rect 53720 30120 53784 30124
rect 53800 30180 53864 30184
rect 53800 30124 53804 30180
rect 53804 30124 53860 30180
rect 53860 30124 53864 30180
rect 53800 30120 53864 30124
rect 53880 30180 53944 30184
rect 53880 30124 53884 30180
rect 53884 30124 53940 30180
rect 53940 30124 53944 30180
rect 53880 30120 53944 30124
rect 53960 30180 54024 30184
rect 53960 30124 53964 30180
rect 53964 30124 54020 30180
rect 54020 30124 54024 30180
rect 53960 30120 54024 30124
rect 54040 30180 54104 30184
rect 54040 30124 54044 30180
rect 54044 30124 54100 30180
rect 54100 30124 54104 30180
rect 54040 30120 54104 30124
rect 54120 30180 54184 30184
rect 54120 30124 54124 30180
rect 54124 30124 54180 30180
rect 54180 30124 54184 30180
rect 54120 30120 54184 30124
rect 54200 30180 54264 30184
rect 54200 30124 54204 30180
rect 54204 30124 54260 30180
rect 54260 30124 54264 30180
rect 54200 30120 54264 30124
rect 54280 30180 54344 30184
rect 54280 30124 54284 30180
rect 54284 30124 54340 30180
rect 54340 30124 54344 30180
rect 54280 30120 54344 30124
rect 54360 30180 54424 30184
rect 54360 30124 54364 30180
rect 54364 30124 54420 30180
rect 54420 30124 54424 30180
rect 54360 30120 54424 30124
rect 54440 30180 54504 30184
rect 54440 30124 54444 30180
rect 54444 30124 54500 30180
rect 54500 30124 54504 30180
rect 54440 30120 54504 30124
rect 54520 30180 54584 30184
rect 54520 30124 54524 30180
rect 54524 30124 54580 30180
rect 54580 30124 54584 30180
rect 54520 30120 54584 30124
rect 54600 30180 54664 30184
rect 54600 30124 54604 30180
rect 54604 30124 54660 30180
rect 54660 30124 54664 30180
rect 54600 30120 54664 30124
rect 54680 30180 54744 30184
rect 54680 30124 54684 30180
rect 54684 30124 54740 30180
rect 54740 30124 54744 30180
rect 54680 30120 54744 30124
rect 54760 30180 54824 30184
rect 54760 30124 54764 30180
rect 54764 30124 54820 30180
rect 54820 30124 54824 30180
rect 54760 30120 54824 30124
rect 54840 30180 54904 30184
rect 54840 30124 54844 30180
rect 54844 30124 54900 30180
rect 54900 30124 54904 30180
rect 54840 30120 54904 30124
rect 54920 30180 54984 30184
rect 54920 30124 54924 30180
rect 54924 30124 54980 30180
rect 54980 30124 54984 30180
rect 54920 30120 54984 30124
rect 55000 30180 55064 30184
rect 55000 30124 55004 30180
rect 55004 30124 55060 30180
rect 55060 30124 55064 30180
rect 55000 30120 55064 30124
rect 30542 29830 30606 29894
rect 31261 29830 31325 29894
rect 31980 29830 32044 29894
rect 32699 29830 32763 29894
rect 33418 29830 33482 29894
rect 34137 29830 34201 29894
rect 34856 29830 34920 29894
rect 35575 29830 35639 29894
rect 36294 29830 36358 29894
rect 37013 29830 37077 29894
rect 30542 29750 30606 29814
rect 31261 29750 31325 29814
rect 31980 29750 32044 29814
rect 32699 29750 32763 29814
rect 33418 29750 33482 29814
rect 34137 29750 34201 29814
rect 34856 29750 34920 29814
rect 35575 29750 35639 29814
rect 36294 29750 36358 29814
rect 37013 29750 37077 29814
rect 30542 29670 30606 29734
rect 31261 29670 31325 29734
rect 31980 29670 32044 29734
rect 32699 29670 32763 29734
rect 33418 29670 33482 29734
rect 34137 29670 34201 29734
rect 34856 29670 34920 29734
rect 35575 29670 35639 29734
rect 36294 29670 36358 29734
rect 37013 29670 37077 29734
rect 30542 29590 30606 29654
rect 31261 29590 31325 29654
rect 31980 29590 32044 29654
rect 32699 29590 32763 29654
rect 33418 29590 33482 29654
rect 34137 29590 34201 29654
rect 34856 29590 34920 29654
rect 35575 29590 35639 29654
rect 36294 29590 36358 29654
rect 37013 29590 37077 29654
rect 30542 29510 30606 29574
rect 31261 29510 31325 29574
rect 31980 29510 32044 29574
rect 32699 29510 32763 29574
rect 33418 29510 33482 29574
rect 34137 29510 34201 29574
rect 34856 29510 34920 29574
rect 35575 29510 35639 29574
rect 36294 29510 36358 29574
rect 37013 29510 37077 29574
rect 30542 29430 30606 29494
rect 31261 29430 31325 29494
rect 31980 29430 32044 29494
rect 32699 29430 32763 29494
rect 33418 29430 33482 29494
rect 34137 29430 34201 29494
rect 34856 29430 34920 29494
rect 35575 29430 35639 29494
rect 36294 29430 36358 29494
rect 37013 29430 37077 29494
rect 30542 29350 30606 29414
rect 31261 29350 31325 29414
rect 31980 29350 32044 29414
rect 32699 29350 32763 29414
rect 33418 29350 33482 29414
rect 34137 29350 34201 29414
rect 34856 29350 34920 29414
rect 35575 29350 35639 29414
rect 36294 29350 36358 29414
rect 37013 29350 37077 29414
rect 30542 29130 30606 29194
rect 31261 29130 31325 29194
rect 31980 29130 32044 29194
rect 32699 29130 32763 29194
rect 33418 29130 33482 29194
rect 34137 29130 34201 29194
rect 34856 29130 34920 29194
rect 35575 29130 35639 29194
rect 36294 29130 36358 29194
rect 37013 29130 37077 29194
rect 30542 29050 30606 29114
rect 31261 29050 31325 29114
rect 31980 29050 32044 29114
rect 32699 29050 32763 29114
rect 33418 29050 33482 29114
rect 34137 29050 34201 29114
rect 34856 29050 34920 29114
rect 35575 29050 35639 29114
rect 36294 29050 36358 29114
rect 37013 29050 37077 29114
rect 30542 28970 30606 29034
rect 31261 28970 31325 29034
rect 31980 28970 32044 29034
rect 32699 28970 32763 29034
rect 33418 28970 33482 29034
rect 34137 28970 34201 29034
rect 34856 28970 34920 29034
rect 35575 28970 35639 29034
rect 36294 28970 36358 29034
rect 37013 28970 37077 29034
rect 30542 28890 30606 28954
rect 31261 28890 31325 28954
rect 31980 28890 32044 28954
rect 32699 28890 32763 28954
rect 33418 28890 33482 28954
rect 34137 28890 34201 28954
rect 34856 28890 34920 28954
rect 35575 28890 35639 28954
rect 36294 28890 36358 28954
rect 37013 28890 37077 28954
rect 30542 28810 30606 28874
rect 31261 28810 31325 28874
rect 31980 28810 32044 28874
rect 32699 28810 32763 28874
rect 33418 28810 33482 28874
rect 34137 28810 34201 28874
rect 34856 28810 34920 28874
rect 35575 28810 35639 28874
rect 36294 28810 36358 28874
rect 37013 28810 37077 28874
rect 30542 28730 30606 28794
rect 31261 28730 31325 28794
rect 31980 28730 32044 28794
rect 32699 28730 32763 28794
rect 33418 28730 33482 28794
rect 34137 28730 34201 28794
rect 34856 28730 34920 28794
rect 35575 28730 35639 28794
rect 36294 28730 36358 28794
rect 37013 28730 37077 28794
rect 30542 28650 30606 28714
rect 31261 28650 31325 28714
rect 31980 28650 32044 28714
rect 32699 28650 32763 28714
rect 33418 28650 33482 28714
rect 34137 28650 34201 28714
rect 34856 28650 34920 28714
rect 35575 28650 35639 28714
rect 36294 28650 36358 28714
rect 37013 28650 37077 28714
rect 29956 28490 30020 28494
rect 30036 28490 30100 28494
rect 29956 28434 30000 28490
rect 30000 28434 30020 28490
rect 30036 28434 30056 28490
rect 30056 28434 30100 28490
rect 29956 28430 30020 28434
rect 30036 28430 30100 28434
rect 924 28300 988 28304
rect 924 28244 928 28300
rect 928 28244 984 28300
rect 984 28244 988 28300
rect 924 28240 988 28244
rect 1004 28300 1068 28304
rect 1004 28244 1008 28300
rect 1008 28244 1064 28300
rect 1064 28244 1068 28300
rect 1004 28240 1068 28244
rect 1084 28300 1148 28304
rect 1084 28244 1088 28300
rect 1088 28244 1144 28300
rect 1144 28244 1148 28300
rect 1084 28240 1148 28244
rect 1164 28300 1228 28304
rect 1164 28244 1168 28300
rect 1168 28244 1224 28300
rect 1224 28244 1228 28300
rect 1164 28240 1228 28244
rect 1244 28300 1308 28304
rect 1244 28244 1248 28300
rect 1248 28244 1304 28300
rect 1304 28244 1308 28300
rect 1244 28240 1308 28244
rect 1324 28300 1388 28304
rect 1324 28244 1328 28300
rect 1328 28244 1384 28300
rect 1384 28244 1388 28300
rect 1324 28240 1388 28244
rect 1404 28300 1468 28304
rect 1404 28244 1408 28300
rect 1408 28244 1464 28300
rect 1464 28244 1468 28300
rect 1404 28240 1468 28244
rect 1484 28300 1548 28304
rect 1484 28244 1488 28300
rect 1488 28244 1544 28300
rect 1544 28244 1548 28300
rect 1484 28240 1548 28244
rect 1564 28300 1628 28304
rect 1564 28244 1568 28300
rect 1568 28244 1624 28300
rect 1624 28244 1628 28300
rect 1564 28240 1628 28244
rect 1644 28300 1708 28304
rect 1644 28244 1648 28300
rect 1648 28244 1704 28300
rect 1704 28244 1708 28300
rect 1644 28240 1708 28244
rect 1724 28300 1788 28304
rect 1724 28244 1728 28300
rect 1728 28244 1784 28300
rect 1784 28244 1788 28300
rect 1724 28240 1788 28244
rect 1804 28300 1868 28304
rect 1804 28244 1808 28300
rect 1808 28244 1864 28300
rect 1864 28244 1868 28300
rect 1804 28240 1868 28244
rect 1884 28300 1948 28304
rect 1884 28244 1888 28300
rect 1888 28244 1944 28300
rect 1944 28244 1948 28300
rect 1884 28240 1948 28244
rect 1964 28300 2028 28304
rect 1964 28244 1968 28300
rect 1968 28244 2024 28300
rect 2024 28244 2028 28300
rect 1964 28240 2028 28244
rect 2044 28300 2108 28304
rect 2044 28244 2048 28300
rect 2048 28244 2104 28300
rect 2104 28244 2108 28300
rect 2044 28240 2108 28244
rect 2124 28300 2188 28304
rect 2124 28244 2128 28300
rect 2128 28244 2184 28300
rect 2184 28244 2188 28300
rect 2124 28240 2188 28244
rect 2204 28300 2268 28304
rect 2204 28244 2208 28300
rect 2208 28244 2264 28300
rect 2264 28244 2268 28300
rect 2204 28240 2268 28244
rect 2284 28300 2348 28304
rect 2284 28244 2288 28300
rect 2288 28244 2344 28300
rect 2344 28244 2348 28300
rect 2284 28240 2348 28244
rect 2364 28300 2428 28304
rect 2364 28244 2368 28300
rect 2368 28244 2424 28300
rect 2424 28244 2428 28300
rect 2364 28240 2428 28244
rect 2444 28300 2508 28304
rect 2444 28244 2448 28300
rect 2448 28244 2504 28300
rect 2504 28244 2508 28300
rect 2444 28240 2508 28244
rect 55928 28300 55992 28304
rect 55928 28244 55932 28300
rect 55932 28244 55988 28300
rect 55988 28244 55992 28300
rect 55928 28240 55992 28244
rect 56008 28300 56072 28304
rect 56008 28244 56012 28300
rect 56012 28244 56068 28300
rect 56068 28244 56072 28300
rect 56008 28240 56072 28244
rect 56088 28300 56152 28304
rect 56088 28244 56092 28300
rect 56092 28244 56148 28300
rect 56148 28244 56152 28300
rect 56088 28240 56152 28244
rect 56168 28300 56232 28304
rect 56168 28244 56172 28300
rect 56172 28244 56228 28300
rect 56228 28244 56232 28300
rect 56168 28240 56232 28244
rect 56248 28300 56312 28304
rect 56248 28244 56252 28300
rect 56252 28244 56308 28300
rect 56308 28244 56312 28300
rect 56248 28240 56312 28244
rect 56328 28300 56392 28304
rect 56328 28244 56332 28300
rect 56332 28244 56388 28300
rect 56388 28244 56392 28300
rect 56328 28240 56392 28244
rect 56408 28300 56472 28304
rect 56408 28244 56412 28300
rect 56412 28244 56468 28300
rect 56468 28244 56472 28300
rect 56408 28240 56472 28244
rect 56488 28300 56552 28304
rect 56488 28244 56492 28300
rect 56492 28244 56548 28300
rect 56548 28244 56552 28300
rect 56488 28240 56552 28244
rect 56568 28300 56632 28304
rect 56568 28244 56572 28300
rect 56572 28244 56628 28300
rect 56628 28244 56632 28300
rect 56568 28240 56632 28244
rect 56648 28300 56712 28304
rect 56648 28244 56652 28300
rect 56652 28244 56708 28300
rect 56708 28244 56712 28300
rect 56648 28240 56712 28244
rect 56728 28300 56792 28304
rect 56728 28244 56732 28300
rect 56732 28244 56788 28300
rect 56788 28244 56792 28300
rect 56728 28240 56792 28244
rect 56808 28300 56872 28304
rect 56808 28244 56812 28300
rect 56812 28244 56868 28300
rect 56868 28244 56872 28300
rect 56808 28240 56872 28244
rect 56888 28300 56952 28304
rect 56888 28244 56892 28300
rect 56892 28244 56948 28300
rect 56948 28244 56952 28300
rect 56888 28240 56952 28244
rect 56968 28300 57032 28304
rect 56968 28244 56972 28300
rect 56972 28244 57028 28300
rect 57028 28244 57032 28300
rect 56968 28240 57032 28244
rect 57048 28300 57112 28304
rect 57048 28244 57052 28300
rect 57052 28244 57108 28300
rect 57108 28244 57112 28300
rect 57048 28240 57112 28244
rect 57128 28300 57192 28304
rect 57128 28244 57132 28300
rect 57132 28244 57188 28300
rect 57188 28244 57192 28300
rect 57128 28240 57192 28244
rect 57208 28300 57272 28304
rect 57208 28244 57212 28300
rect 57212 28244 57268 28300
rect 57268 28244 57272 28300
rect 57208 28240 57272 28244
rect 57288 28300 57352 28304
rect 57288 28244 57292 28300
rect 57292 28244 57348 28300
rect 57348 28244 57352 28300
rect 57288 28240 57352 28244
rect 57368 28300 57432 28304
rect 57368 28244 57372 28300
rect 57372 28244 57428 28300
rect 57428 28244 57432 28300
rect 57368 28240 57432 28244
rect 57448 28300 57512 28304
rect 57448 28244 57452 28300
rect 57452 28244 57508 28300
rect 57508 28244 57512 28300
rect 57448 28240 57512 28244
rect 3372 26420 3436 26424
rect 3372 26364 3376 26420
rect 3376 26364 3432 26420
rect 3432 26364 3436 26420
rect 3372 26360 3436 26364
rect 3452 26420 3516 26424
rect 3452 26364 3456 26420
rect 3456 26364 3512 26420
rect 3512 26364 3516 26420
rect 3452 26360 3516 26364
rect 3532 26420 3596 26424
rect 3532 26364 3536 26420
rect 3536 26364 3592 26420
rect 3592 26364 3596 26420
rect 3532 26360 3596 26364
rect 3612 26420 3676 26424
rect 3612 26364 3616 26420
rect 3616 26364 3672 26420
rect 3672 26364 3676 26420
rect 3612 26360 3676 26364
rect 3692 26420 3756 26424
rect 3692 26364 3696 26420
rect 3696 26364 3752 26420
rect 3752 26364 3756 26420
rect 3692 26360 3756 26364
rect 3772 26420 3836 26424
rect 3772 26364 3776 26420
rect 3776 26364 3832 26420
rect 3832 26364 3836 26420
rect 3772 26360 3836 26364
rect 3852 26420 3916 26424
rect 3852 26364 3856 26420
rect 3856 26364 3912 26420
rect 3912 26364 3916 26420
rect 3852 26360 3916 26364
rect 3932 26420 3996 26424
rect 3932 26364 3936 26420
rect 3936 26364 3992 26420
rect 3992 26364 3996 26420
rect 3932 26360 3996 26364
rect 4012 26420 4076 26424
rect 4012 26364 4016 26420
rect 4016 26364 4072 26420
rect 4072 26364 4076 26420
rect 4012 26360 4076 26364
rect 4092 26420 4156 26424
rect 4092 26364 4096 26420
rect 4096 26364 4152 26420
rect 4152 26364 4156 26420
rect 4092 26360 4156 26364
rect 4172 26420 4236 26424
rect 4172 26364 4176 26420
rect 4176 26364 4232 26420
rect 4232 26364 4236 26420
rect 4172 26360 4236 26364
rect 4252 26420 4316 26424
rect 4252 26364 4256 26420
rect 4256 26364 4312 26420
rect 4312 26364 4316 26420
rect 4252 26360 4316 26364
rect 4332 26420 4396 26424
rect 4332 26364 4336 26420
rect 4336 26364 4392 26420
rect 4392 26364 4396 26420
rect 4332 26360 4396 26364
rect 4412 26420 4476 26424
rect 4412 26364 4416 26420
rect 4416 26364 4472 26420
rect 4472 26364 4476 26420
rect 4412 26360 4476 26364
rect 4492 26420 4556 26424
rect 4492 26364 4496 26420
rect 4496 26364 4552 26420
rect 4552 26364 4556 26420
rect 4492 26360 4556 26364
rect 4572 26420 4636 26424
rect 4572 26364 4576 26420
rect 4576 26364 4632 26420
rect 4632 26364 4636 26420
rect 4572 26360 4636 26364
rect 4652 26420 4716 26424
rect 4652 26364 4656 26420
rect 4656 26364 4712 26420
rect 4712 26364 4716 26420
rect 4652 26360 4716 26364
rect 4732 26420 4796 26424
rect 4732 26364 4736 26420
rect 4736 26364 4792 26420
rect 4792 26364 4796 26420
rect 4732 26360 4796 26364
rect 4812 26420 4876 26424
rect 4812 26364 4816 26420
rect 4816 26364 4872 26420
rect 4872 26364 4876 26420
rect 4812 26360 4876 26364
rect 4892 26420 4956 26424
rect 4892 26364 4896 26420
rect 4896 26364 4952 26420
rect 4952 26364 4956 26420
rect 4892 26360 4956 26364
rect 33410 26392 33474 26396
rect 33410 26336 33414 26392
rect 33414 26336 33470 26392
rect 33470 26336 33474 26392
rect 33410 26332 33474 26336
rect 53480 26420 53544 26424
rect 53480 26364 53484 26420
rect 53484 26364 53540 26420
rect 53540 26364 53544 26420
rect 53480 26360 53544 26364
rect 53560 26420 53624 26424
rect 53560 26364 53564 26420
rect 53564 26364 53620 26420
rect 53620 26364 53624 26420
rect 53560 26360 53624 26364
rect 53640 26420 53704 26424
rect 53640 26364 53644 26420
rect 53644 26364 53700 26420
rect 53700 26364 53704 26420
rect 53640 26360 53704 26364
rect 53720 26420 53784 26424
rect 53720 26364 53724 26420
rect 53724 26364 53780 26420
rect 53780 26364 53784 26420
rect 53720 26360 53784 26364
rect 53800 26420 53864 26424
rect 53800 26364 53804 26420
rect 53804 26364 53860 26420
rect 53860 26364 53864 26420
rect 53800 26360 53864 26364
rect 53880 26420 53944 26424
rect 53880 26364 53884 26420
rect 53884 26364 53940 26420
rect 53940 26364 53944 26420
rect 53880 26360 53944 26364
rect 53960 26420 54024 26424
rect 53960 26364 53964 26420
rect 53964 26364 54020 26420
rect 54020 26364 54024 26420
rect 53960 26360 54024 26364
rect 54040 26420 54104 26424
rect 54040 26364 54044 26420
rect 54044 26364 54100 26420
rect 54100 26364 54104 26420
rect 54040 26360 54104 26364
rect 54120 26420 54184 26424
rect 54120 26364 54124 26420
rect 54124 26364 54180 26420
rect 54180 26364 54184 26420
rect 54120 26360 54184 26364
rect 54200 26420 54264 26424
rect 54200 26364 54204 26420
rect 54204 26364 54260 26420
rect 54260 26364 54264 26420
rect 54200 26360 54264 26364
rect 54280 26420 54344 26424
rect 54280 26364 54284 26420
rect 54284 26364 54340 26420
rect 54340 26364 54344 26420
rect 54280 26360 54344 26364
rect 54360 26420 54424 26424
rect 54360 26364 54364 26420
rect 54364 26364 54420 26420
rect 54420 26364 54424 26420
rect 54360 26360 54424 26364
rect 54440 26420 54504 26424
rect 54440 26364 54444 26420
rect 54444 26364 54500 26420
rect 54500 26364 54504 26420
rect 54440 26360 54504 26364
rect 54520 26420 54584 26424
rect 54520 26364 54524 26420
rect 54524 26364 54580 26420
rect 54580 26364 54584 26420
rect 54520 26360 54584 26364
rect 54600 26420 54664 26424
rect 54600 26364 54604 26420
rect 54604 26364 54660 26420
rect 54660 26364 54664 26420
rect 54600 26360 54664 26364
rect 54680 26420 54744 26424
rect 54680 26364 54684 26420
rect 54684 26364 54740 26420
rect 54740 26364 54744 26420
rect 54680 26360 54744 26364
rect 54760 26420 54824 26424
rect 54760 26364 54764 26420
rect 54764 26364 54820 26420
rect 54820 26364 54824 26420
rect 54760 26360 54824 26364
rect 54840 26420 54904 26424
rect 54840 26364 54844 26420
rect 54844 26364 54900 26420
rect 54900 26364 54904 26420
rect 54840 26360 54904 26364
rect 54920 26420 54984 26424
rect 54920 26364 54924 26420
rect 54924 26364 54980 26420
rect 54980 26364 54984 26420
rect 54920 26360 54984 26364
rect 55000 26420 55064 26424
rect 55000 26364 55004 26420
rect 55004 26364 55060 26420
rect 55060 26364 55064 26420
rect 55000 26360 55064 26364
rect 30542 26070 30606 26134
rect 31261 26070 31325 26134
rect 31980 26070 32044 26134
rect 32699 26070 32763 26134
rect 33418 26070 33482 26134
rect 34137 26070 34201 26134
rect 34856 26070 34920 26134
rect 35575 26070 35639 26134
rect 36294 26070 36358 26134
rect 37013 26070 37077 26134
rect 30542 25990 30606 26054
rect 31261 25990 31325 26054
rect 31980 25990 32044 26054
rect 32699 25990 32763 26054
rect 33418 25990 33482 26054
rect 34137 25990 34201 26054
rect 34856 25990 34920 26054
rect 35575 25990 35639 26054
rect 36294 25990 36358 26054
rect 37013 25990 37077 26054
rect 30542 25910 30606 25974
rect 31261 25910 31325 25974
rect 31980 25910 32044 25974
rect 32699 25910 32763 25974
rect 33418 25910 33482 25974
rect 34137 25910 34201 25974
rect 34856 25910 34920 25974
rect 35575 25910 35639 25974
rect 36294 25910 36358 25974
rect 37013 25910 37077 25974
rect 30542 25830 30606 25894
rect 31261 25830 31325 25894
rect 31980 25830 32044 25894
rect 32699 25830 32763 25894
rect 33418 25830 33482 25894
rect 34137 25830 34201 25894
rect 34856 25830 34920 25894
rect 35575 25830 35639 25894
rect 36294 25830 36358 25894
rect 37013 25830 37077 25894
rect 29684 25722 29748 25786
rect 30542 25750 30606 25814
rect 31261 25750 31325 25814
rect 31980 25750 32044 25814
rect 32699 25750 32763 25814
rect 33418 25750 33482 25814
rect 34137 25750 34201 25814
rect 34856 25750 34920 25814
rect 35575 25750 35639 25814
rect 36294 25750 36358 25814
rect 37013 25750 37077 25814
rect 30542 25670 30606 25734
rect 31261 25670 31325 25734
rect 31980 25670 32044 25734
rect 32699 25670 32763 25734
rect 33418 25670 33482 25734
rect 34137 25670 34201 25734
rect 34856 25670 34920 25734
rect 35575 25670 35639 25734
rect 36294 25670 36358 25734
rect 37013 25670 37077 25734
rect 30542 25590 30606 25654
rect 31261 25590 31325 25654
rect 31980 25590 32044 25654
rect 32699 25590 32763 25654
rect 33418 25590 33482 25654
rect 34137 25590 34201 25654
rect 34856 25590 34920 25654
rect 35575 25590 35639 25654
rect 36294 25590 36358 25654
rect 37013 25590 37077 25654
rect 30542 25370 30606 25434
rect 31261 25370 31325 25434
rect 31980 25370 32044 25434
rect 32699 25370 32763 25434
rect 33418 25370 33482 25434
rect 34137 25370 34201 25434
rect 34856 25370 34920 25434
rect 35575 25370 35639 25434
rect 36294 25370 36358 25434
rect 37013 25370 37077 25434
rect 30542 25290 30606 25354
rect 31261 25290 31325 25354
rect 31980 25290 32044 25354
rect 32699 25290 32763 25354
rect 33418 25290 33482 25354
rect 34137 25290 34201 25354
rect 34856 25290 34920 25354
rect 35575 25290 35639 25354
rect 36294 25290 36358 25354
rect 37013 25290 37077 25354
rect 30542 25210 30606 25274
rect 31261 25210 31325 25274
rect 31980 25210 32044 25274
rect 32699 25210 32763 25274
rect 33418 25210 33482 25274
rect 34137 25210 34201 25274
rect 34856 25210 34920 25274
rect 35575 25210 35639 25274
rect 36294 25210 36358 25274
rect 37013 25210 37077 25274
rect 30542 25130 30606 25194
rect 31261 25130 31325 25194
rect 31980 25130 32044 25194
rect 32699 25130 32763 25194
rect 33418 25130 33482 25194
rect 34137 25130 34201 25194
rect 34856 25130 34920 25194
rect 35575 25130 35639 25194
rect 36294 25130 36358 25194
rect 37013 25130 37077 25194
rect 30542 25050 30606 25114
rect 31261 25050 31325 25114
rect 31980 25050 32044 25114
rect 32699 25050 32763 25114
rect 33418 25050 33482 25114
rect 34137 25050 34201 25114
rect 34856 25050 34920 25114
rect 35575 25050 35639 25114
rect 36294 25050 36358 25114
rect 37013 25050 37077 25114
rect 30542 24970 30606 25034
rect 31261 24970 31325 25034
rect 31980 24970 32044 25034
rect 32699 24970 32763 25034
rect 33418 24970 33482 25034
rect 34137 24970 34201 25034
rect 34856 24970 34920 25034
rect 35575 24970 35639 25034
rect 36294 24970 36358 25034
rect 37013 24970 37077 25034
rect 30542 24890 30606 24954
rect 31261 24890 31325 24954
rect 31980 24890 32044 24954
rect 32699 24890 32763 24954
rect 33418 24890 33482 24954
rect 34137 24890 34201 24954
rect 34856 24890 34920 24954
rect 35575 24890 35639 24954
rect 36294 24890 36358 24954
rect 37013 24890 37077 24954
rect 29956 24730 30020 24734
rect 30036 24730 30100 24734
rect 29956 24674 30000 24730
rect 30000 24674 30020 24730
rect 30036 24674 30056 24730
rect 30056 24674 30100 24730
rect 29956 24670 30020 24674
rect 30036 24670 30100 24674
rect 924 24540 988 24544
rect 924 24484 928 24540
rect 928 24484 984 24540
rect 984 24484 988 24540
rect 924 24480 988 24484
rect 1004 24540 1068 24544
rect 1004 24484 1008 24540
rect 1008 24484 1064 24540
rect 1064 24484 1068 24540
rect 1004 24480 1068 24484
rect 1084 24540 1148 24544
rect 1084 24484 1088 24540
rect 1088 24484 1144 24540
rect 1144 24484 1148 24540
rect 1084 24480 1148 24484
rect 1164 24540 1228 24544
rect 1164 24484 1168 24540
rect 1168 24484 1224 24540
rect 1224 24484 1228 24540
rect 1164 24480 1228 24484
rect 1244 24540 1308 24544
rect 1244 24484 1248 24540
rect 1248 24484 1304 24540
rect 1304 24484 1308 24540
rect 1244 24480 1308 24484
rect 1324 24540 1388 24544
rect 1324 24484 1328 24540
rect 1328 24484 1384 24540
rect 1384 24484 1388 24540
rect 1324 24480 1388 24484
rect 1404 24540 1468 24544
rect 1404 24484 1408 24540
rect 1408 24484 1464 24540
rect 1464 24484 1468 24540
rect 1404 24480 1468 24484
rect 1484 24540 1548 24544
rect 1484 24484 1488 24540
rect 1488 24484 1544 24540
rect 1544 24484 1548 24540
rect 1484 24480 1548 24484
rect 1564 24540 1628 24544
rect 1564 24484 1568 24540
rect 1568 24484 1624 24540
rect 1624 24484 1628 24540
rect 1564 24480 1628 24484
rect 1644 24540 1708 24544
rect 1644 24484 1648 24540
rect 1648 24484 1704 24540
rect 1704 24484 1708 24540
rect 1644 24480 1708 24484
rect 1724 24540 1788 24544
rect 1724 24484 1728 24540
rect 1728 24484 1784 24540
rect 1784 24484 1788 24540
rect 1724 24480 1788 24484
rect 1804 24540 1868 24544
rect 1804 24484 1808 24540
rect 1808 24484 1864 24540
rect 1864 24484 1868 24540
rect 1804 24480 1868 24484
rect 1884 24540 1948 24544
rect 1884 24484 1888 24540
rect 1888 24484 1944 24540
rect 1944 24484 1948 24540
rect 1884 24480 1948 24484
rect 1964 24540 2028 24544
rect 1964 24484 1968 24540
rect 1968 24484 2024 24540
rect 2024 24484 2028 24540
rect 1964 24480 2028 24484
rect 2044 24540 2108 24544
rect 2044 24484 2048 24540
rect 2048 24484 2104 24540
rect 2104 24484 2108 24540
rect 2044 24480 2108 24484
rect 2124 24540 2188 24544
rect 2124 24484 2128 24540
rect 2128 24484 2184 24540
rect 2184 24484 2188 24540
rect 2124 24480 2188 24484
rect 2204 24540 2268 24544
rect 2204 24484 2208 24540
rect 2208 24484 2264 24540
rect 2264 24484 2268 24540
rect 2204 24480 2268 24484
rect 2284 24540 2348 24544
rect 2284 24484 2288 24540
rect 2288 24484 2344 24540
rect 2344 24484 2348 24540
rect 2284 24480 2348 24484
rect 2364 24540 2428 24544
rect 2364 24484 2368 24540
rect 2368 24484 2424 24540
rect 2424 24484 2428 24540
rect 2364 24480 2428 24484
rect 2444 24540 2508 24544
rect 2444 24484 2448 24540
rect 2448 24484 2504 24540
rect 2504 24484 2508 24540
rect 2444 24480 2508 24484
rect 55928 24540 55992 24544
rect 55928 24484 55932 24540
rect 55932 24484 55988 24540
rect 55988 24484 55992 24540
rect 55928 24480 55992 24484
rect 56008 24540 56072 24544
rect 56008 24484 56012 24540
rect 56012 24484 56068 24540
rect 56068 24484 56072 24540
rect 56008 24480 56072 24484
rect 56088 24540 56152 24544
rect 56088 24484 56092 24540
rect 56092 24484 56148 24540
rect 56148 24484 56152 24540
rect 56088 24480 56152 24484
rect 56168 24540 56232 24544
rect 56168 24484 56172 24540
rect 56172 24484 56228 24540
rect 56228 24484 56232 24540
rect 56168 24480 56232 24484
rect 56248 24540 56312 24544
rect 56248 24484 56252 24540
rect 56252 24484 56308 24540
rect 56308 24484 56312 24540
rect 56248 24480 56312 24484
rect 56328 24540 56392 24544
rect 56328 24484 56332 24540
rect 56332 24484 56388 24540
rect 56388 24484 56392 24540
rect 56328 24480 56392 24484
rect 56408 24540 56472 24544
rect 56408 24484 56412 24540
rect 56412 24484 56468 24540
rect 56468 24484 56472 24540
rect 56408 24480 56472 24484
rect 56488 24540 56552 24544
rect 56488 24484 56492 24540
rect 56492 24484 56548 24540
rect 56548 24484 56552 24540
rect 56488 24480 56552 24484
rect 56568 24540 56632 24544
rect 56568 24484 56572 24540
rect 56572 24484 56628 24540
rect 56628 24484 56632 24540
rect 56568 24480 56632 24484
rect 56648 24540 56712 24544
rect 56648 24484 56652 24540
rect 56652 24484 56708 24540
rect 56708 24484 56712 24540
rect 56648 24480 56712 24484
rect 56728 24540 56792 24544
rect 56728 24484 56732 24540
rect 56732 24484 56788 24540
rect 56788 24484 56792 24540
rect 56728 24480 56792 24484
rect 56808 24540 56872 24544
rect 56808 24484 56812 24540
rect 56812 24484 56868 24540
rect 56868 24484 56872 24540
rect 56808 24480 56872 24484
rect 56888 24540 56952 24544
rect 56888 24484 56892 24540
rect 56892 24484 56948 24540
rect 56948 24484 56952 24540
rect 56888 24480 56952 24484
rect 56968 24540 57032 24544
rect 56968 24484 56972 24540
rect 56972 24484 57028 24540
rect 57028 24484 57032 24540
rect 56968 24480 57032 24484
rect 57048 24540 57112 24544
rect 57048 24484 57052 24540
rect 57052 24484 57108 24540
rect 57108 24484 57112 24540
rect 57048 24480 57112 24484
rect 57128 24540 57192 24544
rect 57128 24484 57132 24540
rect 57132 24484 57188 24540
rect 57188 24484 57192 24540
rect 57128 24480 57192 24484
rect 57208 24540 57272 24544
rect 57208 24484 57212 24540
rect 57212 24484 57268 24540
rect 57268 24484 57272 24540
rect 57208 24480 57272 24484
rect 57288 24540 57352 24544
rect 57288 24484 57292 24540
rect 57292 24484 57348 24540
rect 57348 24484 57352 24540
rect 57288 24480 57352 24484
rect 57368 24540 57432 24544
rect 57368 24484 57372 24540
rect 57372 24484 57428 24540
rect 57428 24484 57432 24540
rect 57368 24480 57432 24484
rect 57448 24540 57512 24544
rect 57448 24484 57452 24540
rect 57452 24484 57508 24540
rect 57508 24484 57512 24540
rect 57448 24480 57512 24484
rect 3372 22660 3436 22664
rect 3372 22604 3376 22660
rect 3376 22604 3432 22660
rect 3432 22604 3436 22660
rect 3372 22600 3436 22604
rect 3452 22660 3516 22664
rect 3452 22604 3456 22660
rect 3456 22604 3512 22660
rect 3512 22604 3516 22660
rect 3452 22600 3516 22604
rect 3532 22660 3596 22664
rect 3532 22604 3536 22660
rect 3536 22604 3592 22660
rect 3592 22604 3596 22660
rect 3532 22600 3596 22604
rect 3612 22660 3676 22664
rect 3612 22604 3616 22660
rect 3616 22604 3672 22660
rect 3672 22604 3676 22660
rect 3612 22600 3676 22604
rect 3692 22660 3756 22664
rect 3692 22604 3696 22660
rect 3696 22604 3752 22660
rect 3752 22604 3756 22660
rect 3692 22600 3756 22604
rect 3772 22660 3836 22664
rect 3772 22604 3776 22660
rect 3776 22604 3832 22660
rect 3832 22604 3836 22660
rect 3772 22600 3836 22604
rect 3852 22660 3916 22664
rect 3852 22604 3856 22660
rect 3856 22604 3912 22660
rect 3912 22604 3916 22660
rect 3852 22600 3916 22604
rect 3932 22660 3996 22664
rect 3932 22604 3936 22660
rect 3936 22604 3992 22660
rect 3992 22604 3996 22660
rect 3932 22600 3996 22604
rect 4012 22660 4076 22664
rect 4012 22604 4016 22660
rect 4016 22604 4072 22660
rect 4072 22604 4076 22660
rect 4012 22600 4076 22604
rect 4092 22660 4156 22664
rect 4092 22604 4096 22660
rect 4096 22604 4152 22660
rect 4152 22604 4156 22660
rect 4092 22600 4156 22604
rect 4172 22660 4236 22664
rect 4172 22604 4176 22660
rect 4176 22604 4232 22660
rect 4232 22604 4236 22660
rect 4172 22600 4236 22604
rect 4252 22660 4316 22664
rect 4252 22604 4256 22660
rect 4256 22604 4312 22660
rect 4312 22604 4316 22660
rect 4252 22600 4316 22604
rect 4332 22660 4396 22664
rect 4332 22604 4336 22660
rect 4336 22604 4392 22660
rect 4392 22604 4396 22660
rect 4332 22600 4396 22604
rect 4412 22660 4476 22664
rect 4412 22604 4416 22660
rect 4416 22604 4472 22660
rect 4472 22604 4476 22660
rect 4412 22600 4476 22604
rect 4492 22660 4556 22664
rect 4492 22604 4496 22660
rect 4496 22604 4552 22660
rect 4552 22604 4556 22660
rect 4492 22600 4556 22604
rect 4572 22660 4636 22664
rect 4572 22604 4576 22660
rect 4576 22604 4632 22660
rect 4632 22604 4636 22660
rect 4572 22600 4636 22604
rect 4652 22660 4716 22664
rect 4652 22604 4656 22660
rect 4656 22604 4712 22660
rect 4712 22604 4716 22660
rect 4652 22600 4716 22604
rect 4732 22660 4796 22664
rect 4732 22604 4736 22660
rect 4736 22604 4792 22660
rect 4792 22604 4796 22660
rect 4732 22600 4796 22604
rect 4812 22660 4876 22664
rect 4812 22604 4816 22660
rect 4816 22604 4872 22660
rect 4872 22604 4876 22660
rect 4812 22600 4876 22604
rect 4892 22660 4956 22664
rect 4892 22604 4896 22660
rect 4896 22604 4952 22660
rect 4952 22604 4956 22660
rect 4892 22600 4956 22604
rect 53480 22660 53544 22664
rect 53480 22604 53484 22660
rect 53484 22604 53540 22660
rect 53540 22604 53544 22660
rect 53480 22600 53544 22604
rect 53560 22660 53624 22664
rect 53560 22604 53564 22660
rect 53564 22604 53620 22660
rect 53620 22604 53624 22660
rect 53560 22600 53624 22604
rect 53640 22660 53704 22664
rect 53640 22604 53644 22660
rect 53644 22604 53700 22660
rect 53700 22604 53704 22660
rect 53640 22600 53704 22604
rect 53720 22660 53784 22664
rect 53720 22604 53724 22660
rect 53724 22604 53780 22660
rect 53780 22604 53784 22660
rect 53720 22600 53784 22604
rect 53800 22660 53864 22664
rect 53800 22604 53804 22660
rect 53804 22604 53860 22660
rect 53860 22604 53864 22660
rect 53800 22600 53864 22604
rect 53880 22660 53944 22664
rect 53880 22604 53884 22660
rect 53884 22604 53940 22660
rect 53940 22604 53944 22660
rect 53880 22600 53944 22604
rect 53960 22660 54024 22664
rect 53960 22604 53964 22660
rect 53964 22604 54020 22660
rect 54020 22604 54024 22660
rect 53960 22600 54024 22604
rect 54040 22660 54104 22664
rect 54040 22604 54044 22660
rect 54044 22604 54100 22660
rect 54100 22604 54104 22660
rect 54040 22600 54104 22604
rect 54120 22660 54184 22664
rect 54120 22604 54124 22660
rect 54124 22604 54180 22660
rect 54180 22604 54184 22660
rect 54120 22600 54184 22604
rect 54200 22660 54264 22664
rect 54200 22604 54204 22660
rect 54204 22604 54260 22660
rect 54260 22604 54264 22660
rect 54200 22600 54264 22604
rect 54280 22660 54344 22664
rect 54280 22604 54284 22660
rect 54284 22604 54340 22660
rect 54340 22604 54344 22660
rect 54280 22600 54344 22604
rect 54360 22660 54424 22664
rect 54360 22604 54364 22660
rect 54364 22604 54420 22660
rect 54420 22604 54424 22660
rect 54360 22600 54424 22604
rect 54440 22660 54504 22664
rect 54440 22604 54444 22660
rect 54444 22604 54500 22660
rect 54500 22604 54504 22660
rect 54440 22600 54504 22604
rect 54520 22660 54584 22664
rect 54520 22604 54524 22660
rect 54524 22604 54580 22660
rect 54580 22604 54584 22660
rect 54520 22600 54584 22604
rect 54600 22660 54664 22664
rect 54600 22604 54604 22660
rect 54604 22604 54660 22660
rect 54660 22604 54664 22660
rect 54600 22600 54664 22604
rect 54680 22660 54744 22664
rect 54680 22604 54684 22660
rect 54684 22604 54740 22660
rect 54740 22604 54744 22660
rect 54680 22600 54744 22604
rect 54760 22660 54824 22664
rect 54760 22604 54764 22660
rect 54764 22604 54820 22660
rect 54820 22604 54824 22660
rect 54760 22600 54824 22604
rect 54840 22660 54904 22664
rect 54840 22604 54844 22660
rect 54844 22604 54900 22660
rect 54900 22604 54904 22660
rect 54840 22600 54904 22604
rect 54920 22660 54984 22664
rect 54920 22604 54924 22660
rect 54924 22604 54980 22660
rect 54980 22604 54984 22660
rect 54920 22600 54984 22604
rect 55000 22660 55064 22664
rect 55000 22604 55004 22660
rect 55004 22604 55060 22660
rect 55060 22604 55064 22660
rect 55000 22600 55064 22604
rect 924 20780 988 20784
rect 924 20724 928 20780
rect 928 20724 984 20780
rect 984 20724 988 20780
rect 924 20720 988 20724
rect 1004 20780 1068 20784
rect 1004 20724 1008 20780
rect 1008 20724 1064 20780
rect 1064 20724 1068 20780
rect 1004 20720 1068 20724
rect 1084 20780 1148 20784
rect 1084 20724 1088 20780
rect 1088 20724 1144 20780
rect 1144 20724 1148 20780
rect 1084 20720 1148 20724
rect 1164 20780 1228 20784
rect 1164 20724 1168 20780
rect 1168 20724 1224 20780
rect 1224 20724 1228 20780
rect 1164 20720 1228 20724
rect 1244 20780 1308 20784
rect 1244 20724 1248 20780
rect 1248 20724 1304 20780
rect 1304 20724 1308 20780
rect 1244 20720 1308 20724
rect 1324 20780 1388 20784
rect 1324 20724 1328 20780
rect 1328 20724 1384 20780
rect 1384 20724 1388 20780
rect 1324 20720 1388 20724
rect 1404 20780 1468 20784
rect 1404 20724 1408 20780
rect 1408 20724 1464 20780
rect 1464 20724 1468 20780
rect 1404 20720 1468 20724
rect 1484 20780 1548 20784
rect 1484 20724 1488 20780
rect 1488 20724 1544 20780
rect 1544 20724 1548 20780
rect 1484 20720 1548 20724
rect 1564 20780 1628 20784
rect 1564 20724 1568 20780
rect 1568 20724 1624 20780
rect 1624 20724 1628 20780
rect 1564 20720 1628 20724
rect 1644 20780 1708 20784
rect 1644 20724 1648 20780
rect 1648 20724 1704 20780
rect 1704 20724 1708 20780
rect 1644 20720 1708 20724
rect 1724 20780 1788 20784
rect 1724 20724 1728 20780
rect 1728 20724 1784 20780
rect 1784 20724 1788 20780
rect 1724 20720 1788 20724
rect 1804 20780 1868 20784
rect 1804 20724 1808 20780
rect 1808 20724 1864 20780
rect 1864 20724 1868 20780
rect 1804 20720 1868 20724
rect 1884 20780 1948 20784
rect 1884 20724 1888 20780
rect 1888 20724 1944 20780
rect 1944 20724 1948 20780
rect 1884 20720 1948 20724
rect 1964 20780 2028 20784
rect 1964 20724 1968 20780
rect 1968 20724 2024 20780
rect 2024 20724 2028 20780
rect 1964 20720 2028 20724
rect 2044 20780 2108 20784
rect 2044 20724 2048 20780
rect 2048 20724 2104 20780
rect 2104 20724 2108 20780
rect 2044 20720 2108 20724
rect 2124 20780 2188 20784
rect 2124 20724 2128 20780
rect 2128 20724 2184 20780
rect 2184 20724 2188 20780
rect 2124 20720 2188 20724
rect 2204 20780 2268 20784
rect 2204 20724 2208 20780
rect 2208 20724 2264 20780
rect 2264 20724 2268 20780
rect 2204 20720 2268 20724
rect 2284 20780 2348 20784
rect 2284 20724 2288 20780
rect 2288 20724 2344 20780
rect 2344 20724 2348 20780
rect 2284 20720 2348 20724
rect 2364 20780 2428 20784
rect 2364 20724 2368 20780
rect 2368 20724 2424 20780
rect 2424 20724 2428 20780
rect 2364 20720 2428 20724
rect 2444 20780 2508 20784
rect 2444 20724 2448 20780
rect 2448 20724 2504 20780
rect 2504 20724 2508 20780
rect 2444 20720 2508 20724
rect 55928 20780 55992 20784
rect 55928 20724 55932 20780
rect 55932 20724 55988 20780
rect 55988 20724 55992 20780
rect 55928 20720 55992 20724
rect 56008 20780 56072 20784
rect 56008 20724 56012 20780
rect 56012 20724 56068 20780
rect 56068 20724 56072 20780
rect 56008 20720 56072 20724
rect 56088 20780 56152 20784
rect 56088 20724 56092 20780
rect 56092 20724 56148 20780
rect 56148 20724 56152 20780
rect 56088 20720 56152 20724
rect 56168 20780 56232 20784
rect 56168 20724 56172 20780
rect 56172 20724 56228 20780
rect 56228 20724 56232 20780
rect 56168 20720 56232 20724
rect 56248 20780 56312 20784
rect 56248 20724 56252 20780
rect 56252 20724 56308 20780
rect 56308 20724 56312 20780
rect 56248 20720 56312 20724
rect 56328 20780 56392 20784
rect 56328 20724 56332 20780
rect 56332 20724 56388 20780
rect 56388 20724 56392 20780
rect 56328 20720 56392 20724
rect 56408 20780 56472 20784
rect 56408 20724 56412 20780
rect 56412 20724 56468 20780
rect 56468 20724 56472 20780
rect 56408 20720 56472 20724
rect 56488 20780 56552 20784
rect 56488 20724 56492 20780
rect 56492 20724 56548 20780
rect 56548 20724 56552 20780
rect 56488 20720 56552 20724
rect 56568 20780 56632 20784
rect 56568 20724 56572 20780
rect 56572 20724 56628 20780
rect 56628 20724 56632 20780
rect 56568 20720 56632 20724
rect 56648 20780 56712 20784
rect 56648 20724 56652 20780
rect 56652 20724 56708 20780
rect 56708 20724 56712 20780
rect 56648 20720 56712 20724
rect 56728 20780 56792 20784
rect 56728 20724 56732 20780
rect 56732 20724 56788 20780
rect 56788 20724 56792 20780
rect 56728 20720 56792 20724
rect 56808 20780 56872 20784
rect 56808 20724 56812 20780
rect 56812 20724 56868 20780
rect 56868 20724 56872 20780
rect 56808 20720 56872 20724
rect 56888 20780 56952 20784
rect 56888 20724 56892 20780
rect 56892 20724 56948 20780
rect 56948 20724 56952 20780
rect 56888 20720 56952 20724
rect 56968 20780 57032 20784
rect 56968 20724 56972 20780
rect 56972 20724 57028 20780
rect 57028 20724 57032 20780
rect 56968 20720 57032 20724
rect 57048 20780 57112 20784
rect 57048 20724 57052 20780
rect 57052 20724 57108 20780
rect 57108 20724 57112 20780
rect 57048 20720 57112 20724
rect 57128 20780 57192 20784
rect 57128 20724 57132 20780
rect 57132 20724 57188 20780
rect 57188 20724 57192 20780
rect 57128 20720 57192 20724
rect 57208 20780 57272 20784
rect 57208 20724 57212 20780
rect 57212 20724 57268 20780
rect 57268 20724 57272 20780
rect 57208 20720 57272 20724
rect 57288 20780 57352 20784
rect 57288 20724 57292 20780
rect 57292 20724 57348 20780
rect 57348 20724 57352 20780
rect 57288 20720 57352 20724
rect 57368 20780 57432 20784
rect 57368 20724 57372 20780
rect 57372 20724 57428 20780
rect 57428 20724 57432 20780
rect 57368 20720 57432 20724
rect 57448 20780 57512 20784
rect 57448 20724 57452 20780
rect 57452 20724 57508 20780
rect 57508 20724 57512 20780
rect 57448 20720 57512 20724
rect 3372 18900 3436 18904
rect 3372 18844 3376 18900
rect 3376 18844 3432 18900
rect 3432 18844 3436 18900
rect 3372 18840 3436 18844
rect 3452 18900 3516 18904
rect 3452 18844 3456 18900
rect 3456 18844 3512 18900
rect 3512 18844 3516 18900
rect 3452 18840 3516 18844
rect 3532 18900 3596 18904
rect 3532 18844 3536 18900
rect 3536 18844 3592 18900
rect 3592 18844 3596 18900
rect 3532 18840 3596 18844
rect 3612 18900 3676 18904
rect 3612 18844 3616 18900
rect 3616 18844 3672 18900
rect 3672 18844 3676 18900
rect 3612 18840 3676 18844
rect 3692 18900 3756 18904
rect 3692 18844 3696 18900
rect 3696 18844 3752 18900
rect 3752 18844 3756 18900
rect 3692 18840 3756 18844
rect 3772 18900 3836 18904
rect 3772 18844 3776 18900
rect 3776 18844 3832 18900
rect 3832 18844 3836 18900
rect 3772 18840 3836 18844
rect 3852 18900 3916 18904
rect 3852 18844 3856 18900
rect 3856 18844 3912 18900
rect 3912 18844 3916 18900
rect 3852 18840 3916 18844
rect 3932 18900 3996 18904
rect 3932 18844 3936 18900
rect 3936 18844 3992 18900
rect 3992 18844 3996 18900
rect 3932 18840 3996 18844
rect 4012 18900 4076 18904
rect 4012 18844 4016 18900
rect 4016 18844 4072 18900
rect 4072 18844 4076 18900
rect 4012 18840 4076 18844
rect 4092 18900 4156 18904
rect 4092 18844 4096 18900
rect 4096 18844 4152 18900
rect 4152 18844 4156 18900
rect 4092 18840 4156 18844
rect 4172 18900 4236 18904
rect 4172 18844 4176 18900
rect 4176 18844 4232 18900
rect 4232 18844 4236 18900
rect 4172 18840 4236 18844
rect 4252 18900 4316 18904
rect 4252 18844 4256 18900
rect 4256 18844 4312 18900
rect 4312 18844 4316 18900
rect 4252 18840 4316 18844
rect 4332 18900 4396 18904
rect 4332 18844 4336 18900
rect 4336 18844 4392 18900
rect 4392 18844 4396 18900
rect 4332 18840 4396 18844
rect 4412 18900 4476 18904
rect 4412 18844 4416 18900
rect 4416 18844 4472 18900
rect 4472 18844 4476 18900
rect 4412 18840 4476 18844
rect 4492 18900 4556 18904
rect 4492 18844 4496 18900
rect 4496 18844 4552 18900
rect 4552 18844 4556 18900
rect 4492 18840 4556 18844
rect 4572 18900 4636 18904
rect 4572 18844 4576 18900
rect 4576 18844 4632 18900
rect 4632 18844 4636 18900
rect 4572 18840 4636 18844
rect 4652 18900 4716 18904
rect 4652 18844 4656 18900
rect 4656 18844 4712 18900
rect 4712 18844 4716 18900
rect 4652 18840 4716 18844
rect 4732 18900 4796 18904
rect 4732 18844 4736 18900
rect 4736 18844 4792 18900
rect 4792 18844 4796 18900
rect 4732 18840 4796 18844
rect 4812 18900 4876 18904
rect 4812 18844 4816 18900
rect 4816 18844 4872 18900
rect 4872 18844 4876 18900
rect 4812 18840 4876 18844
rect 4892 18900 4956 18904
rect 4892 18844 4896 18900
rect 4896 18844 4952 18900
rect 4952 18844 4956 18900
rect 4892 18840 4956 18844
rect 53480 18900 53544 18904
rect 53480 18844 53484 18900
rect 53484 18844 53540 18900
rect 53540 18844 53544 18900
rect 53480 18840 53544 18844
rect 53560 18900 53624 18904
rect 53560 18844 53564 18900
rect 53564 18844 53620 18900
rect 53620 18844 53624 18900
rect 53560 18840 53624 18844
rect 53640 18900 53704 18904
rect 53640 18844 53644 18900
rect 53644 18844 53700 18900
rect 53700 18844 53704 18900
rect 53640 18840 53704 18844
rect 53720 18900 53784 18904
rect 53720 18844 53724 18900
rect 53724 18844 53780 18900
rect 53780 18844 53784 18900
rect 53720 18840 53784 18844
rect 53800 18900 53864 18904
rect 53800 18844 53804 18900
rect 53804 18844 53860 18900
rect 53860 18844 53864 18900
rect 53800 18840 53864 18844
rect 53880 18900 53944 18904
rect 53880 18844 53884 18900
rect 53884 18844 53940 18900
rect 53940 18844 53944 18900
rect 53880 18840 53944 18844
rect 53960 18900 54024 18904
rect 53960 18844 53964 18900
rect 53964 18844 54020 18900
rect 54020 18844 54024 18900
rect 53960 18840 54024 18844
rect 54040 18900 54104 18904
rect 54040 18844 54044 18900
rect 54044 18844 54100 18900
rect 54100 18844 54104 18900
rect 54040 18840 54104 18844
rect 54120 18900 54184 18904
rect 54120 18844 54124 18900
rect 54124 18844 54180 18900
rect 54180 18844 54184 18900
rect 54120 18840 54184 18844
rect 54200 18900 54264 18904
rect 54200 18844 54204 18900
rect 54204 18844 54260 18900
rect 54260 18844 54264 18900
rect 54200 18840 54264 18844
rect 54280 18900 54344 18904
rect 54280 18844 54284 18900
rect 54284 18844 54340 18900
rect 54340 18844 54344 18900
rect 54280 18840 54344 18844
rect 54360 18900 54424 18904
rect 54360 18844 54364 18900
rect 54364 18844 54420 18900
rect 54420 18844 54424 18900
rect 54360 18840 54424 18844
rect 54440 18900 54504 18904
rect 54440 18844 54444 18900
rect 54444 18844 54500 18900
rect 54500 18844 54504 18900
rect 54440 18840 54504 18844
rect 54520 18900 54584 18904
rect 54520 18844 54524 18900
rect 54524 18844 54580 18900
rect 54580 18844 54584 18900
rect 54520 18840 54584 18844
rect 54600 18900 54664 18904
rect 54600 18844 54604 18900
rect 54604 18844 54660 18900
rect 54660 18844 54664 18900
rect 54600 18840 54664 18844
rect 54680 18900 54744 18904
rect 54680 18844 54684 18900
rect 54684 18844 54740 18900
rect 54740 18844 54744 18900
rect 54680 18840 54744 18844
rect 54760 18900 54824 18904
rect 54760 18844 54764 18900
rect 54764 18844 54820 18900
rect 54820 18844 54824 18900
rect 54760 18840 54824 18844
rect 54840 18900 54904 18904
rect 54840 18844 54844 18900
rect 54844 18844 54900 18900
rect 54900 18844 54904 18900
rect 54840 18840 54904 18844
rect 54920 18900 54984 18904
rect 54920 18844 54924 18900
rect 54924 18844 54980 18900
rect 54980 18844 54984 18900
rect 54920 18840 54984 18844
rect 55000 18900 55064 18904
rect 55000 18844 55004 18900
rect 55004 18844 55060 18900
rect 55060 18844 55064 18900
rect 55000 18840 55064 18844
rect 924 17020 988 17024
rect 924 16964 928 17020
rect 928 16964 984 17020
rect 984 16964 988 17020
rect 924 16960 988 16964
rect 1004 17020 1068 17024
rect 1004 16964 1008 17020
rect 1008 16964 1064 17020
rect 1064 16964 1068 17020
rect 1004 16960 1068 16964
rect 1084 17020 1148 17024
rect 1084 16964 1088 17020
rect 1088 16964 1144 17020
rect 1144 16964 1148 17020
rect 1084 16960 1148 16964
rect 1164 17020 1228 17024
rect 1164 16964 1168 17020
rect 1168 16964 1224 17020
rect 1224 16964 1228 17020
rect 1164 16960 1228 16964
rect 1244 17020 1308 17024
rect 1244 16964 1248 17020
rect 1248 16964 1304 17020
rect 1304 16964 1308 17020
rect 1244 16960 1308 16964
rect 1324 17020 1388 17024
rect 1324 16964 1328 17020
rect 1328 16964 1384 17020
rect 1384 16964 1388 17020
rect 1324 16960 1388 16964
rect 1404 17020 1468 17024
rect 1404 16964 1408 17020
rect 1408 16964 1464 17020
rect 1464 16964 1468 17020
rect 1404 16960 1468 16964
rect 1484 17020 1548 17024
rect 1484 16964 1488 17020
rect 1488 16964 1544 17020
rect 1544 16964 1548 17020
rect 1484 16960 1548 16964
rect 1564 17020 1628 17024
rect 1564 16964 1568 17020
rect 1568 16964 1624 17020
rect 1624 16964 1628 17020
rect 1564 16960 1628 16964
rect 1644 17020 1708 17024
rect 1644 16964 1648 17020
rect 1648 16964 1704 17020
rect 1704 16964 1708 17020
rect 1644 16960 1708 16964
rect 1724 17020 1788 17024
rect 1724 16964 1728 17020
rect 1728 16964 1784 17020
rect 1784 16964 1788 17020
rect 1724 16960 1788 16964
rect 1804 17020 1868 17024
rect 1804 16964 1808 17020
rect 1808 16964 1864 17020
rect 1864 16964 1868 17020
rect 1804 16960 1868 16964
rect 1884 17020 1948 17024
rect 1884 16964 1888 17020
rect 1888 16964 1944 17020
rect 1944 16964 1948 17020
rect 1884 16960 1948 16964
rect 1964 17020 2028 17024
rect 1964 16964 1968 17020
rect 1968 16964 2024 17020
rect 2024 16964 2028 17020
rect 1964 16960 2028 16964
rect 2044 17020 2108 17024
rect 2044 16964 2048 17020
rect 2048 16964 2104 17020
rect 2104 16964 2108 17020
rect 2044 16960 2108 16964
rect 2124 17020 2188 17024
rect 2124 16964 2128 17020
rect 2128 16964 2184 17020
rect 2184 16964 2188 17020
rect 2124 16960 2188 16964
rect 2204 17020 2268 17024
rect 2204 16964 2208 17020
rect 2208 16964 2264 17020
rect 2264 16964 2268 17020
rect 2204 16960 2268 16964
rect 2284 17020 2348 17024
rect 2284 16964 2288 17020
rect 2288 16964 2344 17020
rect 2344 16964 2348 17020
rect 2284 16960 2348 16964
rect 2364 17020 2428 17024
rect 2364 16964 2368 17020
rect 2368 16964 2424 17020
rect 2424 16964 2428 17020
rect 2364 16960 2428 16964
rect 2444 17020 2508 17024
rect 2444 16964 2448 17020
rect 2448 16964 2504 17020
rect 2504 16964 2508 17020
rect 2444 16960 2508 16964
rect 55928 17020 55992 17024
rect 55928 16964 55932 17020
rect 55932 16964 55988 17020
rect 55988 16964 55992 17020
rect 55928 16960 55992 16964
rect 56008 17020 56072 17024
rect 56008 16964 56012 17020
rect 56012 16964 56068 17020
rect 56068 16964 56072 17020
rect 56008 16960 56072 16964
rect 56088 17020 56152 17024
rect 56088 16964 56092 17020
rect 56092 16964 56148 17020
rect 56148 16964 56152 17020
rect 56088 16960 56152 16964
rect 56168 17020 56232 17024
rect 56168 16964 56172 17020
rect 56172 16964 56228 17020
rect 56228 16964 56232 17020
rect 56168 16960 56232 16964
rect 56248 17020 56312 17024
rect 56248 16964 56252 17020
rect 56252 16964 56308 17020
rect 56308 16964 56312 17020
rect 56248 16960 56312 16964
rect 56328 17020 56392 17024
rect 56328 16964 56332 17020
rect 56332 16964 56388 17020
rect 56388 16964 56392 17020
rect 56328 16960 56392 16964
rect 56408 17020 56472 17024
rect 56408 16964 56412 17020
rect 56412 16964 56468 17020
rect 56468 16964 56472 17020
rect 56408 16960 56472 16964
rect 56488 17020 56552 17024
rect 56488 16964 56492 17020
rect 56492 16964 56548 17020
rect 56548 16964 56552 17020
rect 56488 16960 56552 16964
rect 56568 17020 56632 17024
rect 56568 16964 56572 17020
rect 56572 16964 56628 17020
rect 56628 16964 56632 17020
rect 56568 16960 56632 16964
rect 56648 17020 56712 17024
rect 56648 16964 56652 17020
rect 56652 16964 56708 17020
rect 56708 16964 56712 17020
rect 56648 16960 56712 16964
rect 56728 17020 56792 17024
rect 56728 16964 56732 17020
rect 56732 16964 56788 17020
rect 56788 16964 56792 17020
rect 56728 16960 56792 16964
rect 56808 17020 56872 17024
rect 56808 16964 56812 17020
rect 56812 16964 56868 17020
rect 56868 16964 56872 17020
rect 56808 16960 56872 16964
rect 56888 17020 56952 17024
rect 56888 16964 56892 17020
rect 56892 16964 56948 17020
rect 56948 16964 56952 17020
rect 56888 16960 56952 16964
rect 56968 17020 57032 17024
rect 56968 16964 56972 17020
rect 56972 16964 57028 17020
rect 57028 16964 57032 17020
rect 56968 16960 57032 16964
rect 57048 17020 57112 17024
rect 57048 16964 57052 17020
rect 57052 16964 57108 17020
rect 57108 16964 57112 17020
rect 57048 16960 57112 16964
rect 57128 17020 57192 17024
rect 57128 16964 57132 17020
rect 57132 16964 57188 17020
rect 57188 16964 57192 17020
rect 57128 16960 57192 16964
rect 57208 17020 57272 17024
rect 57208 16964 57212 17020
rect 57212 16964 57268 17020
rect 57268 16964 57272 17020
rect 57208 16960 57272 16964
rect 57288 17020 57352 17024
rect 57288 16964 57292 17020
rect 57292 16964 57348 17020
rect 57348 16964 57352 17020
rect 57288 16960 57352 16964
rect 57368 17020 57432 17024
rect 57368 16964 57372 17020
rect 57372 16964 57428 17020
rect 57428 16964 57432 17020
rect 57368 16960 57432 16964
rect 57448 17020 57512 17024
rect 57448 16964 57452 17020
rect 57452 16964 57508 17020
rect 57508 16964 57512 17020
rect 57448 16960 57512 16964
rect 3372 15140 3436 15144
rect 3372 15084 3376 15140
rect 3376 15084 3432 15140
rect 3432 15084 3436 15140
rect 3372 15080 3436 15084
rect 3452 15140 3516 15144
rect 3452 15084 3456 15140
rect 3456 15084 3512 15140
rect 3512 15084 3516 15140
rect 3452 15080 3516 15084
rect 3532 15140 3596 15144
rect 3532 15084 3536 15140
rect 3536 15084 3592 15140
rect 3592 15084 3596 15140
rect 3532 15080 3596 15084
rect 3612 15140 3676 15144
rect 3612 15084 3616 15140
rect 3616 15084 3672 15140
rect 3672 15084 3676 15140
rect 3612 15080 3676 15084
rect 3692 15140 3756 15144
rect 3692 15084 3696 15140
rect 3696 15084 3752 15140
rect 3752 15084 3756 15140
rect 3692 15080 3756 15084
rect 3772 15140 3836 15144
rect 3772 15084 3776 15140
rect 3776 15084 3832 15140
rect 3832 15084 3836 15140
rect 3772 15080 3836 15084
rect 3852 15140 3916 15144
rect 3852 15084 3856 15140
rect 3856 15084 3912 15140
rect 3912 15084 3916 15140
rect 3852 15080 3916 15084
rect 3932 15140 3996 15144
rect 3932 15084 3936 15140
rect 3936 15084 3992 15140
rect 3992 15084 3996 15140
rect 3932 15080 3996 15084
rect 4012 15140 4076 15144
rect 4012 15084 4016 15140
rect 4016 15084 4072 15140
rect 4072 15084 4076 15140
rect 4012 15080 4076 15084
rect 4092 15140 4156 15144
rect 4092 15084 4096 15140
rect 4096 15084 4152 15140
rect 4152 15084 4156 15140
rect 4092 15080 4156 15084
rect 4172 15140 4236 15144
rect 4172 15084 4176 15140
rect 4176 15084 4232 15140
rect 4232 15084 4236 15140
rect 4172 15080 4236 15084
rect 4252 15140 4316 15144
rect 4252 15084 4256 15140
rect 4256 15084 4312 15140
rect 4312 15084 4316 15140
rect 4252 15080 4316 15084
rect 4332 15140 4396 15144
rect 4332 15084 4336 15140
rect 4336 15084 4392 15140
rect 4392 15084 4396 15140
rect 4332 15080 4396 15084
rect 4412 15140 4476 15144
rect 4412 15084 4416 15140
rect 4416 15084 4472 15140
rect 4472 15084 4476 15140
rect 4412 15080 4476 15084
rect 4492 15140 4556 15144
rect 4492 15084 4496 15140
rect 4496 15084 4552 15140
rect 4552 15084 4556 15140
rect 4492 15080 4556 15084
rect 4572 15140 4636 15144
rect 4572 15084 4576 15140
rect 4576 15084 4632 15140
rect 4632 15084 4636 15140
rect 4572 15080 4636 15084
rect 4652 15140 4716 15144
rect 4652 15084 4656 15140
rect 4656 15084 4712 15140
rect 4712 15084 4716 15140
rect 4652 15080 4716 15084
rect 4732 15140 4796 15144
rect 4732 15084 4736 15140
rect 4736 15084 4792 15140
rect 4792 15084 4796 15140
rect 4732 15080 4796 15084
rect 4812 15140 4876 15144
rect 4812 15084 4816 15140
rect 4816 15084 4872 15140
rect 4872 15084 4876 15140
rect 4812 15080 4876 15084
rect 4892 15140 4956 15144
rect 4892 15084 4896 15140
rect 4896 15084 4952 15140
rect 4952 15084 4956 15140
rect 4892 15080 4956 15084
rect 53480 15140 53544 15144
rect 53480 15084 53484 15140
rect 53484 15084 53540 15140
rect 53540 15084 53544 15140
rect 53480 15080 53544 15084
rect 53560 15140 53624 15144
rect 53560 15084 53564 15140
rect 53564 15084 53620 15140
rect 53620 15084 53624 15140
rect 53560 15080 53624 15084
rect 53640 15140 53704 15144
rect 53640 15084 53644 15140
rect 53644 15084 53700 15140
rect 53700 15084 53704 15140
rect 53640 15080 53704 15084
rect 53720 15140 53784 15144
rect 53720 15084 53724 15140
rect 53724 15084 53780 15140
rect 53780 15084 53784 15140
rect 53720 15080 53784 15084
rect 53800 15140 53864 15144
rect 53800 15084 53804 15140
rect 53804 15084 53860 15140
rect 53860 15084 53864 15140
rect 53800 15080 53864 15084
rect 53880 15140 53944 15144
rect 53880 15084 53884 15140
rect 53884 15084 53940 15140
rect 53940 15084 53944 15140
rect 53880 15080 53944 15084
rect 53960 15140 54024 15144
rect 53960 15084 53964 15140
rect 53964 15084 54020 15140
rect 54020 15084 54024 15140
rect 53960 15080 54024 15084
rect 54040 15140 54104 15144
rect 54040 15084 54044 15140
rect 54044 15084 54100 15140
rect 54100 15084 54104 15140
rect 54040 15080 54104 15084
rect 54120 15140 54184 15144
rect 54120 15084 54124 15140
rect 54124 15084 54180 15140
rect 54180 15084 54184 15140
rect 54120 15080 54184 15084
rect 54200 15140 54264 15144
rect 54200 15084 54204 15140
rect 54204 15084 54260 15140
rect 54260 15084 54264 15140
rect 54200 15080 54264 15084
rect 54280 15140 54344 15144
rect 54280 15084 54284 15140
rect 54284 15084 54340 15140
rect 54340 15084 54344 15140
rect 54280 15080 54344 15084
rect 54360 15140 54424 15144
rect 54360 15084 54364 15140
rect 54364 15084 54420 15140
rect 54420 15084 54424 15140
rect 54360 15080 54424 15084
rect 54440 15140 54504 15144
rect 54440 15084 54444 15140
rect 54444 15084 54500 15140
rect 54500 15084 54504 15140
rect 54440 15080 54504 15084
rect 54520 15140 54584 15144
rect 54520 15084 54524 15140
rect 54524 15084 54580 15140
rect 54580 15084 54584 15140
rect 54520 15080 54584 15084
rect 54600 15140 54664 15144
rect 54600 15084 54604 15140
rect 54604 15084 54660 15140
rect 54660 15084 54664 15140
rect 54600 15080 54664 15084
rect 54680 15140 54744 15144
rect 54680 15084 54684 15140
rect 54684 15084 54740 15140
rect 54740 15084 54744 15140
rect 54680 15080 54744 15084
rect 54760 15140 54824 15144
rect 54760 15084 54764 15140
rect 54764 15084 54820 15140
rect 54820 15084 54824 15140
rect 54760 15080 54824 15084
rect 54840 15140 54904 15144
rect 54840 15084 54844 15140
rect 54844 15084 54900 15140
rect 54900 15084 54904 15140
rect 54840 15080 54904 15084
rect 54920 15140 54984 15144
rect 54920 15084 54924 15140
rect 54924 15084 54980 15140
rect 54980 15084 54984 15140
rect 54920 15080 54984 15084
rect 55000 15140 55064 15144
rect 55000 15084 55004 15140
rect 55004 15084 55060 15140
rect 55060 15084 55064 15140
rect 55000 15080 55064 15084
rect 924 13260 988 13264
rect 924 13204 928 13260
rect 928 13204 984 13260
rect 984 13204 988 13260
rect 924 13200 988 13204
rect 1004 13260 1068 13264
rect 1004 13204 1008 13260
rect 1008 13204 1064 13260
rect 1064 13204 1068 13260
rect 1004 13200 1068 13204
rect 1084 13260 1148 13264
rect 1084 13204 1088 13260
rect 1088 13204 1144 13260
rect 1144 13204 1148 13260
rect 1084 13200 1148 13204
rect 1164 13260 1228 13264
rect 1164 13204 1168 13260
rect 1168 13204 1224 13260
rect 1224 13204 1228 13260
rect 1164 13200 1228 13204
rect 1244 13260 1308 13264
rect 1244 13204 1248 13260
rect 1248 13204 1304 13260
rect 1304 13204 1308 13260
rect 1244 13200 1308 13204
rect 1324 13260 1388 13264
rect 1324 13204 1328 13260
rect 1328 13204 1384 13260
rect 1384 13204 1388 13260
rect 1324 13200 1388 13204
rect 1404 13260 1468 13264
rect 1404 13204 1408 13260
rect 1408 13204 1464 13260
rect 1464 13204 1468 13260
rect 1404 13200 1468 13204
rect 1484 13260 1548 13264
rect 1484 13204 1488 13260
rect 1488 13204 1544 13260
rect 1544 13204 1548 13260
rect 1484 13200 1548 13204
rect 1564 13260 1628 13264
rect 1564 13204 1568 13260
rect 1568 13204 1624 13260
rect 1624 13204 1628 13260
rect 1564 13200 1628 13204
rect 1644 13260 1708 13264
rect 1644 13204 1648 13260
rect 1648 13204 1704 13260
rect 1704 13204 1708 13260
rect 1644 13200 1708 13204
rect 1724 13260 1788 13264
rect 1724 13204 1728 13260
rect 1728 13204 1784 13260
rect 1784 13204 1788 13260
rect 1724 13200 1788 13204
rect 1804 13260 1868 13264
rect 1804 13204 1808 13260
rect 1808 13204 1864 13260
rect 1864 13204 1868 13260
rect 1804 13200 1868 13204
rect 1884 13260 1948 13264
rect 1884 13204 1888 13260
rect 1888 13204 1944 13260
rect 1944 13204 1948 13260
rect 1884 13200 1948 13204
rect 1964 13260 2028 13264
rect 1964 13204 1968 13260
rect 1968 13204 2024 13260
rect 2024 13204 2028 13260
rect 1964 13200 2028 13204
rect 2044 13260 2108 13264
rect 2044 13204 2048 13260
rect 2048 13204 2104 13260
rect 2104 13204 2108 13260
rect 2044 13200 2108 13204
rect 2124 13260 2188 13264
rect 2124 13204 2128 13260
rect 2128 13204 2184 13260
rect 2184 13204 2188 13260
rect 2124 13200 2188 13204
rect 2204 13260 2268 13264
rect 2204 13204 2208 13260
rect 2208 13204 2264 13260
rect 2264 13204 2268 13260
rect 2204 13200 2268 13204
rect 2284 13260 2348 13264
rect 2284 13204 2288 13260
rect 2288 13204 2344 13260
rect 2344 13204 2348 13260
rect 2284 13200 2348 13204
rect 2364 13260 2428 13264
rect 2364 13204 2368 13260
rect 2368 13204 2424 13260
rect 2424 13204 2428 13260
rect 2364 13200 2428 13204
rect 2444 13260 2508 13264
rect 2444 13204 2448 13260
rect 2448 13204 2504 13260
rect 2504 13204 2508 13260
rect 2444 13200 2508 13204
rect 55928 13260 55992 13264
rect 55928 13204 55932 13260
rect 55932 13204 55988 13260
rect 55988 13204 55992 13260
rect 55928 13200 55992 13204
rect 56008 13260 56072 13264
rect 56008 13204 56012 13260
rect 56012 13204 56068 13260
rect 56068 13204 56072 13260
rect 56008 13200 56072 13204
rect 56088 13260 56152 13264
rect 56088 13204 56092 13260
rect 56092 13204 56148 13260
rect 56148 13204 56152 13260
rect 56088 13200 56152 13204
rect 56168 13260 56232 13264
rect 56168 13204 56172 13260
rect 56172 13204 56228 13260
rect 56228 13204 56232 13260
rect 56168 13200 56232 13204
rect 56248 13260 56312 13264
rect 56248 13204 56252 13260
rect 56252 13204 56308 13260
rect 56308 13204 56312 13260
rect 56248 13200 56312 13204
rect 56328 13260 56392 13264
rect 56328 13204 56332 13260
rect 56332 13204 56388 13260
rect 56388 13204 56392 13260
rect 56328 13200 56392 13204
rect 56408 13260 56472 13264
rect 56408 13204 56412 13260
rect 56412 13204 56468 13260
rect 56468 13204 56472 13260
rect 56408 13200 56472 13204
rect 56488 13260 56552 13264
rect 56488 13204 56492 13260
rect 56492 13204 56548 13260
rect 56548 13204 56552 13260
rect 56488 13200 56552 13204
rect 56568 13260 56632 13264
rect 56568 13204 56572 13260
rect 56572 13204 56628 13260
rect 56628 13204 56632 13260
rect 56568 13200 56632 13204
rect 56648 13260 56712 13264
rect 56648 13204 56652 13260
rect 56652 13204 56708 13260
rect 56708 13204 56712 13260
rect 56648 13200 56712 13204
rect 56728 13260 56792 13264
rect 56728 13204 56732 13260
rect 56732 13204 56788 13260
rect 56788 13204 56792 13260
rect 56728 13200 56792 13204
rect 56808 13260 56872 13264
rect 56808 13204 56812 13260
rect 56812 13204 56868 13260
rect 56868 13204 56872 13260
rect 56808 13200 56872 13204
rect 56888 13260 56952 13264
rect 56888 13204 56892 13260
rect 56892 13204 56948 13260
rect 56948 13204 56952 13260
rect 56888 13200 56952 13204
rect 56968 13260 57032 13264
rect 56968 13204 56972 13260
rect 56972 13204 57028 13260
rect 57028 13204 57032 13260
rect 56968 13200 57032 13204
rect 57048 13260 57112 13264
rect 57048 13204 57052 13260
rect 57052 13204 57108 13260
rect 57108 13204 57112 13260
rect 57048 13200 57112 13204
rect 57128 13260 57192 13264
rect 57128 13204 57132 13260
rect 57132 13204 57188 13260
rect 57188 13204 57192 13260
rect 57128 13200 57192 13204
rect 57208 13260 57272 13264
rect 57208 13204 57212 13260
rect 57212 13204 57268 13260
rect 57268 13204 57272 13260
rect 57208 13200 57272 13204
rect 57288 13260 57352 13264
rect 57288 13204 57292 13260
rect 57292 13204 57348 13260
rect 57348 13204 57352 13260
rect 57288 13200 57352 13204
rect 57368 13260 57432 13264
rect 57368 13204 57372 13260
rect 57372 13204 57428 13260
rect 57428 13204 57432 13260
rect 57368 13200 57432 13204
rect 57448 13260 57512 13264
rect 57448 13204 57452 13260
rect 57452 13204 57508 13260
rect 57508 13204 57512 13260
rect 57448 13200 57512 13204
rect 3372 11380 3436 11384
rect 3372 11324 3376 11380
rect 3376 11324 3432 11380
rect 3432 11324 3436 11380
rect 3372 11320 3436 11324
rect 3452 11380 3516 11384
rect 3452 11324 3456 11380
rect 3456 11324 3512 11380
rect 3512 11324 3516 11380
rect 3452 11320 3516 11324
rect 3532 11380 3596 11384
rect 3532 11324 3536 11380
rect 3536 11324 3592 11380
rect 3592 11324 3596 11380
rect 3532 11320 3596 11324
rect 3612 11380 3676 11384
rect 3612 11324 3616 11380
rect 3616 11324 3672 11380
rect 3672 11324 3676 11380
rect 3612 11320 3676 11324
rect 3692 11380 3756 11384
rect 3692 11324 3696 11380
rect 3696 11324 3752 11380
rect 3752 11324 3756 11380
rect 3692 11320 3756 11324
rect 3772 11380 3836 11384
rect 3772 11324 3776 11380
rect 3776 11324 3832 11380
rect 3832 11324 3836 11380
rect 3772 11320 3836 11324
rect 3852 11380 3916 11384
rect 3852 11324 3856 11380
rect 3856 11324 3912 11380
rect 3912 11324 3916 11380
rect 3852 11320 3916 11324
rect 3932 11380 3996 11384
rect 3932 11324 3936 11380
rect 3936 11324 3992 11380
rect 3992 11324 3996 11380
rect 3932 11320 3996 11324
rect 4012 11380 4076 11384
rect 4012 11324 4016 11380
rect 4016 11324 4072 11380
rect 4072 11324 4076 11380
rect 4012 11320 4076 11324
rect 4092 11380 4156 11384
rect 4092 11324 4096 11380
rect 4096 11324 4152 11380
rect 4152 11324 4156 11380
rect 4092 11320 4156 11324
rect 4172 11380 4236 11384
rect 4172 11324 4176 11380
rect 4176 11324 4232 11380
rect 4232 11324 4236 11380
rect 4172 11320 4236 11324
rect 4252 11380 4316 11384
rect 4252 11324 4256 11380
rect 4256 11324 4312 11380
rect 4312 11324 4316 11380
rect 4252 11320 4316 11324
rect 4332 11380 4396 11384
rect 4332 11324 4336 11380
rect 4336 11324 4392 11380
rect 4392 11324 4396 11380
rect 4332 11320 4396 11324
rect 4412 11380 4476 11384
rect 4412 11324 4416 11380
rect 4416 11324 4472 11380
rect 4472 11324 4476 11380
rect 4412 11320 4476 11324
rect 4492 11380 4556 11384
rect 4492 11324 4496 11380
rect 4496 11324 4552 11380
rect 4552 11324 4556 11380
rect 4492 11320 4556 11324
rect 4572 11380 4636 11384
rect 4572 11324 4576 11380
rect 4576 11324 4632 11380
rect 4632 11324 4636 11380
rect 4572 11320 4636 11324
rect 4652 11380 4716 11384
rect 4652 11324 4656 11380
rect 4656 11324 4712 11380
rect 4712 11324 4716 11380
rect 4652 11320 4716 11324
rect 4732 11380 4796 11384
rect 4732 11324 4736 11380
rect 4736 11324 4792 11380
rect 4792 11324 4796 11380
rect 4732 11320 4796 11324
rect 4812 11380 4876 11384
rect 4812 11324 4816 11380
rect 4816 11324 4872 11380
rect 4872 11324 4876 11380
rect 4812 11320 4876 11324
rect 4892 11380 4956 11384
rect 4892 11324 4896 11380
rect 4896 11324 4952 11380
rect 4952 11324 4956 11380
rect 4892 11320 4956 11324
rect 53480 11380 53544 11384
rect 53480 11324 53484 11380
rect 53484 11324 53540 11380
rect 53540 11324 53544 11380
rect 53480 11320 53544 11324
rect 53560 11380 53624 11384
rect 53560 11324 53564 11380
rect 53564 11324 53620 11380
rect 53620 11324 53624 11380
rect 53560 11320 53624 11324
rect 53640 11380 53704 11384
rect 53640 11324 53644 11380
rect 53644 11324 53700 11380
rect 53700 11324 53704 11380
rect 53640 11320 53704 11324
rect 53720 11380 53784 11384
rect 53720 11324 53724 11380
rect 53724 11324 53780 11380
rect 53780 11324 53784 11380
rect 53720 11320 53784 11324
rect 53800 11380 53864 11384
rect 53800 11324 53804 11380
rect 53804 11324 53860 11380
rect 53860 11324 53864 11380
rect 53800 11320 53864 11324
rect 53880 11380 53944 11384
rect 53880 11324 53884 11380
rect 53884 11324 53940 11380
rect 53940 11324 53944 11380
rect 53880 11320 53944 11324
rect 53960 11380 54024 11384
rect 53960 11324 53964 11380
rect 53964 11324 54020 11380
rect 54020 11324 54024 11380
rect 53960 11320 54024 11324
rect 54040 11380 54104 11384
rect 54040 11324 54044 11380
rect 54044 11324 54100 11380
rect 54100 11324 54104 11380
rect 54040 11320 54104 11324
rect 54120 11380 54184 11384
rect 54120 11324 54124 11380
rect 54124 11324 54180 11380
rect 54180 11324 54184 11380
rect 54120 11320 54184 11324
rect 54200 11380 54264 11384
rect 54200 11324 54204 11380
rect 54204 11324 54260 11380
rect 54260 11324 54264 11380
rect 54200 11320 54264 11324
rect 54280 11380 54344 11384
rect 54280 11324 54284 11380
rect 54284 11324 54340 11380
rect 54340 11324 54344 11380
rect 54280 11320 54344 11324
rect 54360 11380 54424 11384
rect 54360 11324 54364 11380
rect 54364 11324 54420 11380
rect 54420 11324 54424 11380
rect 54360 11320 54424 11324
rect 54440 11380 54504 11384
rect 54440 11324 54444 11380
rect 54444 11324 54500 11380
rect 54500 11324 54504 11380
rect 54440 11320 54504 11324
rect 54520 11380 54584 11384
rect 54520 11324 54524 11380
rect 54524 11324 54580 11380
rect 54580 11324 54584 11380
rect 54520 11320 54584 11324
rect 54600 11380 54664 11384
rect 54600 11324 54604 11380
rect 54604 11324 54660 11380
rect 54660 11324 54664 11380
rect 54600 11320 54664 11324
rect 54680 11380 54744 11384
rect 54680 11324 54684 11380
rect 54684 11324 54740 11380
rect 54740 11324 54744 11380
rect 54680 11320 54744 11324
rect 54760 11380 54824 11384
rect 54760 11324 54764 11380
rect 54764 11324 54820 11380
rect 54820 11324 54824 11380
rect 54760 11320 54824 11324
rect 54840 11380 54904 11384
rect 54840 11324 54844 11380
rect 54844 11324 54900 11380
rect 54900 11324 54904 11380
rect 54840 11320 54904 11324
rect 54920 11380 54984 11384
rect 54920 11324 54924 11380
rect 54924 11324 54980 11380
rect 54980 11324 54984 11380
rect 54920 11320 54984 11324
rect 55000 11380 55064 11384
rect 55000 11324 55004 11380
rect 55004 11324 55060 11380
rect 55060 11324 55064 11380
rect 55000 11320 55064 11324
rect 924 9500 988 9504
rect 924 9444 928 9500
rect 928 9444 984 9500
rect 984 9444 988 9500
rect 924 9440 988 9444
rect 1004 9500 1068 9504
rect 1004 9444 1008 9500
rect 1008 9444 1064 9500
rect 1064 9444 1068 9500
rect 1004 9440 1068 9444
rect 1084 9500 1148 9504
rect 1084 9444 1088 9500
rect 1088 9444 1144 9500
rect 1144 9444 1148 9500
rect 1084 9440 1148 9444
rect 1164 9500 1228 9504
rect 1164 9444 1168 9500
rect 1168 9444 1224 9500
rect 1224 9444 1228 9500
rect 1164 9440 1228 9444
rect 1244 9500 1308 9504
rect 1244 9444 1248 9500
rect 1248 9444 1304 9500
rect 1304 9444 1308 9500
rect 1244 9440 1308 9444
rect 1324 9500 1388 9504
rect 1324 9444 1328 9500
rect 1328 9444 1384 9500
rect 1384 9444 1388 9500
rect 1324 9440 1388 9444
rect 1404 9500 1468 9504
rect 1404 9444 1408 9500
rect 1408 9444 1464 9500
rect 1464 9444 1468 9500
rect 1404 9440 1468 9444
rect 1484 9500 1548 9504
rect 1484 9444 1488 9500
rect 1488 9444 1544 9500
rect 1544 9444 1548 9500
rect 1484 9440 1548 9444
rect 1564 9500 1628 9504
rect 1564 9444 1568 9500
rect 1568 9444 1624 9500
rect 1624 9444 1628 9500
rect 1564 9440 1628 9444
rect 1644 9500 1708 9504
rect 1644 9444 1648 9500
rect 1648 9444 1704 9500
rect 1704 9444 1708 9500
rect 1644 9440 1708 9444
rect 1724 9500 1788 9504
rect 1724 9444 1728 9500
rect 1728 9444 1784 9500
rect 1784 9444 1788 9500
rect 1724 9440 1788 9444
rect 1804 9500 1868 9504
rect 1804 9444 1808 9500
rect 1808 9444 1864 9500
rect 1864 9444 1868 9500
rect 1804 9440 1868 9444
rect 1884 9500 1948 9504
rect 1884 9444 1888 9500
rect 1888 9444 1944 9500
rect 1944 9444 1948 9500
rect 1884 9440 1948 9444
rect 1964 9500 2028 9504
rect 1964 9444 1968 9500
rect 1968 9444 2024 9500
rect 2024 9444 2028 9500
rect 1964 9440 2028 9444
rect 2044 9500 2108 9504
rect 2044 9444 2048 9500
rect 2048 9444 2104 9500
rect 2104 9444 2108 9500
rect 2044 9440 2108 9444
rect 2124 9500 2188 9504
rect 2124 9444 2128 9500
rect 2128 9444 2184 9500
rect 2184 9444 2188 9500
rect 2124 9440 2188 9444
rect 2204 9500 2268 9504
rect 2204 9444 2208 9500
rect 2208 9444 2264 9500
rect 2264 9444 2268 9500
rect 2204 9440 2268 9444
rect 2284 9500 2348 9504
rect 2284 9444 2288 9500
rect 2288 9444 2344 9500
rect 2344 9444 2348 9500
rect 2284 9440 2348 9444
rect 2364 9500 2428 9504
rect 2364 9444 2368 9500
rect 2368 9444 2424 9500
rect 2424 9444 2428 9500
rect 2364 9440 2428 9444
rect 2444 9500 2508 9504
rect 2444 9444 2448 9500
rect 2448 9444 2504 9500
rect 2504 9444 2508 9500
rect 2444 9440 2508 9444
rect 55928 9500 55992 9504
rect 55928 9444 55932 9500
rect 55932 9444 55988 9500
rect 55988 9444 55992 9500
rect 55928 9440 55992 9444
rect 56008 9500 56072 9504
rect 56008 9444 56012 9500
rect 56012 9444 56068 9500
rect 56068 9444 56072 9500
rect 56008 9440 56072 9444
rect 56088 9500 56152 9504
rect 56088 9444 56092 9500
rect 56092 9444 56148 9500
rect 56148 9444 56152 9500
rect 56088 9440 56152 9444
rect 56168 9500 56232 9504
rect 56168 9444 56172 9500
rect 56172 9444 56228 9500
rect 56228 9444 56232 9500
rect 56168 9440 56232 9444
rect 56248 9500 56312 9504
rect 56248 9444 56252 9500
rect 56252 9444 56308 9500
rect 56308 9444 56312 9500
rect 56248 9440 56312 9444
rect 56328 9500 56392 9504
rect 56328 9444 56332 9500
rect 56332 9444 56388 9500
rect 56388 9444 56392 9500
rect 56328 9440 56392 9444
rect 56408 9500 56472 9504
rect 56408 9444 56412 9500
rect 56412 9444 56468 9500
rect 56468 9444 56472 9500
rect 56408 9440 56472 9444
rect 56488 9500 56552 9504
rect 56488 9444 56492 9500
rect 56492 9444 56548 9500
rect 56548 9444 56552 9500
rect 56488 9440 56552 9444
rect 56568 9500 56632 9504
rect 56568 9444 56572 9500
rect 56572 9444 56628 9500
rect 56628 9444 56632 9500
rect 56568 9440 56632 9444
rect 56648 9500 56712 9504
rect 56648 9444 56652 9500
rect 56652 9444 56708 9500
rect 56708 9444 56712 9500
rect 56648 9440 56712 9444
rect 56728 9500 56792 9504
rect 56728 9444 56732 9500
rect 56732 9444 56788 9500
rect 56788 9444 56792 9500
rect 56728 9440 56792 9444
rect 56808 9500 56872 9504
rect 56808 9444 56812 9500
rect 56812 9444 56868 9500
rect 56868 9444 56872 9500
rect 56808 9440 56872 9444
rect 56888 9500 56952 9504
rect 56888 9444 56892 9500
rect 56892 9444 56948 9500
rect 56948 9444 56952 9500
rect 56888 9440 56952 9444
rect 56968 9500 57032 9504
rect 56968 9444 56972 9500
rect 56972 9444 57028 9500
rect 57028 9444 57032 9500
rect 56968 9440 57032 9444
rect 57048 9500 57112 9504
rect 57048 9444 57052 9500
rect 57052 9444 57108 9500
rect 57108 9444 57112 9500
rect 57048 9440 57112 9444
rect 57128 9500 57192 9504
rect 57128 9444 57132 9500
rect 57132 9444 57188 9500
rect 57188 9444 57192 9500
rect 57128 9440 57192 9444
rect 57208 9500 57272 9504
rect 57208 9444 57212 9500
rect 57212 9444 57268 9500
rect 57268 9444 57272 9500
rect 57208 9440 57272 9444
rect 57288 9500 57352 9504
rect 57288 9444 57292 9500
rect 57292 9444 57348 9500
rect 57348 9444 57352 9500
rect 57288 9440 57352 9444
rect 57368 9500 57432 9504
rect 57368 9444 57372 9500
rect 57372 9444 57428 9500
rect 57428 9444 57432 9500
rect 57368 9440 57432 9444
rect 57448 9500 57512 9504
rect 57448 9444 57452 9500
rect 57452 9444 57508 9500
rect 57508 9444 57512 9500
rect 57448 9440 57512 9444
rect 3372 7620 3436 7624
rect 3372 7564 3376 7620
rect 3376 7564 3432 7620
rect 3432 7564 3436 7620
rect 3372 7560 3436 7564
rect 3452 7620 3516 7624
rect 3452 7564 3456 7620
rect 3456 7564 3512 7620
rect 3512 7564 3516 7620
rect 3452 7560 3516 7564
rect 3532 7620 3596 7624
rect 3532 7564 3536 7620
rect 3536 7564 3592 7620
rect 3592 7564 3596 7620
rect 3532 7560 3596 7564
rect 3612 7620 3676 7624
rect 3612 7564 3616 7620
rect 3616 7564 3672 7620
rect 3672 7564 3676 7620
rect 3612 7560 3676 7564
rect 3692 7620 3756 7624
rect 3692 7564 3696 7620
rect 3696 7564 3752 7620
rect 3752 7564 3756 7620
rect 3692 7560 3756 7564
rect 3772 7620 3836 7624
rect 3772 7564 3776 7620
rect 3776 7564 3832 7620
rect 3832 7564 3836 7620
rect 3772 7560 3836 7564
rect 3852 7620 3916 7624
rect 3852 7564 3856 7620
rect 3856 7564 3912 7620
rect 3912 7564 3916 7620
rect 3852 7560 3916 7564
rect 3932 7620 3996 7624
rect 3932 7564 3936 7620
rect 3936 7564 3992 7620
rect 3992 7564 3996 7620
rect 3932 7560 3996 7564
rect 4012 7620 4076 7624
rect 4012 7564 4016 7620
rect 4016 7564 4072 7620
rect 4072 7564 4076 7620
rect 4012 7560 4076 7564
rect 4092 7620 4156 7624
rect 4092 7564 4096 7620
rect 4096 7564 4152 7620
rect 4152 7564 4156 7620
rect 4092 7560 4156 7564
rect 4172 7620 4236 7624
rect 4172 7564 4176 7620
rect 4176 7564 4232 7620
rect 4232 7564 4236 7620
rect 4172 7560 4236 7564
rect 4252 7620 4316 7624
rect 4252 7564 4256 7620
rect 4256 7564 4312 7620
rect 4312 7564 4316 7620
rect 4252 7560 4316 7564
rect 4332 7620 4396 7624
rect 4332 7564 4336 7620
rect 4336 7564 4392 7620
rect 4392 7564 4396 7620
rect 4332 7560 4396 7564
rect 4412 7620 4476 7624
rect 4412 7564 4416 7620
rect 4416 7564 4472 7620
rect 4472 7564 4476 7620
rect 4412 7560 4476 7564
rect 4492 7620 4556 7624
rect 4492 7564 4496 7620
rect 4496 7564 4552 7620
rect 4552 7564 4556 7620
rect 4492 7560 4556 7564
rect 4572 7620 4636 7624
rect 4572 7564 4576 7620
rect 4576 7564 4632 7620
rect 4632 7564 4636 7620
rect 4572 7560 4636 7564
rect 4652 7620 4716 7624
rect 4652 7564 4656 7620
rect 4656 7564 4712 7620
rect 4712 7564 4716 7620
rect 4652 7560 4716 7564
rect 4732 7620 4796 7624
rect 4732 7564 4736 7620
rect 4736 7564 4792 7620
rect 4792 7564 4796 7620
rect 4732 7560 4796 7564
rect 4812 7620 4876 7624
rect 4812 7564 4816 7620
rect 4816 7564 4872 7620
rect 4872 7564 4876 7620
rect 4812 7560 4876 7564
rect 4892 7620 4956 7624
rect 4892 7564 4896 7620
rect 4896 7564 4952 7620
rect 4952 7564 4956 7620
rect 4892 7560 4956 7564
rect 53480 7620 53544 7624
rect 53480 7564 53484 7620
rect 53484 7564 53540 7620
rect 53540 7564 53544 7620
rect 53480 7560 53544 7564
rect 53560 7620 53624 7624
rect 53560 7564 53564 7620
rect 53564 7564 53620 7620
rect 53620 7564 53624 7620
rect 53560 7560 53624 7564
rect 53640 7620 53704 7624
rect 53640 7564 53644 7620
rect 53644 7564 53700 7620
rect 53700 7564 53704 7620
rect 53640 7560 53704 7564
rect 53720 7620 53784 7624
rect 53720 7564 53724 7620
rect 53724 7564 53780 7620
rect 53780 7564 53784 7620
rect 53720 7560 53784 7564
rect 53800 7620 53864 7624
rect 53800 7564 53804 7620
rect 53804 7564 53860 7620
rect 53860 7564 53864 7620
rect 53800 7560 53864 7564
rect 53880 7620 53944 7624
rect 53880 7564 53884 7620
rect 53884 7564 53940 7620
rect 53940 7564 53944 7620
rect 53880 7560 53944 7564
rect 53960 7620 54024 7624
rect 53960 7564 53964 7620
rect 53964 7564 54020 7620
rect 54020 7564 54024 7620
rect 53960 7560 54024 7564
rect 54040 7620 54104 7624
rect 54040 7564 54044 7620
rect 54044 7564 54100 7620
rect 54100 7564 54104 7620
rect 54040 7560 54104 7564
rect 54120 7620 54184 7624
rect 54120 7564 54124 7620
rect 54124 7564 54180 7620
rect 54180 7564 54184 7620
rect 54120 7560 54184 7564
rect 54200 7620 54264 7624
rect 54200 7564 54204 7620
rect 54204 7564 54260 7620
rect 54260 7564 54264 7620
rect 54200 7560 54264 7564
rect 54280 7620 54344 7624
rect 54280 7564 54284 7620
rect 54284 7564 54340 7620
rect 54340 7564 54344 7620
rect 54280 7560 54344 7564
rect 54360 7620 54424 7624
rect 54360 7564 54364 7620
rect 54364 7564 54420 7620
rect 54420 7564 54424 7620
rect 54360 7560 54424 7564
rect 54440 7620 54504 7624
rect 54440 7564 54444 7620
rect 54444 7564 54500 7620
rect 54500 7564 54504 7620
rect 54440 7560 54504 7564
rect 54520 7620 54584 7624
rect 54520 7564 54524 7620
rect 54524 7564 54580 7620
rect 54580 7564 54584 7620
rect 54520 7560 54584 7564
rect 54600 7620 54664 7624
rect 54600 7564 54604 7620
rect 54604 7564 54660 7620
rect 54660 7564 54664 7620
rect 54600 7560 54664 7564
rect 54680 7620 54744 7624
rect 54680 7564 54684 7620
rect 54684 7564 54740 7620
rect 54740 7564 54744 7620
rect 54680 7560 54744 7564
rect 54760 7620 54824 7624
rect 54760 7564 54764 7620
rect 54764 7564 54820 7620
rect 54820 7564 54824 7620
rect 54760 7560 54824 7564
rect 54840 7620 54904 7624
rect 54840 7564 54844 7620
rect 54844 7564 54900 7620
rect 54900 7564 54904 7620
rect 54840 7560 54904 7564
rect 54920 7620 54984 7624
rect 54920 7564 54924 7620
rect 54924 7564 54980 7620
rect 54980 7564 54984 7620
rect 54920 7560 54984 7564
rect 55000 7620 55064 7624
rect 55000 7564 55004 7620
rect 55004 7564 55060 7620
rect 55060 7564 55064 7620
rect 55000 7560 55064 7564
rect 924 5740 988 5744
rect 924 5684 928 5740
rect 928 5684 984 5740
rect 984 5684 988 5740
rect 924 5680 988 5684
rect 1004 5740 1068 5744
rect 1004 5684 1008 5740
rect 1008 5684 1064 5740
rect 1064 5684 1068 5740
rect 1004 5680 1068 5684
rect 1084 5740 1148 5744
rect 1084 5684 1088 5740
rect 1088 5684 1144 5740
rect 1144 5684 1148 5740
rect 1084 5680 1148 5684
rect 1164 5740 1228 5744
rect 1164 5684 1168 5740
rect 1168 5684 1224 5740
rect 1224 5684 1228 5740
rect 1164 5680 1228 5684
rect 1244 5740 1308 5744
rect 1244 5684 1248 5740
rect 1248 5684 1304 5740
rect 1304 5684 1308 5740
rect 1244 5680 1308 5684
rect 1324 5740 1388 5744
rect 1324 5684 1328 5740
rect 1328 5684 1384 5740
rect 1384 5684 1388 5740
rect 1324 5680 1388 5684
rect 1404 5740 1468 5744
rect 1404 5684 1408 5740
rect 1408 5684 1464 5740
rect 1464 5684 1468 5740
rect 1404 5680 1468 5684
rect 1484 5740 1548 5744
rect 1484 5684 1488 5740
rect 1488 5684 1544 5740
rect 1544 5684 1548 5740
rect 1484 5680 1548 5684
rect 1564 5740 1628 5744
rect 1564 5684 1568 5740
rect 1568 5684 1624 5740
rect 1624 5684 1628 5740
rect 1564 5680 1628 5684
rect 1644 5740 1708 5744
rect 1644 5684 1648 5740
rect 1648 5684 1704 5740
rect 1704 5684 1708 5740
rect 1644 5680 1708 5684
rect 1724 5740 1788 5744
rect 1724 5684 1728 5740
rect 1728 5684 1784 5740
rect 1784 5684 1788 5740
rect 1724 5680 1788 5684
rect 1804 5740 1868 5744
rect 1804 5684 1808 5740
rect 1808 5684 1864 5740
rect 1864 5684 1868 5740
rect 1804 5680 1868 5684
rect 1884 5740 1948 5744
rect 1884 5684 1888 5740
rect 1888 5684 1944 5740
rect 1944 5684 1948 5740
rect 1884 5680 1948 5684
rect 1964 5740 2028 5744
rect 1964 5684 1968 5740
rect 1968 5684 2024 5740
rect 2024 5684 2028 5740
rect 1964 5680 2028 5684
rect 2044 5740 2108 5744
rect 2044 5684 2048 5740
rect 2048 5684 2104 5740
rect 2104 5684 2108 5740
rect 2044 5680 2108 5684
rect 2124 5740 2188 5744
rect 2124 5684 2128 5740
rect 2128 5684 2184 5740
rect 2184 5684 2188 5740
rect 2124 5680 2188 5684
rect 2204 5740 2268 5744
rect 2204 5684 2208 5740
rect 2208 5684 2264 5740
rect 2264 5684 2268 5740
rect 2204 5680 2268 5684
rect 2284 5740 2348 5744
rect 2284 5684 2288 5740
rect 2288 5684 2344 5740
rect 2344 5684 2348 5740
rect 2284 5680 2348 5684
rect 2364 5740 2428 5744
rect 2364 5684 2368 5740
rect 2368 5684 2424 5740
rect 2424 5684 2428 5740
rect 2364 5680 2428 5684
rect 2444 5740 2508 5744
rect 2444 5684 2448 5740
rect 2448 5684 2504 5740
rect 2504 5684 2508 5740
rect 2444 5680 2508 5684
rect 55928 5740 55992 5744
rect 55928 5684 55932 5740
rect 55932 5684 55988 5740
rect 55988 5684 55992 5740
rect 55928 5680 55992 5684
rect 56008 5740 56072 5744
rect 56008 5684 56012 5740
rect 56012 5684 56068 5740
rect 56068 5684 56072 5740
rect 56008 5680 56072 5684
rect 56088 5740 56152 5744
rect 56088 5684 56092 5740
rect 56092 5684 56148 5740
rect 56148 5684 56152 5740
rect 56088 5680 56152 5684
rect 56168 5740 56232 5744
rect 56168 5684 56172 5740
rect 56172 5684 56228 5740
rect 56228 5684 56232 5740
rect 56168 5680 56232 5684
rect 56248 5740 56312 5744
rect 56248 5684 56252 5740
rect 56252 5684 56308 5740
rect 56308 5684 56312 5740
rect 56248 5680 56312 5684
rect 56328 5740 56392 5744
rect 56328 5684 56332 5740
rect 56332 5684 56388 5740
rect 56388 5684 56392 5740
rect 56328 5680 56392 5684
rect 56408 5740 56472 5744
rect 56408 5684 56412 5740
rect 56412 5684 56468 5740
rect 56468 5684 56472 5740
rect 56408 5680 56472 5684
rect 56488 5740 56552 5744
rect 56488 5684 56492 5740
rect 56492 5684 56548 5740
rect 56548 5684 56552 5740
rect 56488 5680 56552 5684
rect 56568 5740 56632 5744
rect 56568 5684 56572 5740
rect 56572 5684 56628 5740
rect 56628 5684 56632 5740
rect 56568 5680 56632 5684
rect 56648 5740 56712 5744
rect 56648 5684 56652 5740
rect 56652 5684 56708 5740
rect 56708 5684 56712 5740
rect 56648 5680 56712 5684
rect 56728 5740 56792 5744
rect 56728 5684 56732 5740
rect 56732 5684 56788 5740
rect 56788 5684 56792 5740
rect 56728 5680 56792 5684
rect 56808 5740 56872 5744
rect 56808 5684 56812 5740
rect 56812 5684 56868 5740
rect 56868 5684 56872 5740
rect 56808 5680 56872 5684
rect 56888 5740 56952 5744
rect 56888 5684 56892 5740
rect 56892 5684 56948 5740
rect 56948 5684 56952 5740
rect 56888 5680 56952 5684
rect 56968 5740 57032 5744
rect 56968 5684 56972 5740
rect 56972 5684 57028 5740
rect 57028 5684 57032 5740
rect 56968 5680 57032 5684
rect 57048 5740 57112 5744
rect 57048 5684 57052 5740
rect 57052 5684 57108 5740
rect 57108 5684 57112 5740
rect 57048 5680 57112 5684
rect 57128 5740 57192 5744
rect 57128 5684 57132 5740
rect 57132 5684 57188 5740
rect 57188 5684 57192 5740
rect 57128 5680 57192 5684
rect 57208 5740 57272 5744
rect 57208 5684 57212 5740
rect 57212 5684 57268 5740
rect 57268 5684 57272 5740
rect 57208 5680 57272 5684
rect 57288 5740 57352 5744
rect 57288 5684 57292 5740
rect 57292 5684 57348 5740
rect 57348 5684 57352 5740
rect 57288 5680 57352 5684
rect 57368 5740 57432 5744
rect 57368 5684 57372 5740
rect 57372 5684 57428 5740
rect 57428 5684 57432 5740
rect 57368 5680 57432 5684
rect 57448 5740 57512 5744
rect 57448 5684 57452 5740
rect 57452 5684 57508 5740
rect 57508 5684 57512 5740
rect 57448 5680 57512 5684
<< mimcap >>
rect 6017 48574 6417 48622
rect 6017 48270 6065 48574
rect 6369 48270 6417 48574
rect 6017 48222 6417 48270
rect 6736 48574 7136 48622
rect 6736 48270 6784 48574
rect 7088 48270 7136 48574
rect 6736 48222 7136 48270
rect 7455 48574 7855 48622
rect 7455 48270 7503 48574
rect 7807 48270 7855 48574
rect 7455 48222 7855 48270
rect 8174 48574 8574 48622
rect 8174 48270 8222 48574
rect 8526 48270 8574 48574
rect 8174 48222 8574 48270
rect 8893 48574 9293 48622
rect 8893 48270 8941 48574
rect 9245 48270 9293 48574
rect 8893 48222 9293 48270
rect 9612 48574 10012 48622
rect 9612 48270 9660 48574
rect 9964 48270 10012 48574
rect 9612 48222 10012 48270
rect 10331 48574 10731 48622
rect 10331 48270 10379 48574
rect 10683 48270 10731 48574
rect 10331 48222 10731 48270
rect 11050 48574 11450 48622
rect 11050 48270 11098 48574
rect 11402 48270 11450 48574
rect 11050 48222 11450 48270
rect 11769 48574 12169 48622
rect 11769 48270 11817 48574
rect 12121 48270 12169 48574
rect 11769 48222 12169 48270
rect 12488 48574 12888 48622
rect 12488 48270 12536 48574
rect 12840 48270 12888 48574
rect 12488 48222 12888 48270
rect 13465 48574 13865 48622
rect 13465 48270 13513 48574
rect 13817 48270 13865 48574
rect 13465 48222 13865 48270
rect 14184 48574 14584 48622
rect 14184 48270 14232 48574
rect 14536 48270 14584 48574
rect 14184 48222 14584 48270
rect 14903 48574 15303 48622
rect 14903 48270 14951 48574
rect 15255 48270 15303 48574
rect 14903 48222 15303 48270
rect 15622 48574 16022 48622
rect 15622 48270 15670 48574
rect 15974 48270 16022 48574
rect 15622 48222 16022 48270
rect 16341 48574 16741 48622
rect 16341 48270 16389 48574
rect 16693 48270 16741 48574
rect 16341 48222 16741 48270
rect 17060 48574 17460 48622
rect 17060 48270 17108 48574
rect 17412 48270 17460 48574
rect 17060 48222 17460 48270
rect 17779 48574 18179 48622
rect 17779 48270 17827 48574
rect 18131 48270 18179 48574
rect 17779 48222 18179 48270
rect 18498 48574 18898 48622
rect 18498 48270 18546 48574
rect 18850 48270 18898 48574
rect 18498 48222 18898 48270
rect 19217 48574 19617 48622
rect 19217 48270 19265 48574
rect 19569 48270 19617 48574
rect 19217 48222 19617 48270
rect 19936 48574 20336 48622
rect 19936 48270 19984 48574
rect 20288 48270 20336 48574
rect 19936 48222 20336 48270
rect 6017 47874 6417 47922
rect 6017 47570 6065 47874
rect 6369 47570 6417 47874
rect 6017 47522 6417 47570
rect 6736 47874 7136 47922
rect 6736 47570 6784 47874
rect 7088 47570 7136 47874
rect 6736 47522 7136 47570
rect 7455 47874 7855 47922
rect 7455 47570 7503 47874
rect 7807 47570 7855 47874
rect 7455 47522 7855 47570
rect 8174 47874 8574 47922
rect 8174 47570 8222 47874
rect 8526 47570 8574 47874
rect 8174 47522 8574 47570
rect 8893 47874 9293 47922
rect 8893 47570 8941 47874
rect 9245 47570 9293 47874
rect 8893 47522 9293 47570
rect 9612 47874 10012 47922
rect 9612 47570 9660 47874
rect 9964 47570 10012 47874
rect 9612 47522 10012 47570
rect 10331 47874 10731 47922
rect 10331 47570 10379 47874
rect 10683 47570 10731 47874
rect 10331 47522 10731 47570
rect 11050 47874 11450 47922
rect 11050 47570 11098 47874
rect 11402 47570 11450 47874
rect 11050 47522 11450 47570
rect 11769 47874 12169 47922
rect 11769 47570 11817 47874
rect 12121 47570 12169 47874
rect 11769 47522 12169 47570
rect 12488 47874 12888 47922
rect 12488 47570 12536 47874
rect 12840 47570 12888 47874
rect 12488 47522 12888 47570
rect 13465 47874 13865 47922
rect 13465 47570 13513 47874
rect 13817 47570 13865 47874
rect 13465 47522 13865 47570
rect 14184 47874 14584 47922
rect 14184 47570 14232 47874
rect 14536 47570 14584 47874
rect 14184 47522 14584 47570
rect 14903 47874 15303 47922
rect 14903 47570 14951 47874
rect 15255 47570 15303 47874
rect 14903 47522 15303 47570
rect 15622 47874 16022 47922
rect 15622 47570 15670 47874
rect 15974 47570 16022 47874
rect 15622 47522 16022 47570
rect 16341 47874 16741 47922
rect 16341 47570 16389 47874
rect 16693 47570 16741 47874
rect 16341 47522 16741 47570
rect 17060 47874 17460 47922
rect 17060 47570 17108 47874
rect 17412 47570 17460 47874
rect 17060 47522 17460 47570
rect 17779 47874 18179 47922
rect 17779 47570 17827 47874
rect 18131 47570 18179 47874
rect 17779 47522 18179 47570
rect 18498 47874 18898 47922
rect 18498 47570 18546 47874
rect 18850 47570 18898 47874
rect 18498 47522 18898 47570
rect 19217 47874 19617 47922
rect 19217 47570 19265 47874
rect 19569 47570 19617 47874
rect 19217 47522 19617 47570
rect 19936 47874 20336 47922
rect 19936 47570 19984 47874
rect 20288 47570 20336 47874
rect 19936 47522 20336 47570
rect 6017 44814 6417 44862
rect 6017 44510 6065 44814
rect 6369 44510 6417 44814
rect 6017 44462 6417 44510
rect 6736 44814 7136 44862
rect 6736 44510 6784 44814
rect 7088 44510 7136 44814
rect 6736 44462 7136 44510
rect 7455 44814 7855 44862
rect 7455 44510 7503 44814
rect 7807 44510 7855 44814
rect 7455 44462 7855 44510
rect 8174 44814 8574 44862
rect 8174 44510 8222 44814
rect 8526 44510 8574 44814
rect 8174 44462 8574 44510
rect 8893 44814 9293 44862
rect 8893 44510 8941 44814
rect 9245 44510 9293 44814
rect 8893 44462 9293 44510
rect 9612 44814 10012 44862
rect 9612 44510 9660 44814
rect 9964 44510 10012 44814
rect 9612 44462 10012 44510
rect 10331 44814 10731 44862
rect 10331 44510 10379 44814
rect 10683 44510 10731 44814
rect 10331 44462 10731 44510
rect 11050 44814 11450 44862
rect 11050 44510 11098 44814
rect 11402 44510 11450 44814
rect 11050 44462 11450 44510
rect 11769 44814 12169 44862
rect 11769 44510 11817 44814
rect 12121 44510 12169 44814
rect 11769 44462 12169 44510
rect 12488 44814 12888 44862
rect 12488 44510 12536 44814
rect 12840 44510 12888 44814
rect 12488 44462 12888 44510
rect 6017 44114 6417 44162
rect 6017 43810 6065 44114
rect 6369 43810 6417 44114
rect 6017 43762 6417 43810
rect 6736 44114 7136 44162
rect 6736 43810 6784 44114
rect 7088 43810 7136 44114
rect 6736 43762 7136 43810
rect 7455 44114 7855 44162
rect 7455 43810 7503 44114
rect 7807 43810 7855 44114
rect 7455 43762 7855 43810
rect 8174 44114 8574 44162
rect 8174 43810 8222 44114
rect 8526 43810 8574 44114
rect 8174 43762 8574 43810
rect 8893 44114 9293 44162
rect 8893 43810 8941 44114
rect 9245 43810 9293 44114
rect 8893 43762 9293 43810
rect 9612 44114 10012 44162
rect 9612 43810 9660 44114
rect 9964 43810 10012 44114
rect 9612 43762 10012 43810
rect 10331 44114 10731 44162
rect 10331 43810 10379 44114
rect 10683 43810 10731 44114
rect 10331 43762 10731 43810
rect 11050 44114 11450 44162
rect 11050 43810 11098 44114
rect 11402 43810 11450 44114
rect 11050 43762 11450 43810
rect 11769 44114 12169 44162
rect 11769 43810 11817 44114
rect 12121 43810 12169 44114
rect 11769 43762 12169 43810
rect 12488 44114 12888 44162
rect 12488 43810 12536 44114
rect 12840 43810 12888 44114
rect 12488 43762 12888 43810
rect 6409 41054 6809 41102
rect 6409 40750 6457 41054
rect 6761 40750 6809 41054
rect 6409 40702 6809 40750
rect 7128 41054 7528 41102
rect 7128 40750 7176 41054
rect 7480 40750 7528 41054
rect 7128 40702 7528 40750
rect 7847 41054 8247 41102
rect 7847 40750 7895 41054
rect 8199 40750 8247 41054
rect 7847 40702 8247 40750
rect 8566 41054 8966 41102
rect 8566 40750 8614 41054
rect 8918 40750 8966 41054
rect 8566 40702 8966 40750
rect 9285 41054 9685 41102
rect 9285 40750 9333 41054
rect 9637 40750 9685 41054
rect 9285 40702 9685 40750
rect 10004 41054 10404 41102
rect 10004 40750 10052 41054
rect 10356 40750 10404 41054
rect 10004 40702 10404 40750
rect 10723 41054 11123 41102
rect 10723 40750 10771 41054
rect 11075 40750 11123 41054
rect 10723 40702 11123 40750
rect 11442 41054 11842 41102
rect 11442 40750 11490 41054
rect 11794 40750 11842 41054
rect 11442 40702 11842 40750
rect 12161 41054 12561 41102
rect 12161 40750 12209 41054
rect 12513 40750 12561 41054
rect 12161 40702 12561 40750
rect 12880 41054 13280 41102
rect 12880 40750 12928 41054
rect 13232 40750 13280 41054
rect 12880 40702 13280 40750
rect 15229 41054 15629 41102
rect 15229 40750 15277 41054
rect 15581 40750 15629 41054
rect 15229 40702 15629 40750
rect 15948 41054 16348 41102
rect 15948 40750 15996 41054
rect 16300 40750 16348 41054
rect 15948 40702 16348 40750
rect 16667 41054 17067 41102
rect 16667 40750 16715 41054
rect 17019 40750 17067 41054
rect 16667 40702 17067 40750
rect 17386 41054 17786 41102
rect 17386 40750 17434 41054
rect 17738 40750 17786 41054
rect 17386 40702 17786 40750
rect 18105 41054 18505 41102
rect 18105 40750 18153 41054
rect 18457 40750 18505 41054
rect 18105 40702 18505 40750
rect 18824 41054 19224 41102
rect 18824 40750 18872 41054
rect 19176 40750 19224 41054
rect 18824 40702 19224 40750
rect 19543 41054 19943 41102
rect 19543 40750 19591 41054
rect 19895 40750 19943 41054
rect 19543 40702 19943 40750
rect 20262 41054 20662 41102
rect 20262 40750 20310 41054
rect 20614 40750 20662 41054
rect 20262 40702 20662 40750
rect 20981 41054 21381 41102
rect 20981 40750 21029 41054
rect 21333 40750 21381 41054
rect 20981 40702 21381 40750
rect 21700 41054 22100 41102
rect 21700 40750 21748 41054
rect 22052 40750 22100 41054
rect 21700 40702 22100 40750
rect 6409 40354 6809 40402
rect 6409 40050 6457 40354
rect 6761 40050 6809 40354
rect 6409 40002 6809 40050
rect 7128 40354 7528 40402
rect 7128 40050 7176 40354
rect 7480 40050 7528 40354
rect 7128 40002 7528 40050
rect 7847 40354 8247 40402
rect 7847 40050 7895 40354
rect 8199 40050 8247 40354
rect 7847 40002 8247 40050
rect 8566 40354 8966 40402
rect 8566 40050 8614 40354
rect 8918 40050 8966 40354
rect 8566 40002 8966 40050
rect 9285 40354 9685 40402
rect 9285 40050 9333 40354
rect 9637 40050 9685 40354
rect 9285 40002 9685 40050
rect 10004 40354 10404 40402
rect 10004 40050 10052 40354
rect 10356 40050 10404 40354
rect 10004 40002 10404 40050
rect 10723 40354 11123 40402
rect 10723 40050 10771 40354
rect 11075 40050 11123 40354
rect 10723 40002 11123 40050
rect 11442 40354 11842 40402
rect 11442 40050 11490 40354
rect 11794 40050 11842 40354
rect 11442 40002 11842 40050
rect 12161 40354 12561 40402
rect 12161 40050 12209 40354
rect 12513 40050 12561 40354
rect 12161 40002 12561 40050
rect 12880 40354 13280 40402
rect 12880 40050 12928 40354
rect 13232 40050 13280 40354
rect 12880 40002 13280 40050
rect 15229 40354 15629 40402
rect 15229 40050 15277 40354
rect 15581 40050 15629 40354
rect 15229 40002 15629 40050
rect 15948 40354 16348 40402
rect 15948 40050 15996 40354
rect 16300 40050 16348 40354
rect 15948 40002 16348 40050
rect 16667 40354 17067 40402
rect 16667 40050 16715 40354
rect 17019 40050 17067 40354
rect 16667 40002 17067 40050
rect 17386 40354 17786 40402
rect 17386 40050 17434 40354
rect 17738 40050 17786 40354
rect 17386 40002 17786 40050
rect 18105 40354 18505 40402
rect 18105 40050 18153 40354
rect 18457 40050 18505 40354
rect 18105 40002 18505 40050
rect 18824 40354 19224 40402
rect 18824 40050 18872 40354
rect 19176 40050 19224 40354
rect 18824 40002 19224 40050
rect 19543 40354 19943 40402
rect 19543 40050 19591 40354
rect 19895 40050 19943 40354
rect 19543 40002 19943 40050
rect 20262 40354 20662 40402
rect 20262 40050 20310 40354
rect 20614 40050 20662 40354
rect 20262 40002 20662 40050
rect 20981 40354 21381 40402
rect 20981 40050 21029 40354
rect 21333 40050 21381 40354
rect 20981 40002 21381 40050
rect 21700 40354 22100 40402
rect 21700 40050 21748 40354
rect 22052 40050 22100 40354
rect 21700 40002 22100 40050
rect 30027 37294 30427 37342
rect 30027 36990 30075 37294
rect 30379 36990 30427 37294
rect 30027 36942 30427 36990
rect 30746 37294 31146 37342
rect 30746 36990 30794 37294
rect 31098 36990 31146 37294
rect 30746 36942 31146 36990
rect 31465 37294 31865 37342
rect 31465 36990 31513 37294
rect 31817 36990 31865 37294
rect 31465 36942 31865 36990
rect 32184 37294 32584 37342
rect 32184 36990 32232 37294
rect 32536 36990 32584 37294
rect 32184 36942 32584 36990
rect 32903 37294 33303 37342
rect 32903 36990 32951 37294
rect 33255 36990 33303 37294
rect 32903 36942 33303 36990
rect 33622 37294 34022 37342
rect 33622 36990 33670 37294
rect 33974 36990 34022 37294
rect 33622 36942 34022 36990
rect 34341 37294 34741 37342
rect 34341 36990 34389 37294
rect 34693 36990 34741 37294
rect 34341 36942 34741 36990
rect 35060 37294 35460 37342
rect 35060 36990 35108 37294
rect 35412 36990 35460 37294
rect 35060 36942 35460 36990
rect 35779 37294 36179 37342
rect 35779 36990 35827 37294
rect 36131 36990 36179 37294
rect 35779 36942 36179 36990
rect 36498 37294 36898 37342
rect 36498 36990 36546 37294
rect 36850 36990 36898 37294
rect 36498 36942 36898 36990
rect 30027 36594 30427 36642
rect 30027 36290 30075 36594
rect 30379 36290 30427 36594
rect 30027 36242 30427 36290
rect 30746 36594 31146 36642
rect 30746 36290 30794 36594
rect 31098 36290 31146 36594
rect 30746 36242 31146 36290
rect 31465 36594 31865 36642
rect 31465 36290 31513 36594
rect 31817 36290 31865 36594
rect 31465 36242 31865 36290
rect 32184 36594 32584 36642
rect 32184 36290 32232 36594
rect 32536 36290 32584 36594
rect 32184 36242 32584 36290
rect 32903 36594 33303 36642
rect 32903 36290 32951 36594
rect 33255 36290 33303 36594
rect 32903 36242 33303 36290
rect 33622 36594 34022 36642
rect 33622 36290 33670 36594
rect 33974 36290 34022 36594
rect 33622 36242 34022 36290
rect 34341 36594 34741 36642
rect 34341 36290 34389 36594
rect 34693 36290 34741 36594
rect 34341 36242 34741 36290
rect 35060 36594 35460 36642
rect 35060 36290 35108 36594
rect 35412 36290 35460 36594
rect 35060 36242 35460 36290
rect 35779 36594 36179 36642
rect 35779 36290 35827 36594
rect 36131 36290 36179 36594
rect 35779 36242 36179 36290
rect 36498 36594 36898 36642
rect 36498 36290 36546 36594
rect 36850 36290 36898 36594
rect 36498 36242 36898 36290
rect 26303 33534 26703 33582
rect 26303 33230 26351 33534
rect 26655 33230 26703 33534
rect 26303 33182 26703 33230
rect 27022 33534 27422 33582
rect 27022 33230 27070 33534
rect 27374 33230 27422 33534
rect 27022 33182 27422 33230
rect 27741 33534 28141 33582
rect 27741 33230 27789 33534
rect 28093 33230 28141 33534
rect 27741 33182 28141 33230
rect 28460 33534 28860 33582
rect 28460 33230 28508 33534
rect 28812 33230 28860 33534
rect 28460 33182 28860 33230
rect 29179 33534 29579 33582
rect 29179 33230 29227 33534
rect 29531 33230 29579 33534
rect 29179 33182 29579 33230
rect 29898 33534 30298 33582
rect 29898 33230 29946 33534
rect 30250 33230 30298 33534
rect 29898 33182 30298 33230
rect 30617 33534 31017 33582
rect 30617 33230 30665 33534
rect 30969 33230 31017 33534
rect 30617 33182 31017 33230
rect 31336 33534 31736 33582
rect 31336 33230 31384 33534
rect 31688 33230 31736 33534
rect 31336 33182 31736 33230
rect 32055 33534 32455 33582
rect 32055 33230 32103 33534
rect 32407 33230 32455 33534
rect 32055 33182 32455 33230
rect 32774 33534 33174 33582
rect 32774 33230 32822 33534
rect 33126 33230 33174 33534
rect 32774 33182 33174 33230
rect 33751 33534 34151 33582
rect 33751 33230 33799 33534
rect 34103 33230 34151 33534
rect 33751 33182 34151 33230
rect 34470 33534 34870 33582
rect 34470 33230 34518 33534
rect 34822 33230 34870 33534
rect 34470 33182 34870 33230
rect 35189 33534 35589 33582
rect 35189 33230 35237 33534
rect 35541 33230 35589 33534
rect 35189 33182 35589 33230
rect 35908 33534 36308 33582
rect 35908 33230 35956 33534
rect 36260 33230 36308 33534
rect 35908 33182 36308 33230
rect 36627 33534 37027 33582
rect 36627 33230 36675 33534
rect 36979 33230 37027 33534
rect 36627 33182 37027 33230
rect 37346 33534 37746 33582
rect 37346 33230 37394 33534
rect 37698 33230 37746 33534
rect 37346 33182 37746 33230
rect 38065 33534 38465 33582
rect 38065 33230 38113 33534
rect 38417 33230 38465 33534
rect 38065 33182 38465 33230
rect 38784 33534 39184 33582
rect 38784 33230 38832 33534
rect 39136 33230 39184 33534
rect 38784 33182 39184 33230
rect 39503 33534 39903 33582
rect 39503 33230 39551 33534
rect 39855 33230 39903 33534
rect 39503 33182 39903 33230
rect 40222 33534 40622 33582
rect 40222 33230 40270 33534
rect 40574 33230 40622 33534
rect 40222 33182 40622 33230
rect 26303 32834 26703 32882
rect 26303 32530 26351 32834
rect 26655 32530 26703 32834
rect 26303 32482 26703 32530
rect 27022 32834 27422 32882
rect 27022 32530 27070 32834
rect 27374 32530 27422 32834
rect 27022 32482 27422 32530
rect 27741 32834 28141 32882
rect 27741 32530 27789 32834
rect 28093 32530 28141 32834
rect 27741 32482 28141 32530
rect 28460 32834 28860 32882
rect 28460 32530 28508 32834
rect 28812 32530 28860 32834
rect 28460 32482 28860 32530
rect 29179 32834 29579 32882
rect 29179 32530 29227 32834
rect 29531 32530 29579 32834
rect 29179 32482 29579 32530
rect 29898 32834 30298 32882
rect 29898 32530 29946 32834
rect 30250 32530 30298 32834
rect 29898 32482 30298 32530
rect 30617 32834 31017 32882
rect 30617 32530 30665 32834
rect 30969 32530 31017 32834
rect 30617 32482 31017 32530
rect 31336 32834 31736 32882
rect 31336 32530 31384 32834
rect 31688 32530 31736 32834
rect 31336 32482 31736 32530
rect 32055 32834 32455 32882
rect 32055 32530 32103 32834
rect 32407 32530 32455 32834
rect 32055 32482 32455 32530
rect 32774 32834 33174 32882
rect 32774 32530 32822 32834
rect 33126 32530 33174 32834
rect 32774 32482 33174 32530
rect 33751 32834 34151 32882
rect 33751 32530 33799 32834
rect 34103 32530 34151 32834
rect 33751 32482 34151 32530
rect 34470 32834 34870 32882
rect 34470 32530 34518 32834
rect 34822 32530 34870 32834
rect 34470 32482 34870 32530
rect 35189 32834 35589 32882
rect 35189 32530 35237 32834
rect 35541 32530 35589 32834
rect 35189 32482 35589 32530
rect 35908 32834 36308 32882
rect 35908 32530 35956 32834
rect 36260 32530 36308 32834
rect 35908 32482 36308 32530
rect 36627 32834 37027 32882
rect 36627 32530 36675 32834
rect 36979 32530 37027 32834
rect 36627 32482 37027 32530
rect 37346 32834 37746 32882
rect 37346 32530 37394 32834
rect 37698 32530 37746 32834
rect 37346 32482 37746 32530
rect 38065 32834 38465 32882
rect 38065 32530 38113 32834
rect 38417 32530 38465 32834
rect 38065 32482 38465 32530
rect 38784 32834 39184 32882
rect 38784 32530 38832 32834
rect 39136 32530 39184 32834
rect 38784 32482 39184 32530
rect 39503 32834 39903 32882
rect 39503 32530 39551 32834
rect 39855 32530 39903 32834
rect 39503 32482 39903 32530
rect 40222 32834 40622 32882
rect 40222 32530 40270 32834
rect 40574 32530 40622 32834
rect 40222 32482 40622 32530
rect 30027 29774 30427 29822
rect 30027 29470 30075 29774
rect 30379 29470 30427 29774
rect 30027 29422 30427 29470
rect 30746 29774 31146 29822
rect 30746 29470 30794 29774
rect 31098 29470 31146 29774
rect 30746 29422 31146 29470
rect 31465 29774 31865 29822
rect 31465 29470 31513 29774
rect 31817 29470 31865 29774
rect 31465 29422 31865 29470
rect 32184 29774 32584 29822
rect 32184 29470 32232 29774
rect 32536 29470 32584 29774
rect 32184 29422 32584 29470
rect 32903 29774 33303 29822
rect 32903 29470 32951 29774
rect 33255 29470 33303 29774
rect 32903 29422 33303 29470
rect 33622 29774 34022 29822
rect 33622 29470 33670 29774
rect 33974 29470 34022 29774
rect 33622 29422 34022 29470
rect 34341 29774 34741 29822
rect 34341 29470 34389 29774
rect 34693 29470 34741 29774
rect 34341 29422 34741 29470
rect 35060 29774 35460 29822
rect 35060 29470 35108 29774
rect 35412 29470 35460 29774
rect 35060 29422 35460 29470
rect 35779 29774 36179 29822
rect 35779 29470 35827 29774
rect 36131 29470 36179 29774
rect 35779 29422 36179 29470
rect 36498 29774 36898 29822
rect 36498 29470 36546 29774
rect 36850 29470 36898 29774
rect 36498 29422 36898 29470
rect 30027 29074 30427 29122
rect 30027 28770 30075 29074
rect 30379 28770 30427 29074
rect 30027 28722 30427 28770
rect 30746 29074 31146 29122
rect 30746 28770 30794 29074
rect 31098 28770 31146 29074
rect 30746 28722 31146 28770
rect 31465 29074 31865 29122
rect 31465 28770 31513 29074
rect 31817 28770 31865 29074
rect 31465 28722 31865 28770
rect 32184 29074 32584 29122
rect 32184 28770 32232 29074
rect 32536 28770 32584 29074
rect 32184 28722 32584 28770
rect 32903 29074 33303 29122
rect 32903 28770 32951 29074
rect 33255 28770 33303 29074
rect 32903 28722 33303 28770
rect 33622 29074 34022 29122
rect 33622 28770 33670 29074
rect 33974 28770 34022 29074
rect 33622 28722 34022 28770
rect 34341 29074 34741 29122
rect 34341 28770 34389 29074
rect 34693 28770 34741 29074
rect 34341 28722 34741 28770
rect 35060 29074 35460 29122
rect 35060 28770 35108 29074
rect 35412 28770 35460 29074
rect 35060 28722 35460 28770
rect 35779 29074 36179 29122
rect 35779 28770 35827 29074
rect 36131 28770 36179 29074
rect 35779 28722 36179 28770
rect 36498 29074 36898 29122
rect 36498 28770 36546 29074
rect 36850 28770 36898 29074
rect 36498 28722 36898 28770
rect 30027 26014 30427 26062
rect 30027 25710 30075 26014
rect 30379 25710 30427 26014
rect 30027 25662 30427 25710
rect 30746 26014 31146 26062
rect 30746 25710 30794 26014
rect 31098 25710 31146 26014
rect 30746 25662 31146 25710
rect 31465 26014 31865 26062
rect 31465 25710 31513 26014
rect 31817 25710 31865 26014
rect 31465 25662 31865 25710
rect 32184 26014 32584 26062
rect 32184 25710 32232 26014
rect 32536 25710 32584 26014
rect 32184 25662 32584 25710
rect 32903 26014 33303 26062
rect 32903 25710 32951 26014
rect 33255 25710 33303 26014
rect 32903 25662 33303 25710
rect 33622 26014 34022 26062
rect 33622 25710 33670 26014
rect 33974 25710 34022 26014
rect 33622 25662 34022 25710
rect 34341 26014 34741 26062
rect 34341 25710 34389 26014
rect 34693 25710 34741 26014
rect 34341 25662 34741 25710
rect 35060 26014 35460 26062
rect 35060 25710 35108 26014
rect 35412 25710 35460 26014
rect 35060 25662 35460 25710
rect 35779 26014 36179 26062
rect 35779 25710 35827 26014
rect 36131 25710 36179 26014
rect 35779 25662 36179 25710
rect 36498 26014 36898 26062
rect 36498 25710 36546 26014
rect 36850 25710 36898 26014
rect 36498 25662 36898 25710
rect 30027 25314 30427 25362
rect 30027 25010 30075 25314
rect 30379 25010 30427 25314
rect 30027 24962 30427 25010
rect 30746 25314 31146 25362
rect 30746 25010 30794 25314
rect 31098 25010 31146 25314
rect 30746 24962 31146 25010
rect 31465 25314 31865 25362
rect 31465 25010 31513 25314
rect 31817 25010 31865 25314
rect 31465 24962 31865 25010
rect 32184 25314 32584 25362
rect 32184 25010 32232 25314
rect 32536 25010 32584 25314
rect 32184 24962 32584 25010
rect 32903 25314 33303 25362
rect 32903 25010 32951 25314
rect 33255 25010 33303 25314
rect 32903 24962 33303 25010
rect 33622 25314 34022 25362
rect 33622 25010 33670 25314
rect 33974 25010 34022 25314
rect 33622 24962 34022 25010
rect 34341 25314 34741 25362
rect 34341 25010 34389 25314
rect 34693 25010 34741 25314
rect 34341 24962 34741 25010
rect 35060 25314 35460 25362
rect 35060 25010 35108 25314
rect 35412 25010 35460 25314
rect 35060 24962 35460 25010
rect 35779 25314 36179 25362
rect 35779 25010 35827 25314
rect 36131 25010 36179 25314
rect 35779 24962 36179 25010
rect 36498 25314 36898 25362
rect 36498 25010 36546 25314
rect 36850 25010 36898 25314
rect 36498 24962 36898 25010
<< mimcapcontact >>
rect 6065 48270 6369 48574
rect 6784 48270 7088 48574
rect 7503 48270 7807 48574
rect 8222 48270 8526 48574
rect 8941 48270 9245 48574
rect 9660 48270 9964 48574
rect 10379 48270 10683 48574
rect 11098 48270 11402 48574
rect 11817 48270 12121 48574
rect 12536 48270 12840 48574
rect 13513 48270 13817 48574
rect 14232 48270 14536 48574
rect 14951 48270 15255 48574
rect 15670 48270 15974 48574
rect 16389 48270 16693 48574
rect 17108 48270 17412 48574
rect 17827 48270 18131 48574
rect 18546 48270 18850 48574
rect 19265 48270 19569 48574
rect 19984 48270 20288 48574
rect 6065 47570 6369 47874
rect 6784 47570 7088 47874
rect 7503 47570 7807 47874
rect 8222 47570 8526 47874
rect 8941 47570 9245 47874
rect 9660 47570 9964 47874
rect 10379 47570 10683 47874
rect 11098 47570 11402 47874
rect 11817 47570 12121 47874
rect 12536 47570 12840 47874
rect 13513 47570 13817 47874
rect 14232 47570 14536 47874
rect 14951 47570 15255 47874
rect 15670 47570 15974 47874
rect 16389 47570 16693 47874
rect 17108 47570 17412 47874
rect 17827 47570 18131 47874
rect 18546 47570 18850 47874
rect 19265 47570 19569 47874
rect 19984 47570 20288 47874
rect 6065 44510 6369 44814
rect 6784 44510 7088 44814
rect 7503 44510 7807 44814
rect 8222 44510 8526 44814
rect 8941 44510 9245 44814
rect 9660 44510 9964 44814
rect 10379 44510 10683 44814
rect 11098 44510 11402 44814
rect 11817 44510 12121 44814
rect 12536 44510 12840 44814
rect 6065 43810 6369 44114
rect 6784 43810 7088 44114
rect 7503 43810 7807 44114
rect 8222 43810 8526 44114
rect 8941 43810 9245 44114
rect 9660 43810 9964 44114
rect 10379 43810 10683 44114
rect 11098 43810 11402 44114
rect 11817 43810 12121 44114
rect 12536 43810 12840 44114
rect 6457 40750 6761 41054
rect 7176 40750 7480 41054
rect 7895 40750 8199 41054
rect 8614 40750 8918 41054
rect 9333 40750 9637 41054
rect 10052 40750 10356 41054
rect 10771 40750 11075 41054
rect 11490 40750 11794 41054
rect 12209 40750 12513 41054
rect 12928 40750 13232 41054
rect 15277 40750 15581 41054
rect 15996 40750 16300 41054
rect 16715 40750 17019 41054
rect 17434 40750 17738 41054
rect 18153 40750 18457 41054
rect 18872 40750 19176 41054
rect 19591 40750 19895 41054
rect 20310 40750 20614 41054
rect 21029 40750 21333 41054
rect 21748 40750 22052 41054
rect 6457 40050 6761 40354
rect 7176 40050 7480 40354
rect 7895 40050 8199 40354
rect 8614 40050 8918 40354
rect 9333 40050 9637 40354
rect 10052 40050 10356 40354
rect 10771 40050 11075 40354
rect 11490 40050 11794 40354
rect 12209 40050 12513 40354
rect 12928 40050 13232 40354
rect 15277 40050 15581 40354
rect 15996 40050 16300 40354
rect 16715 40050 17019 40354
rect 17434 40050 17738 40354
rect 18153 40050 18457 40354
rect 18872 40050 19176 40354
rect 19591 40050 19895 40354
rect 20310 40050 20614 40354
rect 21029 40050 21333 40354
rect 21748 40050 22052 40354
rect 30075 36990 30379 37294
rect 30794 36990 31098 37294
rect 31513 36990 31817 37294
rect 32232 36990 32536 37294
rect 32951 36990 33255 37294
rect 33670 36990 33974 37294
rect 34389 36990 34693 37294
rect 35108 36990 35412 37294
rect 35827 36990 36131 37294
rect 36546 36990 36850 37294
rect 30075 36290 30379 36594
rect 30794 36290 31098 36594
rect 31513 36290 31817 36594
rect 32232 36290 32536 36594
rect 32951 36290 33255 36594
rect 33670 36290 33974 36594
rect 34389 36290 34693 36594
rect 35108 36290 35412 36594
rect 35827 36290 36131 36594
rect 36546 36290 36850 36594
rect 26351 33230 26655 33534
rect 27070 33230 27374 33534
rect 27789 33230 28093 33534
rect 28508 33230 28812 33534
rect 29227 33230 29531 33534
rect 29946 33230 30250 33534
rect 30665 33230 30969 33534
rect 31384 33230 31688 33534
rect 32103 33230 32407 33534
rect 32822 33230 33126 33534
rect 33799 33230 34103 33534
rect 34518 33230 34822 33534
rect 35237 33230 35541 33534
rect 35956 33230 36260 33534
rect 36675 33230 36979 33534
rect 37394 33230 37698 33534
rect 38113 33230 38417 33534
rect 38832 33230 39136 33534
rect 39551 33230 39855 33534
rect 40270 33230 40574 33534
rect 26351 32530 26655 32834
rect 27070 32530 27374 32834
rect 27789 32530 28093 32834
rect 28508 32530 28812 32834
rect 29227 32530 29531 32834
rect 29946 32530 30250 32834
rect 30665 32530 30969 32834
rect 31384 32530 31688 32834
rect 32103 32530 32407 32834
rect 32822 32530 33126 32834
rect 33799 32530 34103 32834
rect 34518 32530 34822 32834
rect 35237 32530 35541 32834
rect 35956 32530 36260 32834
rect 36675 32530 36979 32834
rect 37394 32530 37698 32834
rect 38113 32530 38417 32834
rect 38832 32530 39136 32834
rect 39551 32530 39855 32834
rect 40270 32530 40574 32834
rect 30075 29470 30379 29774
rect 30794 29470 31098 29774
rect 31513 29470 31817 29774
rect 32232 29470 32536 29774
rect 32951 29470 33255 29774
rect 33670 29470 33974 29774
rect 34389 29470 34693 29774
rect 35108 29470 35412 29774
rect 35827 29470 36131 29774
rect 36546 29470 36850 29774
rect 30075 28770 30379 29074
rect 30794 28770 31098 29074
rect 31513 28770 31817 29074
rect 32232 28770 32536 29074
rect 32951 28770 33255 29074
rect 33670 28770 33974 29074
rect 34389 28770 34693 29074
rect 35108 28770 35412 29074
rect 35827 28770 36131 29074
rect 36546 28770 36850 29074
rect 30075 25710 30379 26014
rect 30794 25710 31098 26014
rect 31513 25710 31817 26014
rect 32232 25710 32536 26014
rect 32951 25710 33255 26014
rect 33670 25710 33974 26014
rect 34389 25710 34693 26014
rect 35108 25710 35412 26014
rect 35827 25710 36131 26014
rect 36546 25710 36850 26014
rect 30075 25010 30379 25314
rect 30794 25010 31098 25314
rect 31513 25010 31817 25314
rect 32232 25010 32536 25314
rect 32951 25010 33255 25314
rect 33670 25010 33974 25314
rect 34389 25010 34693 25314
rect 35108 25010 35412 25314
rect 35827 25010 36131 25314
rect 36546 25010 36850 25314
<< metal4 >>
rect 900 55670 2532 56576
rect 900 54154 958 55670
rect 2474 54154 2532 55670
rect 900 50864 2532 54154
rect 900 50800 924 50864
rect 988 50800 1004 50864
rect 1068 50800 1084 50864
rect 1148 50800 1164 50864
rect 1228 50800 1244 50864
rect 1308 50800 1324 50864
rect 1388 50800 1404 50864
rect 1468 50800 1484 50864
rect 1548 50800 1564 50864
rect 1628 50800 1644 50864
rect 1708 50800 1724 50864
rect 1788 50800 1804 50864
rect 1868 50800 1884 50864
rect 1948 50800 1964 50864
rect 2028 50800 2044 50864
rect 2108 50800 2124 50864
rect 2188 50800 2204 50864
rect 2268 50800 2284 50864
rect 2348 50800 2364 50864
rect 2428 50800 2444 50864
rect 2508 50800 2532 50864
rect 900 47104 2532 50800
rect 900 47040 924 47104
rect 988 47040 1004 47104
rect 1068 47040 1084 47104
rect 1148 47040 1164 47104
rect 1228 47040 1244 47104
rect 1308 47040 1324 47104
rect 1388 47040 1404 47104
rect 1468 47040 1484 47104
rect 1548 47040 1564 47104
rect 1628 47040 1644 47104
rect 1708 47040 1724 47104
rect 1788 47040 1804 47104
rect 1868 47040 1884 47104
rect 1948 47040 1964 47104
rect 2028 47040 2044 47104
rect 2108 47040 2124 47104
rect 2188 47040 2204 47104
rect 2268 47040 2284 47104
rect 2348 47040 2364 47104
rect 2428 47040 2444 47104
rect 2508 47040 2532 47104
rect 900 43344 2532 47040
rect 900 43280 924 43344
rect 988 43280 1004 43344
rect 1068 43280 1084 43344
rect 1148 43280 1164 43344
rect 1228 43280 1244 43344
rect 1308 43280 1324 43344
rect 1388 43280 1404 43344
rect 1468 43280 1484 43344
rect 1548 43280 1564 43344
rect 1628 43280 1644 43344
rect 1708 43280 1724 43344
rect 1788 43280 1804 43344
rect 1868 43280 1884 43344
rect 1948 43280 1964 43344
rect 2028 43280 2044 43344
rect 2108 43280 2124 43344
rect 2188 43280 2204 43344
rect 2268 43280 2284 43344
rect 2348 43280 2364 43344
rect 2428 43280 2444 43344
rect 2508 43280 2532 43344
rect 900 39584 2532 43280
rect 900 39520 924 39584
rect 988 39520 1004 39584
rect 1068 39520 1084 39584
rect 1148 39520 1164 39584
rect 1228 39520 1244 39584
rect 1308 39520 1324 39584
rect 1388 39520 1404 39584
rect 1468 39520 1484 39584
rect 1548 39520 1564 39584
rect 1628 39520 1644 39584
rect 1708 39520 1724 39584
rect 1788 39520 1804 39584
rect 1868 39520 1884 39584
rect 1948 39520 1964 39584
rect 2028 39520 2044 39584
rect 2108 39520 2124 39584
rect 2188 39520 2204 39584
rect 2268 39520 2284 39584
rect 2348 39520 2364 39584
rect 2428 39520 2444 39584
rect 2508 39520 2532 39584
rect 900 35824 2532 39520
rect 900 35760 924 35824
rect 988 35760 1004 35824
rect 1068 35760 1084 35824
rect 1148 35760 1164 35824
rect 1228 35760 1244 35824
rect 1308 35760 1324 35824
rect 1388 35760 1404 35824
rect 1468 35760 1484 35824
rect 1548 35760 1564 35824
rect 1628 35760 1644 35824
rect 1708 35760 1724 35824
rect 1788 35760 1804 35824
rect 1868 35760 1884 35824
rect 1948 35760 1964 35824
rect 2028 35760 2044 35824
rect 2108 35760 2124 35824
rect 2188 35760 2204 35824
rect 2268 35760 2284 35824
rect 2348 35760 2364 35824
rect 2428 35760 2444 35824
rect 2508 35760 2532 35824
rect 900 32064 2532 35760
rect 900 32000 924 32064
rect 988 32000 1004 32064
rect 1068 32000 1084 32064
rect 1148 32000 1164 32064
rect 1228 32000 1244 32064
rect 1308 32000 1324 32064
rect 1388 32000 1404 32064
rect 1468 32000 1484 32064
rect 1548 32000 1564 32064
rect 1628 32000 1644 32064
rect 1708 32000 1724 32064
rect 1788 32000 1804 32064
rect 1868 32000 1884 32064
rect 1948 32000 1964 32064
rect 2028 32000 2044 32064
rect 2108 32000 2124 32064
rect 2188 32000 2204 32064
rect 2268 32000 2284 32064
rect 2348 32000 2364 32064
rect 2428 32000 2444 32064
rect 2508 32000 2532 32064
rect 900 28304 2532 32000
rect 900 28240 924 28304
rect 988 28240 1004 28304
rect 1068 28240 1084 28304
rect 1148 28240 1164 28304
rect 1228 28240 1244 28304
rect 1308 28240 1324 28304
rect 1388 28240 1404 28304
rect 1468 28240 1484 28304
rect 1548 28240 1564 28304
rect 1628 28240 1644 28304
rect 1708 28240 1724 28304
rect 1788 28240 1804 28304
rect 1868 28240 1884 28304
rect 1948 28240 1964 28304
rect 2028 28240 2044 28304
rect 2108 28240 2124 28304
rect 2188 28240 2204 28304
rect 2268 28240 2284 28304
rect 2348 28240 2364 28304
rect 2428 28240 2444 28304
rect 2508 28240 2532 28304
rect 900 24544 2532 28240
rect 900 24480 924 24544
rect 988 24480 1004 24544
rect 1068 24480 1084 24544
rect 1148 24480 1164 24544
rect 1228 24480 1244 24544
rect 1308 24480 1324 24544
rect 1388 24480 1404 24544
rect 1468 24480 1484 24544
rect 1548 24480 1564 24544
rect 1628 24480 1644 24544
rect 1708 24480 1724 24544
rect 1788 24480 1804 24544
rect 1868 24480 1884 24544
rect 1948 24480 1964 24544
rect 2028 24480 2044 24544
rect 2108 24480 2124 24544
rect 2188 24480 2204 24544
rect 2268 24480 2284 24544
rect 2348 24480 2364 24544
rect 2428 24480 2444 24544
rect 2508 24480 2532 24544
rect 900 20784 2532 24480
rect 900 20720 924 20784
rect 988 20720 1004 20784
rect 1068 20720 1084 20784
rect 1148 20720 1164 20784
rect 1228 20720 1244 20784
rect 1308 20720 1324 20784
rect 1388 20720 1404 20784
rect 1468 20720 1484 20784
rect 1548 20720 1564 20784
rect 1628 20720 1644 20784
rect 1708 20720 1724 20784
rect 1788 20720 1804 20784
rect 1868 20720 1884 20784
rect 1948 20720 1964 20784
rect 2028 20720 2044 20784
rect 2108 20720 2124 20784
rect 2188 20720 2204 20784
rect 2268 20720 2284 20784
rect 2348 20720 2364 20784
rect 2428 20720 2444 20784
rect 2508 20720 2532 20784
rect 900 17024 2532 20720
rect 900 16960 924 17024
rect 988 16960 1004 17024
rect 1068 16960 1084 17024
rect 1148 16960 1164 17024
rect 1228 16960 1244 17024
rect 1308 16960 1324 17024
rect 1388 16960 1404 17024
rect 1468 16960 1484 17024
rect 1548 16960 1564 17024
rect 1628 16960 1644 17024
rect 1708 16960 1724 17024
rect 1788 16960 1804 17024
rect 1868 16960 1884 17024
rect 1948 16960 1964 17024
rect 2028 16960 2044 17024
rect 2108 16960 2124 17024
rect 2188 16960 2204 17024
rect 2268 16960 2284 17024
rect 2348 16960 2364 17024
rect 2428 16960 2444 17024
rect 2508 16960 2532 17024
rect 900 13264 2532 16960
rect 900 13200 924 13264
rect 988 13200 1004 13264
rect 1068 13200 1084 13264
rect 1148 13200 1164 13264
rect 1228 13200 1244 13264
rect 1308 13200 1324 13264
rect 1388 13200 1404 13264
rect 1468 13200 1484 13264
rect 1548 13200 1564 13264
rect 1628 13200 1644 13264
rect 1708 13200 1724 13264
rect 1788 13200 1804 13264
rect 1868 13200 1884 13264
rect 1948 13200 1964 13264
rect 2028 13200 2044 13264
rect 2108 13200 2124 13264
rect 2188 13200 2204 13264
rect 2268 13200 2284 13264
rect 2348 13200 2364 13264
rect 2428 13200 2444 13264
rect 2508 13200 2532 13264
rect 900 9504 2532 13200
rect 900 9440 924 9504
rect 988 9440 1004 9504
rect 1068 9440 1084 9504
rect 1148 9440 1164 9504
rect 1228 9440 1244 9504
rect 1308 9440 1324 9504
rect 1388 9440 1404 9504
rect 1468 9440 1484 9504
rect 1548 9440 1564 9504
rect 1628 9440 1644 9504
rect 1708 9440 1724 9504
rect 1788 9440 1804 9504
rect 1868 9440 1884 9504
rect 1948 9440 1964 9504
rect 2028 9440 2044 9504
rect 2108 9440 2124 9504
rect 2188 9440 2204 9504
rect 2268 9440 2284 9504
rect 2348 9440 2364 9504
rect 2428 9440 2444 9504
rect 2508 9440 2532 9504
rect 900 5744 2532 9440
rect 900 5680 924 5744
rect 988 5680 1004 5744
rect 1068 5680 1084 5744
rect 1148 5680 1164 5744
rect 1228 5680 1244 5744
rect 1308 5680 1324 5744
rect 1388 5680 1404 5744
rect 1468 5680 1484 5744
rect 1548 5680 1564 5744
rect 1628 5680 1644 5744
rect 1708 5680 1724 5744
rect 1788 5680 1804 5744
rect 1868 5680 1884 5744
rect 1948 5680 1964 5744
rect 2028 5680 2044 5744
rect 2108 5680 2124 5744
rect 2188 5680 2204 5744
rect 2268 5680 2284 5744
rect 2348 5680 2364 5744
rect 2428 5680 2444 5744
rect 2508 5680 2532 5744
rect 900 2390 2532 5680
rect 900 874 958 2390
rect 2474 874 2532 2390
rect 900 0 2532 874
rect 3348 53222 4980 56576
rect 3348 51706 3406 53222
rect 4922 51706 4980 53222
rect 3348 48984 4980 51706
rect 3348 48920 3372 48984
rect 3436 48920 3452 48984
rect 3516 48920 3532 48984
rect 3596 48920 3612 48984
rect 3676 48920 3692 48984
rect 3756 48920 3772 48984
rect 3836 48920 3852 48984
rect 3916 48920 3932 48984
rect 3996 48920 4012 48984
rect 4076 48920 4092 48984
rect 4156 48920 4172 48984
rect 4236 48920 4252 48984
rect 4316 48920 4332 48984
rect 4396 48920 4412 48984
rect 4476 48920 4492 48984
rect 4556 48920 4572 48984
rect 4636 48920 4652 48984
rect 4716 48920 4732 48984
rect 4796 48920 4812 48984
rect 4876 48920 4892 48984
rect 4956 48920 4980 48984
rect 53456 53222 55088 56576
rect 53456 51706 53514 53222
rect 55030 51706 55088 53222
rect 53456 48984 55088 51706
rect 3348 45224 4980 48920
rect 5674 48904 6596 48964
rect 5674 45304 5734 48904
rect 6536 48710 6596 48904
rect 12988 48904 14048 48964
rect 12988 48710 13048 48904
rect 13988 48710 14048 48904
rect 53456 48920 53480 48984
rect 53544 48920 53560 48984
rect 53624 48920 53640 48984
rect 53704 48920 53720 48984
rect 53784 48920 53800 48984
rect 53864 48920 53880 48984
rect 53944 48920 53960 48984
rect 54024 48920 54040 48984
rect 54104 48920 54120 48984
rect 54184 48920 54200 48984
rect 54264 48920 54280 48984
rect 54344 48920 54360 48984
rect 54424 48920 54440 48984
rect 54504 48920 54520 48984
rect 54584 48920 54600 48984
rect 54664 48920 54680 48984
rect 54744 48920 54760 48984
rect 54824 48920 54840 48984
rect 54904 48920 54920 48984
rect 54984 48920 55000 48984
rect 55064 48920 55088 48984
rect 6516 48694 6612 48710
rect 6516 48630 6532 48694
rect 6596 48630 6612 48694
rect 6516 48614 6612 48630
rect 6056 48583 6376 48602
rect 6056 48574 6378 48583
rect 6056 48270 6065 48574
rect 6369 48270 6378 48574
rect 6056 48261 6378 48270
rect 6516 48550 6532 48614
rect 6596 48550 6612 48614
rect 7235 48694 7331 48710
rect 7235 48630 7251 48694
rect 7315 48630 7331 48694
rect 7235 48614 7331 48630
rect 6776 48583 7096 48602
rect 6516 48534 6612 48550
rect 6516 48470 6532 48534
rect 6596 48470 6612 48534
rect 6516 48454 6612 48470
rect 6516 48390 6532 48454
rect 6596 48390 6612 48454
rect 6516 48374 6612 48390
rect 6516 48310 6532 48374
rect 6596 48310 6612 48374
rect 6516 48294 6612 48310
rect 6056 47883 6376 48261
rect 6516 48230 6532 48294
rect 6596 48230 6612 48294
rect 6775 48574 7097 48583
rect 6775 48270 6784 48574
rect 7088 48270 7097 48574
rect 6775 48261 7097 48270
rect 7235 48550 7251 48614
rect 7315 48550 7331 48614
rect 7954 48694 8050 48710
rect 7954 48630 7970 48694
rect 8034 48630 8050 48694
rect 7954 48614 8050 48630
rect 7496 48583 7816 48602
rect 7235 48534 7331 48550
rect 7235 48470 7251 48534
rect 7315 48470 7331 48534
rect 7235 48454 7331 48470
rect 7235 48390 7251 48454
rect 7315 48390 7331 48454
rect 7235 48374 7331 48390
rect 7235 48310 7251 48374
rect 7315 48310 7331 48374
rect 7235 48294 7331 48310
rect 6516 48214 6612 48230
rect 6516 48150 6532 48214
rect 6596 48150 6612 48214
rect 6516 48134 6612 48150
rect 6516 47994 6612 48010
rect 6516 47930 6532 47994
rect 6596 47930 6612 47994
rect 6516 47914 6612 47930
rect 6056 47874 6378 47883
rect 6056 47570 6065 47874
rect 6369 47570 6378 47874
rect 6056 47561 6378 47570
rect 6516 47850 6532 47914
rect 6596 47850 6612 47914
rect 6776 47883 7096 48261
rect 7235 48230 7251 48294
rect 7315 48230 7331 48294
rect 7494 48574 7816 48583
rect 7494 48270 7503 48574
rect 7807 48270 7816 48574
rect 7494 48261 7816 48270
rect 7235 48214 7331 48230
rect 7235 48150 7251 48214
rect 7315 48150 7331 48214
rect 7235 48134 7331 48150
rect 7235 47994 7331 48010
rect 7235 47930 7251 47994
rect 7315 47930 7331 47994
rect 7235 47914 7331 47930
rect 6516 47834 6612 47850
rect 6516 47770 6532 47834
rect 6596 47770 6612 47834
rect 6516 47754 6612 47770
rect 6516 47690 6532 47754
rect 6596 47690 6612 47754
rect 6516 47674 6612 47690
rect 6516 47610 6532 47674
rect 6596 47610 6612 47674
rect 6516 47594 6612 47610
rect 6056 47322 6376 47561
rect 6516 47530 6532 47594
rect 6596 47530 6612 47594
rect 6775 47874 7097 47883
rect 6775 47570 6784 47874
rect 7088 47570 7097 47874
rect 6775 47561 7097 47570
rect 7235 47850 7251 47914
rect 7315 47850 7331 47914
rect 7496 47883 7816 48261
rect 7954 48550 7970 48614
rect 8034 48550 8050 48614
rect 8673 48694 8769 48710
rect 8673 48630 8689 48694
rect 8753 48630 8769 48694
rect 8673 48614 8769 48630
rect 8216 48583 8536 48602
rect 7954 48534 8050 48550
rect 7954 48470 7970 48534
rect 8034 48470 8050 48534
rect 7954 48454 8050 48470
rect 7954 48390 7970 48454
rect 8034 48390 8050 48454
rect 7954 48374 8050 48390
rect 7954 48310 7970 48374
rect 8034 48310 8050 48374
rect 7954 48294 8050 48310
rect 7954 48230 7970 48294
rect 8034 48230 8050 48294
rect 8213 48574 8536 48583
rect 8213 48270 8222 48574
rect 8526 48270 8536 48574
rect 8213 48261 8536 48270
rect 7954 48214 8050 48230
rect 7954 48150 7970 48214
rect 8034 48150 8050 48214
rect 7954 48134 8050 48150
rect 7235 47834 7331 47850
rect 7235 47770 7251 47834
rect 7315 47770 7331 47834
rect 7235 47754 7331 47770
rect 7235 47690 7251 47754
rect 7315 47690 7331 47754
rect 7235 47674 7331 47690
rect 7235 47610 7251 47674
rect 7315 47610 7331 47674
rect 7235 47594 7331 47610
rect 6516 47514 6612 47530
rect 6516 47450 6532 47514
rect 6596 47450 6612 47514
rect 6516 47434 6612 47450
rect 6776 47322 7096 47561
rect 7235 47530 7251 47594
rect 7315 47530 7331 47594
rect 7494 47874 7816 47883
rect 7494 47570 7503 47874
rect 7807 47570 7816 47874
rect 7494 47561 7816 47570
rect 7235 47514 7331 47530
rect 7235 47450 7251 47514
rect 7315 47450 7331 47514
rect 7235 47434 7331 47450
rect 7496 47322 7816 47561
rect 7954 47994 8050 48010
rect 7954 47930 7970 47994
rect 8034 47930 8050 47994
rect 7954 47914 8050 47930
rect 7954 47850 7970 47914
rect 8034 47850 8050 47914
rect 8216 47883 8536 48261
rect 8673 48550 8689 48614
rect 8753 48550 8769 48614
rect 9392 48694 9488 48710
rect 9392 48630 9408 48694
rect 9472 48630 9488 48694
rect 9392 48614 9488 48630
rect 8936 48583 9256 48602
rect 8673 48534 8769 48550
rect 8673 48470 8689 48534
rect 8753 48470 8769 48534
rect 8673 48454 8769 48470
rect 8673 48390 8689 48454
rect 8753 48390 8769 48454
rect 8673 48374 8769 48390
rect 8673 48310 8689 48374
rect 8753 48310 8769 48374
rect 8673 48294 8769 48310
rect 8673 48230 8689 48294
rect 8753 48230 8769 48294
rect 8932 48574 9256 48583
rect 8932 48270 8941 48574
rect 9245 48270 9256 48574
rect 8932 48261 9256 48270
rect 8673 48214 8769 48230
rect 8673 48150 8689 48214
rect 8753 48150 8769 48214
rect 8673 48134 8769 48150
rect 7954 47834 8050 47850
rect 7954 47770 7970 47834
rect 8034 47770 8050 47834
rect 7954 47754 8050 47770
rect 7954 47690 7970 47754
rect 8034 47690 8050 47754
rect 7954 47674 8050 47690
rect 7954 47610 7970 47674
rect 8034 47610 8050 47674
rect 7954 47594 8050 47610
rect 7954 47530 7970 47594
rect 8034 47530 8050 47594
rect 8213 47874 8536 47883
rect 8213 47570 8222 47874
rect 8526 47570 8536 47874
rect 8213 47561 8536 47570
rect 7954 47514 8050 47530
rect 7954 47450 7970 47514
rect 8034 47450 8050 47514
rect 7954 47434 8050 47450
rect 8216 47322 8536 47561
rect 8673 47994 8769 48010
rect 8673 47930 8689 47994
rect 8753 47930 8769 47994
rect 8673 47914 8769 47930
rect 8673 47850 8689 47914
rect 8753 47850 8769 47914
rect 8936 47883 9256 48261
rect 9392 48550 9408 48614
rect 9472 48550 9488 48614
rect 10111 48694 10207 48710
rect 10111 48630 10127 48694
rect 10191 48630 10207 48694
rect 10111 48614 10207 48630
rect 9656 48583 9976 48602
rect 9392 48534 9488 48550
rect 9392 48470 9408 48534
rect 9472 48470 9488 48534
rect 9392 48454 9488 48470
rect 9392 48390 9408 48454
rect 9472 48390 9488 48454
rect 9392 48374 9488 48390
rect 9392 48310 9408 48374
rect 9472 48310 9488 48374
rect 9392 48294 9488 48310
rect 9392 48230 9408 48294
rect 9472 48230 9488 48294
rect 9651 48574 9976 48583
rect 9651 48270 9660 48574
rect 9964 48270 9976 48574
rect 9651 48261 9976 48270
rect 9392 48214 9488 48230
rect 9392 48150 9408 48214
rect 9472 48150 9488 48214
rect 9392 48134 9488 48150
rect 8673 47834 8769 47850
rect 8673 47770 8689 47834
rect 8753 47770 8769 47834
rect 8673 47754 8769 47770
rect 8673 47690 8689 47754
rect 8753 47690 8769 47754
rect 8673 47674 8769 47690
rect 8673 47610 8689 47674
rect 8753 47610 8769 47674
rect 8673 47594 8769 47610
rect 8673 47530 8689 47594
rect 8753 47530 8769 47594
rect 8932 47874 9256 47883
rect 8932 47570 8941 47874
rect 9245 47570 9256 47874
rect 8932 47561 9256 47570
rect 8673 47514 8769 47530
rect 8673 47450 8689 47514
rect 8753 47450 8769 47514
rect 8673 47434 8769 47450
rect 8936 47322 9256 47561
rect 9392 47994 9488 48010
rect 9392 47930 9408 47994
rect 9472 47930 9488 47994
rect 9392 47914 9488 47930
rect 9392 47850 9408 47914
rect 9472 47850 9488 47914
rect 9656 47883 9976 48261
rect 10111 48550 10127 48614
rect 10191 48550 10207 48614
rect 10830 48694 10926 48710
rect 10830 48630 10846 48694
rect 10910 48630 10926 48694
rect 10830 48614 10926 48630
rect 10376 48583 10696 48602
rect 10111 48534 10207 48550
rect 10111 48470 10127 48534
rect 10191 48470 10207 48534
rect 10111 48454 10207 48470
rect 10111 48390 10127 48454
rect 10191 48390 10207 48454
rect 10111 48374 10207 48390
rect 10111 48310 10127 48374
rect 10191 48310 10207 48374
rect 10111 48294 10207 48310
rect 10111 48230 10127 48294
rect 10191 48230 10207 48294
rect 10370 48574 10696 48583
rect 10370 48270 10379 48574
rect 10683 48270 10696 48574
rect 10370 48261 10696 48270
rect 10111 48214 10207 48230
rect 10111 48150 10127 48214
rect 10191 48150 10207 48214
rect 10111 48134 10207 48150
rect 9392 47834 9488 47850
rect 9392 47770 9408 47834
rect 9472 47770 9488 47834
rect 9392 47754 9488 47770
rect 9392 47690 9408 47754
rect 9472 47690 9488 47754
rect 9392 47674 9488 47690
rect 9392 47610 9408 47674
rect 9472 47610 9488 47674
rect 9392 47594 9488 47610
rect 9392 47530 9408 47594
rect 9472 47530 9488 47594
rect 9651 47874 9976 47883
rect 9651 47570 9660 47874
rect 9964 47570 9976 47874
rect 9651 47561 9976 47570
rect 9392 47514 9488 47530
rect 9392 47450 9408 47514
rect 9472 47450 9488 47514
rect 9392 47434 9488 47450
rect 9656 47322 9976 47561
rect 10111 47994 10207 48010
rect 10111 47930 10127 47994
rect 10191 47930 10207 47994
rect 10111 47914 10207 47930
rect 10111 47850 10127 47914
rect 10191 47850 10207 47914
rect 10376 47883 10696 48261
rect 10830 48550 10846 48614
rect 10910 48550 10926 48614
rect 11549 48694 11645 48710
rect 11549 48630 11565 48694
rect 11629 48630 11645 48694
rect 11549 48614 11645 48630
rect 11096 48583 11416 48602
rect 10830 48534 10926 48550
rect 10830 48470 10846 48534
rect 10910 48470 10926 48534
rect 10830 48454 10926 48470
rect 10830 48390 10846 48454
rect 10910 48390 10926 48454
rect 10830 48374 10926 48390
rect 10830 48310 10846 48374
rect 10910 48310 10926 48374
rect 10830 48294 10926 48310
rect 10830 48230 10846 48294
rect 10910 48230 10926 48294
rect 11089 48574 11416 48583
rect 11089 48270 11098 48574
rect 11402 48270 11416 48574
rect 11089 48261 11416 48270
rect 10830 48214 10926 48230
rect 10830 48150 10846 48214
rect 10910 48150 10926 48214
rect 10830 48134 10926 48150
rect 10111 47834 10207 47850
rect 10111 47770 10127 47834
rect 10191 47770 10207 47834
rect 10111 47754 10207 47770
rect 10111 47690 10127 47754
rect 10191 47690 10207 47754
rect 10111 47674 10207 47690
rect 10111 47610 10127 47674
rect 10191 47610 10207 47674
rect 10111 47594 10207 47610
rect 10111 47530 10127 47594
rect 10191 47530 10207 47594
rect 10370 47874 10696 47883
rect 10370 47570 10379 47874
rect 10683 47570 10696 47874
rect 10370 47561 10696 47570
rect 10111 47514 10207 47530
rect 10111 47450 10127 47514
rect 10191 47450 10207 47514
rect 10111 47434 10207 47450
rect 10376 47322 10696 47561
rect 10830 47994 10926 48010
rect 10830 47930 10846 47994
rect 10910 47930 10926 47994
rect 10830 47914 10926 47930
rect 10830 47850 10846 47914
rect 10910 47850 10926 47914
rect 11096 47883 11416 48261
rect 11549 48550 11565 48614
rect 11629 48550 11645 48614
rect 12268 48694 12364 48710
rect 12268 48630 12284 48694
rect 12348 48630 12364 48694
rect 12268 48614 12364 48630
rect 11816 48583 12136 48602
rect 11549 48534 11645 48550
rect 11549 48470 11565 48534
rect 11629 48470 11645 48534
rect 11549 48454 11645 48470
rect 11549 48390 11565 48454
rect 11629 48390 11645 48454
rect 11549 48374 11645 48390
rect 11549 48310 11565 48374
rect 11629 48310 11645 48374
rect 11549 48294 11645 48310
rect 11549 48230 11565 48294
rect 11629 48230 11645 48294
rect 11808 48574 12136 48583
rect 11808 48270 11817 48574
rect 12121 48270 12136 48574
rect 11808 48261 12136 48270
rect 11549 48214 11645 48230
rect 11549 48150 11565 48214
rect 11629 48150 11645 48214
rect 11549 48134 11645 48150
rect 10830 47834 10926 47850
rect 10830 47770 10846 47834
rect 10910 47770 10926 47834
rect 10830 47754 10926 47770
rect 10830 47690 10846 47754
rect 10910 47690 10926 47754
rect 10830 47674 10926 47690
rect 10830 47610 10846 47674
rect 10910 47610 10926 47674
rect 10830 47594 10926 47610
rect 10830 47530 10846 47594
rect 10910 47530 10926 47594
rect 11089 47874 11416 47883
rect 11089 47570 11098 47874
rect 11402 47570 11416 47874
rect 11089 47561 11416 47570
rect 10830 47514 10926 47530
rect 10830 47450 10846 47514
rect 10910 47450 10926 47514
rect 10830 47434 10926 47450
rect 11096 47322 11416 47561
rect 11549 47994 11645 48010
rect 11549 47930 11565 47994
rect 11629 47930 11645 47994
rect 11549 47914 11645 47930
rect 11549 47850 11565 47914
rect 11629 47850 11645 47914
rect 11816 47883 12136 48261
rect 12268 48550 12284 48614
rect 12348 48550 12364 48614
rect 12987 48694 13083 48710
rect 12987 48630 13003 48694
rect 13067 48630 13083 48694
rect 12987 48614 13083 48630
rect 12536 48583 12856 48602
rect 12268 48534 12364 48550
rect 12268 48470 12284 48534
rect 12348 48470 12364 48534
rect 12268 48454 12364 48470
rect 12268 48390 12284 48454
rect 12348 48390 12364 48454
rect 12268 48374 12364 48390
rect 12268 48310 12284 48374
rect 12348 48310 12364 48374
rect 12268 48294 12364 48310
rect 12268 48230 12284 48294
rect 12348 48230 12364 48294
rect 12527 48574 12856 48583
rect 12527 48270 12536 48574
rect 12840 48270 12856 48574
rect 12527 48261 12856 48270
rect 12268 48214 12364 48230
rect 12268 48150 12284 48214
rect 12348 48150 12364 48214
rect 12268 48134 12364 48150
rect 11549 47834 11645 47850
rect 11549 47770 11565 47834
rect 11629 47770 11645 47834
rect 11549 47754 11645 47770
rect 11549 47690 11565 47754
rect 11629 47690 11645 47754
rect 11549 47674 11645 47690
rect 11549 47610 11565 47674
rect 11629 47610 11645 47674
rect 11549 47594 11645 47610
rect 11549 47530 11565 47594
rect 11629 47530 11645 47594
rect 11808 47874 12136 47883
rect 11808 47570 11817 47874
rect 12121 47570 12136 47874
rect 11808 47561 12136 47570
rect 11549 47514 11645 47530
rect 11549 47450 11565 47514
rect 11629 47450 11645 47514
rect 11549 47434 11645 47450
rect 11816 47322 12136 47561
rect 12268 47994 12364 48010
rect 12268 47930 12284 47994
rect 12348 47930 12364 47994
rect 12268 47914 12364 47930
rect 12268 47850 12284 47914
rect 12348 47850 12364 47914
rect 12536 47883 12856 48261
rect 12987 48550 13003 48614
rect 13067 48550 13083 48614
rect 13964 48694 14060 48710
rect 13964 48630 13980 48694
rect 14044 48630 14060 48694
rect 13964 48614 14060 48630
rect 12987 48534 13083 48550
rect 12987 48470 13003 48534
rect 13067 48470 13083 48534
rect 12987 48454 13083 48470
rect 12987 48390 13003 48454
rect 13067 48390 13083 48454
rect 12987 48374 13083 48390
rect 12987 48310 13003 48374
rect 13067 48310 13083 48374
rect 12987 48294 13083 48310
rect 12987 48230 13003 48294
rect 13067 48230 13083 48294
rect 12987 48214 13083 48230
rect 12987 48150 13003 48214
rect 13067 48150 13083 48214
rect 12987 48134 13083 48150
rect 13504 48583 13824 48602
rect 13504 48574 13826 48583
rect 13504 48270 13513 48574
rect 13817 48270 13826 48574
rect 13504 48261 13826 48270
rect 13964 48550 13980 48614
rect 14044 48550 14060 48614
rect 14683 48694 14779 48710
rect 14683 48630 14699 48694
rect 14763 48630 14779 48694
rect 14683 48614 14779 48630
rect 14224 48583 14544 48602
rect 13964 48534 14060 48550
rect 13964 48470 13980 48534
rect 14044 48470 14060 48534
rect 13964 48454 14060 48470
rect 13964 48390 13980 48454
rect 14044 48390 14060 48454
rect 13964 48374 14060 48390
rect 13964 48310 13980 48374
rect 14044 48310 14060 48374
rect 13964 48294 14060 48310
rect 12268 47834 12364 47850
rect 12268 47770 12284 47834
rect 12348 47770 12364 47834
rect 12268 47754 12364 47770
rect 12268 47690 12284 47754
rect 12348 47690 12364 47754
rect 12268 47674 12364 47690
rect 12268 47610 12284 47674
rect 12348 47610 12364 47674
rect 12268 47594 12364 47610
rect 12268 47530 12284 47594
rect 12348 47530 12364 47594
rect 12527 47874 12856 47883
rect 12527 47570 12536 47874
rect 12840 47570 12856 47874
rect 12527 47561 12856 47570
rect 12268 47514 12364 47530
rect 12268 47450 12284 47514
rect 12348 47450 12364 47514
rect 12268 47434 12364 47450
rect 12536 47322 12856 47561
rect 12987 47994 13083 48010
rect 12987 47930 13003 47994
rect 13067 47930 13083 47994
rect 12987 47914 13083 47930
rect 12987 47850 13003 47914
rect 13067 47850 13083 47914
rect 12987 47834 13083 47850
rect 12987 47770 13003 47834
rect 13067 47770 13083 47834
rect 12987 47754 13083 47770
rect 12987 47690 13003 47754
rect 13067 47690 13083 47754
rect 12987 47674 13083 47690
rect 12987 47610 13003 47674
rect 13067 47610 13083 47674
rect 12987 47594 13083 47610
rect 12987 47530 13003 47594
rect 13067 47530 13083 47594
rect 12987 47514 13083 47530
rect 12987 47450 13003 47514
rect 13067 47450 13083 47514
rect 12987 47434 13083 47450
rect 13504 47883 13824 48261
rect 13964 48230 13980 48294
rect 14044 48230 14060 48294
rect 14223 48574 14545 48583
rect 14223 48270 14232 48574
rect 14536 48270 14545 48574
rect 14223 48261 14545 48270
rect 14683 48550 14699 48614
rect 14763 48550 14779 48614
rect 15402 48694 15498 48710
rect 15402 48630 15418 48694
rect 15482 48630 15498 48694
rect 15402 48614 15498 48630
rect 14944 48583 15264 48602
rect 14683 48534 14779 48550
rect 14683 48470 14699 48534
rect 14763 48470 14779 48534
rect 14683 48454 14779 48470
rect 14683 48390 14699 48454
rect 14763 48390 14779 48454
rect 14683 48374 14779 48390
rect 14683 48310 14699 48374
rect 14763 48310 14779 48374
rect 14683 48294 14779 48310
rect 13964 48214 14060 48230
rect 13964 48150 13980 48214
rect 14044 48150 14060 48214
rect 13964 48134 14060 48150
rect 13964 47994 14060 48010
rect 13964 47930 13980 47994
rect 14044 47930 14060 47994
rect 13964 47914 14060 47930
rect 13504 47874 13826 47883
rect 13504 47570 13513 47874
rect 13817 47570 13826 47874
rect 13504 47561 13826 47570
rect 13964 47850 13980 47914
rect 14044 47850 14060 47914
rect 14224 47883 14544 48261
rect 14683 48230 14699 48294
rect 14763 48230 14779 48294
rect 14942 48574 15264 48583
rect 14942 48270 14951 48574
rect 15255 48270 15264 48574
rect 14942 48261 15264 48270
rect 14683 48214 14779 48230
rect 14683 48150 14699 48214
rect 14763 48150 14779 48214
rect 14683 48134 14779 48150
rect 14683 47994 14779 48010
rect 14683 47930 14699 47994
rect 14763 47930 14779 47994
rect 14683 47914 14779 47930
rect 13964 47834 14060 47850
rect 13964 47770 13980 47834
rect 14044 47770 14060 47834
rect 13964 47754 14060 47770
rect 13964 47690 13980 47754
rect 14044 47690 14060 47754
rect 13964 47674 14060 47690
rect 13964 47610 13980 47674
rect 14044 47610 14060 47674
rect 13964 47594 14060 47610
rect 13504 47322 13824 47561
rect 13964 47530 13980 47594
rect 14044 47530 14060 47594
rect 14223 47874 14545 47883
rect 14223 47570 14232 47874
rect 14536 47570 14545 47874
rect 14223 47561 14545 47570
rect 14683 47850 14699 47914
rect 14763 47850 14779 47914
rect 14944 47883 15264 48261
rect 15402 48550 15418 48614
rect 15482 48550 15498 48614
rect 16121 48694 16217 48710
rect 16121 48630 16137 48694
rect 16201 48630 16217 48694
rect 16121 48614 16217 48630
rect 15664 48583 15984 48602
rect 15402 48534 15498 48550
rect 15402 48470 15418 48534
rect 15482 48470 15498 48534
rect 15402 48454 15498 48470
rect 15402 48390 15418 48454
rect 15482 48390 15498 48454
rect 15402 48374 15498 48390
rect 15402 48310 15418 48374
rect 15482 48310 15498 48374
rect 15402 48294 15498 48310
rect 15402 48230 15418 48294
rect 15482 48230 15498 48294
rect 15661 48574 15984 48583
rect 15661 48270 15670 48574
rect 15974 48270 15984 48574
rect 15661 48261 15984 48270
rect 15402 48214 15498 48230
rect 15402 48150 15418 48214
rect 15482 48150 15498 48214
rect 15402 48134 15498 48150
rect 14683 47834 14779 47850
rect 14683 47770 14699 47834
rect 14763 47770 14779 47834
rect 14683 47754 14779 47770
rect 14683 47690 14699 47754
rect 14763 47690 14779 47754
rect 14683 47674 14779 47690
rect 14683 47610 14699 47674
rect 14763 47610 14779 47674
rect 14683 47594 14779 47610
rect 13964 47514 14060 47530
rect 13964 47450 13980 47514
rect 14044 47450 14060 47514
rect 13964 47434 14060 47450
rect 14224 47322 14544 47561
rect 14683 47530 14699 47594
rect 14763 47530 14779 47594
rect 14942 47874 15264 47883
rect 14942 47570 14951 47874
rect 15255 47570 15264 47874
rect 14942 47561 15264 47570
rect 14683 47514 14779 47530
rect 14683 47450 14699 47514
rect 14763 47450 14779 47514
rect 14683 47434 14779 47450
rect 14944 47322 15264 47561
rect 15402 47994 15498 48010
rect 15402 47930 15418 47994
rect 15482 47930 15498 47994
rect 15402 47914 15498 47930
rect 15402 47850 15418 47914
rect 15482 47850 15498 47914
rect 15664 47883 15984 48261
rect 16121 48550 16137 48614
rect 16201 48550 16217 48614
rect 16840 48694 16936 48710
rect 16840 48630 16856 48694
rect 16920 48630 16936 48694
rect 16840 48614 16936 48630
rect 16384 48583 16704 48602
rect 16121 48534 16217 48550
rect 16121 48470 16137 48534
rect 16201 48470 16217 48534
rect 16121 48454 16217 48470
rect 16121 48390 16137 48454
rect 16201 48390 16217 48454
rect 16121 48374 16217 48390
rect 16121 48310 16137 48374
rect 16201 48310 16217 48374
rect 16121 48294 16217 48310
rect 16121 48230 16137 48294
rect 16201 48230 16217 48294
rect 16380 48574 16704 48583
rect 16380 48270 16389 48574
rect 16693 48270 16704 48574
rect 16380 48261 16704 48270
rect 16121 48214 16217 48230
rect 16121 48150 16137 48214
rect 16201 48150 16217 48214
rect 16121 48134 16217 48150
rect 15402 47834 15498 47850
rect 15402 47770 15418 47834
rect 15482 47770 15498 47834
rect 15402 47754 15498 47770
rect 15402 47690 15418 47754
rect 15482 47690 15498 47754
rect 15402 47674 15498 47690
rect 15402 47610 15418 47674
rect 15482 47610 15498 47674
rect 15402 47594 15498 47610
rect 15402 47530 15418 47594
rect 15482 47530 15498 47594
rect 15661 47874 15984 47883
rect 15661 47570 15670 47874
rect 15974 47570 15984 47874
rect 15661 47561 15984 47570
rect 15402 47514 15498 47530
rect 15402 47450 15418 47514
rect 15482 47450 15498 47514
rect 15402 47434 15498 47450
rect 15664 47322 15984 47561
rect 16121 47994 16217 48010
rect 16121 47930 16137 47994
rect 16201 47930 16217 47994
rect 16121 47914 16217 47930
rect 16121 47850 16137 47914
rect 16201 47850 16217 47914
rect 16384 47883 16704 48261
rect 16840 48550 16856 48614
rect 16920 48550 16936 48614
rect 17559 48694 17655 48710
rect 17559 48630 17575 48694
rect 17639 48630 17655 48694
rect 17559 48614 17655 48630
rect 17104 48583 17424 48602
rect 16840 48534 16936 48550
rect 16840 48470 16856 48534
rect 16920 48470 16936 48534
rect 16840 48454 16936 48470
rect 16840 48390 16856 48454
rect 16920 48390 16936 48454
rect 16840 48374 16936 48390
rect 16840 48310 16856 48374
rect 16920 48310 16936 48374
rect 16840 48294 16936 48310
rect 16840 48230 16856 48294
rect 16920 48230 16936 48294
rect 17099 48574 17424 48583
rect 17099 48270 17108 48574
rect 17412 48270 17424 48574
rect 17099 48261 17424 48270
rect 16840 48214 16936 48230
rect 16840 48150 16856 48214
rect 16920 48150 16936 48214
rect 16840 48134 16936 48150
rect 16121 47834 16217 47850
rect 16121 47770 16137 47834
rect 16201 47770 16217 47834
rect 16121 47754 16217 47770
rect 16121 47690 16137 47754
rect 16201 47690 16217 47754
rect 16121 47674 16217 47690
rect 16121 47610 16137 47674
rect 16201 47610 16217 47674
rect 16121 47594 16217 47610
rect 16121 47530 16137 47594
rect 16201 47530 16217 47594
rect 16380 47874 16704 47883
rect 16380 47570 16389 47874
rect 16693 47570 16704 47874
rect 16380 47561 16704 47570
rect 16121 47514 16217 47530
rect 16121 47450 16137 47514
rect 16201 47450 16217 47514
rect 16121 47434 16217 47450
rect 16384 47322 16704 47561
rect 16840 47994 16936 48010
rect 16840 47930 16856 47994
rect 16920 47930 16936 47994
rect 16840 47914 16936 47930
rect 16840 47850 16856 47914
rect 16920 47850 16936 47914
rect 17104 47883 17424 48261
rect 17559 48550 17575 48614
rect 17639 48550 17655 48614
rect 18278 48694 18374 48710
rect 18278 48630 18294 48694
rect 18358 48630 18374 48694
rect 18278 48614 18374 48630
rect 17824 48583 18144 48602
rect 17559 48534 17655 48550
rect 17559 48470 17575 48534
rect 17639 48470 17655 48534
rect 17559 48454 17655 48470
rect 17559 48390 17575 48454
rect 17639 48390 17655 48454
rect 17559 48374 17655 48390
rect 17559 48310 17575 48374
rect 17639 48310 17655 48374
rect 17559 48294 17655 48310
rect 17559 48230 17575 48294
rect 17639 48230 17655 48294
rect 17818 48574 18144 48583
rect 17818 48270 17827 48574
rect 18131 48270 18144 48574
rect 17818 48261 18144 48270
rect 17559 48214 17655 48230
rect 17559 48150 17575 48214
rect 17639 48150 17655 48214
rect 17559 48134 17655 48150
rect 16840 47834 16936 47850
rect 16840 47770 16856 47834
rect 16920 47770 16936 47834
rect 16840 47754 16936 47770
rect 16840 47690 16856 47754
rect 16920 47690 16936 47754
rect 16840 47674 16936 47690
rect 16840 47610 16856 47674
rect 16920 47610 16936 47674
rect 16840 47594 16936 47610
rect 16840 47530 16856 47594
rect 16920 47530 16936 47594
rect 17099 47874 17424 47883
rect 17099 47570 17108 47874
rect 17412 47570 17424 47874
rect 17099 47561 17424 47570
rect 16840 47514 16936 47530
rect 16840 47450 16856 47514
rect 16920 47450 16936 47514
rect 16840 47434 16936 47450
rect 17104 47322 17424 47561
rect 17559 47994 17655 48010
rect 17559 47930 17575 47994
rect 17639 47930 17655 47994
rect 17559 47914 17655 47930
rect 17559 47850 17575 47914
rect 17639 47850 17655 47914
rect 17824 47883 18144 48261
rect 18278 48550 18294 48614
rect 18358 48550 18374 48614
rect 18997 48694 19093 48710
rect 18997 48630 19013 48694
rect 19077 48630 19093 48694
rect 18997 48614 19093 48630
rect 18544 48583 18864 48602
rect 18278 48534 18374 48550
rect 18278 48470 18294 48534
rect 18358 48470 18374 48534
rect 18278 48454 18374 48470
rect 18278 48390 18294 48454
rect 18358 48390 18374 48454
rect 18278 48374 18374 48390
rect 18278 48310 18294 48374
rect 18358 48310 18374 48374
rect 18278 48294 18374 48310
rect 18278 48230 18294 48294
rect 18358 48230 18374 48294
rect 18537 48574 18864 48583
rect 18537 48270 18546 48574
rect 18850 48270 18864 48574
rect 18537 48261 18864 48270
rect 18278 48214 18374 48230
rect 18278 48150 18294 48214
rect 18358 48150 18374 48214
rect 18278 48134 18374 48150
rect 17559 47834 17655 47850
rect 17559 47770 17575 47834
rect 17639 47770 17655 47834
rect 17559 47754 17655 47770
rect 17559 47690 17575 47754
rect 17639 47690 17655 47754
rect 17559 47674 17655 47690
rect 17559 47610 17575 47674
rect 17639 47610 17655 47674
rect 17559 47594 17655 47610
rect 17559 47530 17575 47594
rect 17639 47530 17655 47594
rect 17818 47874 18144 47883
rect 17818 47570 17827 47874
rect 18131 47570 18144 47874
rect 17818 47561 18144 47570
rect 17559 47514 17655 47530
rect 17559 47450 17575 47514
rect 17639 47450 17655 47514
rect 17559 47434 17655 47450
rect 17824 47322 18144 47561
rect 18278 47994 18374 48010
rect 18278 47930 18294 47994
rect 18358 47930 18374 47994
rect 18278 47914 18374 47930
rect 18278 47850 18294 47914
rect 18358 47850 18374 47914
rect 18544 47883 18864 48261
rect 18997 48550 19013 48614
rect 19077 48550 19093 48614
rect 19716 48694 19812 48710
rect 19716 48630 19732 48694
rect 19796 48630 19812 48694
rect 19716 48614 19812 48630
rect 19264 48583 19584 48602
rect 18997 48534 19093 48550
rect 18997 48470 19013 48534
rect 19077 48470 19093 48534
rect 18997 48454 19093 48470
rect 18997 48390 19013 48454
rect 19077 48390 19093 48454
rect 18997 48374 19093 48390
rect 18997 48310 19013 48374
rect 19077 48310 19093 48374
rect 18997 48294 19093 48310
rect 18997 48230 19013 48294
rect 19077 48230 19093 48294
rect 19256 48574 19584 48583
rect 19256 48270 19265 48574
rect 19569 48270 19584 48574
rect 19256 48261 19584 48270
rect 18997 48214 19093 48230
rect 18997 48150 19013 48214
rect 19077 48150 19093 48214
rect 18997 48134 19093 48150
rect 18278 47834 18374 47850
rect 18278 47770 18294 47834
rect 18358 47770 18374 47834
rect 18278 47754 18374 47770
rect 18278 47690 18294 47754
rect 18358 47690 18374 47754
rect 18278 47674 18374 47690
rect 18278 47610 18294 47674
rect 18358 47610 18374 47674
rect 18278 47594 18374 47610
rect 18278 47530 18294 47594
rect 18358 47530 18374 47594
rect 18537 47874 18864 47883
rect 18537 47570 18546 47874
rect 18850 47570 18864 47874
rect 18537 47561 18864 47570
rect 18278 47514 18374 47530
rect 18278 47450 18294 47514
rect 18358 47450 18374 47514
rect 18278 47434 18374 47450
rect 18544 47322 18864 47561
rect 18997 47994 19093 48010
rect 18997 47930 19013 47994
rect 19077 47930 19093 47994
rect 18997 47914 19093 47930
rect 18997 47850 19013 47914
rect 19077 47850 19093 47914
rect 19264 47883 19584 48261
rect 19716 48550 19732 48614
rect 19796 48550 19812 48614
rect 20435 48694 20531 48710
rect 20435 48630 20451 48694
rect 20515 48630 20531 48694
rect 20435 48614 20531 48630
rect 19984 48583 20304 48602
rect 19716 48534 19812 48550
rect 19716 48470 19732 48534
rect 19796 48470 19812 48534
rect 19716 48454 19812 48470
rect 19716 48390 19732 48454
rect 19796 48390 19812 48454
rect 19716 48374 19812 48390
rect 19716 48310 19732 48374
rect 19796 48310 19812 48374
rect 19716 48294 19812 48310
rect 19716 48230 19732 48294
rect 19796 48230 19812 48294
rect 19975 48574 20304 48583
rect 19975 48270 19984 48574
rect 20288 48270 20304 48574
rect 19975 48261 20304 48270
rect 19716 48214 19812 48230
rect 19716 48150 19732 48214
rect 19796 48150 19812 48214
rect 19716 48134 19812 48150
rect 18997 47834 19093 47850
rect 18997 47770 19013 47834
rect 19077 47770 19093 47834
rect 18997 47754 19093 47770
rect 18997 47690 19013 47754
rect 19077 47690 19093 47754
rect 18997 47674 19093 47690
rect 18997 47610 19013 47674
rect 19077 47610 19093 47674
rect 18997 47594 19093 47610
rect 18997 47530 19013 47594
rect 19077 47530 19093 47594
rect 19256 47874 19584 47883
rect 19256 47570 19265 47874
rect 19569 47570 19584 47874
rect 19256 47561 19584 47570
rect 18997 47514 19093 47530
rect 18997 47450 19013 47514
rect 19077 47450 19093 47514
rect 18997 47434 19093 47450
rect 19264 47322 19584 47561
rect 19716 47994 19812 48010
rect 19716 47930 19732 47994
rect 19796 47930 19812 47994
rect 19716 47914 19812 47930
rect 19716 47850 19732 47914
rect 19796 47850 19812 47914
rect 19984 47883 20304 48261
rect 20435 48550 20451 48614
rect 20515 48550 20531 48614
rect 20435 48534 20531 48550
rect 20435 48470 20451 48534
rect 20515 48470 20531 48534
rect 20435 48454 20531 48470
rect 20435 48390 20451 48454
rect 20515 48390 20531 48454
rect 20435 48374 20531 48390
rect 20435 48310 20451 48374
rect 20515 48310 20531 48374
rect 20435 48294 20531 48310
rect 20435 48230 20451 48294
rect 20515 48230 20531 48294
rect 20435 48214 20531 48230
rect 20435 48150 20451 48214
rect 20515 48150 20531 48214
rect 20435 48134 20531 48150
rect 19716 47834 19812 47850
rect 19716 47770 19732 47834
rect 19796 47770 19812 47834
rect 19716 47754 19812 47770
rect 19716 47690 19732 47754
rect 19796 47690 19812 47754
rect 19716 47674 19812 47690
rect 19716 47610 19732 47674
rect 19796 47610 19812 47674
rect 19716 47594 19812 47610
rect 19716 47530 19732 47594
rect 19796 47530 19812 47594
rect 19975 47874 20304 47883
rect 19975 47570 19984 47874
rect 20288 47570 20304 47874
rect 19975 47561 20304 47570
rect 19716 47514 19812 47530
rect 19716 47450 19732 47514
rect 19796 47450 19812 47514
rect 19716 47434 19812 47450
rect 19984 47322 20304 47561
rect 20435 47994 20531 48010
rect 20435 47930 20451 47994
rect 20515 47930 20531 47994
rect 20435 47914 20531 47930
rect 20435 47850 20451 47914
rect 20515 47850 20531 47914
rect 20435 47834 20531 47850
rect 20435 47770 20451 47834
rect 20515 47770 20531 47834
rect 20435 47754 20531 47770
rect 20435 47690 20451 47754
rect 20515 47690 20531 47754
rect 20435 47674 20531 47690
rect 20435 47610 20451 47674
rect 20515 47610 20531 47674
rect 20435 47594 20531 47610
rect 20435 47530 20451 47594
rect 20515 47530 20531 47594
rect 20435 47514 20531 47530
rect 20435 47450 20451 47514
rect 20515 47450 20531 47514
rect 20435 47434 20531 47450
rect 5918 47294 13086 47322
rect 5918 47230 5946 47294
rect 6010 47230 6026 47294
rect 6090 47230 13086 47294
rect 5918 47202 13086 47230
rect 13366 47294 20534 47322
rect 13366 47230 13394 47294
rect 13458 47230 13474 47294
rect 13538 47230 20534 47294
rect 13366 47202 20534 47230
rect 12988 47012 13048 47202
rect 13402 47012 13462 47202
rect 17680 47137 17740 47202
rect 17677 47136 17743 47137
rect 17677 47072 17678 47136
rect 17742 47072 17743 47136
rect 17677 47071 17743 47072
rect 12988 46952 13462 47012
rect 5674 45244 6596 45304
rect 3348 45160 3372 45224
rect 3436 45160 3452 45224
rect 3516 45160 3532 45224
rect 3596 45160 3612 45224
rect 3676 45160 3692 45224
rect 3756 45160 3772 45224
rect 3836 45160 3852 45224
rect 3916 45160 3932 45224
rect 3996 45160 4012 45224
rect 4076 45160 4092 45224
rect 4156 45160 4172 45224
rect 4236 45160 4252 45224
rect 4316 45160 4332 45224
rect 4396 45160 4412 45224
rect 4476 45160 4492 45224
rect 4556 45160 4572 45224
rect 4636 45160 4652 45224
rect 4716 45160 4732 45224
rect 4796 45160 4812 45224
rect 4876 45160 4892 45224
rect 4956 45160 4980 45224
rect 3348 41464 4980 45160
rect 6536 44950 6596 45244
rect 53456 45224 55088 48920
rect 53456 45160 53480 45224
rect 53544 45160 53560 45224
rect 53624 45160 53640 45224
rect 53704 45160 53720 45224
rect 53784 45160 53800 45224
rect 53864 45160 53880 45224
rect 53944 45160 53960 45224
rect 54024 45160 54040 45224
rect 54104 45160 54120 45224
rect 54184 45160 54200 45224
rect 54264 45160 54280 45224
rect 54344 45160 54360 45224
rect 54424 45160 54440 45224
rect 54504 45160 54520 45224
rect 54584 45160 54600 45224
rect 54664 45160 54680 45224
rect 54744 45160 54760 45224
rect 54824 45160 54840 45224
rect 54904 45160 54920 45224
rect 54984 45160 55000 45224
rect 55064 45160 55088 45224
rect 6516 44934 6612 44950
rect 6516 44870 6532 44934
rect 6596 44870 6612 44934
rect 6516 44854 6612 44870
rect 6056 44823 6376 44842
rect 6056 44814 6378 44823
rect 6056 44510 6065 44814
rect 6369 44510 6378 44814
rect 6056 44501 6378 44510
rect 6516 44790 6532 44854
rect 6596 44790 6612 44854
rect 7235 44934 7331 44950
rect 7235 44870 7251 44934
rect 7315 44870 7331 44934
rect 7235 44854 7331 44870
rect 6776 44823 7096 44842
rect 6516 44774 6612 44790
rect 6516 44710 6532 44774
rect 6596 44710 6612 44774
rect 6516 44694 6612 44710
rect 6516 44630 6532 44694
rect 6596 44630 6612 44694
rect 6516 44614 6612 44630
rect 6516 44550 6532 44614
rect 6596 44550 6612 44614
rect 6516 44534 6612 44550
rect 6056 44123 6376 44501
rect 6516 44470 6532 44534
rect 6596 44470 6612 44534
rect 6775 44814 7097 44823
rect 6775 44510 6784 44814
rect 7088 44510 7097 44814
rect 6775 44501 7097 44510
rect 7235 44790 7251 44854
rect 7315 44790 7331 44854
rect 7954 44934 8050 44950
rect 7954 44870 7970 44934
rect 8034 44870 8050 44934
rect 7954 44854 8050 44870
rect 7496 44823 7816 44842
rect 7235 44774 7331 44790
rect 7235 44710 7251 44774
rect 7315 44710 7331 44774
rect 7235 44694 7331 44710
rect 7235 44630 7251 44694
rect 7315 44630 7331 44694
rect 7235 44614 7331 44630
rect 7235 44550 7251 44614
rect 7315 44550 7331 44614
rect 7235 44534 7331 44550
rect 6516 44454 6612 44470
rect 6516 44390 6532 44454
rect 6596 44390 6612 44454
rect 6516 44374 6612 44390
rect 6516 44234 6612 44250
rect 6516 44170 6532 44234
rect 6596 44170 6612 44234
rect 6516 44154 6612 44170
rect 6056 44114 6378 44123
rect 6056 43810 6065 44114
rect 6369 43810 6378 44114
rect 6056 43801 6378 43810
rect 6516 44090 6532 44154
rect 6596 44090 6612 44154
rect 6776 44123 7096 44501
rect 7235 44470 7251 44534
rect 7315 44470 7331 44534
rect 7494 44814 7816 44823
rect 7494 44510 7503 44814
rect 7807 44510 7816 44814
rect 7494 44501 7816 44510
rect 7235 44454 7331 44470
rect 7235 44390 7251 44454
rect 7315 44390 7331 44454
rect 7235 44374 7331 44390
rect 7235 44234 7331 44250
rect 7235 44170 7251 44234
rect 7315 44170 7331 44234
rect 7235 44154 7331 44170
rect 6516 44074 6612 44090
rect 6516 44010 6532 44074
rect 6596 44010 6612 44074
rect 6516 43994 6612 44010
rect 6516 43930 6532 43994
rect 6596 43930 6612 43994
rect 6516 43914 6612 43930
rect 6516 43850 6532 43914
rect 6596 43850 6612 43914
rect 6516 43834 6612 43850
rect 6056 43562 6376 43801
rect 6516 43770 6532 43834
rect 6596 43770 6612 43834
rect 6775 44114 7097 44123
rect 6775 43810 6784 44114
rect 7088 43810 7097 44114
rect 6775 43801 7097 43810
rect 7235 44090 7251 44154
rect 7315 44090 7331 44154
rect 7496 44123 7816 44501
rect 7954 44790 7970 44854
rect 8034 44790 8050 44854
rect 8673 44934 8769 44950
rect 8673 44870 8689 44934
rect 8753 44870 8769 44934
rect 8673 44854 8769 44870
rect 8216 44823 8536 44842
rect 7954 44774 8050 44790
rect 7954 44710 7970 44774
rect 8034 44710 8050 44774
rect 7954 44694 8050 44710
rect 7954 44630 7970 44694
rect 8034 44630 8050 44694
rect 7954 44614 8050 44630
rect 7954 44550 7970 44614
rect 8034 44550 8050 44614
rect 7954 44534 8050 44550
rect 7954 44470 7970 44534
rect 8034 44470 8050 44534
rect 8213 44814 8536 44823
rect 8213 44510 8222 44814
rect 8526 44510 8536 44814
rect 8213 44501 8536 44510
rect 7954 44454 8050 44470
rect 7954 44390 7970 44454
rect 8034 44390 8050 44454
rect 7954 44374 8050 44390
rect 7235 44074 7331 44090
rect 7235 44010 7251 44074
rect 7315 44010 7331 44074
rect 7235 43994 7331 44010
rect 7235 43930 7251 43994
rect 7315 43930 7331 43994
rect 7235 43914 7331 43930
rect 7235 43850 7251 43914
rect 7315 43850 7331 43914
rect 7235 43834 7331 43850
rect 6516 43754 6612 43770
rect 6516 43690 6532 43754
rect 6596 43690 6612 43754
rect 6516 43674 6612 43690
rect 6776 43562 7096 43801
rect 7235 43770 7251 43834
rect 7315 43770 7331 43834
rect 7494 44114 7816 44123
rect 7494 43810 7503 44114
rect 7807 43810 7816 44114
rect 7494 43801 7816 43810
rect 7235 43754 7331 43770
rect 7235 43690 7251 43754
rect 7315 43690 7331 43754
rect 7235 43674 7331 43690
rect 7496 43562 7816 43801
rect 7954 44234 8050 44250
rect 7954 44170 7970 44234
rect 8034 44170 8050 44234
rect 7954 44154 8050 44170
rect 7954 44090 7970 44154
rect 8034 44090 8050 44154
rect 8216 44123 8536 44501
rect 8673 44790 8689 44854
rect 8753 44790 8769 44854
rect 9392 44934 9488 44950
rect 9392 44870 9408 44934
rect 9472 44870 9488 44934
rect 9392 44854 9488 44870
rect 8936 44823 9256 44842
rect 8673 44774 8769 44790
rect 8673 44710 8689 44774
rect 8753 44710 8769 44774
rect 8673 44694 8769 44710
rect 8673 44630 8689 44694
rect 8753 44630 8769 44694
rect 8673 44614 8769 44630
rect 8673 44550 8689 44614
rect 8753 44550 8769 44614
rect 8673 44534 8769 44550
rect 8673 44470 8689 44534
rect 8753 44470 8769 44534
rect 8932 44814 9256 44823
rect 8932 44510 8941 44814
rect 9245 44510 9256 44814
rect 8932 44501 9256 44510
rect 8673 44454 8769 44470
rect 8673 44390 8689 44454
rect 8753 44390 8769 44454
rect 8673 44374 8769 44390
rect 7954 44074 8050 44090
rect 7954 44010 7970 44074
rect 8034 44010 8050 44074
rect 7954 43994 8050 44010
rect 7954 43930 7970 43994
rect 8034 43930 8050 43994
rect 7954 43914 8050 43930
rect 7954 43850 7970 43914
rect 8034 43850 8050 43914
rect 7954 43834 8050 43850
rect 7954 43770 7970 43834
rect 8034 43770 8050 43834
rect 8213 44114 8536 44123
rect 8213 43810 8222 44114
rect 8526 43810 8536 44114
rect 8213 43801 8536 43810
rect 7954 43754 8050 43770
rect 7954 43690 7970 43754
rect 8034 43690 8050 43754
rect 7954 43674 8050 43690
rect 8216 43562 8536 43801
rect 8673 44234 8769 44250
rect 8673 44170 8689 44234
rect 8753 44170 8769 44234
rect 8673 44154 8769 44170
rect 8673 44090 8689 44154
rect 8753 44090 8769 44154
rect 8936 44123 9256 44501
rect 9392 44790 9408 44854
rect 9472 44790 9488 44854
rect 10111 44934 10207 44950
rect 10111 44870 10127 44934
rect 10191 44870 10207 44934
rect 10111 44854 10207 44870
rect 9656 44823 9976 44842
rect 9392 44774 9488 44790
rect 9392 44710 9408 44774
rect 9472 44710 9488 44774
rect 9392 44694 9488 44710
rect 9392 44630 9408 44694
rect 9472 44630 9488 44694
rect 9392 44614 9488 44630
rect 9392 44550 9408 44614
rect 9472 44550 9488 44614
rect 9392 44534 9488 44550
rect 9392 44470 9408 44534
rect 9472 44470 9488 44534
rect 9651 44814 9976 44823
rect 9651 44510 9660 44814
rect 9964 44510 9976 44814
rect 9651 44501 9976 44510
rect 9392 44454 9488 44470
rect 9392 44390 9408 44454
rect 9472 44390 9488 44454
rect 9392 44374 9488 44390
rect 8673 44074 8769 44090
rect 8673 44010 8689 44074
rect 8753 44010 8769 44074
rect 8673 43994 8769 44010
rect 8673 43930 8689 43994
rect 8753 43930 8769 43994
rect 8673 43914 8769 43930
rect 8673 43850 8689 43914
rect 8753 43850 8769 43914
rect 8673 43834 8769 43850
rect 8673 43770 8689 43834
rect 8753 43770 8769 43834
rect 8932 44114 9256 44123
rect 8932 43810 8941 44114
rect 9245 43810 9256 44114
rect 8932 43801 9256 43810
rect 8673 43754 8769 43770
rect 8673 43690 8689 43754
rect 8753 43690 8769 43754
rect 8673 43674 8769 43690
rect 8936 43562 9256 43801
rect 9392 44234 9488 44250
rect 9392 44170 9408 44234
rect 9472 44170 9488 44234
rect 9392 44154 9488 44170
rect 9392 44090 9408 44154
rect 9472 44090 9488 44154
rect 9656 44123 9976 44501
rect 10111 44790 10127 44854
rect 10191 44790 10207 44854
rect 10830 44934 10926 44950
rect 10830 44870 10846 44934
rect 10910 44870 10926 44934
rect 10830 44854 10926 44870
rect 10376 44823 10696 44842
rect 10111 44774 10207 44790
rect 10111 44710 10127 44774
rect 10191 44710 10207 44774
rect 10111 44694 10207 44710
rect 10111 44630 10127 44694
rect 10191 44630 10207 44694
rect 10111 44614 10207 44630
rect 10111 44550 10127 44614
rect 10191 44550 10207 44614
rect 10111 44534 10207 44550
rect 10111 44470 10127 44534
rect 10191 44470 10207 44534
rect 10370 44814 10696 44823
rect 10370 44510 10379 44814
rect 10683 44510 10696 44814
rect 10370 44501 10696 44510
rect 10111 44454 10207 44470
rect 10111 44390 10127 44454
rect 10191 44390 10207 44454
rect 10111 44374 10207 44390
rect 9392 44074 9488 44090
rect 9392 44010 9408 44074
rect 9472 44010 9488 44074
rect 9392 43994 9488 44010
rect 9392 43930 9408 43994
rect 9472 43930 9488 43994
rect 9392 43914 9488 43930
rect 9392 43850 9408 43914
rect 9472 43850 9488 43914
rect 9392 43834 9488 43850
rect 9392 43770 9408 43834
rect 9472 43770 9488 43834
rect 9651 44114 9976 44123
rect 9651 43810 9660 44114
rect 9964 43810 9976 44114
rect 9651 43801 9976 43810
rect 9392 43754 9488 43770
rect 9392 43690 9408 43754
rect 9472 43690 9488 43754
rect 9392 43674 9488 43690
rect 9656 43562 9976 43801
rect 10111 44234 10207 44250
rect 10111 44170 10127 44234
rect 10191 44170 10207 44234
rect 10111 44154 10207 44170
rect 10111 44090 10127 44154
rect 10191 44090 10207 44154
rect 10376 44123 10696 44501
rect 10830 44790 10846 44854
rect 10910 44790 10926 44854
rect 11549 44934 11645 44950
rect 11549 44870 11565 44934
rect 11629 44870 11645 44934
rect 11549 44854 11645 44870
rect 11096 44823 11416 44842
rect 10830 44774 10926 44790
rect 10830 44710 10846 44774
rect 10910 44710 10926 44774
rect 10830 44694 10926 44710
rect 10830 44630 10846 44694
rect 10910 44630 10926 44694
rect 10830 44614 10926 44630
rect 10830 44550 10846 44614
rect 10910 44550 10926 44614
rect 10830 44534 10926 44550
rect 10830 44470 10846 44534
rect 10910 44470 10926 44534
rect 11089 44814 11416 44823
rect 11089 44510 11098 44814
rect 11402 44510 11416 44814
rect 11089 44501 11416 44510
rect 10830 44454 10926 44470
rect 10830 44390 10846 44454
rect 10910 44390 10926 44454
rect 10830 44374 10926 44390
rect 10111 44074 10207 44090
rect 10111 44010 10127 44074
rect 10191 44010 10207 44074
rect 10111 43994 10207 44010
rect 10111 43930 10127 43994
rect 10191 43930 10207 43994
rect 10111 43914 10207 43930
rect 10111 43850 10127 43914
rect 10191 43850 10207 43914
rect 10111 43834 10207 43850
rect 10111 43770 10127 43834
rect 10191 43770 10207 43834
rect 10370 44114 10696 44123
rect 10370 43810 10379 44114
rect 10683 43810 10696 44114
rect 10370 43801 10696 43810
rect 10111 43754 10207 43770
rect 10111 43690 10127 43754
rect 10191 43690 10207 43754
rect 10111 43674 10207 43690
rect 10376 43562 10696 43801
rect 10830 44234 10926 44250
rect 10830 44170 10846 44234
rect 10910 44170 10926 44234
rect 10830 44154 10926 44170
rect 10830 44090 10846 44154
rect 10910 44090 10926 44154
rect 11096 44123 11416 44501
rect 11549 44790 11565 44854
rect 11629 44790 11645 44854
rect 12268 44934 12364 44950
rect 12268 44870 12284 44934
rect 12348 44870 12364 44934
rect 12268 44854 12364 44870
rect 11816 44823 12136 44842
rect 11549 44774 11645 44790
rect 11549 44710 11565 44774
rect 11629 44710 11645 44774
rect 11549 44694 11645 44710
rect 11549 44630 11565 44694
rect 11629 44630 11645 44694
rect 11549 44614 11645 44630
rect 11549 44550 11565 44614
rect 11629 44550 11645 44614
rect 11549 44534 11645 44550
rect 11549 44470 11565 44534
rect 11629 44470 11645 44534
rect 11808 44814 12136 44823
rect 11808 44510 11817 44814
rect 12121 44510 12136 44814
rect 11808 44501 12136 44510
rect 11549 44454 11645 44470
rect 11549 44390 11565 44454
rect 11629 44390 11645 44454
rect 11549 44374 11645 44390
rect 10830 44074 10926 44090
rect 10830 44010 10846 44074
rect 10910 44010 10926 44074
rect 10830 43994 10926 44010
rect 10830 43930 10846 43994
rect 10910 43930 10926 43994
rect 10830 43914 10926 43930
rect 10830 43850 10846 43914
rect 10910 43850 10926 43914
rect 10830 43834 10926 43850
rect 10830 43770 10846 43834
rect 10910 43770 10926 43834
rect 11089 44114 11416 44123
rect 11089 43810 11098 44114
rect 11402 43810 11416 44114
rect 11089 43801 11416 43810
rect 10830 43754 10926 43770
rect 10830 43690 10846 43754
rect 10910 43690 10926 43754
rect 10830 43674 10926 43690
rect 11096 43562 11416 43801
rect 11549 44234 11645 44250
rect 11549 44170 11565 44234
rect 11629 44170 11645 44234
rect 11549 44154 11645 44170
rect 11549 44090 11565 44154
rect 11629 44090 11645 44154
rect 11816 44123 12136 44501
rect 12268 44790 12284 44854
rect 12348 44790 12364 44854
rect 12987 44934 13083 44950
rect 12987 44870 13003 44934
rect 13067 44870 13083 44934
rect 12987 44854 13083 44870
rect 12536 44823 12856 44842
rect 12268 44774 12364 44790
rect 12268 44710 12284 44774
rect 12348 44710 12364 44774
rect 12268 44694 12364 44710
rect 12268 44630 12284 44694
rect 12348 44630 12364 44694
rect 12268 44614 12364 44630
rect 12268 44550 12284 44614
rect 12348 44550 12364 44614
rect 12268 44534 12364 44550
rect 12268 44470 12284 44534
rect 12348 44470 12364 44534
rect 12527 44814 12856 44823
rect 12527 44510 12536 44814
rect 12840 44510 12856 44814
rect 12527 44501 12856 44510
rect 12268 44454 12364 44470
rect 12268 44390 12284 44454
rect 12348 44390 12364 44454
rect 12268 44374 12364 44390
rect 11549 44074 11645 44090
rect 11549 44010 11565 44074
rect 11629 44010 11645 44074
rect 11549 43994 11645 44010
rect 11549 43930 11565 43994
rect 11629 43930 11645 43994
rect 11549 43914 11645 43930
rect 11549 43850 11565 43914
rect 11629 43850 11645 43914
rect 11549 43834 11645 43850
rect 11549 43770 11565 43834
rect 11629 43770 11645 43834
rect 11808 44114 12136 44123
rect 11808 43810 11817 44114
rect 12121 43810 12136 44114
rect 11808 43801 12136 43810
rect 11549 43754 11645 43770
rect 11549 43690 11565 43754
rect 11629 43690 11645 43754
rect 11549 43674 11645 43690
rect 11816 43562 12136 43801
rect 12268 44234 12364 44250
rect 12268 44170 12284 44234
rect 12348 44170 12364 44234
rect 12268 44154 12364 44170
rect 12268 44090 12284 44154
rect 12348 44090 12364 44154
rect 12536 44123 12856 44501
rect 12987 44790 13003 44854
rect 13067 44790 13083 44854
rect 12987 44774 13083 44790
rect 12987 44710 13003 44774
rect 13067 44710 13083 44774
rect 12987 44694 13083 44710
rect 12987 44630 13003 44694
rect 13067 44630 13083 44694
rect 12987 44614 13083 44630
rect 12987 44550 13003 44614
rect 13067 44550 13083 44614
rect 12987 44534 13083 44550
rect 12987 44470 13003 44534
rect 13067 44470 13083 44534
rect 12987 44454 13083 44470
rect 12987 44390 13003 44454
rect 13067 44390 13083 44454
rect 12987 44374 13083 44390
rect 12268 44074 12364 44090
rect 12268 44010 12284 44074
rect 12348 44010 12364 44074
rect 12268 43994 12364 44010
rect 12268 43930 12284 43994
rect 12348 43930 12364 43994
rect 12268 43914 12364 43930
rect 12268 43850 12284 43914
rect 12348 43850 12364 43914
rect 12268 43834 12364 43850
rect 12268 43770 12284 43834
rect 12348 43770 12364 43834
rect 12527 44114 12856 44123
rect 12527 43810 12536 44114
rect 12840 43810 12856 44114
rect 12527 43801 12856 43810
rect 12268 43754 12364 43770
rect 12268 43690 12284 43754
rect 12348 43690 12364 43754
rect 12268 43674 12364 43690
rect 12536 43562 12856 43801
rect 12987 44234 13083 44250
rect 12987 44170 13003 44234
rect 13067 44170 13083 44234
rect 12987 44154 13083 44170
rect 12987 44090 13003 44154
rect 13067 44090 13083 44154
rect 12987 44074 13083 44090
rect 12987 44010 13003 44074
rect 13067 44010 13083 44074
rect 12987 43994 13083 44010
rect 12987 43930 13003 43994
rect 13067 43930 13083 43994
rect 12987 43914 13083 43930
rect 12987 43850 13003 43914
rect 13067 43850 13083 43914
rect 12987 43840 13083 43850
rect 13399 43842 13465 43843
rect 13399 43840 13400 43842
rect 12987 43834 13400 43840
rect 12987 43770 13003 43834
rect 13067 43780 13400 43834
rect 13067 43770 13083 43780
rect 13399 43778 13400 43780
rect 13464 43778 13465 43842
rect 13399 43777 13465 43778
rect 12987 43754 13083 43770
rect 12987 43690 13003 43754
rect 13067 43690 13083 43754
rect 12987 43674 13083 43690
rect 5918 43534 13086 43562
rect 5918 43470 5946 43534
rect 6010 43470 6026 43534
rect 6090 43470 13086 43534
rect 5918 43442 13086 43470
rect 3348 41400 3372 41464
rect 3436 41400 3452 41464
rect 3516 41400 3532 41464
rect 3596 41400 3612 41464
rect 3676 41400 3692 41464
rect 3756 41400 3772 41464
rect 3836 41400 3852 41464
rect 3916 41400 3932 41464
rect 3996 41400 4012 41464
rect 4076 41400 4092 41464
rect 4156 41400 4172 41464
rect 4236 41400 4252 41464
rect 4316 41400 4332 41464
rect 4396 41400 4412 41464
rect 4476 41400 4492 41464
rect 4556 41400 4572 41464
rect 4636 41400 4652 41464
rect 4716 41400 4732 41464
rect 4796 41400 4812 41464
rect 4876 41400 4892 41464
rect 4956 41400 4980 41464
rect 3348 37704 4980 41400
rect 6640 41082 6700 43442
rect 8296 43355 8356 43442
rect 8293 43354 8359 43355
rect 8293 43290 8294 43354
rect 8358 43290 8359 43354
rect 8293 43289 8359 43290
rect 6913 41402 6979 41403
rect 6913 41338 6914 41402
rect 6978 41338 6979 41402
rect 6913 41337 6979 41338
rect 6916 41190 6976 41337
rect 13402 41190 13462 43777
rect 53456 41464 55088 45160
rect 22231 41402 22297 41403
rect 22231 41338 22232 41402
rect 22296 41338 22297 41402
rect 22231 41337 22297 41338
rect 53456 41400 53480 41464
rect 53544 41400 53560 41464
rect 53624 41400 53640 41464
rect 53704 41400 53720 41464
rect 53784 41400 53800 41464
rect 53864 41400 53880 41464
rect 53944 41400 53960 41464
rect 54024 41400 54040 41464
rect 54104 41400 54120 41464
rect 54184 41400 54200 41464
rect 54264 41400 54280 41464
rect 54344 41400 54360 41464
rect 54424 41400 54440 41464
rect 54504 41400 54520 41464
rect 54584 41400 54600 41464
rect 54664 41400 54680 41464
rect 54744 41400 54760 41464
rect 54824 41400 54840 41464
rect 54904 41400 54920 41464
rect 54984 41400 55000 41464
rect 55064 41400 55088 41464
rect 22234 41190 22294 41337
rect 6908 41174 7004 41190
rect 6908 41110 6924 41174
rect 6988 41110 7004 41174
rect 6908 41094 7004 41110
rect 6448 41063 6768 41082
rect 6448 41054 6770 41063
rect 6448 40750 6457 41054
rect 6761 40750 6770 41054
rect 6448 40741 6770 40750
rect 6908 41030 6924 41094
rect 6988 41030 7004 41094
rect 7627 41174 7723 41190
rect 7627 41110 7643 41174
rect 7707 41110 7723 41174
rect 7627 41094 7723 41110
rect 7168 41063 7488 41082
rect 6908 41014 7004 41030
rect 6908 40950 6924 41014
rect 6988 40950 7004 41014
rect 6908 40934 7004 40950
rect 6908 40870 6924 40934
rect 6988 40870 7004 40934
rect 6908 40854 7004 40870
rect 6908 40790 6924 40854
rect 6988 40790 7004 40854
rect 6908 40774 7004 40790
rect 6448 40363 6768 40741
rect 6908 40710 6924 40774
rect 6988 40710 7004 40774
rect 7167 41054 7489 41063
rect 7167 40750 7176 41054
rect 7480 40750 7489 41054
rect 7167 40741 7489 40750
rect 7627 41030 7643 41094
rect 7707 41030 7723 41094
rect 8346 41174 8442 41190
rect 8346 41110 8362 41174
rect 8426 41110 8442 41174
rect 8346 41094 8442 41110
rect 7888 41063 8208 41082
rect 7627 41014 7723 41030
rect 7627 40950 7643 41014
rect 7707 40950 7723 41014
rect 7627 40934 7723 40950
rect 7627 40870 7643 40934
rect 7707 40870 7723 40934
rect 7627 40854 7723 40870
rect 7627 40790 7643 40854
rect 7707 40790 7723 40854
rect 7627 40774 7723 40790
rect 6908 40694 7004 40710
rect 6908 40630 6924 40694
rect 6988 40630 7004 40694
rect 6908 40614 7004 40630
rect 6908 40474 7004 40490
rect 6908 40410 6924 40474
rect 6988 40410 7004 40474
rect 6908 40394 7004 40410
rect 6448 40354 6770 40363
rect 6448 40050 6457 40354
rect 6761 40050 6770 40354
rect 6448 40041 6770 40050
rect 6908 40330 6924 40394
rect 6988 40330 7004 40394
rect 7168 40363 7488 40741
rect 7627 40710 7643 40774
rect 7707 40710 7723 40774
rect 7886 41054 8208 41063
rect 7886 40750 7895 41054
rect 8199 40750 8208 41054
rect 7886 40741 8208 40750
rect 7627 40694 7723 40710
rect 7627 40630 7643 40694
rect 7707 40630 7723 40694
rect 7627 40614 7723 40630
rect 7627 40474 7723 40490
rect 7627 40410 7643 40474
rect 7707 40410 7723 40474
rect 7627 40394 7723 40410
rect 6908 40314 7004 40330
rect 6908 40250 6924 40314
rect 6988 40250 7004 40314
rect 6908 40234 7004 40250
rect 6908 40170 6924 40234
rect 6988 40170 7004 40234
rect 6908 40154 7004 40170
rect 6908 40090 6924 40154
rect 6988 40090 7004 40154
rect 6908 40074 7004 40090
rect 6448 39802 6768 40041
rect 6908 40010 6924 40074
rect 6988 40010 7004 40074
rect 7167 40354 7489 40363
rect 7167 40050 7176 40354
rect 7480 40050 7489 40354
rect 7167 40041 7489 40050
rect 7627 40330 7643 40394
rect 7707 40330 7723 40394
rect 7888 40363 8208 40741
rect 8346 41030 8362 41094
rect 8426 41030 8442 41094
rect 9065 41174 9161 41190
rect 9065 41110 9081 41174
rect 9145 41110 9161 41174
rect 9065 41094 9161 41110
rect 8608 41063 8928 41082
rect 8346 41014 8442 41030
rect 8346 40950 8362 41014
rect 8426 40950 8442 41014
rect 8346 40934 8442 40950
rect 8346 40870 8362 40934
rect 8426 40870 8442 40934
rect 8346 40854 8442 40870
rect 8346 40790 8362 40854
rect 8426 40790 8442 40854
rect 8346 40774 8442 40790
rect 8346 40710 8362 40774
rect 8426 40710 8442 40774
rect 8605 41054 8928 41063
rect 8605 40750 8614 41054
rect 8918 40750 8928 41054
rect 8605 40741 8928 40750
rect 8346 40694 8442 40710
rect 8346 40630 8362 40694
rect 8426 40630 8442 40694
rect 8346 40614 8442 40630
rect 7627 40314 7723 40330
rect 7627 40250 7643 40314
rect 7707 40250 7723 40314
rect 7627 40234 7723 40250
rect 7627 40170 7643 40234
rect 7707 40170 7723 40234
rect 7627 40154 7723 40170
rect 7627 40090 7643 40154
rect 7707 40090 7723 40154
rect 7627 40074 7723 40090
rect 6908 39994 7004 40010
rect 6908 39930 6924 39994
rect 6988 39930 7004 39994
rect 6908 39914 7004 39930
rect 7168 39802 7488 40041
rect 7627 40010 7643 40074
rect 7707 40010 7723 40074
rect 7886 40354 8208 40363
rect 7886 40050 7895 40354
rect 8199 40050 8208 40354
rect 7886 40041 8208 40050
rect 7627 39994 7723 40010
rect 7627 39930 7643 39994
rect 7707 39930 7723 39994
rect 7627 39914 7723 39930
rect 7888 39802 8208 40041
rect 8346 40474 8442 40490
rect 8346 40410 8362 40474
rect 8426 40410 8442 40474
rect 8346 40394 8442 40410
rect 8346 40330 8362 40394
rect 8426 40330 8442 40394
rect 8608 40363 8928 40741
rect 9065 41030 9081 41094
rect 9145 41030 9161 41094
rect 9784 41174 9880 41190
rect 9784 41110 9800 41174
rect 9864 41110 9880 41174
rect 9784 41094 9880 41110
rect 9328 41063 9648 41082
rect 9065 41014 9161 41030
rect 9065 40950 9081 41014
rect 9145 40950 9161 41014
rect 9065 40934 9161 40950
rect 9065 40870 9081 40934
rect 9145 40870 9161 40934
rect 9065 40854 9161 40870
rect 9065 40790 9081 40854
rect 9145 40790 9161 40854
rect 9065 40774 9161 40790
rect 9065 40710 9081 40774
rect 9145 40710 9161 40774
rect 9324 41054 9648 41063
rect 9324 40750 9333 41054
rect 9637 40750 9648 41054
rect 9324 40741 9648 40750
rect 9065 40694 9161 40710
rect 9065 40630 9081 40694
rect 9145 40630 9161 40694
rect 9065 40614 9161 40630
rect 8346 40314 8442 40330
rect 8346 40250 8362 40314
rect 8426 40250 8442 40314
rect 8346 40234 8442 40250
rect 8346 40170 8362 40234
rect 8426 40170 8442 40234
rect 8346 40154 8442 40170
rect 8346 40090 8362 40154
rect 8426 40090 8442 40154
rect 8346 40074 8442 40090
rect 8346 40010 8362 40074
rect 8426 40010 8442 40074
rect 8605 40354 8928 40363
rect 8605 40050 8614 40354
rect 8918 40050 8928 40354
rect 8605 40041 8928 40050
rect 8346 39994 8442 40010
rect 8346 39930 8362 39994
rect 8426 39930 8442 39994
rect 8346 39914 8442 39930
rect 8608 39802 8928 40041
rect 9065 40474 9161 40490
rect 9065 40410 9081 40474
rect 9145 40410 9161 40474
rect 9065 40394 9161 40410
rect 9065 40330 9081 40394
rect 9145 40330 9161 40394
rect 9328 40363 9648 40741
rect 9784 41030 9800 41094
rect 9864 41030 9880 41094
rect 10503 41174 10599 41190
rect 10503 41110 10519 41174
rect 10583 41110 10599 41174
rect 10503 41094 10599 41110
rect 10048 41063 10368 41082
rect 9784 41014 9880 41030
rect 9784 40950 9800 41014
rect 9864 40950 9880 41014
rect 9784 40934 9880 40950
rect 9784 40870 9800 40934
rect 9864 40870 9880 40934
rect 9784 40854 9880 40870
rect 9784 40790 9800 40854
rect 9864 40790 9880 40854
rect 9784 40774 9880 40790
rect 9784 40710 9800 40774
rect 9864 40710 9880 40774
rect 10043 41054 10368 41063
rect 10043 40750 10052 41054
rect 10356 40750 10368 41054
rect 10043 40741 10368 40750
rect 9784 40694 9880 40710
rect 9784 40630 9800 40694
rect 9864 40630 9880 40694
rect 9784 40614 9880 40630
rect 9065 40314 9161 40330
rect 9065 40250 9081 40314
rect 9145 40250 9161 40314
rect 9065 40234 9161 40250
rect 9065 40170 9081 40234
rect 9145 40170 9161 40234
rect 9065 40154 9161 40170
rect 9065 40090 9081 40154
rect 9145 40090 9161 40154
rect 9065 40074 9161 40090
rect 9065 40010 9081 40074
rect 9145 40010 9161 40074
rect 9324 40354 9648 40363
rect 9324 40050 9333 40354
rect 9637 40050 9648 40354
rect 9324 40041 9648 40050
rect 9065 39994 9161 40010
rect 9065 39930 9081 39994
rect 9145 39930 9161 39994
rect 9065 39914 9161 39930
rect 9328 39802 9648 40041
rect 9784 40474 9880 40490
rect 9784 40410 9800 40474
rect 9864 40410 9880 40474
rect 9784 40394 9880 40410
rect 9784 40330 9800 40394
rect 9864 40330 9880 40394
rect 10048 40363 10368 40741
rect 10503 41030 10519 41094
rect 10583 41030 10599 41094
rect 11222 41174 11318 41190
rect 11222 41110 11238 41174
rect 11302 41110 11318 41174
rect 11222 41094 11318 41110
rect 10768 41063 11088 41082
rect 10503 41014 10599 41030
rect 10503 40950 10519 41014
rect 10583 40950 10599 41014
rect 10503 40934 10599 40950
rect 10503 40870 10519 40934
rect 10583 40870 10599 40934
rect 10503 40854 10599 40870
rect 10503 40790 10519 40854
rect 10583 40790 10599 40854
rect 10503 40774 10599 40790
rect 10503 40710 10519 40774
rect 10583 40710 10599 40774
rect 10762 41054 11088 41063
rect 10762 40750 10771 41054
rect 11075 40750 11088 41054
rect 10762 40741 11088 40750
rect 10503 40694 10599 40710
rect 10503 40630 10519 40694
rect 10583 40630 10599 40694
rect 10503 40614 10599 40630
rect 9784 40314 9880 40330
rect 9784 40250 9800 40314
rect 9864 40250 9880 40314
rect 9784 40234 9880 40250
rect 9784 40170 9800 40234
rect 9864 40170 9880 40234
rect 9784 40154 9880 40170
rect 9784 40090 9800 40154
rect 9864 40090 9880 40154
rect 9784 40074 9880 40090
rect 9784 40010 9800 40074
rect 9864 40010 9880 40074
rect 10043 40354 10368 40363
rect 10043 40050 10052 40354
rect 10356 40050 10368 40354
rect 10043 40041 10368 40050
rect 9784 39994 9880 40010
rect 9784 39930 9800 39994
rect 9864 39930 9880 39994
rect 9784 39914 9880 39930
rect 10048 39802 10368 40041
rect 10503 40474 10599 40490
rect 10503 40410 10519 40474
rect 10583 40410 10599 40474
rect 10503 40394 10599 40410
rect 10503 40330 10519 40394
rect 10583 40330 10599 40394
rect 10768 40363 11088 40741
rect 11222 41030 11238 41094
rect 11302 41030 11318 41094
rect 11941 41174 12037 41190
rect 11941 41110 11957 41174
rect 12021 41110 12037 41174
rect 11941 41094 12037 41110
rect 11488 41063 11808 41082
rect 11222 41014 11318 41030
rect 11222 40950 11238 41014
rect 11302 40950 11318 41014
rect 11222 40934 11318 40950
rect 11222 40870 11238 40934
rect 11302 40870 11318 40934
rect 11222 40854 11318 40870
rect 11222 40790 11238 40854
rect 11302 40790 11318 40854
rect 11222 40774 11318 40790
rect 11222 40710 11238 40774
rect 11302 40710 11318 40774
rect 11481 41054 11808 41063
rect 11481 40750 11490 41054
rect 11794 40750 11808 41054
rect 11481 40741 11808 40750
rect 11222 40694 11318 40710
rect 11222 40630 11238 40694
rect 11302 40630 11318 40694
rect 11222 40614 11318 40630
rect 10503 40314 10599 40330
rect 10503 40250 10519 40314
rect 10583 40250 10599 40314
rect 10503 40234 10599 40250
rect 10503 40170 10519 40234
rect 10583 40170 10599 40234
rect 10503 40154 10599 40170
rect 10503 40090 10519 40154
rect 10583 40090 10599 40154
rect 10503 40074 10599 40090
rect 10503 40010 10519 40074
rect 10583 40010 10599 40074
rect 10762 40354 11088 40363
rect 10762 40050 10771 40354
rect 11075 40050 11088 40354
rect 10762 40041 11088 40050
rect 10503 39994 10599 40010
rect 10503 39930 10519 39994
rect 10583 39930 10599 39994
rect 10503 39914 10599 39930
rect 10768 39802 11088 40041
rect 11222 40474 11318 40490
rect 11222 40410 11238 40474
rect 11302 40410 11318 40474
rect 11222 40394 11318 40410
rect 11222 40330 11238 40394
rect 11302 40330 11318 40394
rect 11488 40363 11808 40741
rect 11941 41030 11957 41094
rect 12021 41030 12037 41094
rect 12660 41174 12756 41190
rect 12660 41110 12676 41174
rect 12740 41110 12756 41174
rect 12660 41094 12756 41110
rect 12208 41063 12528 41082
rect 11941 41014 12037 41030
rect 11941 40950 11957 41014
rect 12021 40950 12037 41014
rect 11941 40934 12037 40950
rect 11941 40870 11957 40934
rect 12021 40870 12037 40934
rect 11941 40854 12037 40870
rect 11941 40790 11957 40854
rect 12021 40790 12037 40854
rect 11941 40774 12037 40790
rect 11941 40710 11957 40774
rect 12021 40710 12037 40774
rect 12200 41054 12528 41063
rect 12200 40750 12209 41054
rect 12513 40750 12528 41054
rect 12200 40741 12528 40750
rect 11941 40694 12037 40710
rect 11941 40630 11957 40694
rect 12021 40630 12037 40694
rect 11941 40614 12037 40630
rect 11222 40314 11318 40330
rect 11222 40250 11238 40314
rect 11302 40250 11318 40314
rect 11222 40234 11318 40250
rect 11222 40170 11238 40234
rect 11302 40170 11318 40234
rect 11222 40154 11318 40170
rect 11222 40090 11238 40154
rect 11302 40090 11318 40154
rect 11222 40074 11318 40090
rect 11222 40010 11238 40074
rect 11302 40010 11318 40074
rect 11481 40354 11808 40363
rect 11481 40050 11490 40354
rect 11794 40050 11808 40354
rect 11481 40041 11808 40050
rect 11222 39994 11318 40010
rect 11222 39930 11238 39994
rect 11302 39930 11318 39994
rect 11222 39914 11318 39930
rect 11488 39802 11808 40041
rect 11941 40474 12037 40490
rect 11941 40410 11957 40474
rect 12021 40410 12037 40474
rect 11941 40394 12037 40410
rect 11941 40330 11957 40394
rect 12021 40330 12037 40394
rect 12208 40363 12528 40741
rect 12660 41030 12676 41094
rect 12740 41030 12756 41094
rect 13379 41174 13475 41190
rect 13379 41110 13395 41174
rect 13459 41110 13475 41174
rect 13379 41094 13475 41110
rect 12928 41063 13248 41082
rect 12660 41014 12756 41030
rect 12660 40950 12676 41014
rect 12740 40950 12756 41014
rect 12660 40934 12756 40950
rect 12660 40870 12676 40934
rect 12740 40870 12756 40934
rect 12660 40854 12756 40870
rect 12660 40790 12676 40854
rect 12740 40790 12756 40854
rect 12660 40774 12756 40790
rect 12660 40710 12676 40774
rect 12740 40710 12756 40774
rect 12919 41054 13248 41063
rect 12919 40750 12928 41054
rect 13232 40750 13248 41054
rect 12919 40741 13248 40750
rect 12660 40694 12756 40710
rect 12660 40630 12676 40694
rect 12740 40630 12756 40694
rect 12660 40614 12756 40630
rect 11941 40314 12037 40330
rect 11941 40250 11957 40314
rect 12021 40250 12037 40314
rect 11941 40234 12037 40250
rect 11941 40170 11957 40234
rect 12021 40170 12037 40234
rect 11941 40154 12037 40170
rect 11941 40090 11957 40154
rect 12021 40090 12037 40154
rect 11941 40074 12037 40090
rect 11941 40010 11957 40074
rect 12021 40010 12037 40074
rect 12200 40354 12528 40363
rect 12200 40050 12209 40354
rect 12513 40050 12528 40354
rect 12200 40041 12528 40050
rect 11941 39994 12037 40010
rect 11941 39930 11957 39994
rect 12021 39930 12037 39994
rect 11941 39914 12037 39930
rect 12208 39802 12528 40041
rect 12660 40474 12756 40490
rect 12660 40410 12676 40474
rect 12740 40410 12756 40474
rect 12660 40394 12756 40410
rect 12660 40330 12676 40394
rect 12740 40330 12756 40394
rect 12928 40363 13248 40741
rect 13379 41030 13395 41094
rect 13459 41030 13475 41094
rect 15728 41174 15824 41190
rect 15728 41110 15744 41174
rect 15808 41110 15824 41174
rect 15728 41094 15824 41110
rect 13379 41014 13475 41030
rect 13379 40950 13395 41014
rect 13459 40950 13475 41014
rect 13379 40934 13475 40950
rect 13379 40870 13395 40934
rect 13459 40870 13475 40934
rect 13379 40854 13475 40870
rect 13379 40790 13395 40854
rect 13459 40790 13475 40854
rect 13379 40774 13475 40790
rect 13379 40710 13395 40774
rect 13459 40710 13475 40774
rect 13379 40694 13475 40710
rect 13379 40630 13395 40694
rect 13459 40630 13475 40694
rect 13379 40614 13475 40630
rect 15268 41063 15588 41082
rect 15268 41054 15590 41063
rect 15268 40750 15277 41054
rect 15581 40750 15590 41054
rect 15268 40741 15590 40750
rect 15728 41030 15744 41094
rect 15808 41030 15824 41094
rect 16447 41174 16543 41190
rect 16447 41110 16463 41174
rect 16527 41110 16543 41174
rect 16447 41094 16543 41110
rect 15988 41063 16308 41082
rect 15728 41014 15824 41030
rect 15728 40950 15744 41014
rect 15808 40950 15824 41014
rect 15728 40934 15824 40950
rect 15728 40870 15744 40934
rect 15808 40870 15824 40934
rect 15728 40854 15824 40870
rect 15728 40790 15744 40854
rect 15808 40790 15824 40854
rect 15728 40774 15824 40790
rect 12660 40314 12756 40330
rect 12660 40250 12676 40314
rect 12740 40250 12756 40314
rect 12660 40234 12756 40250
rect 12660 40170 12676 40234
rect 12740 40170 12756 40234
rect 12660 40154 12756 40170
rect 12660 40090 12676 40154
rect 12740 40090 12756 40154
rect 12660 40074 12756 40090
rect 12660 40010 12676 40074
rect 12740 40010 12756 40074
rect 12919 40354 13248 40363
rect 12919 40050 12928 40354
rect 13232 40050 13248 40354
rect 12919 40041 13248 40050
rect 12660 39994 12756 40010
rect 12660 39930 12676 39994
rect 12740 39930 12756 39994
rect 12660 39914 12756 39930
rect 12928 39802 13248 40041
rect 13379 40474 13475 40490
rect 13379 40410 13395 40474
rect 13459 40410 13475 40474
rect 13379 40394 13475 40410
rect 13379 40330 13395 40394
rect 13459 40330 13475 40394
rect 13379 40314 13475 40330
rect 13379 40250 13395 40314
rect 13459 40250 13475 40314
rect 13379 40234 13475 40250
rect 13379 40170 13395 40234
rect 13459 40170 13475 40234
rect 13379 40154 13475 40170
rect 13379 40090 13395 40154
rect 13459 40090 13475 40154
rect 13379 40074 13475 40090
rect 13379 40010 13395 40074
rect 13459 40010 13475 40074
rect 13379 39994 13475 40010
rect 13379 39930 13395 39994
rect 13459 39936 13475 39994
rect 15268 40363 15588 40741
rect 15728 40710 15744 40774
rect 15808 40710 15824 40774
rect 15987 41054 16309 41063
rect 15987 40750 15996 41054
rect 16300 40750 16309 41054
rect 15987 40741 16309 40750
rect 16447 41030 16463 41094
rect 16527 41030 16543 41094
rect 17166 41174 17262 41190
rect 17166 41110 17182 41174
rect 17246 41110 17262 41174
rect 17166 41094 17262 41110
rect 16708 41063 17028 41082
rect 16447 41014 16543 41030
rect 16447 40950 16463 41014
rect 16527 40950 16543 41014
rect 16447 40934 16543 40950
rect 16447 40870 16463 40934
rect 16527 40870 16543 40934
rect 16447 40854 16543 40870
rect 16447 40790 16463 40854
rect 16527 40790 16543 40854
rect 16447 40774 16543 40790
rect 15728 40694 15824 40710
rect 15728 40630 15744 40694
rect 15808 40630 15824 40694
rect 15728 40614 15824 40630
rect 15728 40474 15824 40490
rect 15728 40410 15744 40474
rect 15808 40410 15824 40474
rect 15728 40394 15824 40410
rect 15268 40354 15590 40363
rect 15268 40050 15277 40354
rect 15581 40050 15590 40354
rect 15268 40041 15590 40050
rect 15728 40330 15744 40394
rect 15808 40330 15824 40394
rect 15988 40363 16308 40741
rect 16447 40710 16463 40774
rect 16527 40710 16543 40774
rect 16706 41054 17028 41063
rect 16706 40750 16715 41054
rect 17019 40750 17028 41054
rect 16706 40741 17028 40750
rect 16447 40694 16543 40710
rect 16447 40630 16463 40694
rect 16527 40630 16543 40694
rect 16447 40614 16543 40630
rect 16447 40474 16543 40490
rect 16447 40410 16463 40474
rect 16527 40410 16543 40474
rect 16447 40394 16543 40410
rect 15728 40314 15824 40330
rect 15728 40250 15744 40314
rect 15808 40250 15824 40314
rect 15728 40234 15824 40250
rect 15728 40170 15744 40234
rect 15808 40170 15824 40234
rect 15728 40154 15824 40170
rect 15728 40090 15744 40154
rect 15808 40090 15824 40154
rect 15728 40074 15824 40090
rect 13459 39930 13600 39936
rect 13379 39914 13600 39930
rect 13402 39876 13600 39914
rect 6310 39774 13478 39802
rect 6310 39710 6338 39774
rect 6402 39710 6418 39774
rect 6482 39710 13478 39774
rect 6310 39682 13478 39710
rect 3348 37640 3372 37704
rect 3436 37640 3452 37704
rect 3516 37640 3532 37704
rect 3596 37640 3612 37704
rect 3676 37640 3692 37704
rect 3756 37640 3772 37704
rect 3836 37640 3852 37704
rect 3916 37640 3932 37704
rect 3996 37640 4012 37704
rect 4076 37640 4092 37704
rect 4156 37640 4172 37704
rect 4236 37640 4252 37704
rect 4316 37640 4332 37704
rect 4396 37640 4412 37704
rect 4476 37640 4492 37704
rect 4556 37640 4572 37704
rect 4636 37640 4652 37704
rect 4716 37640 4732 37704
rect 4796 37640 4812 37704
rect 4876 37640 4892 37704
rect 4956 37640 4980 37704
rect 3348 33944 4980 37640
rect 13540 37255 13600 39876
rect 15268 39802 15588 40041
rect 15728 40010 15744 40074
rect 15808 40010 15824 40074
rect 15987 40354 16309 40363
rect 15987 40050 15996 40354
rect 16300 40050 16309 40354
rect 15987 40041 16309 40050
rect 16447 40330 16463 40394
rect 16527 40330 16543 40394
rect 16708 40363 17028 40741
rect 17166 41030 17182 41094
rect 17246 41030 17262 41094
rect 17885 41174 17981 41190
rect 17885 41110 17901 41174
rect 17965 41110 17981 41174
rect 17885 41094 17981 41110
rect 17428 41063 17748 41082
rect 17166 41014 17262 41030
rect 17166 40950 17182 41014
rect 17246 40950 17262 41014
rect 17166 40934 17262 40950
rect 17166 40870 17182 40934
rect 17246 40870 17262 40934
rect 17166 40854 17262 40870
rect 17166 40790 17182 40854
rect 17246 40790 17262 40854
rect 17166 40774 17262 40790
rect 17166 40710 17182 40774
rect 17246 40710 17262 40774
rect 17425 41054 17748 41063
rect 17425 40750 17434 41054
rect 17738 40750 17748 41054
rect 17425 40741 17748 40750
rect 17166 40694 17262 40710
rect 17166 40630 17182 40694
rect 17246 40630 17262 40694
rect 17166 40614 17262 40630
rect 16447 40314 16543 40330
rect 16447 40250 16463 40314
rect 16527 40250 16543 40314
rect 16447 40234 16543 40250
rect 16447 40170 16463 40234
rect 16527 40170 16543 40234
rect 16447 40154 16543 40170
rect 16447 40090 16463 40154
rect 16527 40090 16543 40154
rect 16447 40074 16543 40090
rect 15728 39994 15824 40010
rect 15728 39930 15744 39994
rect 15808 39930 15824 39994
rect 15728 39914 15824 39930
rect 15988 39802 16308 40041
rect 16447 40010 16463 40074
rect 16527 40010 16543 40074
rect 16706 40354 17028 40363
rect 16706 40050 16715 40354
rect 17019 40050 17028 40354
rect 16706 40041 17028 40050
rect 16447 39994 16543 40010
rect 16447 39930 16463 39994
rect 16527 39930 16543 39994
rect 16447 39914 16543 39930
rect 16708 39802 17028 40041
rect 17166 40474 17262 40490
rect 17166 40410 17182 40474
rect 17246 40410 17262 40474
rect 17166 40394 17262 40410
rect 17166 40330 17182 40394
rect 17246 40330 17262 40394
rect 17428 40363 17748 40741
rect 17885 41030 17901 41094
rect 17965 41030 17981 41094
rect 18604 41174 18700 41190
rect 18604 41110 18620 41174
rect 18684 41110 18700 41174
rect 18604 41094 18700 41110
rect 18148 41063 18468 41082
rect 17885 41014 17981 41030
rect 17885 40950 17901 41014
rect 17965 40950 17981 41014
rect 17885 40934 17981 40950
rect 17885 40870 17901 40934
rect 17965 40870 17981 40934
rect 17885 40854 17981 40870
rect 17885 40790 17901 40854
rect 17965 40790 17981 40854
rect 17885 40774 17981 40790
rect 17885 40710 17901 40774
rect 17965 40710 17981 40774
rect 18144 41054 18468 41063
rect 18144 40750 18153 41054
rect 18457 40750 18468 41054
rect 18144 40741 18468 40750
rect 17885 40694 17981 40710
rect 17885 40630 17901 40694
rect 17965 40630 17981 40694
rect 17885 40614 17981 40630
rect 17166 40314 17262 40330
rect 17166 40250 17182 40314
rect 17246 40250 17262 40314
rect 17166 40234 17262 40250
rect 17166 40170 17182 40234
rect 17246 40170 17262 40234
rect 17166 40154 17262 40170
rect 17166 40090 17182 40154
rect 17246 40090 17262 40154
rect 17166 40074 17262 40090
rect 17166 40010 17182 40074
rect 17246 40010 17262 40074
rect 17425 40354 17748 40363
rect 17425 40050 17434 40354
rect 17738 40050 17748 40354
rect 17425 40041 17748 40050
rect 17166 39994 17262 40010
rect 17166 39930 17182 39994
rect 17246 39930 17262 39994
rect 17166 39914 17262 39930
rect 17428 39802 17748 40041
rect 17885 40474 17981 40490
rect 17885 40410 17901 40474
rect 17965 40410 17981 40474
rect 17885 40394 17981 40410
rect 17885 40330 17901 40394
rect 17965 40330 17981 40394
rect 18148 40363 18468 40741
rect 18604 41030 18620 41094
rect 18684 41030 18700 41094
rect 19323 41174 19419 41190
rect 19323 41110 19339 41174
rect 19403 41110 19419 41174
rect 19323 41094 19419 41110
rect 18868 41063 19188 41082
rect 18604 41014 18700 41030
rect 18604 40950 18620 41014
rect 18684 40950 18700 41014
rect 18604 40934 18700 40950
rect 18604 40870 18620 40934
rect 18684 40870 18700 40934
rect 18604 40854 18700 40870
rect 18604 40790 18620 40854
rect 18684 40790 18700 40854
rect 18604 40774 18700 40790
rect 18604 40710 18620 40774
rect 18684 40710 18700 40774
rect 18863 41054 19188 41063
rect 18863 40750 18872 41054
rect 19176 40750 19188 41054
rect 18863 40741 19188 40750
rect 18604 40694 18700 40710
rect 18604 40630 18620 40694
rect 18684 40630 18700 40694
rect 18604 40614 18700 40630
rect 17885 40314 17981 40330
rect 17885 40250 17901 40314
rect 17965 40250 17981 40314
rect 17885 40234 17981 40250
rect 17885 40170 17901 40234
rect 17965 40170 17981 40234
rect 17885 40154 17981 40170
rect 17885 40090 17901 40154
rect 17965 40090 17981 40154
rect 17885 40074 17981 40090
rect 17885 40010 17901 40074
rect 17965 40010 17981 40074
rect 18144 40354 18468 40363
rect 18144 40050 18153 40354
rect 18457 40050 18468 40354
rect 18144 40041 18468 40050
rect 17885 39994 17981 40010
rect 17885 39930 17901 39994
rect 17965 39930 17981 39994
rect 17885 39914 17981 39930
rect 18148 39802 18468 40041
rect 18604 40474 18700 40490
rect 18604 40410 18620 40474
rect 18684 40410 18700 40474
rect 18604 40394 18700 40410
rect 18604 40330 18620 40394
rect 18684 40330 18700 40394
rect 18868 40363 19188 40741
rect 19323 41030 19339 41094
rect 19403 41030 19419 41094
rect 20042 41174 20138 41190
rect 20042 41110 20058 41174
rect 20122 41110 20138 41174
rect 20042 41094 20138 41110
rect 19588 41063 19908 41082
rect 19323 41014 19419 41030
rect 19323 40950 19339 41014
rect 19403 40950 19419 41014
rect 19323 40934 19419 40950
rect 19323 40870 19339 40934
rect 19403 40870 19419 40934
rect 19323 40854 19419 40870
rect 19323 40790 19339 40854
rect 19403 40790 19419 40854
rect 19323 40774 19419 40790
rect 19323 40710 19339 40774
rect 19403 40710 19419 40774
rect 19582 41054 19908 41063
rect 19582 40750 19591 41054
rect 19895 40750 19908 41054
rect 19582 40741 19908 40750
rect 19323 40694 19419 40710
rect 19323 40630 19339 40694
rect 19403 40630 19419 40694
rect 19323 40614 19419 40630
rect 18604 40314 18700 40330
rect 18604 40250 18620 40314
rect 18684 40250 18700 40314
rect 18604 40234 18700 40250
rect 18604 40170 18620 40234
rect 18684 40170 18700 40234
rect 18604 40154 18700 40170
rect 18604 40090 18620 40154
rect 18684 40090 18700 40154
rect 18604 40074 18700 40090
rect 18604 40010 18620 40074
rect 18684 40010 18700 40074
rect 18863 40354 19188 40363
rect 18863 40050 18872 40354
rect 19176 40050 19188 40354
rect 18863 40041 19188 40050
rect 18604 39994 18700 40010
rect 18604 39930 18620 39994
rect 18684 39930 18700 39994
rect 18604 39914 18700 39930
rect 18868 39802 19188 40041
rect 19323 40474 19419 40490
rect 19323 40410 19339 40474
rect 19403 40410 19419 40474
rect 19323 40394 19419 40410
rect 19323 40330 19339 40394
rect 19403 40330 19419 40394
rect 19588 40363 19908 40741
rect 20042 41030 20058 41094
rect 20122 41030 20138 41094
rect 20761 41174 20857 41190
rect 20761 41110 20777 41174
rect 20841 41110 20857 41174
rect 20761 41094 20857 41110
rect 20308 41063 20628 41082
rect 20042 41014 20138 41030
rect 20042 40950 20058 41014
rect 20122 40950 20138 41014
rect 20042 40934 20138 40950
rect 20042 40870 20058 40934
rect 20122 40870 20138 40934
rect 20042 40854 20138 40870
rect 20042 40790 20058 40854
rect 20122 40790 20138 40854
rect 20042 40774 20138 40790
rect 20042 40710 20058 40774
rect 20122 40710 20138 40774
rect 20301 41054 20628 41063
rect 20301 40750 20310 41054
rect 20614 40750 20628 41054
rect 20301 40741 20628 40750
rect 20042 40694 20138 40710
rect 20042 40630 20058 40694
rect 20122 40630 20138 40694
rect 20042 40614 20138 40630
rect 19323 40314 19419 40330
rect 19323 40250 19339 40314
rect 19403 40250 19419 40314
rect 19323 40234 19419 40250
rect 19323 40170 19339 40234
rect 19403 40170 19419 40234
rect 19323 40154 19419 40170
rect 19323 40090 19339 40154
rect 19403 40090 19419 40154
rect 19323 40074 19419 40090
rect 19323 40010 19339 40074
rect 19403 40010 19419 40074
rect 19582 40354 19908 40363
rect 19582 40050 19591 40354
rect 19895 40050 19908 40354
rect 19582 40041 19908 40050
rect 19323 39994 19419 40010
rect 19323 39930 19339 39994
rect 19403 39930 19419 39994
rect 19323 39914 19419 39930
rect 19588 39802 19908 40041
rect 20042 40474 20138 40490
rect 20042 40410 20058 40474
rect 20122 40410 20138 40474
rect 20042 40394 20138 40410
rect 20042 40330 20058 40394
rect 20122 40330 20138 40394
rect 20308 40363 20628 40741
rect 20761 41030 20777 41094
rect 20841 41030 20857 41094
rect 21480 41174 21576 41190
rect 21480 41110 21496 41174
rect 21560 41110 21576 41174
rect 21480 41094 21576 41110
rect 21028 41063 21348 41082
rect 20761 41014 20857 41030
rect 20761 40950 20777 41014
rect 20841 40950 20857 41014
rect 20761 40934 20857 40950
rect 20761 40870 20777 40934
rect 20841 40870 20857 40934
rect 20761 40854 20857 40870
rect 20761 40790 20777 40854
rect 20841 40790 20857 40854
rect 20761 40774 20857 40790
rect 20761 40710 20777 40774
rect 20841 40710 20857 40774
rect 21020 41054 21348 41063
rect 21020 40750 21029 41054
rect 21333 40750 21348 41054
rect 21020 40741 21348 40750
rect 20761 40694 20857 40710
rect 20761 40630 20777 40694
rect 20841 40630 20857 40694
rect 20761 40614 20857 40630
rect 20042 40314 20138 40330
rect 20042 40250 20058 40314
rect 20122 40250 20138 40314
rect 20042 40234 20138 40250
rect 20042 40170 20058 40234
rect 20122 40170 20138 40234
rect 20042 40154 20138 40170
rect 20042 40090 20058 40154
rect 20122 40090 20138 40154
rect 20042 40074 20138 40090
rect 20042 40010 20058 40074
rect 20122 40010 20138 40074
rect 20301 40354 20628 40363
rect 20301 40050 20310 40354
rect 20614 40050 20628 40354
rect 20301 40041 20628 40050
rect 20042 39994 20138 40010
rect 20042 39930 20058 39994
rect 20122 39930 20138 39994
rect 20042 39914 20138 39930
rect 20308 39802 20628 40041
rect 20761 40474 20857 40490
rect 20761 40410 20777 40474
rect 20841 40410 20857 40474
rect 20761 40394 20857 40410
rect 20761 40330 20777 40394
rect 20841 40330 20857 40394
rect 21028 40363 21348 40741
rect 21480 41030 21496 41094
rect 21560 41030 21576 41094
rect 22199 41174 22295 41190
rect 22199 41110 22215 41174
rect 22279 41110 22295 41174
rect 22199 41094 22295 41110
rect 21748 41063 22068 41082
rect 21480 41014 21576 41030
rect 21480 40950 21496 41014
rect 21560 40950 21576 41014
rect 21480 40934 21576 40950
rect 21480 40870 21496 40934
rect 21560 40870 21576 40934
rect 21480 40854 21576 40870
rect 21480 40790 21496 40854
rect 21560 40790 21576 40854
rect 21480 40774 21576 40790
rect 21480 40710 21496 40774
rect 21560 40710 21576 40774
rect 21739 41054 22068 41063
rect 21739 40750 21748 41054
rect 22052 40750 22068 41054
rect 21739 40741 22068 40750
rect 21480 40694 21576 40710
rect 21480 40630 21496 40694
rect 21560 40630 21576 40694
rect 21480 40614 21576 40630
rect 20761 40314 20857 40330
rect 20761 40250 20777 40314
rect 20841 40250 20857 40314
rect 20761 40234 20857 40250
rect 20761 40170 20777 40234
rect 20841 40170 20857 40234
rect 20761 40154 20857 40170
rect 20761 40090 20777 40154
rect 20841 40090 20857 40154
rect 20761 40074 20857 40090
rect 20761 40010 20777 40074
rect 20841 40010 20857 40074
rect 21020 40354 21348 40363
rect 21020 40050 21029 40354
rect 21333 40050 21348 40354
rect 21020 40041 21348 40050
rect 20761 39994 20857 40010
rect 20761 39930 20777 39994
rect 20841 39930 20857 39994
rect 20761 39914 20857 39930
rect 21028 39802 21348 40041
rect 21480 40474 21576 40490
rect 21480 40410 21496 40474
rect 21560 40410 21576 40474
rect 21480 40394 21576 40410
rect 21480 40330 21496 40394
rect 21560 40330 21576 40394
rect 21748 40363 22068 40741
rect 22199 41030 22215 41094
rect 22279 41030 22295 41094
rect 22199 41014 22295 41030
rect 22199 40950 22215 41014
rect 22279 40950 22295 41014
rect 22199 40934 22295 40950
rect 22199 40870 22215 40934
rect 22279 40870 22295 40934
rect 22199 40854 22295 40870
rect 22199 40790 22215 40854
rect 22279 40790 22295 40854
rect 22199 40774 22295 40790
rect 22199 40710 22215 40774
rect 22279 40710 22295 40774
rect 22199 40694 22295 40710
rect 22199 40630 22215 40694
rect 22279 40630 22295 40694
rect 22199 40614 22295 40630
rect 21480 40314 21576 40330
rect 21480 40250 21496 40314
rect 21560 40250 21576 40314
rect 21480 40234 21576 40250
rect 21480 40170 21496 40234
rect 21560 40170 21576 40234
rect 21480 40154 21576 40170
rect 21480 40090 21496 40154
rect 21560 40090 21576 40154
rect 21480 40074 21576 40090
rect 21480 40010 21496 40074
rect 21560 40010 21576 40074
rect 21739 40354 22068 40363
rect 21739 40050 21748 40354
rect 22052 40050 22068 40354
rect 21739 40041 22068 40050
rect 21480 39994 21576 40010
rect 21480 39930 21496 39994
rect 21560 39930 21576 39994
rect 21480 39914 21576 39930
rect 21748 39802 22068 40041
rect 22199 40474 22295 40490
rect 22199 40410 22215 40474
rect 22279 40410 22295 40474
rect 22199 40394 22295 40410
rect 22199 40330 22215 40394
rect 22279 40330 22295 40394
rect 22199 40314 22295 40330
rect 22199 40250 22215 40314
rect 22279 40250 22295 40314
rect 22199 40234 22295 40250
rect 22199 40170 22215 40234
rect 22279 40170 22295 40234
rect 22199 40154 22295 40170
rect 22199 40090 22215 40154
rect 22279 40090 22295 40154
rect 22199 40074 22295 40090
rect 22199 40010 22215 40074
rect 22279 40010 22295 40074
rect 22199 39994 22295 40010
rect 22199 39930 22215 39994
rect 22279 39930 22295 39994
rect 22199 39914 22295 39930
rect 15130 39774 22298 39802
rect 15130 39710 15158 39774
rect 15222 39710 15238 39774
rect 15302 39710 22298 39774
rect 15130 39694 22298 39710
rect 15130 39682 15470 39694
rect 15469 39630 15470 39682
rect 15534 39682 22298 39694
rect 15534 39630 15535 39682
rect 15469 39629 15535 39630
rect 53456 37704 55088 41400
rect 53456 37640 53480 37704
rect 53544 37640 53560 37704
rect 53624 37640 53640 37704
rect 53704 37640 53720 37704
rect 53784 37640 53800 37704
rect 53864 37640 53880 37704
rect 53944 37640 53960 37704
rect 54024 37640 54040 37704
rect 54104 37640 54120 37704
rect 54184 37640 54200 37704
rect 54264 37640 54280 37704
rect 54344 37640 54360 37704
rect 54424 37640 54440 37704
rect 54504 37640 54520 37704
rect 54584 37640 54600 37704
rect 54664 37640 54680 37704
rect 54744 37640 54760 37704
rect 54824 37640 54840 37704
rect 54904 37640 54920 37704
rect 54984 37640 55000 37704
rect 55064 37640 55088 37704
rect 33409 37620 33475 37621
rect 33409 37556 33410 37620
rect 33474 37556 33475 37620
rect 33409 37555 33475 37556
rect 33412 37430 33472 37555
rect 30526 37414 30622 37430
rect 30526 37350 30542 37414
rect 30606 37350 30622 37414
rect 30526 37334 30622 37350
rect 30066 37303 30386 37322
rect 30066 37294 30388 37303
rect 13537 37254 13603 37255
rect 13537 37190 13538 37254
rect 13602 37190 13603 37254
rect 13537 37189 13603 37190
rect 29683 37010 29749 37011
rect 29683 36946 29684 37010
rect 29748 37008 29749 37010
rect 30066 37008 30075 37294
rect 29748 36990 30075 37008
rect 30379 36990 30388 37294
rect 29748 36981 30388 36990
rect 30526 37270 30542 37334
rect 30606 37270 30622 37334
rect 31245 37414 31341 37430
rect 31245 37350 31261 37414
rect 31325 37350 31341 37414
rect 31245 37334 31341 37350
rect 30786 37303 31106 37322
rect 30526 37254 30622 37270
rect 30526 37190 30542 37254
rect 30606 37190 30622 37254
rect 30526 37174 30622 37190
rect 30526 37110 30542 37174
rect 30606 37110 30622 37174
rect 30526 37094 30622 37110
rect 30526 37030 30542 37094
rect 30606 37030 30622 37094
rect 30526 37014 30622 37030
rect 29748 36948 30386 36981
rect 29748 36946 29749 36948
rect 29683 36945 29749 36946
rect 30066 36603 30386 36948
rect 30526 36950 30542 37014
rect 30606 36950 30622 37014
rect 30785 37294 31107 37303
rect 30785 36990 30794 37294
rect 31098 36990 31107 37294
rect 30785 36981 31107 36990
rect 31245 37270 31261 37334
rect 31325 37270 31341 37334
rect 31964 37414 32060 37430
rect 31964 37350 31980 37414
rect 32044 37350 32060 37414
rect 31964 37334 32060 37350
rect 31506 37303 31826 37322
rect 31245 37254 31341 37270
rect 31245 37190 31261 37254
rect 31325 37190 31341 37254
rect 31245 37174 31341 37190
rect 31245 37110 31261 37174
rect 31325 37110 31341 37174
rect 31245 37094 31341 37110
rect 31245 37030 31261 37094
rect 31325 37030 31341 37094
rect 31245 37014 31341 37030
rect 30526 36934 30622 36950
rect 30526 36870 30542 36934
rect 30606 36870 30622 36934
rect 30526 36854 30622 36870
rect 30526 36714 30622 36730
rect 30526 36650 30542 36714
rect 30606 36650 30622 36714
rect 30526 36634 30622 36650
rect 30066 36594 30388 36603
rect 30066 36290 30075 36594
rect 30379 36290 30388 36594
rect 30066 36281 30388 36290
rect 30526 36570 30542 36634
rect 30606 36570 30622 36634
rect 30786 36603 31106 36981
rect 31245 36950 31261 37014
rect 31325 36950 31341 37014
rect 31504 37294 31826 37303
rect 31504 36990 31513 37294
rect 31817 36990 31826 37294
rect 31504 36981 31826 36990
rect 31245 36934 31341 36950
rect 31245 36870 31261 36934
rect 31325 36870 31341 36934
rect 31245 36854 31341 36870
rect 31245 36714 31341 36730
rect 31245 36650 31261 36714
rect 31325 36650 31341 36714
rect 31245 36634 31341 36650
rect 30526 36554 30622 36570
rect 30526 36490 30542 36554
rect 30606 36490 30622 36554
rect 30526 36474 30622 36490
rect 30526 36410 30542 36474
rect 30606 36410 30622 36474
rect 30526 36394 30622 36410
rect 30526 36330 30542 36394
rect 30606 36330 30622 36394
rect 30526 36314 30622 36330
rect 30066 36042 30386 36281
rect 30526 36250 30542 36314
rect 30606 36250 30622 36314
rect 30785 36594 31107 36603
rect 30785 36290 30794 36594
rect 31098 36290 31107 36594
rect 30785 36281 31107 36290
rect 31245 36570 31261 36634
rect 31325 36570 31341 36634
rect 31506 36603 31826 36981
rect 31964 37270 31980 37334
rect 32044 37270 32060 37334
rect 32683 37414 32779 37430
rect 32683 37350 32699 37414
rect 32763 37350 32779 37414
rect 32683 37334 32779 37350
rect 32226 37303 32546 37322
rect 31964 37254 32060 37270
rect 31964 37190 31980 37254
rect 32044 37190 32060 37254
rect 31964 37174 32060 37190
rect 31964 37110 31980 37174
rect 32044 37110 32060 37174
rect 31964 37094 32060 37110
rect 31964 37030 31980 37094
rect 32044 37030 32060 37094
rect 31964 37014 32060 37030
rect 31964 36950 31980 37014
rect 32044 36950 32060 37014
rect 32223 37294 32546 37303
rect 32223 36990 32232 37294
rect 32536 36990 32546 37294
rect 32223 36981 32546 36990
rect 31964 36934 32060 36950
rect 31964 36870 31980 36934
rect 32044 36870 32060 36934
rect 31964 36854 32060 36870
rect 31245 36554 31341 36570
rect 31245 36490 31261 36554
rect 31325 36490 31341 36554
rect 31245 36474 31341 36490
rect 31245 36410 31261 36474
rect 31325 36410 31341 36474
rect 31245 36394 31341 36410
rect 31245 36330 31261 36394
rect 31325 36330 31341 36394
rect 31245 36314 31341 36330
rect 30526 36234 30622 36250
rect 30526 36170 30542 36234
rect 30606 36170 30622 36234
rect 30526 36154 30622 36170
rect 30786 36042 31106 36281
rect 31245 36250 31261 36314
rect 31325 36250 31341 36314
rect 31504 36594 31826 36603
rect 31504 36290 31513 36594
rect 31817 36290 31826 36594
rect 31504 36281 31826 36290
rect 31245 36234 31341 36250
rect 31245 36170 31261 36234
rect 31325 36170 31341 36234
rect 31245 36154 31341 36170
rect 31506 36042 31826 36281
rect 31964 36714 32060 36730
rect 31964 36650 31980 36714
rect 32044 36650 32060 36714
rect 31964 36634 32060 36650
rect 31964 36570 31980 36634
rect 32044 36570 32060 36634
rect 32226 36603 32546 36981
rect 32683 37270 32699 37334
rect 32763 37270 32779 37334
rect 33402 37414 33498 37430
rect 33402 37350 33418 37414
rect 33482 37350 33498 37414
rect 33402 37334 33498 37350
rect 32946 37303 33266 37322
rect 32683 37254 32779 37270
rect 32683 37190 32699 37254
rect 32763 37190 32779 37254
rect 32683 37174 32779 37190
rect 32683 37110 32699 37174
rect 32763 37110 32779 37174
rect 32683 37094 32779 37110
rect 32683 37030 32699 37094
rect 32763 37030 32779 37094
rect 32683 37014 32779 37030
rect 32683 36950 32699 37014
rect 32763 36950 32779 37014
rect 32942 37294 33266 37303
rect 32942 36990 32951 37294
rect 33255 36990 33266 37294
rect 32942 36981 33266 36990
rect 32683 36934 32779 36950
rect 32683 36870 32699 36934
rect 32763 36870 32779 36934
rect 32683 36854 32779 36870
rect 31964 36554 32060 36570
rect 31964 36490 31980 36554
rect 32044 36490 32060 36554
rect 31964 36474 32060 36490
rect 31964 36410 31980 36474
rect 32044 36410 32060 36474
rect 31964 36394 32060 36410
rect 31964 36330 31980 36394
rect 32044 36330 32060 36394
rect 31964 36314 32060 36330
rect 31964 36250 31980 36314
rect 32044 36250 32060 36314
rect 32223 36594 32546 36603
rect 32223 36290 32232 36594
rect 32536 36290 32546 36594
rect 32223 36281 32546 36290
rect 31964 36234 32060 36250
rect 31964 36170 31980 36234
rect 32044 36170 32060 36234
rect 31964 36154 32060 36170
rect 32226 36042 32546 36281
rect 32683 36714 32779 36730
rect 32683 36650 32699 36714
rect 32763 36650 32779 36714
rect 32683 36634 32779 36650
rect 32683 36570 32699 36634
rect 32763 36570 32779 36634
rect 32946 36603 33266 36981
rect 33402 37270 33418 37334
rect 33482 37270 33498 37334
rect 34121 37414 34217 37430
rect 34121 37350 34137 37414
rect 34201 37350 34217 37414
rect 34121 37334 34217 37350
rect 33666 37303 33986 37322
rect 33402 37254 33498 37270
rect 33402 37190 33418 37254
rect 33482 37190 33498 37254
rect 33402 37174 33498 37190
rect 33402 37110 33418 37174
rect 33482 37110 33498 37174
rect 33402 37094 33498 37110
rect 33402 37030 33418 37094
rect 33482 37030 33498 37094
rect 33402 37014 33498 37030
rect 33402 36950 33418 37014
rect 33482 36950 33498 37014
rect 33661 37294 33986 37303
rect 33661 36990 33670 37294
rect 33974 36990 33986 37294
rect 33661 36981 33986 36990
rect 33402 36934 33498 36950
rect 33402 36870 33418 36934
rect 33482 36870 33498 36934
rect 33402 36854 33498 36870
rect 32683 36554 32779 36570
rect 32683 36490 32699 36554
rect 32763 36490 32779 36554
rect 32683 36474 32779 36490
rect 32683 36410 32699 36474
rect 32763 36410 32779 36474
rect 32683 36394 32779 36410
rect 32683 36330 32699 36394
rect 32763 36330 32779 36394
rect 32683 36314 32779 36330
rect 32683 36250 32699 36314
rect 32763 36250 32779 36314
rect 32942 36594 33266 36603
rect 32942 36290 32951 36594
rect 33255 36290 33266 36594
rect 32942 36281 33266 36290
rect 32683 36234 32779 36250
rect 32683 36170 32699 36234
rect 32763 36170 32779 36234
rect 32683 36154 32779 36170
rect 32946 36042 33266 36281
rect 33402 36714 33498 36730
rect 33402 36650 33418 36714
rect 33482 36650 33498 36714
rect 33402 36634 33498 36650
rect 33402 36570 33418 36634
rect 33482 36570 33498 36634
rect 33666 36603 33986 36981
rect 34121 37270 34137 37334
rect 34201 37270 34217 37334
rect 34840 37414 34936 37430
rect 34840 37350 34856 37414
rect 34920 37350 34936 37414
rect 34840 37334 34936 37350
rect 34386 37303 34706 37322
rect 34121 37254 34217 37270
rect 34121 37190 34137 37254
rect 34201 37190 34217 37254
rect 34121 37174 34217 37190
rect 34121 37110 34137 37174
rect 34201 37110 34217 37174
rect 34121 37094 34217 37110
rect 34121 37030 34137 37094
rect 34201 37030 34217 37094
rect 34121 37014 34217 37030
rect 34121 36950 34137 37014
rect 34201 36950 34217 37014
rect 34380 37294 34706 37303
rect 34380 36990 34389 37294
rect 34693 36990 34706 37294
rect 34380 36981 34706 36990
rect 34121 36934 34217 36950
rect 34121 36870 34137 36934
rect 34201 36870 34217 36934
rect 34121 36854 34217 36870
rect 33402 36554 33498 36570
rect 33402 36490 33418 36554
rect 33482 36490 33498 36554
rect 33402 36474 33498 36490
rect 33402 36410 33418 36474
rect 33482 36410 33498 36474
rect 33402 36394 33498 36410
rect 33402 36330 33418 36394
rect 33482 36330 33498 36394
rect 33402 36314 33498 36330
rect 33402 36250 33418 36314
rect 33482 36250 33498 36314
rect 33661 36594 33986 36603
rect 33661 36290 33670 36594
rect 33974 36290 33986 36594
rect 33661 36281 33986 36290
rect 33402 36234 33498 36250
rect 33402 36170 33418 36234
rect 33482 36170 33498 36234
rect 33402 36154 33498 36170
rect 33666 36042 33986 36281
rect 34121 36714 34217 36730
rect 34121 36650 34137 36714
rect 34201 36650 34217 36714
rect 34121 36634 34217 36650
rect 34121 36570 34137 36634
rect 34201 36570 34217 36634
rect 34386 36603 34706 36981
rect 34840 37270 34856 37334
rect 34920 37270 34936 37334
rect 35559 37414 35655 37430
rect 35559 37350 35575 37414
rect 35639 37350 35655 37414
rect 35559 37334 35655 37350
rect 35106 37303 35426 37322
rect 34840 37254 34936 37270
rect 34840 37190 34856 37254
rect 34920 37190 34936 37254
rect 34840 37174 34936 37190
rect 34840 37110 34856 37174
rect 34920 37110 34936 37174
rect 34840 37094 34936 37110
rect 34840 37030 34856 37094
rect 34920 37030 34936 37094
rect 34840 37014 34936 37030
rect 34840 36950 34856 37014
rect 34920 36950 34936 37014
rect 35099 37294 35426 37303
rect 35099 36990 35108 37294
rect 35412 36990 35426 37294
rect 35099 36981 35426 36990
rect 34840 36934 34936 36950
rect 34840 36870 34856 36934
rect 34920 36870 34936 36934
rect 34840 36854 34936 36870
rect 34121 36554 34217 36570
rect 34121 36490 34137 36554
rect 34201 36490 34217 36554
rect 34121 36474 34217 36490
rect 34121 36410 34137 36474
rect 34201 36410 34217 36474
rect 34121 36394 34217 36410
rect 34121 36330 34137 36394
rect 34201 36330 34217 36394
rect 34121 36314 34217 36330
rect 34121 36250 34137 36314
rect 34201 36250 34217 36314
rect 34380 36594 34706 36603
rect 34380 36290 34389 36594
rect 34693 36290 34706 36594
rect 34380 36281 34706 36290
rect 34121 36234 34217 36250
rect 34121 36170 34137 36234
rect 34201 36170 34217 36234
rect 34121 36154 34217 36170
rect 34386 36042 34706 36281
rect 34840 36714 34936 36730
rect 34840 36650 34856 36714
rect 34920 36650 34936 36714
rect 34840 36634 34936 36650
rect 34840 36570 34856 36634
rect 34920 36570 34936 36634
rect 35106 36603 35426 36981
rect 35559 37270 35575 37334
rect 35639 37270 35655 37334
rect 36278 37414 36374 37430
rect 36278 37350 36294 37414
rect 36358 37350 36374 37414
rect 36278 37334 36374 37350
rect 35826 37303 36146 37322
rect 35559 37254 35655 37270
rect 35559 37190 35575 37254
rect 35639 37190 35655 37254
rect 35559 37174 35655 37190
rect 35559 37110 35575 37174
rect 35639 37110 35655 37174
rect 35559 37094 35655 37110
rect 35559 37030 35575 37094
rect 35639 37030 35655 37094
rect 35559 37014 35655 37030
rect 35559 36950 35575 37014
rect 35639 36950 35655 37014
rect 35818 37294 36146 37303
rect 35818 36990 35827 37294
rect 36131 36990 36146 37294
rect 35818 36981 36146 36990
rect 35559 36934 35655 36950
rect 35559 36870 35575 36934
rect 35639 36870 35655 36934
rect 35559 36854 35655 36870
rect 34840 36554 34936 36570
rect 34840 36490 34856 36554
rect 34920 36490 34936 36554
rect 34840 36474 34936 36490
rect 34840 36410 34856 36474
rect 34920 36410 34936 36474
rect 34840 36394 34936 36410
rect 34840 36330 34856 36394
rect 34920 36330 34936 36394
rect 34840 36314 34936 36330
rect 34840 36250 34856 36314
rect 34920 36250 34936 36314
rect 35099 36594 35426 36603
rect 35099 36290 35108 36594
rect 35412 36290 35426 36594
rect 35099 36281 35426 36290
rect 34840 36234 34936 36250
rect 34840 36170 34856 36234
rect 34920 36170 34936 36234
rect 34840 36154 34936 36170
rect 35106 36042 35426 36281
rect 35559 36714 35655 36730
rect 35559 36650 35575 36714
rect 35639 36650 35655 36714
rect 35559 36634 35655 36650
rect 35559 36570 35575 36634
rect 35639 36570 35655 36634
rect 35826 36603 36146 36981
rect 36278 37270 36294 37334
rect 36358 37270 36374 37334
rect 36997 37414 37093 37430
rect 36997 37350 37013 37414
rect 37077 37350 37093 37414
rect 36997 37334 37093 37350
rect 36546 37303 36866 37322
rect 36278 37254 36374 37270
rect 36278 37190 36294 37254
rect 36358 37190 36374 37254
rect 36278 37174 36374 37190
rect 36278 37110 36294 37174
rect 36358 37110 36374 37174
rect 36278 37094 36374 37110
rect 36278 37030 36294 37094
rect 36358 37030 36374 37094
rect 36278 37014 36374 37030
rect 36278 36950 36294 37014
rect 36358 36950 36374 37014
rect 36537 37294 36866 37303
rect 36537 36990 36546 37294
rect 36850 36990 36866 37294
rect 36537 36981 36866 36990
rect 36278 36934 36374 36950
rect 36278 36870 36294 36934
rect 36358 36870 36374 36934
rect 36278 36854 36374 36870
rect 35559 36554 35655 36570
rect 35559 36490 35575 36554
rect 35639 36490 35655 36554
rect 35559 36474 35655 36490
rect 35559 36410 35575 36474
rect 35639 36410 35655 36474
rect 35559 36394 35655 36410
rect 35559 36330 35575 36394
rect 35639 36330 35655 36394
rect 35559 36314 35655 36330
rect 35559 36250 35575 36314
rect 35639 36250 35655 36314
rect 35818 36594 36146 36603
rect 35818 36290 35827 36594
rect 36131 36290 36146 36594
rect 35818 36281 36146 36290
rect 35559 36234 35655 36250
rect 35559 36170 35575 36234
rect 35639 36170 35655 36234
rect 35559 36154 35655 36170
rect 35826 36042 36146 36281
rect 36278 36714 36374 36730
rect 36278 36650 36294 36714
rect 36358 36650 36374 36714
rect 36278 36634 36374 36650
rect 36278 36570 36294 36634
rect 36358 36570 36374 36634
rect 36546 36603 36866 36981
rect 36997 37270 37013 37334
rect 37077 37270 37093 37334
rect 36997 37254 37093 37270
rect 36997 37190 37013 37254
rect 37077 37190 37093 37254
rect 36997 37174 37093 37190
rect 36997 37110 37013 37174
rect 37077 37110 37093 37174
rect 36997 37094 37093 37110
rect 36997 37030 37013 37094
rect 37077 37030 37093 37094
rect 36997 37014 37093 37030
rect 36997 36950 37013 37014
rect 37077 36950 37093 37014
rect 36997 36934 37093 36950
rect 36997 36870 37013 36934
rect 37077 36870 37093 36934
rect 36997 36854 37093 36870
rect 36278 36554 36374 36570
rect 36278 36490 36294 36554
rect 36358 36490 36374 36554
rect 36278 36474 36374 36490
rect 36278 36410 36294 36474
rect 36358 36410 36374 36474
rect 36278 36394 36374 36410
rect 36278 36330 36294 36394
rect 36358 36330 36374 36394
rect 36278 36314 36374 36330
rect 36278 36250 36294 36314
rect 36358 36250 36374 36314
rect 36537 36594 36866 36603
rect 36537 36290 36546 36594
rect 36850 36290 36866 36594
rect 36537 36281 36866 36290
rect 36278 36234 36374 36250
rect 36278 36170 36294 36234
rect 36358 36170 36374 36234
rect 36278 36154 36374 36170
rect 36546 36042 36866 36281
rect 36997 36714 37093 36730
rect 36997 36650 37013 36714
rect 37077 36650 37093 36714
rect 36997 36634 37093 36650
rect 36997 36570 37013 36634
rect 37077 36570 37093 36634
rect 36997 36554 37093 36570
rect 36997 36490 37013 36554
rect 37077 36490 37093 36554
rect 36997 36474 37093 36490
rect 36997 36410 37013 36474
rect 37077 36410 37093 36474
rect 36997 36394 37093 36410
rect 36997 36330 37013 36394
rect 37077 36330 37093 36394
rect 36997 36314 37093 36330
rect 36997 36250 37013 36314
rect 37077 36250 37093 36314
rect 36997 36234 37093 36250
rect 36997 36170 37013 36234
rect 37077 36170 37093 36234
rect 36997 36154 37093 36170
rect 29928 36014 37096 36042
rect 29928 35950 29956 36014
rect 30020 35950 30036 36014
rect 30100 35950 37096 36014
rect 37549 36034 37615 36035
rect 37549 35970 37550 36034
rect 37614 35970 37615 36034
rect 37549 35969 37615 35970
rect 29928 35922 37096 35950
rect 3348 33880 3372 33944
rect 3436 33880 3452 33944
rect 3516 33880 3532 33944
rect 3596 33880 3612 33944
rect 3676 33880 3692 33944
rect 3756 33880 3772 33944
rect 3836 33880 3852 33944
rect 3916 33880 3932 33944
rect 3996 33880 4012 33944
rect 4076 33880 4092 33944
rect 4156 33880 4172 33944
rect 4236 33880 4252 33944
rect 4316 33880 4332 33944
rect 4396 33880 4412 33944
rect 4476 33880 4492 33944
rect 4556 33880 4572 33944
rect 4636 33880 4652 33944
rect 4716 33880 4732 33944
rect 4796 33880 4812 33944
rect 4876 33880 4892 33944
rect 4956 33880 4980 33944
rect 3348 30184 4980 33880
rect 26802 33654 26898 33670
rect 26802 33590 26818 33654
rect 26882 33590 26898 33654
rect 26802 33574 26898 33590
rect 26342 33543 26662 33562
rect 26342 33534 26664 33543
rect 26342 33230 26351 33534
rect 26655 33230 26664 33534
rect 26342 33221 26664 33230
rect 26802 33510 26818 33574
rect 26882 33510 26898 33574
rect 27521 33654 27617 33670
rect 27521 33590 27537 33654
rect 27601 33590 27617 33654
rect 27521 33574 27617 33590
rect 27062 33543 27382 33562
rect 26802 33494 26898 33510
rect 26802 33430 26818 33494
rect 26882 33430 26898 33494
rect 26802 33414 26898 33430
rect 26802 33350 26818 33414
rect 26882 33350 26898 33414
rect 26802 33334 26898 33350
rect 26802 33270 26818 33334
rect 26882 33270 26898 33334
rect 26802 33254 26898 33270
rect 26342 32843 26662 33221
rect 26802 33190 26818 33254
rect 26882 33190 26898 33254
rect 27061 33534 27383 33543
rect 27061 33230 27070 33534
rect 27374 33230 27383 33534
rect 27061 33221 27383 33230
rect 27521 33510 27537 33574
rect 27601 33510 27617 33574
rect 28240 33654 28336 33670
rect 28240 33590 28256 33654
rect 28320 33590 28336 33654
rect 28240 33574 28336 33590
rect 27782 33543 28102 33562
rect 27521 33494 27617 33510
rect 27521 33430 27537 33494
rect 27601 33430 27617 33494
rect 27521 33414 27617 33430
rect 27521 33350 27537 33414
rect 27601 33350 27617 33414
rect 27521 33334 27617 33350
rect 27521 33270 27537 33334
rect 27601 33270 27617 33334
rect 27521 33254 27617 33270
rect 26802 33174 26898 33190
rect 26802 33110 26818 33174
rect 26882 33110 26898 33174
rect 26802 33094 26898 33110
rect 26802 32954 26898 32970
rect 26802 32890 26818 32954
rect 26882 32890 26898 32954
rect 26802 32874 26898 32890
rect 26342 32834 26664 32843
rect 26342 32530 26351 32834
rect 26655 32530 26664 32834
rect 26342 32521 26664 32530
rect 26802 32810 26818 32874
rect 26882 32810 26898 32874
rect 27062 32843 27382 33221
rect 27521 33190 27537 33254
rect 27601 33190 27617 33254
rect 27780 33534 28102 33543
rect 27780 33230 27789 33534
rect 28093 33230 28102 33534
rect 27780 33221 28102 33230
rect 27521 33174 27617 33190
rect 27521 33110 27537 33174
rect 27601 33110 27617 33174
rect 27521 33094 27617 33110
rect 27521 32954 27617 32970
rect 27521 32890 27537 32954
rect 27601 32890 27617 32954
rect 27521 32874 27617 32890
rect 26802 32794 26898 32810
rect 26802 32730 26818 32794
rect 26882 32730 26898 32794
rect 26802 32714 26898 32730
rect 26802 32650 26818 32714
rect 26882 32650 26898 32714
rect 26802 32634 26898 32650
rect 26802 32570 26818 32634
rect 26882 32570 26898 32634
rect 26802 32554 26898 32570
rect 26342 32282 26662 32521
rect 26802 32490 26818 32554
rect 26882 32490 26898 32554
rect 27061 32834 27383 32843
rect 27061 32530 27070 32834
rect 27374 32530 27383 32834
rect 27061 32521 27383 32530
rect 27521 32810 27537 32874
rect 27601 32810 27617 32874
rect 27782 32843 28102 33221
rect 28240 33510 28256 33574
rect 28320 33510 28336 33574
rect 28959 33654 29055 33670
rect 28959 33590 28975 33654
rect 29039 33590 29055 33654
rect 28959 33574 29055 33590
rect 28502 33543 28822 33562
rect 28240 33494 28336 33510
rect 28240 33430 28256 33494
rect 28320 33430 28336 33494
rect 28240 33414 28336 33430
rect 28240 33350 28256 33414
rect 28320 33350 28336 33414
rect 28240 33334 28336 33350
rect 28240 33270 28256 33334
rect 28320 33270 28336 33334
rect 28240 33254 28336 33270
rect 28240 33190 28256 33254
rect 28320 33190 28336 33254
rect 28499 33534 28822 33543
rect 28499 33230 28508 33534
rect 28812 33230 28822 33534
rect 28499 33221 28822 33230
rect 28240 33174 28336 33190
rect 28240 33110 28256 33174
rect 28320 33110 28336 33174
rect 28240 33094 28336 33110
rect 27521 32794 27617 32810
rect 27521 32730 27537 32794
rect 27601 32730 27617 32794
rect 27521 32714 27617 32730
rect 27521 32650 27537 32714
rect 27601 32650 27617 32714
rect 27521 32634 27617 32650
rect 27521 32570 27537 32634
rect 27601 32570 27617 32634
rect 27521 32554 27617 32570
rect 26802 32474 26898 32490
rect 26802 32410 26818 32474
rect 26882 32410 26898 32474
rect 26802 32394 26898 32410
rect 27062 32282 27382 32521
rect 27521 32490 27537 32554
rect 27601 32490 27617 32554
rect 27780 32834 28102 32843
rect 27780 32530 27789 32834
rect 28093 32530 28102 32834
rect 27780 32521 28102 32530
rect 27521 32474 27617 32490
rect 27521 32410 27537 32474
rect 27601 32410 27617 32474
rect 27521 32394 27617 32410
rect 27782 32282 28102 32521
rect 28240 32954 28336 32970
rect 28240 32890 28256 32954
rect 28320 32890 28336 32954
rect 28240 32874 28336 32890
rect 28240 32810 28256 32874
rect 28320 32810 28336 32874
rect 28502 32843 28822 33221
rect 28959 33510 28975 33574
rect 29039 33510 29055 33574
rect 29678 33654 29774 33670
rect 29678 33590 29694 33654
rect 29758 33590 29774 33654
rect 29678 33574 29774 33590
rect 29222 33543 29542 33562
rect 28959 33494 29055 33510
rect 28959 33430 28975 33494
rect 29039 33430 29055 33494
rect 28959 33414 29055 33430
rect 28959 33350 28975 33414
rect 29039 33350 29055 33414
rect 28959 33334 29055 33350
rect 28959 33270 28975 33334
rect 29039 33270 29055 33334
rect 28959 33254 29055 33270
rect 28959 33190 28975 33254
rect 29039 33190 29055 33254
rect 29218 33534 29542 33543
rect 29218 33230 29227 33534
rect 29531 33230 29542 33534
rect 29218 33221 29542 33230
rect 28959 33174 29055 33190
rect 28959 33110 28975 33174
rect 29039 33110 29055 33174
rect 28959 33094 29055 33110
rect 28240 32794 28336 32810
rect 28240 32730 28256 32794
rect 28320 32730 28336 32794
rect 28240 32714 28336 32730
rect 28240 32650 28256 32714
rect 28320 32650 28336 32714
rect 28240 32634 28336 32650
rect 28240 32570 28256 32634
rect 28320 32570 28336 32634
rect 28240 32554 28336 32570
rect 28240 32490 28256 32554
rect 28320 32490 28336 32554
rect 28499 32834 28822 32843
rect 28499 32530 28508 32834
rect 28812 32530 28822 32834
rect 28499 32521 28822 32530
rect 28240 32474 28336 32490
rect 28240 32410 28256 32474
rect 28320 32410 28336 32474
rect 28240 32394 28336 32410
rect 28502 32282 28822 32521
rect 28959 32954 29055 32970
rect 28959 32890 28975 32954
rect 29039 32890 29055 32954
rect 28959 32874 29055 32890
rect 28959 32810 28975 32874
rect 29039 32810 29055 32874
rect 29222 32843 29542 33221
rect 29678 33510 29694 33574
rect 29758 33510 29774 33574
rect 30397 33654 30493 33670
rect 30397 33590 30413 33654
rect 30477 33590 30493 33654
rect 30397 33574 30493 33590
rect 29942 33543 30262 33562
rect 29678 33494 29774 33510
rect 29678 33430 29694 33494
rect 29758 33430 29774 33494
rect 29678 33414 29774 33430
rect 29678 33350 29694 33414
rect 29758 33350 29774 33414
rect 29678 33334 29774 33350
rect 29678 33270 29694 33334
rect 29758 33270 29774 33334
rect 29678 33254 29774 33270
rect 29678 33190 29694 33254
rect 29758 33190 29774 33254
rect 29937 33534 30262 33543
rect 29937 33230 29946 33534
rect 30250 33230 30262 33534
rect 29937 33221 30262 33230
rect 29678 33174 29774 33190
rect 29678 33110 29694 33174
rect 29758 33110 29774 33174
rect 29678 33094 29774 33110
rect 28959 32794 29055 32810
rect 28959 32730 28975 32794
rect 29039 32730 29055 32794
rect 28959 32714 29055 32730
rect 28959 32650 28975 32714
rect 29039 32650 29055 32714
rect 28959 32634 29055 32650
rect 28959 32570 28975 32634
rect 29039 32570 29055 32634
rect 28959 32554 29055 32570
rect 28959 32490 28975 32554
rect 29039 32490 29055 32554
rect 29218 32834 29542 32843
rect 29218 32530 29227 32834
rect 29531 32530 29542 32834
rect 29218 32521 29542 32530
rect 28959 32474 29055 32490
rect 28959 32410 28975 32474
rect 29039 32410 29055 32474
rect 28959 32394 29055 32410
rect 29222 32282 29542 32521
rect 29678 32954 29774 32970
rect 29678 32890 29694 32954
rect 29758 32890 29774 32954
rect 29678 32874 29774 32890
rect 29678 32810 29694 32874
rect 29758 32810 29774 32874
rect 29942 32843 30262 33221
rect 30397 33510 30413 33574
rect 30477 33510 30493 33574
rect 31116 33654 31212 33670
rect 31116 33590 31132 33654
rect 31196 33590 31212 33654
rect 31116 33574 31212 33590
rect 30662 33543 30982 33562
rect 30397 33494 30493 33510
rect 30397 33430 30413 33494
rect 30477 33430 30493 33494
rect 30397 33414 30493 33430
rect 30397 33350 30413 33414
rect 30477 33350 30493 33414
rect 30397 33334 30493 33350
rect 30397 33270 30413 33334
rect 30477 33270 30493 33334
rect 30397 33254 30493 33270
rect 30397 33190 30413 33254
rect 30477 33190 30493 33254
rect 30656 33534 30982 33543
rect 30656 33230 30665 33534
rect 30969 33230 30982 33534
rect 30656 33221 30982 33230
rect 30397 33174 30493 33190
rect 30397 33110 30413 33174
rect 30477 33110 30493 33174
rect 30397 33094 30493 33110
rect 29678 32794 29774 32810
rect 29678 32730 29694 32794
rect 29758 32730 29774 32794
rect 29678 32714 29774 32730
rect 29678 32650 29694 32714
rect 29758 32650 29774 32714
rect 29678 32634 29774 32650
rect 29678 32570 29694 32634
rect 29758 32570 29774 32634
rect 29678 32554 29774 32570
rect 29678 32490 29694 32554
rect 29758 32490 29774 32554
rect 29937 32834 30262 32843
rect 29937 32530 29946 32834
rect 30250 32530 30262 32834
rect 29937 32521 30262 32530
rect 29678 32474 29774 32490
rect 29678 32410 29694 32474
rect 29758 32410 29774 32474
rect 29678 32394 29774 32410
rect 29942 32282 30262 32521
rect 30397 32954 30493 32970
rect 30397 32890 30413 32954
rect 30477 32890 30493 32954
rect 30397 32874 30493 32890
rect 30397 32810 30413 32874
rect 30477 32810 30493 32874
rect 30662 32843 30982 33221
rect 31116 33510 31132 33574
rect 31196 33510 31212 33574
rect 31835 33654 31931 33670
rect 31835 33590 31851 33654
rect 31915 33590 31931 33654
rect 31835 33574 31931 33590
rect 31382 33543 31702 33562
rect 31116 33494 31212 33510
rect 31116 33430 31132 33494
rect 31196 33430 31212 33494
rect 31116 33414 31212 33430
rect 31116 33350 31132 33414
rect 31196 33350 31212 33414
rect 31116 33334 31212 33350
rect 31116 33270 31132 33334
rect 31196 33270 31212 33334
rect 31116 33254 31212 33270
rect 31116 33190 31132 33254
rect 31196 33190 31212 33254
rect 31375 33534 31702 33543
rect 31375 33230 31384 33534
rect 31688 33230 31702 33534
rect 31375 33221 31702 33230
rect 31116 33174 31212 33190
rect 31116 33110 31132 33174
rect 31196 33110 31212 33174
rect 31116 33094 31212 33110
rect 30397 32794 30493 32810
rect 30397 32730 30413 32794
rect 30477 32730 30493 32794
rect 30397 32714 30493 32730
rect 30397 32650 30413 32714
rect 30477 32650 30493 32714
rect 30397 32634 30493 32650
rect 30397 32570 30413 32634
rect 30477 32570 30493 32634
rect 30397 32554 30493 32570
rect 30397 32490 30413 32554
rect 30477 32490 30493 32554
rect 30656 32834 30982 32843
rect 30656 32530 30665 32834
rect 30969 32530 30982 32834
rect 30656 32521 30982 32530
rect 30397 32474 30493 32490
rect 30397 32410 30413 32474
rect 30477 32410 30493 32474
rect 30397 32394 30493 32410
rect 30662 32282 30982 32521
rect 31116 32954 31212 32970
rect 31116 32890 31132 32954
rect 31196 32890 31212 32954
rect 31116 32874 31212 32890
rect 31116 32810 31132 32874
rect 31196 32810 31212 32874
rect 31382 32843 31702 33221
rect 31835 33510 31851 33574
rect 31915 33510 31931 33574
rect 32554 33654 32650 33670
rect 32554 33590 32570 33654
rect 32634 33590 32650 33654
rect 32554 33574 32650 33590
rect 32102 33543 32422 33562
rect 31835 33494 31931 33510
rect 31835 33430 31851 33494
rect 31915 33430 31931 33494
rect 31835 33414 31931 33430
rect 31835 33350 31851 33414
rect 31915 33350 31931 33414
rect 31835 33334 31931 33350
rect 31835 33270 31851 33334
rect 31915 33270 31931 33334
rect 31835 33254 31931 33270
rect 31835 33190 31851 33254
rect 31915 33190 31931 33254
rect 32094 33534 32422 33543
rect 32094 33230 32103 33534
rect 32407 33230 32422 33534
rect 32094 33221 32422 33230
rect 31835 33174 31931 33190
rect 31835 33110 31851 33174
rect 31915 33110 31931 33174
rect 31835 33094 31931 33110
rect 31116 32794 31212 32810
rect 31116 32730 31132 32794
rect 31196 32730 31212 32794
rect 31116 32714 31212 32730
rect 31116 32650 31132 32714
rect 31196 32650 31212 32714
rect 31116 32634 31212 32650
rect 31116 32570 31132 32634
rect 31196 32570 31212 32634
rect 31116 32554 31212 32570
rect 31116 32490 31132 32554
rect 31196 32490 31212 32554
rect 31375 32834 31702 32843
rect 31375 32530 31384 32834
rect 31688 32530 31702 32834
rect 31375 32521 31702 32530
rect 31116 32474 31212 32490
rect 31116 32410 31132 32474
rect 31196 32410 31212 32474
rect 31116 32394 31212 32410
rect 31382 32282 31702 32521
rect 31835 32954 31931 32970
rect 31835 32890 31851 32954
rect 31915 32890 31931 32954
rect 31835 32874 31931 32890
rect 31835 32810 31851 32874
rect 31915 32810 31931 32874
rect 32102 32843 32422 33221
rect 32554 33510 32570 33574
rect 32634 33510 32650 33574
rect 32998 33562 33058 35922
rect 33271 33838 33337 33839
rect 33271 33774 33272 33838
rect 33336 33774 33337 33838
rect 33271 33773 33337 33774
rect 34099 33838 34165 33839
rect 34099 33774 34100 33838
rect 34164 33836 34165 33838
rect 34164 33776 34334 33836
rect 34164 33774 34165 33776
rect 34099 33773 34165 33774
rect 33274 33670 33334 33773
rect 34274 33670 34334 33776
rect 33273 33654 33369 33670
rect 33273 33590 33289 33654
rect 33353 33590 33369 33654
rect 33273 33574 33369 33590
rect 32822 33543 33142 33562
rect 32554 33494 32650 33510
rect 32554 33430 32570 33494
rect 32634 33430 32650 33494
rect 32554 33414 32650 33430
rect 32554 33350 32570 33414
rect 32634 33350 32650 33414
rect 32554 33334 32650 33350
rect 32554 33270 32570 33334
rect 32634 33270 32650 33334
rect 32554 33254 32650 33270
rect 32554 33190 32570 33254
rect 32634 33190 32650 33254
rect 32813 33534 33142 33543
rect 32813 33230 32822 33534
rect 33126 33230 33142 33534
rect 32813 33221 33142 33230
rect 32554 33174 32650 33190
rect 32554 33110 32570 33174
rect 32634 33110 32650 33174
rect 32554 33094 32650 33110
rect 31835 32794 31931 32810
rect 31835 32730 31851 32794
rect 31915 32730 31931 32794
rect 31835 32714 31931 32730
rect 31835 32650 31851 32714
rect 31915 32650 31931 32714
rect 31835 32634 31931 32650
rect 31835 32570 31851 32634
rect 31915 32570 31931 32634
rect 31835 32554 31931 32570
rect 31835 32490 31851 32554
rect 31915 32490 31931 32554
rect 32094 32834 32422 32843
rect 32094 32530 32103 32834
rect 32407 32530 32422 32834
rect 32094 32521 32422 32530
rect 31835 32474 31931 32490
rect 31835 32410 31851 32474
rect 31915 32410 31931 32474
rect 31835 32394 31931 32410
rect 32102 32282 32422 32521
rect 32554 32954 32650 32970
rect 32554 32890 32570 32954
rect 32634 32890 32650 32954
rect 32554 32874 32650 32890
rect 32554 32810 32570 32874
rect 32634 32810 32650 32874
rect 32822 32843 33142 33221
rect 33273 33510 33289 33574
rect 33353 33510 33369 33574
rect 34250 33654 34346 33670
rect 34250 33590 34266 33654
rect 34330 33590 34346 33654
rect 34250 33574 34346 33590
rect 33273 33494 33369 33510
rect 33273 33430 33289 33494
rect 33353 33430 33369 33494
rect 33273 33414 33369 33430
rect 33273 33350 33289 33414
rect 33353 33350 33369 33414
rect 33273 33334 33369 33350
rect 33273 33270 33289 33334
rect 33353 33270 33369 33334
rect 33273 33254 33369 33270
rect 33273 33190 33289 33254
rect 33353 33190 33369 33254
rect 33273 33174 33369 33190
rect 33273 33110 33289 33174
rect 33353 33110 33369 33174
rect 33273 33094 33369 33110
rect 33790 33543 34110 33562
rect 33790 33534 34112 33543
rect 33790 33230 33799 33534
rect 34103 33230 34112 33534
rect 33790 33221 34112 33230
rect 34250 33510 34266 33574
rect 34330 33510 34346 33574
rect 34969 33654 35065 33670
rect 34969 33590 34985 33654
rect 35049 33590 35065 33654
rect 34969 33574 35065 33590
rect 34510 33543 34830 33562
rect 34250 33494 34346 33510
rect 34250 33430 34266 33494
rect 34330 33430 34346 33494
rect 34250 33414 34346 33430
rect 34250 33350 34266 33414
rect 34330 33350 34346 33414
rect 34250 33334 34346 33350
rect 34250 33270 34266 33334
rect 34330 33270 34346 33334
rect 34250 33254 34346 33270
rect 32554 32794 32650 32810
rect 32554 32730 32570 32794
rect 32634 32730 32650 32794
rect 32554 32714 32650 32730
rect 32554 32650 32570 32714
rect 32634 32650 32650 32714
rect 32554 32634 32650 32650
rect 32554 32570 32570 32634
rect 32634 32570 32650 32634
rect 32554 32554 32650 32570
rect 32554 32490 32570 32554
rect 32634 32490 32650 32554
rect 32813 32834 33142 32843
rect 32813 32530 32822 32834
rect 33126 32530 33142 32834
rect 32813 32521 33142 32530
rect 32554 32474 32650 32490
rect 32554 32410 32570 32474
rect 32634 32410 32650 32474
rect 32554 32394 32650 32410
rect 32822 32282 33142 32521
rect 33273 32954 33369 32970
rect 33273 32890 33289 32954
rect 33353 32890 33369 32954
rect 33273 32874 33369 32890
rect 33273 32810 33289 32874
rect 33353 32810 33369 32874
rect 33273 32794 33369 32810
rect 33273 32730 33289 32794
rect 33353 32730 33369 32794
rect 33273 32714 33369 32730
rect 33273 32650 33289 32714
rect 33353 32650 33369 32714
rect 33273 32634 33369 32650
rect 33273 32570 33289 32634
rect 33353 32570 33369 32634
rect 33273 32554 33369 32570
rect 33273 32490 33289 32554
rect 33353 32490 33369 32554
rect 33273 32474 33369 32490
rect 33273 32410 33289 32474
rect 33353 32410 33369 32474
rect 33273 32394 33369 32410
rect 33790 32843 34110 33221
rect 34250 33190 34266 33254
rect 34330 33190 34346 33254
rect 34509 33534 34831 33543
rect 34509 33230 34518 33534
rect 34822 33230 34831 33534
rect 34509 33221 34831 33230
rect 34969 33510 34985 33574
rect 35049 33510 35065 33574
rect 35688 33654 35784 33670
rect 35688 33590 35704 33654
rect 35768 33590 35784 33654
rect 35688 33574 35784 33590
rect 35230 33543 35550 33562
rect 34969 33494 35065 33510
rect 34969 33430 34985 33494
rect 35049 33430 35065 33494
rect 34969 33414 35065 33430
rect 34969 33350 34985 33414
rect 35049 33350 35065 33414
rect 34969 33334 35065 33350
rect 34969 33270 34985 33334
rect 35049 33270 35065 33334
rect 34969 33254 35065 33270
rect 34250 33174 34346 33190
rect 34250 33110 34266 33174
rect 34330 33110 34346 33174
rect 34250 33094 34346 33110
rect 34250 32954 34346 32970
rect 34250 32890 34266 32954
rect 34330 32890 34346 32954
rect 34250 32874 34346 32890
rect 33790 32834 34112 32843
rect 33790 32530 33799 32834
rect 34103 32530 34112 32834
rect 33790 32521 34112 32530
rect 34250 32810 34266 32874
rect 34330 32810 34346 32874
rect 34510 32843 34830 33221
rect 34969 33190 34985 33254
rect 35049 33190 35065 33254
rect 35228 33534 35550 33543
rect 35228 33230 35237 33534
rect 35541 33230 35550 33534
rect 35228 33221 35550 33230
rect 34969 33174 35065 33190
rect 34969 33110 34985 33174
rect 35049 33110 35065 33174
rect 34969 33094 35065 33110
rect 34969 32954 35065 32970
rect 34969 32890 34985 32954
rect 35049 32890 35065 32954
rect 34969 32874 35065 32890
rect 34250 32794 34346 32810
rect 34250 32730 34266 32794
rect 34330 32730 34346 32794
rect 34250 32714 34346 32730
rect 34250 32650 34266 32714
rect 34330 32650 34346 32714
rect 34250 32634 34346 32650
rect 34250 32570 34266 32634
rect 34330 32570 34346 32634
rect 34250 32554 34346 32570
rect 33790 32282 34110 32521
rect 34250 32490 34266 32554
rect 34330 32490 34346 32554
rect 34509 32834 34831 32843
rect 34509 32530 34518 32834
rect 34822 32530 34831 32834
rect 34509 32521 34831 32530
rect 34969 32810 34985 32874
rect 35049 32810 35065 32874
rect 35230 32843 35550 33221
rect 35688 33510 35704 33574
rect 35768 33510 35784 33574
rect 36407 33654 36503 33670
rect 36407 33590 36423 33654
rect 36487 33590 36503 33654
rect 36407 33574 36503 33590
rect 35950 33543 36270 33562
rect 35688 33494 35784 33510
rect 35688 33430 35704 33494
rect 35768 33430 35784 33494
rect 35688 33414 35784 33430
rect 35688 33350 35704 33414
rect 35768 33350 35784 33414
rect 35688 33334 35784 33350
rect 35688 33270 35704 33334
rect 35768 33270 35784 33334
rect 35688 33254 35784 33270
rect 35688 33190 35704 33254
rect 35768 33190 35784 33254
rect 35947 33534 36270 33543
rect 35947 33230 35956 33534
rect 36260 33230 36270 33534
rect 35947 33221 36270 33230
rect 35688 33174 35784 33190
rect 35688 33110 35704 33174
rect 35768 33110 35784 33174
rect 35688 33094 35784 33110
rect 34969 32794 35065 32810
rect 34969 32730 34985 32794
rect 35049 32730 35065 32794
rect 34969 32714 35065 32730
rect 34969 32650 34985 32714
rect 35049 32650 35065 32714
rect 34969 32634 35065 32650
rect 34969 32570 34985 32634
rect 35049 32570 35065 32634
rect 34969 32554 35065 32570
rect 34250 32474 34346 32490
rect 34250 32410 34266 32474
rect 34330 32410 34346 32474
rect 34250 32394 34346 32410
rect 34510 32282 34830 32521
rect 34969 32490 34985 32554
rect 35049 32490 35065 32554
rect 35228 32834 35550 32843
rect 35228 32530 35237 32834
rect 35541 32530 35550 32834
rect 35228 32521 35550 32530
rect 34969 32474 35065 32490
rect 34969 32410 34985 32474
rect 35049 32410 35065 32474
rect 34969 32394 35065 32410
rect 35230 32282 35550 32521
rect 35688 32954 35784 32970
rect 35688 32890 35704 32954
rect 35768 32890 35784 32954
rect 35688 32874 35784 32890
rect 35688 32810 35704 32874
rect 35768 32810 35784 32874
rect 35950 32843 36270 33221
rect 36407 33510 36423 33574
rect 36487 33510 36503 33574
rect 37126 33654 37222 33670
rect 37126 33590 37142 33654
rect 37206 33590 37222 33654
rect 37126 33574 37222 33590
rect 36670 33543 36990 33562
rect 36407 33494 36503 33510
rect 36407 33430 36423 33494
rect 36487 33430 36503 33494
rect 36407 33414 36503 33430
rect 36407 33350 36423 33414
rect 36487 33350 36503 33414
rect 36407 33334 36503 33350
rect 36407 33270 36423 33334
rect 36487 33270 36503 33334
rect 36407 33254 36503 33270
rect 36407 33190 36423 33254
rect 36487 33190 36503 33254
rect 36666 33534 36990 33543
rect 36666 33230 36675 33534
rect 36979 33230 36990 33534
rect 36666 33221 36990 33230
rect 36407 33174 36503 33190
rect 36407 33110 36423 33174
rect 36487 33110 36503 33174
rect 36407 33094 36503 33110
rect 35688 32794 35784 32810
rect 35688 32730 35704 32794
rect 35768 32730 35784 32794
rect 35688 32714 35784 32730
rect 35688 32650 35704 32714
rect 35768 32650 35784 32714
rect 35688 32634 35784 32650
rect 35688 32570 35704 32634
rect 35768 32570 35784 32634
rect 35688 32554 35784 32570
rect 35688 32490 35704 32554
rect 35768 32490 35784 32554
rect 35947 32834 36270 32843
rect 35947 32530 35956 32834
rect 36260 32530 36270 32834
rect 35947 32521 36270 32530
rect 35688 32474 35784 32490
rect 35688 32410 35704 32474
rect 35768 32410 35784 32474
rect 35688 32394 35784 32410
rect 35950 32282 36270 32521
rect 36407 32954 36503 32970
rect 36407 32890 36423 32954
rect 36487 32890 36503 32954
rect 36407 32874 36503 32890
rect 36407 32810 36423 32874
rect 36487 32810 36503 32874
rect 36670 32843 36990 33221
rect 37126 33510 37142 33574
rect 37206 33510 37222 33574
rect 37552 33562 37612 35969
rect 53456 33944 55088 37640
rect 53456 33880 53480 33944
rect 53544 33880 53560 33944
rect 53624 33880 53640 33944
rect 53704 33880 53720 33944
rect 53784 33880 53800 33944
rect 53864 33880 53880 33944
rect 53944 33880 53960 33944
rect 54024 33880 54040 33944
rect 54104 33880 54120 33944
rect 54184 33880 54200 33944
rect 54264 33880 54280 33944
rect 54344 33880 54360 33944
rect 54424 33880 54440 33944
rect 54504 33880 54520 33944
rect 54584 33880 54600 33944
rect 54664 33880 54680 33944
rect 54744 33880 54760 33944
rect 54824 33880 54840 33944
rect 54904 33880 54920 33944
rect 54984 33880 55000 33944
rect 55064 33880 55088 33944
rect 37845 33654 37941 33670
rect 37845 33590 37861 33654
rect 37925 33590 37941 33654
rect 37845 33574 37941 33590
rect 37390 33543 37710 33562
rect 37126 33494 37222 33510
rect 37126 33430 37142 33494
rect 37206 33430 37222 33494
rect 37126 33414 37222 33430
rect 37126 33350 37142 33414
rect 37206 33350 37222 33414
rect 37126 33334 37222 33350
rect 37126 33270 37142 33334
rect 37206 33270 37222 33334
rect 37126 33254 37222 33270
rect 37126 33190 37142 33254
rect 37206 33190 37222 33254
rect 37385 33534 37710 33543
rect 37385 33230 37394 33534
rect 37698 33230 37710 33534
rect 37385 33221 37710 33230
rect 37126 33174 37222 33190
rect 37126 33110 37142 33174
rect 37206 33110 37222 33174
rect 37126 33094 37222 33110
rect 36407 32794 36503 32810
rect 36407 32730 36423 32794
rect 36487 32730 36503 32794
rect 36407 32714 36503 32730
rect 36407 32650 36423 32714
rect 36487 32650 36503 32714
rect 36407 32634 36503 32650
rect 36407 32570 36423 32634
rect 36487 32570 36503 32634
rect 36407 32554 36503 32570
rect 36407 32490 36423 32554
rect 36487 32490 36503 32554
rect 36666 32834 36990 32843
rect 36666 32530 36675 32834
rect 36979 32530 36990 32834
rect 36666 32521 36990 32530
rect 36407 32474 36503 32490
rect 36407 32410 36423 32474
rect 36487 32410 36503 32474
rect 36407 32394 36503 32410
rect 36670 32282 36990 32521
rect 37126 32954 37222 32970
rect 37126 32890 37142 32954
rect 37206 32890 37222 32954
rect 37126 32874 37222 32890
rect 37126 32810 37142 32874
rect 37206 32810 37222 32874
rect 37390 32843 37710 33221
rect 37845 33510 37861 33574
rect 37925 33510 37941 33574
rect 38564 33654 38660 33670
rect 38564 33590 38580 33654
rect 38644 33590 38660 33654
rect 38564 33574 38660 33590
rect 38110 33543 38430 33562
rect 37845 33494 37941 33510
rect 37845 33430 37861 33494
rect 37925 33430 37941 33494
rect 37845 33414 37941 33430
rect 37845 33350 37861 33414
rect 37925 33350 37941 33414
rect 37845 33334 37941 33350
rect 37845 33270 37861 33334
rect 37925 33270 37941 33334
rect 37845 33254 37941 33270
rect 37845 33190 37861 33254
rect 37925 33190 37941 33254
rect 38104 33534 38430 33543
rect 38104 33230 38113 33534
rect 38417 33230 38430 33534
rect 38104 33221 38430 33230
rect 37845 33174 37941 33190
rect 37845 33110 37861 33174
rect 37925 33110 37941 33174
rect 37845 33094 37941 33110
rect 37126 32794 37222 32810
rect 37126 32730 37142 32794
rect 37206 32730 37222 32794
rect 37126 32714 37222 32730
rect 37126 32650 37142 32714
rect 37206 32650 37222 32714
rect 37126 32634 37222 32650
rect 37126 32570 37142 32634
rect 37206 32570 37222 32634
rect 37126 32554 37222 32570
rect 37126 32490 37142 32554
rect 37206 32490 37222 32554
rect 37385 32834 37710 32843
rect 37385 32530 37394 32834
rect 37698 32530 37710 32834
rect 37385 32521 37710 32530
rect 37126 32474 37222 32490
rect 37126 32410 37142 32474
rect 37206 32410 37222 32474
rect 37126 32394 37222 32410
rect 37390 32282 37710 32521
rect 37845 32954 37941 32970
rect 37845 32890 37861 32954
rect 37925 32890 37941 32954
rect 37845 32874 37941 32890
rect 37845 32810 37861 32874
rect 37925 32810 37941 32874
rect 38110 32843 38430 33221
rect 38564 33510 38580 33574
rect 38644 33510 38660 33574
rect 39283 33654 39379 33670
rect 39283 33590 39299 33654
rect 39363 33590 39379 33654
rect 39283 33574 39379 33590
rect 38830 33543 39150 33562
rect 38564 33494 38660 33510
rect 38564 33430 38580 33494
rect 38644 33430 38660 33494
rect 38564 33414 38660 33430
rect 38564 33350 38580 33414
rect 38644 33350 38660 33414
rect 38564 33334 38660 33350
rect 38564 33270 38580 33334
rect 38644 33270 38660 33334
rect 38564 33254 38660 33270
rect 38564 33190 38580 33254
rect 38644 33190 38660 33254
rect 38823 33534 39150 33543
rect 38823 33230 38832 33534
rect 39136 33230 39150 33534
rect 38823 33221 39150 33230
rect 38564 33174 38660 33190
rect 38564 33110 38580 33174
rect 38644 33110 38660 33174
rect 38564 33094 38660 33110
rect 37845 32794 37941 32810
rect 37845 32730 37861 32794
rect 37925 32730 37941 32794
rect 37845 32714 37941 32730
rect 37845 32650 37861 32714
rect 37925 32650 37941 32714
rect 37845 32634 37941 32650
rect 37845 32570 37861 32634
rect 37925 32570 37941 32634
rect 37845 32554 37941 32570
rect 37845 32490 37861 32554
rect 37925 32490 37941 32554
rect 38104 32834 38430 32843
rect 38104 32530 38113 32834
rect 38417 32530 38430 32834
rect 38104 32521 38430 32530
rect 37845 32474 37941 32490
rect 37845 32410 37861 32474
rect 37925 32410 37941 32474
rect 37845 32394 37941 32410
rect 38110 32282 38430 32521
rect 38564 32954 38660 32970
rect 38564 32890 38580 32954
rect 38644 32890 38660 32954
rect 38564 32874 38660 32890
rect 38564 32810 38580 32874
rect 38644 32810 38660 32874
rect 38830 32843 39150 33221
rect 39283 33510 39299 33574
rect 39363 33510 39379 33574
rect 40002 33654 40098 33670
rect 40002 33590 40018 33654
rect 40082 33590 40098 33654
rect 40002 33574 40098 33590
rect 39550 33543 39870 33562
rect 39283 33494 39379 33510
rect 39283 33430 39299 33494
rect 39363 33430 39379 33494
rect 39283 33414 39379 33430
rect 39283 33350 39299 33414
rect 39363 33350 39379 33414
rect 39283 33334 39379 33350
rect 39283 33270 39299 33334
rect 39363 33270 39379 33334
rect 39283 33254 39379 33270
rect 39283 33190 39299 33254
rect 39363 33190 39379 33254
rect 39542 33534 39870 33543
rect 39542 33230 39551 33534
rect 39855 33230 39870 33534
rect 39542 33221 39870 33230
rect 39283 33174 39379 33190
rect 39283 33110 39299 33174
rect 39363 33110 39379 33174
rect 39283 33094 39379 33110
rect 38564 32794 38660 32810
rect 38564 32730 38580 32794
rect 38644 32730 38660 32794
rect 38564 32714 38660 32730
rect 38564 32650 38580 32714
rect 38644 32650 38660 32714
rect 38564 32634 38660 32650
rect 38564 32570 38580 32634
rect 38644 32570 38660 32634
rect 38564 32554 38660 32570
rect 38564 32490 38580 32554
rect 38644 32490 38660 32554
rect 38823 32834 39150 32843
rect 38823 32530 38832 32834
rect 39136 32530 39150 32834
rect 38823 32521 39150 32530
rect 38564 32474 38660 32490
rect 38564 32410 38580 32474
rect 38644 32410 38660 32474
rect 38564 32394 38660 32410
rect 38830 32282 39150 32521
rect 39283 32954 39379 32970
rect 39283 32890 39299 32954
rect 39363 32890 39379 32954
rect 39283 32874 39379 32890
rect 39283 32810 39299 32874
rect 39363 32810 39379 32874
rect 39550 32843 39870 33221
rect 40002 33510 40018 33574
rect 40082 33510 40098 33574
rect 40721 33654 40817 33670
rect 40721 33590 40737 33654
rect 40801 33590 40817 33654
rect 40721 33574 40817 33590
rect 40270 33543 40590 33562
rect 40002 33494 40098 33510
rect 40002 33430 40018 33494
rect 40082 33430 40098 33494
rect 40002 33414 40098 33430
rect 40002 33350 40018 33414
rect 40082 33350 40098 33414
rect 40002 33334 40098 33350
rect 40002 33270 40018 33334
rect 40082 33270 40098 33334
rect 40002 33254 40098 33270
rect 40002 33190 40018 33254
rect 40082 33190 40098 33254
rect 40261 33534 40590 33543
rect 40261 33230 40270 33534
rect 40574 33230 40590 33534
rect 40261 33221 40590 33230
rect 40002 33174 40098 33190
rect 40002 33110 40018 33174
rect 40082 33110 40098 33174
rect 40002 33094 40098 33110
rect 39283 32794 39379 32810
rect 39283 32730 39299 32794
rect 39363 32730 39379 32794
rect 39283 32714 39379 32730
rect 39283 32650 39299 32714
rect 39363 32650 39379 32714
rect 39283 32634 39379 32650
rect 39283 32570 39299 32634
rect 39363 32570 39379 32634
rect 39283 32554 39379 32570
rect 39283 32490 39299 32554
rect 39363 32490 39379 32554
rect 39542 32834 39870 32843
rect 39542 32530 39551 32834
rect 39855 32530 39870 32834
rect 39542 32521 39870 32530
rect 39283 32474 39379 32490
rect 39283 32410 39299 32474
rect 39363 32410 39379 32474
rect 39283 32394 39379 32410
rect 39550 32282 39870 32521
rect 40002 32954 40098 32970
rect 40002 32890 40018 32954
rect 40082 32890 40098 32954
rect 40002 32874 40098 32890
rect 40002 32810 40018 32874
rect 40082 32810 40098 32874
rect 40270 32843 40590 33221
rect 40721 33510 40737 33574
rect 40801 33510 40817 33574
rect 40721 33494 40817 33510
rect 40721 33430 40737 33494
rect 40801 33430 40817 33494
rect 40721 33414 40817 33430
rect 40721 33350 40737 33414
rect 40801 33350 40817 33414
rect 40721 33334 40817 33350
rect 40721 33270 40737 33334
rect 40801 33270 40817 33334
rect 40721 33254 40817 33270
rect 40721 33190 40737 33254
rect 40801 33190 40817 33254
rect 40721 33174 40817 33190
rect 40721 33110 40737 33174
rect 40801 33110 40817 33174
rect 40721 33094 40817 33110
rect 40002 32794 40098 32810
rect 40002 32730 40018 32794
rect 40082 32730 40098 32794
rect 40002 32714 40098 32730
rect 40002 32650 40018 32714
rect 40082 32650 40098 32714
rect 40002 32634 40098 32650
rect 40002 32570 40018 32634
rect 40082 32570 40098 32634
rect 40002 32554 40098 32570
rect 40002 32490 40018 32554
rect 40082 32490 40098 32554
rect 40261 32834 40590 32843
rect 40261 32530 40270 32834
rect 40574 32530 40590 32834
rect 40261 32521 40590 32530
rect 40002 32474 40098 32490
rect 40002 32410 40018 32474
rect 40082 32410 40098 32474
rect 40002 32394 40098 32410
rect 40270 32282 40590 32521
rect 40721 32954 40817 32970
rect 40721 32890 40737 32954
rect 40801 32890 40817 32954
rect 40721 32874 40817 32890
rect 40721 32810 40737 32874
rect 40801 32810 40817 32874
rect 40721 32794 40817 32810
rect 40721 32730 40737 32794
rect 40801 32730 40817 32794
rect 40721 32714 40817 32730
rect 40721 32650 40737 32714
rect 40801 32650 40817 32714
rect 40721 32634 40817 32650
rect 40721 32570 40737 32634
rect 40801 32570 40817 32634
rect 40721 32554 40817 32570
rect 40721 32490 40737 32554
rect 40801 32490 40817 32554
rect 40721 32474 40817 32490
rect 40721 32410 40737 32474
rect 40801 32410 40817 32474
rect 40721 32394 40817 32410
rect 26204 32254 33372 32282
rect 26204 32190 26232 32254
rect 26296 32190 26312 32254
rect 26376 32250 33372 32254
rect 33652 32254 40820 32282
rect 33652 32250 33680 32254
rect 26376 32190 33680 32250
rect 33744 32190 33760 32254
rect 33824 32190 40820 32254
rect 26204 32162 33372 32190
rect 33652 32162 40820 32190
rect 3348 30120 3372 30184
rect 3436 30120 3452 30184
rect 3516 30120 3532 30184
rect 3596 30120 3612 30184
rect 3676 30120 3692 30184
rect 3756 30120 3772 30184
rect 3836 30120 3852 30184
rect 3916 30120 3932 30184
rect 3996 30120 4012 30184
rect 4076 30120 4092 30184
rect 4156 30120 4172 30184
rect 4236 30120 4252 30184
rect 4316 30120 4332 30184
rect 4396 30120 4412 30184
rect 4476 30120 4492 30184
rect 4556 30120 4572 30184
rect 4636 30120 4652 30184
rect 4716 30120 4732 30184
rect 4796 30120 4812 30184
rect 4876 30120 4892 30184
rect 4956 30120 4980 30184
rect 3348 26424 4980 30120
rect 33409 30178 33475 30179
rect 33409 30114 33410 30178
rect 33474 30114 33475 30178
rect 33409 30113 33475 30114
rect 33412 29910 33472 30113
rect 30526 29894 30622 29910
rect 30526 29830 30542 29894
rect 30606 29830 30622 29894
rect 30526 29814 30622 29830
rect 30066 29783 30386 29802
rect 30066 29774 30388 29783
rect 30066 29470 30075 29774
rect 30379 29470 30388 29774
rect 30066 29461 30388 29470
rect 30526 29750 30542 29814
rect 30606 29750 30622 29814
rect 31245 29894 31341 29910
rect 31245 29830 31261 29894
rect 31325 29830 31341 29894
rect 31245 29814 31341 29830
rect 30786 29783 31106 29802
rect 30526 29734 30622 29750
rect 30526 29670 30542 29734
rect 30606 29670 30622 29734
rect 30526 29654 30622 29670
rect 30526 29590 30542 29654
rect 30606 29590 30622 29654
rect 30526 29574 30622 29590
rect 30526 29510 30542 29574
rect 30606 29510 30622 29574
rect 30526 29494 30622 29510
rect 30066 29083 30386 29461
rect 30526 29430 30542 29494
rect 30606 29430 30622 29494
rect 30785 29774 31107 29783
rect 30785 29470 30794 29774
rect 31098 29470 31107 29774
rect 30785 29461 31107 29470
rect 31245 29750 31261 29814
rect 31325 29750 31341 29814
rect 31964 29894 32060 29910
rect 31964 29830 31980 29894
rect 32044 29830 32060 29894
rect 31964 29814 32060 29830
rect 31506 29783 31826 29802
rect 31245 29734 31341 29750
rect 31245 29670 31261 29734
rect 31325 29670 31341 29734
rect 31245 29654 31341 29670
rect 31245 29590 31261 29654
rect 31325 29590 31341 29654
rect 31245 29574 31341 29590
rect 31245 29510 31261 29574
rect 31325 29510 31341 29574
rect 31245 29494 31341 29510
rect 30526 29414 30622 29430
rect 30526 29350 30542 29414
rect 30606 29350 30622 29414
rect 30526 29334 30622 29350
rect 30526 29194 30622 29210
rect 30526 29130 30542 29194
rect 30606 29130 30622 29194
rect 30526 29114 30622 29130
rect 30066 29074 30388 29083
rect 30066 28770 30075 29074
rect 30379 28770 30388 29074
rect 30066 28761 30388 28770
rect 30526 29050 30542 29114
rect 30606 29050 30622 29114
rect 30786 29083 31106 29461
rect 31245 29430 31261 29494
rect 31325 29430 31341 29494
rect 31504 29774 31826 29783
rect 31504 29470 31513 29774
rect 31817 29470 31826 29774
rect 31504 29461 31826 29470
rect 31245 29414 31341 29430
rect 31245 29350 31261 29414
rect 31325 29350 31341 29414
rect 31245 29334 31341 29350
rect 31245 29194 31341 29210
rect 31245 29130 31261 29194
rect 31325 29130 31341 29194
rect 31245 29114 31341 29130
rect 30526 29034 30622 29050
rect 30526 28970 30542 29034
rect 30606 28970 30622 29034
rect 30526 28954 30622 28970
rect 30526 28890 30542 28954
rect 30606 28890 30622 28954
rect 30526 28874 30622 28890
rect 30526 28810 30542 28874
rect 30606 28810 30622 28874
rect 30526 28794 30622 28810
rect 30066 28522 30386 28761
rect 30526 28730 30542 28794
rect 30606 28730 30622 28794
rect 30785 29074 31107 29083
rect 30785 28770 30794 29074
rect 31098 28770 31107 29074
rect 30785 28761 31107 28770
rect 31245 29050 31261 29114
rect 31325 29050 31341 29114
rect 31506 29083 31826 29461
rect 31964 29750 31980 29814
rect 32044 29750 32060 29814
rect 32683 29894 32779 29910
rect 32683 29830 32699 29894
rect 32763 29830 32779 29894
rect 32683 29814 32779 29830
rect 32226 29783 32546 29802
rect 31964 29734 32060 29750
rect 31964 29670 31980 29734
rect 32044 29670 32060 29734
rect 31964 29654 32060 29670
rect 31964 29590 31980 29654
rect 32044 29590 32060 29654
rect 31964 29574 32060 29590
rect 31964 29510 31980 29574
rect 32044 29510 32060 29574
rect 31964 29494 32060 29510
rect 31964 29430 31980 29494
rect 32044 29430 32060 29494
rect 32223 29774 32546 29783
rect 32223 29470 32232 29774
rect 32536 29470 32546 29774
rect 32223 29461 32546 29470
rect 31964 29414 32060 29430
rect 31964 29350 31980 29414
rect 32044 29350 32060 29414
rect 31964 29334 32060 29350
rect 31245 29034 31341 29050
rect 31245 28970 31261 29034
rect 31325 28970 31341 29034
rect 31245 28954 31341 28970
rect 31245 28890 31261 28954
rect 31325 28890 31341 28954
rect 31245 28874 31341 28890
rect 31245 28810 31261 28874
rect 31325 28810 31341 28874
rect 31245 28794 31341 28810
rect 30526 28714 30622 28730
rect 30526 28650 30542 28714
rect 30606 28650 30622 28714
rect 30526 28634 30622 28650
rect 30786 28522 31106 28761
rect 31245 28730 31261 28794
rect 31325 28730 31341 28794
rect 31504 29074 31826 29083
rect 31504 28770 31513 29074
rect 31817 28770 31826 29074
rect 31504 28761 31826 28770
rect 31245 28714 31341 28730
rect 31245 28650 31261 28714
rect 31325 28650 31341 28714
rect 31245 28634 31341 28650
rect 31506 28522 31826 28761
rect 31964 29194 32060 29210
rect 31964 29130 31980 29194
rect 32044 29130 32060 29194
rect 31964 29114 32060 29130
rect 31964 29050 31980 29114
rect 32044 29050 32060 29114
rect 32226 29083 32546 29461
rect 32683 29750 32699 29814
rect 32763 29750 32779 29814
rect 33402 29894 33498 29910
rect 33402 29830 33418 29894
rect 33482 29830 33498 29894
rect 33402 29814 33498 29830
rect 32946 29783 33266 29802
rect 32683 29734 32779 29750
rect 32683 29670 32699 29734
rect 32763 29670 32779 29734
rect 32683 29654 32779 29670
rect 32683 29590 32699 29654
rect 32763 29590 32779 29654
rect 32683 29574 32779 29590
rect 32683 29510 32699 29574
rect 32763 29510 32779 29574
rect 32683 29494 32779 29510
rect 32683 29430 32699 29494
rect 32763 29430 32779 29494
rect 32942 29774 33266 29783
rect 32942 29470 32951 29774
rect 33255 29470 33266 29774
rect 32942 29461 33266 29470
rect 32683 29414 32779 29430
rect 32683 29350 32699 29414
rect 32763 29350 32779 29414
rect 32683 29334 32779 29350
rect 31964 29034 32060 29050
rect 31964 28970 31980 29034
rect 32044 28970 32060 29034
rect 31964 28954 32060 28970
rect 31964 28890 31980 28954
rect 32044 28890 32060 28954
rect 31964 28874 32060 28890
rect 31964 28810 31980 28874
rect 32044 28810 32060 28874
rect 31964 28794 32060 28810
rect 31964 28730 31980 28794
rect 32044 28730 32060 28794
rect 32223 29074 32546 29083
rect 32223 28770 32232 29074
rect 32536 28770 32546 29074
rect 32223 28761 32546 28770
rect 31964 28714 32060 28730
rect 31964 28650 31980 28714
rect 32044 28650 32060 28714
rect 31964 28634 32060 28650
rect 32226 28522 32546 28761
rect 32683 29194 32779 29210
rect 32683 29130 32699 29194
rect 32763 29130 32779 29194
rect 32683 29114 32779 29130
rect 32683 29050 32699 29114
rect 32763 29050 32779 29114
rect 32946 29083 33266 29461
rect 33402 29750 33418 29814
rect 33482 29750 33498 29814
rect 33826 29802 33886 32162
rect 53456 30184 55088 33880
rect 53456 30120 53480 30184
rect 53544 30120 53560 30184
rect 53624 30120 53640 30184
rect 53704 30120 53720 30184
rect 53784 30120 53800 30184
rect 53864 30120 53880 30184
rect 53944 30120 53960 30184
rect 54024 30120 54040 30184
rect 54104 30120 54120 30184
rect 54184 30120 54200 30184
rect 54264 30120 54280 30184
rect 54344 30120 54360 30184
rect 54424 30120 54440 30184
rect 54504 30120 54520 30184
rect 54584 30120 54600 30184
rect 54664 30120 54680 30184
rect 54744 30120 54760 30184
rect 54824 30120 54840 30184
rect 54904 30120 54920 30184
rect 54984 30120 55000 30184
rect 55064 30120 55088 30184
rect 34121 29894 34217 29910
rect 34121 29830 34137 29894
rect 34201 29830 34217 29894
rect 34121 29814 34217 29830
rect 33666 29783 33986 29802
rect 33402 29734 33498 29750
rect 33402 29670 33418 29734
rect 33482 29670 33498 29734
rect 33402 29654 33498 29670
rect 33402 29590 33418 29654
rect 33482 29590 33498 29654
rect 33402 29574 33498 29590
rect 33402 29510 33418 29574
rect 33482 29510 33498 29574
rect 33402 29494 33498 29510
rect 33402 29430 33418 29494
rect 33482 29430 33498 29494
rect 33661 29774 33986 29783
rect 33661 29470 33670 29774
rect 33974 29470 33986 29774
rect 33661 29461 33986 29470
rect 33402 29414 33498 29430
rect 33402 29350 33418 29414
rect 33482 29350 33498 29414
rect 33402 29334 33498 29350
rect 32683 29034 32779 29050
rect 32683 28970 32699 29034
rect 32763 28970 32779 29034
rect 32683 28954 32779 28970
rect 32683 28890 32699 28954
rect 32763 28890 32779 28954
rect 32683 28874 32779 28890
rect 32683 28810 32699 28874
rect 32763 28810 32779 28874
rect 32683 28794 32779 28810
rect 32683 28730 32699 28794
rect 32763 28730 32779 28794
rect 32942 29074 33266 29083
rect 32942 28770 32951 29074
rect 33255 28770 33266 29074
rect 32942 28761 33266 28770
rect 32683 28714 32779 28730
rect 32683 28650 32699 28714
rect 32763 28650 32779 28714
rect 32683 28634 32779 28650
rect 32946 28522 33266 28761
rect 33402 29194 33498 29210
rect 33402 29130 33418 29194
rect 33482 29130 33498 29194
rect 33402 29114 33498 29130
rect 33402 29050 33418 29114
rect 33482 29050 33498 29114
rect 33666 29083 33986 29461
rect 34121 29750 34137 29814
rect 34201 29750 34217 29814
rect 34840 29894 34936 29910
rect 34840 29830 34856 29894
rect 34920 29830 34936 29894
rect 34840 29814 34936 29830
rect 34386 29783 34706 29802
rect 34121 29734 34217 29750
rect 34121 29670 34137 29734
rect 34201 29670 34217 29734
rect 34121 29654 34217 29670
rect 34121 29590 34137 29654
rect 34201 29590 34217 29654
rect 34121 29574 34217 29590
rect 34121 29510 34137 29574
rect 34201 29510 34217 29574
rect 34121 29494 34217 29510
rect 34121 29430 34137 29494
rect 34201 29430 34217 29494
rect 34380 29774 34706 29783
rect 34380 29470 34389 29774
rect 34693 29470 34706 29774
rect 34380 29461 34706 29470
rect 34121 29414 34217 29430
rect 34121 29350 34137 29414
rect 34201 29350 34217 29414
rect 34121 29334 34217 29350
rect 33402 29034 33498 29050
rect 33402 28970 33418 29034
rect 33482 28970 33498 29034
rect 33402 28954 33498 28970
rect 33402 28890 33418 28954
rect 33482 28890 33498 28954
rect 33402 28874 33498 28890
rect 33402 28810 33418 28874
rect 33482 28810 33498 28874
rect 33402 28794 33498 28810
rect 33402 28730 33418 28794
rect 33482 28730 33498 28794
rect 33661 29074 33986 29083
rect 33661 28770 33670 29074
rect 33974 28770 33986 29074
rect 33661 28761 33986 28770
rect 33402 28714 33498 28730
rect 33402 28650 33418 28714
rect 33482 28650 33498 28714
rect 33402 28634 33498 28650
rect 33666 28522 33986 28761
rect 34121 29194 34217 29210
rect 34121 29130 34137 29194
rect 34201 29130 34217 29194
rect 34121 29114 34217 29130
rect 34121 29050 34137 29114
rect 34201 29050 34217 29114
rect 34386 29083 34706 29461
rect 34840 29750 34856 29814
rect 34920 29750 34936 29814
rect 35559 29894 35655 29910
rect 35559 29830 35575 29894
rect 35639 29830 35655 29894
rect 35559 29814 35655 29830
rect 35106 29783 35426 29802
rect 34840 29734 34936 29750
rect 34840 29670 34856 29734
rect 34920 29670 34936 29734
rect 34840 29654 34936 29670
rect 34840 29590 34856 29654
rect 34920 29590 34936 29654
rect 34840 29574 34936 29590
rect 34840 29510 34856 29574
rect 34920 29510 34936 29574
rect 34840 29494 34936 29510
rect 34840 29430 34856 29494
rect 34920 29430 34936 29494
rect 35099 29774 35426 29783
rect 35099 29470 35108 29774
rect 35412 29470 35426 29774
rect 35099 29461 35426 29470
rect 34840 29414 34936 29430
rect 34840 29350 34856 29414
rect 34920 29350 34936 29414
rect 34840 29334 34936 29350
rect 34121 29034 34217 29050
rect 34121 28970 34137 29034
rect 34201 28970 34217 29034
rect 34121 28954 34217 28970
rect 34121 28890 34137 28954
rect 34201 28890 34217 28954
rect 34121 28874 34217 28890
rect 34121 28810 34137 28874
rect 34201 28810 34217 28874
rect 34121 28794 34217 28810
rect 34121 28730 34137 28794
rect 34201 28730 34217 28794
rect 34380 29074 34706 29083
rect 34380 28770 34389 29074
rect 34693 28770 34706 29074
rect 34380 28761 34706 28770
rect 34121 28714 34217 28730
rect 34121 28650 34137 28714
rect 34201 28650 34217 28714
rect 34121 28634 34217 28650
rect 34386 28522 34706 28761
rect 34840 29194 34936 29210
rect 34840 29130 34856 29194
rect 34920 29130 34936 29194
rect 34840 29114 34936 29130
rect 34840 29050 34856 29114
rect 34920 29050 34936 29114
rect 35106 29083 35426 29461
rect 35559 29750 35575 29814
rect 35639 29750 35655 29814
rect 36278 29894 36374 29910
rect 36278 29830 36294 29894
rect 36358 29830 36374 29894
rect 36278 29814 36374 29830
rect 35826 29783 36146 29802
rect 35559 29734 35655 29750
rect 35559 29670 35575 29734
rect 35639 29670 35655 29734
rect 35559 29654 35655 29670
rect 35559 29590 35575 29654
rect 35639 29590 35655 29654
rect 35559 29574 35655 29590
rect 35559 29510 35575 29574
rect 35639 29510 35655 29574
rect 35559 29494 35655 29510
rect 35559 29430 35575 29494
rect 35639 29430 35655 29494
rect 35818 29774 36146 29783
rect 35818 29470 35827 29774
rect 36131 29470 36146 29774
rect 35818 29461 36146 29470
rect 35559 29414 35655 29430
rect 35559 29350 35575 29414
rect 35639 29350 35655 29414
rect 35559 29334 35655 29350
rect 34840 29034 34936 29050
rect 34840 28970 34856 29034
rect 34920 28970 34936 29034
rect 34840 28954 34936 28970
rect 34840 28890 34856 28954
rect 34920 28890 34936 28954
rect 34840 28874 34936 28890
rect 34840 28810 34856 28874
rect 34920 28810 34936 28874
rect 34840 28794 34936 28810
rect 34840 28730 34856 28794
rect 34920 28730 34936 28794
rect 35099 29074 35426 29083
rect 35099 28770 35108 29074
rect 35412 28770 35426 29074
rect 35099 28761 35426 28770
rect 34840 28714 34936 28730
rect 34840 28650 34856 28714
rect 34920 28650 34936 28714
rect 34840 28634 34936 28650
rect 35106 28522 35426 28761
rect 35559 29194 35655 29210
rect 35559 29130 35575 29194
rect 35639 29130 35655 29194
rect 35559 29114 35655 29130
rect 35559 29050 35575 29114
rect 35639 29050 35655 29114
rect 35826 29083 36146 29461
rect 36278 29750 36294 29814
rect 36358 29750 36374 29814
rect 36997 29894 37093 29910
rect 36997 29830 37013 29894
rect 37077 29830 37093 29894
rect 36997 29814 37093 29830
rect 36546 29783 36866 29802
rect 36278 29734 36374 29750
rect 36278 29670 36294 29734
rect 36358 29670 36374 29734
rect 36278 29654 36374 29670
rect 36278 29590 36294 29654
rect 36358 29590 36374 29654
rect 36278 29574 36374 29590
rect 36278 29510 36294 29574
rect 36358 29510 36374 29574
rect 36278 29494 36374 29510
rect 36278 29430 36294 29494
rect 36358 29430 36374 29494
rect 36537 29774 36866 29783
rect 36537 29470 36546 29774
rect 36850 29470 36866 29774
rect 36537 29461 36866 29470
rect 36278 29414 36374 29430
rect 36278 29350 36294 29414
rect 36358 29350 36374 29414
rect 36278 29334 36374 29350
rect 35559 29034 35655 29050
rect 35559 28970 35575 29034
rect 35639 28970 35655 29034
rect 35559 28954 35655 28970
rect 35559 28890 35575 28954
rect 35639 28890 35655 28954
rect 35559 28874 35655 28890
rect 35559 28810 35575 28874
rect 35639 28810 35655 28874
rect 35559 28794 35655 28810
rect 35559 28730 35575 28794
rect 35639 28730 35655 28794
rect 35818 29074 36146 29083
rect 35818 28770 35827 29074
rect 36131 28770 36146 29074
rect 35818 28761 36146 28770
rect 35559 28714 35655 28730
rect 35559 28650 35575 28714
rect 35639 28650 35655 28714
rect 35559 28634 35655 28650
rect 35826 28522 36146 28761
rect 36278 29194 36374 29210
rect 36278 29130 36294 29194
rect 36358 29130 36374 29194
rect 36278 29114 36374 29130
rect 36278 29050 36294 29114
rect 36358 29050 36374 29114
rect 36546 29083 36866 29461
rect 36997 29750 37013 29814
rect 37077 29750 37093 29814
rect 36997 29734 37093 29750
rect 36997 29670 37013 29734
rect 37077 29670 37093 29734
rect 36997 29654 37093 29670
rect 36997 29590 37013 29654
rect 37077 29590 37093 29654
rect 36997 29574 37093 29590
rect 36997 29510 37013 29574
rect 37077 29510 37093 29574
rect 36997 29494 37093 29510
rect 36997 29430 37013 29494
rect 37077 29430 37093 29494
rect 36997 29414 37093 29430
rect 36997 29350 37013 29414
rect 37077 29350 37093 29414
rect 36997 29334 37093 29350
rect 36278 29034 36374 29050
rect 36278 28970 36294 29034
rect 36358 28970 36374 29034
rect 36278 28954 36374 28970
rect 36278 28890 36294 28954
rect 36358 28890 36374 28954
rect 36278 28874 36374 28890
rect 36278 28810 36294 28874
rect 36358 28810 36374 28874
rect 36278 28794 36374 28810
rect 36278 28730 36294 28794
rect 36358 28730 36374 28794
rect 36537 29074 36866 29083
rect 36537 28770 36546 29074
rect 36850 28770 36866 29074
rect 36537 28761 36866 28770
rect 36278 28714 36374 28730
rect 36278 28650 36294 28714
rect 36358 28650 36374 28714
rect 36278 28634 36374 28650
rect 36546 28522 36866 28761
rect 36997 29194 37093 29210
rect 36997 29130 37013 29194
rect 37077 29130 37093 29194
rect 36997 29114 37093 29130
rect 36997 29050 37013 29114
rect 37077 29050 37093 29114
rect 36997 29034 37093 29050
rect 36997 28970 37013 29034
rect 37077 28970 37093 29034
rect 36997 28954 37093 28970
rect 36997 28890 37013 28954
rect 37077 28890 37093 28954
rect 36997 28874 37093 28890
rect 36997 28810 37013 28874
rect 37077 28810 37093 28874
rect 36997 28794 37093 28810
rect 36997 28730 37013 28794
rect 37077 28730 37093 28794
rect 36997 28714 37093 28730
rect 36997 28650 37013 28714
rect 37077 28650 37093 28714
rect 36997 28634 37093 28650
rect 29928 28494 37096 28522
rect 29928 28430 29956 28494
rect 30020 28430 30036 28494
rect 30100 28430 37096 28494
rect 29928 28402 37096 28430
rect 3348 26360 3372 26424
rect 3436 26360 3452 26424
rect 3516 26360 3532 26424
rect 3596 26360 3612 26424
rect 3676 26360 3692 26424
rect 3756 26360 3772 26424
rect 3836 26360 3852 26424
rect 3916 26360 3932 26424
rect 3996 26360 4012 26424
rect 4076 26360 4092 26424
rect 4156 26360 4172 26424
rect 4236 26360 4252 26424
rect 4316 26360 4332 26424
rect 4396 26360 4412 26424
rect 4476 26360 4492 26424
rect 4556 26360 4572 26424
rect 4636 26360 4652 26424
rect 4716 26360 4732 26424
rect 4796 26360 4812 26424
rect 4876 26360 4892 26424
rect 4956 26360 4980 26424
rect 3348 22664 4980 26360
rect 30526 26134 30622 26150
rect 30526 26070 30542 26134
rect 30606 26070 30622 26134
rect 30526 26054 30622 26070
rect 30066 26023 30386 26042
rect 30066 26014 30388 26023
rect 29683 25786 29749 25787
rect 29683 25722 29684 25786
rect 29748 25784 29749 25786
rect 30066 25784 30075 26014
rect 29748 25724 30075 25784
rect 29748 25722 29749 25724
rect 29683 25721 29749 25722
rect 30066 25710 30075 25724
rect 30379 25710 30388 26014
rect 30066 25701 30388 25710
rect 30526 25990 30542 26054
rect 30606 25990 30622 26054
rect 31245 26134 31341 26150
rect 31245 26070 31261 26134
rect 31325 26070 31341 26134
rect 31245 26054 31341 26070
rect 30786 26023 31106 26042
rect 30526 25974 30622 25990
rect 30526 25910 30542 25974
rect 30606 25910 30622 25974
rect 30526 25894 30622 25910
rect 30526 25830 30542 25894
rect 30606 25830 30622 25894
rect 30526 25814 30622 25830
rect 30526 25750 30542 25814
rect 30606 25750 30622 25814
rect 30526 25734 30622 25750
rect 30066 25323 30386 25701
rect 30526 25670 30542 25734
rect 30606 25670 30622 25734
rect 30785 26014 31107 26023
rect 30785 25710 30794 26014
rect 31098 25710 31107 26014
rect 30785 25701 31107 25710
rect 31245 25990 31261 26054
rect 31325 25990 31341 26054
rect 31618 26042 31678 28402
rect 53456 26424 55088 30120
rect 33409 26396 33475 26397
rect 33409 26332 33410 26396
rect 33474 26332 33475 26396
rect 33409 26331 33475 26332
rect 53456 26360 53480 26424
rect 53544 26360 53560 26424
rect 53624 26360 53640 26424
rect 53704 26360 53720 26424
rect 53784 26360 53800 26424
rect 53864 26360 53880 26424
rect 53944 26360 53960 26424
rect 54024 26360 54040 26424
rect 54104 26360 54120 26424
rect 54184 26360 54200 26424
rect 54264 26360 54280 26424
rect 54344 26360 54360 26424
rect 54424 26360 54440 26424
rect 54504 26360 54520 26424
rect 54584 26360 54600 26424
rect 54664 26360 54680 26424
rect 54744 26360 54760 26424
rect 54824 26360 54840 26424
rect 54904 26360 54920 26424
rect 54984 26360 55000 26424
rect 55064 26360 55088 26424
rect 33412 26150 33472 26331
rect 31964 26134 32060 26150
rect 31964 26070 31980 26134
rect 32044 26070 32060 26134
rect 31964 26054 32060 26070
rect 31506 26023 31826 26042
rect 31245 25974 31341 25990
rect 31245 25910 31261 25974
rect 31325 25910 31341 25974
rect 31245 25894 31341 25910
rect 31245 25830 31261 25894
rect 31325 25830 31341 25894
rect 31245 25814 31341 25830
rect 31245 25750 31261 25814
rect 31325 25750 31341 25814
rect 31245 25734 31341 25750
rect 30526 25654 30622 25670
rect 30526 25590 30542 25654
rect 30606 25590 30622 25654
rect 30526 25574 30622 25590
rect 30526 25434 30622 25450
rect 30526 25370 30542 25434
rect 30606 25370 30622 25434
rect 30526 25354 30622 25370
rect 30066 25314 30388 25323
rect 30066 25010 30075 25314
rect 30379 25010 30388 25314
rect 30066 25001 30388 25010
rect 30526 25290 30542 25354
rect 30606 25290 30622 25354
rect 30786 25323 31106 25701
rect 31245 25670 31261 25734
rect 31325 25670 31341 25734
rect 31504 26014 31826 26023
rect 31504 25710 31513 26014
rect 31817 25710 31826 26014
rect 31504 25701 31826 25710
rect 31245 25654 31341 25670
rect 31245 25590 31261 25654
rect 31325 25590 31341 25654
rect 31245 25574 31341 25590
rect 31245 25434 31341 25450
rect 31245 25370 31261 25434
rect 31325 25370 31341 25434
rect 31245 25354 31341 25370
rect 30526 25274 30622 25290
rect 30526 25210 30542 25274
rect 30606 25210 30622 25274
rect 30526 25194 30622 25210
rect 30526 25130 30542 25194
rect 30606 25130 30622 25194
rect 30526 25114 30622 25130
rect 30526 25050 30542 25114
rect 30606 25050 30622 25114
rect 30526 25034 30622 25050
rect 30066 24762 30386 25001
rect 30526 24970 30542 25034
rect 30606 24970 30622 25034
rect 30785 25314 31107 25323
rect 30785 25010 30794 25314
rect 31098 25010 31107 25314
rect 30785 25001 31107 25010
rect 31245 25290 31261 25354
rect 31325 25290 31341 25354
rect 31506 25323 31826 25701
rect 31964 25990 31980 26054
rect 32044 25990 32060 26054
rect 32683 26134 32779 26150
rect 32683 26070 32699 26134
rect 32763 26070 32779 26134
rect 32683 26054 32779 26070
rect 32226 26023 32546 26042
rect 31964 25974 32060 25990
rect 31964 25910 31980 25974
rect 32044 25910 32060 25974
rect 31964 25894 32060 25910
rect 31964 25830 31980 25894
rect 32044 25830 32060 25894
rect 31964 25814 32060 25830
rect 31964 25750 31980 25814
rect 32044 25750 32060 25814
rect 31964 25734 32060 25750
rect 31964 25670 31980 25734
rect 32044 25670 32060 25734
rect 32223 26014 32546 26023
rect 32223 25710 32232 26014
rect 32536 25710 32546 26014
rect 32223 25701 32546 25710
rect 31964 25654 32060 25670
rect 31964 25590 31980 25654
rect 32044 25590 32060 25654
rect 31964 25574 32060 25590
rect 31245 25274 31341 25290
rect 31245 25210 31261 25274
rect 31325 25210 31341 25274
rect 31245 25194 31341 25210
rect 31245 25130 31261 25194
rect 31325 25130 31341 25194
rect 31245 25114 31341 25130
rect 31245 25050 31261 25114
rect 31325 25050 31341 25114
rect 31245 25034 31341 25050
rect 30526 24954 30622 24970
rect 30526 24890 30542 24954
rect 30606 24890 30622 24954
rect 30526 24874 30622 24890
rect 30786 24762 31106 25001
rect 31245 24970 31261 25034
rect 31325 24970 31341 25034
rect 31504 25314 31826 25323
rect 31504 25010 31513 25314
rect 31817 25010 31826 25314
rect 31504 25001 31826 25010
rect 31245 24954 31341 24970
rect 31245 24890 31261 24954
rect 31325 24890 31341 24954
rect 31245 24874 31341 24890
rect 31506 24762 31826 25001
rect 31964 25434 32060 25450
rect 31964 25370 31980 25434
rect 32044 25370 32060 25434
rect 31964 25354 32060 25370
rect 31964 25290 31980 25354
rect 32044 25290 32060 25354
rect 32226 25323 32546 25701
rect 32683 25990 32699 26054
rect 32763 25990 32779 26054
rect 33402 26134 33498 26150
rect 33402 26070 33418 26134
rect 33482 26070 33498 26134
rect 33402 26054 33498 26070
rect 32946 26023 33266 26042
rect 32683 25974 32779 25990
rect 32683 25910 32699 25974
rect 32763 25910 32779 25974
rect 32683 25894 32779 25910
rect 32683 25830 32699 25894
rect 32763 25830 32779 25894
rect 32683 25814 32779 25830
rect 32683 25750 32699 25814
rect 32763 25750 32779 25814
rect 32683 25734 32779 25750
rect 32683 25670 32699 25734
rect 32763 25670 32779 25734
rect 32942 26014 33266 26023
rect 32942 25710 32951 26014
rect 33255 25710 33266 26014
rect 32942 25701 33266 25710
rect 32683 25654 32779 25670
rect 32683 25590 32699 25654
rect 32763 25590 32779 25654
rect 32683 25574 32779 25590
rect 31964 25274 32060 25290
rect 31964 25210 31980 25274
rect 32044 25210 32060 25274
rect 31964 25194 32060 25210
rect 31964 25130 31980 25194
rect 32044 25130 32060 25194
rect 31964 25114 32060 25130
rect 31964 25050 31980 25114
rect 32044 25050 32060 25114
rect 31964 25034 32060 25050
rect 31964 24970 31980 25034
rect 32044 24970 32060 25034
rect 32223 25314 32546 25323
rect 32223 25010 32232 25314
rect 32536 25010 32546 25314
rect 32223 25001 32546 25010
rect 31964 24954 32060 24970
rect 31964 24890 31980 24954
rect 32044 24890 32060 24954
rect 31964 24874 32060 24890
rect 32226 24762 32546 25001
rect 32683 25434 32779 25450
rect 32683 25370 32699 25434
rect 32763 25370 32779 25434
rect 32683 25354 32779 25370
rect 32683 25290 32699 25354
rect 32763 25290 32779 25354
rect 32946 25323 33266 25701
rect 33402 25990 33418 26054
rect 33482 25990 33498 26054
rect 34121 26134 34217 26150
rect 34121 26070 34137 26134
rect 34201 26070 34217 26134
rect 34121 26054 34217 26070
rect 33666 26023 33986 26042
rect 33402 25974 33498 25990
rect 33402 25910 33418 25974
rect 33482 25910 33498 25974
rect 33402 25894 33498 25910
rect 33402 25830 33418 25894
rect 33482 25830 33498 25894
rect 33402 25814 33498 25830
rect 33402 25750 33418 25814
rect 33482 25750 33498 25814
rect 33402 25734 33498 25750
rect 33402 25670 33418 25734
rect 33482 25670 33498 25734
rect 33661 26014 33986 26023
rect 33661 25710 33670 26014
rect 33974 25710 33986 26014
rect 33661 25701 33986 25710
rect 33402 25654 33498 25670
rect 33402 25590 33418 25654
rect 33482 25590 33498 25654
rect 33402 25574 33498 25590
rect 32683 25274 32779 25290
rect 32683 25210 32699 25274
rect 32763 25210 32779 25274
rect 32683 25194 32779 25210
rect 32683 25130 32699 25194
rect 32763 25130 32779 25194
rect 32683 25114 32779 25130
rect 32683 25050 32699 25114
rect 32763 25050 32779 25114
rect 32683 25034 32779 25050
rect 32683 24970 32699 25034
rect 32763 24970 32779 25034
rect 32942 25314 33266 25323
rect 32942 25010 32951 25314
rect 33255 25010 33266 25314
rect 32942 25001 33266 25010
rect 32683 24954 32779 24970
rect 32683 24890 32699 24954
rect 32763 24890 32779 24954
rect 32683 24874 32779 24890
rect 32946 24762 33266 25001
rect 33402 25434 33498 25450
rect 33402 25370 33418 25434
rect 33482 25370 33498 25434
rect 33402 25354 33498 25370
rect 33402 25290 33418 25354
rect 33482 25290 33498 25354
rect 33666 25323 33986 25701
rect 34121 25990 34137 26054
rect 34201 25990 34217 26054
rect 34840 26134 34936 26150
rect 34840 26070 34856 26134
rect 34920 26070 34936 26134
rect 34840 26054 34936 26070
rect 34386 26023 34706 26042
rect 34121 25974 34217 25990
rect 34121 25910 34137 25974
rect 34201 25910 34217 25974
rect 34121 25894 34217 25910
rect 34121 25830 34137 25894
rect 34201 25830 34217 25894
rect 34121 25814 34217 25830
rect 34121 25750 34137 25814
rect 34201 25750 34217 25814
rect 34121 25734 34217 25750
rect 34121 25670 34137 25734
rect 34201 25670 34217 25734
rect 34380 26014 34706 26023
rect 34380 25710 34389 26014
rect 34693 25710 34706 26014
rect 34380 25701 34706 25710
rect 34121 25654 34217 25670
rect 34121 25590 34137 25654
rect 34201 25590 34217 25654
rect 34121 25574 34217 25590
rect 33402 25274 33498 25290
rect 33402 25210 33418 25274
rect 33482 25210 33498 25274
rect 33402 25194 33498 25210
rect 33402 25130 33418 25194
rect 33482 25130 33498 25194
rect 33402 25114 33498 25130
rect 33402 25050 33418 25114
rect 33482 25050 33498 25114
rect 33402 25034 33498 25050
rect 33402 24970 33418 25034
rect 33482 24970 33498 25034
rect 33661 25314 33986 25323
rect 33661 25010 33670 25314
rect 33974 25010 33986 25314
rect 33661 25001 33986 25010
rect 33402 24954 33498 24970
rect 33402 24890 33418 24954
rect 33482 24890 33498 24954
rect 33402 24874 33498 24890
rect 33666 24762 33986 25001
rect 34121 25434 34217 25450
rect 34121 25370 34137 25434
rect 34201 25370 34217 25434
rect 34121 25354 34217 25370
rect 34121 25290 34137 25354
rect 34201 25290 34217 25354
rect 34386 25323 34706 25701
rect 34840 25990 34856 26054
rect 34920 25990 34936 26054
rect 35559 26134 35655 26150
rect 35559 26070 35575 26134
rect 35639 26070 35655 26134
rect 35559 26054 35655 26070
rect 35106 26023 35426 26042
rect 34840 25974 34936 25990
rect 34840 25910 34856 25974
rect 34920 25910 34936 25974
rect 34840 25894 34936 25910
rect 34840 25830 34856 25894
rect 34920 25830 34936 25894
rect 34840 25814 34936 25830
rect 34840 25750 34856 25814
rect 34920 25750 34936 25814
rect 34840 25734 34936 25750
rect 34840 25670 34856 25734
rect 34920 25670 34936 25734
rect 35099 26014 35426 26023
rect 35099 25710 35108 26014
rect 35412 25710 35426 26014
rect 35099 25701 35426 25710
rect 34840 25654 34936 25670
rect 34840 25590 34856 25654
rect 34920 25590 34936 25654
rect 34840 25574 34936 25590
rect 34121 25274 34217 25290
rect 34121 25210 34137 25274
rect 34201 25210 34217 25274
rect 34121 25194 34217 25210
rect 34121 25130 34137 25194
rect 34201 25130 34217 25194
rect 34121 25114 34217 25130
rect 34121 25050 34137 25114
rect 34201 25050 34217 25114
rect 34121 25034 34217 25050
rect 34121 24970 34137 25034
rect 34201 24970 34217 25034
rect 34380 25314 34706 25323
rect 34380 25010 34389 25314
rect 34693 25010 34706 25314
rect 34380 25001 34706 25010
rect 34121 24954 34217 24970
rect 34121 24890 34137 24954
rect 34201 24890 34217 24954
rect 34121 24874 34217 24890
rect 34386 24762 34706 25001
rect 34840 25434 34936 25450
rect 34840 25370 34856 25434
rect 34920 25370 34936 25434
rect 34840 25354 34936 25370
rect 34840 25290 34856 25354
rect 34920 25290 34936 25354
rect 35106 25323 35426 25701
rect 35559 25990 35575 26054
rect 35639 25990 35655 26054
rect 36278 26134 36374 26150
rect 36278 26070 36294 26134
rect 36358 26070 36374 26134
rect 36278 26054 36374 26070
rect 35826 26023 36146 26042
rect 35559 25974 35655 25990
rect 35559 25910 35575 25974
rect 35639 25910 35655 25974
rect 35559 25894 35655 25910
rect 35559 25830 35575 25894
rect 35639 25830 35655 25894
rect 35559 25814 35655 25830
rect 35559 25750 35575 25814
rect 35639 25750 35655 25814
rect 35559 25734 35655 25750
rect 35559 25670 35575 25734
rect 35639 25670 35655 25734
rect 35818 26014 36146 26023
rect 35818 25710 35827 26014
rect 36131 25710 36146 26014
rect 35818 25701 36146 25710
rect 35559 25654 35655 25670
rect 35559 25590 35575 25654
rect 35639 25590 35655 25654
rect 35559 25574 35655 25590
rect 34840 25274 34936 25290
rect 34840 25210 34856 25274
rect 34920 25210 34936 25274
rect 34840 25194 34936 25210
rect 34840 25130 34856 25194
rect 34920 25130 34936 25194
rect 34840 25114 34936 25130
rect 34840 25050 34856 25114
rect 34920 25050 34936 25114
rect 34840 25034 34936 25050
rect 34840 24970 34856 25034
rect 34920 24970 34936 25034
rect 35099 25314 35426 25323
rect 35099 25010 35108 25314
rect 35412 25010 35426 25314
rect 35099 25001 35426 25010
rect 34840 24954 34936 24970
rect 34840 24890 34856 24954
rect 34920 24890 34936 24954
rect 34840 24874 34936 24890
rect 35106 24762 35426 25001
rect 35559 25434 35655 25450
rect 35559 25370 35575 25434
rect 35639 25370 35655 25434
rect 35559 25354 35655 25370
rect 35559 25290 35575 25354
rect 35639 25290 35655 25354
rect 35826 25323 36146 25701
rect 36278 25990 36294 26054
rect 36358 25990 36374 26054
rect 36997 26134 37093 26150
rect 36997 26070 37013 26134
rect 37077 26070 37093 26134
rect 36997 26054 37093 26070
rect 36546 26023 36866 26042
rect 36278 25974 36374 25990
rect 36278 25910 36294 25974
rect 36358 25910 36374 25974
rect 36278 25894 36374 25910
rect 36278 25830 36294 25894
rect 36358 25830 36374 25894
rect 36278 25814 36374 25830
rect 36278 25750 36294 25814
rect 36358 25750 36374 25814
rect 36278 25734 36374 25750
rect 36278 25670 36294 25734
rect 36358 25670 36374 25734
rect 36537 26014 36866 26023
rect 36537 25710 36546 26014
rect 36850 25710 36866 26014
rect 36537 25701 36866 25710
rect 36278 25654 36374 25670
rect 36278 25590 36294 25654
rect 36358 25590 36374 25654
rect 36278 25574 36374 25590
rect 35559 25274 35655 25290
rect 35559 25210 35575 25274
rect 35639 25210 35655 25274
rect 35559 25194 35655 25210
rect 35559 25130 35575 25194
rect 35639 25130 35655 25194
rect 35559 25114 35655 25130
rect 35559 25050 35575 25114
rect 35639 25050 35655 25114
rect 35559 25034 35655 25050
rect 35559 24970 35575 25034
rect 35639 24970 35655 25034
rect 35818 25314 36146 25323
rect 35818 25010 35827 25314
rect 36131 25010 36146 25314
rect 35818 25001 36146 25010
rect 35559 24954 35655 24970
rect 35559 24890 35575 24954
rect 35639 24890 35655 24954
rect 35559 24874 35655 24890
rect 35826 24762 36146 25001
rect 36278 25434 36374 25450
rect 36278 25370 36294 25434
rect 36358 25370 36374 25434
rect 36278 25354 36374 25370
rect 36278 25290 36294 25354
rect 36358 25290 36374 25354
rect 36546 25323 36866 25701
rect 36997 25990 37013 26054
rect 37077 25990 37093 26054
rect 36997 25974 37093 25990
rect 36997 25910 37013 25974
rect 37077 25910 37093 25974
rect 36997 25894 37093 25910
rect 36997 25830 37013 25894
rect 37077 25830 37093 25894
rect 36997 25814 37093 25830
rect 36997 25750 37013 25814
rect 37077 25750 37093 25814
rect 36997 25734 37093 25750
rect 36997 25670 37013 25734
rect 37077 25670 37093 25734
rect 36997 25654 37093 25670
rect 36997 25590 37013 25654
rect 37077 25590 37093 25654
rect 36997 25574 37093 25590
rect 36278 25274 36374 25290
rect 36278 25210 36294 25274
rect 36358 25210 36374 25274
rect 36278 25194 36374 25210
rect 36278 25130 36294 25194
rect 36358 25130 36374 25194
rect 36278 25114 36374 25130
rect 36278 25050 36294 25114
rect 36358 25050 36374 25114
rect 36278 25034 36374 25050
rect 36278 24970 36294 25034
rect 36358 24970 36374 25034
rect 36537 25314 36866 25323
rect 36537 25010 36546 25314
rect 36850 25010 36866 25314
rect 36537 25001 36866 25010
rect 36278 24954 36374 24970
rect 36278 24890 36294 24954
rect 36358 24890 36374 24954
rect 36278 24874 36374 24890
rect 36546 24762 36866 25001
rect 36997 25434 37093 25450
rect 36997 25370 37013 25434
rect 37077 25370 37093 25434
rect 36997 25354 37093 25370
rect 36997 25290 37013 25354
rect 37077 25290 37093 25354
rect 36997 25274 37093 25290
rect 36997 25210 37013 25274
rect 37077 25210 37093 25274
rect 36997 25194 37093 25210
rect 36997 25130 37013 25194
rect 37077 25130 37093 25194
rect 36997 25114 37093 25130
rect 36997 25050 37013 25114
rect 37077 25050 37093 25114
rect 36997 25034 37093 25050
rect 36997 24970 37013 25034
rect 37077 24970 37093 25034
rect 36997 24954 37093 24970
rect 36997 24890 37013 24954
rect 37077 24890 37093 24954
rect 36997 24874 37093 24890
rect 29928 24734 37096 24762
rect 29928 24670 29956 24734
rect 30020 24670 30036 24734
rect 30100 24670 37096 24734
rect 29928 24642 37096 24670
rect 3348 22600 3372 22664
rect 3436 22600 3452 22664
rect 3516 22600 3532 22664
rect 3596 22600 3612 22664
rect 3676 22600 3692 22664
rect 3756 22600 3772 22664
rect 3836 22600 3852 22664
rect 3916 22600 3932 22664
rect 3996 22600 4012 22664
rect 4076 22600 4092 22664
rect 4156 22600 4172 22664
rect 4236 22600 4252 22664
rect 4316 22600 4332 22664
rect 4396 22600 4412 22664
rect 4476 22600 4492 22664
rect 4556 22600 4572 22664
rect 4636 22600 4652 22664
rect 4716 22600 4732 22664
rect 4796 22600 4812 22664
rect 4876 22600 4892 22664
rect 4956 22600 4980 22664
rect 3348 18904 4980 22600
rect 3348 18840 3372 18904
rect 3436 18840 3452 18904
rect 3516 18840 3532 18904
rect 3596 18840 3612 18904
rect 3676 18840 3692 18904
rect 3756 18840 3772 18904
rect 3836 18840 3852 18904
rect 3916 18840 3932 18904
rect 3996 18840 4012 18904
rect 4076 18840 4092 18904
rect 4156 18840 4172 18904
rect 4236 18840 4252 18904
rect 4316 18840 4332 18904
rect 4396 18840 4412 18904
rect 4476 18840 4492 18904
rect 4556 18840 4572 18904
rect 4636 18840 4652 18904
rect 4716 18840 4732 18904
rect 4796 18840 4812 18904
rect 4876 18840 4892 18904
rect 4956 18840 4980 18904
rect 3348 15144 4980 18840
rect 3348 15080 3372 15144
rect 3436 15080 3452 15144
rect 3516 15080 3532 15144
rect 3596 15080 3612 15144
rect 3676 15080 3692 15144
rect 3756 15080 3772 15144
rect 3836 15080 3852 15144
rect 3916 15080 3932 15144
rect 3996 15080 4012 15144
rect 4076 15080 4092 15144
rect 4156 15080 4172 15144
rect 4236 15080 4252 15144
rect 4316 15080 4332 15144
rect 4396 15080 4412 15144
rect 4476 15080 4492 15144
rect 4556 15080 4572 15144
rect 4636 15080 4652 15144
rect 4716 15080 4732 15144
rect 4796 15080 4812 15144
rect 4876 15080 4892 15144
rect 4956 15080 4980 15144
rect 3348 11384 4980 15080
rect 3348 11320 3372 11384
rect 3436 11320 3452 11384
rect 3516 11320 3532 11384
rect 3596 11320 3612 11384
rect 3676 11320 3692 11384
rect 3756 11320 3772 11384
rect 3836 11320 3852 11384
rect 3916 11320 3932 11384
rect 3996 11320 4012 11384
rect 4076 11320 4092 11384
rect 4156 11320 4172 11384
rect 4236 11320 4252 11384
rect 4316 11320 4332 11384
rect 4396 11320 4412 11384
rect 4476 11320 4492 11384
rect 4556 11320 4572 11384
rect 4636 11320 4652 11384
rect 4716 11320 4732 11384
rect 4796 11320 4812 11384
rect 4876 11320 4892 11384
rect 4956 11320 4980 11384
rect 3348 7624 4980 11320
rect 3348 7560 3372 7624
rect 3436 7560 3452 7624
rect 3516 7560 3532 7624
rect 3596 7560 3612 7624
rect 3676 7560 3692 7624
rect 3756 7560 3772 7624
rect 3836 7560 3852 7624
rect 3916 7560 3932 7624
rect 3996 7560 4012 7624
rect 4076 7560 4092 7624
rect 4156 7560 4172 7624
rect 4236 7560 4252 7624
rect 4316 7560 4332 7624
rect 4396 7560 4412 7624
rect 4476 7560 4492 7624
rect 4556 7560 4572 7624
rect 4636 7560 4652 7624
rect 4716 7560 4732 7624
rect 4796 7560 4812 7624
rect 4876 7560 4892 7624
rect 4956 7560 4980 7624
rect 3348 4838 4980 7560
rect 3348 3322 3406 4838
rect 4922 3322 4980 4838
rect 3348 0 4980 3322
rect 53456 22664 55088 26360
rect 53456 22600 53480 22664
rect 53544 22600 53560 22664
rect 53624 22600 53640 22664
rect 53704 22600 53720 22664
rect 53784 22600 53800 22664
rect 53864 22600 53880 22664
rect 53944 22600 53960 22664
rect 54024 22600 54040 22664
rect 54104 22600 54120 22664
rect 54184 22600 54200 22664
rect 54264 22600 54280 22664
rect 54344 22600 54360 22664
rect 54424 22600 54440 22664
rect 54504 22600 54520 22664
rect 54584 22600 54600 22664
rect 54664 22600 54680 22664
rect 54744 22600 54760 22664
rect 54824 22600 54840 22664
rect 54904 22600 54920 22664
rect 54984 22600 55000 22664
rect 55064 22600 55088 22664
rect 53456 18904 55088 22600
rect 53456 18840 53480 18904
rect 53544 18840 53560 18904
rect 53624 18840 53640 18904
rect 53704 18840 53720 18904
rect 53784 18840 53800 18904
rect 53864 18840 53880 18904
rect 53944 18840 53960 18904
rect 54024 18840 54040 18904
rect 54104 18840 54120 18904
rect 54184 18840 54200 18904
rect 54264 18840 54280 18904
rect 54344 18840 54360 18904
rect 54424 18840 54440 18904
rect 54504 18840 54520 18904
rect 54584 18840 54600 18904
rect 54664 18840 54680 18904
rect 54744 18840 54760 18904
rect 54824 18840 54840 18904
rect 54904 18840 54920 18904
rect 54984 18840 55000 18904
rect 55064 18840 55088 18904
rect 53456 15144 55088 18840
rect 53456 15080 53480 15144
rect 53544 15080 53560 15144
rect 53624 15080 53640 15144
rect 53704 15080 53720 15144
rect 53784 15080 53800 15144
rect 53864 15080 53880 15144
rect 53944 15080 53960 15144
rect 54024 15080 54040 15144
rect 54104 15080 54120 15144
rect 54184 15080 54200 15144
rect 54264 15080 54280 15144
rect 54344 15080 54360 15144
rect 54424 15080 54440 15144
rect 54504 15080 54520 15144
rect 54584 15080 54600 15144
rect 54664 15080 54680 15144
rect 54744 15080 54760 15144
rect 54824 15080 54840 15144
rect 54904 15080 54920 15144
rect 54984 15080 55000 15144
rect 55064 15080 55088 15144
rect 53456 11384 55088 15080
rect 53456 11320 53480 11384
rect 53544 11320 53560 11384
rect 53624 11320 53640 11384
rect 53704 11320 53720 11384
rect 53784 11320 53800 11384
rect 53864 11320 53880 11384
rect 53944 11320 53960 11384
rect 54024 11320 54040 11384
rect 54104 11320 54120 11384
rect 54184 11320 54200 11384
rect 54264 11320 54280 11384
rect 54344 11320 54360 11384
rect 54424 11320 54440 11384
rect 54504 11320 54520 11384
rect 54584 11320 54600 11384
rect 54664 11320 54680 11384
rect 54744 11320 54760 11384
rect 54824 11320 54840 11384
rect 54904 11320 54920 11384
rect 54984 11320 55000 11384
rect 55064 11320 55088 11384
rect 53456 7624 55088 11320
rect 53456 7560 53480 7624
rect 53544 7560 53560 7624
rect 53624 7560 53640 7624
rect 53704 7560 53720 7624
rect 53784 7560 53800 7624
rect 53864 7560 53880 7624
rect 53944 7560 53960 7624
rect 54024 7560 54040 7624
rect 54104 7560 54120 7624
rect 54184 7560 54200 7624
rect 54264 7560 54280 7624
rect 54344 7560 54360 7624
rect 54424 7560 54440 7624
rect 54504 7560 54520 7624
rect 54584 7560 54600 7624
rect 54664 7560 54680 7624
rect 54744 7560 54760 7624
rect 54824 7560 54840 7624
rect 54904 7560 54920 7624
rect 54984 7560 55000 7624
rect 55064 7560 55088 7624
rect 53456 4838 55088 7560
rect 53456 3322 53514 4838
rect 55030 3322 55088 4838
rect 53456 0 55088 3322
rect 55904 55670 57536 56576
rect 55904 54154 55962 55670
rect 57478 54154 57536 55670
rect 55904 50864 57536 54154
rect 55904 50800 55928 50864
rect 55992 50800 56008 50864
rect 56072 50800 56088 50864
rect 56152 50800 56168 50864
rect 56232 50800 56248 50864
rect 56312 50800 56328 50864
rect 56392 50800 56408 50864
rect 56472 50800 56488 50864
rect 56552 50800 56568 50864
rect 56632 50800 56648 50864
rect 56712 50800 56728 50864
rect 56792 50800 56808 50864
rect 56872 50800 56888 50864
rect 56952 50800 56968 50864
rect 57032 50800 57048 50864
rect 57112 50800 57128 50864
rect 57192 50800 57208 50864
rect 57272 50800 57288 50864
rect 57352 50800 57368 50864
rect 57432 50800 57448 50864
rect 57512 50800 57536 50864
rect 55904 47104 57536 50800
rect 55904 47040 55928 47104
rect 55992 47040 56008 47104
rect 56072 47040 56088 47104
rect 56152 47040 56168 47104
rect 56232 47040 56248 47104
rect 56312 47040 56328 47104
rect 56392 47040 56408 47104
rect 56472 47040 56488 47104
rect 56552 47040 56568 47104
rect 56632 47040 56648 47104
rect 56712 47040 56728 47104
rect 56792 47040 56808 47104
rect 56872 47040 56888 47104
rect 56952 47040 56968 47104
rect 57032 47040 57048 47104
rect 57112 47040 57128 47104
rect 57192 47040 57208 47104
rect 57272 47040 57288 47104
rect 57352 47040 57368 47104
rect 57432 47040 57448 47104
rect 57512 47040 57536 47104
rect 55904 43344 57536 47040
rect 55904 43280 55928 43344
rect 55992 43280 56008 43344
rect 56072 43280 56088 43344
rect 56152 43280 56168 43344
rect 56232 43280 56248 43344
rect 56312 43280 56328 43344
rect 56392 43280 56408 43344
rect 56472 43280 56488 43344
rect 56552 43280 56568 43344
rect 56632 43280 56648 43344
rect 56712 43280 56728 43344
rect 56792 43280 56808 43344
rect 56872 43280 56888 43344
rect 56952 43280 56968 43344
rect 57032 43280 57048 43344
rect 57112 43280 57128 43344
rect 57192 43280 57208 43344
rect 57272 43280 57288 43344
rect 57352 43280 57368 43344
rect 57432 43280 57448 43344
rect 57512 43280 57536 43344
rect 55904 39584 57536 43280
rect 55904 39520 55928 39584
rect 55992 39520 56008 39584
rect 56072 39520 56088 39584
rect 56152 39520 56168 39584
rect 56232 39520 56248 39584
rect 56312 39520 56328 39584
rect 56392 39520 56408 39584
rect 56472 39520 56488 39584
rect 56552 39520 56568 39584
rect 56632 39520 56648 39584
rect 56712 39520 56728 39584
rect 56792 39520 56808 39584
rect 56872 39520 56888 39584
rect 56952 39520 56968 39584
rect 57032 39520 57048 39584
rect 57112 39520 57128 39584
rect 57192 39520 57208 39584
rect 57272 39520 57288 39584
rect 57352 39520 57368 39584
rect 57432 39520 57448 39584
rect 57512 39520 57536 39584
rect 55904 35824 57536 39520
rect 55904 35760 55928 35824
rect 55992 35760 56008 35824
rect 56072 35760 56088 35824
rect 56152 35760 56168 35824
rect 56232 35760 56248 35824
rect 56312 35760 56328 35824
rect 56392 35760 56408 35824
rect 56472 35760 56488 35824
rect 56552 35760 56568 35824
rect 56632 35760 56648 35824
rect 56712 35760 56728 35824
rect 56792 35760 56808 35824
rect 56872 35760 56888 35824
rect 56952 35760 56968 35824
rect 57032 35760 57048 35824
rect 57112 35760 57128 35824
rect 57192 35760 57208 35824
rect 57272 35760 57288 35824
rect 57352 35760 57368 35824
rect 57432 35760 57448 35824
rect 57512 35760 57536 35824
rect 55904 32064 57536 35760
rect 55904 32000 55928 32064
rect 55992 32000 56008 32064
rect 56072 32000 56088 32064
rect 56152 32000 56168 32064
rect 56232 32000 56248 32064
rect 56312 32000 56328 32064
rect 56392 32000 56408 32064
rect 56472 32000 56488 32064
rect 56552 32000 56568 32064
rect 56632 32000 56648 32064
rect 56712 32000 56728 32064
rect 56792 32000 56808 32064
rect 56872 32000 56888 32064
rect 56952 32000 56968 32064
rect 57032 32000 57048 32064
rect 57112 32000 57128 32064
rect 57192 32000 57208 32064
rect 57272 32000 57288 32064
rect 57352 32000 57368 32064
rect 57432 32000 57448 32064
rect 57512 32000 57536 32064
rect 55904 28304 57536 32000
rect 55904 28240 55928 28304
rect 55992 28240 56008 28304
rect 56072 28240 56088 28304
rect 56152 28240 56168 28304
rect 56232 28240 56248 28304
rect 56312 28240 56328 28304
rect 56392 28240 56408 28304
rect 56472 28240 56488 28304
rect 56552 28240 56568 28304
rect 56632 28240 56648 28304
rect 56712 28240 56728 28304
rect 56792 28240 56808 28304
rect 56872 28240 56888 28304
rect 56952 28240 56968 28304
rect 57032 28240 57048 28304
rect 57112 28240 57128 28304
rect 57192 28240 57208 28304
rect 57272 28240 57288 28304
rect 57352 28240 57368 28304
rect 57432 28240 57448 28304
rect 57512 28240 57536 28304
rect 55904 24544 57536 28240
rect 55904 24480 55928 24544
rect 55992 24480 56008 24544
rect 56072 24480 56088 24544
rect 56152 24480 56168 24544
rect 56232 24480 56248 24544
rect 56312 24480 56328 24544
rect 56392 24480 56408 24544
rect 56472 24480 56488 24544
rect 56552 24480 56568 24544
rect 56632 24480 56648 24544
rect 56712 24480 56728 24544
rect 56792 24480 56808 24544
rect 56872 24480 56888 24544
rect 56952 24480 56968 24544
rect 57032 24480 57048 24544
rect 57112 24480 57128 24544
rect 57192 24480 57208 24544
rect 57272 24480 57288 24544
rect 57352 24480 57368 24544
rect 57432 24480 57448 24544
rect 57512 24480 57536 24544
rect 55904 20784 57536 24480
rect 55904 20720 55928 20784
rect 55992 20720 56008 20784
rect 56072 20720 56088 20784
rect 56152 20720 56168 20784
rect 56232 20720 56248 20784
rect 56312 20720 56328 20784
rect 56392 20720 56408 20784
rect 56472 20720 56488 20784
rect 56552 20720 56568 20784
rect 56632 20720 56648 20784
rect 56712 20720 56728 20784
rect 56792 20720 56808 20784
rect 56872 20720 56888 20784
rect 56952 20720 56968 20784
rect 57032 20720 57048 20784
rect 57112 20720 57128 20784
rect 57192 20720 57208 20784
rect 57272 20720 57288 20784
rect 57352 20720 57368 20784
rect 57432 20720 57448 20784
rect 57512 20720 57536 20784
rect 55904 17024 57536 20720
rect 55904 16960 55928 17024
rect 55992 16960 56008 17024
rect 56072 16960 56088 17024
rect 56152 16960 56168 17024
rect 56232 16960 56248 17024
rect 56312 16960 56328 17024
rect 56392 16960 56408 17024
rect 56472 16960 56488 17024
rect 56552 16960 56568 17024
rect 56632 16960 56648 17024
rect 56712 16960 56728 17024
rect 56792 16960 56808 17024
rect 56872 16960 56888 17024
rect 56952 16960 56968 17024
rect 57032 16960 57048 17024
rect 57112 16960 57128 17024
rect 57192 16960 57208 17024
rect 57272 16960 57288 17024
rect 57352 16960 57368 17024
rect 57432 16960 57448 17024
rect 57512 16960 57536 17024
rect 55904 13264 57536 16960
rect 55904 13200 55928 13264
rect 55992 13200 56008 13264
rect 56072 13200 56088 13264
rect 56152 13200 56168 13264
rect 56232 13200 56248 13264
rect 56312 13200 56328 13264
rect 56392 13200 56408 13264
rect 56472 13200 56488 13264
rect 56552 13200 56568 13264
rect 56632 13200 56648 13264
rect 56712 13200 56728 13264
rect 56792 13200 56808 13264
rect 56872 13200 56888 13264
rect 56952 13200 56968 13264
rect 57032 13200 57048 13264
rect 57112 13200 57128 13264
rect 57192 13200 57208 13264
rect 57272 13200 57288 13264
rect 57352 13200 57368 13264
rect 57432 13200 57448 13264
rect 57512 13200 57536 13264
rect 55904 9504 57536 13200
rect 55904 9440 55928 9504
rect 55992 9440 56008 9504
rect 56072 9440 56088 9504
rect 56152 9440 56168 9504
rect 56232 9440 56248 9504
rect 56312 9440 56328 9504
rect 56392 9440 56408 9504
rect 56472 9440 56488 9504
rect 56552 9440 56568 9504
rect 56632 9440 56648 9504
rect 56712 9440 56728 9504
rect 56792 9440 56808 9504
rect 56872 9440 56888 9504
rect 56952 9440 56968 9504
rect 57032 9440 57048 9504
rect 57112 9440 57128 9504
rect 57192 9440 57208 9504
rect 57272 9440 57288 9504
rect 57352 9440 57368 9504
rect 57432 9440 57448 9504
rect 57512 9440 57536 9504
rect 55904 5744 57536 9440
rect 55904 5680 55928 5744
rect 55992 5680 56008 5744
rect 56072 5680 56088 5744
rect 56152 5680 56168 5744
rect 56232 5680 56248 5744
rect 56312 5680 56328 5744
rect 56392 5680 56408 5744
rect 56472 5680 56488 5744
rect 56552 5680 56568 5744
rect 56632 5680 56648 5744
rect 56712 5680 56728 5744
rect 56792 5680 56808 5744
rect 56872 5680 56888 5744
rect 56952 5680 56968 5744
rect 57032 5680 57048 5744
rect 57112 5680 57128 5744
rect 57192 5680 57208 5744
rect 57272 5680 57288 5744
rect 57352 5680 57368 5744
rect 57432 5680 57448 5744
rect 57512 5680 57536 5744
rect 55904 2390 57536 5680
rect 55904 874 55962 2390
rect 57478 874 57536 2390
rect 55904 0 57536 874
<< via4 >>
rect 958 54154 2474 55670
rect 958 874 2474 2390
rect 3406 51706 4922 53222
rect 53514 51706 55030 53222
rect 3406 3322 4922 4838
rect 53514 3322 55030 4838
rect 55962 54154 57478 55670
rect 55962 874 57478 2390
<< metal5 >>
rect 0 55670 58512 55728
rect 0 54154 958 55670
rect 2474 54154 55962 55670
rect 57478 54154 58512 55670
rect 0 54096 58512 54154
rect 0 53222 58512 53280
rect 0 51706 3406 53222
rect 4922 51706 53514 53222
rect 55030 51706 58512 53222
rect 0 51648 58512 51706
rect 0 4838 58512 4896
rect 0 3322 3406 4838
rect 4922 3322 53514 4838
rect 55030 3322 58512 4838
rect 0 3264 58512 3322
rect 0 2390 58512 2448
rect 0 874 958 2390
rect 2474 874 55962 2390
rect 57478 874 58512 2390
rect 0 816 58512 874
<< labels >>
rlabel metal2 s 25516 0 25544 97 4 porst
port 1 nsew
rlabel metal3 s 0 40974 160 41034 4 va
port 2 nsew
rlabel metal1 s 58393 33408 58512 33436 4 vb
port 3 nsew
rlabel metal2 s 34348 0 34376 97 4 vbg
port 4 nsew
rlabel metal5 s 0 816 1632 2448 4 VSS
port 5 nsew
rlabel metal5 s 0 3264 1632 4896 4 VDD
port 6 nsew
flabel metal1 50156 7012 50276 7132 1 FreeSans 600 0 0 0 sky130_asc_res_xhigh_po_2p85_1_7/Rin
flabel metal1 50156 6052 50276 6172 1 FreeSans 600 0 0 0 sky130_asc_res_xhigh_po_2p85_1_7/Rout
flabel metal1 50036 7562 50096 7622 1 FreeSans 1000 0 0 0 sky130_asc_res_xhigh_po_2p85_1_7/VPWR
flabel metal1 50036 5682 50096 5742 1 FreeSans 1000 0 0 0 sky130_asc_res_xhigh_po_2p85_1_7/VGND
flabel metal1 44668 7012 44788 7132 1 FreeSans 600 0 0 0 sky130_asc_res_xhigh_po_2p85_1_6/Rin
flabel metal1 44668 6052 44788 6172 1 FreeSans 600 0 0 0 sky130_asc_res_xhigh_po_2p85_1_6/Rout
flabel metal1 44548 7562 44608 7622 1 FreeSans 1000 0 0 0 sky130_asc_res_xhigh_po_2p85_1_6/VPWR
flabel metal1 44548 5682 44608 5742 1 FreeSans 1000 0 0 0 sky130_asc_res_xhigh_po_2p85_1_6/VGND
flabel metal1 47412 7012 47532 7132 1 FreeSans 600 0 0 0 sky130_asc_res_xhigh_po_2p85_1_0/Rin
flabel metal1 47412 6052 47532 6172 1 FreeSans 600 0 0 0 sky130_asc_res_xhigh_po_2p85_1_0/Rout
flabel metal1 47292 7562 47352 7622 1 FreeSans 1000 0 0 0 sky130_asc_res_xhigh_po_2p85_1_0/VPWR
flabel metal1 47292 5682 47352 5742 1 FreeSans 1000 0 0 0 sky130_asc_res_xhigh_po_2p85_1_0/VGND
flabel metal1 43884 10772 44004 10892 1 FreeSans 600 0 0 0 sky130_asc_res_xhigh_po_2p85_1_8/Rin
flabel metal1 43884 9812 44004 9932 1 FreeSans 600 0 0 0 sky130_asc_res_xhigh_po_2p85_1_8/Rout
flabel metal1 43764 11322 43824 11382 1 FreeSans 1000 0 0 0 sky130_asc_res_xhigh_po_2p85_1_8/VPWR
flabel metal1 43764 9442 43824 9502 1 FreeSans 1000 0 0 0 sky130_asc_res_xhigh_po_2p85_1_8/VGND
flabel metal1 46628 10772 46748 10892 1 FreeSans 600 0 0 0 sky130_asc_res_xhigh_po_2p85_1_5/Rin
flabel metal1 46628 9812 46748 9932 1 FreeSans 600 0 0 0 sky130_asc_res_xhigh_po_2p85_1_5/Rout
flabel metal1 46508 11322 46568 11382 1 FreeSans 1000 0 0 0 sky130_asc_res_xhigh_po_2p85_1_5/VPWR
flabel metal1 46508 9442 46568 9502 1 FreeSans 1000 0 0 0 sky130_asc_res_xhigh_po_2p85_1_5/VGND
flabel metal1 49372 10772 49492 10892 1 FreeSans 600 0 0 0 sky130_asc_res_xhigh_po_2p85_1_3/Rin
flabel metal1 49372 9812 49492 9932 1 FreeSans 600 0 0 0 sky130_asc_res_xhigh_po_2p85_1_3/Rout
flabel metal1 49252 11322 49312 11382 1 FreeSans 1000 0 0 0 sky130_asc_res_xhigh_po_2p85_1_3/VPWR
flabel metal1 49252 9442 49312 9502 1 FreeSans 1000 0 0 0 sky130_asc_res_xhigh_po_2p85_1_3/VGND
flabel metal1 43982 14532 44102 14652 1 FreeSans 600 0 0 0 sky130_asc_res_xhigh_po_2p85_1_2/Rin
flabel metal1 43982 13572 44102 13692 1 FreeSans 600 0 0 0 sky130_asc_res_xhigh_po_2p85_1_2/Rout
flabel metal1 43862 15082 43922 15142 1 FreeSans 1000 0 0 0 sky130_asc_res_xhigh_po_2p85_1_2/VPWR
flabel metal1 43862 13202 43922 13262 1 FreeSans 1000 0 0 0 sky130_asc_res_xhigh_po_2p85_1_2/VGND
flabel metal1 46726 14532 46846 14652 1 FreeSans 600 0 0 0 sky130_asc_res_xhigh_po_2p85_1_4/Rin
flabel metal1 46726 13572 46846 13692 1 FreeSans 600 0 0 0 sky130_asc_res_xhigh_po_2p85_1_4/Rout
flabel metal1 46606 15082 46666 15142 1 FreeSans 1000 0 0 0 sky130_asc_res_xhigh_po_2p85_1_4/VPWR
flabel metal1 46606 13202 46666 13262 1 FreeSans 1000 0 0 0 sky130_asc_res_xhigh_po_2p85_1_4/VGND
flabel metal1 49470 14532 49590 14652 1 FreeSans 600 0 0 0 sky130_asc_res_xhigh_po_2p85_1_1/Rin
flabel metal1 49470 13572 49590 13692 1 FreeSans 600 0 0 0 sky130_asc_res_xhigh_po_2p85_1_1/Rout
flabel metal1 49350 15082 49410 15142 1 FreeSans 1000 0 0 0 sky130_asc_res_xhigh_po_2p85_1_1/VPWR
flabel metal1 49350 13202 49410 13262 1 FreeSans 1000 0 0 0 sky130_asc_res_xhigh_po_2p85_1_1/VGND
flabel locali 52378 17096 52438 17156 1 FreeSans 1000 0 0 0 sky130_asc_pfet_01v8_lvt_60_0/GATE
flabel locali 52378 18682 52438 18722 1 FreeSans 1000 0 0 0 sky130_asc_pfet_01v8_lvt_60_0/SOURCE
flabel locali 52378 17202 52438 17262 1 FreeSans 1000 0 0 0 sky130_asc_pfet_01v8_lvt_60_0/DRAIN
flabel nwell 24732 18842 24792 18902 1 FreeSans 1000 0 0 0 sky130_asc_pfet_01v8_lvt_60_0/VPWR
flabel metal1 24732 16962 24890 17022 1 FreeSans 1000 0 0 0 sky130_asc_pfet_01v8_lvt_60_0/VGND
flabel metal1 23990 22052 24110 22172 1 FreeSans 600 0 0 0 sky130_asc_res_xhigh_po_2p85_1_24/Rin
flabel metal1 23990 21092 24110 21212 1 FreeSans 600 0 0 0 sky130_asc_res_xhigh_po_2p85_1_24/Rout
flabel metal1 23870 22602 23930 22662 1 FreeSans 1000 0 0 0 sky130_asc_res_xhigh_po_2p85_1_24/VPWR
flabel metal1 23870 20722 23930 20782 1 FreeSans 1000 0 0 0 sky130_asc_res_xhigh_po_2p85_1_24/VGND
flabel metal1 27322 22052 27442 22172 1 FreeSans 600 0 0 0 sky130_asc_res_xhigh_po_2p85_1_10/Rin
flabel metal1 27322 21092 27442 21212 1 FreeSans 600 0 0 0 sky130_asc_res_xhigh_po_2p85_1_10/Rout
flabel metal1 27202 22602 27262 22662 1 FreeSans 1000 0 0 0 sky130_asc_res_xhigh_po_2p85_1_10/VPWR
flabel metal1 27202 20722 27262 20782 1 FreeSans 1000 0 0 0 sky130_asc_res_xhigh_po_2p85_1_10/VGND
flabel metal1 48490 22052 48610 22172 1 FreeSans 600 0 0 0 sky130_asc_res_xhigh_po_2p85_1_20/Rin
flabel metal1 48490 21092 48610 21212 1 FreeSans 600 0 0 0 sky130_asc_res_xhigh_po_2p85_1_20/Rout
flabel metal1 48370 22602 48430 22662 1 FreeSans 1000 0 0 0 sky130_asc_res_xhigh_po_2p85_1_20/VPWR
flabel metal1 48370 20722 48430 20782 1 FreeSans 1000 0 0 0 sky130_asc_res_xhigh_po_2p85_1_20/VGND
flabel metal1 40258 22052 40378 22172 1 FreeSans 600 0 0 0 sky130_asc_res_xhigh_po_2p85_1_18/Rin
flabel metal1 40258 21092 40378 21212 1 FreeSans 600 0 0 0 sky130_asc_res_xhigh_po_2p85_1_18/Rout
flabel metal1 40138 22602 40198 22662 1 FreeSans 1000 0 0 0 sky130_asc_res_xhigh_po_2p85_1_18/VPWR
flabel metal1 40138 20722 40198 20782 1 FreeSans 1000 0 0 0 sky130_asc_res_xhigh_po_2p85_1_18/VGND
flabel metal1 37514 22052 37634 22172 1 FreeSans 600 0 0 0 sky130_asc_res_xhigh_po_2p85_1_15/Rin
flabel metal1 37514 21092 37634 21212 1 FreeSans 600 0 0 0 sky130_asc_res_xhigh_po_2p85_1_15/Rout
flabel metal1 37394 22602 37454 22662 1 FreeSans 1000 0 0 0 sky130_asc_res_xhigh_po_2p85_1_15/VPWR
flabel metal1 37394 20722 37454 20782 1 FreeSans 1000 0 0 0 sky130_asc_res_xhigh_po_2p85_1_15/VGND
flabel metal1 33300 22052 33420 22172 1 FreeSans 600 0 0 0 sky130_asc_res_xhigh_po_2p85_1_14/Rin
flabel metal1 33300 21092 33420 21212 1 FreeSans 600 0 0 0 sky130_asc_res_xhigh_po_2p85_1_14/Rout
flabel metal1 33180 22602 33240 22662 1 FreeSans 1000 0 0 0 sky130_asc_res_xhigh_po_2p85_1_14/VPWR
flabel metal1 33180 20722 33240 20782 1 FreeSans 1000 0 0 0 sky130_asc_res_xhigh_po_2p85_1_14/VGND
flabel metal1 30066 22052 30186 22172 1 FreeSans 600 0 0 0 sky130_asc_res_xhigh_po_2p85_1_11/Rin
flabel metal1 30066 21092 30186 21212 1 FreeSans 600 0 0 0 sky130_asc_res_xhigh_po_2p85_1_11/Rout
flabel metal1 29946 22602 30006 22662 1 FreeSans 1000 0 0 0 sky130_asc_res_xhigh_po_2p85_1_11/VPWR
flabel metal1 29946 20722 30006 20782 1 FreeSans 1000 0 0 0 sky130_asc_res_xhigh_po_2p85_1_11/VGND
flabel metal1 22520 25812 22640 25932 1 FreeSans 600 0 0 0 sky130_asc_res_xhigh_po_2p85_1_25/Rin
flabel metal1 22520 24852 22640 24972 1 FreeSans 600 0 0 0 sky130_asc_res_xhigh_po_2p85_1_25/Rout
flabel metal1 22400 26362 22460 26422 1 FreeSans 1000 0 0 0 sky130_asc_res_xhigh_po_2p85_1_25/VPWR
flabel metal1 22400 24482 22460 24542 1 FreeSans 1000 0 0 0 sky130_asc_res_xhigh_po_2p85_1_25/VGND
flabel locali 29538 24816 29598 24876 1 FreeSans 1000 0 0 0 sky130_asc_nfet_01v8_lvt_9_0/GATE
flabel locali 29538 26202 29598 26262 1 FreeSans 1000 0 0 0 sky130_asc_nfet_01v8_lvt_9_0/SOURCE
flabel locali 29538 24982 29598 25042 1 FreeSans 1000 0 0 0 sky130_asc_nfet_01v8_lvt_9_0/DRAIN
flabel metal1 25418 26362 25478 26422 1 FreeSans 1000 0 0 0 sky130_asc_nfet_01v8_lvt_9_0/VPWR
flabel metal1 25418 24482 25478 24542 1 FreeSans 1000 0 0 0 sky130_asc_nfet_01v8_lvt_9_0/VGND
flabel metal2 29926 26082 30126 26162 1 FreeSans 1000 0 0 0 sky130_asc_cap_mim_m3_1_0/Cin
flabel metal4 29948 24652 30108 24752 1 FreeSans 1000 0 0 0 sky130_asc_cap_mim_m3_1_0/Cout
flabel metal1 29928 26362 29988 26422 1 FreeSans 1000 0 0 0 sky130_asc_cap_mim_m3_1_0/VPWR
flabel metal1 29928 24482 29988 24542 1 FreeSans 1000 0 0 0 sky130_asc_cap_mim_m3_1_0/VGND
flabel metal1 43002 25812 43122 25932 1 FreeSans 600 0 0 0 sky130_asc_res_xhigh_po_2p85_1_16/Rin
flabel metal1 43002 24852 43122 24972 1 FreeSans 600 0 0 0 sky130_asc_res_xhigh_po_2p85_1_16/Rout
flabel metal1 42882 26362 42942 26422 1 FreeSans 1000 0 0 0 sky130_asc_res_xhigh_po_2p85_1_16/VPWR
flabel metal1 42882 24482 42942 24542 1 FreeSans 1000 0 0 0 sky130_asc_res_xhigh_po_2p85_1_16/VGND
flabel metal1 40258 25812 40378 25932 1 FreeSans 600 0 0 0 sky130_asc_res_xhigh_po_2p85_1_13/Rin
flabel metal1 40258 24852 40378 24972 1 FreeSans 600 0 0 0 sky130_asc_res_xhigh_po_2p85_1_13/Rout
flabel metal1 40138 26362 40198 26422 1 FreeSans 1000 0 0 0 sky130_asc_res_xhigh_po_2p85_1_13/VPWR
flabel metal1 40138 24482 40198 24542 1 FreeSans 1000 0 0 0 sky130_asc_res_xhigh_po_2p85_1_13/VGND
flabel metal1 37514 25812 37634 25932 1 FreeSans 600 0 0 0 sky130_asc_res_xhigh_po_2p85_1_12/Rin
flabel metal1 37514 24852 37634 24972 1 FreeSans 600 0 0 0 sky130_asc_res_xhigh_po_2p85_1_12/Rout
flabel metal1 37394 26362 37454 26422 1 FreeSans 1000 0 0 0 sky130_asc_res_xhigh_po_2p85_1_12/VPWR
flabel metal1 37394 24482 37454 24542 1 FreeSans 1000 0 0 0 sky130_asc_res_xhigh_po_2p85_1_12/VGND
flabel metal1 48490 25812 48610 25932 1 FreeSans 600 0 0 0 sky130_asc_res_xhigh_po_2p85_1_19/Rin
flabel metal1 48490 24852 48610 24972 1 FreeSans 600 0 0 0 sky130_asc_res_xhigh_po_2p85_1_19/Rout
flabel metal1 48370 26362 48430 26422 1 FreeSans 1000 0 0 0 sky130_asc_res_xhigh_po_2p85_1_19/VPWR
flabel metal1 48370 24482 48430 24542 1 FreeSans 1000 0 0 0 sky130_asc_res_xhigh_po_2p85_1_19/VGND
flabel metal1 45746 25812 45866 25932 1 FreeSans 600 0 0 0 sky130_asc_res_xhigh_po_2p85_1_17/Rin
flabel metal1 45746 24852 45866 24972 1 FreeSans 600 0 0 0 sky130_asc_res_xhigh_po_2p85_1_17/Rout
flabel metal1 45626 26362 45686 26422 1 FreeSans 1000 0 0 0 sky130_asc_res_xhigh_po_2p85_1_17/VPWR
flabel metal1 45626 24482 45686 24542 1 FreeSans 1000 0 0 0 sky130_asc_res_xhigh_po_2p85_1_17/VGND
flabel metal1 22128 29572 22248 29692 1 FreeSans 600 0 0 0 sky130_asc_res_xhigh_po_2p85_1_30/Rin
flabel metal1 22128 28612 22248 28732 1 FreeSans 600 0 0 0 sky130_asc_res_xhigh_po_2p85_1_30/Rout
flabel metal1 22008 30122 22068 30182 1 FreeSans 1000 0 0 0 sky130_asc_res_xhigh_po_2p85_1_30/VPWR
flabel metal1 22008 28242 22068 28302 1 FreeSans 1000 0 0 0 sky130_asc_res_xhigh_po_2p85_1_30/VGND
flabel metal1 16640 29572 16760 29692 1 FreeSans 600 0 0 0 sky130_asc_res_xhigh_po_2p85_1_23/Rin
flabel metal1 16640 28612 16760 28732 1 FreeSans 600 0 0 0 sky130_asc_res_xhigh_po_2p85_1_23/Rout
flabel metal1 16520 30122 16580 30182 1 FreeSans 1000 0 0 0 sky130_asc_res_xhigh_po_2p85_1_23/VPWR
flabel metal1 16520 28242 16580 28302 1 FreeSans 1000 0 0 0 sky130_asc_res_xhigh_po_2p85_1_23/VGND
flabel metal1 19384 29572 19504 29692 1 FreeSans 600 0 0 0 sky130_asc_res_xhigh_po_2p85_1_22/Rin
flabel metal1 19384 28612 19504 28732 1 FreeSans 600 0 0 0 sky130_asc_res_xhigh_po_2p85_1_22/Rout
flabel metal1 19264 30122 19324 30182 1 FreeSans 1000 0 0 0 sky130_asc_res_xhigh_po_2p85_1_22/VPWR
flabel metal1 19264 28242 19324 28302 1 FreeSans 1000 0 0 0 sky130_asc_res_xhigh_po_2p85_1_22/VGND
flabel metal1 27322 29572 27442 29692 1 FreeSans 600 0 0 0 sky130_asc_res_xhigh_po_2p85_1_9/Rin
flabel metal1 27322 28612 27442 28732 1 FreeSans 600 0 0 0 sky130_asc_res_xhigh_po_2p85_1_9/Rout
flabel metal1 27202 30122 27262 30182 1 FreeSans 1000 0 0 0 sky130_asc_res_xhigh_po_2p85_1_9/VPWR
flabel metal1 27202 28242 27262 28302 1 FreeSans 1000 0 0 0 sky130_asc_res_xhigh_po_2p85_1_9/VGND
flabel metal2 29926 29842 30126 29922 1 FreeSans 1000 0 0 0 sky130_asc_cap_mim_m3_1_2/Cin
flabel metal4 29948 28412 30108 28512 1 FreeSans 1000 0 0 0 sky130_asc_cap_mim_m3_1_2/Cout
flabel metal1 29928 30122 29988 30182 1 FreeSans 1000 0 0 0 sky130_asc_cap_mim_m3_1_2/VPWR
flabel metal1 29928 28242 29988 28302 1 FreeSans 1000 0 0 0 sky130_asc_cap_mim_m3_1_2/VGND
flabel locali 40288 28376 40348 28436 1 FreeSans 1000 0 0 0 sky130_asc_pfet_01v8_lvt_6_1/GATE
flabel locali 40288 29962 40348 30002 1 FreeSans 1000 0 0 0 sky130_asc_pfet_01v8_lvt_6_1/SOURCE
flabel locali 40288 28482 40348 28542 1 FreeSans 1000 0 0 0 sky130_asc_pfet_01v8_lvt_6_1/DRAIN
flabel nwell 37374 30122 37434 30182 1 FreeSans 1000 0 0 0 sky130_asc_pfet_01v8_lvt_6_1/VPWR
flabel metal1 37374 28242 37532 28302 1 FreeSans 1000 0 0 0 sky130_asc_pfet_01v8_lvt_6_1/VGND
flabel locali 51718 29168 51966 29272 0 FreeSans 500 0 0 0 sky130_asc_pnp_05v5_W3p40L3p40_8_2/sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_6/Emitter
flabel locali 51777 29794 51878 29843 0 FreeSans 500 0 0 0 sky130_asc_pnp_05v5_W3p40L3p40_8_2/sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_6/Collector
flabel locali 51754 29644 51872 29684 0 FreeSans 500 0 0 0 sky130_asc_pnp_05v5_W3p40L3p40_8_2/sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_6/Base
flabel locali 50378 29168 50626 29272 0 FreeSans 500 0 0 0 sky130_asc_pnp_05v5_W3p40L3p40_8_2/sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_5/Emitter
flabel locali 50437 29794 50538 29843 0 FreeSans 500 0 0 0 sky130_asc_pnp_05v5_W3p40L3p40_8_2/sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_5/Collector
flabel locali 50414 29644 50532 29684 0 FreeSans 500 0 0 0 sky130_asc_pnp_05v5_W3p40L3p40_8_2/sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_5/Base
flabel locali 49038 29168 49286 29272 0 FreeSans 500 0 0 0 sky130_asc_pnp_05v5_W3p40L3p40_8_2/sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_4/Emitter
flabel locali 49097 29794 49198 29843 0 FreeSans 500 0 0 0 sky130_asc_pnp_05v5_W3p40L3p40_8_2/sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_4/Collector
flabel locali 49074 29644 49192 29684 0 FreeSans 500 0 0 0 sky130_asc_pnp_05v5_W3p40L3p40_8_2/sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_4/Base
flabel locali 47698 29168 47946 29272 0 FreeSans 500 0 0 0 sky130_asc_pnp_05v5_W3p40L3p40_8_2/sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_3/Emitter
flabel locali 47757 29794 47858 29843 0 FreeSans 500 0 0 0 sky130_asc_pnp_05v5_W3p40L3p40_8_2/sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_3/Collector
flabel locali 47734 29644 47852 29684 0 FreeSans 500 0 0 0 sky130_asc_pnp_05v5_W3p40L3p40_8_2/sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_3/Base
flabel locali 46358 29168 46606 29272 0 FreeSans 500 0 0 0 sky130_asc_pnp_05v5_W3p40L3p40_8_2/sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_2/Emitter
flabel locali 46417 29794 46518 29843 0 FreeSans 500 0 0 0 sky130_asc_pnp_05v5_W3p40L3p40_8_2/sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_2/Collector
flabel locali 46394 29644 46512 29684 0 FreeSans 500 0 0 0 sky130_asc_pnp_05v5_W3p40L3p40_8_2/sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_2/Base
flabel locali 45018 29168 45266 29272 0 FreeSans 500 0 0 0 sky130_asc_pnp_05v5_W3p40L3p40_8_2/sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_1/Emitter
flabel locali 45077 29794 45178 29843 0 FreeSans 500 0 0 0 sky130_asc_pnp_05v5_W3p40L3p40_8_2/sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_1/Collector
flabel locali 45054 29644 45172 29684 0 FreeSans 500 0 0 0 sky130_asc_pnp_05v5_W3p40L3p40_8_2/sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_1/Base
flabel locali 43678 29168 43926 29272 0 FreeSans 500 0 0 0 sky130_asc_pnp_05v5_W3p40L3p40_8_2/sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0/Emitter
flabel locali 43737 29794 43838 29843 0 FreeSans 500 0 0 0 sky130_asc_pnp_05v5_W3p40L3p40_8_2/sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0/Collector
flabel locali 43714 29644 43832 29684 0 FreeSans 500 0 0 0 sky130_asc_pnp_05v5_W3p40L3p40_8_2/sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0/Base
flabel locali 42338 29168 42586 29272 0 FreeSans 500 0 0 0 sky130_asc_pnp_05v5_W3p40L3p40_8_2/xm1/Emitter
flabel locali 42397 29794 42498 29843 0 FreeSans 500 0 0 0 sky130_asc_pnp_05v5_W3p40L3p40_8_2/xm1/Collector
flabel locali 42374 29644 42492 29684 0 FreeSans 500 0 0 0 sky130_asc_pnp_05v5_W3p40L3p40_8_2/xm1/Base
flabel metal1 42324 29282 42564 29412 1 FreeSans 600 0 0 0 sky130_asc_pnp_05v5_W3p40L3p40_8_2/Emitter
flabel metal1 41974 29644 42214 29684 1 FreeSans 600 0 0 0 sky130_asc_pnp_05v5_W3p40L3p40_8_2/Base
flabel metal1 41810 29796 42050 29836 1 FreeSans 600 0 0 0 sky130_asc_pnp_05v5_W3p40L3p40_8_2/Collector
flabel metal1 41784 30122 41844 30182 1 FreeSans 1000 0 0 0 sky130_asc_pnp_05v5_W3p40L3p40_8_2/VPWR
flabel metal1 41784 28242 41844 28302 1 FreeSans 1000 0 0 0 sky130_asc_pnp_05v5_W3p40L3p40_8_2/VGND
flabel metal1 22129 33332 22249 33452 1 FreeSans 600 0 0 0 sky130_asc_res_xhigh_po_2p85_2_0/Rin
flabel metal1 22129 32372 22249 32492 1 FreeSans 600 0 0 0 sky130_asc_res_xhigh_po_2p85_2_0/Rout
flabel metal1 22010 33882 22070 33942 1 FreeSans 1000 0 0 0 sky130_asc_res_xhigh_po_2p85_2_0/VPWR
flabel metal1 22010 32002 22070 32062 1 FreeSans 1000 0 0 0 sky130_asc_res_xhigh_po_2p85_2_0/VGND
flabel metal1 19384 33332 19504 33452 1 FreeSans 600 0 0 0 sky130_asc_res_xhigh_po_2p85_1_28/Rin
flabel metal1 19384 32372 19504 32492 1 FreeSans 600 0 0 0 sky130_asc_res_xhigh_po_2p85_1_28/Rout
flabel metal1 19264 33882 19324 33942 1 FreeSans 1000 0 0 0 sky130_asc_res_xhigh_po_2p85_1_28/VPWR
flabel metal1 19264 32002 19324 32062 1 FreeSans 1000 0 0 0 sky130_asc_res_xhigh_po_2p85_1_28/VGND
flabel metal2 26202 33602 26402 33682 1 FreeSans 1000 0 0 0 sky130_asc_cap_mim_m3_1_4/Cin
flabel metal4 26224 32172 26384 32272 1 FreeSans 1000 0 0 0 sky130_asc_cap_mim_m3_1_4/Cout
flabel metal1 26204 33882 26264 33942 1 FreeSans 1000 0 0 0 sky130_asc_cap_mim_m3_1_4/VPWR
flabel metal1 26204 32002 26264 32062 1 FreeSans 1000 0 0 0 sky130_asc_cap_mim_m3_1_4/VGND
flabel locali 51718 32928 51966 33032 0 FreeSans 500 0 0 0 sky130_asc_pnp_05v5_W3p40L3p40_8_1/sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_6/Emitter
flabel locali 51777 33554 51878 33603 0 FreeSans 500 0 0 0 sky130_asc_pnp_05v5_W3p40L3p40_8_1/sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_6/Collector
flabel locali 51754 33404 51872 33444 0 FreeSans 500 0 0 0 sky130_asc_pnp_05v5_W3p40L3p40_8_1/sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_6/Base
flabel locali 50378 32928 50626 33032 0 FreeSans 500 0 0 0 sky130_asc_pnp_05v5_W3p40L3p40_8_1/sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_5/Emitter
flabel locali 50437 33554 50538 33603 0 FreeSans 500 0 0 0 sky130_asc_pnp_05v5_W3p40L3p40_8_1/sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_5/Collector
flabel locali 50414 33404 50532 33444 0 FreeSans 500 0 0 0 sky130_asc_pnp_05v5_W3p40L3p40_8_1/sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_5/Base
flabel locali 49038 32928 49286 33032 0 FreeSans 500 0 0 0 sky130_asc_pnp_05v5_W3p40L3p40_8_1/sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_4/Emitter
flabel locali 49097 33554 49198 33603 0 FreeSans 500 0 0 0 sky130_asc_pnp_05v5_W3p40L3p40_8_1/sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_4/Collector
flabel locali 49074 33404 49192 33444 0 FreeSans 500 0 0 0 sky130_asc_pnp_05v5_W3p40L3p40_8_1/sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_4/Base
flabel locali 47698 32928 47946 33032 0 FreeSans 500 0 0 0 sky130_asc_pnp_05v5_W3p40L3p40_8_1/sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_3/Emitter
flabel locali 47757 33554 47858 33603 0 FreeSans 500 0 0 0 sky130_asc_pnp_05v5_W3p40L3p40_8_1/sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_3/Collector
flabel locali 47734 33404 47852 33444 0 FreeSans 500 0 0 0 sky130_asc_pnp_05v5_W3p40L3p40_8_1/sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_3/Base
flabel locali 46358 32928 46606 33032 0 FreeSans 500 0 0 0 sky130_asc_pnp_05v5_W3p40L3p40_8_1/sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_2/Emitter
flabel locali 46417 33554 46518 33603 0 FreeSans 500 0 0 0 sky130_asc_pnp_05v5_W3p40L3p40_8_1/sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_2/Collector
flabel locali 46394 33404 46512 33444 0 FreeSans 500 0 0 0 sky130_asc_pnp_05v5_W3p40L3p40_8_1/sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_2/Base
flabel locali 45018 32928 45266 33032 0 FreeSans 500 0 0 0 sky130_asc_pnp_05v5_W3p40L3p40_8_1/sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_1/Emitter
flabel locali 45077 33554 45178 33603 0 FreeSans 500 0 0 0 sky130_asc_pnp_05v5_W3p40L3p40_8_1/sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_1/Collector
flabel locali 45054 33404 45172 33444 0 FreeSans 500 0 0 0 sky130_asc_pnp_05v5_W3p40L3p40_8_1/sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_1/Base
flabel locali 43678 32928 43926 33032 0 FreeSans 500 0 0 0 sky130_asc_pnp_05v5_W3p40L3p40_8_1/sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0/Emitter
flabel locali 43737 33554 43838 33603 0 FreeSans 500 0 0 0 sky130_asc_pnp_05v5_W3p40L3p40_8_1/sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0/Collector
flabel locali 43714 33404 43832 33444 0 FreeSans 500 0 0 0 sky130_asc_pnp_05v5_W3p40L3p40_8_1/sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0/Base
flabel locali 42338 32928 42586 33032 0 FreeSans 500 0 0 0 sky130_asc_pnp_05v5_W3p40L3p40_8_1/xm1/Emitter
flabel locali 42397 33554 42498 33603 0 FreeSans 500 0 0 0 sky130_asc_pnp_05v5_W3p40L3p40_8_1/xm1/Collector
flabel locali 42374 33404 42492 33444 0 FreeSans 500 0 0 0 sky130_asc_pnp_05v5_W3p40L3p40_8_1/xm1/Base
flabel metal1 42324 33042 42564 33172 1 FreeSans 600 0 0 0 sky130_asc_pnp_05v5_W3p40L3p40_8_1/Emitter
flabel metal1 41974 33404 42214 33444 1 FreeSans 600 0 0 0 sky130_asc_pnp_05v5_W3p40L3p40_8_1/Base
flabel metal1 41810 33556 42050 33596 1 FreeSans 600 0 0 0 sky130_asc_pnp_05v5_W3p40L3p40_8_1/Collector
flabel metal1 41784 33882 41844 33942 1 FreeSans 1000 0 0 0 sky130_asc_pnp_05v5_W3p40L3p40_8_1/VPWR
flabel metal1 41784 32002 41844 32062 1 FreeSans 1000 0 0 0 sky130_asc_pnp_05v5_W3p40L3p40_8_1/VGND
flabel metal2 33650 33602 33850 33682 1 FreeSans 1000 0 0 0 sky130_asc_cap_mim_m3_1_3/Cin
flabel metal4 33672 32172 33832 32272 1 FreeSans 1000 0 0 0 sky130_asc_cap_mim_m3_1_3/Cout
flabel metal1 33652 33882 33712 33942 1 FreeSans 1000 0 0 0 sky130_asc_cap_mim_m3_1_3/VPWR
flabel metal1 33652 32002 33712 32062 1 FreeSans 1000 0 0 0 sky130_asc_cap_mim_m3_1_3/VGND
flabel locali 12546 36688 12794 36792 0 FreeSans 500 0 0 0 sky130_asc_pnp_05v5_W3p40L3p40_1_0/xm1/Emitter
flabel locali 12605 37314 12706 37363 0 FreeSans 500 0 0 0 sky130_asc_pnp_05v5_W3p40L3p40_1_0/xm1/Collector
flabel locali 12582 37164 12700 37204 0 FreeSans 500 0 0 0 sky130_asc_pnp_05v5_W3p40L3p40_1_0/xm1/Base
flabel locali 12554 36802 12782 36932 1 FreeSans 600 0 0 0 sky130_asc_pnp_05v5_W3p40L3p40_1_0/Emitter
flabel locali 12766 37164 12886 37204 1 FreeSans 600 0 0 0 sky130_asc_pnp_05v5_W3p40L3p40_1_0/Base
flabel locali 12802 37316 12922 37356 1 FreeSans 600 0 0 0 sky130_asc_pnp_05v5_W3p40L3p40_1_0/Collector
flabel metal1 11992 37642 12052 37702 1 FreeSans 1000 0 0 0 sky130_asc_pnp_05v5_W3p40L3p40_1_0/VPWR
flabel metal1 11992 35762 12052 35822 1 FreeSans 1000 0 0 0 sky130_asc_pnp_05v5_W3p40L3p40_1_0/VGND
flabel metal1 13798 37092 13918 37212 1 FreeSans 600 0 0 0 sky130_asc_res_xhigh_po_2p85_1_26/Rin
flabel metal1 13798 36132 13918 36252 1 FreeSans 600 0 0 0 sky130_asc_res_xhigh_po_2p85_1_26/Rout
flabel metal1 13678 37642 13738 37702 1 FreeSans 1000 0 0 0 sky130_asc_res_xhigh_po_2p85_1_26/VPWR
flabel metal1 13678 35762 13738 35822 1 FreeSans 1000 0 0 0 sky130_asc_res_xhigh_po_2p85_1_26/VGND
flabel metal1 16542 37092 16662 37212 1 FreeSans 600 0 0 0 sky130_asc_res_xhigh_po_2p85_1_27/Rin
flabel metal1 16542 36132 16662 36252 1 FreeSans 600 0 0 0 sky130_asc_res_xhigh_po_2p85_1_27/Rout
flabel metal1 16422 37642 16482 37702 1 FreeSans 1000 0 0 0 sky130_asc_res_xhigh_po_2p85_1_27/VPWR
flabel metal1 16422 35762 16482 35822 1 FreeSans 1000 0 0 0 sky130_asc_res_xhigh_po_2p85_1_27/VGND
flabel metal1 19287 37092 19407 37212 1 FreeSans 600 0 0 0 sky130_asc_res_xhigh_po_2p85_2_1/Rin
flabel metal1 19287 36132 19407 36252 1 FreeSans 600 0 0 0 sky130_asc_res_xhigh_po_2p85_2_1/Rout
flabel metal1 19168 37642 19228 37702 1 FreeSans 1000 0 0 0 sky130_asc_res_xhigh_po_2p85_2_1/VPWR
flabel metal1 19168 35762 19228 35822 1 FreeSans 1000 0 0 0 sky130_asc_res_xhigh_po_2p85_2_1/VGND
flabel metal1 22618 37092 22738 37212 1 FreeSans 600 0 0 0 sky130_asc_res_xhigh_po_2p85_1_21/Rin
flabel metal1 22618 36132 22738 36252 1 FreeSans 600 0 0 0 sky130_asc_res_xhigh_po_2p85_1_21/Rout
flabel metal1 22498 37642 22558 37702 1 FreeSans 1000 0 0 0 sky130_asc_res_xhigh_po_2p85_1_21/VPWR
flabel metal1 22498 35762 22558 35822 1 FreeSans 1000 0 0 0 sky130_asc_res_xhigh_po_2p85_1_21/VGND
flabel locali 29538 36096 29598 36156 1 FreeSans 1000 0 0 0 sky130_asc_nfet_01v8_lvt_9_1/GATE
flabel locali 29538 37482 29598 37542 1 FreeSans 1000 0 0 0 sky130_asc_nfet_01v8_lvt_9_1/SOURCE
flabel locali 29538 36262 29598 36322 1 FreeSans 1000 0 0 0 sky130_asc_nfet_01v8_lvt_9_1/DRAIN
flabel metal1 25418 37642 25478 37702 1 FreeSans 1000 0 0 0 sky130_asc_nfet_01v8_lvt_9_1/VPWR
flabel metal1 25418 35762 25478 35822 1 FreeSans 1000 0 0 0 sky130_asc_nfet_01v8_lvt_9_1/VGND
flabel metal2 29926 37362 30126 37442 1 FreeSans 1000 0 0 0 sky130_asc_cap_mim_m3_1_1/Cin
flabel metal4 29948 35932 30108 36032 1 FreeSans 1000 0 0 0 sky130_asc_cap_mim_m3_1_1/Cout
flabel metal1 29928 37642 29988 37702 1 FreeSans 1000 0 0 0 sky130_asc_cap_mim_m3_1_1/VPWR
flabel metal1 29928 35762 29988 35822 1 FreeSans 1000 0 0 0 sky130_asc_cap_mim_m3_1_1/VGND
flabel locali 40288 35896 40348 35956 1 FreeSans 1000 0 0 0 sky130_asc_pfet_01v8_lvt_6_0/GATE
flabel locali 40288 37482 40348 37522 1 FreeSans 1000 0 0 0 sky130_asc_pfet_01v8_lvt_6_0/SOURCE
flabel locali 40288 36002 40348 36062 1 FreeSans 1000 0 0 0 sky130_asc_pfet_01v8_lvt_6_0/DRAIN
flabel nwell 37374 37642 37434 37702 1 FreeSans 1000 0 0 0 sky130_asc_pfet_01v8_lvt_6_0/VPWR
flabel metal1 37374 35762 37532 35822 1 FreeSans 1000 0 0 0 sky130_asc_pfet_01v8_lvt_6_0/VGND
flabel locali 51718 36688 51966 36792 0 FreeSans 500 0 0 0 sky130_asc_pnp_05v5_W3p40L3p40_8_0/sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_6/Emitter
flabel locali 51777 37314 51878 37363 0 FreeSans 500 0 0 0 sky130_asc_pnp_05v5_W3p40L3p40_8_0/sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_6/Collector
flabel locali 51754 37164 51872 37204 0 FreeSans 500 0 0 0 sky130_asc_pnp_05v5_W3p40L3p40_8_0/sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_6/Base
flabel locali 50378 36688 50626 36792 0 FreeSans 500 0 0 0 sky130_asc_pnp_05v5_W3p40L3p40_8_0/sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_5/Emitter
flabel locali 50437 37314 50538 37363 0 FreeSans 500 0 0 0 sky130_asc_pnp_05v5_W3p40L3p40_8_0/sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_5/Collector
flabel locali 50414 37164 50532 37204 0 FreeSans 500 0 0 0 sky130_asc_pnp_05v5_W3p40L3p40_8_0/sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_5/Base
flabel locali 49038 36688 49286 36792 0 FreeSans 500 0 0 0 sky130_asc_pnp_05v5_W3p40L3p40_8_0/sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_4/Emitter
flabel locali 49097 37314 49198 37363 0 FreeSans 500 0 0 0 sky130_asc_pnp_05v5_W3p40L3p40_8_0/sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_4/Collector
flabel locali 49074 37164 49192 37204 0 FreeSans 500 0 0 0 sky130_asc_pnp_05v5_W3p40L3p40_8_0/sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_4/Base
flabel locali 47698 36688 47946 36792 0 FreeSans 500 0 0 0 sky130_asc_pnp_05v5_W3p40L3p40_8_0/sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_3/Emitter
flabel locali 47757 37314 47858 37363 0 FreeSans 500 0 0 0 sky130_asc_pnp_05v5_W3p40L3p40_8_0/sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_3/Collector
flabel locali 47734 37164 47852 37204 0 FreeSans 500 0 0 0 sky130_asc_pnp_05v5_W3p40L3p40_8_0/sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_3/Base
flabel locali 46358 36688 46606 36792 0 FreeSans 500 0 0 0 sky130_asc_pnp_05v5_W3p40L3p40_8_0/sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_2/Emitter
flabel locali 46417 37314 46518 37363 0 FreeSans 500 0 0 0 sky130_asc_pnp_05v5_W3p40L3p40_8_0/sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_2/Collector
flabel locali 46394 37164 46512 37204 0 FreeSans 500 0 0 0 sky130_asc_pnp_05v5_W3p40L3p40_8_0/sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_2/Base
flabel locali 45018 36688 45266 36792 0 FreeSans 500 0 0 0 sky130_asc_pnp_05v5_W3p40L3p40_8_0/sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_1/Emitter
flabel locali 45077 37314 45178 37363 0 FreeSans 500 0 0 0 sky130_asc_pnp_05v5_W3p40L3p40_8_0/sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_1/Collector
flabel locali 45054 37164 45172 37204 0 FreeSans 500 0 0 0 sky130_asc_pnp_05v5_W3p40L3p40_8_0/sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_1/Base
flabel locali 43678 36688 43926 36792 0 FreeSans 500 0 0 0 sky130_asc_pnp_05v5_W3p40L3p40_8_0/sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0/Emitter
flabel locali 43737 37314 43838 37363 0 FreeSans 500 0 0 0 sky130_asc_pnp_05v5_W3p40L3p40_8_0/sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0/Collector
flabel locali 43714 37164 43832 37204 0 FreeSans 500 0 0 0 sky130_asc_pnp_05v5_W3p40L3p40_8_0/sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0/Base
flabel locali 42338 36688 42586 36792 0 FreeSans 500 0 0 0 sky130_asc_pnp_05v5_W3p40L3p40_8_0/xm1/Emitter
flabel locali 42397 37314 42498 37363 0 FreeSans 500 0 0 0 sky130_asc_pnp_05v5_W3p40L3p40_8_0/xm1/Collector
flabel locali 42374 37164 42492 37204 0 FreeSans 500 0 0 0 sky130_asc_pnp_05v5_W3p40L3p40_8_0/xm1/Base
flabel metal1 42324 36802 42564 36932 1 FreeSans 600 0 0 0 sky130_asc_pnp_05v5_W3p40L3p40_8_0/Emitter
flabel metal1 41974 37164 42214 37204 1 FreeSans 600 0 0 0 sky130_asc_pnp_05v5_W3p40L3p40_8_0/Base
flabel metal1 41810 37316 42050 37356 1 FreeSans 600 0 0 0 sky130_asc_pnp_05v5_W3p40L3p40_8_0/Collector
flabel metal1 41784 37642 41844 37702 1 FreeSans 1000 0 0 0 sky130_asc_pnp_05v5_W3p40L3p40_8_0/VPWR
flabel metal1 41784 35762 41844 35822 1 FreeSans 1000 0 0 0 sky130_asc_pnp_05v5_W3p40L3p40_8_0/VGND
flabel metal2 6308 41122 6508 41202 1 FreeSans 1000 0 0 0 sky130_asc_cap_mim_m3_1_5/Cin
flabel metal4 6330 39692 6490 39792 1 FreeSans 1000 0 0 0 sky130_asc_cap_mim_m3_1_5/Cout
flabel metal1 6310 41402 6370 41462 1 FreeSans 1000 0 0 0 sky130_asc_cap_mim_m3_1_5/VPWR
flabel metal1 6310 39522 6370 39582 1 FreeSans 1000 0 0 0 sky130_asc_cap_mim_m3_1_5/VGND
flabel metal2 15128 41122 15328 41202 1 FreeSans 1000 0 0 0 sky130_asc_cap_mim_m3_1_6/Cin
flabel metal4 15150 39692 15310 39792 1 FreeSans 1000 0 0 0 sky130_asc_cap_mim_m3_1_6/Cout
flabel metal1 15130 41402 15190 41462 1 FreeSans 1000 0 0 0 sky130_asc_cap_mim_m3_1_6/VPWR
flabel metal1 15130 39522 15190 39582 1 FreeSans 1000 0 0 0 sky130_asc_cap_mim_m3_1_6/VGND
flabel locali 28238 39656 28298 39716 1 FreeSans 1000 0 0 0 sky130_asc_pfet_01v8_lvt_12_0/GATE
flabel locali 28238 41242 28298 41282 1 FreeSans 1000 0 0 0 sky130_asc_pfet_01v8_lvt_12_0/SOURCE
flabel locali 28238 39762 28298 39822 1 FreeSans 1000 0 0 0 sky130_asc_pfet_01v8_lvt_12_0/DRAIN
flabel nwell 22576 41402 22636 41462 1 FreeSans 1000 0 0 0 sky130_asc_pfet_01v8_lvt_12_0/VPWR
flabel metal1 22576 39522 22734 39582 1 FreeSans 1000 0 0 0 sky130_asc_pfet_01v8_lvt_12_0/VGND
flabel locali 34902 39656 34962 39716 1 FreeSans 1000 0 0 0 sky130_asc_pfet_01v8_lvt_12_1/GATE
flabel locali 34902 41242 34962 41282 1 FreeSans 1000 0 0 0 sky130_asc_pfet_01v8_lvt_12_1/SOURCE
flabel locali 34902 39762 34962 39822 1 FreeSans 1000 0 0 0 sky130_asc_pfet_01v8_lvt_12_1/DRAIN
flabel nwell 29240 41402 29300 41462 1 FreeSans 1000 0 0 0 sky130_asc_pfet_01v8_lvt_12_1/VPWR
flabel metal1 29240 39522 29398 39582 1 FreeSans 1000 0 0 0 sky130_asc_pfet_01v8_lvt_12_1/VGND
flabel locali 41396 39856 41456 39916 1 FreeSans 1000 0 0 0 sky130_asc_nfet_01v8_lvt_9_2/GATE
flabel locali 41396 41242 41456 41302 1 FreeSans 1000 0 0 0 sky130_asc_nfet_01v8_lvt_9_2/SOURCE
flabel locali 41396 40022 41456 40082 1 FreeSans 1000 0 0 0 sky130_asc_nfet_01v8_lvt_9_2/DRAIN
flabel metal1 37276 41402 37336 41462 1 FreeSans 1000 0 0 0 sky130_asc_nfet_01v8_lvt_9_2/VPWR
flabel metal1 37276 39522 37336 39582 1 FreeSans 1000 0 0 0 sky130_asc_nfet_01v8_lvt_9_2/VGND
flabel locali 51718 40448 51966 40552 0 FreeSans 500 0 0 0 sky130_asc_pnp_05v5_W3p40L3p40_8_3/sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_6/Emitter
flabel locali 51777 41074 51878 41123 0 FreeSans 500 0 0 0 sky130_asc_pnp_05v5_W3p40L3p40_8_3/sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_6/Collector
flabel locali 51754 40924 51872 40964 0 FreeSans 500 0 0 0 sky130_asc_pnp_05v5_W3p40L3p40_8_3/sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_6/Base
flabel locali 50378 40448 50626 40552 0 FreeSans 500 0 0 0 sky130_asc_pnp_05v5_W3p40L3p40_8_3/sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_5/Emitter
flabel locali 50437 41074 50538 41123 0 FreeSans 500 0 0 0 sky130_asc_pnp_05v5_W3p40L3p40_8_3/sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_5/Collector
flabel locali 50414 40924 50532 40964 0 FreeSans 500 0 0 0 sky130_asc_pnp_05v5_W3p40L3p40_8_3/sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_5/Base
flabel locali 49038 40448 49286 40552 0 FreeSans 500 0 0 0 sky130_asc_pnp_05v5_W3p40L3p40_8_3/sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_4/Emitter
flabel locali 49097 41074 49198 41123 0 FreeSans 500 0 0 0 sky130_asc_pnp_05v5_W3p40L3p40_8_3/sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_4/Collector
flabel locali 49074 40924 49192 40964 0 FreeSans 500 0 0 0 sky130_asc_pnp_05v5_W3p40L3p40_8_3/sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_4/Base
flabel locali 47698 40448 47946 40552 0 FreeSans 500 0 0 0 sky130_asc_pnp_05v5_W3p40L3p40_8_3/sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_3/Emitter
flabel locali 47757 41074 47858 41123 0 FreeSans 500 0 0 0 sky130_asc_pnp_05v5_W3p40L3p40_8_3/sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_3/Collector
flabel locali 47734 40924 47852 40964 0 FreeSans 500 0 0 0 sky130_asc_pnp_05v5_W3p40L3p40_8_3/sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_3/Base
flabel locali 46358 40448 46606 40552 0 FreeSans 500 0 0 0 sky130_asc_pnp_05v5_W3p40L3p40_8_3/sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_2/Emitter
flabel locali 46417 41074 46518 41123 0 FreeSans 500 0 0 0 sky130_asc_pnp_05v5_W3p40L3p40_8_3/sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_2/Collector
flabel locali 46394 40924 46512 40964 0 FreeSans 500 0 0 0 sky130_asc_pnp_05v5_W3p40L3p40_8_3/sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_2/Base
flabel locali 45018 40448 45266 40552 0 FreeSans 500 0 0 0 sky130_asc_pnp_05v5_W3p40L3p40_8_3/sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_1/Emitter
flabel locali 45077 41074 45178 41123 0 FreeSans 500 0 0 0 sky130_asc_pnp_05v5_W3p40L3p40_8_3/sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_1/Collector
flabel locali 45054 40924 45172 40964 0 FreeSans 500 0 0 0 sky130_asc_pnp_05v5_W3p40L3p40_8_3/sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_1/Base
flabel locali 43678 40448 43926 40552 0 FreeSans 500 0 0 0 sky130_asc_pnp_05v5_W3p40L3p40_8_3/sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0/Emitter
flabel locali 43737 41074 43838 41123 0 FreeSans 500 0 0 0 sky130_asc_pnp_05v5_W3p40L3p40_8_3/sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0/Collector
flabel locali 43714 40924 43832 40964 0 FreeSans 500 0 0 0 sky130_asc_pnp_05v5_W3p40L3p40_8_3/sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0/Base
flabel locali 42338 40448 42586 40552 0 FreeSans 500 0 0 0 sky130_asc_pnp_05v5_W3p40L3p40_8_3/xm1/Emitter
flabel locali 42397 41074 42498 41123 0 FreeSans 500 0 0 0 sky130_asc_pnp_05v5_W3p40L3p40_8_3/xm1/Collector
flabel locali 42374 40924 42492 40964 0 FreeSans 500 0 0 0 sky130_asc_pnp_05v5_W3p40L3p40_8_3/xm1/Base
flabel metal1 42324 40562 42564 40692 1 FreeSans 600 0 0 0 sky130_asc_pnp_05v5_W3p40L3p40_8_3/Emitter
flabel metal1 41974 40924 42214 40964 1 FreeSans 600 0 0 0 sky130_asc_pnp_05v5_W3p40L3p40_8_3/Base
flabel metal1 41810 41076 42050 41116 1 FreeSans 600 0 0 0 sky130_asc_pnp_05v5_W3p40L3p40_8_3/Collector
flabel metal1 41784 41402 41844 41462 1 FreeSans 1000 0 0 0 sky130_asc_pnp_05v5_W3p40L3p40_8_3/VPWR
flabel metal1 41784 39522 41844 39582 1 FreeSans 1000 0 0 0 sky130_asc_pnp_05v5_W3p40L3p40_8_3/VGND
flabel locali 14574 43456 14634 43516 1 FreeSans 1000 0 0 0 sky130_asc_nfet_01v8_lvt_1_1/GATE
flabel locali 14574 45002 14634 45062 1 FreeSans 1000 0 0 0 sky130_asc_nfet_01v8_lvt_1_1/SOURCE
flabel locali 14574 43682 14634 43742 1 FreeSans 1000 0 0 0 sky130_asc_nfet_01v8_lvt_1_1/DRAIN
flabel metal1 14118 45162 14178 45222 1 FreeSans 1000 0 0 0 sky130_asc_nfet_01v8_lvt_1_1/VPWR
flabel metal1 14118 43282 14178 43342 1 FreeSans 1000 0 0 0 sky130_asc_nfet_01v8_lvt_1_1/VGND
flabel metal2 5916 44882 6116 44962 1 FreeSans 1000 0 0 0 sky130_asc_cap_mim_m3_1_7/Cin
flabel metal4 5938 43452 6098 43552 1 FreeSans 1000 0 0 0 sky130_asc_cap_mim_m3_1_7/Cout
flabel metal1 5918 45162 5978 45222 1 FreeSans 1000 0 0 0 sky130_asc_cap_mim_m3_1_7/VPWR
flabel metal1 5918 43282 5978 43342 1 FreeSans 1000 0 0 0 sky130_asc_cap_mim_m3_1_7/VGND
flabel locali 42578 43416 42638 43476 1 FreeSans 1000 0 0 0 sky130_asc_pfet_01v8_lvt_60_2/GATE
flabel locali 42578 45002 42638 45042 1 FreeSans 1000 0 0 0 sky130_asc_pfet_01v8_lvt_60_2/SOURCE
flabel locali 42578 43522 42638 43582 1 FreeSans 1000 0 0 0 sky130_asc_pfet_01v8_lvt_60_2/DRAIN
flabel nwell 14932 45162 14992 45222 1 FreeSans 1000 0 0 0 sky130_asc_pfet_01v8_lvt_60_2/VPWR
flabel metal1 14932 43282 15090 43342 1 FreeSans 1000 0 0 0 sky130_asc_pfet_01v8_lvt_60_2/VGND
flabel locali 51554 44208 51802 44312 0 FreeSans 500 0 0 0 sky130_asc_pnp_05v5_W3p40L3p40_7_0/sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_5/Emitter
flabel locali 51613 44834 51714 44883 0 FreeSans 500 0 0 0 sky130_asc_pnp_05v5_W3p40L3p40_7_0/sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_5/Collector
flabel locali 51590 44684 51708 44724 0 FreeSans 500 0 0 0 sky130_asc_pnp_05v5_W3p40L3p40_7_0/sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_5/Base
flabel locali 50214 44208 50462 44312 0 FreeSans 500 0 0 0 sky130_asc_pnp_05v5_W3p40L3p40_7_0/sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_4/Emitter
flabel locali 50273 44834 50374 44883 0 FreeSans 500 0 0 0 sky130_asc_pnp_05v5_W3p40L3p40_7_0/sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_4/Collector
flabel locali 50250 44684 50368 44724 0 FreeSans 500 0 0 0 sky130_asc_pnp_05v5_W3p40L3p40_7_0/sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_4/Base
flabel locali 48874 44208 49122 44312 0 FreeSans 500 0 0 0 sky130_asc_pnp_05v5_W3p40L3p40_7_0/sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_3/Emitter
flabel locali 48933 44834 49034 44883 0 FreeSans 500 0 0 0 sky130_asc_pnp_05v5_W3p40L3p40_7_0/sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_3/Collector
flabel locali 48910 44684 49028 44724 0 FreeSans 500 0 0 0 sky130_asc_pnp_05v5_W3p40L3p40_7_0/sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_3/Base
flabel locali 47534 44208 47782 44312 0 FreeSans 500 0 0 0 sky130_asc_pnp_05v5_W3p40L3p40_7_0/sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_2/Emitter
flabel locali 47593 44834 47694 44883 0 FreeSans 500 0 0 0 sky130_asc_pnp_05v5_W3p40L3p40_7_0/sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_2/Collector
flabel locali 47570 44684 47688 44724 0 FreeSans 500 0 0 0 sky130_asc_pnp_05v5_W3p40L3p40_7_0/sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_2/Base
flabel locali 46194 44208 46442 44312 0 FreeSans 500 0 0 0 sky130_asc_pnp_05v5_W3p40L3p40_7_0/sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_1/Emitter
flabel locali 46253 44834 46354 44883 0 FreeSans 500 0 0 0 sky130_asc_pnp_05v5_W3p40L3p40_7_0/sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_1/Collector
flabel locali 46230 44684 46348 44724 0 FreeSans 500 0 0 0 sky130_asc_pnp_05v5_W3p40L3p40_7_0/sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_1/Base
flabel locali 44854 44208 45102 44312 0 FreeSans 500 0 0 0 sky130_asc_pnp_05v5_W3p40L3p40_7_0/sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0/Emitter
flabel locali 44913 44834 45014 44883 0 FreeSans 500 0 0 0 sky130_asc_pnp_05v5_W3p40L3p40_7_0/sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0/Collector
flabel locali 44890 44684 45008 44724 0 FreeSans 500 0 0 0 sky130_asc_pnp_05v5_W3p40L3p40_7_0/sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0/Base
flabel locali 43514 44208 43762 44312 0 FreeSans 500 0 0 0 sky130_asc_pnp_05v5_W3p40L3p40_7_0/xm1/Emitter
flabel locali 43573 44834 43674 44883 0 FreeSans 500 0 0 0 sky130_asc_pnp_05v5_W3p40L3p40_7_0/xm1/Collector
flabel locali 43550 44684 43668 44724 0 FreeSans 500 0 0 0 sky130_asc_pnp_05v5_W3p40L3p40_7_0/xm1/Base
flabel metal1 43500 44322 43740 44452 1 FreeSans 600 0 0 0 sky130_asc_pnp_05v5_W3p40L3p40_7_0/Emitter
flabel metal1 43150 44684 43390 44724 1 FreeSans 600 0 0 0 sky130_asc_pnp_05v5_W3p40L3p40_7_0/Base
flabel metal1 42986 44836 43226 44876 1 FreeSans 600 0 0 0 sky130_asc_pnp_05v5_W3p40L3p40_7_0/Collector
flabel metal1 42960 45162 43020 45222 1 FreeSans 1000 0 0 0 sky130_asc_pnp_05v5_W3p40L3p40_7_0/VPWR
flabel metal1 42960 43282 43020 43342 1 FreeSans 1000 0 0 0 sky130_asc_pnp_05v5_W3p40L3p40_7_0/VGND
flabel metal2 13364 48642 13564 48722 1 FreeSans 1000 0 0 0 sky130_asc_cap_mim_m3_1_9/Cin
flabel metal4 13386 47212 13546 47312 1 FreeSans 1000 0 0 0 sky130_asc_cap_mim_m3_1_9/Cout
flabel metal1 13366 48922 13426 48982 1 FreeSans 1000 0 0 0 sky130_asc_cap_mim_m3_1_9/VPWR
flabel metal1 13366 47042 13426 47102 1 FreeSans 1000 0 0 0 sky130_asc_cap_mim_m3_1_9/VGND
flabel metal2 5916 48642 6116 48722 1 FreeSans 1000 0 0 0 sky130_asc_cap_mim_m3_1_8/Cin
flabel metal4 5938 47212 6098 47312 1 FreeSans 1000 0 0 0 sky130_asc_cap_mim_m3_1_8/Cout
flabel metal1 5918 48922 5978 48982 1 FreeSans 1000 0 0 0 sky130_asc_cap_mim_m3_1_8/VPWR
flabel metal1 5918 47042 5978 47102 1 FreeSans 1000 0 0 0 sky130_asc_cap_mim_m3_1_8/VGND
flabel metal1 20952 48372 21072 48492 1 FreeSans 600 0 0 0 sky130_asc_res_xhigh_po_2p85_1_29/Rin
flabel metal1 20952 47412 21072 47532 1 FreeSans 600 0 0 0 sky130_asc_res_xhigh_po_2p85_1_29/Rout
flabel metal1 20832 48922 20892 48982 1 FreeSans 1000 0 0 0 sky130_asc_res_xhigh_po_2p85_1_29/VPWR
flabel metal1 20832 47042 20892 47102 1 FreeSans 1000 0 0 0 sky130_asc_res_xhigh_po_2p85_1_29/VGND
flabel locali 24374 47216 24434 47276 1 FreeSans 1000 0 0 0 sky130_asc_nfet_01v8_lvt_1_0/GATE
flabel locali 24374 48762 24434 48822 1 FreeSans 1000 0 0 0 sky130_asc_nfet_01v8_lvt_1_0/SOURCE
flabel locali 24374 47442 24434 47502 1 FreeSans 1000 0 0 0 sky130_asc_nfet_01v8_lvt_1_0/DRAIN
flabel metal1 23918 48922 23978 48982 1 FreeSans 1000 0 0 0 sky130_asc_nfet_01v8_lvt_1_0/VPWR
flabel metal1 23918 47042 23978 47102 1 FreeSans 1000 0 0 0 sky130_asc_nfet_01v8_lvt_1_0/VGND
flabel locali 52378 47176 52438 47236 1 FreeSans 1000 0 0 0 sky130_asc_pfet_01v8_lvt_60_1/GATE
flabel locali 52378 48762 52438 48802 1 FreeSans 1000 0 0 0 sky130_asc_pfet_01v8_lvt_60_1/SOURCE
flabel locali 52378 47282 52438 47342 1 FreeSans 1000 0 0 0 sky130_asc_pfet_01v8_lvt_60_1/DRAIN
flabel nwell 24732 48922 24792 48982 1 FreeSans 1000 0 0 0 sky130_asc_pfet_01v8_lvt_60_1/VPWR
flabel metal1 24732 47042 24890 47102 1 FreeSans 1000 0 0 0 sky130_asc_pfet_01v8_lvt_60_1/VGND
<< end >>
