magic
tech sky130A
magscale 1 2
timestamp 1652297564
<< pwell >>
rect 0 1457 1340 1610
rect 0 423 153 1457
rect 1187 423 1340 1457
rect 0 270 1340 423
<< nbase >>
rect 153 423 1187 1457
<< pdiff >>
rect 330 1228 1010 1280
rect 330 1194 384 1228
rect 418 1194 474 1228
rect 508 1194 564 1228
rect 598 1194 654 1228
rect 688 1194 744 1228
rect 778 1194 834 1228
rect 868 1194 924 1228
rect 958 1194 1010 1228
rect 330 1138 1010 1194
rect 330 1104 384 1138
rect 418 1104 474 1138
rect 508 1104 564 1138
rect 598 1104 654 1138
rect 688 1104 744 1138
rect 778 1104 834 1138
rect 868 1104 924 1138
rect 958 1104 1010 1138
rect 330 1048 1010 1104
rect 330 1014 384 1048
rect 418 1014 474 1048
rect 508 1014 564 1048
rect 598 1014 654 1048
rect 688 1014 744 1048
rect 778 1014 834 1048
rect 868 1014 924 1048
rect 958 1014 1010 1048
rect 330 958 1010 1014
rect 330 924 384 958
rect 418 924 474 958
rect 508 924 564 958
rect 598 924 654 958
rect 688 924 744 958
rect 778 924 834 958
rect 868 924 924 958
rect 958 924 1010 958
rect 330 868 1010 924
rect 330 834 384 868
rect 418 834 474 868
rect 508 834 564 868
rect 598 834 654 868
rect 688 834 744 868
rect 778 834 834 868
rect 868 834 924 868
rect 958 834 1010 868
rect 330 778 1010 834
rect 330 744 384 778
rect 418 744 474 778
rect 508 744 564 778
rect 598 744 654 778
rect 688 744 744 778
rect 778 744 834 778
rect 868 744 924 778
rect 958 744 1010 778
rect 330 688 1010 744
rect 330 654 384 688
rect 418 654 474 688
rect 508 654 564 688
rect 598 654 654 688
rect 688 654 744 688
rect 778 654 834 688
rect 868 654 924 688
rect 958 654 1010 688
rect 330 600 1010 654
<< pdiffc >>
rect 384 1194 418 1228
rect 474 1194 508 1228
rect 564 1194 598 1228
rect 654 1194 688 1228
rect 744 1194 778 1228
rect 834 1194 868 1228
rect 924 1194 958 1228
rect 384 1104 418 1138
rect 474 1104 508 1138
rect 564 1104 598 1138
rect 654 1104 688 1138
rect 744 1104 778 1138
rect 834 1104 868 1138
rect 924 1104 958 1138
rect 384 1014 418 1048
rect 474 1014 508 1048
rect 564 1014 598 1048
rect 654 1014 688 1048
rect 744 1014 778 1048
rect 834 1014 868 1048
rect 924 1014 958 1048
rect 384 924 418 958
rect 474 924 508 958
rect 564 924 598 958
rect 654 924 688 958
rect 744 924 778 958
rect 834 924 868 958
rect 924 924 958 958
rect 384 834 418 868
rect 474 834 508 868
rect 564 834 598 868
rect 654 834 688 868
rect 744 834 778 868
rect 834 834 868 868
rect 924 834 958 868
rect 384 744 418 778
rect 474 744 508 778
rect 564 744 598 778
rect 654 744 688 778
rect 744 744 778 778
rect 834 744 868 778
rect 924 744 958 778
rect 384 654 418 688
rect 474 654 508 688
rect 564 654 598 688
rect 654 654 688 688
rect 744 654 778 688
rect 834 654 868 688
rect 924 654 958 688
<< psubdiff >>
rect 26 1549 1314 1584
rect 26 1526 156 1549
rect 26 1492 60 1526
rect 94 1515 156 1526
rect 190 1515 246 1549
rect 280 1515 336 1549
rect 370 1515 426 1549
rect 460 1515 516 1549
rect 550 1515 606 1549
rect 640 1515 696 1549
rect 730 1515 786 1549
rect 820 1515 876 1549
rect 910 1515 966 1549
rect 1000 1515 1056 1549
rect 1090 1515 1146 1549
rect 1180 1526 1314 1549
rect 1180 1515 1247 1526
rect 94 1492 1247 1515
rect 1281 1492 1314 1526
rect 26 1483 1314 1492
rect 26 1436 127 1483
rect 26 1402 60 1436
rect 94 1402 127 1436
rect 1213 1436 1314 1483
rect 26 1346 127 1402
rect 26 1312 60 1346
rect 94 1312 127 1346
rect 26 1256 127 1312
rect 26 1222 60 1256
rect 94 1222 127 1256
rect 26 1166 127 1222
rect 26 1132 60 1166
rect 94 1132 127 1166
rect 26 1076 127 1132
rect 26 1042 60 1076
rect 94 1042 127 1076
rect 26 986 127 1042
rect 26 952 60 986
rect 94 952 127 986
rect 26 896 127 952
rect 26 862 60 896
rect 94 862 127 896
rect 26 806 127 862
rect 26 772 60 806
rect 94 772 127 806
rect 26 716 127 772
rect 26 682 60 716
rect 94 682 127 716
rect 26 626 127 682
rect 26 592 60 626
rect 94 592 127 626
rect 26 536 127 592
rect 26 502 60 536
rect 94 502 127 536
rect 26 446 127 502
rect 1213 1402 1247 1436
rect 1281 1402 1314 1436
rect 1213 1346 1314 1402
rect 1213 1312 1247 1346
rect 1281 1312 1314 1346
rect 1213 1256 1314 1312
rect 1213 1222 1247 1256
rect 1281 1222 1314 1256
rect 1213 1166 1314 1222
rect 1213 1132 1247 1166
rect 1281 1132 1314 1166
rect 1213 1076 1314 1132
rect 1213 1042 1247 1076
rect 1281 1042 1314 1076
rect 1213 986 1314 1042
rect 1213 952 1247 986
rect 1281 952 1314 986
rect 1213 896 1314 952
rect 1213 862 1247 896
rect 1281 862 1314 896
rect 1213 806 1314 862
rect 1213 772 1247 806
rect 1281 772 1314 806
rect 1213 716 1314 772
rect 1213 682 1247 716
rect 1281 682 1314 716
rect 1213 626 1314 682
rect 1213 592 1247 626
rect 1281 592 1314 626
rect 1213 536 1314 592
rect 1213 502 1247 536
rect 1281 502 1314 536
rect 26 412 60 446
rect 94 412 127 446
rect 26 397 127 412
rect 1213 446 1314 502
rect 1213 412 1247 446
rect 1281 412 1314 446
rect 1213 397 1314 412
rect 26 362 1314 397
rect 26 328 156 362
rect 190 328 246 362
rect 280 328 336 362
rect 370 328 426 362
rect 460 328 516 362
rect 550 328 606 362
rect 640 328 696 362
rect 730 328 786 362
rect 820 328 876 362
rect 910 328 966 362
rect 1000 328 1056 362
rect 1090 328 1146 362
rect 1180 328 1314 362
rect 26 296 1314 328
<< nsubdiff >>
rect 189 1402 1151 1421
rect 189 1368 320 1402
rect 354 1368 410 1402
rect 444 1368 500 1402
rect 534 1368 590 1402
rect 624 1368 680 1402
rect 714 1368 770 1402
rect 804 1368 860 1402
rect 894 1368 950 1402
rect 984 1368 1040 1402
rect 1074 1368 1151 1402
rect 189 1349 1151 1368
rect 189 1345 261 1349
rect 189 1311 208 1345
rect 242 1311 261 1345
rect 189 1255 261 1311
rect 1079 1326 1151 1349
rect 1079 1292 1098 1326
rect 1132 1292 1151 1326
rect 189 1221 208 1255
rect 242 1221 261 1255
rect 189 1165 261 1221
rect 189 1131 208 1165
rect 242 1131 261 1165
rect 189 1075 261 1131
rect 189 1041 208 1075
rect 242 1041 261 1075
rect 189 985 261 1041
rect 189 951 208 985
rect 242 951 261 985
rect 189 895 261 951
rect 189 861 208 895
rect 242 861 261 895
rect 189 805 261 861
rect 189 771 208 805
rect 242 771 261 805
rect 189 715 261 771
rect 189 681 208 715
rect 242 681 261 715
rect 189 625 261 681
rect 189 591 208 625
rect 242 591 261 625
rect 1079 1236 1151 1292
rect 1079 1202 1098 1236
rect 1132 1202 1151 1236
rect 1079 1146 1151 1202
rect 1079 1112 1098 1146
rect 1132 1112 1151 1146
rect 1079 1056 1151 1112
rect 1079 1022 1098 1056
rect 1132 1022 1151 1056
rect 1079 966 1151 1022
rect 1079 932 1098 966
rect 1132 932 1151 966
rect 1079 876 1151 932
rect 1079 842 1098 876
rect 1132 842 1151 876
rect 1079 786 1151 842
rect 1079 752 1098 786
rect 1132 752 1151 786
rect 1079 696 1151 752
rect 1079 662 1098 696
rect 1132 662 1151 696
rect 1079 606 1151 662
rect 189 531 261 591
rect 1079 572 1098 606
rect 1132 572 1151 606
rect 1079 531 1151 572
rect 189 512 1151 531
rect 189 478 286 512
rect 320 478 376 512
rect 410 478 466 512
rect 500 478 556 512
rect 590 478 646 512
rect 680 478 736 512
rect 770 478 826 512
rect 860 478 916 512
rect 950 478 1006 512
rect 1040 478 1151 512
rect 189 459 1151 478
<< psubdiffcont >>
rect 60 1492 94 1526
rect 156 1515 190 1549
rect 246 1515 280 1549
rect 336 1515 370 1549
rect 426 1515 460 1549
rect 516 1515 550 1549
rect 606 1515 640 1549
rect 696 1515 730 1549
rect 786 1515 820 1549
rect 876 1515 910 1549
rect 966 1515 1000 1549
rect 1056 1515 1090 1549
rect 1146 1515 1180 1549
rect 1247 1492 1281 1526
rect 60 1402 94 1436
rect 60 1312 94 1346
rect 60 1222 94 1256
rect 60 1132 94 1166
rect 60 1042 94 1076
rect 60 952 94 986
rect 60 862 94 896
rect 60 772 94 806
rect 60 682 94 716
rect 60 592 94 626
rect 60 502 94 536
rect 1247 1402 1281 1436
rect 1247 1312 1281 1346
rect 1247 1222 1281 1256
rect 1247 1132 1281 1166
rect 1247 1042 1281 1076
rect 1247 952 1281 986
rect 1247 862 1281 896
rect 1247 772 1281 806
rect 1247 682 1281 716
rect 1247 592 1281 626
rect 1247 502 1281 536
rect 60 412 94 446
rect 1247 412 1281 446
rect 156 328 190 362
rect 246 328 280 362
rect 336 328 370 362
rect 426 328 460 362
rect 516 328 550 362
rect 606 328 640 362
rect 696 328 730 362
rect 786 328 820 362
rect 876 328 910 362
rect 966 328 1000 362
rect 1056 328 1090 362
rect 1146 328 1180 362
<< nsubdiffcont >>
rect 320 1368 354 1402
rect 410 1368 444 1402
rect 500 1368 534 1402
rect 590 1368 624 1402
rect 680 1368 714 1402
rect 770 1368 804 1402
rect 860 1368 894 1402
rect 950 1368 984 1402
rect 1040 1368 1074 1402
rect 208 1311 242 1345
rect 1098 1292 1132 1326
rect 208 1221 242 1255
rect 208 1131 242 1165
rect 208 1041 242 1075
rect 208 951 242 985
rect 208 861 242 895
rect 208 771 242 805
rect 208 681 242 715
rect 208 591 242 625
rect 1098 1202 1132 1236
rect 1098 1112 1132 1146
rect 1098 1022 1132 1056
rect 1098 932 1132 966
rect 1098 842 1132 876
rect 1098 752 1132 786
rect 1098 662 1132 696
rect 1098 572 1132 606
rect 286 478 320 512
rect 376 478 410 512
rect 466 478 500 512
rect 556 478 590 512
rect 646 478 680 512
rect 736 478 770 512
rect 826 478 860 512
rect 916 478 950 512
rect 1006 478 1040 512
<< locali >>
rect 0 1850 170 1910
rect 230 1850 370 1910
rect 430 1850 570 1910
rect 630 1850 770 1910
rect 830 1850 970 1910
rect 1030 1850 1170 1910
rect 1230 1850 1340 1910
rect 26 1549 1314 1584
rect 26 1526 156 1549
rect 26 1492 60 1526
rect 94 1515 156 1526
rect 190 1515 246 1549
rect 280 1515 336 1549
rect 370 1515 426 1549
rect 460 1515 516 1549
rect 550 1515 606 1549
rect 640 1515 696 1549
rect 730 1515 786 1549
rect 820 1515 876 1549
rect 910 1515 966 1549
rect 1000 1515 1056 1549
rect 1090 1515 1146 1549
rect 1180 1526 1314 1549
rect 1180 1515 1247 1526
rect 94 1492 1247 1515
rect 1281 1492 1314 1526
rect 26 1485 1314 1492
rect 26 1436 125 1485
rect 26 1402 60 1436
rect 94 1402 125 1436
rect 1215 1436 1314 1485
rect 26 1346 125 1402
rect 26 1312 60 1346
rect 94 1312 125 1346
rect 26 1256 125 1312
rect 26 1222 60 1256
rect 94 1222 125 1256
rect 26 1166 125 1222
rect 26 1132 60 1166
rect 94 1132 125 1166
rect 26 1076 125 1132
rect 26 1042 60 1076
rect 94 1042 125 1076
rect 26 986 125 1042
rect 26 952 60 986
rect 94 952 125 986
rect 26 896 125 952
rect 26 862 60 896
rect 94 862 125 896
rect 26 806 125 862
rect 26 772 60 806
rect 94 772 125 806
rect 26 716 125 772
rect 26 682 60 716
rect 94 682 125 716
rect 26 626 125 682
rect 26 592 60 626
rect 94 592 125 626
rect 26 536 125 592
rect 26 502 60 536
rect 94 502 125 536
rect 26 446 125 502
rect 189 1402 1151 1421
rect 189 1368 320 1402
rect 354 1368 410 1402
rect 444 1368 500 1402
rect 534 1368 590 1402
rect 624 1368 680 1402
rect 714 1368 770 1402
rect 804 1368 860 1402
rect 894 1368 950 1402
rect 984 1368 1040 1402
rect 1074 1368 1151 1402
rect 189 1349 1151 1368
rect 189 1345 261 1349
rect 189 1311 208 1345
rect 242 1311 261 1345
rect 189 1255 261 1311
rect 1079 1326 1151 1349
rect 1079 1292 1098 1326
rect 1132 1292 1151 1326
rect 189 1221 208 1255
rect 242 1221 261 1255
rect 189 1165 261 1221
rect 189 1131 208 1165
rect 242 1131 261 1165
rect 189 1075 261 1131
rect 189 1041 208 1075
rect 242 1041 261 1075
rect 189 985 261 1041
rect 189 951 208 985
rect 242 951 261 985
rect 189 895 261 951
rect 189 861 208 895
rect 242 861 261 895
rect 189 805 261 861
rect 189 771 208 805
rect 242 771 261 805
rect 189 715 261 771
rect 189 681 208 715
rect 242 681 261 715
rect 189 625 261 681
rect 189 591 208 625
rect 242 591 261 625
rect 323 1228 1017 1287
rect 323 1194 384 1228
rect 418 1200 474 1228
rect 508 1200 564 1228
rect 598 1200 654 1228
rect 430 1194 474 1200
rect 530 1194 564 1200
rect 630 1194 654 1200
rect 688 1200 744 1228
rect 688 1194 696 1200
rect 323 1166 396 1194
rect 430 1166 496 1194
rect 530 1166 596 1194
rect 630 1166 696 1194
rect 730 1194 744 1200
rect 778 1200 834 1228
rect 778 1194 796 1200
rect 730 1166 796 1194
rect 830 1194 834 1200
rect 868 1200 924 1228
rect 868 1194 896 1200
rect 958 1194 1017 1228
rect 830 1166 896 1194
rect 930 1166 1017 1194
rect 323 1138 1017 1166
rect 323 1104 384 1138
rect 418 1104 474 1138
rect 508 1104 564 1138
rect 598 1104 654 1138
rect 688 1104 744 1138
rect 778 1104 834 1138
rect 868 1104 924 1138
rect 958 1104 1017 1138
rect 323 1100 1017 1104
rect 323 1066 396 1100
rect 430 1066 496 1100
rect 530 1066 596 1100
rect 630 1066 696 1100
rect 730 1066 796 1100
rect 830 1066 896 1100
rect 930 1066 1017 1100
rect 323 1048 1017 1066
rect 323 1014 384 1048
rect 418 1014 474 1048
rect 508 1014 564 1048
rect 598 1014 654 1048
rect 688 1014 744 1048
rect 778 1014 834 1048
rect 868 1014 924 1048
rect 958 1014 1017 1048
rect 323 1000 1017 1014
rect 323 966 396 1000
rect 430 966 496 1000
rect 530 966 596 1000
rect 630 966 696 1000
rect 730 966 796 1000
rect 830 966 896 1000
rect 930 966 1017 1000
rect 323 958 1017 966
rect 323 924 384 958
rect 418 924 474 958
rect 508 924 564 958
rect 598 924 654 958
rect 688 924 744 958
rect 778 924 834 958
rect 868 924 924 958
rect 958 924 1017 958
rect 323 900 1017 924
rect 323 868 396 900
rect 430 868 496 900
rect 530 868 596 900
rect 630 868 696 900
rect 323 834 384 868
rect 430 866 474 868
rect 530 866 564 868
rect 630 866 654 868
rect 418 834 474 866
rect 508 834 564 866
rect 598 834 654 866
rect 688 866 696 868
rect 730 868 796 900
rect 730 866 744 868
rect 688 834 744 866
rect 778 866 796 868
rect 830 868 896 900
rect 930 868 1017 900
rect 830 866 834 868
rect 778 834 834 866
rect 868 866 896 868
rect 868 834 924 866
rect 958 834 1017 868
rect 323 800 1017 834
rect 323 778 396 800
rect 430 778 496 800
rect 530 778 596 800
rect 630 778 696 800
rect 323 744 384 778
rect 430 766 474 778
rect 530 766 564 778
rect 630 766 654 778
rect 418 744 474 766
rect 508 744 564 766
rect 598 744 654 766
rect 688 766 696 778
rect 730 778 796 800
rect 730 766 744 778
rect 688 744 744 766
rect 778 766 796 778
rect 830 778 896 800
rect 930 778 1017 800
rect 830 766 834 778
rect 778 744 834 766
rect 868 766 896 778
rect 868 744 924 766
rect 958 744 1017 778
rect 323 700 1017 744
rect 323 688 396 700
rect 430 688 496 700
rect 530 688 596 700
rect 630 688 696 700
rect 323 654 384 688
rect 430 666 474 688
rect 530 666 564 688
rect 630 666 654 688
rect 418 654 474 666
rect 508 654 564 666
rect 598 654 654 666
rect 688 666 696 688
rect 730 688 796 700
rect 730 666 744 688
rect 688 654 744 666
rect 778 666 796 688
rect 830 688 896 700
rect 930 688 1017 700
rect 830 666 834 688
rect 778 654 834 666
rect 868 666 896 688
rect 868 654 924 666
rect 958 654 1017 688
rect 323 593 1017 654
rect 1079 1236 1151 1292
rect 1079 1202 1098 1236
rect 1132 1202 1151 1236
rect 1079 1146 1151 1202
rect 1079 1112 1098 1146
rect 1132 1112 1151 1146
rect 1079 1056 1151 1112
rect 1079 1022 1098 1056
rect 1132 1022 1151 1056
rect 1079 966 1151 1022
rect 1079 932 1098 966
rect 1132 932 1151 966
rect 1079 876 1151 932
rect 1079 842 1098 876
rect 1132 842 1151 876
rect 1079 786 1151 842
rect 1079 752 1098 786
rect 1132 752 1151 786
rect 1079 696 1151 752
rect 1079 662 1098 696
rect 1132 662 1151 696
rect 1079 606 1151 662
rect 189 531 261 591
rect 1079 572 1098 606
rect 1132 572 1151 606
rect 1079 531 1151 572
rect 189 512 1151 531
rect 189 478 286 512
rect 320 478 376 512
rect 410 478 466 512
rect 500 478 556 512
rect 590 478 646 512
rect 680 478 736 512
rect 770 478 826 512
rect 860 478 916 512
rect 950 478 1006 512
rect 1040 478 1151 512
rect 189 459 1151 478
rect 1215 1402 1247 1436
rect 1281 1402 1314 1436
rect 1215 1346 1314 1402
rect 1215 1312 1247 1346
rect 1281 1312 1314 1346
rect 1215 1256 1314 1312
rect 1215 1222 1247 1256
rect 1281 1222 1314 1256
rect 1215 1166 1314 1222
rect 1215 1132 1247 1166
rect 1281 1132 1314 1166
rect 1215 1076 1314 1132
rect 1215 1042 1247 1076
rect 1281 1042 1314 1076
rect 1215 986 1314 1042
rect 1215 952 1247 986
rect 1281 952 1314 986
rect 1215 896 1314 952
rect 1215 862 1247 896
rect 1281 862 1314 896
rect 1215 806 1314 862
rect 1215 772 1247 806
rect 1281 772 1314 806
rect 1215 716 1314 772
rect 1215 682 1247 716
rect 1281 682 1314 716
rect 1215 626 1314 682
rect 1215 592 1247 626
rect 1281 592 1314 626
rect 1215 536 1314 592
rect 1215 502 1247 536
rect 1281 502 1314 536
rect 26 412 60 446
rect 94 412 125 446
rect 26 395 125 412
rect 1215 446 1314 502
rect 1215 412 1247 446
rect 1281 412 1314 446
rect 1215 395 1314 412
rect 26 362 1314 395
rect 26 328 156 362
rect 190 328 246 362
rect 280 328 336 362
rect 370 328 426 362
rect 460 328 516 362
rect 550 328 606 362
rect 640 328 696 362
rect 730 328 786 362
rect 820 328 876 362
rect 910 328 966 362
rect 1000 328 1056 362
rect 1090 328 1146 362
rect 1180 328 1314 362
rect 26 296 1314 328
rect 0 -30 170 30
rect 230 -30 370 30
rect 430 -30 570 30
rect 630 -30 770 30
rect 830 -30 970 30
rect 1030 -30 1170 30
rect 1230 -30 1340 30
<< viali >>
rect 170 1850 230 1910
rect 370 1850 430 1910
rect 570 1850 630 1910
rect 770 1850 830 1910
rect 970 1850 1030 1910
rect 1170 1850 1230 1910
rect 396 1194 418 1200
rect 418 1194 430 1200
rect 496 1194 508 1200
rect 508 1194 530 1200
rect 596 1194 598 1200
rect 598 1194 630 1200
rect 396 1166 430 1194
rect 496 1166 530 1194
rect 596 1166 630 1194
rect 696 1166 730 1200
rect 796 1166 830 1200
rect 896 1194 924 1200
rect 924 1194 930 1200
rect 896 1166 930 1194
rect 396 1066 430 1100
rect 496 1066 530 1100
rect 596 1066 630 1100
rect 696 1066 730 1100
rect 796 1066 830 1100
rect 896 1066 930 1100
rect 396 966 430 1000
rect 496 966 530 1000
rect 596 966 630 1000
rect 696 966 730 1000
rect 796 966 830 1000
rect 896 966 930 1000
rect 396 868 430 900
rect 496 868 530 900
rect 596 868 630 900
rect 396 866 418 868
rect 418 866 430 868
rect 496 866 508 868
rect 508 866 530 868
rect 596 866 598 868
rect 598 866 630 868
rect 696 866 730 900
rect 796 866 830 900
rect 896 868 930 900
rect 896 866 924 868
rect 924 866 930 868
rect 396 778 430 800
rect 496 778 530 800
rect 596 778 630 800
rect 396 766 418 778
rect 418 766 430 778
rect 496 766 508 778
rect 508 766 530 778
rect 596 766 598 778
rect 598 766 630 778
rect 696 766 730 800
rect 796 766 830 800
rect 896 778 930 800
rect 896 766 924 778
rect 924 766 930 778
rect 396 688 430 700
rect 496 688 530 700
rect 596 688 630 700
rect 396 666 418 688
rect 418 666 430 688
rect 496 666 508 688
rect 508 666 530 688
rect 596 666 598 688
rect 598 666 630 688
rect 696 666 730 700
rect 796 666 830 700
rect 896 688 930 700
rect 896 666 924 688
rect 924 666 930 688
rect 170 -30 230 30
rect 370 -30 430 30
rect 570 -30 630 30
rect 770 -30 830 30
rect 970 -30 1030 30
rect 1170 -30 1230 30
<< metal1 >>
rect 0 1910 1340 1940
rect 0 1850 170 1910
rect 230 1850 370 1910
rect 430 1850 570 1910
rect 630 1850 770 1910
rect 830 1850 970 1910
rect 1030 1850 1170 1910
rect 1230 1850 1340 1910
rect 0 1820 1340 1850
rect 365 1200 975 1245
rect 365 1166 396 1200
rect 430 1166 496 1200
rect 530 1166 596 1200
rect 630 1166 696 1200
rect 730 1166 796 1200
rect 830 1166 896 1200
rect 930 1166 975 1200
rect 365 1100 975 1166
rect 365 1066 396 1100
rect 430 1066 496 1100
rect 530 1066 596 1100
rect 630 1066 696 1100
rect 730 1066 796 1100
rect 830 1066 896 1100
rect 930 1066 975 1100
rect 365 1000 975 1066
rect 365 966 396 1000
rect 430 966 496 1000
rect 530 966 596 1000
rect 630 966 696 1000
rect 730 966 796 1000
rect 830 966 896 1000
rect 930 966 975 1000
rect 365 900 975 966
rect 365 866 396 900
rect 430 866 496 900
rect 530 866 596 900
rect 630 866 696 900
rect 730 866 796 900
rect 830 866 896 900
rect 930 866 975 900
rect 365 800 975 866
rect 365 766 396 800
rect 430 766 496 800
rect 530 766 596 800
rect 630 766 696 800
rect 730 766 796 800
rect 830 766 896 800
rect 930 766 975 800
rect 365 700 975 766
rect 365 666 396 700
rect 430 666 496 700
rect 530 666 596 700
rect 630 666 696 700
rect 730 666 796 700
rect 830 666 896 700
rect 930 666 975 700
rect 365 635 975 666
rect 0 30 1340 60
rect 0 -30 170 30
rect 230 -30 370 30
rect 430 -30 570 30
rect 630 -30 770 30
rect 830 -30 970 30
rect 1030 -30 1170 30
rect 1230 -30 1340 30
rect 0 -60 1340 -30
<< pnp3p40 >>
rect 153 423 1187 1457
<< labels >>
flabel locali 810 1524 930 1564 1 FreeSans 480 0 0 0 Collector
port 3 n default bidirectional
flabel locali 774 1372 894 1412 1 FreeSans 480 0 0 0 Base
port 2 n default bidirectional
flabel locali 562 1010 790 1140 1 FreeSans 480 0 0 0 Emitter
port 1 n default bidirectional
flabel metal1 0 1850 60 1910 1 FreeSans 800 0 0 0 VPWR
port 4 n power bidirectional
flabel metal1 0 -30 60 30 1 FreeSans 800 0 0 0 VGND
port 5 n ground bidirectional
flabel locali 554 896 802 1000 0 FreeSans 400 0 0 0 xm1/Emitter
flabel locali 613 1522 714 1571 0 FreeSans 400 0 0 0 xm1/Collector
flabel locali 590 1372 708 1412 0 FreeSans 400 0 0 0 xm1/Base
<< properties >>
string FIXED_BBOX 0 0 1340 1880
string LEFclass CORE
string LEFsite unitasc
<< end >>
