VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO sky130_asc_pfet_01v8_lvt_60
  CLASS CORE ;
  FOREIGN sky130_asc_pfet_01v8_lvt_60 ;
  ORIGIN 0.000 0.000 ;
  SIZE 138.535 BY 9.400 ;
  SITE unitasc ;
  PIN GATE
    DIRECTION INOUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 774.000000 ;
    PORT
      LAYER li1 ;
        RECT 0.490 0.520 138.530 0.820 ;
    END
  END GATE
  PIN SOURCE
    DIRECTION INOUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 56.114998 ;
    PORT
      LAYER li1 ;
        RECT 0.790 8.650 138.530 8.950 ;
        RECT 3.015 1.755 3.185 8.650 ;
        RECT 7.595 1.755 7.765 8.650 ;
        RECT 12.175 1.755 12.345 8.650 ;
        RECT 16.755 1.755 16.925 8.650 ;
        RECT 21.335 1.755 21.505 8.650 ;
        RECT 25.915 1.755 26.085 8.650 ;
        RECT 30.495 1.755 30.665 8.650 ;
        RECT 35.075 1.755 35.245 8.650 ;
        RECT 39.655 1.755 39.825 8.650 ;
        RECT 44.235 1.755 44.405 8.650 ;
        RECT 48.815 1.755 48.985 8.650 ;
        RECT 53.395 1.755 53.565 8.650 ;
        RECT 57.975 1.755 58.145 8.650 ;
        RECT 62.555 1.755 62.725 8.650 ;
        RECT 67.135 1.755 67.305 8.650 ;
        RECT 71.715 1.755 71.885 8.650 ;
        RECT 76.295 1.755 76.465 8.650 ;
        RECT 80.875 1.755 81.045 8.650 ;
        RECT 85.455 1.755 85.625 8.650 ;
        RECT 90.035 1.755 90.205 8.650 ;
        RECT 94.615 1.755 94.785 8.650 ;
        RECT 99.195 1.755 99.365 8.650 ;
        RECT 103.775 1.755 103.945 8.650 ;
        RECT 108.355 1.755 108.525 8.650 ;
        RECT 112.935 1.755 113.105 8.650 ;
        RECT 117.515 1.755 117.685 8.650 ;
        RECT 122.095 1.755 122.265 8.650 ;
        RECT 126.675 1.755 126.845 8.650 ;
        RECT 131.255 1.755 131.425 8.650 ;
        RECT 135.835 1.755 136.005 8.650 ;
      LAYER mcon ;
        RECT 3.015 1.835 3.185 8.165 ;
        RECT 7.595 1.835 7.765 8.165 ;
        RECT 12.175 1.835 12.345 8.165 ;
        RECT 16.755 1.835 16.925 8.165 ;
        RECT 21.335 1.835 21.505 8.165 ;
        RECT 25.915 1.835 26.085 8.165 ;
        RECT 30.495 1.835 30.665 8.165 ;
        RECT 35.075 1.835 35.245 8.165 ;
        RECT 39.655 1.835 39.825 8.165 ;
        RECT 44.235 1.835 44.405 8.165 ;
        RECT 48.815 1.835 48.985 8.165 ;
        RECT 53.395 1.835 53.565 8.165 ;
        RECT 57.975 1.835 58.145 8.165 ;
        RECT 62.555 1.835 62.725 8.165 ;
        RECT 67.135 1.835 67.305 8.165 ;
        RECT 71.715 1.835 71.885 8.165 ;
        RECT 76.295 1.835 76.465 8.165 ;
        RECT 80.875 1.835 81.045 8.165 ;
        RECT 85.455 1.835 85.625 8.165 ;
        RECT 90.035 1.835 90.205 8.165 ;
        RECT 94.615 1.835 94.785 8.165 ;
        RECT 99.195 1.835 99.365 8.165 ;
        RECT 103.775 1.835 103.945 8.165 ;
        RECT 108.355 1.835 108.525 8.165 ;
        RECT 112.935 1.835 113.105 8.165 ;
        RECT 117.515 1.835 117.685 8.165 ;
        RECT 122.095 1.835 122.265 8.165 ;
        RECT 126.675 1.835 126.845 8.165 ;
        RECT 131.255 1.835 131.425 8.165 ;
        RECT 135.835 1.835 136.005 8.165 ;
      LAYER met1 ;
        RECT 2.985 1.775 3.215 8.225 ;
        RECT 7.565 1.775 7.795 8.225 ;
        RECT 12.145 1.775 12.375 8.225 ;
        RECT 16.725 1.775 16.955 8.225 ;
        RECT 21.305 1.775 21.535 8.225 ;
        RECT 25.885 1.775 26.115 8.225 ;
        RECT 30.465 1.775 30.695 8.225 ;
        RECT 35.045 1.775 35.275 8.225 ;
        RECT 39.625 1.775 39.855 8.225 ;
        RECT 44.205 1.775 44.435 8.225 ;
        RECT 48.785 1.775 49.015 8.225 ;
        RECT 53.365 1.775 53.595 8.225 ;
        RECT 57.945 1.775 58.175 8.225 ;
        RECT 62.525 1.775 62.755 8.225 ;
        RECT 67.105 1.775 67.335 8.225 ;
        RECT 71.685 1.775 71.915 8.225 ;
        RECT 76.265 1.775 76.495 8.225 ;
        RECT 80.845 1.775 81.075 8.225 ;
        RECT 85.425 1.775 85.655 8.225 ;
        RECT 90.005 1.775 90.235 8.225 ;
        RECT 94.585 1.775 94.815 8.225 ;
        RECT 99.165 1.775 99.395 8.225 ;
        RECT 103.745 1.775 103.975 8.225 ;
        RECT 108.325 1.775 108.555 8.225 ;
        RECT 112.905 1.775 113.135 8.225 ;
        RECT 117.485 1.775 117.715 8.225 ;
        RECT 122.065 1.775 122.295 8.225 ;
        RECT 126.645 1.775 126.875 8.225 ;
        RECT 131.225 1.775 131.455 8.225 ;
        RECT 135.805 1.775 136.035 8.225 ;
    END
  END SOURCE
  PIN DRAIN
    DIRECTION INOUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 57.985500 ;
    PORT
      LAYER li1 ;
        RECT 0.725 1.350 0.895 8.245 ;
        RECT 5.305 1.350 5.475 8.245 ;
        RECT 9.885 1.350 10.055 8.245 ;
        RECT 14.465 1.350 14.635 8.245 ;
        RECT 19.045 1.350 19.215 8.245 ;
        RECT 23.625 1.350 23.795 8.245 ;
        RECT 28.205 1.350 28.375 8.245 ;
        RECT 32.785 1.350 32.955 8.245 ;
        RECT 37.365 1.350 37.535 8.245 ;
        RECT 41.945 1.350 42.115 8.245 ;
        RECT 46.525 1.350 46.695 8.245 ;
        RECT 51.105 1.350 51.275 8.245 ;
        RECT 55.685 1.350 55.855 8.245 ;
        RECT 60.265 1.350 60.435 8.245 ;
        RECT 64.845 1.350 65.015 8.245 ;
        RECT 69.425 1.350 69.595 8.245 ;
        RECT 74.005 1.350 74.175 8.245 ;
        RECT 78.585 1.350 78.755 8.245 ;
        RECT 83.165 1.350 83.335 8.245 ;
        RECT 87.745 1.350 87.915 8.245 ;
        RECT 92.325 1.350 92.495 8.245 ;
        RECT 96.905 1.350 97.075 8.245 ;
        RECT 101.485 1.350 101.655 8.245 ;
        RECT 106.065 1.350 106.235 8.245 ;
        RECT 110.645 1.350 110.815 8.245 ;
        RECT 115.225 1.350 115.395 8.245 ;
        RECT 119.805 1.350 119.975 8.245 ;
        RECT 124.385 1.350 124.555 8.245 ;
        RECT 128.965 1.350 129.135 8.245 ;
        RECT 133.545 1.350 133.715 8.245 ;
        RECT 138.125 1.350 138.295 8.245 ;
        RECT 0.490 1.050 138.530 1.350 ;
      LAYER mcon ;
        RECT 0.725 1.835 0.895 8.165 ;
        RECT 5.305 1.835 5.475 8.165 ;
        RECT 9.885 1.835 10.055 8.165 ;
        RECT 14.465 1.835 14.635 8.165 ;
        RECT 19.045 1.835 19.215 8.165 ;
        RECT 23.625 1.835 23.795 8.165 ;
        RECT 28.205 1.835 28.375 8.165 ;
        RECT 32.785 1.835 32.955 8.165 ;
        RECT 37.365 1.835 37.535 8.165 ;
        RECT 41.945 1.835 42.115 8.165 ;
        RECT 46.525 1.835 46.695 8.165 ;
        RECT 51.105 1.835 51.275 8.165 ;
        RECT 55.685 1.835 55.855 8.165 ;
        RECT 60.265 1.835 60.435 8.165 ;
        RECT 64.845 1.835 65.015 8.165 ;
        RECT 69.425 1.835 69.595 8.165 ;
        RECT 74.005 1.835 74.175 8.165 ;
        RECT 78.585 1.835 78.755 8.165 ;
        RECT 83.165 1.835 83.335 8.165 ;
        RECT 87.745 1.835 87.915 8.165 ;
        RECT 92.325 1.835 92.495 8.165 ;
        RECT 96.905 1.835 97.075 8.165 ;
        RECT 101.485 1.835 101.655 8.165 ;
        RECT 106.065 1.835 106.235 8.165 ;
        RECT 110.645 1.835 110.815 8.165 ;
        RECT 115.225 1.835 115.395 8.165 ;
        RECT 119.805 1.835 119.975 8.165 ;
        RECT 124.385 1.835 124.555 8.165 ;
        RECT 128.965 1.835 129.135 8.165 ;
        RECT 133.545 1.835 133.715 8.165 ;
        RECT 138.125 1.835 138.295 8.165 ;
      LAYER met1 ;
        RECT 0.695 1.775 0.925 8.225 ;
        RECT 5.275 1.775 5.505 8.225 ;
        RECT 9.855 1.775 10.085 8.225 ;
        RECT 14.435 1.775 14.665 8.225 ;
        RECT 19.015 1.775 19.245 8.225 ;
        RECT 23.595 1.775 23.825 8.225 ;
        RECT 28.175 1.775 28.405 8.225 ;
        RECT 32.755 1.775 32.985 8.225 ;
        RECT 37.335 1.775 37.565 8.225 ;
        RECT 41.915 1.775 42.145 8.225 ;
        RECT 46.495 1.775 46.725 8.225 ;
        RECT 51.075 1.775 51.305 8.225 ;
        RECT 55.655 1.775 55.885 8.225 ;
        RECT 60.235 1.775 60.465 8.225 ;
        RECT 64.815 1.775 65.045 8.225 ;
        RECT 69.395 1.775 69.625 8.225 ;
        RECT 73.975 1.775 74.205 8.225 ;
        RECT 78.555 1.775 78.785 8.225 ;
        RECT 83.135 1.775 83.365 8.225 ;
        RECT 87.715 1.775 87.945 8.225 ;
        RECT 92.295 1.775 92.525 8.225 ;
        RECT 96.875 1.775 97.105 8.225 ;
        RECT 101.455 1.775 101.685 8.225 ;
        RECT 106.035 1.775 106.265 8.225 ;
        RECT 110.615 1.775 110.845 8.225 ;
        RECT 115.195 1.775 115.425 8.225 ;
        RECT 119.775 1.775 120.005 8.225 ;
        RECT 124.355 1.775 124.585 8.225 ;
        RECT 128.935 1.775 129.165 8.225 ;
        RECT 133.515 1.775 133.745 8.225 ;
        RECT 138.095 1.775 138.325 8.225 ;
    END
  END DRAIN
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT 0.000 8.535 138.530 9.700 ;
        RECT 0.000 1.470 138.535 8.535 ;
        RECT 0.485 1.465 138.535 1.470 ;
      LAYER li1 ;
        RECT 0.000 9.250 138.530 9.550 ;
        RECT 0.140 8.200 0.440 9.250 ;
      LAYER mcon ;
        RECT 1.340 9.250 1.640 9.550 ;
        RECT 3.340 9.250 3.640 9.550 ;
        RECT 5.340 9.250 5.640 9.550 ;
        RECT 7.340 9.250 7.640 9.550 ;
        RECT 9.340 9.250 9.640 9.550 ;
        RECT 11.340 9.250 11.640 9.550 ;
        RECT 13.340 9.250 13.640 9.550 ;
        RECT 15.340 9.250 15.640 9.550 ;
        RECT 17.340 9.250 17.640 9.550 ;
        RECT 19.340 9.250 19.640 9.550 ;
        RECT 21.340 9.250 21.640 9.550 ;
        RECT 23.340 9.250 23.640 9.550 ;
        RECT 25.340 9.250 25.640 9.550 ;
        RECT 27.340 9.250 27.640 9.550 ;
        RECT 29.340 9.250 29.640 9.550 ;
        RECT 31.340 9.250 31.640 9.550 ;
        RECT 33.340 9.250 33.640 9.550 ;
        RECT 35.340 9.250 35.640 9.550 ;
        RECT 37.340 9.250 37.640 9.550 ;
        RECT 39.340 9.250 39.640 9.550 ;
        RECT 41.340 9.250 41.640 9.550 ;
        RECT 43.340 9.250 43.640 9.550 ;
        RECT 45.340 9.250 45.640 9.550 ;
        RECT 47.340 9.250 47.640 9.550 ;
        RECT 49.340 9.250 49.640 9.550 ;
        RECT 51.340 9.250 51.640 9.550 ;
        RECT 53.340 9.250 53.640 9.550 ;
        RECT 55.340 9.250 55.640 9.550 ;
        RECT 57.340 9.250 57.640 9.550 ;
        RECT 59.340 9.250 59.640 9.550 ;
        RECT 61.340 9.250 61.640 9.550 ;
        RECT 63.340 9.250 63.640 9.550 ;
        RECT 65.340 9.250 65.640 9.550 ;
        RECT 67.340 9.250 67.640 9.550 ;
        RECT 69.340 9.250 69.640 9.550 ;
        RECT 71.340 9.250 71.640 9.550 ;
        RECT 73.340 9.250 73.640 9.550 ;
        RECT 75.340 9.250 75.640 9.550 ;
        RECT 77.340 9.250 77.640 9.550 ;
        RECT 79.340 9.250 79.640 9.550 ;
        RECT 81.340 9.250 81.640 9.550 ;
        RECT 83.340 9.250 83.640 9.550 ;
        RECT 85.340 9.250 85.640 9.550 ;
        RECT 87.340 9.250 87.640 9.550 ;
        RECT 89.340 9.250 89.640 9.550 ;
        RECT 91.340 9.250 91.640 9.550 ;
        RECT 93.340 9.250 93.640 9.550 ;
        RECT 95.340 9.250 95.640 9.550 ;
        RECT 97.340 9.250 97.640 9.550 ;
        RECT 99.340 9.250 99.640 9.550 ;
        RECT 101.340 9.250 101.640 9.550 ;
        RECT 103.340 9.250 103.640 9.550 ;
        RECT 105.340 9.250 105.640 9.550 ;
        RECT 107.340 9.250 107.640 9.550 ;
        RECT 109.340 9.250 109.640 9.550 ;
        RECT 111.340 9.250 111.640 9.550 ;
        RECT 113.340 9.250 113.640 9.550 ;
        RECT 115.340 9.250 115.640 9.550 ;
        RECT 117.340 9.250 117.640 9.550 ;
        RECT 119.340 9.250 119.640 9.550 ;
        RECT 121.340 9.250 121.640 9.550 ;
        RECT 123.340 9.250 123.640 9.550 ;
        RECT 125.340 9.250 125.640 9.550 ;
        RECT 127.340 9.250 127.640 9.550 ;
        RECT 129.340 9.250 129.640 9.550 ;
        RECT 131.340 9.250 131.640 9.550 ;
        RECT 133.340 9.250 133.640 9.550 ;
        RECT 135.340 9.250 135.640 9.550 ;
        RECT 137.340 9.250 137.640 9.550 ;
      LAYER met1 ;
        RECT 0.000 9.100 138.530 9.700 ;
    END
  END VPWR
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER li1 ;
        RECT 0.000 -0.150 138.530 0.150 ;
      LAYER mcon ;
        RECT 1.340 -0.150 1.640 0.150 ;
        RECT 3.340 -0.150 3.640 0.150 ;
        RECT 5.340 -0.150 5.640 0.150 ;
        RECT 7.340 -0.150 7.640 0.150 ;
        RECT 9.340 -0.150 9.640 0.150 ;
        RECT 11.340 -0.150 11.640 0.150 ;
        RECT 13.340 -0.150 13.640 0.150 ;
        RECT 15.340 -0.150 15.640 0.150 ;
        RECT 17.340 -0.150 17.640 0.150 ;
        RECT 19.340 -0.150 19.640 0.150 ;
        RECT 21.340 -0.150 21.640 0.150 ;
        RECT 23.340 -0.150 23.640 0.150 ;
        RECT 25.340 -0.150 25.640 0.150 ;
        RECT 27.340 -0.150 27.640 0.150 ;
        RECT 29.340 -0.150 29.640 0.150 ;
        RECT 31.340 -0.150 31.640 0.150 ;
        RECT 33.340 -0.150 33.640 0.150 ;
        RECT 35.340 -0.150 35.640 0.150 ;
        RECT 37.340 -0.150 37.640 0.150 ;
        RECT 39.340 -0.150 39.640 0.150 ;
        RECT 41.340 -0.150 41.640 0.150 ;
        RECT 43.340 -0.150 43.640 0.150 ;
        RECT 45.340 -0.150 45.640 0.150 ;
        RECT 47.340 -0.150 47.640 0.150 ;
        RECT 49.340 -0.150 49.640 0.150 ;
        RECT 51.340 -0.150 51.640 0.150 ;
        RECT 53.340 -0.150 53.640 0.150 ;
        RECT 55.340 -0.150 55.640 0.150 ;
        RECT 57.340 -0.150 57.640 0.150 ;
        RECT 59.340 -0.150 59.640 0.150 ;
        RECT 61.340 -0.150 61.640 0.150 ;
        RECT 63.340 -0.150 63.640 0.150 ;
        RECT 65.340 -0.150 65.640 0.150 ;
        RECT 67.340 -0.150 67.640 0.150 ;
        RECT 69.340 -0.150 69.640 0.150 ;
        RECT 71.340 -0.150 71.640 0.150 ;
        RECT 73.340 -0.150 73.640 0.150 ;
        RECT 75.340 -0.150 75.640 0.150 ;
        RECT 77.340 -0.150 77.640 0.150 ;
        RECT 79.340 -0.150 79.640 0.150 ;
        RECT 81.340 -0.150 81.640 0.150 ;
        RECT 83.340 -0.150 83.640 0.150 ;
        RECT 85.340 -0.150 85.640 0.150 ;
        RECT 87.340 -0.150 87.640 0.150 ;
        RECT 89.340 -0.150 89.640 0.150 ;
        RECT 91.340 -0.150 91.640 0.150 ;
        RECT 93.340 -0.150 93.640 0.150 ;
        RECT 95.340 -0.150 95.640 0.150 ;
        RECT 97.340 -0.150 97.640 0.150 ;
        RECT 99.340 -0.150 99.640 0.150 ;
        RECT 101.340 -0.150 101.640 0.150 ;
        RECT 103.340 -0.150 103.640 0.150 ;
        RECT 105.340 -0.150 105.640 0.150 ;
        RECT 107.340 -0.150 107.640 0.150 ;
        RECT 109.340 -0.150 109.640 0.150 ;
        RECT 111.340 -0.150 111.640 0.150 ;
        RECT 113.340 -0.150 113.640 0.150 ;
        RECT 115.340 -0.150 115.640 0.150 ;
        RECT 117.340 -0.150 117.640 0.150 ;
        RECT 119.340 -0.150 119.640 0.150 ;
        RECT 121.340 -0.150 121.640 0.150 ;
        RECT 123.340 -0.150 123.640 0.150 ;
        RECT 125.340 -0.150 125.640 0.150 ;
        RECT 127.340 -0.150 127.640 0.150 ;
        RECT 129.340 -0.150 129.640 0.150 ;
        RECT 131.340 -0.150 131.640 0.150 ;
        RECT 133.340 -0.150 133.640 0.150 ;
        RECT 135.340 -0.150 135.640 0.150 ;
        RECT 137.340 -0.150 137.640 0.150 ;
      LAYER met1 ;
        RECT 0.000 -0.300 138.530 0.300 ;
    END
  END VGND
END sky130_asc_pfet_01v8_lvt_60
END LIBRARY

