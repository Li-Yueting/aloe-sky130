/home/users/xingyuni/ee372/mflowgen_flow/aloe-sky130/ringosc/build/2-skywater-130nm/view-standard/stdcells.lef