VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO sky130_asc_nfet_01v8_lvt_1
  CLASS CORE ;
  FOREIGN sky130_asc_nfet_01v8_lvt_1 ;
  ORIGIN 0.000 0.000 ;
  SIZE 2.580 BY 9.400 ;
  SITE unitasc ;
  PIN GATE
    DIRECTION INOUT ;
    ANTENNAGATEAREA 8.000000 ;
    PORT
      LAYER li1 ;
        RECT 0.000 0.720 2.580 1.020 ;
    END
  END GATE
  PIN SOURCE
    DIRECTION INOUT ;
    ANTENNADIFFAREA 1.160000 ;
    PORT
      LAYER li1 ;
        RECT 0.000 8.450 2.580 8.750 ;
        RECT 2.345 7.020 2.515 8.450 ;
        RECT 2.345 6.930 2.520 7.020 ;
        RECT 2.350 2.980 2.520 6.930 ;
      LAYER mcon ;
        RECT 2.350 3.060 2.520 6.940 ;
      LAYER met1 ;
        RECT 2.320 3.000 2.550 7.000 ;
    END
  END SOURCE
  PIN DRAIN
    DIRECTION INOUT ;
    ANTENNADIFFAREA 1.160000 ;
    PORT
      LAYER li1 ;
        RECT 0.060 3.270 0.230 7.020 ;
        RECT 0.055 2.980 0.230 3.270 ;
        RECT 0.055 2.150 0.225 2.980 ;
        RECT 0.000 1.850 2.580 2.150 ;
      LAYER mcon ;
        RECT 0.060 3.060 0.230 6.940 ;
      LAYER met1 ;
        RECT 0.030 3.000 0.260 7.000 ;
    END
  END DRAIN
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.000 0.150 2.580 5.000 ;
        RECT 2.280 -0.150 2.580 0.150 ;
    END
  END VNB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER li1 ;
        RECT 0.000 9.250 2.580 9.550 ;
      LAYER mcon ;
        RECT 0.850 9.250 1.150 9.550 ;
      LAYER met1 ;
        RECT 0.000 9.100 2.580 9.700 ;
    END
  END VPWR
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER li1 ;
        RECT 0.000 -0.150 2.580 0.150 ;
      LAYER mcon ;
        RECT 0.850 -0.150 1.150 0.150 ;
      LAYER met1 ;
        RECT 0.000 -0.300 2.580 0.300 ;
    END
  END VGND
END sky130_asc_nfet_01v8_lvt_1
END LIBRARY

