VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO sky130_asc_nfet_01v8_lvt_9
  CLASS CORE ;
  FOREIGN sky130_asc_nfet_01v8_lvt_9 ;
  ORIGIN 0.000 0.000 ;
  SIZE 22.500 BY 9.400 ;
  SITE unitasc ;
  PIN GATE
    DIRECTION INOUT ;
    ANTENNAGATEAREA 72.000000 ;
    PORT
      LAYER li1 ;
        RECT 1.340 0.720 21.840 1.020 ;
    END
  END GATE
  PIN SOURCE
    DIRECTION INOUT ;
    ANTENNADIFFAREA 5.800000 ;
    PORT
      LAYER li1 ;
        RECT 0.940 8.450 21.840 8.750 ;
        RECT 3.285 7.020 3.455 8.450 ;
        RECT 7.865 7.020 8.035 8.450 ;
        RECT 12.445 7.020 12.615 8.450 ;
        RECT 17.025 7.020 17.195 8.450 ;
        RECT 21.605 7.020 21.775 8.450 ;
        RECT 3.285 6.930 3.460 7.020 ;
        RECT 7.865 6.930 8.040 7.020 ;
        RECT 12.445 6.930 12.620 7.020 ;
        RECT 17.025 6.930 17.200 7.020 ;
        RECT 21.605 6.930 21.780 7.020 ;
        RECT 3.290 2.980 3.460 6.930 ;
        RECT 7.870 2.980 8.040 6.930 ;
        RECT 12.450 2.980 12.620 6.930 ;
        RECT 17.030 2.980 17.200 6.930 ;
        RECT 21.610 2.980 21.780 6.930 ;
      LAYER mcon ;
        RECT 3.290 3.060 3.460 6.940 ;
        RECT 7.870 3.060 8.040 6.940 ;
        RECT 12.450 3.060 12.620 6.940 ;
        RECT 17.030 3.060 17.200 6.940 ;
        RECT 21.610 3.060 21.780 6.940 ;
      LAYER met1 ;
        RECT 3.260 3.000 3.490 7.000 ;
        RECT 7.840 3.000 8.070 7.000 ;
        RECT 12.420 3.000 12.650 7.000 ;
        RECT 17.000 3.000 17.230 7.000 ;
        RECT 21.580 3.000 21.810 7.000 ;
    END
  END SOURCE
  PIN DRAIN
    DIRECTION INOUT ;
    ANTENNADIFFAREA 5.800000 ;
    PORT
      LAYER li1 ;
        RECT 1.000 3.270 1.170 7.020 ;
        RECT 5.580 3.270 5.750 7.020 ;
        RECT 10.160 3.270 10.330 7.020 ;
        RECT 14.740 3.270 14.910 7.020 ;
        RECT 19.320 3.270 19.490 7.020 ;
        RECT 0.995 2.980 1.170 3.270 ;
        RECT 5.575 2.980 5.750 3.270 ;
        RECT 10.155 2.980 10.330 3.270 ;
        RECT 14.735 2.980 14.910 3.270 ;
        RECT 19.315 2.980 19.490 3.270 ;
        RECT 0.995 2.150 1.165 2.980 ;
        RECT 5.575 2.150 5.745 2.980 ;
        RECT 10.155 2.150 10.325 2.980 ;
        RECT 14.735 2.150 14.905 2.980 ;
        RECT 19.315 2.150 19.485 2.980 ;
        RECT 0.940 1.850 21.840 2.150 ;
      LAYER mcon ;
        RECT 1.000 3.060 1.170 6.940 ;
        RECT 5.580 3.060 5.750 6.940 ;
        RECT 10.160 3.060 10.330 6.940 ;
        RECT 14.740 3.060 14.910 6.940 ;
        RECT 19.320 3.060 19.490 6.940 ;
      LAYER met1 ;
        RECT 0.970 3.000 1.200 7.000 ;
        RECT 5.550 3.000 5.780 7.000 ;
        RECT 10.130 3.000 10.360 7.000 ;
        RECT 14.710 3.000 14.940 7.000 ;
        RECT 19.290 3.000 19.520 7.000 ;
    END
  END DRAIN
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER li1 ;
        RECT 0.450 9.250 21.840 9.550 ;
      LAYER mcon ;
        RECT 1.790 9.250 2.090 9.550 ;
        RECT 3.790 9.250 4.090 9.550 ;
        RECT 5.790 9.250 6.090 9.550 ;
        RECT 7.790 9.250 8.090 9.550 ;
        RECT 9.790 9.250 10.090 9.550 ;
        RECT 11.790 9.250 12.090 9.550 ;
        RECT 13.790 9.250 14.090 9.550 ;
        RECT 15.790 9.250 16.090 9.550 ;
        RECT 17.790 9.250 18.090 9.550 ;
        RECT 19.790 9.250 20.090 9.550 ;
      LAYER met1 ;
        RECT 0.450 9.100 21.840 9.700 ;
    END
  END VPWR
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.450 0.150 21.840 7.130 ;
      LAYER li1 ;
        RECT 0.590 0.150 0.890 1.200 ;
        RECT 0.450 -0.150 21.840 0.150 ;
      LAYER mcon ;
        RECT 1.790 -0.150 2.090 0.150 ;
        RECT 3.790 -0.150 4.090 0.150 ;
        RECT 5.790 -0.150 6.090 0.150 ;
        RECT 7.790 -0.150 8.090 0.150 ;
        RECT 9.790 -0.150 10.090 0.150 ;
        RECT 11.790 -0.150 12.090 0.150 ;
        RECT 13.790 -0.150 14.090 0.150 ;
        RECT 15.790 -0.150 16.090 0.150 ;
        RECT 17.790 -0.150 18.090 0.150 ;
        RECT 19.790 -0.150 20.090 0.150 ;
      LAYER met1 ;
        RECT 0.450 -0.300 21.840 0.300 ;
    END
  END VGND
END sky130_asc_nfet_01v8_lvt_9
END LIBRARY

