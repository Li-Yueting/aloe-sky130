VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO sky130_asc_pnp_05v5_W3p40L3p40_8
  CLASS CORE ;
  FOREIGN sky130_asc_pnp_05v5_W3p40L3p40_8 ;
  ORIGIN 0.000 0.000 ;
  SIZE 54.800 BY 9.400 ;
  SITE unitasc ;
  PIN Emitter
    DIRECTION INOUT ;
    ANTENNADIFFAREA 92.479996 ;
    PORT
      LAYER met1 ;
        RECT 2.420 3.170 52.380 6.230 ;
    END
  END Emitter
  PIN Base
    DIRECTION INOUT ;
    ANTENNAGATEAREA 213.831192 ;
    ANTENNADIFFAREA 51.264000 ;
    PORT
      LAYER met1 ;
        RECT 1.550 6.750 53.250 7.100 ;
    END
  END Base
  PIN Collector
    DIRECTION INOUT ;
    ANTENNADIFFAREA 107.630394 ;
    PORT
      LAYER pwell ;
        RECT 0.600 7.285 54.200 8.050 ;
        RECT 0.600 2.115 1.365 7.285 ;
        RECT 6.535 2.115 8.065 7.285 ;
        RECT 13.235 2.115 14.765 7.285 ;
        RECT 19.935 2.115 21.465 7.285 ;
        RECT 26.635 2.115 28.165 7.285 ;
        RECT 33.335 2.115 34.865 7.285 ;
        RECT 40.035 2.115 41.565 7.285 ;
        RECT 46.735 2.115 48.265 7.285 ;
        RECT 53.435 2.115 54.200 7.285 ;
        RECT 0.600 1.350 54.200 2.115 ;
      LAYER met1 ;
        RECT 0.730 7.500 54.070 7.850 ;
    END
  END Collector
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.600 9.100 54.200 9.700 ;
    END
  END VPWR
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.600 -0.300 54.200 0.300 ;
    END
  END VGND
  OBS
      LAYER li1 ;
        RECT 0.600 9.250 54.200 9.550 ;
        RECT 0.730 7.425 54.070 7.920 ;
        RECT 0.730 1.975 1.225 7.425 ;
        RECT 1.545 6.745 6.355 7.105 ;
        RECT 1.545 2.655 1.905 6.745 ;
        RECT 2.215 2.965 5.685 6.435 ;
        RECT 5.995 2.655 6.355 6.745 ;
        RECT 1.545 2.295 6.355 2.655 ;
        RECT 6.675 1.975 7.925 7.425 ;
        RECT 8.245 6.745 13.055 7.105 ;
        RECT 8.245 2.655 8.605 6.745 ;
        RECT 8.915 2.965 12.385 6.435 ;
        RECT 12.695 2.655 13.055 6.745 ;
        RECT 8.245 2.295 13.055 2.655 ;
        RECT 13.375 1.975 14.625 7.425 ;
        RECT 14.945 6.745 19.755 7.105 ;
        RECT 14.945 2.655 15.305 6.745 ;
        RECT 15.615 2.965 19.085 6.435 ;
        RECT 19.395 2.655 19.755 6.745 ;
        RECT 14.945 2.295 19.755 2.655 ;
        RECT 20.075 1.975 21.325 7.425 ;
        RECT 21.645 6.745 26.455 7.105 ;
        RECT 21.645 2.655 22.005 6.745 ;
        RECT 22.315 2.965 25.785 6.435 ;
        RECT 26.095 2.655 26.455 6.745 ;
        RECT 21.645 2.295 26.455 2.655 ;
        RECT 26.775 1.975 28.025 7.425 ;
        RECT 28.345 6.745 33.155 7.105 ;
        RECT 28.345 2.655 28.705 6.745 ;
        RECT 29.015 2.965 32.485 6.435 ;
        RECT 32.795 2.655 33.155 6.745 ;
        RECT 28.345 2.295 33.155 2.655 ;
        RECT 33.475 1.975 34.725 7.425 ;
        RECT 35.045 6.745 39.855 7.105 ;
        RECT 35.045 2.655 35.405 6.745 ;
        RECT 35.715 2.965 39.185 6.435 ;
        RECT 39.495 2.655 39.855 6.745 ;
        RECT 35.045 2.295 39.855 2.655 ;
        RECT 40.175 1.975 41.425 7.425 ;
        RECT 41.745 6.745 46.555 7.105 ;
        RECT 41.745 2.655 42.105 6.745 ;
        RECT 42.415 2.965 45.885 6.435 ;
        RECT 46.195 2.655 46.555 6.745 ;
        RECT 41.745 2.295 46.555 2.655 ;
        RECT 46.875 1.975 48.125 7.425 ;
        RECT 48.445 6.745 53.255 7.105 ;
        RECT 48.445 2.655 48.805 6.745 ;
        RECT 49.115 2.965 52.585 6.435 ;
        RECT 52.895 2.655 53.255 6.745 ;
        RECT 48.445 2.295 53.255 2.655 ;
        RECT 53.575 1.975 54.070 7.425 ;
        RECT 0.730 1.480 54.070 1.975 ;
        RECT 0.600 -0.150 54.200 0.150 ;
      LAYER mcon ;
        RECT 1.450 9.250 1.750 9.550 ;
        RECT 2.450 9.250 2.750 9.550 ;
        RECT 3.450 9.250 3.750 9.550 ;
        RECT 4.450 9.250 4.750 9.550 ;
        RECT 5.450 9.250 5.750 9.550 ;
        RECT 6.450 9.250 6.750 9.550 ;
        RECT 7.450 9.250 7.750 9.550 ;
        RECT 8.450 9.250 8.750 9.550 ;
        RECT 9.450 9.250 9.750 9.550 ;
        RECT 10.450 9.250 10.750 9.550 ;
        RECT 11.450 9.250 11.750 9.550 ;
        RECT 12.450 9.250 12.750 9.550 ;
        RECT 13.450 9.250 13.750 9.550 ;
        RECT 14.450 9.250 14.750 9.550 ;
        RECT 15.450 9.250 15.750 9.550 ;
        RECT 16.450 9.250 16.750 9.550 ;
        RECT 17.450 9.250 17.750 9.550 ;
        RECT 18.450 9.250 18.750 9.550 ;
        RECT 19.450 9.250 19.750 9.550 ;
        RECT 20.450 9.250 20.750 9.550 ;
        RECT 21.450 9.250 21.750 9.550 ;
        RECT 22.450 9.250 22.750 9.550 ;
        RECT 23.450 9.250 23.750 9.550 ;
        RECT 24.450 9.250 24.750 9.550 ;
        RECT 25.450 9.250 25.750 9.550 ;
        RECT 26.450 9.250 26.750 9.550 ;
        RECT 27.450 9.250 27.750 9.550 ;
        RECT 28.450 9.250 28.750 9.550 ;
        RECT 29.450 9.250 29.750 9.550 ;
        RECT 30.450 9.250 30.750 9.550 ;
        RECT 31.450 9.250 31.750 9.550 ;
        RECT 32.450 9.250 32.750 9.550 ;
        RECT 33.450 9.250 33.750 9.550 ;
        RECT 34.450 9.250 34.750 9.550 ;
        RECT 35.450 9.250 35.750 9.550 ;
        RECT 36.450 9.250 36.750 9.550 ;
        RECT 37.450 9.250 37.750 9.550 ;
        RECT 38.450 9.250 38.750 9.550 ;
        RECT 39.450 9.250 39.750 9.550 ;
        RECT 40.450 9.250 40.750 9.550 ;
        RECT 41.450 9.250 41.750 9.550 ;
        RECT 42.450 9.250 42.750 9.550 ;
        RECT 43.450 9.250 43.750 9.550 ;
        RECT 44.450 9.250 44.750 9.550 ;
        RECT 45.450 9.250 45.750 9.550 ;
        RECT 46.450 9.250 46.750 9.550 ;
        RECT 47.450 9.250 47.750 9.550 ;
        RECT 48.450 9.250 48.750 9.550 ;
        RECT 49.450 9.250 49.750 9.550 ;
        RECT 50.450 9.250 50.750 9.550 ;
        RECT 51.450 9.250 51.750 9.550 ;
        RECT 52.450 9.250 52.750 9.550 ;
        RECT 53.450 9.250 53.750 9.550 ;
        RECT 0.830 7.650 1.000 7.820 ;
        RECT 1.280 7.650 1.450 7.820 ;
        RECT 1.730 7.650 1.900 7.820 ;
        RECT 2.180 7.650 2.350 7.820 ;
        RECT 2.630 7.650 2.800 7.820 ;
        RECT 3.080 7.650 3.250 7.820 ;
        RECT 3.530 7.650 3.700 7.820 ;
        RECT 3.980 7.650 4.150 7.820 ;
        RECT 4.430 7.650 4.600 7.820 ;
        RECT 4.880 7.650 5.050 7.820 ;
        RECT 5.330 7.650 5.500 7.820 ;
        RECT 5.780 7.650 5.950 7.820 ;
        RECT 6.230 7.650 6.400 7.820 ;
        RECT 6.680 7.650 6.850 7.820 ;
        RECT 7.530 7.650 7.700 7.820 ;
        RECT 7.980 7.650 8.150 7.820 ;
        RECT 8.430 7.650 8.600 7.820 ;
        RECT 8.880 7.650 9.050 7.820 ;
        RECT 9.330 7.650 9.500 7.820 ;
        RECT 9.780 7.650 9.950 7.820 ;
        RECT 10.230 7.650 10.400 7.820 ;
        RECT 10.680 7.650 10.850 7.820 ;
        RECT 11.130 7.650 11.300 7.820 ;
        RECT 11.580 7.650 11.750 7.820 ;
        RECT 12.030 7.650 12.200 7.820 ;
        RECT 12.480 7.650 12.650 7.820 ;
        RECT 12.930 7.650 13.100 7.820 ;
        RECT 13.380 7.650 13.550 7.820 ;
        RECT 14.230 7.650 14.400 7.820 ;
        RECT 14.680 7.650 14.850 7.820 ;
        RECT 15.130 7.650 15.300 7.820 ;
        RECT 15.580 7.650 15.750 7.820 ;
        RECT 16.030 7.650 16.200 7.820 ;
        RECT 16.480 7.650 16.650 7.820 ;
        RECT 16.930 7.650 17.100 7.820 ;
        RECT 17.380 7.650 17.550 7.820 ;
        RECT 17.830 7.650 18.000 7.820 ;
        RECT 18.280 7.650 18.450 7.820 ;
        RECT 18.730 7.650 18.900 7.820 ;
        RECT 19.180 7.650 19.350 7.820 ;
        RECT 19.630 7.650 19.800 7.820 ;
        RECT 20.080 7.650 20.250 7.820 ;
        RECT 20.930 7.650 21.100 7.820 ;
        RECT 21.380 7.650 21.550 7.820 ;
        RECT 21.830 7.650 22.000 7.820 ;
        RECT 22.280 7.650 22.450 7.820 ;
        RECT 22.730 7.650 22.900 7.820 ;
        RECT 23.180 7.650 23.350 7.820 ;
        RECT 23.630 7.650 23.800 7.820 ;
        RECT 24.080 7.650 24.250 7.820 ;
        RECT 24.530 7.650 24.700 7.820 ;
        RECT 24.980 7.650 25.150 7.820 ;
        RECT 25.430 7.650 25.600 7.820 ;
        RECT 25.880 7.650 26.050 7.820 ;
        RECT 26.330 7.650 26.500 7.820 ;
        RECT 26.780 7.650 26.950 7.820 ;
        RECT 27.630 7.650 27.800 7.820 ;
        RECT 28.080 7.650 28.250 7.820 ;
        RECT 28.530 7.650 28.700 7.820 ;
        RECT 28.980 7.650 29.150 7.820 ;
        RECT 29.430 7.650 29.600 7.820 ;
        RECT 29.880 7.650 30.050 7.820 ;
        RECT 30.330 7.650 30.500 7.820 ;
        RECT 30.780 7.650 30.950 7.820 ;
        RECT 31.230 7.650 31.400 7.820 ;
        RECT 31.680 7.650 31.850 7.820 ;
        RECT 32.130 7.650 32.300 7.820 ;
        RECT 32.580 7.650 32.750 7.820 ;
        RECT 33.030 7.650 33.200 7.820 ;
        RECT 33.480 7.650 33.650 7.820 ;
        RECT 34.330 7.650 34.500 7.820 ;
        RECT 34.780 7.650 34.950 7.820 ;
        RECT 35.230 7.650 35.400 7.820 ;
        RECT 35.680 7.650 35.850 7.820 ;
        RECT 36.130 7.650 36.300 7.820 ;
        RECT 36.580 7.650 36.750 7.820 ;
        RECT 37.030 7.650 37.200 7.820 ;
        RECT 37.480 7.650 37.650 7.820 ;
        RECT 37.930 7.650 38.100 7.820 ;
        RECT 38.380 7.650 38.550 7.820 ;
        RECT 38.830 7.650 39.000 7.820 ;
        RECT 39.280 7.650 39.450 7.820 ;
        RECT 39.730 7.650 39.900 7.820 ;
        RECT 40.180 7.650 40.350 7.820 ;
        RECT 41.030 7.650 41.200 7.820 ;
        RECT 41.480 7.650 41.650 7.820 ;
        RECT 41.930 7.650 42.100 7.820 ;
        RECT 42.380 7.650 42.550 7.820 ;
        RECT 42.830 7.650 43.000 7.820 ;
        RECT 43.280 7.650 43.450 7.820 ;
        RECT 43.730 7.650 43.900 7.820 ;
        RECT 44.180 7.650 44.350 7.820 ;
        RECT 44.630 7.650 44.800 7.820 ;
        RECT 45.080 7.650 45.250 7.820 ;
        RECT 45.530 7.650 45.700 7.820 ;
        RECT 45.980 7.650 46.150 7.820 ;
        RECT 46.430 7.650 46.600 7.820 ;
        RECT 46.880 7.650 47.050 7.820 ;
        RECT 47.730 7.650 47.900 7.820 ;
        RECT 48.180 7.650 48.350 7.820 ;
        RECT 48.630 7.650 48.800 7.820 ;
        RECT 49.080 7.650 49.250 7.820 ;
        RECT 49.530 7.650 49.700 7.820 ;
        RECT 49.980 7.650 50.150 7.820 ;
        RECT 50.430 7.650 50.600 7.820 ;
        RECT 50.880 7.650 51.050 7.820 ;
        RECT 51.330 7.650 51.500 7.820 ;
        RECT 51.780 7.650 51.950 7.820 ;
        RECT 52.230 7.650 52.400 7.820 ;
        RECT 52.680 7.650 52.850 7.820 ;
        RECT 53.130 7.650 53.300 7.820 ;
        RECT 53.580 7.650 53.750 7.820 ;
        RECT 1.650 6.850 1.820 7.020 ;
        RECT 2.100 6.850 2.270 7.020 ;
        RECT 2.550 6.850 2.720 7.020 ;
        RECT 3.000 6.850 3.170 7.020 ;
        RECT 3.450 6.850 3.620 7.020 ;
        RECT 3.900 6.850 4.070 7.020 ;
        RECT 4.350 6.850 4.520 7.020 ;
        RECT 4.800 6.850 4.970 7.020 ;
        RECT 5.250 6.850 5.420 7.020 ;
        RECT 5.700 6.850 5.870 7.020 ;
        RECT 6.150 6.850 6.320 7.020 ;
        RECT 2.580 5.830 2.750 6.000 ;
        RECT 3.080 5.830 3.250 6.000 ;
        RECT 3.580 5.830 3.750 6.000 ;
        RECT 4.080 5.830 4.250 6.000 ;
        RECT 4.580 5.830 4.750 6.000 ;
        RECT 5.080 5.830 5.250 6.000 ;
        RECT 2.580 5.330 2.750 5.500 ;
        RECT 3.080 5.330 3.250 5.500 ;
        RECT 3.580 5.330 3.750 5.500 ;
        RECT 4.080 5.330 4.250 5.500 ;
        RECT 4.580 5.330 4.750 5.500 ;
        RECT 5.080 5.330 5.250 5.500 ;
        RECT 2.580 4.830 2.750 5.000 ;
        RECT 3.080 4.830 3.250 5.000 ;
        RECT 3.580 4.830 3.750 5.000 ;
        RECT 4.080 4.830 4.250 5.000 ;
        RECT 4.580 4.830 4.750 5.000 ;
        RECT 5.080 4.830 5.250 5.000 ;
        RECT 2.580 4.330 2.750 4.500 ;
        RECT 3.080 4.330 3.250 4.500 ;
        RECT 3.580 4.330 3.750 4.500 ;
        RECT 4.080 4.330 4.250 4.500 ;
        RECT 4.580 4.330 4.750 4.500 ;
        RECT 5.080 4.330 5.250 4.500 ;
        RECT 2.580 3.830 2.750 4.000 ;
        RECT 3.080 3.830 3.250 4.000 ;
        RECT 3.580 3.830 3.750 4.000 ;
        RECT 4.080 3.830 4.250 4.000 ;
        RECT 4.580 3.830 4.750 4.000 ;
        RECT 5.080 3.830 5.250 4.000 ;
        RECT 2.580 3.330 2.750 3.500 ;
        RECT 3.080 3.330 3.250 3.500 ;
        RECT 3.580 3.330 3.750 3.500 ;
        RECT 4.080 3.330 4.250 3.500 ;
        RECT 4.580 3.330 4.750 3.500 ;
        RECT 5.080 3.330 5.250 3.500 ;
        RECT 8.350 6.850 8.520 7.020 ;
        RECT 8.800 6.850 8.970 7.020 ;
        RECT 9.250 6.850 9.420 7.020 ;
        RECT 9.700 6.850 9.870 7.020 ;
        RECT 10.150 6.850 10.320 7.020 ;
        RECT 10.600 6.850 10.770 7.020 ;
        RECT 11.050 6.850 11.220 7.020 ;
        RECT 11.500 6.850 11.670 7.020 ;
        RECT 11.950 6.850 12.120 7.020 ;
        RECT 12.400 6.850 12.570 7.020 ;
        RECT 12.850 6.850 13.020 7.020 ;
        RECT 9.280 5.830 9.450 6.000 ;
        RECT 9.780 5.830 9.950 6.000 ;
        RECT 10.280 5.830 10.450 6.000 ;
        RECT 10.780 5.830 10.950 6.000 ;
        RECT 11.280 5.830 11.450 6.000 ;
        RECT 11.780 5.830 11.950 6.000 ;
        RECT 9.280 5.330 9.450 5.500 ;
        RECT 9.780 5.330 9.950 5.500 ;
        RECT 10.280 5.330 10.450 5.500 ;
        RECT 10.780 5.330 10.950 5.500 ;
        RECT 11.280 5.330 11.450 5.500 ;
        RECT 11.780 5.330 11.950 5.500 ;
        RECT 9.280 4.830 9.450 5.000 ;
        RECT 9.780 4.830 9.950 5.000 ;
        RECT 10.280 4.830 10.450 5.000 ;
        RECT 10.780 4.830 10.950 5.000 ;
        RECT 11.280 4.830 11.450 5.000 ;
        RECT 11.780 4.830 11.950 5.000 ;
        RECT 9.280 4.330 9.450 4.500 ;
        RECT 9.780 4.330 9.950 4.500 ;
        RECT 10.280 4.330 10.450 4.500 ;
        RECT 10.780 4.330 10.950 4.500 ;
        RECT 11.280 4.330 11.450 4.500 ;
        RECT 11.780 4.330 11.950 4.500 ;
        RECT 9.280 3.830 9.450 4.000 ;
        RECT 9.780 3.830 9.950 4.000 ;
        RECT 10.280 3.830 10.450 4.000 ;
        RECT 10.780 3.830 10.950 4.000 ;
        RECT 11.280 3.830 11.450 4.000 ;
        RECT 11.780 3.830 11.950 4.000 ;
        RECT 9.280 3.330 9.450 3.500 ;
        RECT 9.780 3.330 9.950 3.500 ;
        RECT 10.280 3.330 10.450 3.500 ;
        RECT 10.780 3.330 10.950 3.500 ;
        RECT 11.280 3.330 11.450 3.500 ;
        RECT 11.780 3.330 11.950 3.500 ;
        RECT 15.050 6.850 15.220 7.020 ;
        RECT 15.500 6.850 15.670 7.020 ;
        RECT 15.950 6.850 16.120 7.020 ;
        RECT 16.400 6.850 16.570 7.020 ;
        RECT 16.850 6.850 17.020 7.020 ;
        RECT 17.300 6.850 17.470 7.020 ;
        RECT 17.750 6.850 17.920 7.020 ;
        RECT 18.200 6.850 18.370 7.020 ;
        RECT 18.650 6.850 18.820 7.020 ;
        RECT 19.100 6.850 19.270 7.020 ;
        RECT 19.550 6.850 19.720 7.020 ;
        RECT 15.980 5.830 16.150 6.000 ;
        RECT 16.480 5.830 16.650 6.000 ;
        RECT 16.980 5.830 17.150 6.000 ;
        RECT 17.480 5.830 17.650 6.000 ;
        RECT 17.980 5.830 18.150 6.000 ;
        RECT 18.480 5.830 18.650 6.000 ;
        RECT 15.980 5.330 16.150 5.500 ;
        RECT 16.480 5.330 16.650 5.500 ;
        RECT 16.980 5.330 17.150 5.500 ;
        RECT 17.480 5.330 17.650 5.500 ;
        RECT 17.980 5.330 18.150 5.500 ;
        RECT 18.480 5.330 18.650 5.500 ;
        RECT 15.980 4.830 16.150 5.000 ;
        RECT 16.480 4.830 16.650 5.000 ;
        RECT 16.980 4.830 17.150 5.000 ;
        RECT 17.480 4.830 17.650 5.000 ;
        RECT 17.980 4.830 18.150 5.000 ;
        RECT 18.480 4.830 18.650 5.000 ;
        RECT 15.980 4.330 16.150 4.500 ;
        RECT 16.480 4.330 16.650 4.500 ;
        RECT 16.980 4.330 17.150 4.500 ;
        RECT 17.480 4.330 17.650 4.500 ;
        RECT 17.980 4.330 18.150 4.500 ;
        RECT 18.480 4.330 18.650 4.500 ;
        RECT 15.980 3.830 16.150 4.000 ;
        RECT 16.480 3.830 16.650 4.000 ;
        RECT 16.980 3.830 17.150 4.000 ;
        RECT 17.480 3.830 17.650 4.000 ;
        RECT 17.980 3.830 18.150 4.000 ;
        RECT 18.480 3.830 18.650 4.000 ;
        RECT 15.980 3.330 16.150 3.500 ;
        RECT 16.480 3.330 16.650 3.500 ;
        RECT 16.980 3.330 17.150 3.500 ;
        RECT 17.480 3.330 17.650 3.500 ;
        RECT 17.980 3.330 18.150 3.500 ;
        RECT 18.480 3.330 18.650 3.500 ;
        RECT 21.750 6.850 21.920 7.020 ;
        RECT 22.200 6.850 22.370 7.020 ;
        RECT 22.650 6.850 22.820 7.020 ;
        RECT 23.100 6.850 23.270 7.020 ;
        RECT 23.550 6.850 23.720 7.020 ;
        RECT 24.000 6.850 24.170 7.020 ;
        RECT 24.450 6.850 24.620 7.020 ;
        RECT 24.900 6.850 25.070 7.020 ;
        RECT 25.350 6.850 25.520 7.020 ;
        RECT 25.800 6.850 25.970 7.020 ;
        RECT 26.250 6.850 26.420 7.020 ;
        RECT 22.680 5.830 22.850 6.000 ;
        RECT 23.180 5.830 23.350 6.000 ;
        RECT 23.680 5.830 23.850 6.000 ;
        RECT 24.180 5.830 24.350 6.000 ;
        RECT 24.680 5.830 24.850 6.000 ;
        RECT 25.180 5.830 25.350 6.000 ;
        RECT 22.680 5.330 22.850 5.500 ;
        RECT 23.180 5.330 23.350 5.500 ;
        RECT 23.680 5.330 23.850 5.500 ;
        RECT 24.180 5.330 24.350 5.500 ;
        RECT 24.680 5.330 24.850 5.500 ;
        RECT 25.180 5.330 25.350 5.500 ;
        RECT 22.680 4.830 22.850 5.000 ;
        RECT 23.180 4.830 23.350 5.000 ;
        RECT 23.680 4.830 23.850 5.000 ;
        RECT 24.180 4.830 24.350 5.000 ;
        RECT 24.680 4.830 24.850 5.000 ;
        RECT 25.180 4.830 25.350 5.000 ;
        RECT 22.680 4.330 22.850 4.500 ;
        RECT 23.180 4.330 23.350 4.500 ;
        RECT 23.680 4.330 23.850 4.500 ;
        RECT 24.180 4.330 24.350 4.500 ;
        RECT 24.680 4.330 24.850 4.500 ;
        RECT 25.180 4.330 25.350 4.500 ;
        RECT 22.680 3.830 22.850 4.000 ;
        RECT 23.180 3.830 23.350 4.000 ;
        RECT 23.680 3.830 23.850 4.000 ;
        RECT 24.180 3.830 24.350 4.000 ;
        RECT 24.680 3.830 24.850 4.000 ;
        RECT 25.180 3.830 25.350 4.000 ;
        RECT 22.680 3.330 22.850 3.500 ;
        RECT 23.180 3.330 23.350 3.500 ;
        RECT 23.680 3.330 23.850 3.500 ;
        RECT 24.180 3.330 24.350 3.500 ;
        RECT 24.680 3.330 24.850 3.500 ;
        RECT 25.180 3.330 25.350 3.500 ;
        RECT 28.450 6.850 28.620 7.020 ;
        RECT 28.900 6.850 29.070 7.020 ;
        RECT 29.350 6.850 29.520 7.020 ;
        RECT 29.800 6.850 29.970 7.020 ;
        RECT 30.250 6.850 30.420 7.020 ;
        RECT 30.700 6.850 30.870 7.020 ;
        RECT 31.150 6.850 31.320 7.020 ;
        RECT 31.600 6.850 31.770 7.020 ;
        RECT 32.050 6.850 32.220 7.020 ;
        RECT 32.500 6.850 32.670 7.020 ;
        RECT 32.950 6.850 33.120 7.020 ;
        RECT 29.380 5.830 29.550 6.000 ;
        RECT 29.880 5.830 30.050 6.000 ;
        RECT 30.380 5.830 30.550 6.000 ;
        RECT 30.880 5.830 31.050 6.000 ;
        RECT 31.380 5.830 31.550 6.000 ;
        RECT 31.880 5.830 32.050 6.000 ;
        RECT 29.380 5.330 29.550 5.500 ;
        RECT 29.880 5.330 30.050 5.500 ;
        RECT 30.380 5.330 30.550 5.500 ;
        RECT 30.880 5.330 31.050 5.500 ;
        RECT 31.380 5.330 31.550 5.500 ;
        RECT 31.880 5.330 32.050 5.500 ;
        RECT 29.380 4.830 29.550 5.000 ;
        RECT 29.880 4.830 30.050 5.000 ;
        RECT 30.380 4.830 30.550 5.000 ;
        RECT 30.880 4.830 31.050 5.000 ;
        RECT 31.380 4.830 31.550 5.000 ;
        RECT 31.880 4.830 32.050 5.000 ;
        RECT 29.380 4.330 29.550 4.500 ;
        RECT 29.880 4.330 30.050 4.500 ;
        RECT 30.380 4.330 30.550 4.500 ;
        RECT 30.880 4.330 31.050 4.500 ;
        RECT 31.380 4.330 31.550 4.500 ;
        RECT 31.880 4.330 32.050 4.500 ;
        RECT 29.380 3.830 29.550 4.000 ;
        RECT 29.880 3.830 30.050 4.000 ;
        RECT 30.380 3.830 30.550 4.000 ;
        RECT 30.880 3.830 31.050 4.000 ;
        RECT 31.380 3.830 31.550 4.000 ;
        RECT 31.880 3.830 32.050 4.000 ;
        RECT 29.380 3.330 29.550 3.500 ;
        RECT 29.880 3.330 30.050 3.500 ;
        RECT 30.380 3.330 30.550 3.500 ;
        RECT 30.880 3.330 31.050 3.500 ;
        RECT 31.380 3.330 31.550 3.500 ;
        RECT 31.880 3.330 32.050 3.500 ;
        RECT 35.150 6.850 35.320 7.020 ;
        RECT 35.600 6.850 35.770 7.020 ;
        RECT 36.050 6.850 36.220 7.020 ;
        RECT 36.500 6.850 36.670 7.020 ;
        RECT 36.950 6.850 37.120 7.020 ;
        RECT 37.400 6.850 37.570 7.020 ;
        RECT 37.850 6.850 38.020 7.020 ;
        RECT 38.300 6.850 38.470 7.020 ;
        RECT 38.750 6.850 38.920 7.020 ;
        RECT 39.200 6.850 39.370 7.020 ;
        RECT 39.650 6.850 39.820 7.020 ;
        RECT 36.080 5.830 36.250 6.000 ;
        RECT 36.580 5.830 36.750 6.000 ;
        RECT 37.080 5.830 37.250 6.000 ;
        RECT 37.580 5.830 37.750 6.000 ;
        RECT 38.080 5.830 38.250 6.000 ;
        RECT 38.580 5.830 38.750 6.000 ;
        RECT 36.080 5.330 36.250 5.500 ;
        RECT 36.580 5.330 36.750 5.500 ;
        RECT 37.080 5.330 37.250 5.500 ;
        RECT 37.580 5.330 37.750 5.500 ;
        RECT 38.080 5.330 38.250 5.500 ;
        RECT 38.580 5.330 38.750 5.500 ;
        RECT 36.080 4.830 36.250 5.000 ;
        RECT 36.580 4.830 36.750 5.000 ;
        RECT 37.080 4.830 37.250 5.000 ;
        RECT 37.580 4.830 37.750 5.000 ;
        RECT 38.080 4.830 38.250 5.000 ;
        RECT 38.580 4.830 38.750 5.000 ;
        RECT 36.080 4.330 36.250 4.500 ;
        RECT 36.580 4.330 36.750 4.500 ;
        RECT 37.080 4.330 37.250 4.500 ;
        RECT 37.580 4.330 37.750 4.500 ;
        RECT 38.080 4.330 38.250 4.500 ;
        RECT 38.580 4.330 38.750 4.500 ;
        RECT 36.080 3.830 36.250 4.000 ;
        RECT 36.580 3.830 36.750 4.000 ;
        RECT 37.080 3.830 37.250 4.000 ;
        RECT 37.580 3.830 37.750 4.000 ;
        RECT 38.080 3.830 38.250 4.000 ;
        RECT 38.580 3.830 38.750 4.000 ;
        RECT 36.080 3.330 36.250 3.500 ;
        RECT 36.580 3.330 36.750 3.500 ;
        RECT 37.080 3.330 37.250 3.500 ;
        RECT 37.580 3.330 37.750 3.500 ;
        RECT 38.080 3.330 38.250 3.500 ;
        RECT 38.580 3.330 38.750 3.500 ;
        RECT 41.850 6.850 42.020 7.020 ;
        RECT 42.300 6.850 42.470 7.020 ;
        RECT 42.750 6.850 42.920 7.020 ;
        RECT 43.200 6.850 43.370 7.020 ;
        RECT 43.650 6.850 43.820 7.020 ;
        RECT 44.100 6.850 44.270 7.020 ;
        RECT 44.550 6.850 44.720 7.020 ;
        RECT 45.000 6.850 45.170 7.020 ;
        RECT 45.450 6.850 45.620 7.020 ;
        RECT 45.900 6.850 46.070 7.020 ;
        RECT 46.350 6.850 46.520 7.020 ;
        RECT 42.780 5.830 42.950 6.000 ;
        RECT 43.280 5.830 43.450 6.000 ;
        RECT 43.780 5.830 43.950 6.000 ;
        RECT 44.280 5.830 44.450 6.000 ;
        RECT 44.780 5.830 44.950 6.000 ;
        RECT 45.280 5.830 45.450 6.000 ;
        RECT 42.780 5.330 42.950 5.500 ;
        RECT 43.280 5.330 43.450 5.500 ;
        RECT 43.780 5.330 43.950 5.500 ;
        RECT 44.280 5.330 44.450 5.500 ;
        RECT 44.780 5.330 44.950 5.500 ;
        RECT 45.280 5.330 45.450 5.500 ;
        RECT 42.780 4.830 42.950 5.000 ;
        RECT 43.280 4.830 43.450 5.000 ;
        RECT 43.780 4.830 43.950 5.000 ;
        RECT 44.280 4.830 44.450 5.000 ;
        RECT 44.780 4.830 44.950 5.000 ;
        RECT 45.280 4.830 45.450 5.000 ;
        RECT 42.780 4.330 42.950 4.500 ;
        RECT 43.280 4.330 43.450 4.500 ;
        RECT 43.780 4.330 43.950 4.500 ;
        RECT 44.280 4.330 44.450 4.500 ;
        RECT 44.780 4.330 44.950 4.500 ;
        RECT 45.280 4.330 45.450 4.500 ;
        RECT 42.780 3.830 42.950 4.000 ;
        RECT 43.280 3.830 43.450 4.000 ;
        RECT 43.780 3.830 43.950 4.000 ;
        RECT 44.280 3.830 44.450 4.000 ;
        RECT 44.780 3.830 44.950 4.000 ;
        RECT 45.280 3.830 45.450 4.000 ;
        RECT 42.780 3.330 42.950 3.500 ;
        RECT 43.280 3.330 43.450 3.500 ;
        RECT 43.780 3.330 43.950 3.500 ;
        RECT 44.280 3.330 44.450 3.500 ;
        RECT 44.780 3.330 44.950 3.500 ;
        RECT 45.280 3.330 45.450 3.500 ;
        RECT 48.550 6.850 48.720 7.020 ;
        RECT 49.000 6.850 49.170 7.020 ;
        RECT 49.450 6.850 49.620 7.020 ;
        RECT 49.900 6.850 50.070 7.020 ;
        RECT 50.350 6.850 50.520 7.020 ;
        RECT 50.800 6.850 50.970 7.020 ;
        RECT 51.250 6.850 51.420 7.020 ;
        RECT 51.700 6.850 51.870 7.020 ;
        RECT 52.150 6.850 52.320 7.020 ;
        RECT 52.600 6.850 52.770 7.020 ;
        RECT 53.050 6.850 53.220 7.020 ;
        RECT 49.480 5.830 49.650 6.000 ;
        RECT 49.980 5.830 50.150 6.000 ;
        RECT 50.480 5.830 50.650 6.000 ;
        RECT 50.980 5.830 51.150 6.000 ;
        RECT 51.480 5.830 51.650 6.000 ;
        RECT 51.980 5.830 52.150 6.000 ;
        RECT 49.480 5.330 49.650 5.500 ;
        RECT 49.980 5.330 50.150 5.500 ;
        RECT 50.480 5.330 50.650 5.500 ;
        RECT 50.980 5.330 51.150 5.500 ;
        RECT 51.480 5.330 51.650 5.500 ;
        RECT 51.980 5.330 52.150 5.500 ;
        RECT 49.480 4.830 49.650 5.000 ;
        RECT 49.980 4.830 50.150 5.000 ;
        RECT 50.480 4.830 50.650 5.000 ;
        RECT 50.980 4.830 51.150 5.000 ;
        RECT 51.480 4.830 51.650 5.000 ;
        RECT 51.980 4.830 52.150 5.000 ;
        RECT 49.480 4.330 49.650 4.500 ;
        RECT 49.980 4.330 50.150 4.500 ;
        RECT 50.480 4.330 50.650 4.500 ;
        RECT 50.980 4.330 51.150 4.500 ;
        RECT 51.480 4.330 51.650 4.500 ;
        RECT 51.980 4.330 52.150 4.500 ;
        RECT 49.480 3.830 49.650 4.000 ;
        RECT 49.980 3.830 50.150 4.000 ;
        RECT 50.480 3.830 50.650 4.000 ;
        RECT 50.980 3.830 51.150 4.000 ;
        RECT 51.480 3.830 51.650 4.000 ;
        RECT 51.980 3.830 52.150 4.000 ;
        RECT 49.480 3.330 49.650 3.500 ;
        RECT 49.980 3.330 50.150 3.500 ;
        RECT 50.480 3.330 50.650 3.500 ;
        RECT 50.980 3.330 51.150 3.500 ;
        RECT 51.480 3.330 51.650 3.500 ;
        RECT 51.980 3.330 52.150 3.500 ;
        RECT 1.450 -0.150 1.750 0.150 ;
        RECT 2.450 -0.150 2.750 0.150 ;
        RECT 3.450 -0.150 3.750 0.150 ;
        RECT 4.450 -0.150 4.750 0.150 ;
        RECT 5.450 -0.150 5.750 0.150 ;
        RECT 6.450 -0.150 6.750 0.150 ;
        RECT 7.450 -0.150 7.750 0.150 ;
        RECT 8.450 -0.150 8.750 0.150 ;
        RECT 9.450 -0.150 9.750 0.150 ;
        RECT 10.450 -0.150 10.750 0.150 ;
        RECT 11.450 -0.150 11.750 0.150 ;
        RECT 12.450 -0.150 12.750 0.150 ;
        RECT 13.450 -0.150 13.750 0.150 ;
        RECT 14.450 -0.150 14.750 0.150 ;
        RECT 15.450 -0.150 15.750 0.150 ;
        RECT 16.450 -0.150 16.750 0.150 ;
        RECT 17.450 -0.150 17.750 0.150 ;
        RECT 18.450 -0.150 18.750 0.150 ;
        RECT 19.450 -0.150 19.750 0.150 ;
        RECT 20.450 -0.150 20.750 0.150 ;
        RECT 21.450 -0.150 21.750 0.150 ;
        RECT 22.450 -0.150 22.750 0.150 ;
        RECT 23.450 -0.150 23.750 0.150 ;
        RECT 24.450 -0.150 24.750 0.150 ;
        RECT 25.450 -0.150 25.750 0.150 ;
        RECT 26.450 -0.150 26.750 0.150 ;
        RECT 27.450 -0.150 27.750 0.150 ;
        RECT 28.450 -0.150 28.750 0.150 ;
        RECT 29.450 -0.150 29.750 0.150 ;
        RECT 30.450 -0.150 30.750 0.150 ;
        RECT 31.450 -0.150 31.750 0.150 ;
        RECT 32.450 -0.150 32.750 0.150 ;
        RECT 33.450 -0.150 33.750 0.150 ;
        RECT 34.450 -0.150 34.750 0.150 ;
        RECT 35.450 -0.150 35.750 0.150 ;
        RECT 36.450 -0.150 36.750 0.150 ;
        RECT 37.450 -0.150 37.750 0.150 ;
        RECT 38.450 -0.150 38.750 0.150 ;
        RECT 39.450 -0.150 39.750 0.150 ;
        RECT 40.450 -0.150 40.750 0.150 ;
        RECT 41.450 -0.150 41.750 0.150 ;
        RECT 42.450 -0.150 42.750 0.150 ;
        RECT 43.450 -0.150 43.750 0.150 ;
        RECT 44.450 -0.150 44.750 0.150 ;
        RECT 45.450 -0.150 45.750 0.150 ;
        RECT 46.450 -0.150 46.750 0.150 ;
        RECT 47.450 -0.150 47.750 0.150 ;
        RECT 48.450 -0.150 48.750 0.150 ;
        RECT 49.450 -0.150 49.750 0.150 ;
        RECT 50.450 -0.150 50.750 0.150 ;
        RECT 51.450 -0.150 51.750 0.150 ;
        RECT 52.450 -0.150 52.750 0.150 ;
        RECT 53.450 -0.150 53.750 0.150 ;
  END
END sky130_asc_pnp_05v5_W3p40L3p40_8
END LIBRARY

