VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO sky130_fd_pr__cap_mim_m3_1
  CLASS CORE ;
  FOREIGN sky130_fd_pr__cap_mim_m3_1 ;
  ORIGIN 0.000 0.000 ;
  SIZE 35.855 BY 9.400 ;
  SITE unitasc ;
  PIN c0
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT -0.100 8.250 35.750 8.450 ;
        RECT -0.100 5.250 35.755 8.250 ;
        RECT -0.100 4.750 35.750 5.250 ;
        RECT -0.100 1.750 35.755 4.750 ;
      LAYER via3 ;
        RECT 2.980 5.390 3.300 8.110 ;
        RECT 6.575 5.390 6.895 8.110 ;
        RECT 10.170 5.390 10.490 8.110 ;
        RECT 13.765 5.390 14.085 8.110 ;
        RECT 17.360 5.390 17.680 8.110 ;
        RECT 20.955 5.390 21.275 8.110 ;
        RECT 24.550 5.390 24.870 8.110 ;
        RECT 28.145 5.390 28.465 8.110 ;
        RECT 31.740 5.390 32.060 8.110 ;
        RECT 35.335 5.390 35.655 8.110 ;
        RECT 2.980 1.890 3.300 4.610 ;
        RECT 6.575 1.890 6.895 4.610 ;
        RECT 10.170 1.890 10.490 4.610 ;
        RECT 13.765 1.890 14.085 4.610 ;
        RECT 17.360 1.890 17.680 4.610 ;
        RECT 20.955 1.890 21.275 4.610 ;
        RECT 24.550 1.890 24.870 4.610 ;
        RECT 28.145 1.890 28.465 4.610 ;
        RECT 31.740 1.890 32.060 4.610 ;
        RECT 35.335 1.890 35.655 4.610 ;
      LAYER met4 ;
        RECT 2.900 5.310 3.380 8.190 ;
        RECT 6.495 5.310 6.975 8.190 ;
        RECT 10.090 5.310 10.570 8.190 ;
        RECT 13.685 5.310 14.165 8.190 ;
        RECT 17.280 5.310 17.760 8.190 ;
        RECT 20.875 5.310 21.355 8.190 ;
        RECT 24.470 5.310 24.950 8.190 ;
        RECT 28.065 5.310 28.545 8.190 ;
        RECT 31.660 5.310 32.140 8.190 ;
        RECT 35.255 5.310 35.735 8.190 ;
        RECT 2.900 1.810 3.380 4.690 ;
        RECT 6.495 1.810 6.975 4.690 ;
        RECT 10.090 1.810 10.570 4.690 ;
        RECT 13.685 1.810 14.165 4.690 ;
        RECT 17.280 1.810 17.760 4.690 ;
        RECT 20.875 1.810 21.355 4.690 ;
        RECT 24.470 1.810 24.950 4.690 ;
        RECT 28.065 1.810 28.545 4.690 ;
        RECT 31.660 1.810 32.140 4.690 ;
        RECT 35.255 1.810 35.735 4.690 ;
    END
  END c0
  PIN c1
    DIRECTION INOUT ;
    PORT
      LAYER met4 ;
        RECT 0.600 7.555 2.200 7.650 ;
        RECT 4.200 7.555 5.800 7.650 ;
        RECT 7.800 7.555 9.400 7.650 ;
        RECT 11.400 7.555 13.000 7.650 ;
        RECT 15.000 7.555 16.600 7.650 ;
        RECT 18.600 7.555 20.200 7.650 ;
        RECT 22.200 7.555 23.800 7.650 ;
        RECT 25.800 7.555 27.400 7.650 ;
        RECT 29.400 7.555 31.000 7.650 ;
        RECT 33.000 7.555 34.600 7.650 ;
        RECT 0.600 5.945 2.210 7.555 ;
        RECT 4.195 5.945 5.805 7.555 ;
        RECT 7.790 5.945 9.400 7.555 ;
        RECT 11.385 5.945 13.000 7.555 ;
        RECT 14.980 5.945 16.600 7.555 ;
        RECT 18.575 5.945 20.200 7.555 ;
        RECT 22.170 5.945 23.800 7.555 ;
        RECT 25.765 5.945 27.400 7.555 ;
        RECT 29.360 5.945 31.000 7.555 ;
        RECT 32.955 5.945 34.600 7.555 ;
        RECT 0.600 4.055 2.200 5.945 ;
        RECT 4.200 4.055 5.800 5.945 ;
        RECT 7.800 4.055 9.400 5.945 ;
        RECT 11.400 4.055 13.000 5.945 ;
        RECT 15.000 4.055 16.600 5.945 ;
        RECT 18.600 4.055 20.200 5.945 ;
        RECT 22.200 4.055 23.800 5.945 ;
        RECT 25.800 4.055 27.400 5.945 ;
        RECT 29.400 4.055 31.000 5.945 ;
        RECT 33.000 4.055 34.600 5.945 ;
        RECT 0.600 2.445 2.210 4.055 ;
        RECT 4.195 2.445 5.805 4.055 ;
        RECT 7.790 2.445 9.400 4.055 ;
        RECT 11.385 2.445 13.000 4.055 ;
        RECT 14.980 2.445 16.600 4.055 ;
        RECT 18.575 2.445 20.200 4.055 ;
        RECT 22.170 2.445 23.800 4.055 ;
        RECT 25.765 2.445 27.400 4.055 ;
        RECT 29.360 2.445 31.000 4.055 ;
        RECT 32.955 2.445 34.600 4.055 ;
        RECT 0.600 1.450 2.200 2.445 ;
        RECT 4.200 1.450 5.800 2.445 ;
        RECT 7.800 1.450 9.400 2.445 ;
        RECT 11.400 1.450 13.000 2.445 ;
        RECT 15.000 1.450 16.600 2.445 ;
        RECT 18.600 1.450 20.200 2.445 ;
        RECT 22.200 1.450 23.800 2.445 ;
        RECT 25.800 1.450 27.400 2.445 ;
        RECT 29.400 1.450 31.000 2.445 ;
        RECT 33.000 1.450 34.600 2.445 ;
        RECT -0.090 0.950 35.750 1.450 ;
    END
  END c1
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER li1 ;
        RECT -0.090 9.250 35.750 9.550 ;
      LAYER mcon ;
        RECT 0.760 9.250 1.060 9.550 ;
        RECT 2.760 9.250 3.060 9.550 ;
        RECT 4.760 9.250 5.060 9.550 ;
        RECT 6.760 9.250 7.060 9.550 ;
        RECT 8.760 9.250 9.060 9.550 ;
        RECT 10.760 9.250 11.060 9.550 ;
        RECT 12.760 9.250 13.060 9.550 ;
        RECT 14.760 9.250 15.060 9.550 ;
        RECT 16.760 9.250 17.060 9.550 ;
        RECT 18.760 9.250 19.060 9.550 ;
        RECT 20.760 9.250 21.060 9.550 ;
        RECT 22.760 9.250 23.060 9.550 ;
        RECT 24.760 9.250 25.060 9.550 ;
        RECT 26.760 9.250 27.060 9.550 ;
        RECT 28.760 9.250 29.060 9.550 ;
        RECT 30.760 9.250 31.060 9.550 ;
        RECT 32.760 9.250 33.060 9.550 ;
        RECT 34.760 9.250 35.060 9.550 ;
      LAYER met1 ;
        RECT -0.090 9.100 35.750 9.700 ;
    END
  END VPWR
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER li1 ;
        RECT -0.090 -0.150 35.750 0.150 ;
      LAYER mcon ;
        RECT 0.760 -0.150 1.060 0.150 ;
        RECT 2.760 -0.150 3.060 0.150 ;
        RECT 4.760 -0.150 5.060 0.150 ;
        RECT 6.760 -0.150 7.060 0.150 ;
        RECT 8.760 -0.150 9.060 0.150 ;
        RECT 10.760 -0.150 11.060 0.150 ;
        RECT 12.760 -0.150 13.060 0.150 ;
        RECT 14.760 -0.150 15.060 0.150 ;
        RECT 16.760 -0.150 17.060 0.150 ;
        RECT 18.760 -0.150 19.060 0.150 ;
        RECT 20.760 -0.150 21.060 0.150 ;
        RECT 22.760 -0.150 23.060 0.150 ;
        RECT 24.760 -0.150 25.060 0.150 ;
        RECT 26.760 -0.150 27.060 0.150 ;
        RECT 28.760 -0.150 29.060 0.150 ;
        RECT 30.760 -0.150 31.060 0.150 ;
        RECT 32.760 -0.150 33.060 0.150 ;
        RECT 34.760 -0.150 35.060 0.150 ;
      LAYER met1 ;
        RECT -0.090 -0.300 35.750 0.300 ;
    END
  END VGND
END sky130_fd_pr__cap_mim_m3_1
END LIBRARY

