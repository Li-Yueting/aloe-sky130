* NGSPICE file created from sky130_asc_pfet_01v8_lvt_1.ext - technology: sky130A

.subckt sky130_asc_pfet_01v8_lvt_1 GATE SOURCE DRAIN VPWR VGND
X0 SOURCE GATE DRAIN w_130_293# sky130_fd_pr__pfet_01v8_lvt ad=1.8705e+12p pd=1.348e+07u as=1.8705e+12p ps=1.348e+07u w=6.45e+06u l=2e+06u
.ends

