magic
tech sky130A
magscale 1 2
timestamp 1658609783
<< nwell >>
rect 130 293 4382 1940
<< pmoslvt >>
rect 224 355 624 1645
rect 682 355 1082 1645
rect 1140 355 1540 1645
rect 1598 355 1998 1645
rect 2056 355 2456 1645
rect 2514 355 2914 1645
rect 2972 355 3372 1645
rect 3430 355 3830 1645
rect 3888 355 4288 1645
<< pdiff >>
rect 166 1633 224 1645
rect 166 367 178 1633
rect 212 367 224 1633
rect 166 355 224 367
rect 624 1633 682 1645
rect 624 367 636 1633
rect 670 367 682 1633
rect 624 355 682 367
rect 1082 1633 1140 1645
rect 1082 367 1094 1633
rect 1128 367 1140 1633
rect 1082 355 1140 367
rect 1540 1633 1598 1645
rect 1540 367 1552 1633
rect 1586 367 1598 1633
rect 1540 355 1598 367
rect 1998 1633 2056 1645
rect 1998 367 2010 1633
rect 2044 367 2056 1633
rect 1998 355 2056 367
rect 2456 1633 2514 1645
rect 2456 367 2468 1633
rect 2502 367 2514 1633
rect 2456 355 2514 367
rect 2914 1633 2972 1645
rect 2914 367 2926 1633
rect 2960 367 2972 1633
rect 2914 355 2972 367
rect 3372 1633 3430 1645
rect 3372 367 3384 1633
rect 3418 367 3430 1633
rect 3372 355 3430 367
rect 3830 1633 3888 1645
rect 3830 367 3842 1633
rect 3876 367 3888 1633
rect 3830 355 3888 367
rect 4288 1633 4346 1645
rect 4288 367 4300 1633
rect 4334 367 4346 1633
rect 4288 355 4346 367
<< pdiffc >>
rect 178 367 212 1633
rect 636 367 670 1633
rect 1094 367 1128 1633
rect 1552 367 1586 1633
rect 2010 367 2044 1633
rect 2468 367 2502 1633
rect 2926 367 2960 1633
rect 3384 367 3418 1633
rect 3842 367 3876 1633
rect 4300 367 4334 1633
<< poly >>
rect 224 1645 624 1671
rect 682 1645 1082 1671
rect 1140 1645 1540 1671
rect 1598 1645 1998 1671
rect 2056 1645 2456 1671
rect 2514 1645 2914 1671
rect 2972 1645 3372 1671
rect 3430 1645 3830 1671
rect 3888 1645 4288 1671
rect 224 329 624 355
rect 682 329 1082 355
rect 1140 329 1540 355
rect 1598 329 1998 355
rect 2056 329 2456 355
rect 2514 329 2914 355
rect 2972 329 3372 355
rect 3430 329 3830 355
rect 3888 329 4288 355
rect 370 182 490 329
rect 826 182 946 329
rect 1282 182 1402 329
rect 1738 182 1858 329
rect 2194 182 2314 329
rect 2650 182 2770 329
rect 3106 182 3226 329
rect 3562 182 3682 329
rect 4018 182 4138 329
rect 130 162 4382 182
rect 130 102 300 162
rect 360 102 700 162
rect 760 102 1100 162
rect 1160 102 1500 162
rect 1560 102 1900 162
rect 1960 102 2300 162
rect 2360 102 2700 162
rect 2760 102 3100 162
rect 3160 102 3500 162
rect 3560 102 3900 162
rect 3960 102 4382 162
rect 130 82 4382 102
<< polycont >>
rect 300 102 360 162
rect 700 102 760 162
rect 1100 102 1160 162
rect 1500 102 1560 162
rect 1900 102 1960 162
rect 2300 102 2360 162
rect 2700 102 2760 162
rect 3100 102 3160 162
rect 3500 102 3560 162
rect 3900 102 3960 162
<< locali >>
rect 130 1850 300 1910
rect 360 1850 700 1910
rect 760 1850 1100 1910
rect 1160 1850 1500 1910
rect 1560 1850 1900 1910
rect 1960 1850 2300 1910
rect 2360 1850 2700 1910
rect 2760 1850 3100 1910
rect 3160 1850 3500 1910
rect 3560 1850 3900 1910
rect 3960 1850 4382 1910
rect 130 1730 4382 1790
rect 635 1649 669 1730
rect 1551 1649 1585 1730
rect 2467 1649 2501 1730
rect 3383 1649 3417 1730
rect 4299 1649 4333 1730
rect 178 1633 212 1649
rect 177 367 178 372
rect 635 1633 670 1649
rect 635 1626 636 1633
rect 177 351 212 367
rect 1094 1633 1128 1649
rect 636 351 670 367
rect 1093 367 1094 372
rect 1551 1633 1586 1649
rect 1551 1626 1552 1633
rect 1093 351 1128 367
rect 2010 1633 2044 1649
rect 1552 351 1586 367
rect 2009 367 2010 372
rect 2467 1633 2502 1649
rect 2467 1626 2468 1633
rect 2009 351 2044 367
rect 2926 1633 2960 1649
rect 2468 351 2502 367
rect 2925 367 2926 372
rect 3383 1633 3418 1649
rect 3383 1626 3384 1633
rect 2925 351 2960 367
rect 3842 1633 3876 1649
rect 3384 351 3418 367
rect 3841 367 3842 372
rect 4299 1633 4334 1649
rect 4299 1626 4300 1633
rect 3841 351 3876 367
rect 4300 351 4334 367
rect 177 270 211 351
rect 1093 270 1127 351
rect 2009 270 2043 351
rect 2925 270 2959 351
rect 3841 270 3875 351
rect 130 210 4382 270
rect 130 102 300 162
rect 360 102 700 162
rect 760 102 1100 162
rect 1160 102 1500 162
rect 1560 102 1900 162
rect 1960 102 2300 162
rect 2360 102 2700 162
rect 2760 102 3100 162
rect 3160 102 3500 162
rect 3560 102 3900 162
rect 3960 102 4382 162
rect 130 -30 300 30
rect 360 -30 700 30
rect 760 -30 1100 30
rect 1160 -30 1500 30
rect 1560 -30 1900 30
rect 1960 -30 2300 30
rect 2360 -30 2700 30
rect 2760 -30 3100 30
rect 3160 -30 3500 30
rect 3560 -30 3900 30
rect 3960 -30 4382 30
<< viali >>
rect 300 1850 360 1910
rect 700 1850 760 1910
rect 1100 1850 1160 1910
rect 1500 1850 1560 1910
rect 1900 1850 1960 1910
rect 2300 1850 2360 1910
rect 2700 1850 2760 1910
rect 3100 1850 3160 1910
rect 3500 1850 3560 1910
rect 3900 1850 3960 1910
rect 178 367 212 1633
rect 636 367 670 1633
rect 1094 367 1128 1633
rect 1552 367 1586 1633
rect 2010 367 2044 1633
rect 2468 367 2502 1633
rect 2926 367 2960 1633
rect 3384 367 3418 1633
rect 3842 367 3876 1633
rect 4300 367 4334 1633
rect 300 -30 360 30
rect 700 -30 760 30
rect 1100 -30 1160 30
rect 1500 -30 1560 30
rect 1900 -30 1960 30
rect 2300 -30 2360 30
rect 2700 -30 2760 30
rect 3100 -30 3160 30
rect 3500 -30 3560 30
rect 3900 -30 3960 30
<< metal1 >>
rect 130 1910 4382 1940
rect 130 1850 300 1910
rect 360 1850 700 1910
rect 760 1850 1100 1910
rect 1160 1850 1500 1910
rect 1560 1850 1900 1910
rect 1960 1850 2300 1910
rect 2360 1850 2700 1910
rect 2760 1850 3100 1910
rect 3160 1850 3500 1910
rect 3560 1850 3900 1910
rect 3960 1850 4382 1910
rect 130 1820 4382 1850
rect 172 1633 218 1645
rect 172 367 178 1633
rect 212 367 218 1633
rect 172 355 218 367
rect 630 1633 676 1645
rect 630 367 636 1633
rect 670 367 676 1633
rect 630 355 676 367
rect 1088 1633 1134 1645
rect 1088 367 1094 1633
rect 1128 367 1134 1633
rect 1088 355 1134 367
rect 1546 1633 1592 1645
rect 1546 367 1552 1633
rect 1586 367 1592 1633
rect 1546 355 1592 367
rect 2004 1633 2050 1645
rect 2004 367 2010 1633
rect 2044 367 2050 1633
rect 2004 355 2050 367
rect 2462 1633 2508 1645
rect 2462 367 2468 1633
rect 2502 367 2508 1633
rect 2462 355 2508 367
rect 2920 1633 2966 1645
rect 2920 367 2926 1633
rect 2960 367 2966 1633
rect 2920 355 2966 367
rect 3378 1633 3424 1645
rect 3378 367 3384 1633
rect 3418 367 3424 1633
rect 3378 355 3424 367
rect 3836 1633 3882 1645
rect 3836 367 3842 1633
rect 3876 367 3882 1633
rect 3836 355 3882 367
rect 4294 1633 4340 1645
rect 4294 367 4300 1633
rect 4334 367 4340 1633
rect 4294 355 4340 367
rect 130 30 4382 60
rect 130 -30 300 30
rect 360 -30 700 30
rect 760 -30 1100 30
rect 1160 -30 1500 30
rect 1560 -30 1900 30
rect 1960 -30 2300 30
rect 2360 -30 2700 30
rect 2760 -30 3100 30
rect 3160 -30 3500 30
rect 3560 -30 3900 30
rect 3960 -30 4382 30
rect 130 -60 4382 -30
<< labels >>
flabel metal1 130 1850 190 1910 1 FreeSans 480 0 0 0 VPWR
port 4 n power bidirectional
flabel space 120 1850 180 1910 1 FreeSans 480 0 0 0 VPB
flabel metal1 130 -30 190 30 1 FreeSans 480 0 0 0 VGND
port 5 n ground bidirectional
flabel locali 4322 1730 4382 1790 1 FreeSans 480 0 0 0 SOURCE
port 2 n signal bidirectional
flabel locali 4322 210 4382 270 1 FreeSans 480 0 0 0 DRAIN
port 3 n signal bidirectional
flabel locali 4322 102 4382 162 1 FreeSans 480 0 0 0 GATE
port 1 n signal bidirectional
<< properties >>
string FIXED_BBOX 0 0 4770 1880
string LEFclass CORE
string LEFsite unitasc
<< end >>
