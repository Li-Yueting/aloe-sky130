magic
tech sky130A
magscale 1 2
timestamp 1653530608
<< locali >>
rect 122 1850 292 1910
rect 352 1850 692 1910
rect 752 1850 1092 1910
rect 1152 1850 1492 1910
rect 1552 1850 1892 1910
rect 1952 1850 2292 1910
rect 2352 1850 2692 1910
rect 2752 1850 3092 1910
rect 3152 1850 3492 1910
rect 3552 1850 3892 1910
rect 3952 1850 4292 1910
rect 4352 1850 4692 1910
rect 4752 1850 5092 1910
rect 5152 1850 5492 1910
rect 5552 1850 5892 1910
rect 5952 1850 6292 1910
rect 6352 1850 6692 1910
rect 6752 1850 7092 1910
rect 7152 1850 7290 1910
rect 122 -30 292 30
rect 352 -30 692 30
rect 752 -30 1092 30
rect 1152 -30 1492 30
rect 1552 -30 1892 30
rect 1952 -30 2292 30
rect 2352 -30 2692 30
rect 2752 -30 3092 30
rect 3152 -30 3492 30
rect 3552 -30 3892 30
rect 3952 -30 4292 30
rect 4352 -30 4692 30
rect 4752 -30 5092 30
rect 5152 -30 5492 30
rect 5552 -30 5892 30
rect 5952 -30 6292 30
rect 6352 -30 6692 30
rect 6752 -30 7092 30
rect 7152 -30 7290 30
<< viali >>
rect 292 1850 352 1910
rect 692 1850 752 1910
rect 1092 1850 1152 1910
rect 1492 1850 1552 1910
rect 1892 1850 1952 1910
rect 2292 1850 2352 1910
rect 2692 1850 2752 1910
rect 3092 1850 3152 1910
rect 3492 1850 3552 1910
rect 3892 1850 3952 1910
rect 4292 1850 4352 1910
rect 4692 1850 4752 1910
rect 5092 1850 5152 1910
rect 5492 1850 5552 1910
rect 5892 1850 5952 1910
rect 6292 1850 6352 1910
rect 6692 1850 6752 1910
rect 7092 1850 7152 1910
rect 292 -30 352 30
rect 692 -30 752 30
rect 1092 -30 1152 30
rect 1492 -30 1552 30
rect 1892 -30 1952 30
rect 2292 -30 2352 30
rect 2692 -30 2752 30
rect 3092 -30 3152 30
rect 3492 -30 3552 30
rect 3892 -30 3952 30
rect 4292 -30 4352 30
rect 4692 -30 4752 30
rect 5092 -30 5152 30
rect 5492 -30 5552 30
rect 5892 -30 5952 30
rect 6292 -30 6352 30
rect 6692 -30 6752 30
rect 7092 -30 7152 30
<< metal1 >>
rect 122 1910 7290 1940
rect 122 1850 292 1910
rect 352 1850 692 1910
rect 752 1850 1092 1910
rect 1152 1850 1492 1910
rect 1552 1850 1892 1910
rect 1952 1850 2292 1910
rect 2352 1850 2692 1910
rect 2752 1850 3092 1910
rect 3152 1850 3492 1910
rect 3552 1850 3892 1910
rect 3952 1850 4292 1910
rect 4352 1850 4692 1910
rect 4752 1850 5092 1910
rect 5152 1850 5492 1910
rect 5552 1850 5892 1910
rect 5952 1850 6292 1910
rect 6352 1850 6692 1910
rect 6752 1850 7092 1910
rect 7152 1850 7290 1910
rect 122 1820 7290 1850
rect 122 30 7290 60
rect 122 -30 292 30
rect 352 -30 692 30
rect 752 -30 1092 30
rect 1152 -30 1492 30
rect 1552 -30 1892 30
rect 1952 -30 2292 30
rect 2352 -30 2692 30
rect 2752 -30 3092 30
rect 3152 -30 3492 30
rect 3552 -30 3892 30
rect 3952 -30 4292 30
rect 4352 -30 4692 30
rect 4752 -30 5092 30
rect 5152 -30 5492 30
rect 5552 -30 5892 30
rect 5952 -30 6292 30
rect 6352 -30 6692 30
rect 6752 -30 7092 30
rect 7152 -30 7290 30
rect 122 -60 7290 -30
<< metal2 >>
rect 120 1640 320 1650
rect 120 1580 140 1640
rect 300 1580 320 1640
rect 120 1570 320 1580
rect 142 230 302 240
rect 142 150 162 230
rect 282 150 302 230
rect 142 140 302 150
<< via2 >>
rect 140 1580 300 1640
rect 162 150 282 230
<< metal3 >>
rect 120 1640 7292 1650
rect 120 1580 140 1640
rect 300 1622 7292 1640
rect 300 1580 736 1622
rect 120 1078 736 1580
rect 800 1078 1455 1622
rect 1519 1078 2174 1622
rect 2238 1078 2893 1622
rect 2957 1078 3612 1622
rect 3676 1078 4331 1622
rect 4395 1078 5050 1622
rect 5114 1078 5769 1622
rect 5833 1078 6488 1622
rect 6552 1078 7207 1622
rect 7271 1078 7292 1622
rect 120 922 7292 1078
rect 120 378 736 922
rect 800 378 1455 922
rect 1519 378 2174 922
rect 2238 378 2893 922
rect 2957 378 3612 922
rect 3676 378 4331 922
rect 4395 378 5050 922
rect 5114 378 5769 922
rect 5833 378 6488 922
rect 6552 378 7207 922
rect 7271 378 7292 922
rect 120 350 7292 378
rect 122 240 322 250
rect 122 140 142 240
rect 302 140 322 240
rect 122 130 322 140
<< via3 >>
rect 736 1078 800 1622
rect 1455 1078 1519 1622
rect 2174 1078 2238 1622
rect 2893 1078 2957 1622
rect 3612 1078 3676 1622
rect 4331 1078 4395 1622
rect 5050 1078 5114 1622
rect 5769 1078 5833 1622
rect 6488 1078 6552 1622
rect 7207 1078 7271 1622
rect 736 378 800 922
rect 1455 378 1519 922
rect 2174 378 2238 922
rect 2893 378 2957 922
rect 3612 378 3676 922
rect 4331 378 4395 922
rect 5050 378 5114 922
rect 5769 378 5833 922
rect 6488 378 6552 922
rect 7207 378 7271 922
rect 142 230 302 240
rect 142 150 162 230
rect 162 150 282 230
rect 282 150 302 230
rect 142 140 302 150
<< mimcap >>
rect 221 1510 621 1550
rect 221 1190 261 1510
rect 581 1190 621 1510
rect 221 1150 621 1190
rect 940 1510 1340 1550
rect 940 1190 980 1510
rect 1300 1190 1340 1510
rect 940 1150 1340 1190
rect 1659 1510 2059 1550
rect 1659 1190 1699 1510
rect 2019 1190 2059 1510
rect 1659 1150 2059 1190
rect 2378 1510 2778 1550
rect 2378 1190 2418 1510
rect 2738 1190 2778 1510
rect 2378 1150 2778 1190
rect 3097 1510 3497 1550
rect 3097 1190 3137 1510
rect 3457 1190 3497 1510
rect 3097 1150 3497 1190
rect 3816 1510 4216 1550
rect 3816 1190 3856 1510
rect 4176 1190 4216 1510
rect 3816 1150 4216 1190
rect 4535 1510 4935 1550
rect 4535 1190 4575 1510
rect 4895 1190 4935 1510
rect 4535 1150 4935 1190
rect 5254 1510 5654 1550
rect 5254 1190 5294 1510
rect 5614 1190 5654 1510
rect 5254 1150 5654 1190
rect 5973 1510 6373 1550
rect 5973 1190 6013 1510
rect 6333 1190 6373 1510
rect 5973 1150 6373 1190
rect 6692 1510 7092 1550
rect 6692 1190 6732 1510
rect 7052 1190 7092 1510
rect 6692 1150 7092 1190
rect 221 810 621 850
rect 221 490 261 810
rect 581 490 621 810
rect 221 450 621 490
rect 940 810 1340 850
rect 940 490 980 810
rect 1300 490 1340 810
rect 940 450 1340 490
rect 1659 810 2059 850
rect 1659 490 1699 810
rect 2019 490 2059 810
rect 1659 450 2059 490
rect 2378 810 2778 850
rect 2378 490 2418 810
rect 2738 490 2778 810
rect 2378 450 2778 490
rect 3097 810 3497 850
rect 3097 490 3137 810
rect 3457 490 3497 810
rect 3097 450 3497 490
rect 3816 810 4216 850
rect 3816 490 3856 810
rect 4176 490 4216 810
rect 3816 450 4216 490
rect 4535 810 4935 850
rect 4535 490 4575 810
rect 4895 490 4935 810
rect 4535 450 4935 490
rect 5254 810 5654 850
rect 5254 490 5294 810
rect 5614 490 5654 810
rect 5254 450 5654 490
rect 5973 810 6373 850
rect 5973 490 6013 810
rect 6333 490 6373 810
rect 5973 450 6373 490
rect 6692 810 7092 850
rect 6692 490 6732 810
rect 7052 490 7092 810
rect 6692 450 7092 490
<< mimcapcontact >>
rect 261 1190 581 1510
rect 980 1190 1300 1510
rect 1699 1190 2019 1510
rect 2418 1190 2738 1510
rect 3137 1190 3457 1510
rect 3856 1190 4176 1510
rect 4575 1190 4895 1510
rect 5294 1190 5614 1510
rect 6013 1190 6333 1510
rect 6732 1190 7052 1510
rect 261 490 581 810
rect 980 490 1300 810
rect 1699 490 2019 810
rect 2418 490 2738 810
rect 3137 490 3457 810
rect 3856 490 4176 810
rect 4575 490 4895 810
rect 5294 490 5614 810
rect 6013 490 6333 810
rect 6732 490 7052 810
<< metal4 >>
rect 720 1622 816 1638
rect 260 1511 580 1530
rect 260 1510 582 1511
rect 260 1190 261 1510
rect 581 1190 582 1510
rect 260 1189 582 1190
rect 260 811 580 1189
rect 720 1078 736 1622
rect 800 1078 816 1622
rect 1439 1622 1535 1638
rect 980 1511 1300 1530
rect 979 1510 1301 1511
rect 979 1190 980 1510
rect 1300 1190 1301 1510
rect 979 1189 1301 1190
rect 720 1062 816 1078
rect 720 922 816 938
rect 260 810 582 811
rect 260 490 261 810
rect 581 490 582 810
rect 260 489 582 490
rect 260 250 580 489
rect 720 378 736 922
rect 800 378 816 922
rect 980 811 1300 1189
rect 1439 1078 1455 1622
rect 1519 1078 1535 1622
rect 2158 1622 2254 1638
rect 1700 1511 2020 1530
rect 1698 1510 2020 1511
rect 1698 1190 1699 1510
rect 2019 1190 2020 1510
rect 1698 1189 2020 1190
rect 1439 1062 1535 1078
rect 1439 922 1535 938
rect 979 810 1301 811
rect 979 490 980 810
rect 1300 490 1301 810
rect 979 489 1301 490
rect 720 362 816 378
rect 980 250 1300 489
rect 1439 378 1455 922
rect 1519 378 1535 922
rect 1700 811 2020 1189
rect 2158 1078 2174 1622
rect 2238 1078 2254 1622
rect 2877 1622 2973 1638
rect 2420 1511 2740 1530
rect 2417 1510 2740 1511
rect 2417 1190 2418 1510
rect 2738 1190 2740 1510
rect 2417 1189 2740 1190
rect 2158 1062 2254 1078
rect 1698 810 2020 811
rect 1698 490 1699 810
rect 2019 490 2020 810
rect 1698 489 2020 490
rect 1439 362 1535 378
rect 1700 250 2020 489
rect 2158 922 2254 938
rect 2158 378 2174 922
rect 2238 378 2254 922
rect 2420 811 2740 1189
rect 2877 1078 2893 1622
rect 2957 1078 2973 1622
rect 3596 1622 3692 1638
rect 3140 1511 3460 1530
rect 3136 1510 3460 1511
rect 3136 1190 3137 1510
rect 3457 1190 3460 1510
rect 3136 1189 3460 1190
rect 2877 1062 2973 1078
rect 2417 810 2740 811
rect 2417 490 2418 810
rect 2738 490 2740 810
rect 2417 489 2740 490
rect 2158 362 2254 378
rect 2420 250 2740 489
rect 2877 922 2973 938
rect 2877 378 2893 922
rect 2957 378 2973 922
rect 3140 811 3460 1189
rect 3596 1078 3612 1622
rect 3676 1078 3692 1622
rect 4315 1622 4411 1638
rect 3860 1511 4180 1530
rect 3855 1510 4180 1511
rect 3855 1190 3856 1510
rect 4176 1190 4180 1510
rect 3855 1189 4180 1190
rect 3596 1062 3692 1078
rect 3136 810 3460 811
rect 3136 490 3137 810
rect 3457 490 3460 810
rect 3136 489 3460 490
rect 2877 362 2973 378
rect 3140 250 3460 489
rect 3596 922 3692 938
rect 3596 378 3612 922
rect 3676 378 3692 922
rect 3860 811 4180 1189
rect 4315 1078 4331 1622
rect 4395 1078 4411 1622
rect 5034 1622 5130 1638
rect 4580 1511 4900 1530
rect 4574 1510 4900 1511
rect 4574 1190 4575 1510
rect 4895 1190 4900 1510
rect 4574 1189 4900 1190
rect 4315 1062 4411 1078
rect 3855 810 4180 811
rect 3855 490 3856 810
rect 4176 490 4180 810
rect 3855 489 4180 490
rect 3596 362 3692 378
rect 3860 250 4180 489
rect 4315 922 4411 938
rect 4315 378 4331 922
rect 4395 378 4411 922
rect 4580 811 4900 1189
rect 5034 1078 5050 1622
rect 5114 1078 5130 1622
rect 5753 1622 5849 1638
rect 5300 1511 5620 1530
rect 5293 1510 5620 1511
rect 5293 1190 5294 1510
rect 5614 1190 5620 1510
rect 5293 1189 5620 1190
rect 5034 1062 5130 1078
rect 4574 810 4900 811
rect 4574 490 4575 810
rect 4895 490 4900 810
rect 4574 489 4900 490
rect 4315 362 4411 378
rect 4580 250 4900 489
rect 5034 922 5130 938
rect 5034 378 5050 922
rect 5114 378 5130 922
rect 5300 811 5620 1189
rect 5753 1078 5769 1622
rect 5833 1078 5849 1622
rect 6472 1622 6568 1638
rect 6020 1511 6340 1530
rect 6012 1510 6340 1511
rect 6012 1190 6013 1510
rect 6333 1190 6340 1510
rect 6012 1189 6340 1190
rect 5753 1062 5849 1078
rect 5293 810 5620 811
rect 5293 490 5294 810
rect 5614 490 5620 810
rect 5293 489 5620 490
rect 5034 362 5130 378
rect 5300 250 5620 489
rect 5753 922 5849 938
rect 5753 378 5769 922
rect 5833 378 5849 922
rect 6020 811 6340 1189
rect 6472 1078 6488 1622
rect 6552 1078 6568 1622
rect 7191 1622 7287 1638
rect 6740 1511 7060 1530
rect 6731 1510 7060 1511
rect 6731 1190 6732 1510
rect 7052 1190 7060 1510
rect 6731 1189 7060 1190
rect 6472 1062 6568 1078
rect 6012 810 6340 811
rect 6012 490 6013 810
rect 6333 490 6340 810
rect 6012 489 6340 490
rect 5753 362 5849 378
rect 6020 250 6340 489
rect 6472 922 6568 938
rect 6472 378 6488 922
rect 6552 378 6568 922
rect 6740 811 7060 1189
rect 7191 1078 7207 1622
rect 7271 1078 7287 1622
rect 7191 1062 7287 1078
rect 6731 810 7060 811
rect 6731 490 6732 810
rect 7052 490 7060 810
rect 6731 489 7060 490
rect 6472 362 6568 378
rect 6740 250 7060 489
rect 7191 922 7287 938
rect 7191 378 7207 922
rect 7271 378 7287 922
rect 7191 362 7287 378
rect 122 240 7290 250
rect 122 140 142 240
rect 302 140 7290 240
rect 122 130 7290 140
<< labels >>
flabel metal2 120 1570 320 1650 1 FreeSans 800 0 0 0 Cin
port 1 n default bidirectional
flabel metal4 142 140 302 240 1 FreeSans 800 0 0 0 Cout
port 2 n default bidirectional
flabel metal1 122 1850 182 1910 1 FreeSans 800 0 0 0 VPWR
port 3 n power bidirectional
flabel metal1 122 -30 182 30 1 FreeSans 800 0 0 0 VGND
port 4 n ground bidirectional
<< properties >>
string FIXED_BBOX 0 0 7411 1880
string LEFclass CORE
string LEFsite unitasc
<< end >>
