VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO sky130_asc_pfet_01v8_lvt_60
  CLASS CORE ;
  FOREIGN sky130_asc_pfet_01v8_lvt_60 ;
  ORIGIN 0.000 0.000 ;
  SIZE 139.735 BY 9.400 ;
  SITE unitasc ;
  PIN GATE
    DIRECTION INOUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 774.000000 ;
    PORT
      LAYER li1 ;
        RECT 0.650 0.510 138.700 0.810 ;
    END
  END GATE
  PIN SOURCE
    DIRECTION INOUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 56.114998 ;
    PORT
      LAYER li1 ;
        RECT 0.650 8.650 138.700 8.950 ;
        RECT 3.175 8.245 3.345 8.650 ;
        RECT 7.755 8.245 7.925 8.650 ;
        RECT 12.335 8.245 12.505 8.650 ;
        RECT 16.915 8.245 17.085 8.650 ;
        RECT 21.495 8.245 21.665 8.650 ;
        RECT 26.075 8.245 26.245 8.650 ;
        RECT 30.655 8.245 30.825 8.650 ;
        RECT 35.235 8.245 35.405 8.650 ;
        RECT 39.815 8.245 39.985 8.650 ;
        RECT 44.395 8.245 44.565 8.650 ;
        RECT 48.975 8.245 49.145 8.650 ;
        RECT 53.555 8.245 53.725 8.650 ;
        RECT 58.135 8.245 58.305 8.650 ;
        RECT 62.715 8.245 62.885 8.650 ;
        RECT 67.295 8.245 67.465 8.650 ;
        RECT 71.875 8.245 72.045 8.650 ;
        RECT 76.455 8.245 76.625 8.650 ;
        RECT 81.035 8.245 81.205 8.650 ;
        RECT 85.615 8.245 85.785 8.650 ;
        RECT 90.195 8.245 90.365 8.650 ;
        RECT 94.775 8.245 94.945 8.650 ;
        RECT 99.355 8.245 99.525 8.650 ;
        RECT 103.935 8.245 104.105 8.650 ;
        RECT 108.515 8.245 108.685 8.650 ;
        RECT 113.095 8.245 113.265 8.650 ;
        RECT 117.675 8.245 117.845 8.650 ;
        RECT 122.255 8.245 122.425 8.650 ;
        RECT 126.835 8.245 127.005 8.650 ;
        RECT 131.415 8.245 131.585 8.650 ;
        RECT 135.995 8.245 136.165 8.650 ;
        RECT 3.175 8.130 3.355 8.245 ;
        RECT 7.755 8.130 7.935 8.245 ;
        RECT 12.335 8.130 12.515 8.245 ;
        RECT 16.915 8.130 17.095 8.245 ;
        RECT 21.495 8.130 21.675 8.245 ;
        RECT 26.075 8.130 26.255 8.245 ;
        RECT 30.655 8.130 30.835 8.245 ;
        RECT 35.235 8.130 35.415 8.245 ;
        RECT 39.815 8.130 39.995 8.245 ;
        RECT 44.395 8.130 44.575 8.245 ;
        RECT 48.975 8.130 49.155 8.245 ;
        RECT 53.555 8.130 53.735 8.245 ;
        RECT 58.135 8.130 58.315 8.245 ;
        RECT 62.715 8.130 62.895 8.245 ;
        RECT 67.295 8.130 67.475 8.245 ;
        RECT 71.875 8.130 72.055 8.245 ;
        RECT 76.455 8.130 76.635 8.245 ;
        RECT 81.035 8.130 81.215 8.245 ;
        RECT 85.615 8.130 85.795 8.245 ;
        RECT 90.195 8.130 90.375 8.245 ;
        RECT 94.775 8.130 94.955 8.245 ;
        RECT 99.355 8.130 99.535 8.245 ;
        RECT 103.935 8.130 104.115 8.245 ;
        RECT 108.515 8.130 108.695 8.245 ;
        RECT 113.095 8.130 113.275 8.245 ;
        RECT 117.675 8.130 117.855 8.245 ;
        RECT 122.255 8.130 122.435 8.245 ;
        RECT 126.835 8.130 127.015 8.245 ;
        RECT 131.415 8.130 131.595 8.245 ;
        RECT 135.995 8.130 136.175 8.245 ;
        RECT 3.185 1.755 3.355 8.130 ;
        RECT 7.765 1.755 7.935 8.130 ;
        RECT 12.345 1.755 12.515 8.130 ;
        RECT 16.925 1.755 17.095 8.130 ;
        RECT 21.505 1.755 21.675 8.130 ;
        RECT 26.085 1.755 26.255 8.130 ;
        RECT 30.665 1.755 30.835 8.130 ;
        RECT 35.245 1.755 35.415 8.130 ;
        RECT 39.825 1.755 39.995 8.130 ;
        RECT 44.405 1.755 44.575 8.130 ;
        RECT 48.985 1.755 49.155 8.130 ;
        RECT 53.565 1.755 53.735 8.130 ;
        RECT 58.145 1.755 58.315 8.130 ;
        RECT 62.725 1.755 62.895 8.130 ;
        RECT 67.305 1.755 67.475 8.130 ;
        RECT 71.885 1.755 72.055 8.130 ;
        RECT 76.465 1.755 76.635 8.130 ;
        RECT 81.045 1.755 81.215 8.130 ;
        RECT 85.625 1.755 85.795 8.130 ;
        RECT 90.205 1.755 90.375 8.130 ;
        RECT 94.785 1.755 94.955 8.130 ;
        RECT 99.365 1.755 99.535 8.130 ;
        RECT 103.945 1.755 104.115 8.130 ;
        RECT 108.525 1.755 108.695 8.130 ;
        RECT 113.105 1.755 113.275 8.130 ;
        RECT 117.685 1.755 117.855 8.130 ;
        RECT 122.265 1.755 122.435 8.130 ;
        RECT 126.845 1.755 127.015 8.130 ;
        RECT 131.425 1.755 131.595 8.130 ;
        RECT 136.005 1.755 136.175 8.130 ;
      LAYER mcon ;
        RECT 3.185 1.835 3.355 8.165 ;
        RECT 7.765 1.835 7.935 8.165 ;
        RECT 12.345 1.835 12.515 8.165 ;
        RECT 16.925 1.835 17.095 8.165 ;
        RECT 21.505 1.835 21.675 8.165 ;
        RECT 26.085 1.835 26.255 8.165 ;
        RECT 30.665 1.835 30.835 8.165 ;
        RECT 35.245 1.835 35.415 8.165 ;
        RECT 39.825 1.835 39.995 8.165 ;
        RECT 44.405 1.835 44.575 8.165 ;
        RECT 48.985 1.835 49.155 8.165 ;
        RECT 53.565 1.835 53.735 8.165 ;
        RECT 58.145 1.835 58.315 8.165 ;
        RECT 62.725 1.835 62.895 8.165 ;
        RECT 67.305 1.835 67.475 8.165 ;
        RECT 71.885 1.835 72.055 8.165 ;
        RECT 76.465 1.835 76.635 8.165 ;
        RECT 81.045 1.835 81.215 8.165 ;
        RECT 85.625 1.835 85.795 8.165 ;
        RECT 90.205 1.835 90.375 8.165 ;
        RECT 94.785 1.835 94.955 8.165 ;
        RECT 99.365 1.835 99.535 8.165 ;
        RECT 103.945 1.835 104.115 8.165 ;
        RECT 108.525 1.835 108.695 8.165 ;
        RECT 113.105 1.835 113.275 8.165 ;
        RECT 117.685 1.835 117.855 8.165 ;
        RECT 122.265 1.835 122.435 8.165 ;
        RECT 126.845 1.835 127.015 8.165 ;
        RECT 131.425 1.835 131.595 8.165 ;
        RECT 136.005 1.835 136.175 8.165 ;
      LAYER met1 ;
        RECT 3.155 1.775 3.385 8.225 ;
        RECT 7.735 1.775 7.965 8.225 ;
        RECT 12.315 1.775 12.545 8.225 ;
        RECT 16.895 1.775 17.125 8.225 ;
        RECT 21.475 1.775 21.705 8.225 ;
        RECT 26.055 1.775 26.285 8.225 ;
        RECT 30.635 1.775 30.865 8.225 ;
        RECT 35.215 1.775 35.445 8.225 ;
        RECT 39.795 1.775 40.025 8.225 ;
        RECT 44.375 1.775 44.605 8.225 ;
        RECT 48.955 1.775 49.185 8.225 ;
        RECT 53.535 1.775 53.765 8.225 ;
        RECT 58.115 1.775 58.345 8.225 ;
        RECT 62.695 1.775 62.925 8.225 ;
        RECT 67.275 1.775 67.505 8.225 ;
        RECT 71.855 1.775 72.085 8.225 ;
        RECT 76.435 1.775 76.665 8.225 ;
        RECT 81.015 1.775 81.245 8.225 ;
        RECT 85.595 1.775 85.825 8.225 ;
        RECT 90.175 1.775 90.405 8.225 ;
        RECT 94.755 1.775 94.985 8.225 ;
        RECT 99.335 1.775 99.565 8.225 ;
        RECT 103.915 1.775 104.145 8.225 ;
        RECT 108.495 1.775 108.725 8.225 ;
        RECT 113.075 1.775 113.305 8.225 ;
        RECT 117.655 1.775 117.885 8.225 ;
        RECT 122.235 1.775 122.465 8.225 ;
        RECT 126.815 1.775 127.045 8.225 ;
        RECT 131.395 1.775 131.625 8.225 ;
        RECT 135.975 1.775 136.205 8.225 ;
    END
  END SOURCE
  PIN DRAIN
    DIRECTION INOUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 57.985500 ;
    PORT
      LAYER li1 ;
        RECT 0.895 1.860 1.065 8.245 ;
        RECT 5.475 1.860 5.645 8.245 ;
        RECT 10.055 1.860 10.225 8.245 ;
        RECT 14.635 1.860 14.805 8.245 ;
        RECT 19.215 1.860 19.385 8.245 ;
        RECT 23.795 1.860 23.965 8.245 ;
        RECT 28.375 1.860 28.545 8.245 ;
        RECT 32.955 1.860 33.125 8.245 ;
        RECT 37.535 1.860 37.705 8.245 ;
        RECT 42.115 1.860 42.285 8.245 ;
        RECT 46.695 1.860 46.865 8.245 ;
        RECT 51.275 1.860 51.445 8.245 ;
        RECT 55.855 1.860 56.025 8.245 ;
        RECT 60.435 1.860 60.605 8.245 ;
        RECT 65.015 1.860 65.185 8.245 ;
        RECT 69.595 1.860 69.765 8.245 ;
        RECT 74.175 1.860 74.345 8.245 ;
        RECT 78.755 1.860 78.925 8.245 ;
        RECT 83.335 1.860 83.505 8.245 ;
        RECT 87.915 1.860 88.085 8.245 ;
        RECT 92.495 1.860 92.665 8.245 ;
        RECT 97.075 1.860 97.245 8.245 ;
        RECT 101.655 1.860 101.825 8.245 ;
        RECT 106.235 1.860 106.405 8.245 ;
        RECT 110.815 1.860 110.985 8.245 ;
        RECT 115.395 1.860 115.565 8.245 ;
        RECT 119.975 1.860 120.145 8.245 ;
        RECT 124.555 1.860 124.725 8.245 ;
        RECT 129.135 1.860 129.305 8.245 ;
        RECT 133.715 1.860 133.885 8.245 ;
        RECT 138.295 1.860 138.465 8.245 ;
        RECT 0.885 1.755 1.065 1.860 ;
        RECT 5.465 1.755 5.645 1.860 ;
        RECT 10.045 1.755 10.225 1.860 ;
        RECT 14.625 1.755 14.805 1.860 ;
        RECT 19.205 1.755 19.385 1.860 ;
        RECT 23.785 1.755 23.965 1.860 ;
        RECT 28.365 1.755 28.545 1.860 ;
        RECT 32.945 1.755 33.125 1.860 ;
        RECT 37.525 1.755 37.705 1.860 ;
        RECT 42.105 1.755 42.285 1.860 ;
        RECT 46.685 1.755 46.865 1.860 ;
        RECT 51.265 1.755 51.445 1.860 ;
        RECT 55.845 1.755 56.025 1.860 ;
        RECT 60.425 1.755 60.605 1.860 ;
        RECT 65.005 1.755 65.185 1.860 ;
        RECT 69.585 1.755 69.765 1.860 ;
        RECT 74.165 1.755 74.345 1.860 ;
        RECT 78.745 1.755 78.925 1.860 ;
        RECT 83.325 1.755 83.505 1.860 ;
        RECT 87.905 1.755 88.085 1.860 ;
        RECT 92.485 1.755 92.665 1.860 ;
        RECT 97.065 1.755 97.245 1.860 ;
        RECT 101.645 1.755 101.825 1.860 ;
        RECT 106.225 1.755 106.405 1.860 ;
        RECT 110.805 1.755 110.985 1.860 ;
        RECT 115.385 1.755 115.565 1.860 ;
        RECT 119.965 1.755 120.145 1.860 ;
        RECT 124.545 1.755 124.725 1.860 ;
        RECT 129.125 1.755 129.305 1.860 ;
        RECT 133.705 1.755 133.885 1.860 ;
        RECT 138.285 1.755 138.465 1.860 ;
        RECT 0.885 1.350 1.055 1.755 ;
        RECT 5.465 1.350 5.635 1.755 ;
        RECT 10.045 1.350 10.215 1.755 ;
        RECT 14.625 1.350 14.795 1.755 ;
        RECT 19.205 1.350 19.375 1.755 ;
        RECT 23.785 1.350 23.955 1.755 ;
        RECT 28.365 1.350 28.535 1.755 ;
        RECT 32.945 1.350 33.115 1.755 ;
        RECT 37.525 1.350 37.695 1.755 ;
        RECT 42.105 1.350 42.275 1.755 ;
        RECT 46.685 1.350 46.855 1.755 ;
        RECT 51.265 1.350 51.435 1.755 ;
        RECT 55.845 1.350 56.015 1.755 ;
        RECT 60.425 1.350 60.595 1.755 ;
        RECT 65.005 1.350 65.175 1.755 ;
        RECT 69.585 1.350 69.755 1.755 ;
        RECT 74.165 1.350 74.335 1.755 ;
        RECT 78.745 1.350 78.915 1.755 ;
        RECT 83.325 1.350 83.495 1.755 ;
        RECT 87.905 1.350 88.075 1.755 ;
        RECT 92.485 1.350 92.655 1.755 ;
        RECT 97.065 1.350 97.235 1.755 ;
        RECT 101.645 1.350 101.815 1.755 ;
        RECT 106.225 1.350 106.395 1.755 ;
        RECT 110.805 1.350 110.975 1.755 ;
        RECT 115.385 1.350 115.555 1.755 ;
        RECT 119.965 1.350 120.135 1.755 ;
        RECT 124.545 1.350 124.715 1.755 ;
        RECT 129.125 1.350 129.295 1.755 ;
        RECT 133.705 1.350 133.875 1.755 ;
        RECT 138.285 1.350 138.455 1.755 ;
        RECT 0.650 1.050 138.700 1.350 ;
      LAYER mcon ;
        RECT 0.895 1.835 1.065 8.165 ;
        RECT 5.475 1.835 5.645 8.165 ;
        RECT 10.055 1.835 10.225 8.165 ;
        RECT 14.635 1.835 14.805 8.165 ;
        RECT 19.215 1.835 19.385 8.165 ;
        RECT 23.795 1.835 23.965 8.165 ;
        RECT 28.375 1.835 28.545 8.165 ;
        RECT 32.955 1.835 33.125 8.165 ;
        RECT 37.535 1.835 37.705 8.165 ;
        RECT 42.115 1.835 42.285 8.165 ;
        RECT 46.695 1.835 46.865 8.165 ;
        RECT 51.275 1.835 51.445 8.165 ;
        RECT 55.855 1.835 56.025 8.165 ;
        RECT 60.435 1.835 60.605 8.165 ;
        RECT 65.015 1.835 65.185 8.165 ;
        RECT 69.595 1.835 69.765 8.165 ;
        RECT 74.175 1.835 74.345 8.165 ;
        RECT 78.755 1.835 78.925 8.165 ;
        RECT 83.335 1.835 83.505 8.165 ;
        RECT 87.915 1.835 88.085 8.165 ;
        RECT 92.495 1.835 92.665 8.165 ;
        RECT 97.075 1.835 97.245 8.165 ;
        RECT 101.655 1.835 101.825 8.165 ;
        RECT 106.235 1.835 106.405 8.165 ;
        RECT 110.815 1.835 110.985 8.165 ;
        RECT 115.395 1.835 115.565 8.165 ;
        RECT 119.975 1.835 120.145 8.165 ;
        RECT 124.555 1.835 124.725 8.165 ;
        RECT 129.135 1.835 129.305 8.165 ;
        RECT 133.715 1.835 133.885 8.165 ;
        RECT 138.295 1.835 138.465 8.165 ;
      LAYER met1 ;
        RECT 0.865 1.775 1.095 8.225 ;
        RECT 5.445 1.775 5.675 8.225 ;
        RECT 10.025 1.775 10.255 8.225 ;
        RECT 14.605 1.775 14.835 8.225 ;
        RECT 19.185 1.775 19.415 8.225 ;
        RECT 23.765 1.775 23.995 8.225 ;
        RECT 28.345 1.775 28.575 8.225 ;
        RECT 32.925 1.775 33.155 8.225 ;
        RECT 37.505 1.775 37.735 8.225 ;
        RECT 42.085 1.775 42.315 8.225 ;
        RECT 46.665 1.775 46.895 8.225 ;
        RECT 51.245 1.775 51.475 8.225 ;
        RECT 55.825 1.775 56.055 8.225 ;
        RECT 60.405 1.775 60.635 8.225 ;
        RECT 64.985 1.775 65.215 8.225 ;
        RECT 69.565 1.775 69.795 8.225 ;
        RECT 74.145 1.775 74.375 8.225 ;
        RECT 78.725 1.775 78.955 8.225 ;
        RECT 83.305 1.775 83.535 8.225 ;
        RECT 87.885 1.775 88.115 8.225 ;
        RECT 92.465 1.775 92.695 8.225 ;
        RECT 97.045 1.775 97.275 8.225 ;
        RECT 101.625 1.775 101.855 8.225 ;
        RECT 106.205 1.775 106.435 8.225 ;
        RECT 110.785 1.775 111.015 8.225 ;
        RECT 115.365 1.775 115.595 8.225 ;
        RECT 119.945 1.775 120.175 8.225 ;
        RECT 124.525 1.775 124.755 8.225 ;
        RECT 129.105 1.775 129.335 8.225 ;
        RECT 133.685 1.775 133.915 8.225 ;
        RECT 138.265 1.775 138.495 8.225 ;
    END
  END DRAIN
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER li1 ;
        RECT 0.650 9.250 138.700 9.550 ;
      LAYER mcon ;
        RECT 1.500 9.250 1.800 9.550 ;
        RECT 3.500 9.250 3.800 9.550 ;
        RECT 5.500 9.250 5.800 9.550 ;
        RECT 7.500 9.250 7.800 9.550 ;
        RECT 9.500 9.250 9.800 9.550 ;
        RECT 11.500 9.250 11.800 9.550 ;
        RECT 13.500 9.250 13.800 9.550 ;
        RECT 15.500 9.250 15.800 9.550 ;
        RECT 17.500 9.250 17.800 9.550 ;
        RECT 19.500 9.250 19.800 9.550 ;
        RECT 21.500 9.250 21.800 9.550 ;
        RECT 23.500 9.250 23.800 9.550 ;
        RECT 25.500 9.250 25.800 9.550 ;
        RECT 27.500 9.250 27.800 9.550 ;
        RECT 29.500 9.250 29.800 9.550 ;
        RECT 31.500 9.250 31.800 9.550 ;
        RECT 33.500 9.250 33.800 9.550 ;
        RECT 35.500 9.250 35.800 9.550 ;
        RECT 37.500 9.250 37.800 9.550 ;
        RECT 39.500 9.250 39.800 9.550 ;
        RECT 41.500 9.250 41.800 9.550 ;
        RECT 43.500 9.250 43.800 9.550 ;
        RECT 45.500 9.250 45.800 9.550 ;
        RECT 47.500 9.250 47.800 9.550 ;
        RECT 49.500 9.250 49.800 9.550 ;
        RECT 51.500 9.250 51.800 9.550 ;
        RECT 53.500 9.250 53.800 9.550 ;
        RECT 55.500 9.250 55.800 9.550 ;
        RECT 57.500 9.250 57.800 9.550 ;
        RECT 59.500 9.250 59.800 9.550 ;
        RECT 61.500 9.250 61.800 9.550 ;
        RECT 63.500 9.250 63.800 9.550 ;
        RECT 65.500 9.250 65.800 9.550 ;
        RECT 67.500 9.250 67.800 9.550 ;
        RECT 69.500 9.250 69.800 9.550 ;
        RECT 71.500 9.250 71.800 9.550 ;
        RECT 73.500 9.250 73.800 9.550 ;
        RECT 75.500 9.250 75.800 9.550 ;
        RECT 77.500 9.250 77.800 9.550 ;
        RECT 79.500 9.250 79.800 9.550 ;
        RECT 81.500 9.250 81.800 9.550 ;
        RECT 83.500 9.250 83.800 9.550 ;
        RECT 85.500 9.250 85.800 9.550 ;
        RECT 87.500 9.250 87.800 9.550 ;
        RECT 89.500 9.250 89.800 9.550 ;
        RECT 91.500 9.250 91.800 9.550 ;
        RECT 93.500 9.250 93.800 9.550 ;
        RECT 95.500 9.250 95.800 9.550 ;
        RECT 97.500 9.250 97.800 9.550 ;
        RECT 99.500 9.250 99.800 9.550 ;
        RECT 101.500 9.250 101.800 9.550 ;
        RECT 103.500 9.250 103.800 9.550 ;
        RECT 105.500 9.250 105.800 9.550 ;
        RECT 107.500 9.250 107.800 9.550 ;
        RECT 109.500 9.250 109.800 9.550 ;
        RECT 111.500 9.250 111.800 9.550 ;
        RECT 113.500 9.250 113.800 9.550 ;
        RECT 115.500 9.250 115.800 9.550 ;
        RECT 117.500 9.250 117.800 9.550 ;
        RECT 119.500 9.250 119.800 9.550 ;
        RECT 121.500 9.250 121.800 9.550 ;
        RECT 123.500 9.250 123.800 9.550 ;
        RECT 125.500 9.250 125.800 9.550 ;
        RECT 127.500 9.250 127.800 9.550 ;
        RECT 129.500 9.250 129.800 9.550 ;
        RECT 131.500 9.250 131.800 9.550 ;
        RECT 133.500 9.250 133.800 9.550 ;
        RECT 135.500 9.250 135.800 9.550 ;
        RECT 137.500 9.250 137.800 9.550 ;
      LAYER met1 ;
        RECT 0.650 9.100 138.700 9.700 ;
    END
  END VPWR
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER li1 ;
        RECT 0.650 -0.150 138.700 0.150 ;
      LAYER mcon ;
        RECT 1.500 -0.150 1.800 0.150 ;
        RECT 3.500 -0.150 3.800 0.150 ;
        RECT 5.500 -0.150 5.800 0.150 ;
        RECT 7.500 -0.150 7.800 0.150 ;
        RECT 9.500 -0.150 9.800 0.150 ;
        RECT 11.500 -0.150 11.800 0.150 ;
        RECT 13.500 -0.150 13.800 0.150 ;
        RECT 15.500 -0.150 15.800 0.150 ;
        RECT 17.500 -0.150 17.800 0.150 ;
        RECT 19.500 -0.150 19.800 0.150 ;
        RECT 21.500 -0.150 21.800 0.150 ;
        RECT 23.500 -0.150 23.800 0.150 ;
        RECT 25.500 -0.150 25.800 0.150 ;
        RECT 27.500 -0.150 27.800 0.150 ;
        RECT 29.500 -0.150 29.800 0.150 ;
        RECT 31.500 -0.150 31.800 0.150 ;
        RECT 33.500 -0.150 33.800 0.150 ;
        RECT 35.500 -0.150 35.800 0.150 ;
        RECT 37.500 -0.150 37.800 0.150 ;
        RECT 39.500 -0.150 39.800 0.150 ;
        RECT 41.500 -0.150 41.800 0.150 ;
        RECT 43.500 -0.150 43.800 0.150 ;
        RECT 45.500 -0.150 45.800 0.150 ;
        RECT 47.500 -0.150 47.800 0.150 ;
        RECT 49.500 -0.150 49.800 0.150 ;
        RECT 51.500 -0.150 51.800 0.150 ;
        RECT 53.500 -0.150 53.800 0.150 ;
        RECT 55.500 -0.150 55.800 0.150 ;
        RECT 57.500 -0.150 57.800 0.150 ;
        RECT 59.500 -0.150 59.800 0.150 ;
        RECT 61.500 -0.150 61.800 0.150 ;
        RECT 63.500 -0.150 63.800 0.150 ;
        RECT 65.500 -0.150 65.800 0.150 ;
        RECT 67.500 -0.150 67.800 0.150 ;
        RECT 69.500 -0.150 69.800 0.150 ;
        RECT 71.500 -0.150 71.800 0.150 ;
        RECT 73.500 -0.150 73.800 0.150 ;
        RECT 75.500 -0.150 75.800 0.150 ;
        RECT 77.500 -0.150 77.800 0.150 ;
        RECT 79.500 -0.150 79.800 0.150 ;
        RECT 81.500 -0.150 81.800 0.150 ;
        RECT 83.500 -0.150 83.800 0.150 ;
        RECT 85.500 -0.150 85.800 0.150 ;
        RECT 87.500 -0.150 87.800 0.150 ;
        RECT 89.500 -0.150 89.800 0.150 ;
        RECT 91.500 -0.150 91.800 0.150 ;
        RECT 93.500 -0.150 93.800 0.150 ;
        RECT 95.500 -0.150 95.800 0.150 ;
        RECT 97.500 -0.150 97.800 0.150 ;
        RECT 99.500 -0.150 99.800 0.150 ;
        RECT 101.500 -0.150 101.800 0.150 ;
        RECT 103.500 -0.150 103.800 0.150 ;
        RECT 105.500 -0.150 105.800 0.150 ;
        RECT 107.500 -0.150 107.800 0.150 ;
        RECT 109.500 -0.150 109.800 0.150 ;
        RECT 111.500 -0.150 111.800 0.150 ;
        RECT 113.500 -0.150 113.800 0.150 ;
        RECT 115.500 -0.150 115.800 0.150 ;
        RECT 117.500 -0.150 117.800 0.150 ;
        RECT 119.500 -0.150 119.800 0.150 ;
        RECT 121.500 -0.150 121.800 0.150 ;
        RECT 123.500 -0.150 123.800 0.150 ;
        RECT 125.500 -0.150 125.800 0.150 ;
        RECT 127.500 -0.150 127.800 0.150 ;
        RECT 129.500 -0.150 129.800 0.150 ;
        RECT 131.500 -0.150 131.800 0.150 ;
        RECT 133.500 -0.150 133.800 0.150 ;
        RECT 135.500 -0.150 135.800 0.150 ;
        RECT 137.500 -0.150 137.800 0.150 ;
      LAYER met1 ;
        RECT 0.650 -0.300 138.700 0.300 ;
    END
  END VGND
  OBS
      LAYER nwell ;
        RECT 0.650 8.535 138.700 9.700 ;
        RECT 0.650 5.000 138.705 8.535 ;
        RECT 0.655 1.465 138.705 5.000 ;
  END
END sky130_asc_pfet_01v8_lvt_60
END LIBRARY

