VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO sky130_asc_pfet_01v8_lvt_6
  CLASS CORE ;
  FOREIGN sky130_asc_pfet_01v8_lvt_6 ;
  ORIGIN 0.000 0.000 ;
  SIZE 16.975 BY 9.400 ;
  SITE unitasc ;
  PIN GATE
    DIRECTION INOUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 77.400002 ;
    PORT
      LAYER li1 ;
        RECT 0.650 0.510 15.040 0.810 ;
    END
  END GATE
  PIN SOURCE
    DIRECTION INOUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 5.611500 ;
    PORT
      LAYER li1 ;
        RECT 0.650 8.650 15.040 8.950 ;
        RECT 3.175 8.245 3.345 8.650 ;
        RECT 7.755 8.245 7.925 8.650 ;
        RECT 12.335 8.245 12.505 8.650 ;
        RECT 3.175 8.130 3.355 8.245 ;
        RECT 7.755 8.130 7.935 8.245 ;
        RECT 12.335 8.130 12.515 8.245 ;
        RECT 3.185 1.755 3.355 8.130 ;
        RECT 7.765 1.755 7.935 8.130 ;
        RECT 12.345 1.755 12.515 8.130 ;
      LAYER mcon ;
        RECT 3.185 1.835 3.355 8.165 ;
        RECT 7.765 1.835 7.935 8.165 ;
        RECT 12.345 1.835 12.515 8.165 ;
      LAYER met1 ;
        RECT 3.155 1.775 3.385 8.225 ;
        RECT 7.735 1.775 7.965 8.225 ;
        RECT 12.315 1.775 12.545 8.225 ;
    END
  END SOURCE
  PIN DRAIN
    DIRECTION INOUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 7.482000 ;
    PORT
      LAYER li1 ;
        RECT 0.895 1.860 1.065 8.245 ;
        RECT 5.475 1.860 5.645 8.245 ;
        RECT 10.055 1.860 10.225 8.245 ;
        RECT 14.635 1.860 14.805 8.245 ;
        RECT 0.885 1.755 1.065 1.860 ;
        RECT 5.465 1.755 5.645 1.860 ;
        RECT 10.045 1.755 10.225 1.860 ;
        RECT 14.625 1.755 14.805 1.860 ;
        RECT 0.885 1.350 1.055 1.755 ;
        RECT 5.465 1.350 5.635 1.755 ;
        RECT 10.045 1.350 10.215 1.755 ;
        RECT 14.625 1.350 14.795 1.755 ;
        RECT 0.650 1.050 15.040 1.350 ;
      LAYER mcon ;
        RECT 0.895 1.835 1.065 8.165 ;
        RECT 5.475 1.835 5.645 8.165 ;
        RECT 10.055 1.835 10.225 8.165 ;
        RECT 14.635 1.835 14.805 8.165 ;
      LAYER met1 ;
        RECT 0.865 1.775 1.095 8.225 ;
        RECT 5.445 1.775 5.675 8.225 ;
        RECT 10.025 1.775 10.255 8.225 ;
        RECT 14.605 1.775 14.835 8.225 ;
    END
  END DRAIN
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER li1 ;
        RECT 0.650 9.250 15.040 9.550 ;
      LAYER mcon ;
        RECT 1.500 9.250 1.800 9.550 ;
        RECT 3.500 9.250 3.800 9.550 ;
        RECT 5.500 9.250 5.800 9.550 ;
        RECT 7.500 9.250 7.800 9.550 ;
        RECT 9.500 9.250 9.800 9.550 ;
        RECT 11.500 9.250 11.800 9.550 ;
        RECT 13.500 9.250 13.800 9.550 ;
      LAYER met1 ;
        RECT 0.650 9.100 15.040 9.700 ;
    END
  END VPWR
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER li1 ;
        RECT 0.650 -0.150 15.040 0.150 ;
      LAYER mcon ;
        RECT 1.500 -0.150 1.800 0.150 ;
        RECT 3.500 -0.150 3.800 0.150 ;
        RECT 5.500 -0.150 5.800 0.150 ;
        RECT 7.500 -0.150 7.800 0.150 ;
        RECT 9.500 -0.150 9.800 0.150 ;
        RECT 11.500 -0.150 11.800 0.150 ;
        RECT 13.500 -0.150 13.800 0.150 ;
      LAYER met1 ;
        RECT 0.650 -0.300 15.040 0.300 ;
    END
  END VGND
  OBS
      LAYER nwell ;
        RECT 0.650 8.535 15.040 9.700 ;
        RECT 0.650 5.000 15.045 8.535 ;
        RECT 0.655 1.465 15.045 5.000 ;
  END
END sky130_asc_pfet_01v8_lvt_6
END LIBRARY

