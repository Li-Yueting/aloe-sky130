magic
tech sky130A
magscale 1 2
timestamp 1652136261
<< nwell >>
rect 0 1707 27706 1940
rect 0 294 27707 1707
rect 97 293 27707 294
<< pmoslvt >>
rect 191 355 591 1645
rect 649 355 1049 1645
rect 1107 355 1507 1645
rect 1565 355 1965 1645
rect 2023 355 2423 1645
rect 2481 355 2881 1645
rect 2939 355 3339 1645
rect 3397 355 3797 1645
rect 3855 355 4255 1645
rect 4313 355 4713 1645
rect 4771 355 5171 1645
rect 5229 355 5629 1645
rect 5687 355 6087 1645
rect 6145 355 6545 1645
rect 6603 355 7003 1645
rect 7061 355 7461 1645
rect 7519 355 7919 1645
rect 7977 355 8377 1645
rect 8435 355 8835 1645
rect 8893 355 9293 1645
rect 9351 355 9751 1645
rect 9809 355 10209 1645
rect 10267 355 10667 1645
rect 10725 355 11125 1645
rect 11183 355 11583 1645
rect 11641 355 12041 1645
rect 12099 355 12499 1645
rect 12557 355 12957 1645
rect 13015 355 13415 1645
rect 13473 355 13873 1645
rect 13931 355 14331 1645
rect 14389 355 14789 1645
rect 14847 355 15247 1645
rect 15305 355 15705 1645
rect 15763 355 16163 1645
rect 16221 355 16621 1645
rect 16679 355 17079 1645
rect 17137 355 17537 1645
rect 17595 355 17995 1645
rect 18053 355 18453 1645
rect 18511 355 18911 1645
rect 18969 355 19369 1645
rect 19427 355 19827 1645
rect 19885 355 20285 1645
rect 20343 355 20743 1645
rect 20801 355 21201 1645
rect 21259 355 21659 1645
rect 21717 355 22117 1645
rect 22175 355 22575 1645
rect 22633 355 23033 1645
rect 23091 355 23491 1645
rect 23549 355 23949 1645
rect 24007 355 24407 1645
rect 24465 355 24865 1645
rect 24923 355 25323 1645
rect 25381 355 25781 1645
rect 25839 355 26239 1645
rect 26297 355 26697 1645
rect 26755 355 27155 1645
rect 27213 355 27613 1645
<< pdiff >>
rect 133 1633 191 1645
rect 133 367 145 1633
rect 179 367 191 1633
rect 133 355 191 367
rect 591 1633 649 1645
rect 591 367 603 1633
rect 637 367 649 1633
rect 591 355 649 367
rect 1049 1633 1107 1645
rect 1049 367 1061 1633
rect 1095 367 1107 1633
rect 1049 355 1107 367
rect 1507 1633 1565 1645
rect 1507 367 1519 1633
rect 1553 367 1565 1633
rect 1507 355 1565 367
rect 1965 1633 2023 1645
rect 1965 367 1977 1633
rect 2011 367 2023 1633
rect 1965 355 2023 367
rect 2423 1633 2481 1645
rect 2423 367 2435 1633
rect 2469 367 2481 1633
rect 2423 355 2481 367
rect 2881 1633 2939 1645
rect 2881 367 2893 1633
rect 2927 367 2939 1633
rect 2881 355 2939 367
rect 3339 1633 3397 1645
rect 3339 367 3351 1633
rect 3385 367 3397 1633
rect 3339 355 3397 367
rect 3797 1633 3855 1645
rect 3797 367 3809 1633
rect 3843 367 3855 1633
rect 3797 355 3855 367
rect 4255 1633 4313 1645
rect 4255 367 4267 1633
rect 4301 367 4313 1633
rect 4255 355 4313 367
rect 4713 1633 4771 1645
rect 4713 367 4725 1633
rect 4759 367 4771 1633
rect 4713 355 4771 367
rect 5171 1633 5229 1645
rect 5171 367 5183 1633
rect 5217 367 5229 1633
rect 5171 355 5229 367
rect 5629 1633 5687 1645
rect 5629 367 5641 1633
rect 5675 367 5687 1633
rect 5629 355 5687 367
rect 6087 1633 6145 1645
rect 6087 367 6099 1633
rect 6133 367 6145 1633
rect 6087 355 6145 367
rect 6545 1633 6603 1645
rect 6545 367 6557 1633
rect 6591 367 6603 1633
rect 6545 355 6603 367
rect 7003 1633 7061 1645
rect 7003 367 7015 1633
rect 7049 367 7061 1633
rect 7003 355 7061 367
rect 7461 1633 7519 1645
rect 7461 367 7473 1633
rect 7507 367 7519 1633
rect 7461 355 7519 367
rect 7919 1633 7977 1645
rect 7919 367 7931 1633
rect 7965 367 7977 1633
rect 7919 355 7977 367
rect 8377 1633 8435 1645
rect 8377 367 8389 1633
rect 8423 367 8435 1633
rect 8377 355 8435 367
rect 8835 1633 8893 1645
rect 8835 367 8847 1633
rect 8881 367 8893 1633
rect 8835 355 8893 367
rect 9293 1633 9351 1645
rect 9293 367 9305 1633
rect 9339 367 9351 1633
rect 9293 355 9351 367
rect 9751 1633 9809 1645
rect 9751 367 9763 1633
rect 9797 367 9809 1633
rect 9751 355 9809 367
rect 10209 1633 10267 1645
rect 10209 367 10221 1633
rect 10255 367 10267 1633
rect 10209 355 10267 367
rect 10667 1633 10725 1645
rect 10667 367 10679 1633
rect 10713 367 10725 1633
rect 10667 355 10725 367
rect 11125 1633 11183 1645
rect 11125 367 11137 1633
rect 11171 367 11183 1633
rect 11125 355 11183 367
rect 11583 1633 11641 1645
rect 11583 367 11595 1633
rect 11629 367 11641 1633
rect 11583 355 11641 367
rect 12041 1633 12099 1645
rect 12041 367 12053 1633
rect 12087 367 12099 1633
rect 12041 355 12099 367
rect 12499 1633 12557 1645
rect 12499 367 12511 1633
rect 12545 367 12557 1633
rect 12499 355 12557 367
rect 12957 1633 13015 1645
rect 12957 367 12969 1633
rect 13003 367 13015 1633
rect 12957 355 13015 367
rect 13415 1633 13473 1645
rect 13415 367 13427 1633
rect 13461 367 13473 1633
rect 13415 355 13473 367
rect 13873 1633 13931 1645
rect 13873 367 13885 1633
rect 13919 367 13931 1633
rect 13873 355 13931 367
rect 14331 1633 14389 1645
rect 14331 367 14343 1633
rect 14377 367 14389 1633
rect 14331 355 14389 367
rect 14789 1633 14847 1645
rect 14789 367 14801 1633
rect 14835 367 14847 1633
rect 14789 355 14847 367
rect 15247 1633 15305 1645
rect 15247 367 15259 1633
rect 15293 367 15305 1633
rect 15247 355 15305 367
rect 15705 1633 15763 1645
rect 15705 367 15717 1633
rect 15751 367 15763 1633
rect 15705 355 15763 367
rect 16163 1633 16221 1645
rect 16163 367 16175 1633
rect 16209 367 16221 1633
rect 16163 355 16221 367
rect 16621 1633 16679 1645
rect 16621 367 16633 1633
rect 16667 367 16679 1633
rect 16621 355 16679 367
rect 17079 1633 17137 1645
rect 17079 367 17091 1633
rect 17125 367 17137 1633
rect 17079 355 17137 367
rect 17537 1633 17595 1645
rect 17537 367 17549 1633
rect 17583 367 17595 1633
rect 17537 355 17595 367
rect 17995 1633 18053 1645
rect 17995 367 18007 1633
rect 18041 367 18053 1633
rect 17995 355 18053 367
rect 18453 1633 18511 1645
rect 18453 367 18465 1633
rect 18499 367 18511 1633
rect 18453 355 18511 367
rect 18911 1633 18969 1645
rect 18911 367 18923 1633
rect 18957 367 18969 1633
rect 18911 355 18969 367
rect 19369 1633 19427 1645
rect 19369 367 19381 1633
rect 19415 367 19427 1633
rect 19369 355 19427 367
rect 19827 1633 19885 1645
rect 19827 367 19839 1633
rect 19873 367 19885 1633
rect 19827 355 19885 367
rect 20285 1633 20343 1645
rect 20285 367 20297 1633
rect 20331 367 20343 1633
rect 20285 355 20343 367
rect 20743 1633 20801 1645
rect 20743 367 20755 1633
rect 20789 367 20801 1633
rect 20743 355 20801 367
rect 21201 1633 21259 1645
rect 21201 367 21213 1633
rect 21247 367 21259 1633
rect 21201 355 21259 367
rect 21659 1633 21717 1645
rect 21659 367 21671 1633
rect 21705 367 21717 1633
rect 21659 355 21717 367
rect 22117 1633 22175 1645
rect 22117 367 22129 1633
rect 22163 367 22175 1633
rect 22117 355 22175 367
rect 22575 1633 22633 1645
rect 22575 367 22587 1633
rect 22621 367 22633 1633
rect 22575 355 22633 367
rect 23033 1633 23091 1645
rect 23033 367 23045 1633
rect 23079 367 23091 1633
rect 23033 355 23091 367
rect 23491 1633 23549 1645
rect 23491 367 23503 1633
rect 23537 367 23549 1633
rect 23491 355 23549 367
rect 23949 1633 24007 1645
rect 23949 367 23961 1633
rect 23995 367 24007 1633
rect 23949 355 24007 367
rect 24407 1633 24465 1645
rect 24407 367 24419 1633
rect 24453 367 24465 1633
rect 24407 355 24465 367
rect 24865 1633 24923 1645
rect 24865 367 24877 1633
rect 24911 367 24923 1633
rect 24865 355 24923 367
rect 25323 1633 25381 1645
rect 25323 367 25335 1633
rect 25369 367 25381 1633
rect 25323 355 25381 367
rect 25781 1633 25839 1645
rect 25781 367 25793 1633
rect 25827 367 25839 1633
rect 25781 355 25839 367
rect 26239 1633 26297 1645
rect 26239 367 26251 1633
rect 26285 367 26297 1633
rect 26239 355 26297 367
rect 26697 1633 26755 1645
rect 26697 367 26709 1633
rect 26743 367 26755 1633
rect 26697 355 26755 367
rect 27155 1633 27213 1645
rect 27155 367 27167 1633
rect 27201 367 27213 1633
rect 27155 355 27213 367
rect 27613 1633 27671 1645
rect 27613 367 27625 1633
rect 27659 367 27671 1633
rect 27613 355 27671 367
<< pdiffc >>
rect 145 367 179 1633
rect 603 367 637 1633
rect 1061 367 1095 1633
rect 1519 367 1553 1633
rect 1977 367 2011 1633
rect 2435 367 2469 1633
rect 2893 367 2927 1633
rect 3351 367 3385 1633
rect 3809 367 3843 1633
rect 4267 367 4301 1633
rect 4725 367 4759 1633
rect 5183 367 5217 1633
rect 5641 367 5675 1633
rect 6099 367 6133 1633
rect 6557 367 6591 1633
rect 7015 367 7049 1633
rect 7473 367 7507 1633
rect 7931 367 7965 1633
rect 8389 367 8423 1633
rect 8847 367 8881 1633
rect 9305 367 9339 1633
rect 9763 367 9797 1633
rect 10221 367 10255 1633
rect 10679 367 10713 1633
rect 11137 367 11171 1633
rect 11595 367 11629 1633
rect 12053 367 12087 1633
rect 12511 367 12545 1633
rect 12969 367 13003 1633
rect 13427 367 13461 1633
rect 13885 367 13919 1633
rect 14343 367 14377 1633
rect 14801 367 14835 1633
rect 15259 367 15293 1633
rect 15717 367 15751 1633
rect 16175 367 16209 1633
rect 16633 367 16667 1633
rect 17091 367 17125 1633
rect 17549 367 17583 1633
rect 18007 367 18041 1633
rect 18465 367 18499 1633
rect 18923 367 18957 1633
rect 19381 367 19415 1633
rect 19839 367 19873 1633
rect 20297 367 20331 1633
rect 20755 367 20789 1633
rect 21213 367 21247 1633
rect 21671 367 21705 1633
rect 22129 367 22163 1633
rect 22587 367 22621 1633
rect 23045 367 23079 1633
rect 23503 367 23537 1633
rect 23961 367 23995 1633
rect 24419 367 24453 1633
rect 24877 367 24911 1633
rect 25335 367 25369 1633
rect 25793 367 25827 1633
rect 26251 367 26285 1633
rect 26709 367 26743 1633
rect 27167 367 27201 1633
rect 27625 367 27659 1633
<< nsubdiff >>
rect 38 1760 78 1800
rect 38 1680 78 1720
<< nsubdiffcont >>
rect 38 1720 78 1760
<< poly >>
rect 191 1645 591 1671
rect 649 1645 1049 1671
rect 1107 1645 1507 1671
rect 1565 1645 1965 1671
rect 2023 1645 2423 1671
rect 2481 1645 2881 1671
rect 2939 1645 3339 1671
rect 3397 1645 3797 1671
rect 3855 1645 4255 1671
rect 4313 1645 4713 1671
rect 4771 1645 5171 1671
rect 5229 1645 5629 1671
rect 5687 1645 6087 1671
rect 6145 1645 6545 1671
rect 6603 1645 7003 1671
rect 7061 1645 7461 1671
rect 7519 1645 7919 1671
rect 7977 1645 8377 1671
rect 8435 1645 8835 1671
rect 8893 1645 9293 1671
rect 9351 1645 9751 1671
rect 9809 1645 10209 1671
rect 10267 1645 10667 1671
rect 10725 1645 11125 1671
rect 11183 1645 11583 1671
rect 11641 1645 12041 1671
rect 12099 1645 12499 1671
rect 12557 1645 12957 1671
rect 13015 1645 13415 1671
rect 13473 1645 13873 1671
rect 13931 1645 14331 1671
rect 14389 1645 14789 1671
rect 14847 1645 15247 1671
rect 15305 1645 15705 1671
rect 15763 1645 16163 1671
rect 16221 1645 16621 1671
rect 16679 1645 17079 1671
rect 17137 1645 17537 1671
rect 17595 1645 17995 1671
rect 18053 1645 18453 1671
rect 18511 1645 18911 1671
rect 18969 1645 19369 1671
rect 19427 1645 19827 1671
rect 19885 1645 20285 1671
rect 20343 1645 20743 1671
rect 20801 1645 21201 1671
rect 21259 1645 21659 1671
rect 21717 1645 22117 1671
rect 22175 1645 22575 1671
rect 22633 1645 23033 1671
rect 23091 1645 23491 1671
rect 23549 1645 23949 1671
rect 24007 1645 24407 1671
rect 24465 1645 24865 1671
rect 24923 1645 25323 1671
rect 25381 1645 25781 1671
rect 25839 1645 26239 1671
rect 26297 1645 26697 1671
rect 26755 1645 27155 1671
rect 27213 1645 27613 1671
rect 191 329 591 355
rect 649 329 1049 355
rect 1107 329 1507 355
rect 1565 329 1965 355
rect 2023 329 2423 355
rect 2481 329 2881 355
rect 2939 329 3339 355
rect 3397 329 3797 355
rect 3855 329 4255 355
rect 4313 329 4713 355
rect 4771 329 5171 355
rect 5229 329 5629 355
rect 5687 329 6087 355
rect 6145 329 6545 355
rect 6603 329 7003 355
rect 7061 329 7461 355
rect 7519 329 7919 355
rect 7977 329 8377 355
rect 8435 329 8835 355
rect 8893 329 9293 355
rect 9351 329 9751 355
rect 9809 329 10209 355
rect 10267 329 10667 355
rect 10725 329 11125 355
rect 11183 329 11583 355
rect 11641 329 12041 355
rect 12099 329 12499 355
rect 12557 329 12957 355
rect 13015 329 13415 355
rect 13473 329 13873 355
rect 13931 329 14331 355
rect 14389 329 14789 355
rect 14847 329 15247 355
rect 15305 329 15705 355
rect 15763 329 16163 355
rect 16221 329 16621 355
rect 16679 329 17079 355
rect 17137 329 17537 355
rect 17595 329 17995 355
rect 18053 329 18453 355
rect 18511 329 18911 355
rect 18969 329 19369 355
rect 19427 329 19827 355
rect 19885 329 20285 355
rect 20343 329 20743 355
rect 20801 329 21201 355
rect 21259 329 21659 355
rect 21717 329 22117 355
rect 22175 329 22575 355
rect 22633 329 23033 355
rect 23091 329 23491 355
rect 23549 329 23949 355
rect 24007 329 24407 355
rect 24465 329 24865 355
rect 24923 329 25323 355
rect 25381 329 25781 355
rect 25839 329 26239 355
rect 26297 329 26697 355
rect 26755 329 27155 355
rect 27213 329 27613 355
rect 338 184 458 329
rect 794 184 914 329
rect 1250 184 1370 329
rect 1706 184 1826 329
rect 2162 184 2282 329
rect 2618 184 2738 329
rect 3074 184 3194 329
rect 3530 184 3650 329
rect 3986 184 4106 329
rect 4442 184 4562 329
rect 4898 184 5018 329
rect 5354 184 5474 329
rect 5810 184 5930 329
rect 6266 184 6386 329
rect 6722 184 6842 329
rect 7178 184 7298 329
rect 7634 184 7754 329
rect 8090 184 8210 329
rect 8546 184 8666 329
rect 9002 184 9122 329
rect 9458 184 9578 329
rect 9914 184 10034 329
rect 10370 184 10490 329
rect 10826 184 10946 329
rect 11282 184 11402 329
rect 11738 184 11858 329
rect 12194 184 12314 329
rect 12650 184 12770 329
rect 13106 184 13226 329
rect 13562 184 13682 329
rect 14018 184 14138 329
rect 14474 184 14594 329
rect 14930 184 15050 329
rect 15386 184 15506 329
rect 15842 184 15962 329
rect 16298 184 16418 329
rect 16754 184 16874 329
rect 17210 184 17330 329
rect 17666 184 17786 329
rect 18122 184 18242 329
rect 18578 184 18698 329
rect 19034 184 19154 329
rect 19490 184 19610 329
rect 19946 184 20066 329
rect 20402 184 20522 329
rect 20858 184 20978 329
rect 21314 184 21434 329
rect 21770 184 21890 329
rect 22226 184 22346 329
rect 22682 184 22802 329
rect 23138 184 23258 329
rect 23594 184 23714 329
rect 24050 184 24170 329
rect 24506 184 24626 329
rect 24962 184 25082 329
rect 25418 184 25538 329
rect 25874 184 25994 329
rect 26330 184 26450 329
rect 26786 184 26906 329
rect 27242 184 27362 329
rect 98 164 27706 184
rect 98 104 268 164
rect 328 104 668 164
rect 728 104 1068 164
rect 1128 104 1468 164
rect 1528 104 1868 164
rect 1928 104 2268 164
rect 2328 104 2668 164
rect 2728 104 3068 164
rect 3128 104 3468 164
rect 3528 104 3868 164
rect 3928 104 4268 164
rect 4328 104 4668 164
rect 4728 104 5068 164
rect 5128 104 5468 164
rect 5528 104 5868 164
rect 5928 104 6268 164
rect 6328 104 6668 164
rect 6728 104 7068 164
rect 7128 104 7468 164
rect 7528 104 7868 164
rect 7928 104 8268 164
rect 8328 104 8668 164
rect 8728 104 9068 164
rect 9128 104 9468 164
rect 9528 104 9868 164
rect 9928 104 10268 164
rect 10328 104 10668 164
rect 10728 104 11068 164
rect 11128 104 11468 164
rect 11528 104 11868 164
rect 11928 104 12268 164
rect 12328 104 12668 164
rect 12728 104 13068 164
rect 13128 104 13468 164
rect 13528 104 13868 164
rect 13928 104 14268 164
rect 14328 104 14668 164
rect 14728 104 15068 164
rect 15128 104 15468 164
rect 15528 104 15868 164
rect 15928 104 16268 164
rect 16328 104 16668 164
rect 16728 104 17068 164
rect 17128 104 17468 164
rect 17528 104 17868 164
rect 17928 104 18268 164
rect 18328 104 18668 164
rect 18728 104 19068 164
rect 19128 104 19468 164
rect 19528 104 19868 164
rect 19928 104 20268 164
rect 20328 104 20668 164
rect 20728 104 21068 164
rect 21128 104 21468 164
rect 21528 104 21868 164
rect 21928 104 22268 164
rect 22328 104 22668 164
rect 22728 104 23068 164
rect 23128 104 23468 164
rect 23528 104 23868 164
rect 23928 104 24268 164
rect 24328 104 24668 164
rect 24728 104 25068 164
rect 25128 104 25468 164
rect 25528 104 25868 164
rect 25928 104 26268 164
rect 26328 104 26668 164
rect 26728 104 27068 164
rect 27128 104 27468 164
rect 27528 104 27706 164
rect 98 84 27706 104
<< polycont >>
rect 268 104 328 164
rect 668 104 728 164
rect 1068 104 1128 164
rect 1468 104 1528 164
rect 1868 104 1928 164
rect 2268 104 2328 164
rect 2668 104 2728 164
rect 3068 104 3128 164
rect 3468 104 3528 164
rect 3868 104 3928 164
rect 4268 104 4328 164
rect 4668 104 4728 164
rect 5068 104 5128 164
rect 5468 104 5528 164
rect 5868 104 5928 164
rect 6268 104 6328 164
rect 6668 104 6728 164
rect 7068 104 7128 164
rect 7468 104 7528 164
rect 7868 104 7928 164
rect 8268 104 8328 164
rect 8668 104 8728 164
rect 9068 104 9128 164
rect 9468 104 9528 164
rect 9868 104 9928 164
rect 10268 104 10328 164
rect 10668 104 10728 164
rect 11068 104 11128 164
rect 11468 104 11528 164
rect 11868 104 11928 164
rect 12268 104 12328 164
rect 12668 104 12728 164
rect 13068 104 13128 164
rect 13468 104 13528 164
rect 13868 104 13928 164
rect 14268 104 14328 164
rect 14668 104 14728 164
rect 15068 104 15128 164
rect 15468 104 15528 164
rect 15868 104 15928 164
rect 16268 104 16328 164
rect 16668 104 16728 164
rect 17068 104 17128 164
rect 17468 104 17528 164
rect 17868 104 17928 164
rect 18268 104 18328 164
rect 18668 104 18728 164
rect 19068 104 19128 164
rect 19468 104 19528 164
rect 19868 104 19928 164
rect 20268 104 20328 164
rect 20668 104 20728 164
rect 21068 104 21128 164
rect 21468 104 21528 164
rect 21868 104 21928 164
rect 22268 104 22328 164
rect 22668 104 22728 164
rect 23068 104 23128 164
rect 23468 104 23528 164
rect 23868 104 23928 164
rect 24268 104 24328 164
rect 24668 104 24728 164
rect 25068 104 25128 164
rect 25468 104 25528 164
rect 25868 104 25928 164
rect 26268 104 26328 164
rect 26668 104 26728 164
rect 27068 104 27128 164
rect 27468 104 27528 164
<< locali >>
rect 0 1850 268 1910
rect 328 1850 668 1910
rect 728 1850 1068 1910
rect 1128 1850 1468 1910
rect 1528 1850 1868 1910
rect 1928 1850 2268 1910
rect 2328 1850 2668 1910
rect 2728 1850 3068 1910
rect 3128 1850 3468 1910
rect 3528 1850 3868 1910
rect 3928 1850 4268 1910
rect 4328 1850 4668 1910
rect 4728 1850 5068 1910
rect 5128 1850 5468 1910
rect 5528 1850 5868 1910
rect 5928 1850 6268 1910
rect 6328 1850 6668 1910
rect 6728 1850 7068 1910
rect 7128 1850 7468 1910
rect 7528 1850 7868 1910
rect 7928 1850 8268 1910
rect 8328 1850 8668 1910
rect 8728 1850 9068 1910
rect 9128 1850 9468 1910
rect 9528 1850 9868 1910
rect 9928 1850 10268 1910
rect 10328 1850 10668 1910
rect 10728 1850 11068 1910
rect 11128 1850 11468 1910
rect 11528 1850 11868 1910
rect 11928 1850 12268 1910
rect 12328 1850 12668 1910
rect 12728 1850 13068 1910
rect 13128 1850 13468 1910
rect 13528 1850 13868 1910
rect 13928 1850 14268 1910
rect 14328 1850 14668 1910
rect 14728 1850 15068 1910
rect 15128 1850 15468 1910
rect 15528 1850 15868 1910
rect 15928 1850 16268 1910
rect 16328 1850 16668 1910
rect 16728 1850 17068 1910
rect 17128 1850 17468 1910
rect 17528 1850 17868 1910
rect 17928 1850 18268 1910
rect 18328 1850 18668 1910
rect 18728 1850 19068 1910
rect 19128 1850 19468 1910
rect 19528 1850 19868 1910
rect 19928 1850 20268 1910
rect 20328 1850 20668 1910
rect 20728 1850 21068 1910
rect 21128 1850 21468 1910
rect 21528 1850 21868 1910
rect 21928 1850 22268 1910
rect 22328 1850 22668 1910
rect 22728 1850 23068 1910
rect 23128 1850 23468 1910
rect 23528 1850 23868 1910
rect 23928 1850 24268 1910
rect 24328 1850 24668 1910
rect 24728 1850 25068 1910
rect 25128 1850 25468 1910
rect 25528 1850 25868 1910
rect 25928 1850 26268 1910
rect 26328 1850 26668 1910
rect 26728 1850 27068 1910
rect 27128 1850 27468 1910
rect 27528 1850 27706 1910
rect 28 1760 88 1850
rect 28 1720 38 1760
rect 78 1720 88 1760
rect 158 1730 27706 1790
rect 28 1640 88 1720
rect 145 1633 179 1649
rect 145 270 179 367
rect 603 1633 637 1730
rect 603 351 637 367
rect 1061 1633 1095 1649
rect 1061 270 1095 367
rect 1519 1633 1553 1730
rect 1519 351 1553 367
rect 1977 1633 2011 1649
rect 1977 270 2011 367
rect 2435 1633 2469 1730
rect 2435 351 2469 367
rect 2893 1633 2927 1649
rect 2893 270 2927 367
rect 3351 1633 3385 1730
rect 3351 351 3385 367
rect 3809 1633 3843 1649
rect 3809 270 3843 367
rect 4267 1633 4301 1730
rect 4267 351 4301 367
rect 4725 1633 4759 1649
rect 4725 270 4759 367
rect 5183 1633 5217 1730
rect 5183 351 5217 367
rect 5641 1633 5675 1649
rect 5641 270 5675 367
rect 6099 1633 6133 1730
rect 6099 351 6133 367
rect 6557 1633 6591 1649
rect 6557 270 6591 367
rect 7015 1633 7049 1730
rect 7015 351 7049 367
rect 7473 1633 7507 1649
rect 7473 270 7507 367
rect 7931 1633 7965 1730
rect 7931 351 7965 367
rect 8389 1633 8423 1649
rect 8389 270 8423 367
rect 8847 1633 8881 1730
rect 8847 351 8881 367
rect 9305 1633 9339 1649
rect 9305 270 9339 367
rect 9763 1633 9797 1730
rect 9763 351 9797 367
rect 10221 1633 10255 1649
rect 10221 270 10255 367
rect 10679 1633 10713 1730
rect 10679 351 10713 367
rect 11137 1633 11171 1649
rect 11137 270 11171 367
rect 11595 1633 11629 1730
rect 11595 351 11629 367
rect 12053 1633 12087 1649
rect 12053 270 12087 367
rect 12511 1633 12545 1730
rect 12511 351 12545 367
rect 12969 1633 13003 1649
rect 12969 270 13003 367
rect 13427 1633 13461 1730
rect 13427 351 13461 367
rect 13885 1633 13919 1649
rect 13885 270 13919 367
rect 14343 1633 14377 1730
rect 14343 351 14377 367
rect 14801 1633 14835 1649
rect 14801 270 14835 367
rect 15259 1633 15293 1730
rect 15259 351 15293 367
rect 15717 1633 15751 1649
rect 15717 270 15751 367
rect 16175 1633 16209 1730
rect 16175 351 16209 367
rect 16633 1633 16667 1649
rect 16633 270 16667 367
rect 17091 1633 17125 1730
rect 17091 351 17125 367
rect 17549 1633 17583 1649
rect 17549 270 17583 367
rect 18007 1633 18041 1730
rect 18007 351 18041 367
rect 18465 1633 18499 1649
rect 18465 270 18499 367
rect 18923 1633 18957 1730
rect 18923 351 18957 367
rect 19381 1633 19415 1649
rect 19381 270 19415 367
rect 19839 1633 19873 1730
rect 19839 351 19873 367
rect 20297 1633 20331 1649
rect 20297 270 20331 367
rect 20755 1633 20789 1730
rect 20755 351 20789 367
rect 21213 1633 21247 1649
rect 21213 270 21247 367
rect 21671 1633 21705 1730
rect 21671 351 21705 367
rect 22129 1633 22163 1649
rect 22129 270 22163 367
rect 22587 1633 22621 1730
rect 22587 351 22621 367
rect 23045 1633 23079 1649
rect 23045 270 23079 367
rect 23503 1633 23537 1730
rect 23503 351 23537 367
rect 23961 1633 23995 1649
rect 23961 270 23995 367
rect 24419 1633 24453 1730
rect 24419 351 24453 367
rect 24877 1633 24911 1649
rect 24877 270 24911 367
rect 25335 1633 25369 1730
rect 25335 351 25369 367
rect 25793 1633 25827 1649
rect 25793 270 25827 367
rect 26251 1633 26285 1730
rect 26251 351 26285 367
rect 26709 1633 26743 1649
rect 26709 270 26743 367
rect 27167 1633 27201 1730
rect 27167 351 27201 367
rect 27625 1633 27659 1649
rect 27625 270 27659 367
rect 98 210 27706 270
rect 98 104 268 164
rect 328 104 668 164
rect 728 104 1068 164
rect 1128 104 1468 164
rect 1528 104 1868 164
rect 1928 104 2268 164
rect 2328 104 2668 164
rect 2728 104 3068 164
rect 3128 104 3468 164
rect 3528 104 3868 164
rect 3928 104 4268 164
rect 4328 104 4668 164
rect 4728 104 5068 164
rect 5128 104 5468 164
rect 5528 104 5868 164
rect 5928 104 6268 164
rect 6328 104 6668 164
rect 6728 104 7068 164
rect 7128 104 7468 164
rect 7528 104 7868 164
rect 7928 104 8268 164
rect 8328 104 8668 164
rect 8728 104 9068 164
rect 9128 104 9468 164
rect 9528 104 9868 164
rect 9928 104 10268 164
rect 10328 104 10668 164
rect 10728 104 11068 164
rect 11128 104 11468 164
rect 11528 104 11868 164
rect 11928 104 12268 164
rect 12328 104 12668 164
rect 12728 104 13068 164
rect 13128 104 13468 164
rect 13528 104 13868 164
rect 13928 104 14268 164
rect 14328 104 14668 164
rect 14728 104 15068 164
rect 15128 104 15468 164
rect 15528 104 15868 164
rect 15928 104 16268 164
rect 16328 104 16668 164
rect 16728 104 17068 164
rect 17128 104 17468 164
rect 17528 104 17868 164
rect 17928 104 18268 164
rect 18328 104 18668 164
rect 18728 104 19068 164
rect 19128 104 19468 164
rect 19528 104 19868 164
rect 19928 104 20268 164
rect 20328 104 20668 164
rect 20728 104 21068 164
rect 21128 104 21468 164
rect 21528 104 21868 164
rect 21928 104 22268 164
rect 22328 104 22668 164
rect 22728 104 23068 164
rect 23128 104 23468 164
rect 23528 104 23868 164
rect 23928 104 24268 164
rect 24328 104 24668 164
rect 24728 104 25068 164
rect 25128 104 25468 164
rect 25528 104 25868 164
rect 25928 104 26268 164
rect 26328 104 26668 164
rect 26728 104 27068 164
rect 27128 104 27468 164
rect 27528 104 27706 164
rect 0 -30 268 30
rect 328 -30 668 30
rect 728 -30 1068 30
rect 1128 -30 1468 30
rect 1528 -30 1868 30
rect 1928 -30 2268 30
rect 2328 -30 2668 30
rect 2728 -30 3068 30
rect 3128 -30 3468 30
rect 3528 -30 3868 30
rect 3928 -30 4268 30
rect 4328 -30 4668 30
rect 4728 -30 5068 30
rect 5128 -30 5468 30
rect 5528 -30 5868 30
rect 5928 -30 6268 30
rect 6328 -30 6668 30
rect 6728 -30 7068 30
rect 7128 -30 7468 30
rect 7528 -30 7868 30
rect 7928 -30 8268 30
rect 8328 -30 8668 30
rect 8728 -30 9068 30
rect 9128 -30 9468 30
rect 9528 -30 9868 30
rect 9928 -30 10268 30
rect 10328 -30 10668 30
rect 10728 -30 11068 30
rect 11128 -30 11468 30
rect 11528 -30 11868 30
rect 11928 -30 12268 30
rect 12328 -30 12668 30
rect 12728 -30 13068 30
rect 13128 -30 13468 30
rect 13528 -30 13868 30
rect 13928 -30 14268 30
rect 14328 -30 14668 30
rect 14728 -30 15068 30
rect 15128 -30 15468 30
rect 15528 -30 15868 30
rect 15928 -30 16268 30
rect 16328 -30 16668 30
rect 16728 -30 17068 30
rect 17128 -30 17468 30
rect 17528 -30 17868 30
rect 17928 -30 18268 30
rect 18328 -30 18668 30
rect 18728 -30 19068 30
rect 19128 -30 19468 30
rect 19528 -30 19868 30
rect 19928 -30 20268 30
rect 20328 -30 20668 30
rect 20728 -30 21068 30
rect 21128 -30 21468 30
rect 21528 -30 21868 30
rect 21928 -30 22268 30
rect 22328 -30 22668 30
rect 22728 -30 23068 30
rect 23128 -30 23468 30
rect 23528 -30 23868 30
rect 23928 -30 24268 30
rect 24328 -30 24668 30
rect 24728 -30 25068 30
rect 25128 -30 25468 30
rect 25528 -30 25868 30
rect 25928 -30 26268 30
rect 26328 -30 26668 30
rect 26728 -30 27068 30
rect 27128 -30 27468 30
rect 27528 -30 27706 30
<< viali >>
rect 268 1850 328 1910
rect 668 1850 728 1910
rect 1068 1850 1128 1910
rect 1468 1850 1528 1910
rect 1868 1850 1928 1910
rect 2268 1850 2328 1910
rect 2668 1850 2728 1910
rect 3068 1850 3128 1910
rect 3468 1850 3528 1910
rect 3868 1850 3928 1910
rect 4268 1850 4328 1910
rect 4668 1850 4728 1910
rect 5068 1850 5128 1910
rect 5468 1850 5528 1910
rect 5868 1850 5928 1910
rect 6268 1850 6328 1910
rect 6668 1850 6728 1910
rect 7068 1850 7128 1910
rect 7468 1850 7528 1910
rect 7868 1850 7928 1910
rect 8268 1850 8328 1910
rect 8668 1850 8728 1910
rect 9068 1850 9128 1910
rect 9468 1850 9528 1910
rect 9868 1850 9928 1910
rect 10268 1850 10328 1910
rect 10668 1850 10728 1910
rect 11068 1850 11128 1910
rect 11468 1850 11528 1910
rect 11868 1850 11928 1910
rect 12268 1850 12328 1910
rect 12668 1850 12728 1910
rect 13068 1850 13128 1910
rect 13468 1850 13528 1910
rect 13868 1850 13928 1910
rect 14268 1850 14328 1910
rect 14668 1850 14728 1910
rect 15068 1850 15128 1910
rect 15468 1850 15528 1910
rect 15868 1850 15928 1910
rect 16268 1850 16328 1910
rect 16668 1850 16728 1910
rect 17068 1850 17128 1910
rect 17468 1850 17528 1910
rect 17868 1850 17928 1910
rect 18268 1850 18328 1910
rect 18668 1850 18728 1910
rect 19068 1850 19128 1910
rect 19468 1850 19528 1910
rect 19868 1850 19928 1910
rect 20268 1850 20328 1910
rect 20668 1850 20728 1910
rect 21068 1850 21128 1910
rect 21468 1850 21528 1910
rect 21868 1850 21928 1910
rect 22268 1850 22328 1910
rect 22668 1850 22728 1910
rect 23068 1850 23128 1910
rect 23468 1850 23528 1910
rect 23868 1850 23928 1910
rect 24268 1850 24328 1910
rect 24668 1850 24728 1910
rect 25068 1850 25128 1910
rect 25468 1850 25528 1910
rect 25868 1850 25928 1910
rect 26268 1850 26328 1910
rect 26668 1850 26728 1910
rect 27068 1850 27128 1910
rect 27468 1850 27528 1910
rect 145 367 179 1633
rect 603 367 637 1633
rect 1061 367 1095 1633
rect 1519 367 1553 1633
rect 1977 367 2011 1633
rect 2435 367 2469 1633
rect 2893 367 2927 1633
rect 3351 367 3385 1633
rect 3809 367 3843 1633
rect 4267 367 4301 1633
rect 4725 367 4759 1633
rect 5183 367 5217 1633
rect 5641 367 5675 1633
rect 6099 367 6133 1633
rect 6557 367 6591 1633
rect 7015 367 7049 1633
rect 7473 367 7507 1633
rect 7931 367 7965 1633
rect 8389 367 8423 1633
rect 8847 367 8881 1633
rect 9305 367 9339 1633
rect 9763 367 9797 1633
rect 10221 367 10255 1633
rect 10679 367 10713 1633
rect 11137 367 11171 1633
rect 11595 367 11629 1633
rect 12053 367 12087 1633
rect 12511 367 12545 1633
rect 12969 367 13003 1633
rect 13427 367 13461 1633
rect 13885 367 13919 1633
rect 14343 367 14377 1633
rect 14801 367 14835 1633
rect 15259 367 15293 1633
rect 15717 367 15751 1633
rect 16175 367 16209 1633
rect 16633 367 16667 1633
rect 17091 367 17125 1633
rect 17549 367 17583 1633
rect 18007 367 18041 1633
rect 18465 367 18499 1633
rect 18923 367 18957 1633
rect 19381 367 19415 1633
rect 19839 367 19873 1633
rect 20297 367 20331 1633
rect 20755 367 20789 1633
rect 21213 367 21247 1633
rect 21671 367 21705 1633
rect 22129 367 22163 1633
rect 22587 367 22621 1633
rect 23045 367 23079 1633
rect 23503 367 23537 1633
rect 23961 367 23995 1633
rect 24419 367 24453 1633
rect 24877 367 24911 1633
rect 25335 367 25369 1633
rect 25793 367 25827 1633
rect 26251 367 26285 1633
rect 26709 367 26743 1633
rect 27167 367 27201 1633
rect 27625 367 27659 1633
rect 268 -30 328 30
rect 668 -30 728 30
rect 1068 -30 1128 30
rect 1468 -30 1528 30
rect 1868 -30 1928 30
rect 2268 -30 2328 30
rect 2668 -30 2728 30
rect 3068 -30 3128 30
rect 3468 -30 3528 30
rect 3868 -30 3928 30
rect 4268 -30 4328 30
rect 4668 -30 4728 30
rect 5068 -30 5128 30
rect 5468 -30 5528 30
rect 5868 -30 5928 30
rect 6268 -30 6328 30
rect 6668 -30 6728 30
rect 7068 -30 7128 30
rect 7468 -30 7528 30
rect 7868 -30 7928 30
rect 8268 -30 8328 30
rect 8668 -30 8728 30
rect 9068 -30 9128 30
rect 9468 -30 9528 30
rect 9868 -30 9928 30
rect 10268 -30 10328 30
rect 10668 -30 10728 30
rect 11068 -30 11128 30
rect 11468 -30 11528 30
rect 11868 -30 11928 30
rect 12268 -30 12328 30
rect 12668 -30 12728 30
rect 13068 -30 13128 30
rect 13468 -30 13528 30
rect 13868 -30 13928 30
rect 14268 -30 14328 30
rect 14668 -30 14728 30
rect 15068 -30 15128 30
rect 15468 -30 15528 30
rect 15868 -30 15928 30
rect 16268 -30 16328 30
rect 16668 -30 16728 30
rect 17068 -30 17128 30
rect 17468 -30 17528 30
rect 17868 -30 17928 30
rect 18268 -30 18328 30
rect 18668 -30 18728 30
rect 19068 -30 19128 30
rect 19468 -30 19528 30
rect 19868 -30 19928 30
rect 20268 -30 20328 30
rect 20668 -30 20728 30
rect 21068 -30 21128 30
rect 21468 -30 21528 30
rect 21868 -30 21928 30
rect 22268 -30 22328 30
rect 22668 -30 22728 30
rect 23068 -30 23128 30
rect 23468 -30 23528 30
rect 23868 -30 23928 30
rect 24268 -30 24328 30
rect 24668 -30 24728 30
rect 25068 -30 25128 30
rect 25468 -30 25528 30
rect 25868 -30 25928 30
rect 26268 -30 26328 30
rect 26668 -30 26728 30
rect 27068 -30 27128 30
rect 27468 -30 27528 30
<< metal1 >>
rect 0 1910 27706 1940
rect 0 1850 268 1910
rect 328 1850 668 1910
rect 728 1850 1068 1910
rect 1128 1850 1468 1910
rect 1528 1850 1868 1910
rect 1928 1850 2268 1910
rect 2328 1850 2668 1910
rect 2728 1850 3068 1910
rect 3128 1850 3468 1910
rect 3528 1850 3868 1910
rect 3928 1850 4268 1910
rect 4328 1850 4668 1910
rect 4728 1850 5068 1910
rect 5128 1850 5468 1910
rect 5528 1850 5868 1910
rect 5928 1850 6268 1910
rect 6328 1850 6668 1910
rect 6728 1850 7068 1910
rect 7128 1850 7468 1910
rect 7528 1850 7868 1910
rect 7928 1850 8268 1910
rect 8328 1850 8668 1910
rect 8728 1850 9068 1910
rect 9128 1850 9468 1910
rect 9528 1850 9868 1910
rect 9928 1850 10268 1910
rect 10328 1850 10668 1910
rect 10728 1850 11068 1910
rect 11128 1850 11468 1910
rect 11528 1850 11868 1910
rect 11928 1850 12268 1910
rect 12328 1850 12668 1910
rect 12728 1850 13068 1910
rect 13128 1850 13468 1910
rect 13528 1850 13868 1910
rect 13928 1850 14268 1910
rect 14328 1850 14668 1910
rect 14728 1850 15068 1910
rect 15128 1850 15468 1910
rect 15528 1850 15868 1910
rect 15928 1850 16268 1910
rect 16328 1850 16668 1910
rect 16728 1850 17068 1910
rect 17128 1850 17468 1910
rect 17528 1850 17868 1910
rect 17928 1850 18268 1910
rect 18328 1850 18668 1910
rect 18728 1850 19068 1910
rect 19128 1850 19468 1910
rect 19528 1850 19868 1910
rect 19928 1850 20268 1910
rect 20328 1850 20668 1910
rect 20728 1850 21068 1910
rect 21128 1850 21468 1910
rect 21528 1850 21868 1910
rect 21928 1850 22268 1910
rect 22328 1850 22668 1910
rect 22728 1850 23068 1910
rect 23128 1850 23468 1910
rect 23528 1850 23868 1910
rect 23928 1850 24268 1910
rect 24328 1850 24668 1910
rect 24728 1850 25068 1910
rect 25128 1850 25468 1910
rect 25528 1850 25868 1910
rect 25928 1850 26268 1910
rect 26328 1850 26668 1910
rect 26728 1850 27068 1910
rect 27128 1850 27468 1910
rect 27528 1850 27706 1910
rect 0 1820 27706 1850
rect 139 1633 185 1645
rect 139 367 145 1633
rect 179 367 185 1633
rect 139 355 185 367
rect 597 1633 643 1645
rect 597 367 603 1633
rect 637 367 643 1633
rect 597 355 643 367
rect 1055 1633 1101 1645
rect 1055 367 1061 1633
rect 1095 367 1101 1633
rect 1055 355 1101 367
rect 1513 1633 1559 1645
rect 1513 367 1519 1633
rect 1553 367 1559 1633
rect 1513 355 1559 367
rect 1971 1633 2017 1645
rect 1971 367 1977 1633
rect 2011 367 2017 1633
rect 1971 355 2017 367
rect 2429 1633 2475 1645
rect 2429 367 2435 1633
rect 2469 367 2475 1633
rect 2429 355 2475 367
rect 2887 1633 2933 1645
rect 2887 367 2893 1633
rect 2927 367 2933 1633
rect 2887 355 2933 367
rect 3345 1633 3391 1645
rect 3345 367 3351 1633
rect 3385 367 3391 1633
rect 3345 355 3391 367
rect 3803 1633 3849 1645
rect 3803 367 3809 1633
rect 3843 367 3849 1633
rect 3803 355 3849 367
rect 4261 1633 4307 1645
rect 4261 367 4267 1633
rect 4301 367 4307 1633
rect 4261 355 4307 367
rect 4719 1633 4765 1645
rect 4719 367 4725 1633
rect 4759 367 4765 1633
rect 4719 355 4765 367
rect 5177 1633 5223 1645
rect 5177 367 5183 1633
rect 5217 367 5223 1633
rect 5177 355 5223 367
rect 5635 1633 5681 1645
rect 5635 367 5641 1633
rect 5675 367 5681 1633
rect 5635 355 5681 367
rect 6093 1633 6139 1645
rect 6093 367 6099 1633
rect 6133 367 6139 1633
rect 6093 355 6139 367
rect 6551 1633 6597 1645
rect 6551 367 6557 1633
rect 6591 367 6597 1633
rect 6551 355 6597 367
rect 7009 1633 7055 1645
rect 7009 367 7015 1633
rect 7049 367 7055 1633
rect 7009 355 7055 367
rect 7467 1633 7513 1645
rect 7467 367 7473 1633
rect 7507 367 7513 1633
rect 7467 355 7513 367
rect 7925 1633 7971 1645
rect 7925 367 7931 1633
rect 7965 367 7971 1633
rect 7925 355 7971 367
rect 8383 1633 8429 1645
rect 8383 367 8389 1633
rect 8423 367 8429 1633
rect 8383 355 8429 367
rect 8841 1633 8887 1645
rect 8841 367 8847 1633
rect 8881 367 8887 1633
rect 8841 355 8887 367
rect 9299 1633 9345 1645
rect 9299 367 9305 1633
rect 9339 367 9345 1633
rect 9299 355 9345 367
rect 9757 1633 9803 1645
rect 9757 367 9763 1633
rect 9797 367 9803 1633
rect 9757 355 9803 367
rect 10215 1633 10261 1645
rect 10215 367 10221 1633
rect 10255 367 10261 1633
rect 10215 355 10261 367
rect 10673 1633 10719 1645
rect 10673 367 10679 1633
rect 10713 367 10719 1633
rect 10673 355 10719 367
rect 11131 1633 11177 1645
rect 11131 367 11137 1633
rect 11171 367 11177 1633
rect 11131 355 11177 367
rect 11589 1633 11635 1645
rect 11589 367 11595 1633
rect 11629 367 11635 1633
rect 11589 355 11635 367
rect 12047 1633 12093 1645
rect 12047 367 12053 1633
rect 12087 367 12093 1633
rect 12047 355 12093 367
rect 12505 1633 12551 1645
rect 12505 367 12511 1633
rect 12545 367 12551 1633
rect 12505 355 12551 367
rect 12963 1633 13009 1645
rect 12963 367 12969 1633
rect 13003 367 13009 1633
rect 12963 355 13009 367
rect 13421 1633 13467 1645
rect 13421 367 13427 1633
rect 13461 367 13467 1633
rect 13421 355 13467 367
rect 13879 1633 13925 1645
rect 13879 367 13885 1633
rect 13919 367 13925 1633
rect 13879 355 13925 367
rect 14337 1633 14383 1645
rect 14337 367 14343 1633
rect 14377 367 14383 1633
rect 14337 355 14383 367
rect 14795 1633 14841 1645
rect 14795 367 14801 1633
rect 14835 367 14841 1633
rect 14795 355 14841 367
rect 15253 1633 15299 1645
rect 15253 367 15259 1633
rect 15293 367 15299 1633
rect 15253 355 15299 367
rect 15711 1633 15757 1645
rect 15711 367 15717 1633
rect 15751 367 15757 1633
rect 15711 355 15757 367
rect 16169 1633 16215 1645
rect 16169 367 16175 1633
rect 16209 367 16215 1633
rect 16169 355 16215 367
rect 16627 1633 16673 1645
rect 16627 367 16633 1633
rect 16667 367 16673 1633
rect 16627 355 16673 367
rect 17085 1633 17131 1645
rect 17085 367 17091 1633
rect 17125 367 17131 1633
rect 17085 355 17131 367
rect 17543 1633 17589 1645
rect 17543 367 17549 1633
rect 17583 367 17589 1633
rect 17543 355 17589 367
rect 18001 1633 18047 1645
rect 18001 367 18007 1633
rect 18041 367 18047 1633
rect 18001 355 18047 367
rect 18459 1633 18505 1645
rect 18459 367 18465 1633
rect 18499 367 18505 1633
rect 18459 355 18505 367
rect 18917 1633 18963 1645
rect 18917 367 18923 1633
rect 18957 367 18963 1633
rect 18917 355 18963 367
rect 19375 1633 19421 1645
rect 19375 367 19381 1633
rect 19415 367 19421 1633
rect 19375 355 19421 367
rect 19833 1633 19879 1645
rect 19833 367 19839 1633
rect 19873 367 19879 1633
rect 19833 355 19879 367
rect 20291 1633 20337 1645
rect 20291 367 20297 1633
rect 20331 367 20337 1633
rect 20291 355 20337 367
rect 20749 1633 20795 1645
rect 20749 367 20755 1633
rect 20789 367 20795 1633
rect 20749 355 20795 367
rect 21207 1633 21253 1645
rect 21207 367 21213 1633
rect 21247 367 21253 1633
rect 21207 355 21253 367
rect 21665 1633 21711 1645
rect 21665 367 21671 1633
rect 21705 367 21711 1633
rect 21665 355 21711 367
rect 22123 1633 22169 1645
rect 22123 367 22129 1633
rect 22163 367 22169 1633
rect 22123 355 22169 367
rect 22581 1633 22627 1645
rect 22581 367 22587 1633
rect 22621 367 22627 1633
rect 22581 355 22627 367
rect 23039 1633 23085 1645
rect 23039 367 23045 1633
rect 23079 367 23085 1633
rect 23039 355 23085 367
rect 23497 1633 23543 1645
rect 23497 367 23503 1633
rect 23537 367 23543 1633
rect 23497 355 23543 367
rect 23955 1633 24001 1645
rect 23955 367 23961 1633
rect 23995 367 24001 1633
rect 23955 355 24001 367
rect 24413 1633 24459 1645
rect 24413 367 24419 1633
rect 24453 367 24459 1633
rect 24413 355 24459 367
rect 24871 1633 24917 1645
rect 24871 367 24877 1633
rect 24911 367 24917 1633
rect 24871 355 24917 367
rect 25329 1633 25375 1645
rect 25329 367 25335 1633
rect 25369 367 25375 1633
rect 25329 355 25375 367
rect 25787 1633 25833 1645
rect 25787 367 25793 1633
rect 25827 367 25833 1633
rect 25787 355 25833 367
rect 26245 1633 26291 1645
rect 26245 367 26251 1633
rect 26285 367 26291 1633
rect 26245 355 26291 367
rect 26703 1633 26749 1645
rect 26703 367 26709 1633
rect 26743 367 26749 1633
rect 26703 355 26749 367
rect 27161 1633 27207 1645
rect 27161 367 27167 1633
rect 27201 367 27207 1633
rect 27161 355 27207 367
rect 27619 1633 27665 1645
rect 27619 367 27625 1633
rect 27659 367 27665 1633
rect 27619 355 27665 367
rect 0 30 27706 60
rect 0 -30 268 30
rect 328 -30 668 30
rect 728 -30 1068 30
rect 1128 -30 1468 30
rect 1528 -30 1868 30
rect 1928 -30 2268 30
rect 2328 -30 2668 30
rect 2728 -30 3068 30
rect 3128 -30 3468 30
rect 3528 -30 3868 30
rect 3928 -30 4268 30
rect 4328 -30 4668 30
rect 4728 -30 5068 30
rect 5128 -30 5468 30
rect 5528 -30 5868 30
rect 5928 -30 6268 30
rect 6328 -30 6668 30
rect 6728 -30 7068 30
rect 7128 -30 7468 30
rect 7528 -30 7868 30
rect 7928 -30 8268 30
rect 8328 -30 8668 30
rect 8728 -30 9068 30
rect 9128 -30 9468 30
rect 9528 -30 9868 30
rect 9928 -30 10268 30
rect 10328 -30 10668 30
rect 10728 -30 11068 30
rect 11128 -30 11468 30
rect 11528 -30 11868 30
rect 11928 -30 12268 30
rect 12328 -30 12668 30
rect 12728 -30 13068 30
rect 13128 -30 13468 30
rect 13528 -30 13868 30
rect 13928 -30 14268 30
rect 14328 -30 14668 30
rect 14728 -30 15068 30
rect 15128 -30 15468 30
rect 15528 -30 15868 30
rect 15928 -30 16268 30
rect 16328 -30 16668 30
rect 16728 -30 17068 30
rect 17128 -30 17468 30
rect 17528 -30 17868 30
rect 17928 -30 18268 30
rect 18328 -30 18668 30
rect 18728 -30 19068 30
rect 19128 -30 19468 30
rect 19528 -30 19868 30
rect 19928 -30 20268 30
rect 20328 -30 20668 30
rect 20728 -30 21068 30
rect 21128 -30 21468 30
rect 21528 -30 21868 30
rect 21928 -30 22268 30
rect 22328 -30 22668 30
rect 22728 -30 23068 30
rect 23128 -30 23468 30
rect 23528 -30 23868 30
rect 23928 -30 24268 30
rect 24328 -30 24668 30
rect 24728 -30 25068 30
rect 25128 -30 25468 30
rect 25528 -30 25868 30
rect 25928 -30 26268 30
rect 26328 -30 26668 30
rect 26728 -30 27068 30
rect 27128 -30 27468 30
rect 27528 -30 27706 30
rect 0 -60 27706 -30
<< labels >>
flabel nwell 0 1850 60 1910 1 FreeSans 800 0 0 0 VPWR
port 4 n power bidirectional
flabel metal1 0 -30 158 30 1 FreeSans 800 0 0 0 VGND
port 5 n ground bidirectional
flabel locali 27646 1730 27706 1790 1 FreeSans 800 0 0 0 SOURCE
port 2 n signal bidirectional
flabel locali 27646 210 27706 270 1 FreeSans 800 0 0 0 DRAIN
port 3 n signal bidirectional
flabel locali 27646 104 27706 164 1 FreeSans 800 0 0 0 GATE
port 1 n signal bidirectional
<< properties >>
string FIXED_BBOX 0 0 27707 1880
string LEFclass CORE
string LEFsite unitasc
<< end >>
