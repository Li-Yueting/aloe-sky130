magic
tech sky130A
magscale 1 2
timestamp 1654939146
<< pwell >>
rect -356 -970 258 526
<< nmoslvt >>
rect -200 -500 200 500
<< ndiff >>
rect -258 488 -200 500
rect -258 -488 -246 488
rect -212 -488 -200 488
rect -258 -500 -200 -488
rect 200 488 258 500
rect 200 -488 212 488
rect 246 -488 258 488
rect 200 -500 258 -488
<< ndiffc >>
rect -246 -488 -212 488
rect 212 -488 246 488
<< psubdiff >>
rect -318 -840 -278 -800
rect -318 -920 -278 -880
<< psubdiffcont >>
rect -318 -880 -278 -840
<< poly >>
rect -200 500 200 526
rect -200 -526 200 -500
rect -138 -716 -18 -526
rect -178 -736 258 -716
rect -178 -796 -88 -736
rect -28 -796 258 -736
rect -178 -816 258 -796
<< polycont >>
rect -88 -796 -28 -736
<< locali >>
rect -356 850 -88 910
rect -28 850 258 910
rect -258 690 258 750
rect 211 504 245 690
rect -246 488 -212 504
rect -247 -488 -246 -446
rect 211 488 246 504
rect 211 486 212 488
rect -247 -504 -212 -488
rect 212 -504 246 -488
rect -247 -570 -213 -504
rect -258 -630 258 -570
rect -328 -840 -268 -760
rect -178 -796 -88 -736
rect -28 -796 258 -736
rect -328 -880 -318 -840
rect -278 -880 -268 -840
rect -328 -970 -268 -880
rect -356 -1030 -88 -970
rect -28 -1030 258 -970
<< viali >>
rect -88 850 -28 910
rect -246 -488 -212 488
rect 212 -488 246 488
rect -88 -1030 -28 -970
<< metal1 >>
rect -356 910 258 940
rect -356 850 -88 910
rect -28 850 258 910
rect -356 820 258 850
rect -252 488 -206 500
rect -252 -488 -246 488
rect -212 -488 -206 488
rect -252 -500 -206 -488
rect 206 488 252 500
rect 206 -488 212 488
rect 246 -488 252 488
rect 206 -500 252 -488
rect -356 -970 258 -940
rect -356 -1030 -88 -970
rect -28 -1030 258 -970
rect -356 -1060 258 -1030
<< labels >>
flabel metal1 -258 850 -198 910 1 FreeSans 800 0 0 0 VPWR
flabel metal1 -258 -1030 -198 -970 1 FreeSans 800 0 0 0 VGND
flabel locali 198 690 258 750 1 FreeSans 800 0 0 0 SOURCE
flabel locali 198 -630 258 -570 1 FreeSans 800 0 0 0 DRAIN
flabel locali 198 -796 258 -736 1 FreeSans 800 0 0 0 GATE
<< end >>
