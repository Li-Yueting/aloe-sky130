* NGSPICE file created from analog_mux_ready.ext - technology: sky130A

.subckt analog_mux_ready out en31_b in_31 en30_b in_30 en29_b in_29 en28_b in_28 en27_b
+ in_27 en26_b in_26 en25_b in_25 en24_b in_24 en23_b in_23 en22_b in_22 en21_b in_21
+ en20_b in_20 en19_b in_19 en18_b in_18 en17_b in_17 en16_b in_16 en15_b in_15 en14_b
+ in_14 en13_b in_13 en12_b in_12 en11_b in_11 en10_b in_10 en9_b in_9 en8_b in_8
+ en7_b in_7 en6_b in_6 en5_b in_5 en4_b in_4 en3_b in_3 en2_b in_2 en1_b in_1 en0_b
+ in_0 en_b en VPWR VGND
X0 a_301_6438# en27_b a_2454_6442# VPWR sky130_fd_pr__pfet_01v8 ad=4.8824e+12p pd=3.71e+07u as=4.8824e+12p ps=3.71e+07u w=1.36e+06u l=150000u
X1 a_301_18021# en18_b a_2454_18025# VPWR sky130_fd_pr__pfet_01v8 ad=4.8824e+12p pd=3.71e+07u as=4.8824e+12p ps=3.71e+07u w=1.36e+06u l=150000u
X2 a_301_1290# en31_b a_2454_1294# VPWR sky130_fd_pr__pfet_01v8 ad=4.8824e+12p pd=3.71e+07u as=4.8824e+12p ps=3.71e+07u w=1.36e+06u l=150000u
X3 out a_2450_12789# a_2454_12877# VGND sky130_fd_pr__nfet_01v8 ad=3.22816e+13p pd=3.2384e+08u as=2.0118e+12p ps=2.02e+07u w=520000u l=150000u
X4 a_301_5151# en_b in_28 VPWR sky130_fd_pr__pfet_01v8 ad=4.8824e+12p pd=3.71e+07u as=2.244e+12p ps=1.69e+07u w=1.36e+06u l=150000u
X5 a_2454_11590# a_2450_11502# out VGND sky130_fd_pr__nfet_01v8 ad=2.0118e+12p pd=2.02e+07u as=0p ps=0u w=520000u l=150000u
X6 VGND en14_b a_2450_23085# VGND sky130_fd_pr__nfet_01v8 ad=1.0048e+13p pd=1.088e+08u as=1.69e+11p ps=1.82e+06u w=650000u l=150000u
X7 a_2454_5155# a_2450_5067# a_301_5151# VGND sky130_fd_pr__nfet_01v8 ad=2.0118e+12p pd=2.02e+07u as=1.8668e+12p ps=1.862e+07u w=520000u l=150000u
X8 a_301_16734# a_2450_16650# a_2454_16738# VGND sky130_fd_pr__nfet_01v8 ad=1.8668e+12p pd=1.862e+07u as=2.0118e+12p ps=2.02e+07u w=520000u l=150000u
X9 out a_2450_10215# a_2454_10303# VGND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.0118e+12p ps=2.02e+07u w=520000u l=150000u
X10 a_301_24456# a_2450_24372# a_2454_24460# VGND sky130_fd_pr__nfet_01v8 ad=1.8668e+12p pd=1.862e+07u as=2.0118e+12p ps=2.02e+07u w=520000u l=150000u
X11 out a_2450_33381# a_2454_33469# VGND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.0118e+12p ps=2.02e+07u w=520000u l=150000u
X12 a_2454_18025# a_2450_17937# out VGND sky130_fd_pr__nfet_01v8 ad=2.0118e+12p pd=2.02e+07u as=0p ps=0u w=520000u l=150000u
X13 a_2454_15451# en20_b out VPWR sky130_fd_pr__pfet_01v8 ad=4.8824e+12p pd=3.71e+07u as=8.44288e+13p ps=6.464e+08u w=1.36e+06u l=150000u
X14 out a_2450_28233# a_2454_28321# VGND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.0118e+12p ps=2.02e+07u w=520000u l=150000u
X15 out a_2450_41103# a_2454_41191# VGND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.0118e+12p ps=2.02e+07u w=520000u l=150000u
X16 in_27 en a_301_6438# VGND sky130_fd_pr__nfet_01v8 ad=8.58e+11p pd=8.5e+06u as=1.8668e+12p ps=1.862e+07u w=520000u l=150000u
X17 a_2454_19312# a_2450_19224# out VGND sky130_fd_pr__nfet_01v8 ad=2.0118e+12p pd=2.02e+07u as=0p ps=0u w=520000u l=150000u
X18 a_2454_32182# a_2450_32094# out VGND sky130_fd_pr__nfet_01v8 ad=2.0118e+12p pd=2.02e+07u as=0p ps=0u w=520000u l=150000u
X19 in_14 en a_301_23169# VGND sky130_fd_pr__nfet_01v8 ad=8.58e+11p pd=8.5e+06u as=1.8668e+12p ps=1.862e+07u w=520000u l=150000u
X20 a_301_33465# en in_6 VGND sky130_fd_pr__nfet_01v8 ad=1.8668e+12p pd=1.862e+07u as=8.58e+11p ps=8.5e+06u w=520000u l=150000u
X21 in_18 en a_301_18021# VGND sky130_fd_pr__nfet_01v8 ad=8.58e+11p pd=8.5e+06u as=1.8668e+12p ps=1.862e+07u w=520000u l=150000u
X22 a_301_18021# en18_b a_2454_18025# VPWR sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.36e+06u l=150000u
X23 a_2454_7729# en26_b a_301_7725# VPWR sky130_fd_pr__pfet_01v8 ad=4.8824e+12p pd=3.71e+07u as=4.8824e+12p ps=3.71e+07u w=1.36e+06u l=150000u
X24 a_301_9012# en_b in_25 VPWR sky130_fd_pr__pfet_01v8 ad=4.8824e+12p pd=3.71e+07u as=2.244e+12p ps=1.69e+07u w=1.36e+06u l=150000u
X25 out en11_b a_2454_27034# VPWR sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=4.8824e+12p ps=3.71e+07u w=1.36e+06u l=150000u
X26 a_2454_37330# en3_b out VPWR sky130_fd_pr__pfet_01v8 ad=4.8824e+12p pd=3.71e+07u as=0p ps=0u w=1.36e+06u l=150000u
X27 in_10 en_b a_301_28317# VPWR sky130_fd_pr__pfet_01v8 ad=2.244e+12p pd=1.69e+07u as=4.8824e+12p ps=3.71e+07u w=1.36e+06u l=150000u
X28 in_0 en_b a_301_41187# VPWR sky130_fd_pr__pfet_01v8 ad=2.244e+12p pd=1.69e+07u as=4.8824e+12p ps=3.71e+07u w=1.36e+06u l=150000u
X29 in_25 en a_301_9012# VGND sky130_fd_pr__nfet_01v8 ad=8.58e+11p pd=8.5e+06u as=1.8668e+12p ps=1.862e+07u w=520000u l=150000u
X30 a_301_10299# en in_24 VGND sky130_fd_pr__nfet_01v8 ad=1.8668e+12p pd=1.862e+07u as=8.58e+11p ps=8.5e+06u w=520000u l=150000u
X31 in_4 en_b a_301_36039# VPWR sky130_fd_pr__pfet_01v8 ad=2.244e+12p pd=1.69e+07u as=4.8824e+12p ps=3.71e+07u w=1.36e+06u l=150000u
X32 in_19 en_b a_301_16734# VPWR sky130_fd_pr__pfet_01v8 ad=2.244e+12p pd=1.69e+07u as=4.8824e+12p ps=3.71e+07u w=1.36e+06u l=150000u
X33 a_301_10299# en_b in_24 VPWR sky130_fd_pr__pfet_01v8 ad=4.8824e+12p pd=3.71e+07u as=2.244e+12p ps=1.69e+07u w=1.36e+06u l=150000u
X34 a_301_38613# en2_b a_2454_38617# VPWR sky130_fd_pr__pfet_01v8 ad=4.8824e+12p pd=3.71e+07u as=4.8824e+12p ps=3.71e+07u w=1.36e+06u l=150000u
X35 out a_2450_6354# a_2454_6442# VGND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.0118e+12p ps=2.02e+07u w=520000u l=150000u
X36 a_2454_5155# en28_b out VPWR sky130_fd_pr__pfet_01v8 ad=4.8824e+12p pd=3.71e+07u as=0p ps=0u w=1.36e+06u l=150000u
X37 a_301_15447# en_b in_20 VPWR sky130_fd_pr__pfet_01v8 ad=4.8824e+12p pd=3.71e+07u as=2.244e+12p ps=1.69e+07u w=1.36e+06u l=150000u
X38 in_10 en a_301_28317# VGND sky130_fd_pr__nfet_01v8 ad=8.58e+11p pd=8.5e+06u as=1.8668e+12p ps=1.862e+07u w=520000u l=150000u
X39 a_2454_15451# a_2450_15363# a_301_15447# VGND sky130_fd_pr__nfet_01v8 ad=2.0118e+12p pd=2.02e+07u as=1.8668e+12p ps=1.862e+07u w=520000u l=150000u
X40 a_2454_18025# en18_b a_301_18021# VPWR sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.36e+06u l=150000u
X41 in_19 en a_301_16734# VGND sky130_fd_pr__nfet_01v8 ad=8.58e+11p pd=8.5e+06u as=0p ps=0u w=520000u l=150000u
X42 a_301_38613# a_2450_38529# a_2454_38617# VGND sky130_fd_pr__nfet_01v8 ad=1.8668e+12p pd=1.862e+07u as=2.0118e+12p ps=2.02e+07u w=520000u l=150000u
X43 a_301_2577# en30_b a_2454_2581# VPWR sky130_fd_pr__pfet_01v8 ad=4.8824e+12p pd=3.71e+07u as=4.8824e+12p ps=3.71e+07u w=1.36e+06u l=150000u
X44 a_2454_30895# en8_b VGND VGND sky130_fd_pr__nfet_01v8 ad=2.0118e+12p pd=2.02e+07u as=0p ps=0u w=500000u l=150000u
X45 a_2454_7729# en26_b out VPWR sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.36e+06u l=150000u
X46 out a_2450_8928# a_2454_9016# VGND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.0118e+12p ps=2.02e+07u w=520000u l=150000u
X47 a_2454_15451# en20_b a_301_15447# VPWR sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.36e+06u l=150000u
X48 a_301_41187# a_2450_41103# a_2454_41191# VGND sky130_fd_pr__nfet_01v8 ad=1.8668e+12p pd=1.862e+07u as=0p ps=0u w=520000u l=150000u
X49 a_301_1290# en in_31 VGND sky130_fd_pr__nfet_01v8 ad=1.8668e+12p pd=1.862e+07u as=8.58e+11p ps=8.5e+06u w=520000u l=150000u
X50 a_301_20595# en16_b a_2454_20599# VPWR sky130_fd_pr__pfet_01v8 ad=4.8824e+12p pd=3.71e+07u as=4.8824e+12p ps=3.71e+07u w=1.36e+06u l=150000u
X51 out en15_b a_2454_21886# VPWR sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=4.8824e+12p ps=3.71e+07u w=1.36e+06u l=150000u
X52 a_2454_32182# en7_b out VPWR sky130_fd_pr__pfet_01v8 ad=4.8824e+12p pd=3.71e+07u as=0p ps=0u w=1.36e+06u l=150000u
X53 in_26 en_b a_301_7725# VPWR sky130_fd_pr__pfet_01v8 ad=2.244e+12p pd=1.69e+07u as=0p ps=0u w=1.36e+06u l=150000u
X54 out en19_b a_2454_16738# VPWR sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=4.8824e+12p ps=3.71e+07u w=1.36e+06u l=150000u
X55 a_2454_39904# en1_b out VPWR sky130_fd_pr__pfet_01v8 ad=4.8824e+12p pd=3.71e+07u as=0p ps=0u w=1.36e+06u l=150000u
X56 a_2454_12877# en22_b out VPWR sky130_fd_pr__pfet_01v8 ad=4.8824e+12p pd=3.71e+07u as=0p ps=0u w=1.36e+06u l=150000u
X57 a_301_21882# en_b in_15 VPWR sky130_fd_pr__pfet_01v8 ad=4.8824e+12p pd=3.71e+07u as=2.244e+12p ps=1.69e+07u w=1.36e+06u l=150000u
X58 a_301_25743# en12_b a_2454_25747# VPWR sky130_fd_pr__pfet_01v8 ad=4.8824e+12p pd=3.71e+07u as=4.8824e+12p ps=3.71e+07u w=1.36e+06u l=150000u
X59 a_2454_36043# en4_b a_301_36039# VPWR sky130_fd_pr__pfet_01v8 ad=4.8824e+12p pd=3.71e+07u as=0p ps=0u w=1.36e+06u l=150000u
X60 a_301_29604# en_b in_9 VPWR sky130_fd_pr__pfet_01v8 ad=4.8824e+12p pd=3.71e+07u as=2.244e+12p ps=1.69e+07u w=1.36e+06u l=150000u
X61 a_301_6438# en_b in_27 VPWR sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.244e+12p ps=1.69e+07u w=1.36e+06u l=150000u
X62 a_301_5151# a_2450_5067# a_2454_5155# VGND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X63 a_301_1290# en_b in_31 VPWR sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.244e+12p ps=1.69e+07u w=1.36e+06u l=150000u
X64 a_2454_30895# a_2450_30807# out VGND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X65 out a_2450_21798# a_2454_21886# VGND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.0118e+12p ps=2.02e+07u w=520000u l=150000u
X66 in_26 en a_301_7725# VGND sky130_fd_pr__nfet_01v8 ad=8.58e+11p pd=8.5e+06u as=1.8668e+12p ps=1.862e+07u w=520000u l=150000u
X67 a_2454_12877# a_2450_12789# out VGND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X68 in_8 en a_301_30891# VGND sky130_fd_pr__nfet_01v8 ad=8.58e+11p pd=8.5e+06u as=1.8668e+12p ps=1.862e+07u w=520000u l=150000u
X69 in_23 en a_301_11586# VGND sky130_fd_pr__nfet_01v8 ad=8.58e+11p pd=8.5e+06u as=1.8668e+12p ps=1.862e+07u w=520000u l=150000u
X70 a_301_25743# a_2450_25659# a_2454_25747# VGND sky130_fd_pr__nfet_01v8 ad=1.8668e+12p pd=1.862e+07u as=2.0118e+12p ps=2.02e+07u w=520000u l=150000u
X71 a_301_21882# en in_15 VGND sky130_fd_pr__nfet_01v8 ad=1.8668e+12p pd=1.862e+07u as=8.58e+11p ps=8.5e+06u w=520000u l=150000u
X72 in_0 en_b a_301_41187# VPWR sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.36e+06u l=150000u
X73 out a_2450_29520# a_2454_29608# VGND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.0118e+12p ps=2.02e+07u w=520000u l=150000u
X74 a_301_41187# a_2450_41103# a_2454_41191# VGND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X75 in_19 en_b a_301_16734# VPWR sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.36e+06u l=150000u
X76 a_2454_27034# a_2450_26946# out VGND sky130_fd_pr__nfet_01v8 ad=2.0118e+12p pd=2.02e+07u as=0p ps=0u w=520000u l=150000u
X77 out a_2450_37242# a_2454_37330# VGND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.0118e+12p ps=2.02e+07u w=520000u l=150000u
X78 a_2454_33469# a_2450_33381# out VGND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X79 a_2454_1294# a_2450_1206# out VGND sky130_fd_pr__nfet_01v8 ad=2.0118e+12p pd=2.02e+07u as=0p ps=0u w=520000u l=150000u
X80 a_2454_32182# a_2450_32094# a_301_32178# VGND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.8668e+12p ps=1.862e+07u w=520000u l=150000u
X81 a_301_41187# en in_0 VGND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=8.58e+11p ps=8.5e+06u w=520000u l=150000u
X82 out a_2450_17937# a_2454_18025# VGND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X83 a_2454_28321# a_2450_28233# out VGND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X84 a_2454_11590# en23_b a_301_11586# VPWR sky130_fd_pr__pfet_01v8 ad=4.8824e+12p pd=3.71e+07u as=4.8824e+12p ps=3.71e+07u w=1.36e+06u l=150000u
X85 out en20_b a_2454_15451# VPWR sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.36e+06u l=150000u
X86 in_17 en a_301_19308# VGND sky130_fd_pr__nfet_01v8 ad=8.58e+11p pd=8.5e+06u as=1.8668e+12p ps=1.862e+07u w=520000u l=150000u
X87 in_7 en a_301_32178# VGND sky130_fd_pr__nfet_01v8 ad=8.58e+11p pd=8.5e+06u as=0p ps=0u w=520000u l=150000u
X88 out a_2450_19224# a_2454_19312# VGND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X89 in_11 en a_301_27030# VGND sky130_fd_pr__nfet_01v8 ad=8.58e+11p pd=8.5e+06u as=1.8668e+12p ps=1.862e+07u w=520000u l=150000u
X90 a_301_18021# en in_18 VGND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X91 a_2454_9016# en25_b a_301_9012# VPWR sky130_fd_pr__pfet_01v8 ad=4.8824e+12p pd=3.71e+07u as=0p ps=0u w=1.36e+06u l=150000u
X92 a_301_27030# en11_b a_2454_27034# VPWR sky130_fd_pr__pfet_01v8 ad=4.8824e+12p pd=3.71e+07u as=0p ps=0u w=1.36e+06u l=150000u
X93 a_2454_37330# en3_b a_301_37326# VPWR sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=4.8824e+12p ps=3.71e+07u w=1.36e+06u l=150000u
X94 VPWR en7_b a_2450_32094# VPWR sky130_fd_pr__pfet_01v8_hvt ad=8.32e+12p pd=8.064e+07u as=2.6e+11p ps=2.52e+06u w=1e+06u l=150000u
X95 a_2454_6442# en27_b out VPWR sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.36e+06u l=150000u
X96 in_3 en_b a_301_37326# VPWR sky130_fd_pr__pfet_01v8 ad=2.244e+12p pd=1.69e+07u as=0p ps=0u w=1.36e+06u l=150000u
X97 a_2454_1294# en31_b out VPWR sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.36e+06u l=150000u
X98 in_19 en a_301_16734# VGND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X99 a_2454_41191# a_2450_41103# a_301_41187# VGND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X100 a_301_14160# en in_21 VGND sky130_fd_pr__nfet_01v8 ad=1.8668e+12p pd=1.862e+07u as=8.58e+11p ps=8.5e+06u w=520000u l=150000u
X101 out a_2450_7641# a_2454_7729# VGND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.0118e+12p ps=2.02e+07u w=520000u l=150000u
X102 a_2454_16738# a_2450_16650# a_301_16734# VGND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X103 a_2454_2581# en30_b a_301_2577# VPWR sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.36e+06u l=150000u
X104 a_301_19308# en_b in_17 VPWR sky130_fd_pr__pfet_01v8 ad=4.8824e+12p pd=3.71e+07u as=2.244e+12p ps=1.69e+07u w=1.36e+06u l=150000u
X105 a_2454_9016# en25_b out VPWR sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.36e+06u l=150000u
X106 a_301_1290# a_2450_1206# a_2454_1294# VGND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X107 a_2454_39904# en1_b VGND VGND sky130_fd_pr__nfet_01v8 ad=2.0118e+12p pd=2.02e+07u as=0p ps=0u w=500000u l=150000u
X108 a_301_33465# en6_b a_2454_33469# VPWR sky130_fd_pr__pfet_01v8 ad=4.8824e+12p pd=3.71e+07u as=4.8824e+12p ps=3.71e+07u w=1.36e+06u l=150000u
X109 a_301_2577# en in_30 VGND sky130_fd_pr__nfet_01v8 ad=1.8668e+12p pd=1.862e+07u as=8.58e+11p ps=8.5e+06u w=520000u l=150000u
X110 a_2454_27034# a_2450_26946# a_301_27030# VGND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X111 a_301_41187# en0_b a_2454_41191# VPWR sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=4.8824e+12p ps=3.71e+07u w=1.36e+06u l=150000u
X112 a_301_14160# en21_b a_2454_14164# VPWR sky130_fd_pr__pfet_01v8 ad=4.8824e+12p pd=3.71e+07u as=4.8824e+12p ps=3.71e+07u w=1.36e+06u l=150000u
X113 a_2454_24460# en13_b a_301_24456# VPWR sky130_fd_pr__pfet_01v8 ad=4.8824e+12p pd=3.71e+07u as=4.8824e+12p ps=3.71e+07u w=1.36e+06u l=150000u
X114 a_301_6438# en27_b a_2454_6442# VPWR sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.36e+06u l=150000u
X115 a_301_18021# a_2450_17937# a_2454_18025# VGND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X116 a_301_6438# a_2450_6354# a_2454_6442# VGND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X117 out en18_b a_2454_18025# VPWR sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.36e+06u l=150000u
X118 VPWR en27_b a_2450_6354# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.6e+11p ps=2.52e+06u w=1e+06u l=150000u
X119 out en7_b a_2454_32182# VPWR sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.36e+06u l=150000u
X120 a_2454_21886# en15_b out VPWR sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.36e+06u l=150000u
X121 out en1_b a_2454_39904# VPWR sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.36e+06u l=150000u
X122 a_2454_16738# en19_b out VPWR sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.36e+06u l=150000u
X123 in_28 en_b a_301_5151# VPWR sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.36e+06u l=150000u
X124 VGND en22_b a_2450_12789# VGND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.69e+11p ps=1.82e+06u w=650000u l=150000u
X125 out en2_b a_2454_38617# VPWR sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.36e+06u l=150000u
X126 a_301_5151# en in_28 VGND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=8.58e+11p ps=8.5e+06u w=520000u l=150000u
X127 a_301_38613# en_b in_2 VPWR sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.244e+12p ps=1.69e+07u w=1.36e+06u l=150000u
X128 out a_2450_30807# a_2454_30895# VGND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X129 a_2454_15451# a_2450_15363# out VGND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X130 a_2454_21886# a_2450_21798# out VGND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X131 VGND en10_b a_2450_28233# VGND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.69e+11p ps=1.82e+06u w=650000u l=150000u
X132 in_16 en a_301_20595# VGND sky130_fd_pr__nfet_01v8 ad=8.58e+11p pd=8.5e+06u as=1.8668e+12p ps=1.862e+07u w=520000u l=150000u
X133 a_301_30891# en in_8 VGND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X134 out a_2450_38529# a_2454_38617# VGND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X135 a_301_34752# en_b in_5 VPWR sky130_fd_pr__pfet_01v8 ad=4.8824e+12p pd=3.71e+07u as=2.244e+12p ps=1.69e+07u w=1.36e+06u l=150000u
X136 a_2454_33469# a_2450_33381# a_301_33465# VGND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X137 a_301_18021# a_2450_17937# a_2454_18025# VGND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X138 a_2454_29608# a_2450_29520# out VGND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X139 a_301_9012# en in_25 VGND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X140 a_301_15447# en20_b a_2454_15451# VPWR sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.36e+06u l=150000u
X141 VPWR en16_b a_2450_20511# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.6e+11p ps=2.52e+06u w=1e+06u l=150000u
X142 a_2454_37330# a_2450_37242# out VGND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X143 out a_2450_26946# a_2454_27034# VGND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X144 out en29_b a_2454_3868# VPWR sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=4.8824e+12p ps=3.71e+07u w=1.36e+06u l=150000u
X145 in_10 en a_301_28317# VGND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X146 in_0 en a_301_41187# VGND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X147 a_301_38613# en in_2 VGND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=8.58e+11p ps=8.5e+06u w=520000u l=150000u
X148 a_301_19308# en in_17 VGND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X149 a_2454_23173# en14_b VGND VGND sky130_fd_pr__nfet_01v8 ad=2.0118e+12p pd=2.02e+07u as=0p ps=0u w=500000u l=150000u
X150 a_2454_5155# a_2450_5067# out VGND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X151 a_301_34752# en in_5 VGND sky130_fd_pr__nfet_01v8 ad=1.8668e+12p pd=1.862e+07u as=8.58e+11p ps=8.5e+06u w=520000u l=150000u
X152 a_301_15447# en in_20 VGND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=8.58e+11p ps=8.5e+06u w=520000u l=150000u
X153 a_2454_18025# a_2450_17937# a_301_18021# VGND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X154 a_301_2577# a_2450_2493# a_2454_2581# VGND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.0118e+12p ps=2.02e+07u w=520000u l=150000u
X155 a_2454_1294# a_2450_1206# a_301_1290# VGND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X156 a_2454_2581# en30_b VGND VGND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X157 a_2454_20599# a_2450_20511# a_301_20595# VGND sky130_fd_pr__nfet_01v8 ad=2.0118e+12p pd=2.02e+07u as=0p ps=0u w=520000u l=150000u
X158 a_2454_15451# a_2450_15363# a_301_15447# VGND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X159 a_301_30891# a_2450_30807# a_2454_30895# VGND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X160 a_301_10299# en24_b a_2454_10303# VPWR sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=4.8824e+12p ps=3.71e+07u w=1.36e+06u l=150000u
X161 out a_2450_41103# a_2454_41191# VGND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X162 a_2454_6442# en27_b a_301_6438# VPWR sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.36e+06u l=150000u
X163 a_2454_32182# a_2450_32094# out VGND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X164 a_2454_11590# en23_b out VPWR sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.36e+06u l=150000u
X165 a_301_11586# en_b in_23 VPWR sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.244e+12p ps=1.69e+07u w=1.36e+06u l=150000u
X166 a_2454_36043# a_2450_35955# a_301_36039# VGND sky130_fd_pr__nfet_01v8 ad=2.0118e+12p pd=2.02e+07u as=1.8668e+12p ps=1.862e+07u w=520000u l=150000u
X167 a_2454_36043# en4_b out VPWR sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.36e+06u l=150000u
X168 a_301_7725# a_2450_7641# a_2454_7729# VGND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X169 in_31 en_b a_301_1290# VPWR sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.36e+06u l=150000u
X170 out en11_b a_2454_27034# VPWR sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.36e+06u l=150000u
X171 a_2454_37330# en3_b out VPWR sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.36e+06u l=150000u
X172 a_2454_21886# en15_b a_301_21882# VPWR sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.36e+06u l=150000u
X173 in_0 en_b a_301_41187# VPWR sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.36e+06u l=150000u
X174 a_2454_18025# en18_b out VPWR sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.36e+06u l=150000u
X175 in_4 en_b a_301_36039# VPWR sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.36e+06u l=150000u
X176 in_19 en_b a_301_16734# VPWR sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.36e+06u l=150000u
X177 a_301_27030# en_b in_11 VPWR sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.244e+12p ps=1.69e+07u w=1.36e+06u l=150000u
X178 a_301_6438# en in_27 VGND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X179 a_2454_38617# en2_b out VPWR sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.36e+06u l=150000u
X180 in_0 en a_301_41187# VGND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X181 a_2454_16738# a_2450_16650# out VGND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X182 a_301_30891# a_2450_30807# a_2454_30895# VGND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X183 a_301_23169# en_b in_14 VPWR sky130_fd_pr__pfet_01v8 ad=4.8824e+12p pd=3.71e+07u as=2.244e+12p ps=1.69e+07u w=1.36e+06u l=150000u
X184 a_2454_21886# a_2450_21798# a_301_21882# VGND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X185 VGND en9_b a_2450_29520# VGND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.69e+11p ps=1.82e+06u w=650000u l=150000u
X186 a_301_30891# en_b in_8 VPWR sky130_fd_pr__pfet_01v8 ad=4.8824e+12p pd=3.71e+07u as=2.244e+12p ps=1.69e+07u w=1.36e+06u l=150000u
X187 out a_2450_15363# a_2454_15451# VGND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X188 in_19 en a_301_16734# VGND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X189 a_2454_33469# en6_b a_301_33465# VPWR sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.36e+06u l=150000u
X190 a_2454_9016# a_2450_8928# a_301_9012# VGND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X191 a_2454_41191# en0_b a_301_41187# VPWR sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.36e+06u l=150000u
X192 a_2454_38617# a_2450_38529# out VGND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X193 a_2454_37330# a_2450_37242# a_301_37326# VGND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.8668e+12p ps=1.862e+07u w=520000u l=150000u
X194 a_2454_6442# a_2450_6354# out VGND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X195 a_301_27030# a_2450_26946# a_2454_27034# VGND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X196 out en28_b a_2454_5155# VPWR sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.36e+06u l=150000u
X197 in_3 en a_301_37326# VGND sky130_fd_pr__nfet_01v8 ad=8.58e+11p pd=8.5e+06u as=0p ps=0u w=520000u l=150000u
X198 a_2454_30895# a_2450_30807# a_301_30891# VGND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X199 a_2454_24460# en13_b VGND VGND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X200 VPWR en3_b a_2450_37242# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.6e+11p ps=2.52e+06u w=1e+06u l=150000u
X201 a_2454_11590# en23_b a_301_11586# VPWR sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.36e+06u l=150000u
X202 a_2454_2581# en30_b a_301_2577# VPWR sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.36e+06u l=150000u
X203 a_2454_2581# a_2450_2493# a_301_2577# VGND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X204 a_301_3864# a_2450_3780# a_2454_3868# VGND sky130_fd_pr__nfet_01v8 ad=1.8668e+12p pd=1.862e+07u as=2.0118e+12p ps=2.02e+07u w=520000u l=150000u
X205 a_2454_9016# a_2450_8928# out VGND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X206 a_301_7725# en_b in_26 VPWR sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.36e+06u l=150000u
X207 a_2454_6442# en27_b VGND VGND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X208 a_2454_16738# a_2450_16650# a_301_16734# VGND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X209 a_301_14160# a_2450_14076# a_2454_14164# VGND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.0118e+12p ps=2.02e+07u w=520000u l=150000u
X210 a_301_6438# a_2450_6354# a_2454_6442# VGND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X211 a_2454_24460# a_2450_24372# a_301_24456# VGND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X212 a_2454_33469# a_2450_33381# out VGND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X213 a_2454_24460# en13_b out VPWR sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.36e+06u l=150000u
X214 out a_2450_17937# a_2454_18025# VGND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X215 a_2454_41191# a_2450_41103# out VGND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X216 out en20_b a_2454_15451# VPWR sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.36e+06u l=150000u
X217 in_7 en a_301_32178# VGND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X218 out a_2450_32094# a_2454_32182# VGND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X219 a_301_23169# en in_14 VGND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X220 a_301_7725# en in_26 VGND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X221 in_28 en a_301_5151# VGND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X222 out en23_b a_2454_11590# VPWR sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.36e+06u l=150000u
X223 a_301_19308# en17_b a_2454_19312# VPWR sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=4.8824e+12p ps=3.71e+07u w=1.36e+06u l=150000u
X224 out en4_b a_2454_36043# VPWR sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.36e+06u l=150000u
X225 in_3 en_b a_301_37326# VPWR sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.36e+06u l=150000u
X226 out en3_b a_2454_37330# VPWR sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.36e+06u l=150000u
X227 a_2454_27034# en11_b out VPWR sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.36e+06u l=150000u
X228 a_301_34752# en_b in_5 VPWR sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.36e+06u l=150000u
X229 a_301_28317# en_b in_10 VPWR sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.36e+06u l=150000u
X230 in_12 en_b a_301_25743# VPWR sky130_fd_pr__pfet_01v8 ad=2.244e+12p pd=1.69e+07u as=0p ps=0u w=1.36e+06u l=150000u
X231 a_301_36039# en_b in_4 VPWR sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.36e+06u l=150000u
X232 a_2454_38617# en2_b a_301_38613# VPWR sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.36e+06u l=150000u
X233 a_301_24456# en_b in_13 VPWR sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.244e+12p ps=1.69e+07u w=1.36e+06u l=150000u
X234 a_301_32178# en_b in_7 VPWR sky130_fd_pr__pfet_01v8 ad=4.8824e+12p pd=3.71e+07u as=2.244e+12p ps=1.69e+07u w=1.36e+06u l=150000u
X235 a_301_39900# en_b in_1 VPWR sky130_fd_pr__pfet_01v8 ad=4.8824e+12p pd=3.71e+07u as=2.244e+12p ps=1.69e+07u w=1.36e+06u l=150000u
X236 a_301_15447# a_2450_15363# a_2454_15451# VGND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X237 out a_2450_16650# a_2454_16738# VGND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X238 a_301_34752# en in_5 VGND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X239 a_2454_3868# en29_b out VPWR sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.36e+06u l=150000u
X240 out en31_b a_2454_1294# VPWR sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.36e+06u l=150000u
X241 in_12 en a_301_25743# VGND sky130_fd_pr__nfet_01v8 ad=8.58e+11p pd=8.5e+06u as=0p ps=0u w=520000u l=150000u
X242 a_2454_12877# en22_b VGND VGND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X243 a_2454_38617# a_2450_38529# a_301_38613# VGND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X244 a_2454_7729# a_2450_7641# out VGND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X245 a_2454_20599# en16_b VGND VGND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X246 a_301_2577# en30_b a_2454_2581# VPWR sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.36e+06u l=150000u
X247 a_301_7725# en26_b a_2454_7729# VPWR sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.36e+06u l=150000u
X248 out en30_b a_2454_2581# VPWR sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.36e+06u l=150000u
X249 a_301_29604# en9_b a_2454_29608# VPWR sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=4.8824e+12p ps=3.71e+07u w=1.36e+06u l=150000u
X250 a_301_39900# en in_1 VGND sky130_fd_pr__nfet_01v8 ad=1.8668e+12p pd=1.862e+07u as=8.58e+11p ps=8.5e+06u w=520000u l=150000u
X251 a_2454_20599# en16_b a_301_20595# VPWR sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.36e+06u l=150000u
X252 a_2454_21886# en15_b out VPWR sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.36e+06u l=150000u
X253 a_2454_3868# a_2450_3780# a_301_3864# VGND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X254 a_301_34752# en5_b a_2454_34756# VPWR sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=4.8824e+12p ps=3.71e+07u w=1.36e+06u l=150000u
X255 a_301_36039# en4_b a_2454_36043# VPWR sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.36e+06u l=150000u
X256 a_2454_25747# en12_b a_301_25743# VPWR sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.36e+06u l=150000u
X257 a_2454_20599# a_2450_20511# out VGND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X258 out a_2450_30807# a_2454_30895# VGND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X259 a_301_10299# a_2450_10215# a_2454_10303# VGND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X260 a_2454_6442# a_2450_6354# a_301_6438# VGND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X261 a_2454_21886# a_2450_21798# out VGND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X262 a_301_34752# a_2450_34668# a_2454_34756# VGND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.0118e+12p ps=2.02e+07u w=520000u l=150000u
X263 a_2454_7729# en26_b VGND VGND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X264 in_16 en a_301_20595# VGND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X265 a_301_7725# a_2450_7641# a_2454_7729# VGND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X266 a_301_11586# en in_23 VGND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X267 a_2454_25747# a_2450_25659# a_301_25743# VGND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X268 a_2454_36043# a_2450_35955# out VGND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X269 a_301_5151# en_b in_28 VPWR sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.36e+06u l=150000u
X270 a_2454_33469# en6_b out VPWR sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.36e+06u l=150000u
X271 a_2454_41191# en0_b out VPWR sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.36e+06u l=150000u
X272 a_2454_37330# a_2450_37242# out VGND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X273 out a_2450_26946# a_2454_27034# VGND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X274 out a_2450_33381# a_2454_33469# VGND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X275 a_2454_18025# a_2450_17937# out VGND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X276 out en13_b a_2454_24460# VPWR sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.36e+06u l=150000u
X277 in_0 en a_301_41187# VGND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X278 a_2454_15451# en20_b out VPWR sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.36e+06u l=150000u
X279 in_27 en a_301_6438# VGND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X280 a_301_11586# en23_b a_2454_11590# VPWR sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.36e+06u l=150000u
X281 a_301_23169# en_b in_14 VPWR sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.36e+06u l=150000u
X282 a_301_32178# en in_7 VGND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X283 a_301_30891# en_b in_8 VPWR sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.36e+06u l=150000u
X284 in_21 en_b a_301_14160# VPWR sky130_fd_pr__pfet_01v8 ad=2.244e+12p pd=1.69e+07u as=0p ps=0u w=1.36e+06u l=150000u
X285 a_301_27030# en in_11 VGND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X286 a_301_36039# en4_b a_2454_36043# VPWR sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.36e+06u l=150000u
X287 VPWR en15_b a_2450_21798# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.6e+11p ps=2.52e+06u w=1e+06u l=150000u
X288 a_2454_27034# en11_b a_301_27030# VPWR sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.36e+06u l=150000u
X289 a_301_37326# en_b in_3 VPWR sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.36e+06u l=150000u
X290 in_5 en_b a_301_34752# VPWR sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.36e+06u l=150000u
X291 a_301_36039# en in_4 VGND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=8.58e+11p ps=8.5e+06u w=520000u l=150000u
X292 a_301_33465# en_b in_6 VPWR sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.244e+12p ps=1.69e+07u w=1.36e+06u l=150000u
X293 a_301_16734# a_2450_16650# a_2454_16738# VGND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X294 a_2454_36043# en4_b a_301_36039# VPWR sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.36e+06u l=150000u
X295 a_2454_5155# en28_b out VPWR sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.36e+06u l=150000u
X296 out a_2450_5067# a_2454_5155# VGND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X297 in_5 en a_301_34752# VGND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X298 a_2454_7729# en26_b a_301_7725# VPWR sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.36e+06u l=150000u
X299 a_2454_2581# a_2450_2493# a_301_2577# VGND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X300 a_2454_29608# en9_b VGND VGND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X301 a_2454_33469# en6_b a_301_33465# VPWR sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.36e+06u l=150000u
X302 a_301_9012# en25_b a_2454_9016# VPWR sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.36e+06u l=150000u
X303 a_301_23169# en14_b a_2454_23173# VPWR sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=4.8824e+12p ps=3.71e+07u w=1.36e+06u l=150000u
X304 a_2454_41191# en0_b a_301_41187# VPWR sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.36e+06u l=150000u
X305 a_2454_14164# en21_b a_301_14160# VPWR sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.36e+06u l=150000u
X306 a_301_30891# en8_b a_2454_30895# VPWR sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=4.8824e+12p ps=3.71e+07u w=1.36e+06u l=150000u
X307 a_301_24456# en13_b a_2454_24460# VPWR sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.36e+06u l=150000u
X308 out en15_b a_2454_21886# VPWR sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.36e+06u l=150000u
X309 a_2454_38617# en2_b out VPWR sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.36e+06u l=150000u
X310 a_2454_7729# a_2450_7641# a_301_7725# VGND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X311 a_2454_24460# a_2450_24372# out VGND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X312 out a_2450_20511# a_2454_20599# VGND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X313 a_301_1290# en_b in_31 VPWR sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.36e+06u l=150000u
X314 out a_2450_15363# a_2454_15451# VGND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X315 a_2454_30895# a_2450_30807# out VGND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X316 VGND en18_b a_2450_17937# VGND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.69e+11p ps=1.82e+06u w=650000u l=150000u
X317 out a_2450_21798# a_2454_21886# VGND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X318 in_24 en a_301_10299# VGND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X319 a_301_19308# a_2450_19224# a_2454_19312# VGND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X320 a_301_20595# en in_16 VGND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X321 a_2454_38617# a_2450_38529# out VGND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X322 in_5 en_b a_301_34752# VPWR sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.36e+06u l=150000u
X323 in_24 en_b a_301_10299# VPWR sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.36e+06u l=150000u
X324 a_301_24456# en13_b a_2454_24460# VPWR sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.36e+06u l=150000u
X325 out a_2450_35955# a_2454_36043# VGND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X326 VPWR en24_b a_2450_10215# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.6e+11p ps=2.52e+06u w=1e+06u l=150000u
X327 a_2454_15451# en20_b a_301_15447# VPWR sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.36e+06u l=150000u
X328 in_3 en a_301_37326# VGND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X329 out en6_b a_2454_33469# VPWR sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.36e+06u l=150000u
X330 a_301_24456# en_b in_13 VPWR sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.36e+06u l=150000u
X331 a_2454_27034# a_2450_26946# out VGND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X332 a_2454_29608# en9_b a_301_29604# VPWR sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.36e+06u l=150000u
X333 out en0_b a_2454_41191# VPWR sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.36e+06u l=150000u
X334 out a_2450_37242# a_2454_37330# VGND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X335 in_20 en_b a_301_15447# VPWR sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.36e+06u l=150000u
X336 a_301_28317# en in_10 VGND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X337 a_2454_1294# a_2450_1206# out VGND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X338 in_14 en_b a_301_23169# VPWR sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.36e+06u l=150000u
X339 a_2454_34756# en5_b a_301_34752# VPWR sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.36e+06u l=150000u
X340 in_8 en_b a_301_30891# VPWR sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.36e+06u l=150000u
X341 a_301_24456# en in_13 VGND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=8.58e+11p ps=8.5e+06u w=520000u l=150000u
X342 in_5 en a_301_34752# VGND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X343 a_2454_6442# en27_b out VPWR sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.36e+06u l=150000u
X344 a_2454_24460# en13_b a_301_24456# VPWR sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.36e+06u l=150000u
X345 a_2454_1294# en31_b out VPWR sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.36e+06u l=150000u
X346 a_2454_34756# a_2450_34668# a_301_34752# VGND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X347 a_301_39900# en in_1 VGND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X348 a_301_2577# a_2450_2493# a_2454_2581# VGND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X349 a_2454_9016# en25_b a_301_9012# VPWR sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.36e+06u l=150000u
X350 a_301_20595# a_2450_20511# a_2454_20599# VGND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X351 out a_2450_2493# a_2454_2581# VGND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X352 a_2454_10303# en24_b a_301_10299# VPWR sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.36e+06u l=150000u
X353 a_2454_3868# a_2450_3780# a_301_3864# VGND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X354 a_2454_20599# en16_b out VPWR sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.36e+06u l=150000u
X355 out en23_b a_2454_11590# VPWR sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.36e+06u l=150000u
X356 a_301_32178# en7_b a_2454_32182# VPWR sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.36e+06u l=150000u
X357 a_301_39900# en1_b a_2454_39904# VPWR sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.36e+06u l=150000u
X358 a_301_36039# a_2450_35955# a_2454_36043# VGND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X359 a_2454_25747# en12_b out VPWR sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.36e+06u l=150000u
X360 out en4_b a_2454_36043# VPWR sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.36e+06u l=150000u
X361 a_2454_27034# en11_b out VPWR sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.36e+06u l=150000u
X362 a_301_41187# en_b in_0 VPWR sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.36e+06u l=150000u
X363 in_12 en_b a_301_25743# VPWR sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.36e+06u l=150000u
X364 a_301_16734# en_b in_19 VPWR sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.36e+06u l=150000u
X365 a_2454_25747# a_2450_25659# out VGND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X366 out en2_b a_2454_38617# VPWR sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.36e+06u l=150000u
X367 a_301_20595# a_2450_20511# a_2454_20599# VGND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X368 a_301_5151# en in_28 VGND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X369 a_301_12873# en_b in_22 VPWR sky130_fd_pr__pfet_01v8 ad=4.8824e+12p pd=3.71e+07u as=2.244e+12p ps=1.69e+07u w=1.36e+06u l=150000u
X370 out a_2450_16650# a_2454_16738# VGND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X371 in_29 en_b a_301_3864# VPWR sky130_fd_pr__pfet_01v8 ad=2.244e+12p pd=1.69e+07u as=4.8824e+12p ps=3.71e+07u w=1.36e+06u l=150000u
X372 a_301_20595# en_b in_16 VPWR sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.244e+12p ps=1.69e+07u w=1.36e+06u l=150000u
X373 in_14 en_b a_301_23169# VPWR sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.36e+06u l=150000u
X374 out a_2450_24372# a_2454_24460# VGND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X375 in_8 en_b a_301_30891# VPWR sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.36e+06u l=150000u
X376 a_301_39900# a_2450_39816# a_2454_39904# VGND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X377 a_2454_15451# a_2450_15363# out VGND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X378 in_12 en a_301_25743# VGND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X379 a_301_16734# en in_19 VGND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X380 in_21 en a_301_14160# VGND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X381 a_301_36039# a_2450_35955# a_2454_36043# VGND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X382 a_2454_23173# en14_b a_301_23169# VPWR sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.36e+06u l=150000u
X383 a_301_33465# en6_b a_2454_33469# VPWR sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.36e+06u l=150000u
X384 a_2454_27034# a_2450_26946# a_301_27030# VGND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X385 a_2454_30895# en8_b a_301_30891# VPWR sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.36e+06u l=150000u
X386 a_301_41187# en0_b a_2454_41191# VPWR sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.36e+06u l=150000u
X387 out a_2450_38529# a_2454_38617# VGND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X388 a_301_36039# en in_4 VGND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X389 a_301_12873# en in_22 VGND sky130_fd_pr__nfet_01v8 ad=1.8668e+12p pd=1.862e+07u as=8.58e+11p ps=8.5e+06u w=520000u l=150000u
X390 a_2454_20599# a_2450_20511# a_301_20595# VGND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X391 a_301_37326# en in_3 VGND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X392 in_29 en a_301_3864# VGND sky130_fd_pr__nfet_01v8 ad=8.58e+11p pd=8.5e+06u as=0p ps=0u w=520000u l=150000u
X393 in_13 en_b a_301_24456# VPWR sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.36e+06u l=150000u
X394 in_17 en_b a_301_19308# VPWR sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.36e+06u l=150000u
X395 out en29_b a_2454_3868# VPWR sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.36e+06u l=150000u
X396 VPWR en17_b a_2450_19224# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.6e+11p ps=2.52e+06u w=1e+06u l=150000u
X397 VPWR en11_b a_2450_26946# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.6e+11p ps=2.52e+06u w=1e+06u l=150000u
X398 a_301_33465# en in_6 VGND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X399 a_2454_36043# a_2450_35955# a_301_36039# VGND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X400 a_2454_5155# a_2450_5067# out VGND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X401 a_2454_7729# en26_b a_301_7725# VPWR sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.36e+06u l=150000u
X402 a_301_3864# a_2450_3780# a_2454_3868# VGND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X403 in_1 en a_301_39900# VGND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X404 a_301_23169# a_2450_23085# a_2454_23173# VGND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X405 out a_2450_3780# a_2454_3868# VGND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X406 a_301_9012# a_2450_8928# a_2454_9016# VGND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X407 a_2454_14164# a_2450_14076# a_301_14160# VGND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X408 a_2454_14164# en21_b out VPWR sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.36e+06u l=150000u
X409 a_301_24456# a_2450_24372# a_2454_24460# VGND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X410 out en13_b a_2454_24460# VPWR sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.36e+06u l=150000u
X411 in_30 en_b a_301_2577# VPWR sky130_fd_pr__pfet_01v8 ad=2.244e+12p pd=1.69e+07u as=0p ps=0u w=1.36e+06u l=150000u
X412 a_2454_15451# en20_b out VPWR sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.36e+06u l=150000u
X413 a_2454_29608# en9_b out VPWR sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.36e+06u l=150000u
X414 in_21 en_b a_301_14160# VPWR sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.36e+06u l=150000u
X415 out en16_b a_2454_20599# VPWR sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.36e+06u l=150000u
X416 a_301_28317# en10_b a_2454_28321# VPWR sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=4.8824e+12p ps=3.71e+07u w=1.36e+06u l=150000u
X417 a_2454_11590# en23_b out VPWR sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.36e+06u l=150000u
X418 a_2454_19312# en17_b a_301_19308# VPWR sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.36e+06u l=150000u
X419 a_2454_34756# en5_b out VPWR sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.36e+06u l=150000u
X420 out en12_b a_2454_25747# VPWR sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.36e+06u l=150000u
X421 a_2454_36043# en4_b out VPWR sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.36e+06u l=150000u
X422 out en11_b a_2454_27034# VPWR sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.36e+06u l=150000u
X423 in_5 en_b a_301_34752# VPWR sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.36e+06u l=150000u
X424 in_28 en_b a_301_5151# VPWR sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.36e+06u l=150000u
X425 a_301_25743# en_b in_12 VPWR sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.36e+06u l=150000u
X426 out en30_b a_2454_2581# VPWR sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.36e+06u l=150000u
X427 a_2454_34756# a_2450_34668# out VGND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X428 a_301_6438# en in_27 VGND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X429 in_13 en_b a_301_24456# VPWR sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.36e+06u l=150000u
X430 a_301_21882# en_b in_15 VPWR sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.36e+06u l=150000u
X431 a_301_24456# a_2450_24372# a_2454_24460# VGND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X432 out a_2450_25659# a_2454_25747# VGND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X433 a_301_29604# en_b in_9 VPWR sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.36e+06u l=150000u
X434 a_2454_15451# a_2450_15363# a_301_15447# VGND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X435 a_2454_16738# a_2450_16650# out VGND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X436 a_301_24456# en in_13 VGND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X437 in_5 en a_301_34752# VGND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X438 in_20 en a_301_15447# VGND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X439 a_301_25743# en in_12 VGND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X440 VPWR en20_b a_2450_15363# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.6e+11p ps=2.52e+06u w=1e+06u l=150000u
X441 a_301_21882# en in_15 VGND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X442 in_4 en a_301_36039# VGND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X443 a_2454_6442# a_2450_6354# out VGND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X444 out en28_b a_2454_5155# VPWR sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.36e+06u l=150000u
X445 a_2454_24460# a_2450_24372# a_301_24456# VGND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X446 a_2454_18025# en18_b VGND VGND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X447 a_2454_29608# en9_b a_301_29604# VPWR sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.36e+06u l=150000u
X448 a_301_29604# en in_9 VGND sky130_fd_pr__nfet_01v8 ad=1.8668e+12p pd=1.862e+07u as=8.58e+11p ps=8.5e+06u w=520000u l=150000u
X449 in_1 en a_301_39900# VGND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X450 a_301_20595# en16_b a_2454_20599# VPWR sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.36e+06u l=150000u
X451 a_301_7725# en26_b a_2454_7729# VPWR sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.36e+06u l=150000u
X452 a_2454_34756# en5_b a_301_34752# VPWR sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.36e+06u l=150000u
X453 a_301_25743# en12_b a_2454_25747# VPWR sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.36e+06u l=150000u
X454 out en26_b a_2454_7729# VPWR sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.36e+06u l=150000u
X455 a_2454_39904# a_2450_39816# a_301_39900# VGND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X456 a_2454_9016# en25_b a_301_9012# VPWR sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.36e+06u l=150000u
X457 a_301_11586# a_2450_11502# a_2454_11590# VGND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X458 a_2454_9016# a_2450_8928# a_301_9012# VGND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X459 out a_2450_20511# a_2454_20599# VGND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X460 a_2454_10303# a_2450_10215# a_301_10299# VGND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X461 a_2454_10303# en24_b out VPWR sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.36e+06u l=150000u
X462 in_31 en a_301_1290# VGND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X463 in_24 en a_301_10299# VGND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X464 a_2454_34756# a_2450_34668# a_301_34752# VGND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X465 a_301_32178# a_2450_32094# a_2454_32182# VGND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X466 in_24 en_b a_301_10299# VPWR sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.36e+06u l=150000u
X467 a_301_25743# a_2450_25659# a_2454_25747# VGND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X468 out a_2450_35955# a_2454_36043# VGND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X469 out en6_b a_2454_33469# VPWR sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.36e+06u l=150000u
X470 a_2454_23173# en14_b out VPWR sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.36e+06u l=150000u
X471 out en0_b a_2454_41191# VPWR sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.36e+06u l=150000u
X472 out en21_b a_2454_14164# VPWR sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.36e+06u l=150000u
X473 a_2454_27034# a_2450_26946# out VGND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X474 a_2454_30895# en8_b out VPWR sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.36e+06u l=150000u
X475 a_2454_24460# en13_b out VPWR sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.36e+06u l=150000u
X476 in_27 en_b a_301_6438# VPWR sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.36e+06u l=150000u
X477 in_20 en_b a_301_15447# VPWR sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.36e+06u l=150000u
X478 a_301_20595# en16_b a_2454_20599# VPWR sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.36e+06u l=150000u
X479 a_301_41187# en in_0 VGND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X480 a_2454_11590# en23_b a_301_11586# VPWR sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.36e+06u l=150000u
X481 a_301_12873# en_b in_22 VPWR sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.36e+06u l=150000u
X482 out en20_b a_2454_15451# VPWR sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.36e+06u l=150000u
X483 a_301_20595# en_b in_16 VPWR sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.36e+06u l=150000u
X484 in_14 en_b a_301_23169# VPWR sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.36e+06u l=150000u
X485 out en9_b a_2454_29608# VPWR sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.36e+06u l=150000u
X486 a_301_37326# en3_b a_2454_37330# VPWR sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.36e+06u l=150000u
X487 in_31 en_b a_301_1290# VPWR sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.36e+06u l=150000u
X488 in_8 en_b a_301_30891# VPWR sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.36e+06u l=150000u
X489 a_301_14160# en_b in_21 VPWR sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.36e+06u l=150000u
X490 a_301_25743# en12_b a_2454_25747# VPWR sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.36e+06u l=150000u
X491 out en5_b a_2454_34756# VPWR sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.36e+06u l=150000u
X492 a_301_3864# en_b in_29 VPWR sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.36e+06u l=150000u
X493 a_301_12873# en in_22 VGND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X494 a_2454_20599# en16_b a_301_20595# VPWR sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.36e+06u l=150000u
X495 in_4 en a_301_36039# VGND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X496 out a_2450_1206# a_2454_1294# VGND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X497 a_301_25743# a_2450_25659# a_2454_25747# VGND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X498 a_301_18021# en_b in_18 VPWR sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.244e+12p ps=1.69e+07u w=1.36e+06u l=150000u
X499 out a_2450_34668# a_2454_34756# VGND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X500 in_25 en_b a_301_9012# VPWR sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.36e+06u l=150000u
X501 a_2454_16738# a_2450_16650# a_301_16734# VGND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X502 a_2454_23173# a_2450_23085# a_301_23169# VGND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X503 a_2454_25747# en12_b a_301_25743# VPWR sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.36e+06u l=150000u
X504 a_301_3864# en in_29 VGND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X505 VGND en28_b a_2450_5067# VGND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.69e+11p ps=1.82e+06u w=650000u l=150000u
X506 out en27_b a_2454_6442# VPWR sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.36e+06u l=150000u
X507 in_13 en a_301_24456# VGND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X508 a_301_38613# en_b in_2 VPWR sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.36e+06u l=150000u
X509 out en31_b a_2454_1294# VPWR sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.36e+06u l=150000u
X510 a_2454_28321# en10_b a_301_28317# VPWR sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.36e+06u l=150000u
X511 a_2454_7729# a_2450_7641# out VGND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X512 a_2454_25747# a_2450_25659# a_301_25743# VGND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X513 a_301_12873# en22_b a_2454_12877# VPWR sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.36e+06u l=150000u
X514 a_2454_23173# en14_b a_301_23169# VPWR sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.36e+06u l=150000u
X515 a_2454_30895# en8_b a_301_30891# VPWR sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.36e+06u l=150000u
X516 a_301_14160# en21_b a_2454_14164# VPWR sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.36e+06u l=150000u
X517 a_301_2577# en30_b a_2454_2581# VPWR sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.36e+06u l=150000u
X518 a_301_38613# en in_2 VGND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X519 a_301_9012# en25_b a_2454_9016# VPWR sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.36e+06u l=150000u
X520 out en25_b a_2454_9016# VPWR sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.36e+06u l=150000u
X521 a_2454_1294# a_2450_1206# a_301_1290# VGND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X522 a_301_12873# a_2450_12789# a_2454_12877# VGND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X523 a_2454_14164# a_2450_14076# out VGND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X524 out a_2450_24372# a_2454_24460# VGND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X525 a_2454_20599# a_2450_20511# out VGND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X526 in_30 en a_301_2577# VGND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X527 a_2454_15451# a_2450_15363# out VGND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X528 a_2454_6442# en27_b a_301_6438# VPWR sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.36e+06u l=150000u
X529 out en24_b a_2454_10303# VPWR sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.36e+06u l=150000u
X530 a_301_33465# a_2450_33381# a_2454_33469# VGND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X531 in_21 en a_301_14160# VGND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X532 a_301_28317# a_2450_28233# a_2454_28321# VGND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X533 a_301_10299# en in_24 VGND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X534 a_2454_19312# a_2450_19224# a_301_19308# VGND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X535 a_301_14160# en21_b a_2454_14164# VPWR sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.36e+06u l=150000u
X536 a_2454_19312# en17_b out VPWR sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.36e+06u l=150000u
X537 a_301_10299# en_b in_24 VPWR sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.36e+06u l=150000u
X538 a_2454_36043# a_2450_35955# out VGND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X539 a_301_5151# en_b in_28 VPWR sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.36e+06u l=150000u
X540 a_2454_3868# en29_b a_301_3864# VPWR sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.36e+06u l=150000u
X541 out en14_b a_2454_23173# VPWR sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.36e+06u l=150000u
X542 a_2454_33469# en6_b out VPWR sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.36e+06u l=150000u
X543 a_2454_41191# en0_b out VPWR sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.36e+06u l=150000u
X544 in_13 en_b a_301_24456# VPWR sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.36e+06u l=150000u
X545 out a_2450_26946# a_2454_27034# VGND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X546 a_301_29604# en9_b a_2454_29608# VPWR sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.36e+06u l=150000u
X547 out en8_b a_2454_30895# VPWR sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.36e+06u l=150000u
X548 in_28 en a_301_5151# VGND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X549 in_17 en_b a_301_19308# VPWR sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.36e+06u l=150000u
X550 in_7 en_b a_301_32178# VPWR sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.36e+06u l=150000u
X551 a_301_15447# en_b in_20 VPWR sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.36e+06u l=150000u
X552 in_1 en_b a_301_39900# VPWR sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.36e+06u l=150000u
X553 in_22 en_b a_301_12873# VPWR sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.36e+06u l=150000u
X554 in_16 en_b a_301_20595# VPWR sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.36e+06u l=150000u
X555 VPWR en1_b a_2450_39816# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.6e+11p ps=2.52e+06u w=1e+06u l=150000u
X556 a_301_34752# en5_b a_2454_34756# VPWR sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.36e+06u l=150000u
X557 out a_2450_2493# a_2454_2581# VGND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X558 a_301_11586# en_b in_23 VPWR sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.36e+06u l=150000u
X559 in_13 en a_301_24456# VGND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X560 a_2454_11590# a_2450_11502# a_301_11586# VGND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X561 a_2454_14164# en21_b a_301_14160# VPWR sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.36e+06u l=150000u
X562 VGND en31_b a_2450_1206# VGND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.69e+11p ps=1.82e+06u w=650000u l=150000u
X563 a_2454_39904# a_2450_39816# out VGND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X564 in_22 en a_301_12873# VGND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X565 a_301_34752# a_2450_34668# a_2454_34756# VGND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X566 a_2454_3868# en29_b out VPWR sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.36e+06u l=150000u
X567 a_301_27030# en_b in_11 VPWR sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.36e+06u l=150000u
X568 a_301_29604# en in_9 VGND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X569 in_1 en a_301_39900# VGND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X570 out a_2450_5067# a_2454_5155# VGND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X571 a_301_10299# en24_b a_2454_10303# VPWR sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.36e+06u l=150000u
X572 in_29 en_b a_301_3864# VPWR sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.36e+06u l=150000u
X573 out en16_b a_2454_20599# VPWR sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.36e+06u l=150000u
X574 a_2454_11590# en23_b out VPWR sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.36e+06u l=150000u
X575 a_2454_32182# en7_b a_301_32178# VPWR sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.36e+06u l=150000u
X576 a_301_21882# en15_b a_2454_21886# VPWR sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.36e+06u l=150000u
X577 a_2454_39904# en1_b a_301_39900# VPWR sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.36e+06u l=150000u
X578 a_301_16734# en19_b a_2454_16738# VPWR sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.36e+06u l=150000u
X579 out en12_b a_2454_25747# VPWR sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.36e+06u l=150000u
X580 a_301_1290# a_2450_1206# a_2454_1294# VGND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X581 a_2454_9016# a_2450_8928# a_301_9012# VGND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X582 in_29 en a_301_3864# VGND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X583 a_2454_10303# a_2450_10215# out VGND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X584 a_301_2577# en_b in_30 VPWR sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.36e+06u l=150000u
X585 a_301_6438# en27_b a_2454_6442# VPWR sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.36e+06u l=150000u
X586 a_301_21882# a_2450_21798# a_2454_21886# VGND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X587 out a_2450_25659# a_2454_25747# VGND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X588 a_2454_23173# a_2450_23085# out VGND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X589 in_22 en_b a_301_12873# VPWR sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.36e+06u l=150000u
X590 a_2454_16738# a_2450_16650# out VGND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X591 VGND en4_b a_2450_35955# VGND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.69e+11p ps=1.82e+06u w=650000u l=150000u
X592 a_301_10299# en24_b a_2454_10303# VPWR sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.36e+06u l=150000u
X593 out a_2450_14076# a_2454_14164# VGND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X594 in_16 en_b a_301_20595# VPWR sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.36e+06u l=150000u
X595 a_2454_24460# a_2450_24372# out VGND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X596 a_301_1290# en_b in_31 VPWR sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.36e+06u l=150000u
X597 in_20 en a_301_15447# VGND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X598 a_301_29604# a_2450_29520# a_2454_29608# VGND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X599 a_2454_39904# a_2450_39816# a_301_39900# VGND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X600 out a_2450_15363# a_2454_15451# VGND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X601 a_301_37326# a_2450_37242# a_2454_37330# VGND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X602 a_301_14160# en in_21 VGND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X603 a_2454_5155# en28_b a_301_5151# VPWR sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.36e+06u l=150000u
X604 a_2454_12877# en22_b a_301_12873# VPWR sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.36e+06u l=150000u
X605 a_301_23169# en14_b a_2454_23173# VPWR sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.36e+06u l=150000u
X606 a_2454_28321# en10_b out VPWR sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.36e+06u l=150000u
X607 a_2454_33469# en6_b a_301_33465# VPWR sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.36e+06u l=150000u
X608 a_2454_2581# en30_b out VPWR sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.36e+06u l=150000u
X609 out en17_b a_2454_19312# VPWR sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.36e+06u l=150000u
X610 a_301_30891# en8_b a_2454_30895# VPWR sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.36e+06u l=150000u
X611 a_2454_41191# en0_b a_301_41187# VPWR sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.36e+06u l=150000u
X612 in_4 en a_301_36039# VGND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X613 in_27 en a_301_6438# VGND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X614 in_6 en_b a_301_33465# VPWR sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.36e+06u l=150000u
X615 in_22 en a_301_12873# VGND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X616 a_301_18021# en_b in_18 VPWR sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.36e+06u l=150000u
X617 a_301_19308# en_b in_17 VPWR sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.36e+06u l=150000u
X618 out a_2450_3780# a_2454_3868# VGND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X619 a_2454_10303# en24_b a_301_10299# VPWR sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.36e+06u l=150000u
X620 VPWR en19_b a_2450_16650# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.6e+11p ps=2.52e+06u w=1e+06u l=150000u
X621 a_301_9012# en_b in_25 VPWR sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.36e+06u l=150000u
X622 a_301_23169# en in_14 VGND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X623 a_2454_12877# a_2450_12789# a_301_12873# VGND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X624 a_301_18021# en in_18 VGND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X625 in_25 en a_301_9012# VGND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X626 out a_2450_6354# a_2454_6442# VGND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X627 a_2454_5155# en28_b out VPWR sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.36e+06u l=150000u
X628 a_301_28317# en_b in_10 VPWR sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.36e+06u l=150000u
X629 a_2454_28321# a_2450_28233# a_301_28317# VGND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X630 out a_2450_39816# a_2454_39904# VGND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X631 in_9 en a_301_29604# VGND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X632 a_2454_23173# a_2450_23085# a_301_23169# VGND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X633 a_301_2577# en30_b a_2454_2581# VPWR sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.36e+06u l=150000u
X634 a_301_14160# a_2450_14076# a_2454_14164# VGND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X635 out en21_b a_2454_14164# VPWR sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.36e+06u l=150000u
X636 a_301_2577# a_2450_2493# a_2454_2581# VGND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X637 VPWR en30_b a_2450_2493# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.6e+11p ps=2.52e+06u w=1e+06u l=150000u
X638 a_301_9012# a_2450_8928# a_2454_9016# VGND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X639 out en9_b a_2454_29608# VPWR sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.36e+06u l=150000u
X640 a_301_18021# en18_b a_2454_18025# VPWR sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.36e+06u l=150000u
X641 a_2454_20599# en16_b out VPWR sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.36e+06u l=150000u
X642 a_2454_28321# en10_b a_301_28317# VPWR sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.36e+06u l=150000u
X643 out a_2450_8928# a_2454_9016# VGND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X644 out en23_b a_2454_11590# VPWR sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.36e+06u l=150000u
X645 a_301_19308# en17_b a_2454_19312# VPWR sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.36e+06u l=150000u
X646 out en5_b a_2454_34756# VPWR sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.36e+06u l=150000u
X647 a_301_1290# en in_31 VGND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X648 a_2454_25747# en12_b out VPWR sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.36e+06u l=150000u
X649 in_26 en_b a_301_7725# VPWR sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.36e+06u l=150000u
X650 a_301_38613# en2_b a_2454_38617# VPWR sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.36e+06u l=150000u
X651 a_301_34752# en_b in_5 VPWR sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.36e+06u l=150000u
X652 a_2454_11590# a_2450_11502# out VGND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X653 VGND en13_b a_2450_24372# VGND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.69e+11p ps=1.82e+06u w=650000u l=150000u
X654 a_301_6438# en_b in_27 VPWR sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.36e+06u l=150000u
X655 a_2454_6442# a_2450_6354# a_301_6438# VGND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X656 out a_2450_10215# a_2454_10303# VGND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X657 VGND en7_b a_2450_32094# VGND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.69e+11p ps=1.82e+06u w=650000u l=150000u
X658 out a_2450_34668# a_2454_34756# VGND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X659 a_2454_19312# a_2450_19224# out VGND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X660 a_301_14160# a_2450_14076# a_2454_14164# VGND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X661 a_2454_25747# a_2450_25659# out VGND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X662 in_26 en a_301_7725# VGND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X663 a_301_5151# en in_28 VGND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X664 a_2454_1294# en31_b a_301_1290# VPWR sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.36e+06u l=150000u
X665 out a_2450_23085# a_2454_23173# VGND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X666 out a_2450_16650# a_2454_16738# VGND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X667 a_301_38613# a_2450_38529# a_2454_38617# VGND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X668 in_13 en a_301_24456# VGND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X669 a_301_34752# en in_5 VGND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X670 out en26_b a_2454_7729# VPWR sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.36e+06u l=150000u
X671 a_301_15447# en in_20 VGND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X672 a_301_19308# en17_b a_2454_19312# VPWR sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.36e+06u l=150000u
X673 a_2454_16738# en19_b a_301_16734# VPWR sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.36e+06u l=150000u
X674 out en10_b a_2454_28321# VPWR sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.36e+06u l=150000u
X675 a_2454_1294# a_2450_1206# out VGND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X676 a_301_30891# en in_8 VGND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X677 a_301_11586# en in_23 VGND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X678 a_2454_14164# a_2450_14076# a_301_14160# VGND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X679 in_18 en_b a_301_18021# VPWR sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.36e+06u l=150000u
X680 a_2454_6442# en27_b out VPWR sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.36e+06u l=150000u
X681 a_301_19308# en in_17 VGND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X682 in_9 en a_301_29604# VGND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X683 a_2454_1294# en31_b out VPWR sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.36e+06u l=150000u
X684 a_301_27030# en in_11 VGND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X685 a_2454_19312# en17_b a_301_19308# VPWR sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.36e+06u l=150000u
X686 out a_2450_7641# a_2454_7729# VGND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X687 a_2454_29608# a_2450_29520# a_301_29604# VGND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X688 a_301_39900# a_2450_39816# a_2454_39904# VGND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X689 a_2454_11590# a_2450_11502# a_301_11586# VGND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X690 a_2454_2581# en30_b a_301_2577# VPWR sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.36e+06u l=150000u
X691 a_301_10299# a_2450_10215# a_2454_10303# VGND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X692 out en24_b a_2454_10303# VPWR sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.36e+06u l=150000u
X693 a_301_41187# a_2450_41103# a_2454_41191# VGND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X694 a_2454_32182# a_2450_32094# a_301_32178# VGND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X695 a_2454_32182# en7_b out VPWR sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.36e+06u l=150000u
X696 a_301_3864# a_2450_3780# a_2454_3868# VGND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X697 a_2454_39904# en1_b out VPWR sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.36e+06u l=150000u
X698 a_2454_12877# en22_b out VPWR sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.36e+06u l=150000u
X699 out en14_b a_2454_23173# VPWR sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.36e+06u l=150000u
X700 a_2454_33469# en6_b out VPWR sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.36e+06u l=150000u
X701 out en8_b a_2454_30895# VPWR sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.36e+06u l=150000u
X702 a_2454_41191# en0_b out VPWR sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.36e+06u l=150000u
X703 in_25 en_b a_301_9012# VPWR sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.36e+06u l=150000u
X704 a_2454_14164# en21_b out VPWR sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.36e+06u l=150000u
X705 in_7 en_b a_301_32178# VPWR sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.36e+06u l=150000u
X706 in_30 en_b a_301_2577# VPWR sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.36e+06u l=150000u
X707 in_1 en_b a_301_39900# VPWR sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.36e+06u l=150000u
X708 in_22 en_b a_301_12873# VPWR sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.36e+06u l=150000u
X709 a_301_27030# en11_b a_2454_27034# VPWR sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.36e+06u l=150000u
X710 a_2454_29608# en9_b out VPWR sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.36e+06u l=150000u
X711 a_2454_37330# en3_b a_301_37326# VPWR sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.36e+06u l=150000u
X712 in_16 en_b a_301_20595# VPWR sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.36e+06u l=150000u
X713 a_301_23169# en_b in_14 VPWR sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.36e+06u l=150000u
X714 a_301_2577# en in_30 VGND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X715 a_301_30891# en_b in_8 VPWR sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.36e+06u l=150000u
X716 VGND en16_b a_2450_20511# VGND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.69e+11p ps=1.82e+06u w=650000u l=150000u
X717 a_2454_34756# en5_b out VPWR sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.36e+06u l=150000u
X718 a_301_6438# a_2450_6354# a_2454_6442# VGND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X719 a_2454_12877# a_2450_12789# out VGND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X720 VGND en12_b a_2450_25659# VGND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.69e+11p ps=1.82e+06u w=650000u l=150000u
X721 a_2454_7729# a_2450_7641# a_301_7725# VGND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X722 a_301_10299# a_2450_10215# a_2454_10303# VGND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X723 out a_2450_11502# a_2454_11590# VGND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X724 in_22 en a_301_12873# VGND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X725 a_2454_28321# a_2450_28233# out VGND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X726 a_301_6438# en in_27 VGND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X727 a_2454_5155# a_2450_5067# a_301_5151# VGND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X728 in_18 en_b a_301_18021# VPWR sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.36e+06u l=150000u
X729 a_301_23169# a_2450_23085# a_2454_23173# VGND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X730 a_2454_34756# a_2450_34668# out VGND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X731 a_2454_2581# a_2450_2493# out VGND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X732 out a_2450_19224# a_2454_19312# VGND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X733 in_6 en a_301_33465# VGND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X734 out en25_b a_2454_9016# VPWR sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.36e+06u l=150000u
X735 a_301_18021# en in_18 VGND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X736 a_2454_10303# a_2450_10215# a_301_10299# VGND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X737 a_2454_18025# en18_b a_301_18021# VPWR sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.36e+06u l=150000u
X738 a_301_28317# en10_b a_2454_28321# VPWR sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.36e+06u l=150000u
X739 VPWR en6_b a_2450_33381# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.6e+11p ps=2.52e+06u w=1e+06u l=150000u
X740 a_301_9012# en in_25 VGND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X741 VPWR en2_b a_2450_38529# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.6e+11p ps=2.52e+06u w=1e+06u l=150000u
X742 a_2454_36043# en4_b VGND VGND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X743 a_2454_12877# en22_b a_301_12873# VPWR sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.36e+06u l=150000u
X744 a_301_28317# en in_10 VGND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X745 a_2454_5155# a_2450_5067# out VGND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X746 a_301_3864# en_b in_29 VPWR sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.36e+06u l=150000u
X747 a_301_7725# en26_b a_2454_7729# VPWR sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.36e+06u l=150000u
X748 a_2454_12877# a_2450_12789# a_301_12873# VGND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X749 a_301_2577# a_2450_2493# a_2454_2581# VGND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X750 out a_2450_14076# a_2454_14164# VGND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X751 a_2454_10303# en24_b out VPWR sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.36e+06u l=150000u
X752 a_2454_33469# a_2450_33381# a_301_33465# VGND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X753 a_301_18021# a_2450_17937# a_2454_18025# VGND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X754 a_301_3864# en in_29 VGND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X755 in_31 en a_301_1290# VGND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X756 a_301_15447# en20_b a_2454_15451# VPWR sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.36e+06u l=150000u
X757 a_2454_28321# a_2450_28233# a_301_28317# VGND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X758 a_301_19308# a_2450_19224# a_2454_19312# VGND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X759 out en17_b a_2454_19312# VPWR sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.36e+06u l=150000u
X760 out en7_b a_2454_32182# VPWR sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.36e+06u l=150000u
X761 out en1_b a_2454_39904# VPWR sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.36e+06u l=150000u
X762 out en22_b a_2454_12877# VPWR sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.36e+06u l=150000u
X763 a_2454_16738# en19_b out VPWR sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.36e+06u l=150000u
X764 in_6 en_b a_301_33465# VPWR sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.36e+06u l=150000u
X765 a_2454_23173# en14_b out VPWR sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.36e+06u l=150000u
X766 out en6_b a_2454_33469# VPWR sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.36e+06u l=150000u
X767 a_2454_29608# en9_b a_301_29604# VPWR sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.36e+06u l=150000u
X768 a_2454_30895# en8_b out VPWR sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.36e+06u l=150000u
X769 out en0_b a_2454_41191# VPWR sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.36e+06u l=150000u
X770 a_301_24456# en_b in_13 VPWR sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.36e+06u l=150000u
X771 in_27 en_b a_301_6438# VPWR sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.36e+06u l=150000u
X772 in_15 en_b a_301_21882# VPWR sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.36e+06u l=150000u
X773 a_301_32178# en_b in_7 VPWR sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.36e+06u l=150000u
X774 in_9 en_b a_301_29604# VPWR sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.36e+06u l=150000u
X775 a_301_39900# en_b in_1 VPWR sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.36e+06u l=150000u
X776 VGND en15_b a_2450_21798# VGND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.69e+11p ps=1.82e+06u w=650000u l=150000u
X777 a_2454_34756# en5_b a_301_34752# VPWR sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.36e+06u l=150000u
X778 a_301_7725# a_2450_7641# a_2454_7729# VGND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X779 a_301_11586# a_2450_11502# a_2454_11590# VGND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X780 out a_2450_12789# a_2454_12877# VGND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X781 a_301_30891# en in_8 VGND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X782 in_15 en a_301_21882# VGND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X783 a_301_41187# en_b in_0 VPWR sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.36e+06u l=150000u
X784 a_2454_29608# a_2450_29520# out VGND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X785 a_2454_41191# a_2450_41103# a_301_41187# VGND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X786 out a_2450_39816# a_2454_39904# VGND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X787 a_301_36039# en_b in_4 VPWR sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.36e+06u l=150000u
X788 a_2454_34756# a_2450_34668# a_301_34752# VGND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X789 a_2454_3868# a_2450_3780# out VGND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X790 a_301_16734# en_b in_19 VPWR sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.36e+06u l=150000u
X791 a_301_19308# a_2450_19224# a_2454_19312# VGND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X792 out a_2450_28233# a_2454_28321# VGND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X793 a_301_19308# en in_17 VGND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X794 a_301_39900# en in_1 VGND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X795 in_9 en a_301_29604# VGND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X796 in_18 en a_301_18021# VGND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X797 a_301_3864# en29_b a_2454_3868# VPWR sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.36e+06u l=150000u
X798 a_2454_6442# a_2450_6354# out VGND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X799 a_301_16734# en in_19 VGND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X800 a_2454_37330# en3_b VGND VGND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X801 a_2454_19312# a_2450_19224# a_301_19308# VGND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X802 a_2454_21886# en15_b a_301_21882# VPWR sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.36e+06u l=150000u
X803 a_301_32178# en7_b a_2454_32182# VPWR sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.36e+06u l=150000u
X804 a_2454_16738# en19_b a_301_16734# VPWR sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.36e+06u l=150000u
X805 a_301_39900# en1_b a_2454_39904# VPWR sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.36e+06u l=150000u
X806 VPWR en29_b a_2450_3780# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.6e+11p ps=2.52e+06u w=1e+06u l=150000u
X807 a_2454_2581# a_2450_2493# a_301_2577# VGND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X808 out a_2450_10215# a_2454_10303# VGND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X809 a_2454_3868# en29_b VGND VGND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X810 a_301_9012# en25_b a_2454_9016# VPWR sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.36e+06u l=150000u
X811 a_301_30891# a_2450_30807# a_2454_30895# VGND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X812 a_301_3864# a_2450_3780# a_2454_3868# VGND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X813 a_2454_21886# a_2450_21798# a_301_21882# VGND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X814 a_2454_32182# a_2450_32094# out VGND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X815 out a_2450_23085# a_2454_23173# VGND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X816 in_25 en a_301_9012# VGND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X817 a_301_7725# en_b in_26 VPWR sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.36e+06u l=150000u
X818 a_2454_14164# a_2450_14076# out VGND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X819 in_30 en a_301_2577# VGND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X820 a_2454_29608# a_2450_29520# a_301_29604# VGND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X821 a_301_27030# a_2450_26946# a_2454_27034# VGND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X822 a_2454_37330# a_2450_37242# a_301_37326# VGND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X823 a_2454_37330# en3_b out VPWR sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.36e+06u l=150000u
X824 a_301_32178# en7_b a_2454_32182# VPWR sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.36e+06u l=150000u
X825 a_301_39900# en1_b a_2454_39904# VPWR sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.36e+06u l=150000u
X826 a_301_12873# en22_b a_2454_12877# VPWR sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.36e+06u l=150000u
X827 a_2454_18025# en18_b out VPWR sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.36e+06u l=150000u
X828 out en10_b a_2454_28321# VPWR sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.36e+06u l=150000u
X829 a_2454_23173# en14_b a_301_23169# VPWR sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.36e+06u l=150000u
X830 a_2454_19312# en17_b out VPWR sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.36e+06u l=150000u
X831 a_2454_30895# en8_b a_301_30891# VPWR sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.36e+06u l=150000u
X832 a_301_36039# en in_4 VGND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X833 out en19_b a_2454_16738# VPWR sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.36e+06u l=150000u
X834 a_301_33465# en_b in_6 VPWR sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.36e+06u l=150000u
X835 in_18 en_b a_301_18021# VPWR sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.36e+06u l=150000u
X836 a_301_7725# en in_26 VGND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X837 a_301_32178# en in_7 VGND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X838 a_2454_7729# en26_b out VPWR sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.36e+06u l=150000u
X839 in_2 en_b a_301_38613# VPWR sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.36e+06u l=150000u
X840 a_301_12873# a_2450_12789# a_2454_12877# VGND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X841 in_18 en a_301_18021# VGND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X842 a_2454_32182# en7_b a_301_32178# VPWR sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.36e+06u l=150000u
X843 a_2454_39904# en1_b a_301_39900# VPWR sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.36e+06u l=150000u
X844 out a_2450_1206# a_2454_1294# VGND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X845 out a_2450_8928# a_2454_9016# VGND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X846 in_8 en a_301_30891# VGND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X847 a_301_37326# en_b in_3 VPWR sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.36e+06u l=150000u
X848 a_2454_18025# a_2450_17937# a_301_18021# VGND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X849 a_301_28317# a_2450_28233# a_2454_28321# VGND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X850 out a_2450_29520# a_2454_29608# VGND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X851 a_2454_39904# a_2450_39816# out VGND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X852 a_2454_3868# en29_b a_301_3864# VPWR sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.36e+06u l=150000u
X853 out en27_b a_2454_6442# VPWR sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.36e+06u l=150000u
X854 in_2 en a_301_38613# VGND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X855 in_17 en a_301_19308# VGND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X856 a_2454_25747# en12_b VGND VGND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X857 a_301_5151# en28_b a_2454_5155# VPWR sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.36e+06u l=150000u
X858 a_2454_7729# a_2450_7641# out VGND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X859 a_2454_29608# en9_b out VPWR sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.36e+06u l=150000u
X860 a_2454_18025# en18_b a_301_18021# VPWR sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.36e+06u l=150000u
X861 a_2454_34756# en5_b out VPWR sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.36e+06u l=150000u
X862 a_301_7725# en26_b a_2454_7729# VPWR sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.36e+06u l=150000u
X863 VPWR en26_b a_2450_7641# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.6e+11p ps=2.52e+06u w=1e+06u l=150000u
X864 a_2454_3868# a_2450_3780# a_301_3864# VGND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X865 a_2454_38617# en2_b a_301_38613# VPWR sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.36e+06u l=150000u
X866 a_301_9012# en_b in_25 VPWR sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.36e+06u l=150000u
X867 out a_2450_11502# a_2454_11590# VGND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X868 VGND en21_b a_2450_14076# VGND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.69e+11p ps=1.82e+06u w=650000u l=150000u
X869 a_2454_10303# a_2450_10215# out VGND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X870 a_2454_33469# a_2450_33381# out VGND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X871 a_301_2577# en_b in_30 VPWR sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.36e+06u l=150000u
X872 a_301_15447# a_2450_15363# a_2454_15451# VGND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X873 a_2454_41191# a_2450_41103# out VGND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X874 a_2454_34756# a_2450_34668# out VGND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X875 out a_2450_19224# a_2454_19312# VGND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X876 out a_2450_32094# a_2454_32182# VGND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X877 in_6 en a_301_33465# VGND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X878 a_2454_23173# a_2450_23085# out VGND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X879 a_301_24456# en in_13 VGND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X880 a_2454_38617# a_2450_38529# a_301_38613# VGND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X881 in_23 en_b a_301_11586# VPWR sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.36e+06u l=150000u
X882 out en3_b a_2454_37330# VPWR sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.36e+06u l=150000u
X883 out en18_b a_2454_18025# VPWR sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.36e+06u l=150000u
X884 a_301_16734# en19_b a_2454_16738# VPWR sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.36e+06u l=150000u
X885 a_301_20595# en in_16 VGND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X886 a_2454_28321# en10_b out VPWR sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.36e+06u l=150000u
X887 a_301_36039# en_b in_4 VPWR sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.36e+06u l=150000u
X888 in_8 en a_301_30891# VGND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X889 a_2454_2581# en30_b out VPWR sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.36e+06u l=150000u
X890 in_11 en_b a_301_27030# VPWR sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.36e+06u l=150000u
X891 VPWR en5_b a_2450_34668# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.6e+11p ps=2.52e+06u w=1e+06u l=150000u
X892 a_2454_9016# en25_b out VPWR sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.36e+06u l=150000u
X893 a_301_41187# en in_0 VGND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X894 in_17 en a_301_19308# VGND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X895 a_2454_30895# a_2450_30807# a_301_30891# VGND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X896 a_301_29604# a_2450_29520# a_2454_29608# VGND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X897 a_2454_39904# a_2450_39816# a_301_39900# VGND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X898 a_2454_5155# en28_b a_301_5151# VPWR sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.36e+06u l=150000u
X899 a_301_1290# en31_b a_2454_1294# VPWR sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.36e+06u l=150000u
X900 a_2454_41191# a_2450_41103# a_301_41187# VGND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X901 out en7_b a_2454_32182# VPWR sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.36e+06u l=150000u
X902 a_2454_21886# en15_b out VPWR sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.36e+06u l=150000u
X903 a_301_32178# a_2450_32094# a_2454_32182# VGND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X904 out en1_b a_2454_39904# VPWR sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.36e+06u l=150000u
X905 a_301_11586# en23_b a_2454_11590# VPWR sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.36e+06u l=150000u
X906 out en22_b a_2454_12877# VPWR sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.36e+06u l=150000u
X907 a_2454_7729# en26_b a_301_7725# VPWR sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.36e+06u l=150000u
X908 a_2454_23173# en14_b out VPWR sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.36e+06u l=150000u
X909 a_2454_30895# en8_b out VPWR sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.36e+06u l=150000u
X910 a_301_36039# en4_b a_2454_36043# VPWR sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.36e+06u l=150000u
X911 in_15 en_b a_301_21882# VPWR sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.36e+06u l=150000u
X912 in_9 en_b a_301_29604# VPWR sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.36e+06u l=150000u
X913 a_301_9012# en25_b a_2454_9016# VPWR sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.36e+06u l=150000u
X914 a_301_12873# en_b in_22 VPWR sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.36e+06u l=150000u
X915 a_2454_27034# en11_b a_301_27030# VPWR sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.36e+06u l=150000u
X916 out en9_b a_2454_29608# VPWR sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.36e+06u l=150000u
X917 a_301_37326# en3_b a_2454_37330# VPWR sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.36e+06u l=150000u
X918 a_301_20595# en_b in_16 VPWR sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.36e+06u l=150000u
X919 a_301_9012# a_2450_8928# a_2454_9016# VGND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X920 VGND en24_b a_2450_10215# VGND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.69e+11p ps=1.82e+06u w=650000u l=150000u
X921 out en5_b a_2454_34756# VPWR sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.36e+06u l=150000u
X922 a_2454_21886# a_2450_21798# out VGND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X923 in_26 en_b a_301_7725# VPWR sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.36e+06u l=150000u
X924 a_301_1290# en in_31 VGND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X925 out a_2450_12789# a_2454_12877# VGND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X926 in_15 en a_301_21882# VGND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X927 a_2454_11590# a_2450_11502# out VGND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X928 a_301_12873# en in_22 VGND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X929 a_301_16734# a_2450_16650# a_2454_16738# VGND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X930 a_2454_37330# a_2450_37242# out VGND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X931 out a_2450_33381# a_2454_33469# VGND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X932 a_301_6438# en_b in_27 VPWR sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.36e+06u l=150000u
X933 a_2454_18025# a_2450_17937# out VGND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X934 a_301_32178# a_2450_32094# a_2454_32182# VGND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X935 out a_2450_28233# a_2454_28321# VGND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X936 out a_2450_41103# a_2454_41191# VGND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X937 a_2454_23173# a_2450_23085# a_301_23169# VGND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X938 out a_2450_34668# a_2454_34756# VGND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X939 a_301_32178# en in_7 VGND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X940 a_2454_19312# a_2450_19224# out VGND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X941 a_301_33465# en in_6 VGND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X942 in_26 en a_301_7725# VGND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X943 in_14 en a_301_23169# VGND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X944 in_18 en a_301_18021# VGND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X945 a_301_37326# en3_b a_2454_37330# VPWR sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.36e+06u l=150000u
X946 a_301_18021# en18_b a_2454_18025# VPWR sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.36e+06u l=150000u
X947 VPWR en14_b a_2450_23085# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.6e+11p ps=2.52e+06u w=1e+06u l=150000u
X948 a_2454_28321# en10_b a_301_28317# VPWR sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.36e+06u l=150000u
X949 a_301_37326# en_b in_3 VPWR sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.36e+06u l=150000u
X950 in_10 en_b a_301_28317# VPWR sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.36e+06u l=150000u
X951 a_2454_32182# a_2450_32094# a_301_32178# VGND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X952 in_4 en_b a_301_36039# VPWR sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.36e+06u l=150000u
X953 a_2454_1294# a_2450_1206# out VGND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X954 a_301_37326# en in_3 VGND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X955 a_2454_37330# en3_b a_301_37326# VPWR sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.36e+06u l=150000u
X956 a_2454_3868# en29_b a_301_3864# VPWR sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.36e+06u l=150000u
X957 a_2454_6442# en27_b out VPWR sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.36e+06u l=150000u
X958 a_2454_1294# en31_b a_301_1290# VPWR sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.36e+06u l=150000u
X959 out a_2450_6354# a_2454_6442# VGND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X960 a_301_5151# a_2450_5067# a_2454_5155# VGND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X961 a_301_24456# en13_b a_2454_24460# VPWR sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.36e+06u l=150000u
X962 a_301_33465# a_2450_33381# a_2454_33469# VGND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X963 a_2454_18025# a_2450_17937# a_301_18021# VGND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X964 a_2454_15451# en20_b a_301_15447# VPWR sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.36e+06u l=150000u
X965 a_2454_9016# en25_b a_301_9012# VPWR sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.36e+06u l=150000u
X966 out en15_b a_2454_21886# VPWR sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.36e+06u l=150000u
X967 a_2454_32182# en7_b out VPWR sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.36e+06u l=150000u
X968 out en19_b a_2454_16738# VPWR sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.36e+06u l=150000u
X969 a_2454_39904# en1_b out VPWR sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.36e+06u l=150000u
X970 a_2454_12877# en22_b out VPWR sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.36e+06u l=150000u
X971 out en14_b a_2454_23173# VPWR sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.36e+06u l=150000u
X972 out en8_b a_2454_30895# VPWR sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.36e+06u l=150000u
X973 a_2454_38617# en2_b out VPWR sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.36e+06u l=150000u
X974 a_301_9012# en in_25 VGND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X975 a_301_21882# en_b in_15 VPWR sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.36e+06u l=150000u
X976 a_301_29604# en_b in_9 VPWR sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.36e+06u l=150000u
X977 in_2 en_b a_301_38613# VPWR sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.36e+06u l=150000u
X978 a_301_2577# en in_30 VGND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X979 a_2454_30895# a_2450_30807# out VGND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X980 out a_2450_21798# a_2454_21886# VGND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X981 a_2454_11590# a_2450_11502# a_301_11586# VGND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X982 a_2454_12877# a_2450_12789# out VGND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X983 VGND en17_b a_2450_19224# VGND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.69e+11p ps=1.82e+06u w=650000u l=150000u
X984 a_301_20595# en in_16 VGND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X985 in_8 en a_301_30891# VGND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X986 in_23 en a_301_11586# VGND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X987 a_2454_38617# a_2450_38529# out VGND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X988 a_301_21882# en in_15 VGND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X989 a_301_33465# a_2450_33381# a_2454_33469# VGND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X990 in_4 en_b a_301_36039# VPWR sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.36e+06u l=150000u
X991 a_301_25743# en_b in_12 VPWR sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.36e+06u l=150000u
X992 out a_2450_29520# a_2454_29608# VGND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X993 a_301_41187# a_2450_41103# a_2454_41191# VGND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X994 a_2454_39904# a_2450_39816# out VGND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X995 out a_2450_37242# a_2454_37330# VGND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X996 VPWR en23_b a_2450_11502# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.6e+11p ps=2.52e+06u w=1e+06u l=150000u
X997 out a_2450_17937# a_2454_18025# VGND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X998 in_2 en a_301_38613# VGND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X999 a_2454_28321# a_2450_28233# out VGND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X1000 in_17 en a_301_19308# VGND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X1001 a_301_29604# en in_9 VGND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X1002 in_7 en a_301_32178# VGND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X1003 a_2454_2581# a_2450_2493# out VGND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X1004 in_11 en a_301_27030# VGND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X1005 a_2454_36043# en4_b a_301_36039# VPWR sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.36e+06u l=150000u
X1006 a_2454_14164# en21_b VGND VGND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X1007 a_2454_9016# a_2450_8928# out VGND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X1008 a_301_25743# en in_12 VGND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X1009 a_2454_33469# a_2450_33381# a_301_33465# VGND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X1010 in_3 en_b a_301_37326# VPWR sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.36e+06u l=150000u
X1011 a_301_3864# en29_b a_2454_3868# VPWR sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.36e+06u l=150000u
X1012 a_301_21882# en15_b a_2454_21886# VPWR sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.36e+06u l=150000u
X1013 out en29_b a_2454_3868# VPWR sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.36e+06u l=150000u
X1014 a_2454_5155# en28_b a_301_5151# VPWR sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.36e+06u l=150000u
X1015 out a_2450_7641# a_2454_7729# VGND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X1016 a_2454_5155# a_2450_5067# a_301_5151# VGND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X1017 a_301_20595# a_2450_20511# a_2454_20599# VGND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X1018 a_2454_30895# a_2450_30807# a_301_30891# VGND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X1019 a_301_21882# a_2450_21798# a_2454_21886# VGND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X1020 out a_2450_32094# a_2454_32182# VGND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X1021 a_2454_23173# a_2450_23085# out VGND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X1022 in_23 en_b a_301_11586# VPWR sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.36e+06u l=150000u
X1023 a_301_36039# a_2450_35955# a_2454_36043# VGND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X1024 a_2454_9016# en25_b VGND VGND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X1025 a_301_33465# en6_b a_2454_33469# VPWR sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.36e+06u l=150000u
X1026 a_301_41187# en0_b a_2454_41191# VPWR sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.36e+06u l=150000u
X1027 a_301_9012# a_2450_8928# a_2454_9016# VGND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X1028 a_2454_27034# a_2450_26946# a_301_27030# VGND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X1029 a_2454_27034# en11_b out VPWR sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.36e+06u l=150000u
X1030 out en3_b a_2454_37330# VPWR sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.36e+06u l=150000u
X1031 a_301_37326# a_2450_37242# a_2454_37330# VGND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X1032 a_301_21882# en15_b a_2454_21886# VPWR sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.36e+06u l=150000u
X1033 out en18_b a_2454_18025# VPWR sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.36e+06u l=150000u
X1034 a_2454_12877# en22_b a_301_12873# VPWR sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.36e+06u l=150000u
X1035 a_2454_28321# en10_b out VPWR sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.36e+06u l=150000u
X1036 in_30 en_b a_301_2577# VPWR sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.36e+06u l=150000u
X1037 a_2454_16738# en19_b out VPWR sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.36e+06u l=150000u
X1038 in_11 en_b a_301_27030# VPWR sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.36e+06u l=150000u
X1039 a_301_18021# en_b in_18 VPWR sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.36e+06u l=150000u
X1040 out en2_b a_2454_38617# VPWR sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.36e+06u l=150000u
X1041 in_7 en a_301_32178# VGND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X1042 a_301_14160# en_b in_21 VPWR sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.36e+06u l=150000u
X1043 a_301_21882# a_2450_21798# a_2454_21886# VGND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X1044 a_301_38613# en_b in_2 VPWR sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.36e+06u l=150000u
X1045 in_28 en_b a_301_5151# VPWR sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.36e+06u l=150000u
X1046 a_2454_12877# a_2450_12789# a_301_12873# VGND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X1047 a_2454_21886# en15_b a_301_21882# VPWR sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.36e+06u l=150000u
X1048 out a_2450_30807# a_2454_30895# VGND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X1049 in_16 en a_301_20595# VGND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X1050 in_3 en_b a_301_37326# VPWR sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.36e+06u l=150000u
X1051 out en30_b a_2454_2581# VPWR sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.36e+06u l=150000u
X1052 out a_2450_38529# a_2454_38617# VGND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X1053 a_301_37326# a_2450_37242# a_2454_37330# VGND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X1054 a_301_34752# en_b in_5 VPWR sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.36e+06u l=150000u
X1055 a_2454_24460# en13_b a_301_24456# VPWR sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.36e+06u l=150000u
X1056 a_2454_10303# en24_b VGND VGND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X1057 a_301_18021# a_2450_17937# a_2454_18025# VGND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X1058 a_2454_28321# a_2450_28233# a_301_28317# VGND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X1059 a_2454_29608# a_2450_29520# out VGND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X1060 out a_2450_39816# a_2454_39904# VGND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X1061 a_301_37326# en in_3 VGND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X1062 a_301_38613# en in_2 VGND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X1063 a_2454_3868# a_2450_3780# out VGND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X1064 a_2454_21886# a_2450_21798# a_301_21882# VGND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X1065 in_10 en a_301_28317# VGND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X1066 a_2454_15451# en20_b VGND VGND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X1067 a_301_34752# en in_5 VGND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X1068 a_2454_37330# a_2450_37242# a_301_37326# VGND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X1069 a_301_5151# en28_b a_2454_5155# VPWR sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.36e+06u l=150000u
X1070 a_2454_1294# en31_b a_301_1290# VPWR sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.36e+06u l=150000u
X1071 a_2454_6442# a_2450_6354# out VGND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X1072 out en28_b a_2454_5155# VPWR sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.36e+06u l=150000u
X1073 a_301_38613# en2_b a_2454_38617# VPWR sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.36e+06u l=150000u
X1074 a_2454_11590# a_2450_11502# out VGND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X1075 a_2454_2581# en30_b a_301_2577# VPWR sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.36e+06u l=150000u
X1076 a_301_24456# a_2450_24372# a_2454_24460# VGND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X1077 out a_2450_33381# a_2454_33469# VGND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X1078 a_2454_15451# a_2450_15363# a_301_15447# VGND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X1079 a_2454_15451# en20_b out VPWR sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.36e+06u l=150000u
X1080 out a_2450_41103# a_2454_41191# VGND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X1081 a_2454_9016# a_2450_8928# a_301_9012# VGND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X1082 a_2454_32182# a_2450_32094# out VGND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X1083 in_14 en a_301_23169# VGND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X1084 out a_2450_23085# a_2454_23173# VGND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X1085 in_31 en a_301_1290# VGND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X1086 a_301_11586# en_b in_23 VPWR sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.36e+06u l=150000u
X1087 a_301_38613# a_2450_38529# a_2454_38617# VGND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X1088 a_2454_36043# en4_b out VPWR sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.36e+06u l=150000u
X1089 a_301_7725# en_b in_26 VPWR sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.36e+06u l=150000u
X1090 out en11_b a_2454_27034# VPWR sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.36e+06u l=150000u
X1091 a_2454_37330# en3_b out VPWR sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.36e+06u l=150000u
X1092 a_301_10299# en in_24 VGND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X1093 a_2454_16738# en19_b a_301_16734# VPWR sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.36e+06u l=150000u
X1094 a_2454_18025# en18_b out VPWR sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.36e+06u l=150000u
X1095 in_10 en_b a_301_28317# VPWR sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.36e+06u l=150000u
X1096 in_0 en_b a_301_41187# VPWR sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.36e+06u l=150000u
X1097 in_16 en a_301_20595# VGND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X1098 a_301_25743# en_b in_12 VPWR sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.36e+06u l=150000u
X1099 out en10_b a_2454_28321# VPWR sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.36e+06u l=150000u
X1100 in_4 en_b a_301_36039# VPWR sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.36e+06u l=150000u
X1101 in_27 en_b a_301_6438# VPWR sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.36e+06u l=150000u
X1102 a_301_10299# en_b in_24 VPWR sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.36e+06u l=150000u
X1103 in_19 en_b a_301_16734# VPWR sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.36e+06u l=150000u
X1104 a_301_27030# en_b in_11 VPWR sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.36e+06u l=150000u
X1105 a_301_38613# en2_b a_2454_38617# VPWR sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.36e+06u l=150000u
X1106 in_31 en_b a_301_1290# VPWR sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.36e+06u l=150000u
X1107 a_301_15447# en_b in_20 VPWR sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.36e+06u l=150000u
X1108 a_301_7725# en in_26 VGND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X1109 a_2454_20599# a_2450_20511# a_301_20595# VGND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X1110 a_301_23169# en_b in_14 VPWR sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.36e+06u l=150000u
X1111 a_301_30891# a_2450_30807# a_2454_30895# VGND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X1112 a_301_30891# en_b in_8 VPWR sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.36e+06u l=150000u
X1113 a_2454_7729# en26_b out VPWR sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.36e+06u l=150000u
X1114 a_301_25743# en in_12 VGND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X1115 in_19 en a_301_16734# VGND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X1116 a_301_38613# a_2450_38529# a_2454_38617# VGND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X1117 a_2454_36043# a_2450_35955# a_301_36039# VGND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X1118 out a_2450_1206# a_2454_1294# VGND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X1119 a_2454_38617# en2_b a_301_38613# VPWR sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.36e+06u l=150000u
X1120 a_2454_29608# a_2450_29520# a_301_29604# VGND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X1121 in_3 en a_301_37326# VGND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X1122 out en27_b a_2454_6442# VPWR sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.36e+06u l=150000u
X1123 a_301_1290# en31_b a_2454_1294# VPWR sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.36e+06u l=150000u
X1124 a_2454_19312# en17_b VGND VGND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X1125 a_301_20595# en16_b a_2454_20599# VPWR sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.36e+06u l=150000u
X1126 out en15_b a_2454_21886# VPWR sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.36e+06u l=150000u
X1127 out en31_b a_2454_1294# VPWR sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.36e+06u l=150000u
X1128 a_2454_11590# en23_b a_301_11586# VPWR sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.36e+06u l=150000u
X1129 a_2454_12877# en22_b out VPWR sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.36e+06u l=150000u
X1130 a_2454_38617# a_2450_38529# a_301_38613# VGND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X1131 a_2454_5155# a_2450_5067# a_301_5151# VGND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X1132 a_2454_7729# a_2450_7641# out VGND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X1133 a_301_25743# en12_b a_2454_25747# VPWR sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.36e+06u l=150000u
X1134 a_2454_36043# en4_b a_301_36039# VPWR sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.36e+06u l=150000u
X1135 a_301_27030# en11_b a_2454_27034# VPWR sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.36e+06u l=150000u
X1136 a_301_2577# en30_b a_2454_2581# VPWR sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.36e+06u l=150000u
X1137 out a_2450_21798# a_2454_21886# VGND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X1138 a_2454_12877# a_2450_12789# out VGND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X1139 in_23 en a_301_11586# VGND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X1140 a_301_25743# a_2450_25659# a_2454_25747# VGND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X1141 out a_2450_11502# a_2454_11590# VGND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X1142 a_2454_16738# a_2450_16650# a_301_16734# VGND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X1143 a_2454_27034# a_2450_26946# out VGND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X1144 out a_2450_37242# a_2454_37330# VGND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X1145 a_2454_24460# en13_b out VPWR sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.36e+06u l=150000u
X1146 a_2454_33469# a_2450_33381# out VGND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X1147 a_301_2577# en_b in_30 VPWR sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.36e+06u l=150000u
X1148 out a_2450_17937# a_2454_18025# VGND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X1149 out en20_b a_2454_15451# VPWR sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.36e+06u l=150000u
X1150 a_2454_28321# a_2450_28233# out VGND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X1151 a_2454_41191# a_2450_41103# out VGND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X1152 in_30 en a_301_2577# VGND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X1153 in_7 en a_301_32178# VGND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X1154 a_301_14160# en_b in_21 VPWR sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.36e+06u l=150000u
X1155 a_301_23169# en in_14 VGND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X1156 in_11 en a_301_27030# VGND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X1157 a_301_18021# en in_18 VGND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X1158 a_301_27030# en11_b a_2454_27034# VPWR sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.36e+06u l=150000u
X1159 out en4_b a_2454_36043# VPWR sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.36e+06u l=150000u
X1160 VPWR en22_b a_2450_12789# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.6e+11p ps=2.52e+06u w=1e+06u l=150000u
X1161 a_2454_18025# en18_b a_301_18021# VPWR sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.36e+06u l=150000u
X1162 in_3 en_b a_301_37326# VPWR sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.36e+06u l=150000u
X1163 a_301_5151# en_b in_28 VPWR sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.36e+06u l=150000u
X1164 a_301_14160# en in_21 VGND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X1165 a_301_28317# en_b in_10 VPWR sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.36e+06u l=150000u
X1166 in_28 en a_301_5151# VGND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X1167 in_12 en_b a_301_25743# VPWR sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.36e+06u l=150000u
X1168 in_3 en a_301_37326# VGND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X1169 out a_2450_2493# a_2454_2581# VGND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X1170 a_301_24456# en_b in_13 VPWR sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.36e+06u l=150000u
X1171 a_301_19308# en_b in_17 VPWR sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.36e+06u l=150000u
X1172 a_2454_9016# en25_b out VPWR sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.36e+06u l=150000u
X1173 a_2454_24460# a_2450_24372# a_301_24456# VGND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X1174 a_2454_27034# en11_b a_301_27030# VPWR sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.36e+06u l=150000u
X1175 VGND en27_b a_2450_6354# VGND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.69e+11p ps=1.82e+06u w=650000u l=150000u
X1176 in_12 en a_301_25743# VGND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X1177 a_301_5151# a_2450_5067# a_2454_5155# VGND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X1178 a_301_14160# en21_b a_2454_14164# VPWR sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.36e+06u l=150000u
X1179 a_2454_24460# en13_b a_301_24456# VPWR sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.36e+06u l=150000u
X1180 out a_2450_5067# a_2454_5155# VGND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X1181 a_301_15447# en20_b a_2454_15451# VPWR sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.36e+06u l=150000u
X1182 a_301_29604# en9_b a_2454_29608# VPWR sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.36e+06u l=150000u
X1183 a_301_39900# en in_1 VGND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X1184 a_2454_21886# en15_b out VPWR sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.36e+06u l=150000u
X1185 in_29 en_b a_301_3864# VPWR sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.36e+06u l=150000u
X1186 a_2454_16738# en19_b out VPWR sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.36e+06u l=150000u
X1187 out en22_b a_2454_12877# VPWR sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.36e+06u l=150000u
X1188 a_301_34752# en5_b a_2454_34756# VPWR sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.36e+06u l=150000u
X1189 out en2_b a_2454_38617# VPWR sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.36e+06u l=150000u
X1190 a_2454_2581# a_2450_2493# a_301_2577# VGND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X1191 a_2454_20599# a_2450_20511# out VGND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X1192 a_2454_15451# a_2450_15363# out VGND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X1193 out a_2450_30807# a_2454_30895# VGND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X1194 a_2454_21886# a_2450_21798# out VGND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X1195 in_29 en a_301_3864# VGND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X1196 a_301_1290# en in_31 VGND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X1197 out a_2450_12789# a_2454_12877# VGND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X1198 a_301_10299# en in_24 VGND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X1199 in_16 en a_301_20595# VGND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X1200 a_301_34752# a_2450_34668# a_2454_34756# VGND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X1201 a_301_30891# en in_8 VGND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X1202 out en29_b a_2454_3868# VPWR sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.36e+06u l=150000u
X1203 a_301_11586# en in_23 VGND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X1204 out a_2450_38529# a_2454_38617# VGND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X1205 a_301_10299# en_b in_24 VPWR sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.36e+06u l=150000u
X1206 a_2454_36043# a_2450_35955# out VGND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X1207 in_12 en_b a_301_25743# VPWR sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.36e+06u l=150000u
X1208 a_301_15447# en20_b a_2454_15451# VPWR sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.36e+06u l=150000u
X1209 a_2454_29608# a_2450_29520# out VGND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X1210 a_2454_41191# a_2450_41103# a_301_41187# VGND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X1211 out a_2450_26946# a_2454_27034# VGND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X1212 a_2454_37330# a_2450_37242# out VGND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X1213 a_301_6438# en_b in_27 VPWR sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.36e+06u l=150000u
X1214 a_2454_20599# en16_b a_301_20595# VPWR sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.36e+06u l=150000u
X1215 out en13_b a_2454_24460# VPWR sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.36e+06u l=150000u
X1216 a_301_15447# en_b in_20 VPWR sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.36e+06u l=150000u
X1217 a_2454_18025# a_2450_17937# out VGND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X1218 in_10 en a_301_28317# VGND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X1219 in_0 en a_301_41187# VGND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X1220 a_301_19308# en in_17 VGND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X1221 out a_2450_28233# a_2454_28321# VGND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X1222 a_301_1290# en_b in_31 VPWR sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.36e+06u l=150000u
X1223 in_21 en_b a_301_14160# VPWR sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.36e+06u l=150000u
X1224 a_301_27030# en in_11 VGND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X1225 a_301_36039# en4_b a_2454_36043# VPWR sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.36e+06u l=150000u
X1226 a_2454_25747# en12_b a_301_25743# VPWR sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.36e+06u l=150000u
X1227 VPWR en0_b a_2450_41103# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.6e+11p ps=2.52e+06u w=1e+06u l=150000u
X1228 a_2454_2581# en30_b out VPWR sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.36e+06u l=150000u
X1229 a_301_15447# en in_20 VGND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X1230 in_27 en a_301_6438# VGND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X1231 in_12 en a_301_25743# VGND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X1232 a_2454_15451# en20_b a_301_15447# VPWR sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.36e+06u l=150000u
X1233 out a_2450_3780# a_2454_3868# VGND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X1234 VGND en30_b a_2450_2493# VGND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.69e+11p ps=1.82e+06u w=650000u l=150000u
X1235 a_301_36039# en in_4 VGND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X1236 a_2454_25747# a_2450_25659# a_301_25743# VGND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X1237 a_2454_20599# a_2450_20511# a_301_20595# VGND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X1238 out a_2450_6354# a_2454_6442# VGND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X1239 a_301_10299# en24_b a_2454_10303# VPWR sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.36e+06u l=150000u
X1240 in_28 en_b a_301_5151# VPWR sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.36e+06u l=150000u
X1241 a_2454_11590# en23_b out VPWR sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.36e+06u l=150000u
X1242 a_2454_36043# a_2450_35955# a_301_36039# VGND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X1243 a_301_23169# en14_b a_2454_23173# VPWR sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.36e+06u l=150000u
X1244 a_2454_33469# en6_b a_301_33465# VPWR sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.36e+06u l=150000u
X1245 a_301_30891# en8_b a_2454_30895# VPWR sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.36e+06u l=150000u
X1246 a_2454_41191# en0_b a_301_41187# VPWR sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.36e+06u l=150000u
X1247 a_301_27030# a_2450_26946# a_2454_27034# VGND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X1248 out en11_b a_2454_27034# VPWR sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.36e+06u l=150000u
X1249 a_301_2577# a_2450_2493# a_2454_2581# VGND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X1250 a_2454_18025# en18_b out VPWR sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.36e+06u l=150000u
X1251 in_0 en_b a_301_41187# VPWR sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.36e+06u l=150000u
X1252 in_19 en_b a_301_16734# VPWR sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.36e+06u l=150000u
X1253 out en19_b a_2454_16738# VPWR sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.36e+06u l=150000u
X1254 a_2454_3868# a_2450_3780# a_301_3864# VGND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X1255 a_2454_38617# en2_b out VPWR sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.36e+06u l=150000u
X1256 a_2454_16738# a_2450_16650# out VGND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X1257 in_26 en_b a_301_7725# VPWR sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.36e+06u l=150000u
X1258 in_21 en_b a_301_14160# VPWR sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.36e+06u l=150000u
X1259 a_2454_24460# a_2450_24372# out VGND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X1260 a_2454_1294# a_2450_1206# a_301_1290# VGND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X1261 a_301_2577# en in_30 VGND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X1262 out a_2450_20511# a_2454_20599# VGND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X1263 VGND en3_b a_2450_37242# VGND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.69e+11p ps=1.82e+06u w=650000u l=150000u
X1264 out a_2450_15363# a_2454_15451# VGND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X1265 a_2454_30895# a_2450_30807# out VGND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X1266 in_19 en a_301_16734# VGND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X1267 out en28_b a_2454_5155# VPWR sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.36e+06u l=150000u
X1268 in_24 en a_301_10299# VGND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X1269 a_301_14160# en in_21 VGND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X1270 in_24 en_b a_301_10299# VPWR sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.36e+06u l=150000u
X1271 a_2454_14164# en21_b a_301_14160# VPWR sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.36e+06u l=150000u
X1272 a_301_27030# a_2450_26946# a_2454_27034# VGND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X1273 a_2454_38617# a_2450_38529# out VGND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X1274 a_2454_6442# en27_b a_301_6438# VPWR sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.36e+06u l=150000u
X1275 a_301_24456# en13_b a_2454_24460# VPWR sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.36e+06u l=150000u
X1276 out a_2450_35955# a_2454_36043# VGND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X1277 a_2454_18025# a_2450_17937# a_301_18021# VGND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X1278 in_26 en a_301_7725# VGND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X1279 out a_2450_29520# a_2454_29608# VGND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X1280 in_3 en a_301_37326# VGND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X1281 a_301_5151# en in_28 VGND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X1282 a_301_19308# en_b in_17 VPWR sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.36e+06u l=150000u
X1283 a_301_28317# en in_10 VGND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X1284 in_20 en_b a_301_15447# VPWR sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.36e+06u l=150000u
X1285 out en26_b a_2454_7729# VPWR sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.36e+06u l=150000u
X1286 a_2454_32182# en7_b VGND VGND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X1287 a_2454_1294# a_2450_1206# out VGND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X1288 a_301_24456# en in_13 VGND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X1289 a_2454_9016# a_2450_8928# out VGND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X1290 a_2454_27034# a_2450_26946# a_301_27030# VGND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X1291 a_301_3864# en29_b a_2454_3868# VPWR sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.36e+06u l=150000u
X1292 a_2454_6442# en27_b out VPWR sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.36e+06u l=150000u
X1293 out a_2450_7641# a_2454_7729# VGND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X1294 in_31 en_b a_301_1290# VPWR sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.36e+06u l=150000u
X1295 a_301_14160# a_2450_14076# a_2454_14164# VGND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X1296 a_2454_24460# a_2450_24372# a_301_24456# VGND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X1297 a_301_15447# a_2450_15363# a_2454_15451# VGND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X1298 out en20_b a_2454_15451# VPWR sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.36e+06u l=150000u
X1299 a_2454_41191# a_2450_41103# out VGND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X1300 a_2454_20599# en16_b out VPWR sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.36e+06u l=150000u
X1301 a_2454_7729# en26_b a_301_7725# VPWR sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.36e+06u l=150000u
X1302 out en23_b a_2454_11590# VPWR sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.36e+06u l=150000u
X1303 a_301_19308# en17_b a_2454_19312# VPWR sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.36e+06u l=150000u
X1304 a_2454_25747# en12_b out VPWR sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.36e+06u l=150000u
X1305 out en4_b a_2454_36043# VPWR sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.36e+06u l=150000u
X1306 a_301_3864# a_2450_3780# a_2454_3868# VGND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X1307 a_2454_27034# en11_b out VPWR sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.36e+06u l=150000u
X1308 in_25 en_b a_301_9012# VPWR sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.36e+06u l=150000u
X1309 in_24 en a_301_10299# VGND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X1310 out en18_b a_2454_18025# VPWR sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.36e+06u l=150000u
X1311 a_301_41187# en_b in_0 VPWR sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.36e+06u l=150000u
X1312 in_12 en_b a_301_25743# VPWR sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.36e+06u l=150000u
X1313 a_301_36039# en_b in_4 VPWR sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.36e+06u l=150000u
X1314 in_24 en_b a_301_10299# VPWR sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.36e+06u l=150000u
X1315 a_301_16734# en_b in_19 VPWR sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.36e+06u l=150000u
X1316 out en31_b a_2454_1294# VPWR sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.36e+06u l=150000u
X1317 a_301_32178# en_b in_7 VPWR sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.36e+06u l=150000u
X1318 in_20 en_b a_301_15447# VPWR sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.36e+06u l=150000u
X1319 a_2454_25747# a_2450_25659# out VGND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X1320 a_301_39900# en_b in_1 VPWR sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.36e+06u l=150000u
X1321 a_301_12873# en_b in_22 VPWR sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.36e+06u l=150000u
X1322 a_301_20595# a_2450_20511# a_2454_20599# VGND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X1323 VGND en2_b a_2450_38529# VGND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.69e+11p ps=1.82e+06u w=650000u l=150000u
X1324 a_301_15447# a_2450_15363# a_2454_15451# VGND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X1325 out a_2450_16650# a_2454_16738# VGND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X1326 a_301_20595# en_b in_16 VPWR sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.36e+06u l=150000u
X1327 a_2454_30895# a_2450_30807# a_301_30891# VGND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X1328 a_2454_10303# en24_b a_301_10299# VPWR sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.36e+06u l=150000u
X1329 a_301_15447# en in_20 VGND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X1330 out a_2450_24372# a_2454_24460# VGND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X1331 in_12 en a_301_25743# VGND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X1332 a_301_39900# a_2450_39816# a_2454_39904# VGND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X1333 a_301_16734# en in_19 VGND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X1334 in_21 en a_301_14160# VGND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X1335 a_301_36039# a_2450_35955# a_2454_36043# VGND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X1336 a_301_6438# en in_27 VGND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X1337 a_2454_2581# a_2450_2493# out VGND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X1338 a_301_12873# en in_22 VGND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X1339 a_2454_33469# en6_b VGND VGND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X1340 out en25_b a_2454_9016# VPWR sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.36e+06u l=150000u
X1341 a_2454_15451# a_2450_15363# a_301_15447# VGND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X1342 in_17 en_b a_301_19308# VPWR sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.36e+06u l=150000u
X1343 a_2454_20599# en16_b a_301_20595# VPWR sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.36e+06u l=150000u
X1344 a_301_11586# en23_b a_2454_11590# VPWR sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.36e+06u l=150000u
X1345 a_2454_25747# en12_b a_301_25743# VPWR sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.36e+06u l=150000u
X1346 a_301_5151# en28_b a_2454_5155# VPWR sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.36e+06u l=150000u
X1347 a_301_10299# a_2450_10215# a_2454_10303# VGND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X1348 in_28 en a_301_5151# VGND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X1349 a_301_3864# en_b in_29 VPWR sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.36e+06u l=150000u
X1350 a_2454_25747# a_2450_25659# a_301_25743# VGND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X1351 a_301_7725# en26_b a_2454_7729# VPWR sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.36e+06u l=150000u
X1352 a_301_16734# a_2450_16650# a_2454_16738# VGND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X1353 a_301_23169# a_2450_23085# a_2454_23173# VGND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X1354 a_2454_33469# en6_b out VPWR sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.36e+06u l=150000u
X1355 a_2454_41191# en0_b out VPWR sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.36e+06u l=150000u
X1356 a_2454_14164# en21_b out VPWR sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.36e+06u l=150000u
X1357 out a_2450_26946# a_2454_27034# VGND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X1358 out en13_b a_2454_24460# VPWR sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.36e+06u l=150000u
X1359 a_2454_18025# a_2450_17937# out VGND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X1360 in_0 en a_301_41187# VGND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X1361 a_2454_9016# en25_b a_301_9012# VPWR sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.36e+06u l=150000u
X1362 a_301_11586# en23_b a_2454_11590# VPWR sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.36e+06u l=150000u
X1363 a_2454_15451# en20_b out VPWR sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.36e+06u l=150000u
X1364 out a_2450_41103# a_2454_41191# VGND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X1365 a_301_32178# en in_7 VGND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X1366 out en16_b a_2454_20599# VPWR sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.36e+06u l=150000u
X1367 in_21 en_b a_301_14160# VPWR sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.36e+06u l=150000u
X1368 a_301_28317# en10_b a_2454_28321# VPWR sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.36e+06u l=150000u
X1369 a_301_3864# en in_29 VGND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X1370 a_301_7725# en_b in_26 VPWR sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.36e+06u l=150000u
X1371 out en12_b a_2454_25747# VPWR sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.36e+06u l=150000u
X1372 a_2454_36043# en4_b out VPWR sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.36e+06u l=150000u
X1373 a_2454_3868# en29_b out VPWR sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.36e+06u l=150000u
X1374 a_301_37326# en_b in_3 VPWR sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.36e+06u l=150000u
X1375 in_5 en_b a_301_34752# VPWR sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.36e+06u l=150000u
X1376 in_21 en a_301_14160# VGND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X1377 a_2454_11590# en23_b a_301_11586# VPWR sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.36e+06u l=150000u
X1378 out a_2450_5067# a_2454_5155# VGND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X1379 a_301_33465# en_b in_6 VPWR sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.36e+06u l=150000u
X1380 a_301_16734# a_2450_16650# a_2454_16738# VGND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X1381 a_301_7725# en in_26 VGND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X1382 a_2454_6442# a_2450_6354# a_301_6438# VGND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X1383 a_2454_14164# a_2450_14076# a_301_14160# VGND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X1384 in_17 en_b a_301_19308# VPWR sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.36e+06u l=150000u
X1385 a_301_24456# a_2450_24372# a_2454_24460# VGND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X1386 out a_2450_25659# a_2454_25747# VGND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X1387 out en30_b a_2454_2581# VPWR sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.36e+06u l=150000u
X1388 in_5 en a_301_34752# VGND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X1389 in_20 en a_301_15447# VGND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X1390 a_2454_21886# en15_b VGND VGND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X1391 a_2454_19312# en17_b a_301_19308# VPWR sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.36e+06u l=150000u
X1392 a_2454_3868# a_2450_3780# out VGND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X1393 a_2454_16738# a_2450_16650# a_301_16734# VGND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X1394 a_2454_14164# en21_b a_301_14160# VPWR sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.36e+06u l=150000u
X1395 a_301_3864# en29_b a_2454_3868# VPWR sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.36e+06u l=150000u
X1396 a_2454_29608# en9_b a_301_29604# VPWR sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.36e+06u l=150000u
X1397 a_2454_6442# a_2450_6354# out VGND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X1398 a_301_1290# en31_b a_2454_1294# VPWR sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.36e+06u l=150000u
X1399 a_301_29604# en in_9 VGND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X1400 a_2454_34756# en5_b a_301_34752# VPWR sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.36e+06u l=150000u
X1401 a_301_5151# en_b in_28 VPWR sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.36e+06u l=150000u
X1402 VPWR en25_b a_2450_8928# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.6e+11p ps=2.52e+06u w=1e+06u l=150000u
X1403 a_301_11586# a_2450_11502# a_2454_11590# VGND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X1404 out a_2450_20511# a_2454_20599# VGND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X1405 a_2454_30895# a_2450_30807# out VGND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X1406 in_27 en a_301_6438# VGND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X1407 out a_2450_15363# a_2454_15451# VGND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X1408 a_2454_10303# en24_b out VPWR sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.36e+06u l=150000u
X1409 in_24 en a_301_10299# VGND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X1410 a_301_9012# en25_b a_2454_9016# VPWR sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.36e+06u l=150000u
X1411 a_301_20595# en in_16 VGND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X1412 a_2454_34756# a_2450_34668# a_301_34752# VGND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X1413 a_301_19308# a_2450_19224# a_2454_19312# VGND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X1414 in_24 en_b a_301_10299# VPWR sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.36e+06u l=150000u
X1415 out a_2450_35955# a_2454_36043# VGND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X1416 out en6_b a_2454_33469# VPWR sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.36e+06u l=150000u
X1417 out en0_b a_2454_41191# VPWR sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.36e+06u l=150000u
X1418 out en21_b a_2454_14164# VPWR sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.36e+06u l=150000u
X1419 a_2454_27034# a_2450_26946# out VGND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X1420 in_25 en a_301_9012# VGND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X1421 in_20 en_b a_301_15447# VPWR sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.36e+06u l=150000u
X1422 a_301_20595# en16_b a_2454_20599# VPWR sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.36e+06u l=150000u
X1423 a_2454_24460# en13_b out VPWR sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.36e+06u l=150000u
X1424 a_301_41187# en in_0 VGND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X1425 a_301_32178# en_b in_7 VPWR sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.36e+06u l=150000u
X1426 out a_2450_17937# a_2454_18025# VGND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X1427 a_301_39900# en_b in_1 VPWR sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.36e+06u l=150000u
X1428 in_14 en_b a_301_23169# VPWR sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.36e+06u l=150000u
X1429 in_8 en_b a_301_30891# VPWR sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.36e+06u l=150000u
X1430 a_301_25743# en12_b a_2454_25747# VPWR sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.36e+06u l=150000u
X1431 a_2454_36043# en4_b a_301_36039# VPWR sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.36e+06u l=150000u
X1432 a_2454_5155# en28_b out VPWR sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.36e+06u l=150000u
X1433 VPWR en8_b a_2450_30807# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.6e+11p ps=2.52e+06u w=1e+06u l=150000u
X1434 in_20 en a_301_15447# VGND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X1435 a_2454_10303# a_2450_10215# a_301_10299# VGND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X1436 a_2454_7729# en26_b out VPWR sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.36e+06u l=150000u
X1437 a_2454_7729# a_2450_7641# a_301_7725# VGND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X1438 a_301_18021# en_b in_18 VPWR sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.36e+06u l=150000u
X1439 a_301_25743# a_2450_25659# a_2454_25747# VGND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X1440 out a_2450_8928# a_2454_9016# VGND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X1441 a_2454_10303# en24_b a_301_10299# VPWR sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.36e+06u l=150000u
X1442 a_2454_3868# en29_b a_301_3864# VPWR sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.36e+06u l=150000u
X1443 out en23_b a_2454_11590# VPWR sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.36e+06u l=150000u
X1444 a_2454_38617# en2_b VGND VGND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X1445 a_301_32178# en7_b a_2454_32182# VPWR sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.36e+06u l=150000u
X1446 a_301_39900# en1_b a_2454_39904# VPWR sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.36e+06u l=150000u
X1447 a_301_12873# en22_b a_2454_12877# VPWR sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.36e+06u l=150000u
X1448 a_301_5151# en28_b a_2454_5155# VPWR sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.36e+06u l=150000u
X1449 a_2454_23173# en14_b a_301_23169# VPWR sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.36e+06u l=150000u
X1450 a_301_33465# en6_b a_2454_33469# VPWR sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.36e+06u l=150000u
X1451 a_2454_30895# en8_b a_301_30891# VPWR sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.36e+06u l=150000u
X1452 a_301_41187# en0_b a_2454_41191# VPWR sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.36e+06u l=150000u
X1453 a_2454_7729# a_2450_7641# out VGND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X1454 VPWR en28_b a_2450_5067# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.6e+11p ps=2.52e+06u w=1e+06u l=150000u
X1455 a_301_5151# a_2450_5067# a_2454_5155# VGND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X1456 a_301_1290# en_b in_31 VPWR sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.36e+06u l=150000u
X1457 in_29 en_b a_301_3864# VPWR sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.36e+06u l=150000u
X1458 a_301_12873# a_2450_12789# a_2454_12877# VGND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X1459 out a_2450_16650# a_2454_16738# VGND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X1460 a_2454_14164# a_2450_14076# out VGND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X1461 out a_2450_24372# a_2454_24460# VGND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X1462 a_2454_20599# a_2450_20511# out VGND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X1463 VGND en11_b a_2450_26946# VGND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.69e+11p ps=1.82e+06u w=650000u l=150000u
X1464 out a_2450_30807# a_2454_30895# VGND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X1465 a_2454_9016# a_2450_8928# a_301_9012# VGND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X1466 a_301_9012# en_b in_25 VPWR sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.36e+06u l=150000u
X1467 a_2454_15451# a_2450_15363# out VGND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X1468 in_29 en a_301_3864# VGND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X1469 out en24_b a_2454_10303# VPWR sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.36e+06u l=150000u
X1470 in_21 en a_301_14160# VGND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X1471 a_301_28317# a_2450_28233# a_2454_28321# VGND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X1472 a_301_33465# en6_b a_2454_33469# VPWR sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.36e+06u l=150000u
X1473 a_2454_19312# en17_b out VPWR sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.36e+06u l=150000u
X1474 a_301_41187# en0_b a_2454_41191# VPWR sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.36e+06u l=150000u
X1475 a_301_14160# en21_b a_2454_14164# VPWR sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.36e+06u l=150000u
X1476 a_2454_24460# en13_b a_301_24456# VPWR sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.36e+06u l=150000u
X1477 a_2454_36043# a_2450_35955# out VGND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X1478 a_301_33465# en_b in_6 VPWR sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.36e+06u l=150000u
X1479 a_2454_1294# en31_b out VPWR sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.36e+06u l=150000u
X1480 a_301_37326# en in_3 VGND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X1481 in_13 en_b a_301_24456# VPWR sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.36e+06u l=150000u
X1482 in_17 en_b a_301_19308# VPWR sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.36e+06u l=150000u
X1483 in_7 en_b a_301_32178# VPWR sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.36e+06u l=150000u
X1484 in_1 en_b a_301_39900# VPWR sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.36e+06u l=150000u
X1485 a_301_33465# en in_6 VGND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X1486 a_2454_33469# en6_b a_301_33465# VPWR sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.36e+06u l=150000u
X1487 a_2454_41191# en0_b a_301_41187# VPWR sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.36e+06u l=150000u
X1488 a_2454_2581# en30_b out VPWR sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.36e+06u l=150000u
X1489 out a_2450_2493# a_2454_2581# VGND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X1490 a_2454_9016# en25_b out VPWR sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.36e+06u l=150000u
X1491 a_301_1290# a_2450_1206# a_2454_1294# VGND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X1492 a_2454_19312# a_2450_19224# a_301_19308# VGND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X1493 in_1 en a_301_39900# VGND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X1494 a_301_6438# en27_b a_2454_6442# VPWR sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.36e+06u l=150000u
X1495 a_2454_14164# a_2450_14076# a_301_14160# VGND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X1496 a_2454_5155# en28_b a_301_5151# VPWR sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.36e+06u l=150000u
X1497 a_301_1290# en31_b a_2454_1294# VPWR sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.36e+06u l=150000u
X1498 a_2454_29608# en9_b out VPWR sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.36e+06u l=150000u
X1499 out en16_b a_2454_20599# VPWR sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.36e+06u l=150000u
X1500 a_2454_11590# en23_b out VPWR sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.36e+06u l=150000u
X1501 a_2454_34756# en5_b out VPWR sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.36e+06u l=150000u
X1502 a_2454_19312# en17_b a_301_19308# VPWR sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.36e+06u l=150000u
X1503 a_301_5151# en in_28 VGND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X1504 a_301_16734# en19_b a_2454_16738# VPWR sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.36e+06u l=150000u
X1505 out en12_b a_2454_25747# VPWR sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.36e+06u l=150000u
X1506 a_2454_36043# en4_b out VPWR sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.36e+06u l=150000u
X1507 in_5 en_b a_301_34752# VPWR sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.36e+06u l=150000u
X1508 a_301_25743# en_b in_12 VPWR sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.36e+06u l=150000u
X1509 a_2454_10303# a_2450_10215# out VGND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X1510 VGND en20_b a_2450_15363# VGND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.69e+11p ps=1.82e+06u w=650000u l=150000u
X1511 a_301_9012# a_2450_8928# a_2454_9016# VGND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X1512 a_2454_34756# a_2450_34668# out VGND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X1513 a_301_21882# en_b in_15 VPWR sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.36e+06u l=150000u
X1514 in_7 en_b a_301_32178# VPWR sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.36e+06u l=150000u
X1515 a_2454_20599# a_2450_20511# a_301_20595# VGND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X1516 out a_2450_25659# a_2454_25747# VGND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X1517 a_301_29604# en_b in_9 VPWR sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.36e+06u l=150000u
X1518 in_1 en_b a_301_39900# VPWR sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.36e+06u l=150000u
X1519 a_2454_16738# a_2450_16650# out VGND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X1520 in_5 en a_301_34752# VGND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X1521 a_301_10299# en24_b a_2454_10303# VPWR sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.36e+06u l=150000u
X1522 out a_2450_14076# a_2454_14164# VGND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X1523 in_20 en a_301_15447# VGND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X1524 a_2454_24460# a_2450_24372# out VGND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X1525 a_2454_39904# a_2450_39816# a_301_39900# VGND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X1526 a_301_25743# en in_12 VGND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X1527 a_301_29604# a_2450_29520# a_2454_29608# VGND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X1528 a_2454_32182# en7_b a_301_32178# VPWR sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.36e+06u l=150000u
X1529 a_2454_39904# en1_b a_301_39900# VPWR sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.36e+06u l=150000u
X1530 a_2454_36043# a_2450_35955# a_301_36039# VGND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X1531 a_2454_5155# a_2450_5067# out VGND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X1532 out en17_b a_2454_19312# VPWR sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.36e+06u l=150000u
X1533 in_4 en a_301_36039# VGND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X1534 a_301_21882# en in_15 VGND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X1535 in_6 en_b a_301_33465# VPWR sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.36e+06u l=150000u
X1536 VPWR en10_b a_2450_28233# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.6e+11p ps=2.52e+06u w=1e+06u l=150000u
X1537 VPWR en4_b a_2450_35955# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.6e+11p ps=2.52e+06u w=1e+06u l=150000u
X1538 a_2454_1294# a_2450_1206# a_301_1290# VGND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X1539 a_301_18021# en in_18 VGND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X1540 out a_2450_3780# a_2454_3868# VGND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X1541 a_2454_6442# en27_b a_301_6438# VPWR sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.36e+06u l=150000u
X1542 a_2454_10303# a_2450_10215# a_301_10299# VGND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X1543 a_2454_1294# en31_b a_301_1290# VPWR sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.36e+06u l=150000u
X1544 a_2454_5155# en28_b VGND VGND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X1545 a_301_32178# a_2450_32094# a_2454_32182# VGND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X1546 a_301_5151# a_2450_5067# a_2454_5155# VGND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X1547 a_2454_23173# a_2450_23085# a_301_23169# VGND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X1548 a_2454_23173# en14_b out VPWR sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.36e+06u l=150000u
X1549 out en6_b a_2454_33469# VPWR sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.36e+06u l=150000u
X1550 a_2454_30895# en8_b out VPWR sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.36e+06u l=150000u
X1551 out en0_b a_2454_41191# VPWR sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.36e+06u l=150000u
X1552 out en21_b a_2454_14164# VPWR sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.36e+06u l=150000u
X1553 a_2454_24460# en13_b out VPWR sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.36e+06u l=150000u
X1554 out en9_b a_2454_29608# VPWR sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.36e+06u l=150000u
X1555 a_301_37326# en3_b a_2454_37330# VPWR sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.36e+06u l=150000u
X1556 in_14 en_b a_301_23169# VPWR sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.36e+06u l=150000u
X1557 a_301_6438# en in_27 VGND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X1558 a_301_14160# en_b in_21 VPWR sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.36e+06u l=150000u
X1559 a_301_18021# en18_b a_2454_18025# VPWR sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.36e+06u l=150000u
X1560 a_2454_20599# en16_b out VPWR sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.36e+06u l=150000u
X1561 in_8 en_b a_301_30891# VPWR sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.36e+06u l=150000u
X1562 a_2454_28321# en10_b a_301_28317# VPWR sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.36e+06u l=150000u
X1563 out en5_b a_2454_34756# VPWR sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.36e+06u l=150000u
X1564 VGND en23_b a_2450_11502# VGND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.69e+11p ps=1.82e+06u w=650000u l=150000u
X1565 a_2454_25747# en12_b out VPWR sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.36e+06u l=150000u
X1566 out en4_b a_2454_36043# VPWR sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.36e+06u l=150000u
X1567 in_25 en_b a_301_9012# VPWR sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.36e+06u l=150000u
X1568 a_301_34752# en_b in_5 VPWR sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.36e+06u l=150000u
X1569 VGND en19_b a_2450_16650# VGND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.69e+11p ps=1.82e+06u w=650000u l=150000u
X1570 a_301_9012# en in_25 VGND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X1571 out a_2450_10215# a_2454_10303# VGND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X1572 in_6 en_b a_301_33465# VPWR sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.36e+06u l=150000u
X1573 out a_2450_34668# a_2454_34756# VGND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X1574 a_2454_19312# a_2450_19224# out VGND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X1575 a_301_14160# a_2450_14076# a_2454_14164# VGND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X1576 a_2454_25747# a_2450_25659# out VGND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X1577 a_301_33465# en in_6 VGND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X1578 a_2454_24460# a_2450_24372# a_301_24456# VGND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X1579 in_13 en a_301_24456# VGND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X1580 a_301_34752# en in_5 VGND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X1581 a_301_38613# en_b in_2 VPWR sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.36e+06u l=150000u
X1582 a_2454_11590# en23_b VGND VGND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X1583 a_301_19308# en17_b a_2454_19312# VPWR sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.36e+06u l=150000u
X1584 VPWR en13_b a_2450_24372# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.6e+11p ps=2.52e+06u w=1e+06u l=150000u
X1585 out en26_b a_2454_7729# VPWR sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.36e+06u l=150000u
X1586 a_301_30891# en in_8 VGND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X1587 a_2454_27034# en11_b VGND VGND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X1588 VPWR en9_b a_2450_29520# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.6e+11p ps=2.52e+06u w=1e+06u l=150000u
X1589 a_2454_2581# a_2450_2493# out VGND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X1590 a_301_38613# en in_2 VGND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X1591 a_2454_9016# a_2450_8928# out VGND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X1592 a_301_19308# en in_17 VGND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X1593 a_301_29604# en9_b a_2454_29608# VPWR sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.36e+06u l=150000u
X1594 a_301_34752# en5_b a_2454_34756# VPWR sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.36e+06u l=150000u
X1595 a_301_6438# a_2450_6354# a_2454_6442# VGND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X1596 a_2454_1294# en31_b VGND VGND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X1597 a_2454_11590# a_2450_11502# a_301_11586# VGND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X1598 a_2454_5155# a_2450_5067# a_301_5151# VGND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X1599 a_2454_20599# a_2450_20511# out VGND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X1600 out en24_b a_2454_10303# VPWR sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.36e+06u l=150000u
X1601 a_301_33465# a_2450_33381# a_2454_33469# VGND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X1602 a_301_10299# en in_24 VGND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X1603 a_301_41187# a_2450_41103# a_2454_41191# VGND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X1604 a_301_34752# a_2450_34668# a_2454_34756# VGND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X1605 a_2454_19312# a_2450_19224# a_301_19308# VGND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X1606 a_2454_32182# en7_b out VPWR sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.36e+06u l=150000u
X1607 a_301_3864# en_b in_29 VPWR sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.36e+06u l=150000u
X1608 a_301_10299# en_b in_24 VPWR sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.36e+06u l=150000u
X1609 a_2454_39904# en1_b out VPWR sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.36e+06u l=150000u
X1610 a_2454_36043# a_2450_35955# out VGND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X1611 out en14_b a_2454_23173# VPWR sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.36e+06u l=150000u
X1612 a_2454_33469# en6_b out VPWR sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.36e+06u l=150000u
X1613 in_13 en_b a_301_24456# VPWR sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.36e+06u l=150000u
X1614 a_301_29604# en9_b a_2454_29608# VPWR sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.36e+06u l=150000u
X1615 out en8_b a_2454_30895# VPWR sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.36e+06u l=150000u
X1616 a_2454_41191# en0_b out VPWR sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.36e+06u l=150000u
X1617 a_2454_14164# en21_b out VPWR sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.36e+06u l=150000u
X1618 a_301_15447# en_b in_20 VPWR sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.36e+06u l=150000u
X1619 a_2454_20599# en16_b a_301_20595# VPWR sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.36e+06u l=150000u
X1620 a_301_21882# en_b in_15 VPWR sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.36e+06u l=150000u
X1621 out en13_b a_2454_24460# VPWR sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.36e+06u l=150000u
X1622 in_7 en_b a_301_32178# VPWR sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.36e+06u l=150000u
X1623 a_301_29604# en_b in_9 VPWR sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.36e+06u l=150000u
X1624 in_1 en_b a_301_39900# VPWR sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.36e+06u l=150000u
X1625 in_22 en_b a_301_12873# VPWR sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.36e+06u l=150000u
X1626 a_301_23169# en_b in_14 VPWR sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.36e+06u l=150000u
X1627 a_301_34752# en5_b a_2454_34756# VPWR sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.36e+06u l=150000u
X1628 in_16 en_b a_301_20595# VPWR sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.36e+06u l=150000u
X1629 a_301_30891# en_b in_8 VPWR sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.36e+06u l=150000u
X1630 a_2454_25747# en12_b a_301_25743# VPWR sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.36e+06u l=150000u
X1631 a_301_3864# en in_29 VGND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X1632 a_301_11586# en_b in_23 VPWR sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.36e+06u l=150000u
X1633 in_30 en_b a_301_2577# VPWR sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.36e+06u l=150000u
X1634 a_2454_3868# en29_b out VPWR sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.36e+06u l=150000u
X1635 a_301_10299# a_2450_10215# a_2454_10303# VGND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X1636 a_301_21882# en in_15 VGND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X1637 a_2454_29608# en9_b a_301_29604# VPWR sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.36e+06u l=150000u
X1638 in_22 en a_301_12873# VGND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X1639 a_2454_39904# a_2450_39816# out VGND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X1640 a_301_34752# a_2450_34668# a_2454_34756# VGND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X1641 a_301_27030# en_b in_11 VPWR sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.36e+06u l=150000u
X1642 a_2454_34756# en5_b a_301_34752# VPWR sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.36e+06u l=150000u
X1643 a_2454_25747# a_2450_25659# a_301_25743# VGND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X1644 a_2454_32182# a_2450_32094# a_301_32178# VGND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X1645 in_1 en a_301_39900# VGND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X1646 out a_2450_19224# a_2454_19312# VGND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X1647 in_6 en a_301_33465# VGND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X1648 out en30_b a_2454_2581# VPWR sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.36e+06u l=150000u
X1649 a_2454_37330# en3_b a_301_37326# VPWR sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.36e+06u l=150000u
X1650 out en25_b a_2454_9016# VPWR sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.36e+06u l=150000u
X1651 a_2454_34756# a_2450_34668# a_301_34752# VGND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X1652 a_2454_1294# a_2450_1206# a_301_1290# VGND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X1653 a_2454_3868# a_2450_3780# out VGND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X1654 a_2454_28321# en10_b VGND VGND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X1655 a_301_21882# en15_b a_2454_21886# VPWR sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.36e+06u l=150000u
X1656 a_2454_32182# en7_b a_301_32178# VPWR sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.36e+06u l=150000u
X1657 a_2454_39904# en1_b a_301_39900# VPWR sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.36e+06u l=150000u
X1658 a_2454_12877# en22_b a_301_12873# VPWR sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.36e+06u l=150000u
X1659 a_301_23169# en14_b a_2454_23173# VPWR sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.36e+06u l=150000u
X1660 a_301_30891# en8_b a_2454_30895# VPWR sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.36e+06u l=150000u
X1661 a_2454_6442# en27_b a_301_6438# VPWR sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.36e+06u l=150000u
X1662 a_2454_6442# a_2450_6354# a_301_6438# VGND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X1663 a_301_21882# a_2450_21798# a_2454_21886# VGND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X1664 a_301_7725# a_2450_7641# a_2454_7729# VGND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X1665 a_2454_12877# a_2450_12789# a_301_12873# VGND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X1666 a_2454_23173# a_2450_23085# out VGND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X1667 out a_2450_14076# a_2454_14164# VGND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X1668 out a_2450_20511# a_2454_20599# VGND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X1669 a_2454_24460# a_2450_24372# out VGND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X1670 a_301_37326# a_2450_37242# a_2454_37330# VGND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X1671 a_2454_10303# en24_b out VPWR sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.36e+06u l=150000u
X1672 a_301_14160# en in_21 VGND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X1673 a_301_18021# a_2450_17937# a_2454_18025# VGND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X1674 a_2454_28321# a_2450_28233# a_301_28317# VGND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X1675 a_2454_28321# en10_b out VPWR sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.36e+06u l=150000u
X1676 a_301_23169# en14_b a_2454_23173# VPWR sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.36e+06u l=150000u
X1677 out en17_b a_2454_19312# VPWR sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.36e+06u l=150000u
X1678 a_301_30891# en8_b a_2454_30895# VPWR sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.36e+06u l=150000u
X1679 in_4 en a_301_36039# VGND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X1680 out en7_b a_2454_32182# VPWR sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.36e+06u l=150000u
X1681 a_2454_14164# en21_b a_301_14160# VPWR sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.36e+06u l=150000u
X1682 out en1_b a_2454_39904# VPWR sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.36e+06u l=150000u
X1683 in_6 en_b a_301_33465# VPWR sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.36e+06u l=150000u
X1684 out a_2450_35955# a_2454_36043# VGND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X1685 a_301_24456# en_b in_13 VPWR sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.36e+06u l=150000u
X1686 in_31 en a_301_1290# VGND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X1687 in_25 en a_301_9012# VGND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X1688 a_301_19308# en_b in_17 VPWR sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.36e+06u l=150000u
X1689 in_15 en_b a_301_21882# VPWR sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.36e+06u l=150000u
X1690 in_9 en_b a_301_29604# VPWR sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.36e+06u l=150000u
X1691 a_301_23169# en in_14 VGND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X1692 a_301_38613# en_b in_2 VPWR sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.36e+06u l=150000u
X1693 in_6 en a_301_33465# VGND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X1694 in_27 en_b a_301_6438# VPWR sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.36e+06u l=150000u
X1695 a_2454_5155# en28_b out VPWR sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.36e+06u l=150000u
X1696 a_2454_23173# en14_b a_301_23169# VPWR sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.36e+06u l=150000u
X1697 a_2454_30895# en8_b a_301_30891# VPWR sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.36e+06u l=150000u
X1698 in_15 en a_301_21882# VGND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X1699 a_301_28317# en_b in_10 VPWR sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.36e+06u l=150000u
X1700 a_2454_33469# a_2450_33381# a_301_33465# VGND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X1701 a_301_36039# en_b in_4 VPWR sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.36e+06u l=150000u
X1702 out a_2450_39816# a_2454_39904# VGND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X1703 a_301_19308# a_2450_19224# a_2454_19312# VGND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X1704 a_301_38613# en in_2 VGND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X1705 a_2454_7729# en26_b out VPWR sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.36e+06u l=150000u
X1706 in_9 en a_301_29604# VGND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X1707 a_301_39900# en in_1 VGND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X1708 a_301_1290# a_2450_1206# a_2454_1294# VGND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X1709 a_2454_16738# en19_b VGND VGND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X1710 out a_2450_1206# a_2454_1294# VGND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X1711 out en9_b a_2454_29608# VPWR sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.36e+06u l=150000u
X1712 a_301_6438# en27_b a_2454_6442# VPWR sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.36e+06u l=150000u
X1713 a_2454_20599# en16_b out VPWR sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.36e+06u l=150000u
X1714 out en27_b a_2454_6442# VPWR sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.36e+06u l=150000u
X1715 out en5_b a_2454_34756# VPWR sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.36e+06u l=150000u
X1716 a_2454_16738# en19_b a_301_16734# VPWR sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.36e+06u l=150000u
X1717 a_2454_25747# en12_b out VPWR sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.36e+06u l=150000u
X1718 a_2454_7729# a_2450_7641# a_301_7725# VGND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X1719 a_301_38613# en2_b a_2454_38617# VPWR sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.36e+06u l=150000u
X1720 a_2454_11590# a_2450_11502# out VGND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X1721 out a_2450_10215# a_2454_10303# VGND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X1722 a_301_30891# a_2450_30807# a_2454_30895# VGND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X1723 out a_2450_34668# a_2454_34756# VGND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X1724 in_15 en_b a_301_21882# VPWR sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.36e+06u l=150000u
X1725 a_2454_25747# a_2450_25659# out VGND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X1726 a_2454_32182# a_2450_32094# out VGND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X1727 in_9 en_b a_301_29604# VPWR sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.36e+06u l=150000u
X1728 out a_2450_23085# a_2454_23173# VGND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X1729 a_301_11586# en_b in_23 VPWR sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.36e+06u l=150000u
X1730 in_13 en a_301_24456# VGND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X1731 a_301_38613# a_2450_38529# a_2454_38617# VGND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X1732 a_2454_10303# en24_b a_301_10299# VPWR sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.36e+06u l=150000u
X1733 a_2454_14164# a_2450_14076# out VGND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X1734 out a_2450_24372# a_2454_24460# VGND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X1735 a_301_15447# en in_20 VGND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X1736 a_2454_29608# a_2450_29520# a_301_29604# VGND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X1737 a_301_39900# a_2450_39816# a_2454_39904# VGND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X1738 a_2454_37330# en3_b out VPWR sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.36e+06u l=150000u
X1739 a_301_9012# en_b in_25 VPWR sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.36e+06u l=150000u
X1740 a_2454_21886# en15_b a_301_21882# VPWR sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.36e+06u l=150000u
X1741 a_301_32178# en7_b a_2454_32182# VPWR sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.36e+06u l=150000u
X1742 a_301_39900# en1_b a_2454_39904# VPWR sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.36e+06u l=150000u
X1743 a_301_2577# en_b in_30 VPWR sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.36e+06u l=150000u
X1744 out en10_b a_2454_28321# VPWR sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.36e+06u l=150000u
X1745 a_301_11586# en in_23 VGND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X1746 a_2454_19312# en17_b out VPWR sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.36e+06u l=150000u
X1747 in_15 en a_301_21882# VGND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X1748 a_301_36039# en in_4 VGND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X1749 in_30 en a_301_2577# VGND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X1750 a_301_27030# en_b in_11 VPWR sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.36e+06u l=150000u
X1751 in_18 en_b a_301_18021# VPWR sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.36e+06u l=150000u
X1752 a_2454_1294# en31_b out VPWR sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.36e+06u l=150000u
X1753 VPWR en18_b a_2450_17937# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.6e+11p ps=2.52e+06u w=1e+06u l=150000u
X1754 VPWR en12_b a_2450_25659# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.6e+11p ps=2.52e+06u w=1e+06u l=150000u
X1755 a_301_32178# en in_7 VGND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X1756 a_2454_21886# a_2450_21798# a_301_21882# VGND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X1757 a_301_27030# en in_11 VGND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X1758 in_2 en_b a_301_38613# VPWR sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.36e+06u l=150000u
X1759 VGND en29_b a_2450_3780# VGND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.69e+11p ps=1.82e+06u w=650000u l=150000u
X1760 a_301_37326# en_b in_3 VPWR sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.36e+06u l=150000u
X1761 a_301_39900# a_2450_39816# a_2454_39904# VGND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X1762 out a_2450_2493# a_2454_2581# VGND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X1763 a_2454_37330# a_2450_37242# a_301_37326# VGND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X1764 out a_2450_8928# a_2454_9016# VGND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X1765 a_2454_9016# en25_b out VPWR sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.36e+06u l=150000u
X1766 in_2 en a_301_38613# VGND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X1767 a_2454_32182# a_2450_32094# a_301_32178# VGND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X1768 a_2454_12877# en22_b out VPWR sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.36e+06u l=150000u
X1769 a_301_23169# a_2450_23085# a_2454_23173# VGND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X1770 out en14_b a_2454_23173# VPWR sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.36e+06u l=150000u
X1771 out en8_b a_2454_30895# VPWR sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.36e+06u l=150000u
X1772 a_2454_14164# en21_b out VPWR sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.36e+06u l=150000u
X1773 a_2454_39904# a_2450_39816# a_301_39900# VGND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X1774 a_2454_6442# a_2450_6354# a_301_6438# VGND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X1775 in_22 en_b a_301_12873# VPWR sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.36e+06u l=150000u
X1776 a_301_27030# en11_b a_2454_27034# VPWR sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.36e+06u l=150000u
X1777 a_2454_29608# en9_b out VPWR sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.36e+06u l=150000u
X1778 a_2454_37330# en3_b a_301_37326# VPWR sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.36e+06u l=150000u
X1779 in_16 en_b a_301_20595# VPWR sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.36e+06u l=150000u
X1780 a_2454_18025# en18_b a_301_18021# VPWR sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.36e+06u l=150000u
X1781 out en16_b a_2454_20599# VPWR sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.36e+06u l=150000u
X1782 a_301_28317# en10_b a_2454_28321# VPWR sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.36e+06u l=150000u
X1783 a_2454_34756# en5_b out VPWR sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.36e+06u l=150000u
X1784 a_2454_12877# a_2450_12789# out VGND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X1785 out en12_b a_2454_25747# VPWR sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.36e+06u l=150000u
X1786 in_29 en_b a_301_3864# VPWR sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.36e+06u l=150000u
X1787 out a_2450_11502# a_2454_11590# VGND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X1788 VGND en6_b a_2450_33381# VGND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.69e+11p ps=1.82e+06u w=650000u l=150000u
X1789 VGND en0_b a_2450_41103# VGND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.69e+11p ps=1.82e+06u w=650000u l=150000u
X1790 in_22 en a_301_12873# VGND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X1791 a_2454_10303# a_2450_10215# out VGND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X1792 a_2454_33469# a_2450_33381# out VGND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X1793 a_2454_28321# a_2450_28233# out VGND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X1794 a_2454_34756# a_2450_34668# out VGND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X1795 a_2454_2581# en30_b a_301_2577# VPWR sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.36e+06u l=150000u
X1796 a_301_23169# a_2450_23085# a_2454_23173# VGND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X1797 out a_2450_19224# a_2454_19312# VGND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X1798 a_2454_14164# a_2450_14076# a_301_14160# VGND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X1799 a_301_23169# en in_14 VGND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X1800 out a_2450_25659# a_2454_25747# VGND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X1801 out a_2450_32094# a_2454_32182# VGND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X1802 in_6 en a_301_33465# VGND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X1803 in_29 en a_301_3864# VGND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X1804 a_301_1290# en in_31 VGND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X1805 in_23 en_b a_301_11586# VPWR sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.36e+06u l=150000u
X1806 a_301_24456# en in_13 VGND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X1807 in_2 en_b a_301_38613# VPWR sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.36e+06u l=150000u
X1808 out en29_b a_2454_3868# VPWR sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.36e+06u l=150000u
X1809 a_301_28317# en10_b a_2454_28321# VPWR sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.36e+06u l=150000u
X1810 out en3_b a_2454_37330# VPWR sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.36e+06u l=150000u
X1811 VPWR en21_b a_2450_14076# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.6e+11p ps=2.52e+06u w=1e+06u l=150000u
X1812 a_2454_19312# en17_b a_301_19308# VPWR sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.36e+06u l=150000u
X1813 a_301_6438# en_b in_27 VPWR sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.36e+06u l=150000u
X1814 a_301_28317# en_b in_10 VPWR sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.36e+06u l=150000u
X1815 a_301_20595# en in_16 VGND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X1816 a_2454_41191# en0_b VGND VGND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X1817 a_2454_5155# a_2450_5067# out VGND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X1818 a_2454_23173# a_2450_23085# a_301_23169# VGND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X1819 a_2454_38617# en2_b a_301_38613# VPWR sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.36e+06u l=150000u
X1820 in_11 en_b a_301_27030# VPWR sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.36e+06u l=150000u
X1821 a_301_28317# en in_10 VGND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X1822 in_2 en a_301_38613# VGND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X1823 a_2454_2581# en30_b out VPWR sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.36e+06u l=150000u
X1824 a_2454_28321# en10_b a_301_28317# VPWR sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.36e+06u l=150000u
X1825 VGND en26_b a_2450_7641# VGND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.69e+11p ps=1.82e+06u w=650000u l=150000u
X1826 out a_2450_3780# a_2454_3868# VGND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X1827 a_2454_38617# a_2450_38529# a_301_38613# VGND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X1828 a_301_11586# a_2450_11502# a_2454_11590# VGND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X1829 in_30 en_b a_301_2577# VPWR sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.36e+06u l=150000u
X1830 a_2454_10303# en24_b out VPWR sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.36e+06u l=150000u
X1831 a_2454_33469# a_2450_33381# a_301_33465# VGND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X1832 a_301_6438# a_2450_6354# a_2454_6442# VGND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X1833 a_2454_3868# en29_b a_301_3864# VPWR sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.36e+06u l=150000u
X1834 a_301_15447# en20_b a_2454_15451# VPWR sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.36e+06u l=150000u
X1835 a_2454_41191# a_2450_41103# a_301_41187# VGND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X1836 out a_2450_6354# a_2454_6442# VGND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X1837 a_2454_21886# en15_b out VPWR sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.36e+06u l=150000u
X1838 out en7_b a_2454_32182# VPWR sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.36e+06u l=150000u
X1839 a_2454_16738# en19_b out VPWR sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.36e+06u l=150000u
X1840 out en1_b a_2454_39904# VPWR sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.36e+06u l=150000u
X1841 a_2454_7729# a_2450_7641# a_301_7725# VGND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X1842 out en22_b a_2454_12877# VPWR sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.36e+06u l=150000u
X1843 a_2454_23173# en14_b out VPWR sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.36e+06u l=150000u
X1844 in_28 en_b a_301_5151# VPWR sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.36e+06u l=150000u
X1845 a_2454_30895# en8_b out VPWR sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.36e+06u l=150000u
X1846 out en21_b a_2454_14164# VPWR sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.36e+06u l=150000u
X1847 a_301_36039# en4_b a_2454_36043# VPWR sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.36e+06u l=150000u
X1848 a_301_32178# en_b in_7 VPWR sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.36e+06u l=150000u
X1849 in_15 en_b a_301_21882# VPWR sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.36e+06u l=150000u
X1850 a_301_39900# en_b in_1 VPWR sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.36e+06u l=150000u
X1851 a_301_12873# en_b in_22 VPWR sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.36e+06u l=150000u
X1852 in_9 en_b a_301_29604# VPWR sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.36e+06u l=150000u
X1853 a_301_20595# en_b in_16 VPWR sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.36e+06u l=150000u
X1854 a_2454_21886# a_2450_21798# out VGND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X1855 in_23 en_b a_301_11586# VPWR sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.36e+06u l=150000u
X1856 a_301_11586# a_2450_11502# a_2454_11590# VGND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X1857 out a_2450_12789# a_2454_12877# VGND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X1858 VGND en5_b a_2450_34668# VGND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.69e+11p ps=1.82e+06u w=650000u l=150000u
X1859 a_2454_10303# a_2450_10215# a_301_10299# VGND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X1860 a_301_11586# en in_23 VGND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X1861 in_15 en a_301_21882# VGND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X1862 a_301_41187# en_b in_0 VPWR sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.36e+06u l=150000u
X1863 out a_2450_39816# a_2454_39904# VGND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X1864 a_301_12873# en in_22 VGND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X1865 a_2454_29608# a_2450_29520# out VGND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X1866 a_301_16734# en_b in_19 VPWR sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.36e+06u l=150000u
X1867 a_2454_37330# a_2450_37242# out VGND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X1868 a_301_9012# en in_25 VGND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X1869 in_11 en_b a_301_27030# VPWR sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.36e+06u l=150000u
X1870 out a_2450_33381# a_2454_33469# VGND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X1871 in_26 en_b a_301_7725# VPWR sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.36e+06u l=150000u
X1872 a_301_32178# a_2450_32094# a_2454_32182# VGND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X1873 a_301_2577# en in_30 VGND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X1874 out a_2450_28233# a_2454_28321# VGND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X1875 in_9 en a_301_29604# VGND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X1876 a_2454_19312# a_2450_19224# out VGND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X1877 a_301_27030# en in_11 VGND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X1878 in_14 en a_301_23169# VGND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X1879 out en28_b a_2454_5155# VPWR sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.36e+06u l=150000u
X1880 in_18 en a_301_18021# VGND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X1881 a_2454_11590# a_2450_11502# a_301_11586# VGND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X1882 a_2454_27034# en11_b a_301_27030# VPWR sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.36e+06u l=150000u
X1883 a_301_37326# en3_b a_2454_37330# VPWR sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.36e+06u l=150000u
X1884 a_301_16734# en in_19 VGND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X1885 in_26 en a_301_7725# VGND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X1886 in_10 en_b a_301_28317# VPWR sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.36e+06u l=150000u
X1887 a_2454_21886# en15_b a_301_21882# VPWR sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.36e+06u l=150000u
X1888 out en26_b a_2454_7729# VPWR sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.36e+06u l=150000u
X1889 a_301_12873# en22_b a_2454_12877# VPWR sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.36e+06u l=150000u
X1890 a_301_37326# en in_3 VGND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X1891 a_2454_9016# a_2450_8928# out VGND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X1892 in_31 en a_301_1290# VGND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X1893 a_2454_21886# a_2450_21798# a_301_21882# VGND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X1894 a_301_3864# en29_b a_2454_3868# VPWR sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.36e+06u l=150000u
X1895 a_301_12873# a_2450_12789# a_2454_12877# VGND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X1896 out a_2450_23085# a_2454_23173# VGND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X1897 a_2454_14164# a_2450_14076# out VGND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X1898 a_301_7725# a_2450_7641# a_2454_7729# VGND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X1899 in_27 en_b a_301_6438# VPWR sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.36e+06u l=150000u
X1900 a_2454_5155# en28_b a_301_5151# VPWR sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.36e+06u l=150000u
X1901 in_31 en_b a_301_1290# VPWR sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.36e+06u l=150000u
X1902 a_2454_37330# a_2450_37242# a_301_37326# VGND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X1903 out a_2450_7641# a_2454_7729# VGND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X1904 out en24_b a_2454_10303# VPWR sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.36e+06u l=150000u
X1905 a_301_27030# a_2450_26946# a_2454_27034# VGND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X1906 a_301_24456# en13_b a_2454_24460# VPWR sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.36e+06u l=150000u
X1907 a_2454_18025# a_2450_17937# a_301_18021# VGND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X1908 a_2454_18025# en18_b out VPWR sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.36e+06u l=150000u
X1909 a_301_28317# a_2450_28233# a_2454_28321# VGND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X1910 a_301_12873# en22_b a_2454_12877# VPWR sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.36e+06u l=150000u
X1911 out en10_b a_2454_28321# VPWR sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.36e+06u l=150000u
X1912 a_301_3864# en_b in_29 VPWR sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.36e+06u l=150000u
X1913 a_2454_19312# en17_b out VPWR sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.36e+06u l=150000u
X1914 out en15_b a_2454_21886# VPWR sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.36e+06u l=150000u
X1915 a_2454_32182# en7_b out VPWR sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.36e+06u l=150000u
X1916 out en19_b a_2454_16738# VPWR sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.36e+06u l=150000u
X1917 a_2454_39904# en1_b out VPWR sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.36e+06u l=150000u
X1918 a_301_33465# en_b in_6 VPWR sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.36e+06u l=150000u
X1919 in_18 en_b a_301_18021# VPWR sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.36e+06u l=150000u
X1920 a_2454_38617# en2_b out VPWR sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.36e+06u l=150000u
X1921 VGND en8_b a_2450_30807# VGND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.69e+11p ps=1.82e+06u w=650000u l=150000u
X1922 out a_2450_1206# a_2454_1294# VGND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X1923 a_301_12873# a_2450_12789# a_2454_12877# VGND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X1924 in_14 en a_301_23169# VGND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X1925 in_2 en_b a_301_38613# VPWR sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.36e+06u l=150000u
X1926 in_25 en_b a_301_9012# VPWR sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.36e+06u l=150000u
X1927 a_301_3864# en in_29 VGND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X1928 a_2454_2581# a_2450_2493# a_301_2577# VGND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X1929 a_2454_12877# en22_b a_301_12873# VPWR sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.36e+06u l=150000u
X1930 out a_2450_21798# a_2454_21886# VGND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X1931 out en27_b a_2454_6442# VPWR sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.36e+06u l=150000u
X1932 in_8 en a_301_30891# VGND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X1933 in_23 en a_301_11586# VGND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X1934 a_2454_38617# a_2450_38529# out VGND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X1935 in_10 en_b a_301_28317# VPWR sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.36e+06u l=150000u
X1936 a_301_33465# a_2450_33381# a_2454_33469# VGND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X1937 out en31_b a_2454_1294# VPWR sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.36e+06u l=150000u
X1938 a_301_25743# en_b in_12 VPWR sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.36e+06u l=150000u
X1939 a_2454_39904# a_2450_39816# out VGND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X1940 a_2454_15451# en20_b a_301_15447# VPWR sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.36e+06u l=150000u
X1941 a_301_28317# a_2450_28233# a_2454_28321# VGND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X1942 out a_2450_29520# a_2454_29608# VGND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X1943 out a_2450_37242# a_2454_37330# VGND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X1944 a_2454_19312# a_2450_19224# a_301_19308# VGND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X1945 a_301_28317# en in_10 VGND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X1946 in_2 en a_301_38613# VGND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X1947 in_17 en a_301_19308# VGND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X1948 a_2454_12877# a_2450_12789# a_301_12873# VGND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X1949 a_301_29604# en in_9 VGND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X1950 in_11 en a_301_27030# VGND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X1951 a_2454_2581# a_2450_2493# out VGND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X1952 a_301_25743# en in_12 VGND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X1953 a_2454_28321# a_2450_28233# a_301_28317# VGND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X1954 out en25_b a_2454_9016# VPWR sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.36e+06u l=150000u
X1955 a_301_16734# en19_b a_2454_16738# VPWR sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.36e+06u l=150000u
X1956 a_2454_38617# en2_b a_301_38613# VPWR sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.36e+06u l=150000u
X1957 in_30 en a_301_2577# VGND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X1958 out a_2450_11502# a_2454_11590# VGND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X1959 a_2454_10303# a_2450_10215# out VGND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X1960 a_301_5151# en28_b a_2454_5155# VPWR sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.36e+06u l=150000u
X1961 a_301_20595# a_2450_20511# a_2454_20599# VGND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X1962 a_2454_1294# en31_b a_301_1290# VPWR sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.36e+06u l=150000u
X1963 a_301_15447# a_2450_15363# a_2454_15451# VGND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X1964 a_2454_30895# a_2450_30807# a_301_30891# VGND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X1965 a_2454_41191# a_2450_41103# out VGND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X1966 out a_2450_32094# a_2454_32182# VGND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X1967 a_2454_23173# a_2450_23085# out VGND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X1968 a_2454_38617# a_2450_38529# a_301_38613# VGND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X1969 in_28 en a_301_5151# VGND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X1970 in_23 en_b a_301_11586# VPWR sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.36e+06u l=150000u
X1971 out a_2450_14076# a_2454_14164# VGND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X1972 a_301_36039# a_2450_35955# a_2454_36043# VGND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X1973 a_301_29604# a_2450_29520# a_2454_29608# VGND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X1974 a_2454_27034# en11_b out VPWR sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.36e+06u l=150000u
X1975 out en3_b a_2454_37330# VPWR sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.36e+06u l=150000u
X1976 a_301_21882# en15_b a_2454_21886# VPWR sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.36e+06u l=150000u
X1977 a_2454_32182# en7_b a_301_32178# VPWR sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.36e+06u l=150000u
X1978 a_301_16734# en19_b a_2454_16738# VPWR sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.36e+06u l=150000u
X1979 out en18_b a_2454_18025# VPWR sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.36e+06u l=150000u
X1980 a_301_41187# en_b in_0 VPWR sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.36e+06u l=150000u
X1981 a_2454_39904# en1_b a_301_39900# VPWR sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.36e+06u l=150000u
X1982 a_2454_28321# en10_b out VPWR sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.36e+06u l=150000u
X1983 in_23 en a_301_11586# VGND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X1984 out en17_b a_2454_19312# VPWR sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.36e+06u l=150000u
X1985 a_301_16734# en_b in_19 VPWR sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.36e+06u l=150000u
X1986 in_11 en_b a_301_27030# VPWR sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.36e+06u l=150000u
X1987 a_301_18021# en_b in_18 VPWR sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.36e+06u l=150000u
X1988 out en2_b a_2454_38617# VPWR sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.36e+06u l=150000u
X1989 a_301_41187# en in_0 VGND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X1990 a_301_7725# en_b in_26 VPWR sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.36e+06u l=150000u
X1991 a_2454_3868# en29_b out VPWR sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.36e+06u l=150000u
X1992 a_2454_3868# a_2450_3780# a_301_3864# VGND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X1993 a_301_21882# a_2450_21798# a_2454_21886# VGND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X1994 VGND en1_b a_2450_39816# VGND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.69e+11p ps=1.82e+06u w=650000u l=150000u
X1995 a_301_14160# en_b in_21 VPWR sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.36e+06u l=150000u
X1996 in_11 en a_301_27030# VGND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X1997 a_2454_16738# en19_b a_301_16734# VPWR sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.36e+06u l=150000u
X1998 a_301_16734# en in_19 VGND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X1999 out a_2450_5067# a_2454_5155# VGND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X2000 a_301_29604# a_2450_29520# a_2454_29608# VGND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X2001 a_2454_27034# a_2450_26946# a_301_27030# VGND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X2002 out a_2450_38529# a_2454_38617# VGND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X2003 a_301_37326# a_2450_37242# a_2454_37330# VGND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X2004 a_301_7725# en in_26 VGND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X2005 VGND en25_b a_2450_8928# VGND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.69e+11p ps=1.82e+06u w=650000u l=150000u
X2006 in_10 en a_301_28317# VGND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X2007 a_2454_34756# en5_b VGND VGND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X2008 a_301_1290# a_2450_1206# a_2454_1294# VGND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X2009 a_301_11586# en23_b a_2454_11590# VPWR sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.36e+06u l=150000u
X2010 out en22_b a_2454_12877# VPWR sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.36e+06u l=150000u
X2011 a_2454_3868# a_2450_3780# out VGND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X2012 VPWR en31_b a_2450_1206# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.6e+11p ps=2.52e+06u w=1e+06u l=150000u
X2013 a_2454_29608# a_2450_29520# a_301_29604# VGND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X2014 a_301_2577# en_b in_30 VPWR sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.36e+06u l=150000u
X2015 a_2454_27034# en11_b a_301_27030# VPWR sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.36e+06u l=150000u
C0 en2_b a_2450_39816# 0.49fF
C1 a_301_7725# a_2454_7729# 7.45fF
C2 a_301_34752# in_4 0.07fF
C3 en en17_b 0.01fF
C4 a_301_23169# en14_b 1.19fF
C5 a_2450_32094# a_301_33465# 0.01fF
C6 a_2450_23085# VPWR 0.55fF
C7 a_2450_5067# a_301_6438# 0.01fF
C8 en31_b a_2450_1206# 0.51fF
C9 a_301_20595# in_16 6.75fF
C10 a_2454_21886# a_2454_23173# 0.37fF
C11 in_17 VPWR 1.24fF
C12 out a_2454_10303# 7.60fF
C13 a_2450_6354# en26_b 0.01fF
C14 in_25 a_301_10299# 0.08fF
C15 a_301_9012# en 0.79fF
C16 en30_b en29_b 0.22fF
C17 a_301_23169# a_301_25743# 0.03fF
C18 a_301_2577# a_2450_3780# 0.05fF
C19 en27_b en26_b 0.22fF
C20 a_301_3864# in_30 0.08fF
C21 a_2450_28233# en 0.06fF
C22 in_29 in_31 0.03fF
C23 a_301_37326# VPWR 3.21fF
C24 a_301_11586# in_22 0.07fF
C25 en15_b en 0.01fF
C26 a_2450_7641# en_b 0.01fF
C27 a_301_1290# VPWR 2.94fF
C28 a_301_19308# in_18 0.08fF
C29 a_2454_21886# a_301_23169# 0.07fF
C30 out a_2450_35955# 0.78fF
C31 en5_b a_2450_35955# 0.49fF
C32 in_24 a_301_9012# 0.07fF
C33 en13_b out 0.70fF
C34 en21_b VPWR 3.16fF
C35 en20_b a_2450_15363# 0.51fF
C36 out a_301_3864# 0.43fF
C37 out a_301_5151# 0.43fF
C38 a_2450_30807# a_301_30891# 1.32fF
C39 a_2454_38617# VPWR 2.95fF
C40 in_12 a_301_27030# 0.08fF
C41 en19_b a_301_18021# 0.05fF
C42 in_14 a_301_21882# 0.07fF
C43 en6_b en 0.01fF
C44 a_2454_19312# VPWR 2.95fF
C45 en4_b en 0.01fF
C46 en28_b en 0.01fF
C47 en_b en19_b 0.05fF
C48 a_2454_36043# en4_b 1.80fF
C49 a_2450_26946# a_2450_25659# 0.18fF
C50 en a_301_7725# 0.79fF
C51 en13_b in_13 0.00fF
C52 en_b in_4 1.24fF
C53 en a_301_38613# 0.79fF
C54 en en29_b 0.01fF
C55 en in_20 1.38fF
C56 a_301_16734# a_2454_15451# 0.07fF
C57 en0_b a_2450_39816# 0.01fF
C58 a_2450_11502# a_301_12873# 0.01fF
C59 a_2454_30895# en9_b 0.10fF
C60 in_26 in_27 0.28fF
C61 a_2454_37330# a_2454_36043# 0.37fF
C62 in_14 en_b 1.24fF
C63 en9_b a_301_28317# 0.01fF
C64 out a_2450_1206# 0.70fF
C65 en9_b in_9 0.00fF
C66 a_2450_25659# a_2450_24372# 0.18fF
C67 en_b a_301_28317# 0.58fF
C68 a_2450_32094# en 0.06fF
C69 a_2450_17937# in_18 0.00fF
C70 in_9 en_b 1.24fF
C71 a_2454_21886# en14_b 0.03fF
C72 a_2454_34756# a_2454_33469# 0.37fF
C73 a_301_12873# en_b 0.58fF
C74 en30_b a_2454_2581# 1.80fF
C75 in_26 a_2454_7729# 0.05fF
C76 out a_2450_38529# 0.78fF
C77 a_301_6438# a_2454_6442# 7.45fF
C78 a_301_20595# a_2450_19224# 0.01fF
C79 a_301_27030# en10_b 0.01fF
C80 in_14 a_2450_23085# 0.00fF
C81 in_31 VPWR 1.16fF
C82 a_2454_10303# a_2450_8928# 0.03fF
C83 a_301_20595# a_301_19308# 0.39fF
C84 a_2454_34756# VPWR 2.95fF
C85 in_22 in_21 0.28fF
C86 en15_b in_15 0.00fF
C87 a_301_37326# in_4 0.08fF
C88 in_11 a_301_25743# 0.07fF
C89 a_2454_29608# a_2450_30807# 0.10fF
C90 a_2454_24460# a_301_24456# 7.45fF
C91 a_2450_16650# a_301_18021# 0.01fF
C92 in_19 en 1.38fF
C93 a_2450_29520# a_301_30891# 0.01fF
C94 a_2450_15363# VPWR 0.55fF
C95 a_301_29604# in_10 0.08fF
C96 a_2450_16650# en_b 0.01fF
C97 a_301_2577# a_2454_3868# 0.08fF
C98 out a_2450_3780# 0.78fF
C99 a_301_20595# a_301_23169# 0.03fF
C100 en13_b a_2454_25747# 0.10fF
C101 a_301_33465# a_2454_32182# 0.07fF
C102 a_2454_29608# en10_b 0.10fF
C103 a_2450_12789# a_301_14160# 0.01fF
C104 a_301_24456# VPWR 3.21fF
C105 out a_2450_6354# 0.78fF
C106 a_301_36039# a_2450_37242# 0.05fF
C107 a_2454_1294# a_301_1290# 7.45fF
C108 out en27_b 0.70fF
C109 a_2450_2493# a_301_3864# 0.01fF
C110 a_2454_5155# a_2454_7729# 0.03fF
C111 en7_b en6_b 0.22fF
C112 a_2450_12789# a_2450_14076# 0.18fF
C113 a_2450_28233# en11_b 0.49fF
C114 en_b a_2450_25659# 0.01fF
C115 a_301_12873# en21_b 0.01fF
C116 out a_2450_30807# 0.78fF
C117 a_2450_5067# a_2454_6442# 0.03fF
C118 in_26 en 1.38fF
C119 in_12 in_13 0.28fF
C120 a_301_29604# en 0.79fF
C121 a_2454_39904# a_301_38613# 0.08fF
C122 in_28 a_301_3864# 0.07fF
C123 in_28 a_301_5151# 6.75fF
C124 en8_b en 0.01fF
C125 a_2454_37330# a_2454_39904# 0.03fF
C126 en13_b a_2454_23173# 0.03fF
C127 in_1 en 1.38fF
C128 a_2454_16738# in_19 0.05fF
C129 a_2450_34668# in_5 0.00fF
C130 out a_2450_33381# 0.78fF
C131 a_301_11586# a_2450_11502# 1.32fF
C132 en2_b a_2450_38529# 0.51fF
C133 out en10_b 0.70fF
C134 en5_b a_2450_33381# 0.01fF
C135 en7_b a_2450_32094# 0.51fF
C136 a_2454_9016# a_2454_7729# 0.37fF
C137 in_24 in_26 0.03fF
C138 a_2450_2493# a_2450_1206# 0.18fF
C139 a_301_16734# en 0.79fF
C140 a_2450_29520# a_2454_29608# 1.92fF
C141 a_2454_27034# en10_b 0.03fF
C142 a_2450_26946# a_301_27030# 1.32fF
C143 in_10 in_8 0.03fF
C144 en12_b en 0.01fF
C145 en13_b a_301_23169# 0.01fF
C146 a_301_6438# a_301_5151# 0.39fF
C147 en16_b VPWR 3.16fF
C148 a_301_6438# a_301_3864# 0.03fF
C149 a_2454_18025# a_301_18021# 7.45fF
C150 in_3 en_b 1.24fF
C151 a_301_11586# en_b 0.58fF
C152 a_2454_15451# a_2454_12877# 0.03fF
C153 en23_b a_2454_12877# 0.10fF
C154 a_2450_15363# en19_b 0.01fF
C155 a_301_36039# in_5 0.08fF
C156 a_301_38613# a_301_41187# 0.03fF
C157 a_301_39900# a_301_38613# 0.39fF
C158 a_2450_11502# a_301_10299# 0.05fF
C159 a_2454_1294# in_31 0.05fF
C160 a_2450_10215# a_301_9012# 0.05fF
C161 en20_b in_20 0.00fF
C162 in_29 en29_b 0.00fF
C163 en25_b a_301_9012# 1.19fF
C164 a_301_20595# a_2454_21886# 0.08fF
C165 a_301_14160# a_301_15447# 0.39fF
C166 en17_b VPWR 3.16fF
C167 en18_b a_301_18021# 1.19fF
C168 in_8 en 1.38fF
C169 a_2450_29520# out 0.78fF
C170 en_b a_301_10299# 0.58fF
C171 in_12 a_2454_25747# 0.05fF
C172 a_2450_34668# a_301_36039# 0.01fF
C173 a_301_15447# a_2450_14076# 0.01fF
C174 a_2450_35955# a_2450_37242# 0.18fF
C175 in_14 a_301_24456# 0.08fF
C176 out a_2454_3868# 7.60fF
C177 in_0 in_2 0.03fF
C178 en18_b en_b 0.05fF
C179 a_2450_2493# a_2450_3780# 0.18fF
C180 a_301_9012# VPWR 3.21fF
C181 in_3 a_301_37326# 6.75fF
C182 en13_b en14_b 0.22fF
C183 in_25 a_2450_8928# 0.00fF
C184 en_b en26_b 0.05fF
C185 in_2 en_b 1.24fF
C186 a_301_16734# a_2454_16738# 7.45fF
C187 a_2454_9016# a_2454_11590# 0.03fF
C188 a_2450_28233# VPWR 0.55fF
C189 en6_b a_2454_33469# 1.80fF
C190 en15_b VPWR 3.16fF
C191 a_2450_5067# a_301_3864# 0.05fF
C192 a_2450_5067# a_301_5151# 1.32fF
C193 en3_b en 0.01fF
C194 en25_b a_301_7725# 0.01fF
C195 a_301_2577# en_b 0.58fF
C196 en9_b a_301_30891# 0.05fF
C197 a_301_30891# en_b 0.58fF
C198 a_2454_36043# en3_b 0.03fF
C199 en13_b a_301_25743# 0.05fF
C200 en7_b en8_b 0.22fF
C201 a_2450_16650# a_2450_15363# 0.18fF
C202 en6_b VPWR 3.16fF
C203 in_1 a_2454_39904# 0.05fF
C204 en6_b in_6 0.00fF
C205 out a_2450_26946# 0.78fF
C206 en4_b VPWR 3.16fF
C207 en_b in_21 1.24fF
C208 a_2454_18025# a_2454_19312# 0.37fF
C209 a_2450_32094# a_2454_33469# 0.03fF
C210 en28_b VPWR 3.16fF
C211 a_301_32178# a_2450_30807# 0.01fF
C212 a_2450_26946# a_2454_27034# 1.92fF
C213 a_301_7725# VPWR 3.21fF
C214 en_b a_301_27030# 0.58fF
C215 a_301_38613# VPWR 3.21fF
C216 a_2454_37330# VPWR 2.95fF
C217 en29_b VPWR 3.16fF
C218 en24_b a_2450_11502# 0.49fF
C219 in_2 a_301_37326# 0.07fF
C220 en a_2450_20511# 0.06fF
C221 a_301_6438# a_2450_6354# 1.32fF
C222 a_2450_38529# a_2450_37242# 0.18fF
C223 in_20 VPWR 1.24fF
C224 a_301_9012# a_2450_7641# 0.01fF
C225 out a_2450_24372# 0.78fF
C226 en31_b en_b 0.05fF
C227 en23_b a_2454_11590# 1.80fF
C228 a_301_6438# en27_b 1.19fF
C229 en23_b en 0.01fF
C230 a_2450_32094# VPWR 0.55fF
C231 out a_301_34752# 0.43fF
C232 en24_b en_b 0.05fF
C233 a_301_32178# a_2450_33381# 0.05fF
C234 en5_b a_301_34752# 1.19fF
C235 a_2454_15451# a_2454_14164# 0.37fF
C236 a_301_14160# a_2450_14076# 1.32fF
C237 en18_b a_2454_19312# 0.10fF
C238 in_1 a_301_41187# 0.08fF
C239 in_2 a_2454_38617# 0.05fF
C240 a_2454_12877# a_2454_11590# 0.37fF
C241 in_1 a_301_39900# 6.75fF
C242 en7_b a_2454_32182# 1.80fF
C243 a_301_2577# a_301_1290# 0.39fF
C244 a_301_24456# a_2450_25659# 0.05fF
C245 in_13 a_2450_24372# 0.00fF
C246 a_2450_34668# a_2450_35955# 0.18fF
C247 in_0 a_2454_41191# 0.05fF
C248 en12_b en11_b 0.22fF
C249 a_2454_12877# a_2454_14164# 0.37fF
C250 a_301_16734# en20_b 0.05fF
C251 a_2454_29608# en9_b 1.80fF
C252 in_27 en 1.38fF
C253 en1_b a_2454_41191# 0.10fF
C254 in_19 VPWR 1.24fF
C255 a_2450_7641# a_301_7725# 1.32fF
C256 a_301_33465# en 0.79fF
C257 a_2454_20599# VPWR 2.95fF
C258 a_2450_5067# a_2450_3780# 0.18fF
C259 en21_b in_21 0.00fF
C260 a_2450_2493# a_2454_3868# 0.03fF
C261 a_2450_35955# a_301_36039# 1.32fF
C262 a_2450_28233# a_301_28317# 1.32fF
C263 a_301_5151# a_2454_6442# 0.08fF
C264 out a_301_21882# 0.43fF
C265 en_b in_30 1.24fF
C266 en31_b a_301_1290# 1.17fF
C267 a_2450_5067# a_2450_6354# 0.18fF
C268 out a_2450_11502# 0.78fF
C269 a_2454_16738# a_2454_15451# 0.37fF
C270 a_2450_39816# a_2450_38529# 0.18fF
C271 in_12 a_301_25743# 6.75fF
C272 a_2454_2581# VPWR 2.95fF
C273 en4_b in_4 0.00fF
C274 out a_301_18021# 0.43fF
C275 a_2450_5067# en27_b 0.01fF
C276 out en9_b 0.70fF
C277 a_2450_26946# a_2454_25747# 0.10fF
C278 a_2450_21798# out 0.78fF
C279 en30_b en 0.01fF
C280 a_2450_12789# in_22 0.00fF
C281 in_16 a_301_21882# 0.08fF
C282 en5_b en_b 0.05fF
C283 in_10 en 1.38fF
C284 en1_b out 0.70fF
C285 a_301_2577# in_31 0.08fF
C286 in_11 in_12 0.28fF
C287 in_26 VPWR 1.24fF
C288 in_25 in_23 0.03fF
C289 a_2454_24460# en12_b 0.03fF
C290 a_301_29604# VPWR 3.21fF
C291 a_2454_25747# a_2450_24372# 0.03fF
C292 en8_b VPWR 3.16fF
C293 in_1 VPWR 1.24fF
C294 in_16 en_b 1.24fF
C295 out a_2450_23085# 0.78fF
C296 a_2454_41191# a_2454_38617# 0.03fF
C297 en_b in_13 1.24fF
C298 a_2450_32094# a_2454_30895# 0.10fF
C299 in_30 a_301_1290# 0.07fF
C300 a_301_16734# VPWR 3.21fF
C301 en22_b en23_b 0.22fF
C302 en12_b VPWR 3.16fF
C303 a_2450_41103# in_0 0.00fF
C304 en31_b in_31 0.00fF
C305 a_2454_32182# a_2454_33469# 0.37fF
C306 out a_301_37326# 0.43fF
C307 a_2450_41103# en_b 0.01fF
C308 in_19 en19_b 0.00fF
C309 a_2454_23173# a_2450_24372# 0.10fF
C310 a_2454_11590# a_2454_14164# 0.03fF
C311 a_2454_28321# en10_b 1.80fF
C312 en22_b a_2454_12877# 1.80fF
C313 a_2450_41103# en1_b 0.49fF
C314 out a_301_1290# 0.43fF
C315 in_16 in_17 0.28fF
C316 in_7 en_b 1.24fF
C317 in_23 in_22 0.28fF
C318 a_301_32178# a_301_34752# 0.03fF
C319 in_26 a_2450_7641# 0.00fF
C320 out en21_b 0.70fF
C321 a_2454_32182# VPWR 2.95fF
C322 in_24 en 1.38fF
C323 en7_b a_301_33465# 0.05fF
C324 out a_2454_38617# 7.60fF
C325 a_2454_9016# a_2450_10215# 0.10fF
C326 a_2454_5155# VPWR 2.95fF
C327 a_301_23169# a_2450_24372# 0.05fF
C328 a_2454_6442# a_2450_6354# 1.92fF
C329 a_2454_9016# en25_b 1.80fF
C330 en20_b a_2454_15451# 1.80fF
C331 out a_2454_19312# 7.60fF
C332 a_2454_18025# en17_b 0.03fF
C333 a_2450_5067# a_2454_3868# 0.10fF
C334 a_301_3864# a_301_5151# 0.39fF
C335 a_301_24456# a_301_27030# 0.03fF
C336 in_8 VPWR 1.24fF
C337 a_2454_6442# en27_b 1.80fF
C338 in_8 in_6 0.03fF
C339 en2_b en_b 0.05fF
C340 a_2450_34668# a_2450_33381# 0.18fF
C341 a_301_11586# a_301_9012# 0.03fF
C342 en_b a_2450_8928# 0.01fF
C343 en2_b en1_b 0.22fF
C344 a_2454_9016# VPWR 2.95fF
C345 in_30 in_31 0.28fF
C346 a_301_19308# a_301_21882# 0.03fF
C347 a_2450_19224# a_301_18021# 0.05fF
C348 a_2450_29520# a_2454_28321# 0.10fF
C349 a_2454_2581# a_2454_1294# 0.37fF
C350 a_2454_23173# a_301_21882# 0.08fF
C351 en18_b en17_b 0.22fF
C352 en3_b VPWR 3.16fF
C353 in_29 in_27 0.03fF
C354 a_2450_2493# en_b 0.01fF
C355 a_301_29604# a_2454_30895# 0.08fF
C356 a_2454_16738# a_2454_14164# 0.03fF
C357 a_2450_16650# in_19 0.00fF
C358 en_b a_2450_19224# 0.01fF
C359 a_2454_30895# en8_b 1.80fF
C360 a_301_29604# in_9 6.75fF
C361 a_301_19308# a_301_18021# 0.39fF
C362 a_301_29604# a_301_28317# 0.39fF
C363 a_301_16734# en19_b 1.19fF
C364 a_301_9012# a_301_10299# 0.39fF
C365 in_28 en_b 1.24fF
C366 en14_b a_2450_24372# 0.49fF
C367 a_2450_10215# en23_b 0.01fF
C368 a_301_19308# en_b 0.58fF
C369 in_15 en 1.38fF
C370 a_301_32178# en_b 0.58fF
C371 a_2450_21798# a_2454_23173# 0.03fF
C372 a_301_23169# a_301_21882# 0.39fF
C373 a_2454_34756# out 7.60fF
C374 a_2454_34756# en5_b 1.80fF
C375 a_2450_26946# a_301_25743# 0.05fF
C376 en2_b a_301_37326# 0.01fF
C377 a_2454_37330# in_3 0.05fF
C378 a_301_9012# en26_b 0.05fF
C379 in_3 a_301_38613# 0.08fF
C380 a_2450_20511# VPWR 0.55fF
C381 out a_2450_15363# 0.78fF
C382 in_17 a_2450_19224# 0.00fF
C383 a_2450_24372# a_301_25743# 0.01fF
C384 a_301_6438# en_b 0.58fF
C385 in_11 a_2450_26946# 0.00fF
C386 a_2450_26946# a_2454_28321# 0.03fF
C387 a_2450_21798# a_301_23169# 0.01fF
C388 en7_b en 0.01fF
C389 a_2454_15451# VPWR 2.95fF
C390 a_301_23169# en_b 0.58fF
C391 a_2454_9016# a_2450_7641# 0.03fF
C392 a_2450_12789# a_2450_11502# 0.18fF
C393 a_2450_23085# a_2454_23173# 1.92fF
C394 en22_b a_2454_11590# 0.03fF
C395 en23_b VPWR 3.16fF
C396 a_301_14160# in_22 0.08fF
C397 en0_b in_0 0.00fF
C398 en2_b a_2454_38617# 1.80fF
C399 a_301_19308# in_17 6.75fF
C400 en22_b en 0.01fF
C401 en0_b en_b 0.05fF
C402 a_2450_3780# a_301_3864# 1.32fF
C403 a_2450_3780# a_301_5151# 0.01fF
C404 a_2450_17937# a_301_18021# 1.32fF
C405 a_2454_30895# a_2454_32182# 0.37fF
C406 out a_301_24456# 0.43fF
C407 a_2450_2493# a_301_1290# 0.05fF
C408 a_301_10299# a_301_7725# 0.03fF
C409 en22_b a_2454_14164# 0.10fF
C410 a_2454_12877# VPWR 2.95fF
C411 a_2454_6442# a_2454_3868# 0.03fF
C412 en_b a_2450_17937# 0.01fF
C413 en0_b en1_b 0.22fF
C414 a_301_33465# a_2454_33469# 7.45fF
C415 a_2450_12789# en_b 0.01fF
C416 a_301_5151# a_2450_6354# 0.05fF
C417 a_301_23169# a_2450_23085# 1.32fF
C418 en en11_b 0.01fF
C419 en14_b a_301_21882# 0.01fF
C420 en25_b a_2454_7729# 0.03fF
C421 a_2454_30895# in_8 0.05fF
C422 a_301_7725# en26_b 1.19fF
C423 in_2 a_301_38613# 6.75fF
C424 a_301_16734# a_2450_16650# 1.32fF
C425 a_2450_28233# a_301_27030# 0.05fF
C426 in_9 in_8 0.28fF
C427 a_301_5151# en27_b 0.01fF
C428 a_301_34752# in_5 6.75fF
C429 in_27 VPWR 1.24fF
C430 a_301_24456# in_13 6.75fF
C431 a_2454_19312# a_2450_19224# 1.92fF
C432 en a_301_41187# 0.73fF
C433 a_301_33465# VPWR 3.21fF
C434 en a_301_39900# 0.79fF
C435 en20_b en 0.01fF
C436 a_2454_20599# a_2454_18025# 0.03fF
C437 in_29 en 1.38fF
C438 a_301_33465# in_6 6.75fF
C439 en_b a_2450_37242# 0.01fF
C440 en24_b a_301_9012# 0.01fF
C441 a_2450_21798# en14_b 0.01fF
C442 en20_b a_2454_14164# 0.03fF
C443 a_301_19308# a_2454_19312# 7.45fF
C444 a_301_2577# en29_b 0.01fF
C445 en14_b en_b 0.05fF
C446 VPWR a_2454_7729# 2.95fF
C447 a_2450_5067# en_b 0.01fF
C448 out en16_b 0.70fF
C449 a_2450_11502# in_23 0.00fF
C450 a_2450_32094# a_301_30891# 0.05fF
C451 a_2450_34668# a_301_34752# 1.32fF
C452 a_2454_21886# a_301_21882# 7.45fF
C453 en12_b a_2450_25659# 0.51fF
C454 in_21 in_20 0.28fF
C455 en30_b VPWR 3.16fF
C456 a_2454_29608# a_2450_28233# 0.03fF
C457 en_b a_301_25743# 0.58fF
C458 en14_b a_2450_23085# 0.51fF
C459 in_10 VPWR 1.24fF
C460 in_23 en_b 1.24fF
C461 a_2454_15451# en19_b 0.03fF
C462 a_2450_21798# a_2454_21886# 1.92fF
C463 in_16 en16_b 0.00fF
C464 a_2450_12789# en21_b 0.01fF
C465 a_2450_10215# a_2454_11590# 0.03fF
C466 out en17_b 0.70fF
C467 a_301_15447# a_301_18021# 0.03fF
C468 in_3 in_1 0.03fF
C469 a_2450_10215# en 0.06fF
C470 a_301_37326# a_2450_37242# 1.32fF
C471 a_301_36039# a_301_34752# 0.39fF
C472 en9_b a_2454_28321# 0.03fF
C473 a_2450_17937# a_2454_19312# 0.03fF
C474 en25_b en 0.01fF
C475 in_11 en_b 1.24fF
C476 en20_b a_2454_16738# 0.10fF
C477 en_b in_5 1.24fF
C478 a_301_15447# en_b 0.58fF
C479 a_301_18021# in_18 6.75fF
C480 a_2454_36043# a_2454_33469# 0.03fF
C481 a_301_24456# a_2454_25747# 0.08fF
C482 a_2450_7641# a_2454_7729# 1.92fF
C483 a_2454_21886# a_2450_23085# 0.10fF
C484 a_2450_39816# en_b 0.01fF
C485 out a_301_9012# 0.43fF
C486 en23_b a_301_12873# 0.05fF
C487 a_301_16734# a_2454_18025# 0.08fF
C488 in_19 in_21 0.03fF
C489 a_2454_11590# VPWR 2.95fF
C490 in_24 a_2450_10215# 0.00fF
C491 en_b in_18 1.24fF
C492 a_2450_37242# a_2454_38617# 0.03fF
C493 a_301_5151# a_2454_3868# 0.07fF
C494 a_301_3864# a_2454_3868# 7.45fF
C495 out a_2450_28233# 0.78fF
C496 en VPWR 32.43fF
C497 a_301_2577# a_2454_2581# 7.45fF
C498 en1_b a_2450_39816# 0.51fF
C499 en in_6 1.38fF
C500 in_26 en26_b 0.00fF
C501 out en15_b 0.70fF
C502 a_2454_36043# VPWR 2.95fF
C503 a_2450_6354# en27_b 0.51fF
C504 a_2454_14164# VPWR 2.95fF
C505 a_301_12873# a_2454_12877# 7.45fF
C506 a_2454_27034# a_2450_28233# 0.10fF
C507 a_2450_34668# en_b 0.01fF
C508 in_2 in_1 0.28fF
C509 a_2454_39904# a_301_41187# 0.07fF
C510 a_2454_23173# a_301_24456# 0.07fF
C511 in_24 VPWR 1.24fF
C512 a_2454_39904# a_301_39900# 7.45fF
C513 out en6_b 0.70fF
C514 a_301_16734# en18_b 0.01fF
C515 out en4_b 0.70fF
C516 en5_b en6_b 0.22fF
C517 en5_b en4_b 0.22fF
C518 in_17 in_18 0.28fF
C519 a_2450_16650# a_2454_15451# 0.10fF
C520 a_301_29604# a_301_30891# 0.39fF
C521 a_301_30891# en8_b 1.19fF
C522 out en28_b 0.70fF
C523 out a_301_7725# 0.43fF
C524 en31_b a_2454_2581# 0.10fF
C525 out a_301_38613# 0.43fF
C526 a_301_36039# en_b 0.58fF
C527 out en29_b 0.70fF
C528 a_2454_21886# a_2454_19312# 0.03fF
C529 a_2454_37330# out 7.60fF
C530 a_301_20595# a_301_21882# 0.39fF
C531 a_301_23169# a_301_24456# 0.39fF
C532 a_301_15447# en21_b 0.05fF
C533 en13_b a_2450_24372# 0.51fF
C534 a_2450_7641# en 0.06fF
C535 out a_2450_32094# 0.78fF
C536 a_301_29604# a_301_27030# 0.03fF
C537 a_2454_16738# VPWR 2.95fF
C538 a_301_14160# en_b 0.58fF
C539 en16_b a_2450_19224# 0.01fF
C540 in_3 en3_b 0.00fF
C541 a_301_20595# a_301_18021# 0.03fF
C542 in_10 a_301_28317# 6.75fF
C543 a_2450_35955# a_301_34752# 0.05fF
C544 in_10 in_9 0.28fF
C545 a_301_20595# a_2450_21798# 0.05fF
C546 a_301_39900# a_301_41187# 0.39fF
C547 a_2450_39816# a_2454_38617# 0.10fF
C548 a_301_20595# en_b 0.58fF
C549 a_301_19308# en16_b 0.01fF
C550 en_b a_2450_14076# 0.01fF
C551 en30_b a_2454_1294# 0.03fF
C552 in_15 VPWR 1.24fF
C553 a_301_30891# a_2454_32182# 0.08fF
C554 en12_b a_301_27030# 0.05fF
C555 en en19_b 0.01fF
C556 a_2454_9016# a_301_10299# 0.07fF
C557 a_2450_11502# a_2454_10303# 0.10fF
C558 a_301_9012# a_2450_8928# 1.32fF
C559 en7_b a_2454_33469# 0.10fF
C560 a_2450_3780# a_2454_3868# 1.92fF
C561 en17_b a_2450_19224# 0.51fF
C562 a_301_36039# a_301_37326# 0.39fF
C563 en in_4 1.38fF
C564 out a_2454_20599# 7.60fF
C565 a_2454_2581# in_30 0.05fF
C566 a_2454_9016# en26_b 0.10fF
C567 en14_b a_301_24456# 0.05fF
C568 a_2454_36043# in_4 0.05fF
C569 a_301_19308# en17_b 1.19fF
C570 in_14 en 1.38fF
C571 a_2454_29608# a_301_29604# 7.45fF
C572 in_8 a_301_30891# 6.75fF
C573 a_301_20595# in_17 0.08fF
C574 a_2454_29608# en8_b 0.03fF
C575 in_9 en 1.38fF
C576 en a_301_28317# 0.79fF
C577 a_301_11586# en23_b 1.19fF
C578 en7_b VPWR 3.16fF
C579 a_2454_39904# VPWR 2.95fF
C580 a_2450_29520# a_2450_30807# 0.18fF
C581 a_301_12873# a_2454_11590# 0.07fF
C582 a_2454_34756# in_5 0.05fF
C583 a_2454_15451# a_2454_18025# 0.03fF
C584 a_301_12873# en 0.79fF
C585 en22_b VPWR 3.16fF
C586 in_7 a_2450_32094# 0.00fF
C587 out a_2454_2581# 7.60fF
C588 a_301_11586# a_2454_12877# 0.08fF
C589 in_16 a_2454_20599# 0.05fF
C590 a_301_24456# a_301_25743# 0.39fF
C591 a_301_12873# a_2454_14164# 0.08fF
C592 a_301_14160# en21_b 1.19fF
C593 a_2450_15363# a_301_15447# 1.32fF
C594 a_301_7725# a_2450_8928# 0.05fF
C595 en2_b a_301_38613# 1.19fF
C596 a_2450_35955# en_b 0.01fF
C597 a_2450_29520# en10_b 0.49fF
C598 en13_b en_b 0.05fF
C599 a_2454_37330# en2_b 0.03fF
C600 en11_b VPWR 3.16fF
C601 a_301_3864# en_b 0.58fF
C602 en_b a_301_5151# 0.58fF
C603 en15_b a_2454_23173# 0.10fF
C604 en23_b a_301_10299# 0.01fF
C605 en21_b a_2450_14076# 0.51fF
C606 a_2454_16738# en19_b 1.80fF
C607 a_301_6438# a_301_9012# 0.03fF
C608 a_2454_34756# a_2450_34668# 1.92fF
C609 a_2450_17937# en17_b 0.01fF
C610 out en8_b 0.70fF
C611 out a_301_29604# 0.43fF
C612 a_301_20595# a_2454_19312# 0.07fF
C613 a_301_41187# VPWR 3.33fF
C614 en20_b VPWR 3.16fF
C615 a_2450_16650# en 0.06fF
C616 a_301_39900# VPWR 3.21fF
C617 a_2454_29608# a_2454_32182# 0.03fF
C618 in_29 VPWR 1.24fF
C619 a_2450_2493# en29_b 0.01fF
C620 en13_b a_2450_23085# 0.01fF
C621 en6_b a_301_32178# 0.01fF
C622 in_28 en28_b 0.00fF
C623 a_301_23169# en15_b 0.05fF
C624 en24_b a_2454_9016# 0.03fF
C625 a_301_16734# out 0.43fF
C626 en_b a_2450_1206# 0.01fF
C627 a_2454_34756# a_301_36039# 0.07fF
C628 out en12_b 0.70fF
C629 a_2450_10215# en25_b 0.49fF
C630 a_2450_35955# a_301_37326# 0.01fF
C631 a_2450_26946# en10_b 0.01fF
C632 in_14 in_15 0.28fF
C633 en a_2450_25659# 0.06fF
C634 a_2454_27034# en12_b 0.10fF
C635 a_2454_21886# en16_b 0.10fF
C636 en_b a_2450_38529# 0.01fF
C637 en28_b a_301_6438# 0.05fF
C638 a_2450_32094# a_301_32178# 1.32fF
C639 a_301_6438# a_301_7725# 0.39fF
C640 en1_b a_2450_38529# 0.01fF
C641 out a_2454_32182# 7.60fF
C642 a_301_3864# a_301_1290# 0.03fF
C643 a_2450_10215# VPWR 0.55fF
C644 a_2454_5155# out 7.60fF
C645 a_2454_24460# VPWR 2.95fF
C646 en25_b VPWR 3.16fF
C647 a_2450_33381# a_301_34752# 0.01fF
C648 en26_b a_2454_7729# 1.80fF
C649 a_301_14160# a_2450_15363# 0.05fF
C650 en7_b a_2454_30895# 0.03fF
C651 a_2454_33469# VPWR 2.95fF
C652 a_2450_16650# a_2454_16738# 1.92fF
C653 a_2454_20599# a_2450_19224# 0.03fF
C654 en15_b en14_b 0.22fF
C655 a_301_33465# a_301_30891# 0.03fF
C656 in_6 a_2454_33469# 0.05fF
C657 en24_b en23_b 0.22fF
C658 a_2450_15363# a_2450_14076# 0.18fF
C659 a_301_11586# a_2454_11590# 7.45fF
C660 in_3 en 1.38fF
C661 a_301_19308# a_2454_20599# 0.08fF
C662 a_2450_1206# a_301_1290# 1.33fF
C663 a_301_11586# en 0.79fF
C664 a_2450_3780# en_b 0.01fF
C665 a_2450_2493# a_2454_2581# 1.92fF
C666 en22_b a_301_12873# 1.19fF
C667 a_2454_23173# a_2454_20599# 0.03fF
C668 in_12 en_b 1.24fF
C669 out a_2454_9016# 7.60fF
C670 en20_b en19_b 0.22fF
C671 en4_b a_2450_37242# 0.49fF
C672 a_301_37326# a_2450_38529# 0.05fF
C673 in_6 VPWR 1.24fF
C674 en11_b a_301_28317# 0.05fF
C675 en_b a_2450_6354# 0.01fF
C676 out en3_b 0.70fF
C677 en30_b a_301_2577# 1.19fF
C678 a_2450_37242# a_301_38613# 0.01fF
C679 a_2454_37330# a_2450_37242# 1.92fF
C680 en_b en27_b 0.05fF
C681 a_2450_28233# a_2454_28321# 1.92fF
C682 in_25 en_b 1.24fF
C683 en9_b a_2450_30807# 0.49fF
C684 a_2454_21886# en15_b 1.80fF
C685 a_301_11586# in_24 0.08fF
C686 a_2450_30807# en_b 0.01fF
C687 a_2450_5067# en28_b 0.51fF
C688 a_2454_11590# a_301_10299# 0.08fF
C689 in_7 a_2454_32182# 0.05fF
C690 en25_b a_2450_7641# 0.01fF
C691 a_2450_5067# en29_b 0.49fF
C692 a_2450_38529# a_2454_38617# 1.92fF
C693 en a_301_10299# 0.79fF
C694 a_2454_34756# a_2450_35955# 0.10fF
C695 in_28 in_26 0.03fF
C696 en18_b en 0.01fF
C697 en12_b a_2454_25747# 1.80fF
C698 out a_2450_20511# 0.78fF
C699 en en26_b 0.01fF
C700 in_2 en 1.38fF
C701 a_2450_33381# en_b 0.01fF
C702 en9_b en10_b 0.22fF
C703 en_b en10_b 0.05fF
C704 in_10 a_301_27030# 0.07fF
C705 in_7 in_8 0.28fF
C706 a_301_32178# en8_b 0.05fF
C707 a_301_29604# a_301_32178# 0.03fF
C708 en31_b en30_b 0.22fF
C709 a_2450_7641# VPWR 0.55fF
C710 out en23_b 0.70fF
C711 out a_2454_15451# 7.60fF
C712 in_24 a_301_10299# 6.75fF
C713 a_301_20595# en16_b 1.19fF
C714 a_301_2577# en 0.79fF
C715 a_2450_1206# in_31 0.00fF
C716 a_301_6438# in_26 0.07fF
C717 a_301_30891# en 0.79fF
C718 a_2454_16738# a_2454_18025# 0.37fF
C719 a_301_16734# a_301_19308# 0.03fF
C720 in_22 en_b 1.24fF
C721 in_16 a_2450_20511# 0.00fF
C722 en20_b a_2450_16650# 0.49fF
C723 out a_2454_12877# 7.60fF
C724 en13_b a_301_24456# 1.19fF
C725 a_301_15447# in_20 6.75fF
C726 a_2454_30895# a_2454_33469# 0.03fF
C727 en in_21 1.38fF
C728 en19_b VPWR 3.16fF
C729 a_2450_39816# a_301_38613# 0.05fF
C730 en a_301_27030# 0.79fF
C731 en6_b a_2450_34668# 0.49fF
C732 in_4 VPWR 1.24fF
C733 a_301_20595# en17_b 0.05fF
C734 en11_b a_2450_25659# 0.01fF
C735 in_21 a_2454_14164# 0.05fF
C736 in_20 in_18 0.03fF
C737 a_2450_34668# en4_b 0.01fF
C738 in_6 in_4 0.03fF
C739 a_2454_9016# a_2450_8928# 1.92fF
C740 out a_301_33465# 0.43fF
C741 a_301_32178# a_2454_32182# 7.45fF
C742 a_2454_5155# in_28 0.05fF
C743 a_2454_16738# en18_b 0.03fF
C744 en5_b a_301_33465# 0.01fF
C745 a_2450_29520# en9_b 0.51fF
C746 en2_b en3_b 0.22fF
C747 in_14 VPWR 1.24fF
C748 a_2454_30895# VPWR 2.95fF
C749 en31_b en 0.01fF
C750 a_2450_29520# en_b 0.01fF
C751 a_301_28317# VPWR 3.21fF
C752 in_9 VPWR 1.24fF
C753 en24_b a_2454_11590# 0.10fF
C754 en30_b in_30 0.00fF
C755 out a_2454_7729# 7.60fF
C756 en24_b en 0.01fF
C757 a_2454_21886# a_2454_20599# 0.37fF
C758 a_301_11586# en22_b 0.01fF
C759 a_301_16734# a_2450_17937# 0.05fF
C760 a_301_32178# in_8 0.08fF
C761 a_301_12873# VPWR 3.21fF
C762 a_301_36039# en4_b 1.19fF
C763 en28_b a_2454_6442# 0.10fF
C764 a_2454_6442# a_301_7725# 0.07fF
C765 a_2454_1294# VPWR 2.78fF
C766 a_301_20595# en15_b 0.01fF
C767 in_19 a_301_15447# 0.07fF
C768 a_2454_5155# a_301_6438# 0.07fF
C769 a_301_36039# a_301_38613# 0.03fF
C770 out en30_b 0.70fF
C771 a_2454_37330# a_301_36039# 0.08fF
C772 en24_b in_24 0.00fF
C773 in_19 in_18 0.28fF
C774 a_301_9012# a_2454_10303# 0.08fF
C775 a_2450_26946# en_b 0.01fF
C776 a_2450_16650# VPWR 0.55fF
C777 a_301_14160# in_20 0.07fF
C778 en in_30 1.38fF
C779 in_7 a_301_33465# 0.08fF
C780 a_2454_24460# a_2450_25659# 0.10fF
C781 a_2450_20511# a_2450_19224# 0.18fF
C782 en_b a_2450_24372# 0.01fF
C783 in_12 a_301_24456# 0.07fF
C784 a_301_29604# a_2454_28321# 0.07fF
C785 en7_b a_301_30891# 0.01fF
C786 out a_2454_11590# 7.60fF
C787 a_301_19308# a_2450_20511# 0.05fF
C788 en12_b a_301_25743# 1.19fF
C789 a_301_34752# en_b 0.58fF
C790 a_2454_34756# a_2450_33381# 0.03fF
C791 en5_b en 0.01fF
C792 a_2450_25659# VPWR 0.55fF
C793 out a_2454_14164# 7.60fF
C794 out a_2454_36043# 7.60fF
C795 en5_b a_2454_36043# 0.10fF
C796 a_2450_23085# a_2450_24372# 0.18fF
C797 a_2454_5155# a_2450_5067# 1.92fF
C798 a_301_16734# a_301_15447# 0.39fF
C799 in_1 a_2450_39816# 0.00fF
C800 in_2 a_301_39900# 0.08fF
C801 a_301_11586# a_2450_10215# 0.01fF
C802 a_2450_8928# a_2454_7729# 0.10fF
C803 en in_13 1.38fF
C804 in_16 en 1.38fF
C805 in_9 a_301_28317# 0.07fF
C806 a_2450_35955# en4_b 0.51fF
C807 in_28 in_27 0.28fF
C808 a_301_20595# a_2454_20599# 7.45fF
C809 a_301_16734# in_18 0.07fF
C810 en3_b a_2450_37242# 0.51fF
C811 in_29 a_301_2577# 0.07fF
C812 a_2450_21798# a_301_21882# 1.32fF
C813 en_b a_301_21882# 0.58fF
C814 a_2454_37330# a_2450_35955# 0.03fF
C815 en28_b a_301_3864# 0.01fF
C816 en28_b a_301_5151# 1.19fF
C817 a_301_34752# a_301_37326# 0.03fF
C818 a_301_5151# a_301_7725# 0.03fF
C819 en11_b a_301_27030# 1.19fF
C820 a_2450_11502# en_b 0.01fF
C821 in_3 VPWR 1.24fF
C822 a_2450_41103# en 0.06fF
C823 a_301_33465# a_301_32178# 0.39fF
C824 a_301_3864# en29_b 1.19fF
C825 a_301_5151# en29_b 0.05fF
C826 a_301_11586# VPWR 3.21fF
C827 a_2450_10215# a_301_10299# 1.32fF
C828 a_2450_16650# en19_b 0.51fF
C829 a_2450_12789# en23_b 0.49fF
C830 en25_b a_301_10299# 0.05fF
C831 a_2454_16738# out 7.60fF
C832 a_2454_18025# VPWR 2.95fF
C833 en_b a_301_18021# 0.58fF
C834 a_2454_41191# a_2454_39904# 0.37fF
C835 in_0 en_b 1.28fF
C836 in_7 en 1.38fF
C837 en30_b a_2450_2493# 0.51fF
C838 a_301_6438# in_27 6.75fF
C839 a_2450_21798# en_b 0.01fF
C840 en9_b en_b 0.05fF
C841 a_2450_23085# a_301_21882# 0.05fF
C842 en25_b en26_b 0.22fF
C843 a_2450_12789# a_2454_12877# 1.92fF
C844 en1_b en_b 0.05fF
C845 a_301_6438# a_2454_7729# 0.08fF
C846 a_301_10299# VPWR 3.21fF
C847 en2_b en 0.01fF
C848 en a_2450_8928# 0.06fF
C849 a_2450_21798# a_2450_23085# 0.18fF
C850 a_2450_23085# en_b 0.01fF
C851 en18_b VPWR 3.16fF
C852 in_17 a_301_18021# 0.07fF
C853 en26_b VPWR 3.16fF
C854 in_2 VPWR 1.24fF
C855 a_301_16734# a_301_14160# 0.03fF
C856 a_2450_38529# a_301_38613# 1.32fF
C857 a_2454_37330# a_2450_38529# 0.10fF
C858 in_17 en_b 1.24fF
C859 a_2454_41191# a_301_41187# 7.45fF
C860 a_2454_41191# a_301_39900# 0.08fF
C861 in_15 in_13 0.03fF
C862 out a_2454_39904# 7.60fF
C863 in_16 in_15 0.28fF
C864 en7_b out 0.70fF
C865 a_2454_5155# a_2454_6442# 0.37fF
C866 a_2450_2493# en 0.06fF
C867 a_2454_21886# a_2450_20511# 0.03fF
C868 a_301_37326# en_b 0.58fF
C869 in_25 a_301_9012# 6.75fF
C870 out en22_b 0.70fF
C871 a_301_2577# VPWR 3.21fF
C872 a_301_30891# VPWR 3.21fF
C873 in_23 en23_b 0.00fF
C874 en a_2450_19224# 0.06fF
C875 in_28 en 1.38fF
C876 en_b a_301_1290# 0.51fF
C877 a_2454_2581# a_301_3864# 0.07fF
C878 a_301_19308# en 0.79fF
C879 a_2454_34756# a_301_34752# 7.45fF
C880 en24_b a_2450_10215# 0.51fF
C881 in_29 in_30 0.28fF
C882 a_301_32178# en 0.79fF
C883 in_21 VPWR 1.24fF
C884 out en11_b 0.70fF
C885 en28_b a_2450_3780# 0.01fF
C886 a_2454_19312# a_301_18021# 0.08fF
C887 in_3 in_4 0.28fF
C888 en24_b en25_b 0.22fF
C889 a_2454_15451# a_301_15447# 7.45fF
C890 en21_b en_b 0.05fF
C891 a_2454_9016# a_2454_6442# 0.03fF
C892 a_2454_18025# en19_b 0.10fF
C893 a_2450_3780# en29_b 0.51fF
C894 a_301_27030# VPWR 3.21fF
C895 en28_b a_2450_6354# 0.49fF
C896 en1_b a_2454_38617# 0.03fF
C897 a_2454_27034# en11_b 1.80fF
C898 out a_301_41187# 0.43fF
C899 a_2450_28233# en10_b 0.51fF
C900 en20_b out 0.70fF
C901 a_2450_6354# a_301_7725# 0.01fF
C902 out a_301_39900# 0.43fF
C903 a_2450_7641# en26_b 0.51fF
C904 a_301_6438# en 0.79fF
C905 en31_b VPWR 2.84fF
C906 en3_b a_301_36039# 0.01fF
C907 a_301_24456# a_2450_24372# 1.32fF
C908 a_2450_41103# a_2454_39904# 0.10fF
C909 a_301_23169# en 0.79fF
C910 en28_b en27_b 0.22fF
C911 a_301_7725# en27_b 0.05fF
C912 a_2454_2581# a_2450_1206# 0.03fF
C913 en24_b VPWR 3.16fF
C914 in_25 a_301_7725# 0.07fF
C915 a_301_11586# a_301_12873# 0.39fF
C916 en0_b en 0.01fF
C917 en7_b in_7 0.00fF
C918 en6_b a_2450_33381# 0.51fF
C919 a_2450_12789# a_2454_11590# 0.10fF
C920 en18_b en19_b 0.22fF
C921 en a_2450_17937# 0.06fF
C922 in_17 a_2454_19312# 0.05fF
C923 a_2450_12789# en 0.06fF
C924 a_301_33465# in_5 0.07fF
C925 en13_b en12_b 0.22fF
C926 a_2450_32094# a_2450_30807# 0.18fF
C927 a_2454_41191# VPWR 3.05fF
C928 a_2454_29608# VPWR 2.95fF
C929 a_301_37326# a_2454_38617# 0.08fF
C930 in_2 in_4 0.03fF
C931 a_2450_12789# a_2454_14164# 0.03fF
C932 en_b in_31 1.17fF
C933 en2_b a_2454_39904# 0.10fF
C934 a_2450_41103# a_301_41187# 1.32fF
C935 a_301_12873# a_301_10299# 0.03fF
C936 a_2450_41103# a_301_39900# 0.05fF
C937 out a_2450_10215# 0.78fF
C938 a_2450_29520# a_2450_28233# 0.18fF
C939 a_2454_24460# out 7.60fF
C940 a_2450_32094# a_2450_33381# 0.18fF
C941 en a_2450_37242# 0.06fF
C942 a_2454_9016# a_2454_10303# 0.37fF
C943 out en25_b 0.70fF
C944 en14_b en 0.01fF
C945 in_30 VPWR 1.24fF
C946 in_10 a_2454_28321# 0.05fF
C947 a_2450_16650# a_2454_18025# 0.03fF
C948 out a_2454_33469# 7.60fF
C949 a_2454_5155# a_301_3864# 0.08fF
C950 a_2454_5155# a_301_5151# 7.45fF
C951 a_301_33465# a_2450_34668# 0.05fF
C952 a_301_24456# a_301_21882# 0.03fF
C953 in_11 in_10 0.28fF
C954 en5_b a_2454_33469# 0.03fF
C955 a_2454_36043# a_2450_37242# 0.10fF
C956 a_2454_24460# a_2454_27034# 0.03fF
C957 a_2454_2581# a_2450_3780# 0.10fF
C958 a_301_20595# a_2450_20511# 1.32fF
C959 a_2450_15363# en_b 0.01fF
C960 in_22 in_20 0.03fF
C961 a_2450_5067# en 0.06fF
C962 a_301_14160# a_2454_15451# 0.08fF
C963 a_2454_30895# a_301_30891# 7.45fF
C964 a_301_30891# a_301_28317# 0.03fF
C965 in_9 a_301_30891# 0.08fF
C966 in_27 a_2454_6442# 0.05fF
C967 a_2454_15451# a_2450_14076# 0.03fF
C968 a_2454_24460# in_13 0.05fF
C969 a_301_14160# a_2454_12877# 0.07fF
C970 out VPWR 53.27fF
C971 in_23 a_2454_11590# 0.05fF
C972 a_2454_25747# en11_b 0.03fF
C973 en a_301_25743# 0.79fF
C974 en5_b VPWR 3.16fF
C975 a_2454_16738# a_2450_17937# 0.10fF
C976 a_301_24456# en_b 0.58fF
C977 a_301_33465# a_301_36039# 0.03fF
C978 a_301_23169# in_15 0.08fF
C979 in_23 en 1.38fF
C980 en7_b a_301_32178# 1.19fF
C981 a_301_2577# a_2454_1294# 0.07fF
C982 en2_b a_301_39900# 0.05fF
C983 en3_b a_2450_35955# 0.01fF
C984 a_2450_16650# en18_b 0.01fF
C985 a_2454_27034# VPWR 2.95fF
C986 a_2454_6442# a_2454_7729# 0.37fF
C987 a_301_28317# a_301_27030# 0.39fF
C988 en28_b a_2454_3868# 0.03fF
C989 a_2454_12877# a_2450_14076# 0.10fF
C990 a_301_1290# in_31 6.75fF
C991 a_301_12873# in_21 0.07fF
C992 a_2450_26946# a_2450_28233# 0.18fF
C993 en29_b a_2454_3868# 1.80fF
C994 in_11 en 1.38fF
C995 in_13 VPWR 1.24fF
C996 in_16 VPWR 1.24fF
C997 en in_5 1.38fF
C998 a_301_15447# en 0.79fF
C999 a_2454_10303# en23_b 0.03fF
C1000 a_2450_23085# a_301_24456# 0.01fF
C1001 in_25 in_26 0.28fF
C1002 in_24 in_23 0.28fF
C1003 en16_b a_301_21882# 0.05fF
C1004 a_301_15447# a_2454_14164# 0.07fF
C1005 a_2450_30807# en8_b 0.51fF
C1006 a_301_29604# a_2450_30807# 0.05fF
C1007 en a_2450_39816# 0.06fF
C1008 en0_b a_2454_39904# 0.03fF
C1009 en31_b a_2454_1294# 1.77fF
C1010 in_12 en12_b 0.00fF
C1011 en in_18 1.38fF
C1012 a_2454_10303# a_2454_12877# 0.03fF
C1013 a_2450_41103# VPWR 0.54fF
C1014 in_28 in_29 0.28fF
C1015 a_2450_15363# en21_b 0.49fF
C1016 out a_2450_7641# 0.78fF
C1017 a_2450_21798# en16_b 0.49fF
C1018 a_2454_29608# a_2454_30895# 0.37fF
C1019 en16_b en_b 0.05fF
C1020 a_2454_29608# in_9 0.05fF
C1021 a_2450_34668# en 0.06fF
C1022 a_2454_29608# a_301_28317# 0.08fF
C1023 in_7 VPWR 1.24fF
C1024 a_2450_12789# en22_b 0.51fF
C1025 a_2450_10215# a_2450_8928# 0.18fF
C1026 a_301_29604# en10_b 0.05fF
C1027 in_7 in_6 0.28fF
C1028 en25_b a_2450_8928# 0.51fF
C1029 a_2454_5155# a_2450_3780# 0.03fF
C1030 a_2454_36043# a_2450_34668# 0.03fF
C1031 a_2454_24460# a_2454_25747# 0.37fF
C1032 en3_b a_2450_38529# 0.49fF
C1033 en6_b a_301_34752# 0.05fF
C1034 en17_b a_301_18021# 0.01fF
C1035 en4_b a_301_34752# 0.01fF
C1036 a_2454_5155# a_2450_6354# 0.10fF
C1037 a_301_11586# a_301_10299# 0.39fF
C1038 a_2454_10303# a_2454_7729# 0.03fF
C1039 out en19_b 0.70fF
C1040 en0_b a_301_41187# 1.24fF
C1041 a_2454_16738# a_301_15447# 0.08fF
C1042 en0_b a_301_39900# 0.01fF
C1043 en_b en17_b 0.05fF
C1044 en2_b VPWR 3.16fF
C1045 a_301_36039# en 0.79fF
C1046 a_2450_30807# a_2454_32182# 0.03fF
C1047 a_2450_8928# VPWR 0.55fF
C1048 a_2454_5155# en27_b 0.03fF
C1049 in_3 in_2 0.28fF
C1050 a_2450_25659# a_301_27030# 0.01fF
C1051 in_27 a_301_5151# 0.07fF
C1052 a_2454_2581# a_2454_3868# 0.37fF
C1053 a_2454_36043# a_301_36039# 7.45fF
C1054 a_2454_21886# in_15 0.05fF
C1055 en18_b a_2454_18025# 1.80fF
C1056 en15_b a_301_21882# 1.19fF
C1057 a_2454_25747# VPWR 2.95fF
C1058 out a_2454_30895# 7.60fF
C1059 out a_301_28317# 0.43fF
C1060 a_2454_24460# a_2454_23173# 0.37fF
C1061 in_8 a_2450_30807# 0.00fF
C1062 a_301_14160# en 0.79fF
C1063 a_301_9012# en_b 0.58fF
C1064 a_301_32178# a_2454_33469# 0.08fF
C1065 a_2450_33381# a_2454_32182# 0.10fF
C1066 a_2454_27034# a_301_28317# 0.07fF
C1067 a_2450_2493# VPWR 0.55fF
C1068 out a_301_12873# 0.43fF
C1069 en9_b a_2450_28233# 0.01fF
C1070 a_2450_28233# en_b 0.01fF
C1071 a_301_14160# a_2454_14164# 7.45fF
C1072 a_2450_29520# a_301_29604# 1.32fF
C1073 a_2450_19224# VPWR 0.55fF
C1074 a_2450_29520# en8_b 0.01fF
C1075 a_301_20595# en 0.79fF
C1076 a_2450_21798# en15_b 0.51fF
C1077 out a_2454_1294# 7.49fF
C1078 en15_b en_b 0.05fF
C1079 en a_2450_14076# 0.06fF
C1080 in_17 en17_b 0.00fF
C1081 a_2454_9016# in_25 0.05fF
C1082 in_14 in_13 0.28fF
C1083 in_14 in_16 0.03fF
C1084 in_28 VPWR 1.24fF
C1085 a_301_19308# VPWR 3.21fF
C1086 a_2454_24460# a_301_23169# 0.08fF
C1087 a_2450_14076# a_2454_14164# 1.92fF
C1088 en16_b a_2454_19312# 0.03fF
C1089 a_301_32178# VPWR 3.21fF
C1090 a_2454_23173# VPWR 2.95fF
C1091 en30_b a_301_3864# 0.05fF
C1092 en11_b a_301_25743# 0.01fF
C1093 a_301_32178# in_6 0.07fF
C1094 en6_b en_b 0.05fF
C1095 en15_b a_2450_23085# 0.49fF
C1096 en4_b en_b 0.05fF
C1097 a_2454_10303# a_2454_11590# 0.37fF
C1098 a_2450_7641# a_2450_8928# 0.18fF
C1099 a_2454_39904# a_2450_39816# 1.92fF
C1100 a_2450_16650# out 0.78fF
C1101 en28_b en_b 0.05fF
C1102 a_301_6438# VPWR 3.21fF
C1103 en_b a_301_7725# 0.58fF
C1104 a_2454_28321# en11_b 0.10fF
C1105 en_b a_301_38613# 0.58fF
C1106 a_301_23169# VPWR 3.21fF
C1107 in_11 en11_b 0.00fF
C1108 a_301_11586# en24_b 0.05fF
C1109 en_b en29_b 0.05fF
C1110 a_2454_19312# en17_b 1.80fF
C1111 en_b in_20 1.24fF
C1112 en1_b a_301_38613# 0.01fF
C1113 in_7 in_9 0.03fF
C1114 en0_b VPWR 3.67fF
C1115 en30_b a_2450_1206# 0.01fF
C1116 a_2450_32094# en_b 0.01fF
C1117 a_2450_17937# VPWR 0.55fF
C1118 in_24 a_2454_10303# 0.05fF
C1119 en20_b a_301_15447# 1.19fF
C1120 a_2450_35955# en 0.06fF
C1121 a_2450_12789# VPWR 0.55fF
C1122 a_2454_5155# a_2454_3868# 0.37fF
C1123 en13_b en 0.01fF
C1124 a_2454_24460# en14_b 0.10fF
C1125 out a_2450_25659# 0.78fF
C1126 a_301_3864# en 0.79fF
C1127 a_2454_20599# a_301_21882# 0.07fF
C1128 en a_301_5151# 0.79fF
C1129 a_2454_36043# a_2450_35955# 1.92fF
C1130 a_2450_39816# a_301_41187# 0.01fF
C1131 a_2450_26946# en12_b 0.49fF
C1132 a_2450_39816# a_301_39900# 1.32fF
C1133 en4_b a_301_37326# 0.05fF
C1134 en24_b a_301_10299# 1.19fF
C1135 a_2454_27034# a_2450_25659# 0.03fF
C1136 in_27 a_2450_6354# 0.00fF
C1137 a_301_20595# in_15 0.07fF
C1138 in_19 a_301_18021# 0.08fF
C1139 a_301_37326# a_301_38613# 0.39fF
C1140 a_2450_37242# VPWR 0.55fF
C1141 a_2454_37330# a_301_37326# 7.45fF
C1142 en12_b a_2450_24372# 0.01fF
C1143 a_2454_24460# a_301_25743# 0.07fF
C1144 in_27 en27_b 0.00fF
C1145 a_301_6438# a_2450_7641# 0.05fF
C1146 a_2450_21798# a_2454_20599# 0.10fF
C1147 en14_b VPWR 3.16fF
C1148 in_19 en_b 1.24fF
C1149 in_25 in_27 0.03fF
C1150 en a_2450_1206# 0.05fF
C1151 en31_b a_301_2577# 0.05fF
C1152 a_2450_6354# a_2454_7729# 0.03fF
C1153 a_2454_24460# a_2454_21886# 0.03fF
C1154 a_2450_5067# VPWR 0.55fF
C1155 a_301_14160# en22_b 0.05fF
C1156 a_301_11586# out 0.43fF
C1157 en30_b a_2450_3780# 0.49fF
C1158 en27_b a_2454_7729# 0.10fF
C1159 a_301_38613# a_2454_38617# 7.45fF
C1160 a_2454_37330# a_2454_38617# 0.37fF
C1161 in_14 a_2454_23173# 0.05fF
C1162 a_301_32178# a_2454_30895# 0.07fF
C1163 a_2450_2493# a_2454_1294# 0.10fF
C1164 out a_2454_18025# 7.60fF
C1165 VPWR a_301_25743# 3.21fF
C1166 en22_b a_2450_14076# 0.49fF
C1167 in_12 in_10 0.03fF
C1168 en a_2450_38529# 0.06fF
C1169 in_23 VPWR 1.24fF
C1170 in_22 a_2454_12877# 0.05fF
C1171 a_301_33465# a_2450_33381# 1.32fF
C1172 in_19 in_17 0.03fF
C1173 a_2454_21886# VPWR 2.95fF
C1174 a_2454_29608# a_301_30891# 0.07fF
C1175 a_2454_28321# VPWR 2.95fF
C1176 in_11 VPWR 1.24fF
C1177 in_14 a_301_23169# 6.75fF
C1178 in_26 en_b 1.24fF
C1179 en20_b a_301_14160# 0.01fF
C1180 in_5 VPWR 1.24fF
C1181 en19_b a_2450_17937# 0.49fF
C1182 a_301_15447# VPWR 3.21fF
C1183 a_301_29604# en_b 0.58fF
C1184 out a_301_10299# 0.43fF
C1185 in_0 in_1 0.28fF
C1186 en9_b en8_b 0.22fF
C1187 a_301_29604# en9_b 1.19fF
C1188 in_6 in_5 0.28fF
C1189 en8_b en_b 0.05fF
C1190 in_1 en_b 1.24fF
C1191 a_2450_34668# a_2454_33469# 0.10fF
C1192 out en18_b 0.70fF
C1193 en20_b a_2450_14076# 0.01fF
C1194 a_301_2577# in_30 6.75fF
C1195 a_2450_39816# VPWR 0.55fF
C1196 a_301_16734# a_301_18021# 0.39fF
C1197 VPWR in_18 1.24fF
C1198 a_2450_3780# en 0.06fF
C1199 out en26_b 0.70fF
C1200 a_2454_34756# en6_b 0.10fF
C1201 en1_b in_1 0.00fF
C1202 a_2454_34756# en4_b 0.03fF
C1203 in_12 en 1.38fF
C1204 a_2454_25747# a_2450_25659# 1.92fF
C1205 a_301_16734# en_b 0.58fF
C1206 in_10 en10_b 0.00fF
C1207 en a_2450_6354# 0.06fF
C1208 a_2454_20599# a_2454_19312# 0.37fF
C1209 en12_b en_b 0.05fF
C1210 a_2450_12789# a_301_12873# 1.32fF
C1211 a_2454_2581# a_301_1290# 0.08fF
C1212 a_2450_34668# VPWR 0.55fF
C1213 a_2454_37330# a_2454_34756# 0.03fF
C1214 out a_301_2577# 0.43fF
C1215 en en27_b 0.01fF
C1216 out a_301_30891# 0.43fF
C1217 in_25 en 1.38fF
C1218 a_2450_30807# en 0.06fF
C1219 en16_b en17_b 0.22fF
C1220 in_14 en14_b 0.00fF
C1221 a_2450_15363# in_20 0.00fF
C1222 a_2454_6442# VPWR 2.95fF
C1223 out a_301_27030# 0.43fF
C1224 a_301_36039# VPWR 3.21fF
C1225 a_2450_33381# en 0.06fF
C1226 in_24 in_25 0.28fF
C1227 en en10_b 0.01fF
C1228 a_2450_16650# a_2450_17937# 0.18fF
C1229 en31_b out 0.66fF
C1230 in_8 en_b 1.24fF
C1231 a_2454_27034# a_301_27030# 7.45fF
C1232 a_301_28317# a_301_25743# 0.03fF
C1233 en30_b a_2454_3868# 0.10fF
C1234 a_301_14160# VPWR 3.21fF
C1235 en24_b out 0.70fF
C1236 a_301_15447# en19_b 0.01fF
C1237 in_29 a_301_3864# 6.75fF
C1238 in_29 a_301_5151# 0.08fF
C1239 a_2454_39904# a_2450_38529# 0.03fF
C1240 en15_b en16_b 0.22fF
C1241 in_22 en 1.38fF
C1242 in_5 in_4 0.28fF
C1243 a_301_20595# VPWR 3.21fF
C1244 a_2454_18025# a_2450_19224# 0.10fF
C1245 a_301_10299# a_2450_8928# 0.01fF
C1246 a_2450_10215# a_2454_10303# 1.92fF
C1247 in_23 a_301_12873# 0.08fF
C1248 a_2454_30895# a_2454_28321# 0.03fF
C1249 a_2450_14076# VPWR 0.55fF
C1250 in_7 a_301_30891# 0.07fF
C1251 in_11 a_301_28317# 0.08fF
C1252 en25_b a_2454_10303# 0.10fF
C1253 a_2454_28321# a_301_28317# 7.45fF
C1254 en3_b en_b 0.05fF
C1255 in_11 in_9 0.03fF
C1256 out a_2454_41191# 7.45fF
C1257 a_301_19308# a_2454_18025# 0.07fF
C1258 en2_b in_2 0.00fF
C1259 a_2454_29608# out 7.60fF
C1260 a_2450_8928# en26_b 0.49fF
C1261 a_301_21882# a_2450_20511# 0.01fF
C1262 a_2450_7641# a_2454_6442# 0.10fF
C1263 in_24 in_22 0.03fF
C1264 a_301_33465# a_301_34752# 0.39fF
C1265 a_301_15447# a_301_12873# 0.03fF
C1266 a_2454_29608# a_2454_27034# 0.03fF
C1267 a_2450_29520# en 0.06fF
C1268 a_2454_10303# VPWR 2.95fF
C1269 a_2454_24460# en13_b 1.80fF
C1270 a_2450_11502# en23_b 0.51fF
C1271 a_301_39900# a_2450_38529# 0.01fF
C1272 en18_b a_2450_19224# 0.49fF
C1273 a_2450_21798# a_2450_20511# 0.18fF
C1274 en_b a_2450_20511# 0.01fF
C1275 a_301_19308# en18_b 0.05fF
C1276 a_2450_11502# a_2454_12877# 0.03fF
C1277 en23_b en_b 0.05fF
C1278 a_2450_12789# a_301_11586# 0.05fF
C1279 en3_b a_301_37326# 1.19fF
C1280 a_2450_2493# a_301_2577# 1.32fF
C1281 a_301_36039# in_4 6.75fF
C1282 en7_b a_2450_30807# 0.01fF
C1283 en5_b out 0.70fF
C1284 a_2450_35955# VPWR 0.55fF
C1285 a_2450_16650# a_301_15447# 0.05fF
C1286 a_2450_41103# a_2454_41191# 1.92fF
C1287 en13_b VPWR 3.16fF
C1288 a_2454_18025# a_2450_17937# 1.92fF
C1289 a_301_5151# VPWR 3.21fF
C1290 out a_2454_27034# 7.60fF
C1291 a_2450_25659# a_301_25743# 1.32fF
C1292 a_301_3864# VPWR 3.21fF
C1293 a_2454_25747# a_301_27030# 0.07fF
C1294 a_2450_26946# en 0.06fF
C1295 a_301_6438# en26_b 0.01fF
C1296 a_301_32178# a_301_30891# 0.39fF
C1297 a_301_9012# a_301_7725# 0.39fF
C1298 in_3 a_2450_37242# 0.00fF
C1299 in_29 a_2450_3780# 0.00fF
C1300 en7_b a_2450_33381# 0.49fF
C1301 en3_b a_2454_38617# 0.10fF
C1302 a_301_16734# a_2450_15363# 0.01fF
C1303 en24_b a_2450_8928# 0.01fF
C1304 en16_b a_2454_20599# 1.80fF
C1305 in_27 en_b 1.24fF
C1306 a_301_33465# en_b 0.58fF
C1307 en a_2450_24372# 0.06fF
C1308 en31_b a_2450_2493# 0.49fF
C1309 en18_b a_2450_17937# 0.51fF
C1310 a_2454_34756# a_2454_32182# 0.03fF
C1311 a_2450_1206# VPWR 0.39fF
C1312 a_301_14160# a_301_12873# 0.39fF
C1313 en a_301_34752# 0.79fF
C1314 a_2450_41103# out 0.76fF
C1315 a_301_24456# en12_b 0.01fF
C1316 en11_b en10_b 0.22fF
C1317 en22_b in_22 0.00fF
C1318 a_2454_20599# en17_b 0.10fF
C1319 a_2454_36043# a_301_34752# 0.08fF
C1320 a_2454_19312# a_2450_20511# 0.10fF
C1321 a_2450_38529# VPWR 0.55fF
C1322 a_2454_37330# en4_b 0.10fF
C1323 a_301_11586# in_23 6.75fF
C1324 a_301_12873# a_2450_14076# 0.05fF
C1325 a_2454_15451# en21_b 0.10fF
C1326 en30_b en_b 0.05fF
C1327 en28_b en29_b 0.22fF
C1328 a_2450_32094# en6_b 0.01fF
C1329 a_2454_37330# a_301_38613# 0.07fF
C1330 in_10 en_b 1.24fF
C1331 in_3 in_5 0.03fF
C1332 en21_b a_2454_12877# 0.03fF
C1333 en15_b a_2454_20599# 0.03fF
C1334 a_2450_35955# in_4 0.00fF
C1335 a_2450_2493# in_30 0.00fF
C1336 en2_b out 0.70fF
C1337 out a_2450_8928# 0.78fF
C1338 en a_301_21882# 0.79fF
C1339 a_2450_11502# a_2454_11590# 1.92fF
C1340 in_23 a_301_10299# 0.07fF
C1341 a_2450_11502# en 0.06fF
C1342 out a_2454_25747# 7.60fF
C1343 in_25 en25_b 0.00fF
C1344 a_2450_3780# VPWR 0.55fF
C1345 a_2454_18025# in_18 0.05fF
C1346 in_12 VPWR 1.24fF
C1347 in_28 in_30 0.03fF
C1348 en a_301_18021# 0.79fF
C1349 a_2450_6354# VPWR 0.55fF
C1350 a_2454_27034# a_2454_25747# 0.37fF
C1351 in_0 en 1.33fF
C1352 out a_2450_2493# 0.78fF
C1353 a_2450_21798# en 0.06fF
C1354 en9_b en 0.01fF
C1355 en en_b 36.55fF
C1356 out a_2450_19224# 0.78fF
C1357 en27_b VPWR 3.16fF
C1358 a_301_9012# in_26 0.08fF
C1359 en0_b a_2454_41191# 1.80fF
C1360 a_2450_33381# a_2454_33469# 1.92fF
C1361 in_25 VPWR 1.24fF
C1362 en1_b en 0.01fF
C1363 a_2450_30807# VPWR 0.55fF
C1364 en30_b a_301_1290# 0.01fF
C1365 in_19 in_20 0.28fF
C1366 out a_301_19308# 0.43fF
C1367 out a_301_32178# 0.43fF
C1368 in_29 a_2454_3868# 0.05fF
C1369 out a_2454_23173# 7.60fF
C1370 a_301_29604# a_2450_28233# 0.01fF
C1371 en18_b in_18 0.00fF
C1372 in_3 a_301_36039# 0.07fF
C1373 in_24 en_b 1.24fF
C1374 a_2450_23085# en 0.06fF
C1375 in_23 in_21 0.03fF
C1376 a_2454_15451# a_2450_15363# 1.92fF
C1377 a_301_27030# a_301_25743# 0.39fF
C1378 a_2450_33381# VPWR 0.55fF
C1379 a_2454_2581# en29_b 0.03fF
C1380 VPWR en10_b 3.16fF
C1381 in_17 en 1.38fF
C1382 a_2450_33381# in_6 0.00fF
C1383 a_2450_26946# en11_b 0.51fF
C1384 out a_301_6438# 0.43fF
C1385 out a_301_23169# 0.43fF
C1386 in_16 a_301_19308# 0.07fF
C1387 a_301_11586# a_301_14160# 0.03fF
C1388 a_301_15447# in_21 0.08fF
C1389 en a_301_37326# 0.79fF
C1390 a_2450_1206# a_2454_1294# 1.88fF
C1391 a_2454_28321# a_301_27030# 0.08fF
C1392 a_2450_7641# a_2450_6354# 0.18fF
C1393 in_11 a_301_27030# 6.75fF
C1394 in_26 a_301_7725# 6.75fF
C1395 a_2454_34756# a_301_33465# 0.08fF
C1396 a_2454_16738# a_301_18021# 0.07fF
C1397 en0_b out 0.58fF
C1398 in_22 VPWR 1.24fF
C1399 a_2454_36043# a_301_37326# 0.07fF
C1400 in_15 a_301_21882# 6.75fF
C1401 en a_301_1290# 0.76fF
C1402 a_2450_7641# en27_b 0.49fF
C1403 out a_2450_17937# 0.78fF
C1404 a_2450_12789# out 0.78fF
C1405 a_2454_6442# en26_b 0.03fF
C1406 in_1 a_301_38613# 0.07fF
C1407 a_301_23169# in_13 0.07fF
C1408 en21_b en 0.01fF
C1409 en13_b a_2450_25659# 0.49fF
C1410 a_2450_32094# en8_b 0.49fF
C1411 en21_b a_2454_14164# 1.80fF
C1412 in_7 a_301_32178# 6.75fF
C1413 a_2450_21798# in_15 0.00fF
C1414 in_15 en_b 1.24fF
C1415 a_2454_36043# a_2454_38617# 0.03fF
C1416 a_301_16734# in_20 0.08fF
C1417 a_301_11586# a_2454_10303# 0.07fF
C1418 a_2450_29520# VPWR 0.55fF
C1419 in_14 in_12 0.03fF
C1420 out a_2450_37242# 0.78fF
C1421 en16_b a_2450_20511# 0.51fF
C1422 a_2454_3868# VPWR 2.95fF
C1423 out en14_b 0.70fF
C1424 a_2454_29608# a_2454_28321# 0.37fF
C1425 en6_b a_2454_32182# 0.03fF
C1426 a_2454_9016# a_301_9012# 7.45fF
C1427 a_2450_11502# en22_b 0.01fF
C1428 a_2450_5067# out 0.78fF
C1429 a_2450_41103# en0_b 0.51fF
C1430 en7_b en_b 0.05fF
C1431 a_2454_30895# a_2450_30807# 1.92fF
C1432 a_2454_5155# en28_b 1.80fF
C1433 a_2454_41191# a_2450_39816# 0.03fF
C1434 en1_b a_2454_39904# 1.80fF
C1435 in_17 in_15 0.03fF
C1436 en22_b en_b 0.05fF
C1437 en17_b a_2450_20511# 0.49fF
C1438 a_2454_5155# en29_b 0.10fF
C1439 out a_301_25743# 0.43fF
C1440 a_2454_23173# a_2454_25747# 0.03fF
C1441 a_2454_10303# a_301_10299# 7.45fF
C1442 a_2454_24460# a_2450_24372# 1.92fF
C1443 a_2450_32094# a_2454_32182# 1.92fF
C1444 en in_31 1.37fF
C1445 a_301_14160# in_21 6.75fF
C1446 a_2454_27034# a_301_25743# 0.08fF
C1447 out a_2454_21886# 7.60fF
C1448 a_301_19308# a_2450_19224# 1.32fF
C1449 a_2450_26946# VPWR 0.55fF
C1450 a_301_16734# in_19 6.75fF
C1451 a_2454_16738# a_2454_19312# 0.03fF
C1452 en_b en11_b 0.05fF
C1453 a_301_28317# en10_b 1.19fF
C1454 out a_2454_28321# 7.60fF
C1455 a_301_34752# a_2454_33469# 0.07fF
C1456 in_21 a_2450_14076# 0.00fF
C1457 out a_301_15447# 0.43fF
C1458 a_2454_9016# a_301_7725# 0.08fF
C1459 a_2454_34756# a_2454_36043# 0.37fF
C1460 en3_b en4_b 0.22fF
C1461 in_0 a_301_41187# 6.75fF
C1462 in_13 a_301_25743# 0.08fF
C1463 in_0 a_301_39900# 0.07fF
C1464 en5_b in_5 0.00fF
C1465 a_2450_15363# en 0.06fF
C1466 a_2454_27034# a_2454_28321# 0.37fF
C1467 en_b a_301_41187# 0.57fF
C1468 en20_b en_b 0.05fF
C1469 in_11 a_2454_27034# 0.05fF
C1470 a_301_39900# en_b 0.58fF
C1471 a_2450_24372# VPWR 0.55fF
C1472 en15_b a_2450_20511# 0.01fF
C1473 in_29 en_b 1.24fF
C1474 en3_b a_301_38613# 0.05fF
C1475 a_2454_37330# en3_b 1.80fF
C1476 en1_b a_301_41187# 0.05fF
C1477 en1_b a_301_39900# 1.19fF
C1478 a_2450_15363# a_2454_14164# 0.10fF
C1479 out a_2450_39816# 0.78fF
C1480 a_301_34752# VPWR 3.21fF
C1481 a_301_29604# en8_b 0.01fF
C1482 in_28 a_301_6438# 0.08fF
C1483 in_11 in_13 0.03fF
C1484 a_301_34752# in_6 0.08fF
C1485 a_301_12873# in_22 6.75fF
C1486 a_301_24456# en 0.79fF
C1487 in_12 a_2450_25659# 0.00fF
C1488 out a_2450_34668# 0.78fF
C1489 en2_b a_2450_37242# 0.01fF
C1490 a_301_23169# a_2454_23173# 7.45fF
C1491 a_2454_39904# a_2454_38617# 0.37fF
C1492 a_2450_17937# a_2450_19224# 0.18fF
C1493 en5_b a_2450_34668# 0.51fF
C1494 a_2450_11502# a_2450_10215# 0.18fF
C1495 en22_b en21_b 0.22fF
C1496 in_16 in_18 0.03fF
C1497 a_2450_29520# a_2454_30895# 0.03fF
C1498 a_301_2577# a_301_3864# 0.39fF
C1499 a_301_2577# a_301_5151# 0.03fF
C1500 a_2450_29520# a_301_28317# 0.05fF
C1501 a_2450_29520# in_9 0.00fF
C1502 a_2454_5155# a_2454_2581# 0.03fF
C1503 a_301_19308# a_2450_17937# 0.01fF
C1504 out a_2454_6442# 7.60fF
C1505 a_301_37326# a_301_39900# 0.03fF
C1506 en24_b a_2454_10303# 1.80fF
C1507 a_2450_10215# en_b 0.01fF
C1508 out a_301_36039# 0.43fF
C1509 a_2454_15451# in_20 0.05fF
C1510 en25_b en_b 0.05fF
C1511 a_301_9012# a_2454_7729# 0.07fF
C1512 in_7 in_5 0.03fF
C1513 en5_b a_301_36039# 0.05fF
C1514 a_301_21882# VPWR 3.21fF
C1515 a_2450_41103# a_2450_39816# 0.18fF
C1516 a_2454_16738# a_2450_15363# 0.03fF
C1517 a_2450_11502# VPWR 0.55fF
C1518 a_2454_3868# a_2454_1294# 0.03fF
C1519 en8_b a_2454_32182# 0.10fF
C1520 a_2454_25747# a_301_25743# 7.45fF
C1521 en20_b en21_b 0.22fF
C1522 a_301_2577# a_2450_1206# 0.01fF
C1523 in_2 a_2450_38529# 0.00fF
C1524 a_301_39900# a_2454_38617# 0.07fF
C1525 en16_b en 0.01fF
C1526 a_301_33465# en6_b 1.19fF
C1527 out a_301_14160# 0.43fF
C1528 VPWR a_301_18021# 3.21fF
C1529 in_0 VPWR 1.40fF
C1530 a_2450_5067# in_28 0.00fF
C1531 en14_b a_2454_23173# 1.80fF
C1532 in_27 a_301_7725# 0.08fF
C1533 a_2450_21798# VPWR 0.55fF
C1534 a_2454_24460# a_2450_23085# 0.03fF
C1535 en9_b VPWR 3.16fF
C1536 in_8 en8_b 0.00fF
C1537 a_301_29604# in_8 0.07fF
C1538 en_b VPWR 63.19fF
C1539 a_301_20595# out 0.43fF
C1540 a_2450_26946# a_301_28317# 0.01fF
C1541 en_b in_6 1.24fF
C1542 a_2454_25747# a_2454_28321# 0.03fF
C1543 in_10 a_2450_28233# 0.00fF
C1544 out a_2450_14076# 0.78fF
C1545 en1_b VPWR 3.16fF
C1546 a_2454_20599# a_2450_20511# 1.92fF
.ends

