VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO sky130_asc_pfet_01v8_lvt_1
  CLASS CORE ;
  FOREIGN sky130_asc_pfet_01v8_lvt_1 ;
  ORIGIN 0.000 0.000 ;
  SIZE 2.940 BY 9.400 ;
  SITE unitasc ;
  PIN GATE
    DIRECTION INOUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 12.900000 ;
    PORT
      LAYER li1 ;
        RECT 0.000 0.520 2.940 0.820 ;
    END
  END GATE
  PIN SOURCE
    DIRECTION INOUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.870500 ;
    PORT
      LAYER li1 ;
        RECT 0.000 8.650 2.940 8.950 ;
        RECT 2.525 8.245 2.695 8.650 ;
        RECT 2.525 8.130 2.700 8.245 ;
        RECT 2.530 1.755 2.700 8.130 ;
      LAYER mcon ;
        RECT 2.530 1.835 2.700 8.165 ;
      LAYER met1 ;
        RECT 2.500 1.775 2.730 8.225 ;
    END
  END SOURCE
  PIN DRAIN
    DIRECTION INOUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.870500 ;
    PORT
      LAYER li1 ;
        RECT 0.240 1.870 0.410 8.245 ;
        RECT 0.235 1.755 0.410 1.870 ;
        RECT 0.235 1.350 0.405 1.755 ;
        RECT 0.000 1.050 2.940 1.350 ;
      LAYER mcon ;
        RECT 0.240 1.835 0.410 8.165 ;
      LAYER met1 ;
        RECT 0.210 1.775 0.440 8.225 ;
    END
  END DRAIN
  PIN VPB
    DIRECTION INPUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT 0.000 1.465 2.940 9.700 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER li1 ;
        RECT 0.000 9.250 2.940 9.550 ;
      LAYER mcon ;
        RECT 0.850 9.250 1.150 9.550 ;
      LAYER met1 ;
        RECT 0.000 9.100 2.940 9.700 ;
    END
  END VPWR
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER li1 ;
        RECT 0.000 -0.150 2.940 0.150 ;
      LAYER mcon ;
        RECT 0.850 -0.150 1.150 0.150 ;
      LAYER met1 ;
        RECT 0.000 -0.300 2.940 0.300 ;
    END
  END VGND
END sky130_asc_pfet_01v8_lvt_1

#--------EOF---------

MACRO sky130_asc_nfet_01v8_lvt_1
  CLASS CORE ;
  FOREIGN sky130_asc_nfet_01v8_lvt_1 ;
  ORIGIN 0.000 0.000 ;
  SIZE 2.580 BY 9.400 ;
  SITE unitasc ;
  PIN VNB
    DIRECTION INPUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.000 0.150 2.580 5.000 ;
        RECT 0.150 -0.150 0.450 0.150 ;
    END
  END VNB
  PIN GATE
    DIRECTION INOUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 8.000000 ;
    PORT
      LAYER li1 ;
        RECT 0.000 0.720 2.580 1.020 ;
    END
  END GATE
  PIN SOURCE
    DIRECTION INOUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.160000 ;
    PORT
      LAYER li1 ;
        RECT 0.000 8.250 2.580 8.550 ;
        RECT 2.345 7.020 2.515 8.250 ;
        RECT 2.345 6.730 2.520 7.020 ;
        RECT 2.350 2.980 2.520 6.730 ;
      LAYER mcon ;
        RECT 2.350 3.060 2.520 6.940 ;
      LAYER met1 ;
        RECT 2.320 3.000 2.550 7.000 ;
    END
  END SOURCE
  PIN DRAIN
    DIRECTION INOUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.160000 ;
    PORT
      LAYER li1 ;
        RECT 0.060 3.270 0.230 7.020 ;
        RECT 0.055 2.980 0.230 3.270 ;
        RECT 0.055 2.520 0.225 2.980 ;
        RECT 0.000 2.220 2.580 2.520 ;
      LAYER mcon ;
        RECT 0.060 3.060 0.230 6.940 ;
      LAYER met1 ;
        RECT 0.030 3.000 0.260 7.000 ;
    END
  END DRAIN
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER li1 ;
        RECT 0.000 9.250 2.580 9.550 ;
      LAYER mcon ;
        RECT 0.850 9.250 1.150 9.550 ;
      LAYER met1 ;
        RECT 0.000 9.100 2.580 9.700 ;
    END
  END VPWR
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER li1 ;
        RECT 0.000 -0.150 2.580 0.150 ;
      LAYER mcon ;
        RECT 0.850 -0.150 1.150 0.150 ;
      LAYER met1 ;
        RECT 0.000 -0.300 2.580 0.300 ;
    END
  END VGND
END sky130_asc_nfet_01v8_lvt_1
END LIBRARY





