** A_MUX_TB flat netlist

V2 VDD GND 1.8
V4 IN0 GND 0.1
V5 IN1 GND 0.2
V6 IN2 GND 0.3
V7 IN3 GND 0.4
R2 OUT32 GND 1E9 M=1
*--------BEGIN_X3->LINE_SWITCHES
*.PININFO IN5:I IN6:I IN7:I IN8:I IN9:I IN10:I IN11:I IN12:I IN13:I IN14:I IN15:I IN16:I IN17:I
*+ IN18:I IN19:I OUT:O IN0:I IN1:I IN2:I IN3:I IN4:I EN0_B:I EN1_B:I EN2_B:I EN3_B:I EN4_B:I EN5_B:I EN6_B:I
*+ EN7_B:I EN8_B:I EN9_B:I EN10_B:I EN11_B:I EN12_B:I EN13_B:I EN14_B:I EN15_B:I EN16_B:I EN17_B:I EN18_B:I
*+ EN19_B:I EN20_B:I EN21_B:I EN22_B:I EN23_B:I EN24_B:I EN25_B:I EN26_B:I EN27_B:I EN28_B:I EN29_B:I EN30_B:I
*+ EN31_B:I EN_B:I EN:I
*--------BEGIN_X3_X28->TRANSMISSION_GATE
*.PININFO IN:B OUT:B EN:I EN_B:I
*--------BEGIN_X3_X28_XM1->W'
XM1_X3_X28 X3_NET1 VDD IN10 X3_VSS X3_X28_SKY130_FD_PR__NFET_01V8 X3_X28_* X3_X28_W/NF X3_X28_* X3_X28_0.29'
+ X3_X28_* X3_X28_W/NF X3_X28_* X3_X28_0.29' X3_X28_* X3_X28_(W/NF X3_X28_+ X3_X28_0.29)' X3_X28_* X3_X28_(W/NF
+ X3_X28_+ X3_X28_0.29)' X3_X28_/ X3_X28_W' X3_X28_/  W' L='L_N' W='W_N' NF=1 AD='INT((NF+1)/2) AS='INT((NF+2)/2) PD='2*INT((NF+1)/2)
+ PS='2*INT((NF+2)/2) NRD='0.29 NRS='0.29 SA=0 SB=0 SD=0 MULT='N' M='N' 
*--------END___X3_X28_XM1->W'
*--------BEGIN_X3_X28_XM2->W'
XM2_X3_X28 X3_NET1 GND IN10 VDD X3_X28_SKY130_FD_PR__PFET_01V8 X3_X28_* X3_X28_W/NF X3_X28_* X3_X28_0.29'
+ X3_X28_* X3_X28_W/NF X3_X28_* X3_X28_0.29' X3_X28_* X3_X28_(W/NF X3_X28_+ X3_X28_0.29)' X3_X28_* X3_X28_(W/NF
+ X3_X28_+ X3_X28_0.29)' X3_X28_/ X3_X28_W' X3_X28_/  W' L='L_P' W='W_P' NF=1 AD='INT((NF+1)/2) AS='INT((NF+2)/2) PD='2*INT((NF+1)/2)
+ PS='2*INT((NF+2)/2) NRD='0.29 NRS='0.29 SA=0 SB=0 SD=0 MULT='N' M='N' 
*--------END___X3_X28_XM2->W'
*--------END___X3_X28->TRANSMISSION_GATE
*--------BEGIN_X3_X29->SWITCH_5T
*.PININFO IN:B OUT:B EN:I EN_B:I
*--------BEGIN_X3_X29_X1->TRANSMISSION_GATE
*.PININFO IN:B OUT:B EN:I EN_B:I
*--------BEGIN_X3_X29_X1_XM1->W'
XM1_X3_X29_X1 X3_X29_NET1 X3_NET21 X3_NET1 X3_VSS X3_X29_X1_SKY130_FD_PR__NFET_01V8 X3_X29_X1_* X3_X29_X1_W/NF X3_X29_X1_* X3_X29_X1_0.29'
+ X3_X29_X1_* X3_X29_X1_W/NF X3_X29_X1_* X3_X29_X1_0.29' X3_X29_X1_* X3_X29_X1_(W/NF X3_X29_X1_+ X3_X29_X1_0.29)'
+ X3_X29_X1_* X3_X29_X1_(W/NF X3_X29_X1_+ X3_X29_X1_0.29)' X3_X29_X1_/ X3_X29_X1_W' X3_X29_X1_/  W' L='L_N' W='W_N' NF=1 AD='INT((NF+1)/2)
+ AS='INT((NF+2)/2) PD='2*INT((NF+1)/2) PS='2*INT((NF+2)/2) NRD='0.29 NRS='0.29 SA=0 SB=0 SD=0 MULT='N' M='N' 
*--------END___X3_X29_X1_XM1->W'
*--------BEGIN_X3_X29_X1_XM2->W'
XM2_X3_X29_X1 X3_X29_NET1 VDD X3_NET1 VDD X3_X29_X1_SKY130_FD_PR__PFET_01V8 X3_X29_X1_* X3_X29_X1_W/NF X3_X29_X1_* X3_X29_X1_0.29'
+ X3_X29_X1_* X3_X29_X1_W/NF X3_X29_X1_* X3_X29_X1_0.29' X3_X29_X1_* X3_X29_X1_(W/NF X3_X29_X1_+ X3_X29_X1_0.29)'
+ X3_X29_X1_* X3_X29_X1_(W/NF X3_X29_X1_+ X3_X29_X1_0.29)' X3_X29_X1_/ X3_X29_X1_W' X3_X29_X1_/  W' L='L_P' W='W_P' NF=1 AD='INT((NF+1)/2)
+ AS='INT((NF+2)/2) PD='2*INT((NF+1)/2) PS='2*INT((NF+2)/2) NRD='0.29 NRS='0.29 SA=0 SB=0 SD=0 MULT='N' M='N' 
*--------END___X3_X29_X1_XM2->W'
*--------END___X3_X29_X1->TRANSMISSION_GATE
*--------BEGIN_X3_X29_X2->TRANSMISSION_GATE
*.PININFO IN:B OUT:B EN:I EN_B:I
*--------BEGIN_X3_X29_X2_XM1->W'
XM1_X3_X29_X2 OUT32 X3_NET21 X3_X29_NET1 X3_VSS X3_X29_X2_SKY130_FD_PR__NFET_01V8 X3_X29_X2_* X3_X29_X2_W/NF X3_X29_X2_* X3_X29_X2_0.29'
+ X3_X29_X2_* X3_X29_X2_W/NF X3_X29_X2_* X3_X29_X2_0.29' X3_X29_X2_* X3_X29_X2_(W/NF X3_X29_X2_+ X3_X29_X2_0.29)'
+ X3_X29_X2_* X3_X29_X2_(W/NF X3_X29_X2_+ X3_X29_X2_0.29)' X3_X29_X2_/ X3_X29_X2_W' X3_X29_X2_/  W' L='L_N' W='W_N' NF=1 AD='INT((NF+1)/2)
+ AS='INT((NF+2)/2) PD='2*INT((NF+1)/2) PS='2*INT((NF+2)/2) NRD='0.29 NRS='0.29 SA=0 SB=0 SD=0 MULT='N' M='N' 
*--------END___X3_X29_X2_XM1->W'
*--------BEGIN_X3_X29_X2_XM2->W'
XM2_X3_X29_X2 OUT32 VDD X3_X29_NET1 VDD X3_X29_X2_SKY130_FD_PR__PFET_01V8 X3_X29_X2_* X3_X29_X2_W/NF X3_X29_X2_* X3_X29_X2_0.29'
+ X3_X29_X2_* X3_X29_X2_W/NF X3_X29_X2_* X3_X29_X2_0.29' X3_X29_X2_* X3_X29_X2_(W/NF X3_X29_X2_+ X3_X29_X2_0.29)'
+ X3_X29_X2_* X3_X29_X2_(W/NF X3_X29_X2_+ X3_X29_X2_0.29)' X3_X29_X2_/ X3_X29_X2_W' X3_X29_X2_/  W' L='L_P' W='W_P' NF=1 AD='INT((NF+1)/2)
+ AS='INT((NF+2)/2) PD='2*INT((NF+1)/2) PS='2*INT((NF+2)/2) NRD='0.29 NRS='0.29 SA=0 SB=0 SD=0 MULT='N' M='N' 
*--------END___X3_X29_X2_XM2->W'
*--------END___X3_X29_X2->TRANSMISSION_GATE
*--------BEGIN_X3_X29_XM1->W'
XM1_X3_X29 X3_X29_NET1 VDD X3_VSS X3_VSS X3_X29_SKY130_FD_PR__NFET_01V8 X3_X29_* X3_X29_W/NF X3_X29_* X3_X29_0.29'
+ X3_X29_* X3_X29_W/NF X3_X29_* X3_X29_0.29' X3_X29_* X3_X29_(W/NF X3_X29_+ X3_X29_0.29)' X3_X29_* X3_X29_(W/NF
+ X3_X29_+ X3_X29_0.29)' X3_X29_/ X3_X29_W' X3_X29_/  W' L=0.15 W=0.5 NF=1 AD='INT((NF+1)/2) AS='INT((NF+2)/2) PD='2*INT((NF+1)/2)
+ PS='2*INT((NF+2)/2) NRD='0.29 NRS='0.29 SA=0 SB=0 SD=0 MULT=1 M=1 
*--------END___X3_X29_XM1->W'
*--------END___X3_X29->SWITCH_5T
*--------BEGIN_X3_X30->SKY130_FD_SC_HD__INV_1
X30_X3 VDD X3_VGND X3_VNB X3_VPB X3_VPWR X3_NET21  SKY130_FD_SC_HD__INV_1
*--------END___X3_X30->SKY130_FD_SC_HD__INV_1
*--------BEGIN_X3_X31->TRANSMISSION_GATE
*.PININFO IN:B OUT:B EN:I EN_B:I
*--------BEGIN_X3_X31_XM1->W'
XM1_X3_X31 X3_NET2 VDD IN11 X3_VSS X3_X31_SKY130_FD_PR__NFET_01V8 X3_X31_* X3_X31_W/NF X3_X31_* X3_X31_0.29'
+ X3_X31_* X3_X31_W/NF X3_X31_* X3_X31_0.29' X3_X31_* X3_X31_(W/NF X3_X31_+ X3_X31_0.29)' X3_X31_* X3_X31_(W/NF
+ X3_X31_+ X3_X31_0.29)' X3_X31_/ X3_X31_W' X3_X31_/  W' L='L_N' W='W_N' NF=1 AD='INT((NF+1)/2) AS='INT((NF+2)/2) PD='2*INT((NF+1)/2)
+ PS='2*INT((NF+2)/2) NRD='0.29 NRS='0.29 SA=0 SB=0 SD=0 MULT='N' M='N' 
*--------END___X3_X31_XM1->W'
*--------BEGIN_X3_X31_XM2->W'
XM2_X3_X31 X3_NET2 GND IN11 VDD X3_X31_SKY130_FD_PR__PFET_01V8 X3_X31_* X3_X31_W/NF X3_X31_* X3_X31_0.29'
+ X3_X31_* X3_X31_W/NF X3_X31_* X3_X31_0.29' X3_X31_* X3_X31_(W/NF X3_X31_+ X3_X31_0.29)' X3_X31_* X3_X31_(W/NF
+ X3_X31_+ X3_X31_0.29)' X3_X31_/ X3_X31_W' X3_X31_/  W' L='L_P' W='W_P' NF=1 AD='INT((NF+1)/2) AS='INT((NF+2)/2) PD='2*INT((NF+1)/2)
+ PS='2*INT((NF+2)/2) NRD='0.29 NRS='0.29 SA=0 SB=0 SD=0 MULT='N' M='N' 
*--------END___X3_X31_XM2->W'
*--------END___X3_X31->TRANSMISSION_GATE
*--------BEGIN_X3_X32->SWITCH_5T
*.PININFO IN:B OUT:B EN:I EN_B:I
*--------BEGIN_X3_X32_X1->TRANSMISSION_GATE
*.PININFO IN:B OUT:B EN:I EN_B:I
*--------BEGIN_X3_X32_X1_XM1->W'
XM1_X3_X32_X1 X3_X32_NET1 X3_NET22 X3_NET2 X3_VSS X3_X32_X1_SKY130_FD_PR__NFET_01V8 X3_X32_X1_* X3_X32_X1_W/NF X3_X32_X1_* X3_X32_X1_0.29'
+ X3_X32_X1_* X3_X32_X1_W/NF X3_X32_X1_* X3_X32_X1_0.29' X3_X32_X1_* X3_X32_X1_(W/NF X3_X32_X1_+ X3_X32_X1_0.29)'
+ X3_X32_X1_* X3_X32_X1_(W/NF X3_X32_X1_+ X3_X32_X1_0.29)' X3_X32_X1_/ X3_X32_X1_W' X3_X32_X1_/  W' L='L_N' W='W_N' NF=1 AD='INT((NF+1)/2)
+ AS='INT((NF+2)/2) PD='2*INT((NF+1)/2) PS='2*INT((NF+2)/2) NRD='0.29 NRS='0.29 SA=0 SB=0 SD=0 MULT='N' M='N' 
*--------END___X3_X32_X1_XM1->W'
*--------BEGIN_X3_X32_X1_XM2->W'
XM2_X3_X32_X1 X3_X32_NET1 VDD X3_NET2 VDD X3_X32_X1_SKY130_FD_PR__PFET_01V8 X3_X32_X1_* X3_X32_X1_W/NF X3_X32_X1_* X3_X32_X1_0.29'
+ X3_X32_X1_* X3_X32_X1_W/NF X3_X32_X1_* X3_X32_X1_0.29' X3_X32_X1_* X3_X32_X1_(W/NF X3_X32_X1_+ X3_X32_X1_0.29)'
+ X3_X32_X1_* X3_X32_X1_(W/NF X3_X32_X1_+ X3_X32_X1_0.29)' X3_X32_X1_/ X3_X32_X1_W' X3_X32_X1_/  W' L='L_P' W='W_P' NF=1 AD='INT((NF+1)/2)
+ AS='INT((NF+2)/2) PD='2*INT((NF+1)/2) PS='2*INT((NF+2)/2) NRD='0.29 NRS='0.29 SA=0 SB=0 SD=0 MULT='N' M='N' 
*--------END___X3_X32_X1_XM2->W'
*--------END___X3_X32_X1->TRANSMISSION_GATE
*--------BEGIN_X3_X32_X2->TRANSMISSION_GATE
*.PININFO IN:B OUT:B EN:I EN_B:I
*--------BEGIN_X3_X32_X2_XM1->W'
XM1_X3_X32_X2 OUT32 X3_NET22 X3_X32_NET1 X3_VSS X3_X32_X2_SKY130_FD_PR__NFET_01V8 X3_X32_X2_* X3_X32_X2_W/NF X3_X32_X2_* X3_X32_X2_0.29'
+ X3_X32_X2_* X3_X32_X2_W/NF X3_X32_X2_* X3_X32_X2_0.29' X3_X32_X2_* X3_X32_X2_(W/NF X3_X32_X2_+ X3_X32_X2_0.29)'
+ X3_X32_X2_* X3_X32_X2_(W/NF X3_X32_X2_+ X3_X32_X2_0.29)' X3_X32_X2_/ X3_X32_X2_W' X3_X32_X2_/  W' L='L_N' W='W_N' NF=1 AD='INT((NF+1)/2)
+ AS='INT((NF+2)/2) PD='2*INT((NF+1)/2) PS='2*INT((NF+2)/2) NRD='0.29 NRS='0.29 SA=0 SB=0 SD=0 MULT='N' M='N' 
*--------END___X3_X32_X2_XM1->W'
*--------BEGIN_X3_X32_X2_XM2->W'
XM2_X3_X32_X2 OUT32 VDD X3_X32_NET1 VDD X3_X32_X2_SKY130_FD_PR__PFET_01V8 X3_X32_X2_* X3_X32_X2_W/NF X3_X32_X2_* X3_X32_X2_0.29'
+ X3_X32_X2_* X3_X32_X2_W/NF X3_X32_X2_* X3_X32_X2_0.29' X3_X32_X2_* X3_X32_X2_(W/NF X3_X32_X2_+ X3_X32_X2_0.29)'
+ X3_X32_X2_* X3_X32_X2_(W/NF X3_X32_X2_+ X3_X32_X2_0.29)' X3_X32_X2_/ X3_X32_X2_W' X3_X32_X2_/  W' L='L_P' W='W_P' NF=1 AD='INT((NF+1)/2)
+ AS='INT((NF+2)/2) PD='2*INT((NF+1)/2) PS='2*INT((NF+2)/2) NRD='0.29 NRS='0.29 SA=0 SB=0 SD=0 MULT='N' M='N' 
*--------END___X3_X32_X2_XM2->W'
*--------END___X3_X32_X2->TRANSMISSION_GATE
*--------BEGIN_X3_X32_XM1->W'
XM1_X3_X32 X3_X32_NET1 VDD X3_VSS X3_VSS X3_X32_SKY130_FD_PR__NFET_01V8 X3_X32_* X3_X32_W/NF X3_X32_* X3_X32_0.29'
+ X3_X32_* X3_X32_W/NF X3_X32_* X3_X32_0.29' X3_X32_* X3_X32_(W/NF X3_X32_+ X3_X32_0.29)' X3_X32_* X3_X32_(W/NF
+ X3_X32_+ X3_X32_0.29)' X3_X32_/ X3_X32_W' X3_X32_/  W' L=0.15 W=0.5 NF=1 AD='INT((NF+1)/2) AS='INT((NF+2)/2) PD='2*INT((NF+1)/2)
+ PS='2*INT((NF+2)/2) NRD='0.29 NRS='0.29 SA=0 SB=0 SD=0 MULT=1 M=1 
*--------END___X3_X32_XM1->W'
*--------END___X3_X32->SWITCH_5T
*--------BEGIN_X3_X33->SKY130_FD_SC_HD__INV_1
X33_X3 VDD X3_VGND X3_VNB X3_VPB X3_VPWR X3_NET22  SKY130_FD_SC_HD__INV_1
*--------END___X3_X33->SKY130_FD_SC_HD__INV_1
*--------BEGIN_X3_X34->TRANSMISSION_GATE
*.PININFO IN:B OUT:B EN:I EN_B:I
*--------BEGIN_X3_X34_XM1->W'
XM1_X3_X34 X3_NET3 VDD IN12 X3_VSS X3_X34_SKY130_FD_PR__NFET_01V8 X3_X34_* X3_X34_W/NF X3_X34_* X3_X34_0.29'
+ X3_X34_* X3_X34_W/NF X3_X34_* X3_X34_0.29' X3_X34_* X3_X34_(W/NF X3_X34_+ X3_X34_0.29)' X3_X34_* X3_X34_(W/NF
+ X3_X34_+ X3_X34_0.29)' X3_X34_/ X3_X34_W' X3_X34_/  W' L='L_N' W='W_N' NF=1 AD='INT((NF+1)/2) AS='INT((NF+2)/2) PD='2*INT((NF+1)/2)
+ PS='2*INT((NF+2)/2) NRD='0.29 NRS='0.29 SA=0 SB=0 SD=0 MULT='N' M='N' 
*--------END___X3_X34_XM1->W'
*--------BEGIN_X3_X34_XM2->W'
XM2_X3_X34 X3_NET3 GND IN12 VDD X3_X34_SKY130_FD_PR__PFET_01V8 X3_X34_* X3_X34_W/NF X3_X34_* X3_X34_0.29'
+ X3_X34_* X3_X34_W/NF X3_X34_* X3_X34_0.29' X3_X34_* X3_X34_(W/NF X3_X34_+ X3_X34_0.29)' X3_X34_* X3_X34_(W/NF
+ X3_X34_+ X3_X34_0.29)' X3_X34_/ X3_X34_W' X3_X34_/  W' L='L_P' W='W_P' NF=1 AD='INT((NF+1)/2) AS='INT((NF+2)/2) PD='2*INT((NF+1)/2)
+ PS='2*INT((NF+2)/2) NRD='0.29 NRS='0.29 SA=0 SB=0 SD=0 MULT='N' M='N' 
*--------END___X3_X34_XM2->W'
*--------END___X3_X34->TRANSMISSION_GATE
*--------BEGIN_X3_X35->SWITCH_5T
*.PININFO IN:B OUT:B EN:I EN_B:I
*--------BEGIN_X3_X35_X1->TRANSMISSION_GATE
*.PININFO IN:B OUT:B EN:I EN_B:I
*--------BEGIN_X3_X35_X1_XM1->W'
XM1_X3_X35_X1 X3_X35_NET1 X3_NET23 X3_NET3 X3_VSS X3_X35_X1_SKY130_FD_PR__NFET_01V8 X3_X35_X1_* X3_X35_X1_W/NF X3_X35_X1_* X3_X35_X1_0.29'
+ X3_X35_X1_* X3_X35_X1_W/NF X3_X35_X1_* X3_X35_X1_0.29' X3_X35_X1_* X3_X35_X1_(W/NF X3_X35_X1_+ X3_X35_X1_0.29)'
+ X3_X35_X1_* X3_X35_X1_(W/NF X3_X35_X1_+ X3_X35_X1_0.29)' X3_X35_X1_/ X3_X35_X1_W' X3_X35_X1_/  W' L='L_N' W='W_N' NF=1 AD='INT((NF+1)/2)
+ AS='INT((NF+2)/2) PD='2*INT((NF+1)/2) PS='2*INT((NF+2)/2) NRD='0.29 NRS='0.29 SA=0 SB=0 SD=0 MULT='N' M='N' 
*--------END___X3_X35_X1_XM1->W'
*--------BEGIN_X3_X35_X1_XM2->W'
XM2_X3_X35_X1 X3_X35_NET1 VDD X3_NET3 VDD X3_X35_X1_SKY130_FD_PR__PFET_01V8 X3_X35_X1_* X3_X35_X1_W/NF X3_X35_X1_* X3_X35_X1_0.29'
+ X3_X35_X1_* X3_X35_X1_W/NF X3_X35_X1_* X3_X35_X1_0.29' X3_X35_X1_* X3_X35_X1_(W/NF X3_X35_X1_+ X3_X35_X1_0.29)'
+ X3_X35_X1_* X3_X35_X1_(W/NF X3_X35_X1_+ X3_X35_X1_0.29)' X3_X35_X1_/ X3_X35_X1_W' X3_X35_X1_/  W' L='L_P' W='W_P' NF=1 AD='INT((NF+1)/2)
+ AS='INT((NF+2)/2) PD='2*INT((NF+1)/2) PS='2*INT((NF+2)/2) NRD='0.29 NRS='0.29 SA=0 SB=0 SD=0 MULT='N' M='N' 
*--------END___X3_X35_X1_XM2->W'
*--------END___X3_X35_X1->TRANSMISSION_GATE
*--------BEGIN_X3_X35_X2->TRANSMISSION_GATE
*.PININFO IN:B OUT:B EN:I EN_B:I
*--------BEGIN_X3_X35_X2_XM1->W'
XM1_X3_X35_X2 OUT32 X3_NET23 X3_X35_NET1 X3_VSS X3_X35_X2_SKY130_FD_PR__NFET_01V8 X3_X35_X2_* X3_X35_X2_W/NF X3_X35_X2_* X3_X35_X2_0.29'
+ X3_X35_X2_* X3_X35_X2_W/NF X3_X35_X2_* X3_X35_X2_0.29' X3_X35_X2_* X3_X35_X2_(W/NF X3_X35_X2_+ X3_X35_X2_0.29)'
+ X3_X35_X2_* X3_X35_X2_(W/NF X3_X35_X2_+ X3_X35_X2_0.29)' X3_X35_X2_/ X3_X35_X2_W' X3_X35_X2_/  W' L='L_N' W='W_N' NF=1 AD='INT((NF+1)/2)
+ AS='INT((NF+2)/2) PD='2*INT((NF+1)/2) PS='2*INT((NF+2)/2) NRD='0.29 NRS='0.29 SA=0 SB=0 SD=0 MULT='N' M='N' 
*--------END___X3_X35_X2_XM1->W'
*--------BEGIN_X3_X35_X2_XM2->W'
XM2_X3_X35_X2 OUT32 VDD X3_X35_NET1 VDD X3_X35_X2_SKY130_FD_PR__PFET_01V8 X3_X35_X2_* X3_X35_X2_W/NF X3_X35_X2_* X3_X35_X2_0.29'
+ X3_X35_X2_* X3_X35_X2_W/NF X3_X35_X2_* X3_X35_X2_0.29' X3_X35_X2_* X3_X35_X2_(W/NF X3_X35_X2_+ X3_X35_X2_0.29)'
+ X3_X35_X2_* X3_X35_X2_(W/NF X3_X35_X2_+ X3_X35_X2_0.29)' X3_X35_X2_/ X3_X35_X2_W' X3_X35_X2_/  W' L='L_P' W='W_P' NF=1 AD='INT((NF+1)/2)
+ AS='INT((NF+2)/2) PD='2*INT((NF+1)/2) PS='2*INT((NF+2)/2) NRD='0.29 NRS='0.29 SA=0 SB=0 SD=0 MULT='N' M='N' 
*--------END___X3_X35_X2_XM2->W'
*--------END___X3_X35_X2->TRANSMISSION_GATE
*--------BEGIN_X3_X35_XM1->W'
XM1_X3_X35 X3_X35_NET1 VDD X3_VSS X3_VSS X3_X35_SKY130_FD_PR__NFET_01V8 X3_X35_* X3_X35_W/NF X3_X35_* X3_X35_0.29'
+ X3_X35_* X3_X35_W/NF X3_X35_* X3_X35_0.29' X3_X35_* X3_X35_(W/NF X3_X35_+ X3_X35_0.29)' X3_X35_* X3_X35_(W/NF
+ X3_X35_+ X3_X35_0.29)' X3_X35_/ X3_X35_W' X3_X35_/  W' L=0.15 W=0.5 NF=1 AD='INT((NF+1)/2) AS='INT((NF+2)/2) PD='2*INT((NF+1)/2)
+ PS='2*INT((NF+2)/2) NRD='0.29 NRS='0.29 SA=0 SB=0 SD=0 MULT=1 M=1 
*--------END___X3_X35_XM1->W'
*--------END___X3_X35->SWITCH_5T
*--------BEGIN_X3_X36->SKY130_FD_SC_HD__INV_1
X36_X3 VDD X3_VGND X3_VNB X3_VPB X3_VPWR X3_NET23  SKY130_FD_SC_HD__INV_1
*--------END___X3_X36->SKY130_FD_SC_HD__INV_1
*--------BEGIN_X3_X37->TRANSMISSION_GATE
*.PININFO IN:B OUT:B EN:I EN_B:I
*--------BEGIN_X3_X37_XM1->W'
XM1_X3_X37 X3_NET4 VDD IN13 X3_VSS X3_X37_SKY130_FD_PR__NFET_01V8 X3_X37_* X3_X37_W/NF X3_X37_* X3_X37_0.29'
+ X3_X37_* X3_X37_W/NF X3_X37_* X3_X37_0.29' X3_X37_* X3_X37_(W/NF X3_X37_+ X3_X37_0.29)' X3_X37_* X3_X37_(W/NF
+ X3_X37_+ X3_X37_0.29)' X3_X37_/ X3_X37_W' X3_X37_/  W' L='L_N' W='W_N' NF=1 AD='INT((NF+1)/2) AS='INT((NF+2)/2) PD='2*INT((NF+1)/2)
+ PS='2*INT((NF+2)/2) NRD='0.29 NRS='0.29 SA=0 SB=0 SD=0 MULT='N' M='N' 
*--------END___X3_X37_XM1->W'
*--------BEGIN_X3_X37_XM2->W'
XM2_X3_X37 X3_NET4 GND IN13 VDD X3_X37_SKY130_FD_PR__PFET_01V8 X3_X37_* X3_X37_W/NF X3_X37_* X3_X37_0.29'
+ X3_X37_* X3_X37_W/NF X3_X37_* X3_X37_0.29' X3_X37_* X3_X37_(W/NF X3_X37_+ X3_X37_0.29)' X3_X37_* X3_X37_(W/NF
+ X3_X37_+ X3_X37_0.29)' X3_X37_/ X3_X37_W' X3_X37_/  W' L='L_P' W='W_P' NF=1 AD='INT((NF+1)/2) AS='INT((NF+2)/2) PD='2*INT((NF+1)/2)
+ PS='2*INT((NF+2)/2) NRD='0.29 NRS='0.29 SA=0 SB=0 SD=0 MULT='N' M='N' 
*--------END___X3_X37_XM2->W'
*--------END___X3_X37->TRANSMISSION_GATE
*--------BEGIN_X3_X38->SWITCH_5T
*.PININFO IN:B OUT:B EN:I EN_B:I
*--------BEGIN_X3_X38_X1->TRANSMISSION_GATE
*.PININFO IN:B OUT:B EN:I EN_B:I
*--------BEGIN_X3_X38_X1_XM1->W'
XM1_X3_X38_X1 X3_X38_NET1 X3_NET24 X3_NET4 X3_VSS X3_X38_X1_SKY130_FD_PR__NFET_01V8 X3_X38_X1_* X3_X38_X1_W/NF X3_X38_X1_* X3_X38_X1_0.29'
+ X3_X38_X1_* X3_X38_X1_W/NF X3_X38_X1_* X3_X38_X1_0.29' X3_X38_X1_* X3_X38_X1_(W/NF X3_X38_X1_+ X3_X38_X1_0.29)'
+ X3_X38_X1_* X3_X38_X1_(W/NF X3_X38_X1_+ X3_X38_X1_0.29)' X3_X38_X1_/ X3_X38_X1_W' X3_X38_X1_/  W' L='L_N' W='W_N' NF=1 AD='INT((NF+1)/2)
+ AS='INT((NF+2)/2) PD='2*INT((NF+1)/2) PS='2*INT((NF+2)/2) NRD='0.29 NRS='0.29 SA=0 SB=0 SD=0 MULT='N' M='N' 
*--------END___X3_X38_X1_XM1->W'
*--------BEGIN_X3_X38_X1_XM2->W'
XM2_X3_X38_X1 X3_X38_NET1 VDD X3_NET4 VDD X3_X38_X1_SKY130_FD_PR__PFET_01V8 X3_X38_X1_* X3_X38_X1_W/NF X3_X38_X1_* X3_X38_X1_0.29'
+ X3_X38_X1_* X3_X38_X1_W/NF X3_X38_X1_* X3_X38_X1_0.29' X3_X38_X1_* X3_X38_X1_(W/NF X3_X38_X1_+ X3_X38_X1_0.29)'
+ X3_X38_X1_* X3_X38_X1_(W/NF X3_X38_X1_+ X3_X38_X1_0.29)' X3_X38_X1_/ X3_X38_X1_W' X3_X38_X1_/  W' L='L_P' W='W_P' NF=1 AD='INT((NF+1)/2)
+ AS='INT((NF+2)/2) PD='2*INT((NF+1)/2) PS='2*INT((NF+2)/2) NRD='0.29 NRS='0.29 SA=0 SB=0 SD=0 MULT='N' M='N' 
*--------END___X3_X38_X1_XM2->W'
*--------END___X3_X38_X1->TRANSMISSION_GATE
*--------BEGIN_X3_X38_X2->TRANSMISSION_GATE
*.PININFO IN:B OUT:B EN:I EN_B:I
*--------BEGIN_X3_X38_X2_XM1->W'
XM1_X3_X38_X2 OUT32 X3_NET24 X3_X38_NET1 X3_VSS X3_X38_X2_SKY130_FD_PR__NFET_01V8 X3_X38_X2_* X3_X38_X2_W/NF X3_X38_X2_* X3_X38_X2_0.29'
+ X3_X38_X2_* X3_X38_X2_W/NF X3_X38_X2_* X3_X38_X2_0.29' X3_X38_X2_* X3_X38_X2_(W/NF X3_X38_X2_+ X3_X38_X2_0.29)'
+ X3_X38_X2_* X3_X38_X2_(W/NF X3_X38_X2_+ X3_X38_X2_0.29)' X3_X38_X2_/ X3_X38_X2_W' X3_X38_X2_/  W' L='L_N' W='W_N' NF=1 AD='INT((NF+1)/2)
+ AS='INT((NF+2)/2) PD='2*INT((NF+1)/2) PS='2*INT((NF+2)/2) NRD='0.29 NRS='0.29 SA=0 SB=0 SD=0 MULT='N' M='N' 
*--------END___X3_X38_X2_XM1->W'
*--------BEGIN_X3_X38_X2_XM2->W'
XM2_X3_X38_X2 OUT32 VDD X3_X38_NET1 VDD X3_X38_X2_SKY130_FD_PR__PFET_01V8 X3_X38_X2_* X3_X38_X2_W/NF X3_X38_X2_* X3_X38_X2_0.29'
+ X3_X38_X2_* X3_X38_X2_W/NF X3_X38_X2_* X3_X38_X2_0.29' X3_X38_X2_* X3_X38_X2_(W/NF X3_X38_X2_+ X3_X38_X2_0.29)'
+ X3_X38_X2_* X3_X38_X2_(W/NF X3_X38_X2_+ X3_X38_X2_0.29)' X3_X38_X2_/ X3_X38_X2_W' X3_X38_X2_/  W' L='L_P' W='W_P' NF=1 AD='INT((NF+1)/2)
+ AS='INT((NF+2)/2) PD='2*INT((NF+1)/2) PS='2*INT((NF+2)/2) NRD='0.29 NRS='0.29 SA=0 SB=0 SD=0 MULT='N' M='N' 
*--------END___X3_X38_X2_XM2->W'
*--------END___X3_X38_X2->TRANSMISSION_GATE
*--------BEGIN_X3_X38_XM1->W'
XM1_X3_X38 X3_X38_NET1 VDD X3_VSS X3_VSS X3_X38_SKY130_FD_PR__NFET_01V8 X3_X38_* X3_X38_W/NF X3_X38_* X3_X38_0.29'
+ X3_X38_* X3_X38_W/NF X3_X38_* X3_X38_0.29' X3_X38_* X3_X38_(W/NF X3_X38_+ X3_X38_0.29)' X3_X38_* X3_X38_(W/NF
+ X3_X38_+ X3_X38_0.29)' X3_X38_/ X3_X38_W' X3_X38_/  W' L=0.15 W=0.5 NF=1 AD='INT((NF+1)/2) AS='INT((NF+2)/2) PD='2*INT((NF+1)/2)
+ PS='2*INT((NF+2)/2) NRD='0.29 NRS='0.29 SA=0 SB=0 SD=0 MULT=1 M=1 
*--------END___X3_X38_XM1->W'
*--------END___X3_X38->SWITCH_5T
*--------BEGIN_X3_X39->SKY130_FD_SC_HD__INV_1
X39_X3 VDD X3_VGND X3_VNB X3_VPB X3_VPWR X3_NET24  SKY130_FD_SC_HD__INV_1
*--------END___X3_X39->SKY130_FD_SC_HD__INV_1
*--------BEGIN_X3_X40->TRANSMISSION_GATE
*.PININFO IN:B OUT:B EN:I EN_B:I
*--------BEGIN_X3_X40_XM1->W'
XM1_X3_X40 X3_NET5 VDD IN14 X3_VSS X3_X40_SKY130_FD_PR__NFET_01V8 X3_X40_* X3_X40_W/NF X3_X40_* X3_X40_0.29'
+ X3_X40_* X3_X40_W/NF X3_X40_* X3_X40_0.29' X3_X40_* X3_X40_(W/NF X3_X40_+ X3_X40_0.29)' X3_X40_* X3_X40_(W/NF
+ X3_X40_+ X3_X40_0.29)' X3_X40_/ X3_X40_W' X3_X40_/  W' L='L_N' W='W_N' NF=1 AD='INT((NF+1)/2) AS='INT((NF+2)/2) PD='2*INT((NF+1)/2)
+ PS='2*INT((NF+2)/2) NRD='0.29 NRS='0.29 SA=0 SB=0 SD=0 MULT='N' M='N' 
*--------END___X3_X40_XM1->W'
*--------BEGIN_X3_X40_XM2->W'
XM2_X3_X40 X3_NET5 GND IN14 VDD X3_X40_SKY130_FD_PR__PFET_01V8 X3_X40_* X3_X40_W/NF X3_X40_* X3_X40_0.29'
+ X3_X40_* X3_X40_W/NF X3_X40_* X3_X40_0.29' X3_X40_* X3_X40_(W/NF X3_X40_+ X3_X40_0.29)' X3_X40_* X3_X40_(W/NF
+ X3_X40_+ X3_X40_0.29)' X3_X40_/ X3_X40_W' X3_X40_/  W' L='L_P' W='W_P' NF=1 AD='INT((NF+1)/2) AS='INT((NF+2)/2) PD='2*INT((NF+1)/2)
+ PS='2*INT((NF+2)/2) NRD='0.29 NRS='0.29 SA=0 SB=0 SD=0 MULT='N' M='N' 
*--------END___X3_X40_XM2->W'
*--------END___X3_X40->TRANSMISSION_GATE
*--------BEGIN_X3_X41->SWITCH_5T
*.PININFO IN:B OUT:B EN:I EN_B:I
*--------BEGIN_X3_X41_X1->TRANSMISSION_GATE
*.PININFO IN:B OUT:B EN:I EN_B:I
*--------BEGIN_X3_X41_X1_XM1->W'
XM1_X3_X41_X1 X3_X41_NET1 X3_NET25 X3_NET5 X3_VSS X3_X41_X1_SKY130_FD_PR__NFET_01V8 X3_X41_X1_* X3_X41_X1_W/NF X3_X41_X1_* X3_X41_X1_0.29'
+ X3_X41_X1_* X3_X41_X1_W/NF X3_X41_X1_* X3_X41_X1_0.29' X3_X41_X1_* X3_X41_X1_(W/NF X3_X41_X1_+ X3_X41_X1_0.29)'
+ X3_X41_X1_* X3_X41_X1_(W/NF X3_X41_X1_+ X3_X41_X1_0.29)' X3_X41_X1_/ X3_X41_X1_W' X3_X41_X1_/  W' L='L_N' W='W_N' NF=1 AD='INT((NF+1)/2)
+ AS='INT((NF+2)/2) PD='2*INT((NF+1)/2) PS='2*INT((NF+2)/2) NRD='0.29 NRS='0.29 SA=0 SB=0 SD=0 MULT='N' M='N' 
*--------END___X3_X41_X1_XM1->W'
*--------BEGIN_X3_X41_X1_XM2->W'
XM2_X3_X41_X1 X3_X41_NET1 VDD X3_NET5 VDD X3_X41_X1_SKY130_FD_PR__PFET_01V8 X3_X41_X1_* X3_X41_X1_W/NF X3_X41_X1_* X3_X41_X1_0.29'
+ X3_X41_X1_* X3_X41_X1_W/NF X3_X41_X1_* X3_X41_X1_0.29' X3_X41_X1_* X3_X41_X1_(W/NF X3_X41_X1_+ X3_X41_X1_0.29)'
+ X3_X41_X1_* X3_X41_X1_(W/NF X3_X41_X1_+ X3_X41_X1_0.29)' X3_X41_X1_/ X3_X41_X1_W' X3_X41_X1_/  W' L='L_P' W='W_P' NF=1 AD='INT((NF+1)/2)
+ AS='INT((NF+2)/2) PD='2*INT((NF+1)/2) PS='2*INT((NF+2)/2) NRD='0.29 NRS='0.29 SA=0 SB=0 SD=0 MULT='N' M='N' 
*--------END___X3_X41_X1_XM2->W'
*--------END___X3_X41_X1->TRANSMISSION_GATE
*--------BEGIN_X3_X41_X2->TRANSMISSION_GATE
*.PININFO IN:B OUT:B EN:I EN_B:I
*--------BEGIN_X3_X41_X2_XM1->W'
XM1_X3_X41_X2 OUT32 X3_NET25 X3_X41_NET1 X3_VSS X3_X41_X2_SKY130_FD_PR__NFET_01V8 X3_X41_X2_* X3_X41_X2_W/NF X3_X41_X2_* X3_X41_X2_0.29'
+ X3_X41_X2_* X3_X41_X2_W/NF X3_X41_X2_* X3_X41_X2_0.29' X3_X41_X2_* X3_X41_X2_(W/NF X3_X41_X2_+ X3_X41_X2_0.29)'
+ X3_X41_X2_* X3_X41_X2_(W/NF X3_X41_X2_+ X3_X41_X2_0.29)' X3_X41_X2_/ X3_X41_X2_W' X3_X41_X2_/  W' L='L_N' W='W_N' NF=1 AD='INT((NF+1)/2)
+ AS='INT((NF+2)/2) PD='2*INT((NF+1)/2) PS='2*INT((NF+2)/2) NRD='0.29 NRS='0.29 SA=0 SB=0 SD=0 MULT='N' M='N' 
*--------END___X3_X41_X2_XM1->W'
*--------BEGIN_X3_X41_X2_XM2->W'
XM2_X3_X41_X2 OUT32 VDD X3_X41_NET1 VDD X3_X41_X2_SKY130_FD_PR__PFET_01V8 X3_X41_X2_* X3_X41_X2_W/NF X3_X41_X2_* X3_X41_X2_0.29'
+ X3_X41_X2_* X3_X41_X2_W/NF X3_X41_X2_* X3_X41_X2_0.29' X3_X41_X2_* X3_X41_X2_(W/NF X3_X41_X2_+ X3_X41_X2_0.29)'
+ X3_X41_X2_* X3_X41_X2_(W/NF X3_X41_X2_+ X3_X41_X2_0.29)' X3_X41_X2_/ X3_X41_X2_W' X3_X41_X2_/  W' L='L_P' W='W_P' NF=1 AD='INT((NF+1)/2)
+ AS='INT((NF+2)/2) PD='2*INT((NF+1)/2) PS='2*INT((NF+2)/2) NRD='0.29 NRS='0.29 SA=0 SB=0 SD=0 MULT='N' M='N' 
*--------END___X3_X41_X2_XM2->W'
*--------END___X3_X41_X2->TRANSMISSION_GATE
*--------BEGIN_X3_X41_XM1->W'
XM1_X3_X41 X3_X41_NET1 VDD X3_VSS X3_VSS X3_X41_SKY130_FD_PR__NFET_01V8 X3_X41_* X3_X41_W/NF X3_X41_* X3_X41_0.29'
+ X3_X41_* X3_X41_W/NF X3_X41_* X3_X41_0.29' X3_X41_* X3_X41_(W/NF X3_X41_+ X3_X41_0.29)' X3_X41_* X3_X41_(W/NF
+ X3_X41_+ X3_X41_0.29)' X3_X41_/ X3_X41_W' X3_X41_/  W' L=0.15 W=0.5 NF=1 AD='INT((NF+1)/2) AS='INT((NF+2)/2) PD='2*INT((NF+1)/2)
+ PS='2*INT((NF+2)/2) NRD='0.29 NRS='0.29 SA=0 SB=0 SD=0 MULT=1 M=1 
*--------END___X3_X41_XM1->W'
*--------END___X3_X41->SWITCH_5T
*--------BEGIN_X3_X42->SKY130_FD_SC_HD__INV_1
X42_X3 VDD X3_VGND X3_VNB X3_VPB X3_VPWR X3_NET25  SKY130_FD_SC_HD__INV_1
*--------END___X3_X42->SKY130_FD_SC_HD__INV_1
*--------BEGIN_X3_X43->TRANSMISSION_GATE
*.PININFO IN:B OUT:B EN:I EN_B:I
*--------BEGIN_X3_X43_XM1->W'
XM1_X3_X43 X3_NET6 VDD IN15 X3_VSS X3_X43_SKY130_FD_PR__NFET_01V8 X3_X43_* X3_X43_W/NF X3_X43_* X3_X43_0.29'
+ X3_X43_* X3_X43_W/NF X3_X43_* X3_X43_0.29' X3_X43_* X3_X43_(W/NF X3_X43_+ X3_X43_0.29)' X3_X43_* X3_X43_(W/NF
+ X3_X43_+ X3_X43_0.29)' X3_X43_/ X3_X43_W' X3_X43_/  W' L='L_N' W='W_N' NF=1 AD='INT((NF+1)/2) AS='INT((NF+2)/2) PD='2*INT((NF+1)/2)
+ PS='2*INT((NF+2)/2) NRD='0.29 NRS='0.29 SA=0 SB=0 SD=0 MULT='N' M='N' 
*--------END___X3_X43_XM1->W'
*--------BEGIN_X3_X43_XM2->W'
XM2_X3_X43 X3_NET6 GND IN15 VDD X3_X43_SKY130_FD_PR__PFET_01V8 X3_X43_* X3_X43_W/NF X3_X43_* X3_X43_0.29'
+ X3_X43_* X3_X43_W/NF X3_X43_* X3_X43_0.29' X3_X43_* X3_X43_(W/NF X3_X43_+ X3_X43_0.29)' X3_X43_* X3_X43_(W/NF
+ X3_X43_+ X3_X43_0.29)' X3_X43_/ X3_X43_W' X3_X43_/  W' L='L_P' W='W_P' NF=1 AD='INT((NF+1)/2) AS='INT((NF+2)/2) PD='2*INT((NF+1)/2)
+ PS='2*INT((NF+2)/2) NRD='0.29 NRS='0.29 SA=0 SB=0 SD=0 MULT='N' M='N' 
*--------END___X3_X43_XM2->W'
*--------END___X3_X43->TRANSMISSION_GATE
*--------BEGIN_X3_X44->SWITCH_5T
*.PININFO IN:B OUT:B EN:I EN_B:I
*--------BEGIN_X3_X44_X1->TRANSMISSION_GATE
*.PININFO IN:B OUT:B EN:I EN_B:I
*--------BEGIN_X3_X44_X1_XM1->W'
XM1_X3_X44_X1 X3_X44_NET1 X3_NET26 X3_NET6 X3_VSS X3_X44_X1_SKY130_FD_PR__NFET_01V8 X3_X44_X1_* X3_X44_X1_W/NF X3_X44_X1_* X3_X44_X1_0.29'
+ X3_X44_X1_* X3_X44_X1_W/NF X3_X44_X1_* X3_X44_X1_0.29' X3_X44_X1_* X3_X44_X1_(W/NF X3_X44_X1_+ X3_X44_X1_0.29)'
+ X3_X44_X1_* X3_X44_X1_(W/NF X3_X44_X1_+ X3_X44_X1_0.29)' X3_X44_X1_/ X3_X44_X1_W' X3_X44_X1_/  W' L='L_N' W='W_N' NF=1 AD='INT((NF+1)/2)
+ AS='INT((NF+2)/2) PD='2*INT((NF+1)/2) PS='2*INT((NF+2)/2) NRD='0.29 NRS='0.29 SA=0 SB=0 SD=0 MULT='N' M='N' 
*--------END___X3_X44_X1_XM1->W'
*--------BEGIN_X3_X44_X1_XM2->W'
XM2_X3_X44_X1 X3_X44_NET1 VDD X3_NET6 VDD X3_X44_X1_SKY130_FD_PR__PFET_01V8 X3_X44_X1_* X3_X44_X1_W/NF X3_X44_X1_* X3_X44_X1_0.29'
+ X3_X44_X1_* X3_X44_X1_W/NF X3_X44_X1_* X3_X44_X1_0.29' X3_X44_X1_* X3_X44_X1_(W/NF X3_X44_X1_+ X3_X44_X1_0.29)'
+ X3_X44_X1_* X3_X44_X1_(W/NF X3_X44_X1_+ X3_X44_X1_0.29)' X3_X44_X1_/ X3_X44_X1_W' X3_X44_X1_/  W' L='L_P' W='W_P' NF=1 AD='INT((NF+1)/2)
+ AS='INT((NF+2)/2) PD='2*INT((NF+1)/2) PS='2*INT((NF+2)/2) NRD='0.29 NRS='0.29 SA=0 SB=0 SD=0 MULT='N' M='N' 
*--------END___X3_X44_X1_XM2->W'
*--------END___X3_X44_X1->TRANSMISSION_GATE
*--------BEGIN_X3_X44_X2->TRANSMISSION_GATE
*.PININFO IN:B OUT:B EN:I EN_B:I
*--------BEGIN_X3_X44_X2_XM1->W'
XM1_X3_X44_X2 OUT32 X3_NET26 X3_X44_NET1 X3_VSS X3_X44_X2_SKY130_FD_PR__NFET_01V8 X3_X44_X2_* X3_X44_X2_W/NF X3_X44_X2_* X3_X44_X2_0.29'
+ X3_X44_X2_* X3_X44_X2_W/NF X3_X44_X2_* X3_X44_X2_0.29' X3_X44_X2_* X3_X44_X2_(W/NF X3_X44_X2_+ X3_X44_X2_0.29)'
+ X3_X44_X2_* X3_X44_X2_(W/NF X3_X44_X2_+ X3_X44_X2_0.29)' X3_X44_X2_/ X3_X44_X2_W' X3_X44_X2_/  W' L='L_N' W='W_N' NF=1 AD='INT((NF+1)/2)
+ AS='INT((NF+2)/2) PD='2*INT((NF+1)/2) PS='2*INT((NF+2)/2) NRD='0.29 NRS='0.29 SA=0 SB=0 SD=0 MULT='N' M='N' 
*--------END___X3_X44_X2_XM1->W'
*--------BEGIN_X3_X44_X2_XM2->W'
XM2_X3_X44_X2 OUT32 VDD X3_X44_NET1 VDD X3_X44_X2_SKY130_FD_PR__PFET_01V8 X3_X44_X2_* X3_X44_X2_W/NF X3_X44_X2_* X3_X44_X2_0.29'
+ X3_X44_X2_* X3_X44_X2_W/NF X3_X44_X2_* X3_X44_X2_0.29' X3_X44_X2_* X3_X44_X2_(W/NF X3_X44_X2_+ X3_X44_X2_0.29)'
+ X3_X44_X2_* X3_X44_X2_(W/NF X3_X44_X2_+ X3_X44_X2_0.29)' X3_X44_X2_/ X3_X44_X2_W' X3_X44_X2_/  W' L='L_P' W='W_P' NF=1 AD='INT((NF+1)/2)
+ AS='INT((NF+2)/2) PD='2*INT((NF+1)/2) PS='2*INT((NF+2)/2) NRD='0.29 NRS='0.29 SA=0 SB=0 SD=0 MULT='N' M='N' 
*--------END___X3_X44_X2_XM2->W'
*--------END___X3_X44_X2->TRANSMISSION_GATE
*--------BEGIN_X3_X44_XM1->W'
XM1_X3_X44 X3_X44_NET1 VDD X3_VSS X3_VSS X3_X44_SKY130_FD_PR__NFET_01V8 X3_X44_* X3_X44_W/NF X3_X44_* X3_X44_0.29'
+ X3_X44_* X3_X44_W/NF X3_X44_* X3_X44_0.29' X3_X44_* X3_X44_(W/NF X3_X44_+ X3_X44_0.29)' X3_X44_* X3_X44_(W/NF
+ X3_X44_+ X3_X44_0.29)' X3_X44_/ X3_X44_W' X3_X44_/  W' L=0.15 W=0.5 NF=1 AD='INT((NF+1)/2) AS='INT((NF+2)/2) PD='2*INT((NF+1)/2)
+ PS='2*INT((NF+2)/2) NRD='0.29 NRS='0.29 SA=0 SB=0 SD=0 MULT=1 M=1 
*--------END___X3_X44_XM1->W'
*--------END___X3_X44->SWITCH_5T
*--------BEGIN_X3_X45->SKY130_FD_SC_HD__INV_1
X45_X3 VDD X3_VGND X3_VNB X3_VPB X3_VPWR X3_NET26  SKY130_FD_SC_HD__INV_1
*--------END___X3_X45->SKY130_FD_SC_HD__INV_1
*--------BEGIN_X3_X46->TRANSMISSION_GATE
*.PININFO IN:B OUT:B EN:I EN_B:I
*--------BEGIN_X3_X46_XM1->W'
XM1_X3_X46 X3_NET7 VDD IN16 X3_VSS X3_X46_SKY130_FD_PR__NFET_01V8 X3_X46_* X3_X46_W/NF X3_X46_* X3_X46_0.29'
+ X3_X46_* X3_X46_W/NF X3_X46_* X3_X46_0.29' X3_X46_* X3_X46_(W/NF X3_X46_+ X3_X46_0.29)' X3_X46_* X3_X46_(W/NF
+ X3_X46_+ X3_X46_0.29)' X3_X46_/ X3_X46_W' X3_X46_/  W' L='L_N' W='W_N' NF=1 AD='INT((NF+1)/2) AS='INT((NF+2)/2) PD='2*INT((NF+1)/2)
+ PS='2*INT((NF+2)/2) NRD='0.29 NRS='0.29 SA=0 SB=0 SD=0 MULT='N' M='N' 
*--------END___X3_X46_XM1->W'
*--------BEGIN_X3_X46_XM2->W'
XM2_X3_X46 X3_NET7 GND IN16 VDD X3_X46_SKY130_FD_PR__PFET_01V8 X3_X46_* X3_X46_W/NF X3_X46_* X3_X46_0.29'
+ X3_X46_* X3_X46_W/NF X3_X46_* X3_X46_0.29' X3_X46_* X3_X46_(W/NF X3_X46_+ X3_X46_0.29)' X3_X46_* X3_X46_(W/NF
+ X3_X46_+ X3_X46_0.29)' X3_X46_/ X3_X46_W' X3_X46_/  W' L='L_P' W='W_P' NF=1 AD='INT((NF+1)/2) AS='INT((NF+2)/2) PD='2*INT((NF+1)/2)
+ PS='2*INT((NF+2)/2) NRD='0.29 NRS='0.29 SA=0 SB=0 SD=0 MULT='N' M='N' 
*--------END___X3_X46_XM2->W'
*--------END___X3_X46->TRANSMISSION_GATE
*--------BEGIN_X3_X47->SWITCH_5T
*.PININFO IN:B OUT:B EN:I EN_B:I
*--------BEGIN_X3_X47_X1->TRANSMISSION_GATE
*.PININFO IN:B OUT:B EN:I EN_B:I
*--------BEGIN_X3_X47_X1_XM1->W'
XM1_X3_X47_X1 X3_X47_NET1 X3_NET27 X3_NET7 X3_VSS X3_X47_X1_SKY130_FD_PR__NFET_01V8 X3_X47_X1_* X3_X47_X1_W/NF X3_X47_X1_* X3_X47_X1_0.29'
+ X3_X47_X1_* X3_X47_X1_W/NF X3_X47_X1_* X3_X47_X1_0.29' X3_X47_X1_* X3_X47_X1_(W/NF X3_X47_X1_+ X3_X47_X1_0.29)'
+ X3_X47_X1_* X3_X47_X1_(W/NF X3_X47_X1_+ X3_X47_X1_0.29)' X3_X47_X1_/ X3_X47_X1_W' X3_X47_X1_/  W' L='L_N' W='W_N' NF=1 AD='INT((NF+1)/2)
+ AS='INT((NF+2)/2) PD='2*INT((NF+1)/2) PS='2*INT((NF+2)/2) NRD='0.29 NRS='0.29 SA=0 SB=0 SD=0 MULT='N' M='N' 
*--------END___X3_X47_X1_XM1->W'
*--------BEGIN_X3_X47_X1_XM2->W'
XM2_X3_X47_X1 X3_X47_NET1 VDD X3_NET7 VDD X3_X47_X1_SKY130_FD_PR__PFET_01V8 X3_X47_X1_* X3_X47_X1_W/NF X3_X47_X1_* X3_X47_X1_0.29'
+ X3_X47_X1_* X3_X47_X1_W/NF X3_X47_X1_* X3_X47_X1_0.29' X3_X47_X1_* X3_X47_X1_(W/NF X3_X47_X1_+ X3_X47_X1_0.29)'
+ X3_X47_X1_* X3_X47_X1_(W/NF X3_X47_X1_+ X3_X47_X1_0.29)' X3_X47_X1_/ X3_X47_X1_W' X3_X47_X1_/  W' L='L_P' W='W_P' NF=1 AD='INT((NF+1)/2)
+ AS='INT((NF+2)/2) PD='2*INT((NF+1)/2) PS='2*INT((NF+2)/2) NRD='0.29 NRS='0.29 SA=0 SB=0 SD=0 MULT='N' M='N' 
*--------END___X3_X47_X1_XM2->W'
*--------END___X3_X47_X1->TRANSMISSION_GATE
*--------BEGIN_X3_X47_X2->TRANSMISSION_GATE
*.PININFO IN:B OUT:B EN:I EN_B:I
*--------BEGIN_X3_X47_X2_XM1->W'
XM1_X3_X47_X2 OUT32 X3_NET27 X3_X47_NET1 X3_VSS X3_X47_X2_SKY130_FD_PR__NFET_01V8 X3_X47_X2_* X3_X47_X2_W/NF X3_X47_X2_* X3_X47_X2_0.29'
+ X3_X47_X2_* X3_X47_X2_W/NF X3_X47_X2_* X3_X47_X2_0.29' X3_X47_X2_* X3_X47_X2_(W/NF X3_X47_X2_+ X3_X47_X2_0.29)'
+ X3_X47_X2_* X3_X47_X2_(W/NF X3_X47_X2_+ X3_X47_X2_0.29)' X3_X47_X2_/ X3_X47_X2_W' X3_X47_X2_/  W' L='L_N' W='W_N' NF=1 AD='INT((NF+1)/2)
+ AS='INT((NF+2)/2) PD='2*INT((NF+1)/2) PS='2*INT((NF+2)/2) NRD='0.29 NRS='0.29 SA=0 SB=0 SD=0 MULT='N' M='N' 
*--------END___X3_X47_X2_XM1->W'
*--------BEGIN_X3_X47_X2_XM2->W'
XM2_X3_X47_X2 OUT32 VDD X3_X47_NET1 VDD X3_X47_X2_SKY130_FD_PR__PFET_01V8 X3_X47_X2_* X3_X47_X2_W/NF X3_X47_X2_* X3_X47_X2_0.29'
+ X3_X47_X2_* X3_X47_X2_W/NF X3_X47_X2_* X3_X47_X2_0.29' X3_X47_X2_* X3_X47_X2_(W/NF X3_X47_X2_+ X3_X47_X2_0.29)'
+ X3_X47_X2_* X3_X47_X2_(W/NF X3_X47_X2_+ X3_X47_X2_0.29)' X3_X47_X2_/ X3_X47_X2_W' X3_X47_X2_/  W' L='L_P' W='W_P' NF=1 AD='INT((NF+1)/2)
+ AS='INT((NF+2)/2) PD='2*INT((NF+1)/2) PS='2*INT((NF+2)/2) NRD='0.29 NRS='0.29 SA=0 SB=0 SD=0 MULT='N' M='N' 
*--------END___X3_X47_X2_XM2->W'
*--------END___X3_X47_X2->TRANSMISSION_GATE
*--------BEGIN_X3_X47_XM1->W'
XM1_X3_X47 X3_X47_NET1 VDD X3_VSS X3_VSS X3_X47_SKY130_FD_PR__NFET_01V8 X3_X47_* X3_X47_W/NF X3_X47_* X3_X47_0.29'
+ X3_X47_* X3_X47_W/NF X3_X47_* X3_X47_0.29' X3_X47_* X3_X47_(W/NF X3_X47_+ X3_X47_0.29)' X3_X47_* X3_X47_(W/NF
+ X3_X47_+ X3_X47_0.29)' X3_X47_/ X3_X47_W' X3_X47_/  W' L=0.15 W=0.5 NF=1 AD='INT((NF+1)/2) AS='INT((NF+2)/2) PD='2*INT((NF+1)/2)
+ PS='2*INT((NF+2)/2) NRD='0.29 NRS='0.29 SA=0 SB=0 SD=0 MULT=1 M=1 
*--------END___X3_X47_XM1->W'
*--------END___X3_X47->SWITCH_5T
*--------BEGIN_X3_X48->SKY130_FD_SC_HD__INV_1
X48_X3 VDD X3_VGND X3_VNB X3_VPB X3_VPWR X3_NET27  SKY130_FD_SC_HD__INV_1
*--------END___X3_X48->SKY130_FD_SC_HD__INV_1
*--------BEGIN_X3_X49->TRANSMISSION_GATE
*.PININFO IN:B OUT:B EN:I EN_B:I
*--------BEGIN_X3_X49_XM1->W'
XM1_X3_X49 X3_NET8 VDD IN17 X3_VSS X3_X49_SKY130_FD_PR__NFET_01V8 X3_X49_* X3_X49_W/NF X3_X49_* X3_X49_0.29'
+ X3_X49_* X3_X49_W/NF X3_X49_* X3_X49_0.29' X3_X49_* X3_X49_(W/NF X3_X49_+ X3_X49_0.29)' X3_X49_* X3_X49_(W/NF
+ X3_X49_+ X3_X49_0.29)' X3_X49_/ X3_X49_W' X3_X49_/  W' L='L_N' W='W_N' NF=1 AD='INT((NF+1)/2) AS='INT((NF+2)/2) PD='2*INT((NF+1)/2)
+ PS='2*INT((NF+2)/2) NRD='0.29 NRS='0.29 SA=0 SB=0 SD=0 MULT='N' M='N' 
*--------END___X3_X49_XM1->W'
*--------BEGIN_X3_X49_XM2->W'
XM2_X3_X49 X3_NET8 GND IN17 VDD X3_X49_SKY130_FD_PR__PFET_01V8 X3_X49_* X3_X49_W/NF X3_X49_* X3_X49_0.29'
+ X3_X49_* X3_X49_W/NF X3_X49_* X3_X49_0.29' X3_X49_* X3_X49_(W/NF X3_X49_+ X3_X49_0.29)' X3_X49_* X3_X49_(W/NF
+ X3_X49_+ X3_X49_0.29)' X3_X49_/ X3_X49_W' X3_X49_/  W' L='L_P' W='W_P' NF=1 AD='INT((NF+1)/2) AS='INT((NF+2)/2) PD='2*INT((NF+1)/2)
+ PS='2*INT((NF+2)/2) NRD='0.29 NRS='0.29 SA=0 SB=0 SD=0 MULT='N' M='N' 
*--------END___X3_X49_XM2->W'
*--------END___X3_X49->TRANSMISSION_GATE
*--------BEGIN_X3_X50->SWITCH_5T
*.PININFO IN:B OUT:B EN:I EN_B:I
*--------BEGIN_X3_X50_X1->TRANSMISSION_GATE
*.PININFO IN:B OUT:B EN:I EN_B:I
*--------BEGIN_X3_X50_X1_XM1->W'
XM1_X3_X50_X1 X3_X50_NET1 X3_NET28 X3_NET8 X3_VSS X3_X50_X1_SKY130_FD_PR__NFET_01V8 X3_X50_X1_* X3_X50_X1_W/NF X3_X50_X1_* X3_X50_X1_0.29'
+ X3_X50_X1_* X3_X50_X1_W/NF X3_X50_X1_* X3_X50_X1_0.29' X3_X50_X1_* X3_X50_X1_(W/NF X3_X50_X1_+ X3_X50_X1_0.29)'
+ X3_X50_X1_* X3_X50_X1_(W/NF X3_X50_X1_+ X3_X50_X1_0.29)' X3_X50_X1_/ X3_X50_X1_W' X3_X50_X1_/  W' L='L_N' W='W_N' NF=1 AD='INT((NF+1)/2)
+ AS='INT((NF+2)/2) PD='2*INT((NF+1)/2) PS='2*INT((NF+2)/2) NRD='0.29 NRS='0.29 SA=0 SB=0 SD=0 MULT='N' M='N' 
*--------END___X3_X50_X1_XM1->W'
*--------BEGIN_X3_X50_X1_XM2->W'
XM2_X3_X50_X1 X3_X50_NET1 VDD X3_NET8 VDD X3_X50_X1_SKY130_FD_PR__PFET_01V8 X3_X50_X1_* X3_X50_X1_W/NF X3_X50_X1_* X3_X50_X1_0.29'
+ X3_X50_X1_* X3_X50_X1_W/NF X3_X50_X1_* X3_X50_X1_0.29' X3_X50_X1_* X3_X50_X1_(W/NF X3_X50_X1_+ X3_X50_X1_0.29)'
+ X3_X50_X1_* X3_X50_X1_(W/NF X3_X50_X1_+ X3_X50_X1_0.29)' X3_X50_X1_/ X3_X50_X1_W' X3_X50_X1_/  W' L='L_P' W='W_P' NF=1 AD='INT((NF+1)/2)
+ AS='INT((NF+2)/2) PD='2*INT((NF+1)/2) PS='2*INT((NF+2)/2) NRD='0.29 NRS='0.29 SA=0 SB=0 SD=0 MULT='N' M='N' 
*--------END___X3_X50_X1_XM2->W'
*--------END___X3_X50_X1->TRANSMISSION_GATE
*--------BEGIN_X3_X50_X2->TRANSMISSION_GATE
*.PININFO IN:B OUT:B EN:I EN_B:I
*--------BEGIN_X3_X50_X2_XM1->W'
XM1_X3_X50_X2 OUT32 X3_NET28 X3_X50_NET1 X3_VSS X3_X50_X2_SKY130_FD_PR__NFET_01V8 X3_X50_X2_* X3_X50_X2_W/NF X3_X50_X2_* X3_X50_X2_0.29'
+ X3_X50_X2_* X3_X50_X2_W/NF X3_X50_X2_* X3_X50_X2_0.29' X3_X50_X2_* X3_X50_X2_(W/NF X3_X50_X2_+ X3_X50_X2_0.29)'
+ X3_X50_X2_* X3_X50_X2_(W/NF X3_X50_X2_+ X3_X50_X2_0.29)' X3_X50_X2_/ X3_X50_X2_W' X3_X50_X2_/  W' L='L_N' W='W_N' NF=1 AD='INT((NF+1)/2)
+ AS='INT((NF+2)/2) PD='2*INT((NF+1)/2) PS='2*INT((NF+2)/2) NRD='0.29 NRS='0.29 SA=0 SB=0 SD=0 MULT='N' M='N' 
*--------END___X3_X50_X2_XM1->W'
*--------BEGIN_X3_X50_X2_XM2->W'
XM2_X3_X50_X2 OUT32 VDD X3_X50_NET1 VDD X3_X50_X2_SKY130_FD_PR__PFET_01V8 X3_X50_X2_* X3_X50_X2_W/NF X3_X50_X2_* X3_X50_X2_0.29'
+ X3_X50_X2_* X3_X50_X2_W/NF X3_X50_X2_* X3_X50_X2_0.29' X3_X50_X2_* X3_X50_X2_(W/NF X3_X50_X2_+ X3_X50_X2_0.29)'
+ X3_X50_X2_* X3_X50_X2_(W/NF X3_X50_X2_+ X3_X50_X2_0.29)' X3_X50_X2_/ X3_X50_X2_W' X3_X50_X2_/  W' L='L_P' W='W_P' NF=1 AD='INT((NF+1)/2)
+ AS='INT((NF+2)/2) PD='2*INT((NF+1)/2) PS='2*INT((NF+2)/2) NRD='0.29 NRS='0.29 SA=0 SB=0 SD=0 MULT='N' M='N' 
*--------END___X3_X50_X2_XM2->W'
*--------END___X3_X50_X2->TRANSMISSION_GATE
*--------BEGIN_X3_X50_XM1->W'
XM1_X3_X50 X3_X50_NET1 VDD X3_VSS X3_VSS X3_X50_SKY130_FD_PR__NFET_01V8 X3_X50_* X3_X50_W/NF X3_X50_* X3_X50_0.29'
+ X3_X50_* X3_X50_W/NF X3_X50_* X3_X50_0.29' X3_X50_* X3_X50_(W/NF X3_X50_+ X3_X50_0.29)' X3_X50_* X3_X50_(W/NF
+ X3_X50_+ X3_X50_0.29)' X3_X50_/ X3_X50_W' X3_X50_/  W' L=0.15 W=0.5 NF=1 AD='INT((NF+1)/2) AS='INT((NF+2)/2) PD='2*INT((NF+1)/2)
+ PS='2*INT((NF+2)/2) NRD='0.29 NRS='0.29 SA=0 SB=0 SD=0 MULT=1 M=1 
*--------END___X3_X50_XM1->W'
*--------END___X3_X50->SWITCH_5T
*--------BEGIN_X3_X51->SKY130_FD_SC_HD__INV_1
X51_X3 VDD X3_VGND X3_VNB X3_VPB X3_VPWR X3_NET28  SKY130_FD_SC_HD__INV_1
*--------END___X3_X51->SKY130_FD_SC_HD__INV_1
*--------BEGIN_X3_X52->TRANSMISSION_GATE
*.PININFO IN:B OUT:B EN:I EN_B:I
*--------BEGIN_X3_X52_XM1->W'
XM1_X3_X52 X3_NET9 VDD IN18 X3_VSS X3_X52_SKY130_FD_PR__NFET_01V8 X3_X52_* X3_X52_W/NF X3_X52_* X3_X52_0.29'
+ X3_X52_* X3_X52_W/NF X3_X52_* X3_X52_0.29' X3_X52_* X3_X52_(W/NF X3_X52_+ X3_X52_0.29)' X3_X52_* X3_X52_(W/NF
+ X3_X52_+ X3_X52_0.29)' X3_X52_/ X3_X52_W' X3_X52_/  W' L='L_N' W='W_N' NF=1 AD='INT((NF+1)/2) AS='INT((NF+2)/2) PD='2*INT((NF+1)/2)
+ PS='2*INT((NF+2)/2) NRD='0.29 NRS='0.29 SA=0 SB=0 SD=0 MULT='N' M='N' 
*--------END___X3_X52_XM1->W'
*--------BEGIN_X3_X52_XM2->W'
XM2_X3_X52 X3_NET9 GND IN18 VDD X3_X52_SKY130_FD_PR__PFET_01V8 X3_X52_* X3_X52_W/NF X3_X52_* X3_X52_0.29'
+ X3_X52_* X3_X52_W/NF X3_X52_* X3_X52_0.29' X3_X52_* X3_X52_(W/NF X3_X52_+ X3_X52_0.29)' X3_X52_* X3_X52_(W/NF
+ X3_X52_+ X3_X52_0.29)' X3_X52_/ X3_X52_W' X3_X52_/  W' L='L_P' W='W_P' NF=1 AD='INT((NF+1)/2) AS='INT((NF+2)/2) PD='2*INT((NF+1)/2)
+ PS='2*INT((NF+2)/2) NRD='0.29 NRS='0.29 SA=0 SB=0 SD=0 MULT='N' M='N' 
*--------END___X3_X52_XM2->W'
*--------END___X3_X52->TRANSMISSION_GATE
*--------BEGIN_X3_X53->SWITCH_5T
*.PININFO IN:B OUT:B EN:I EN_B:I
*--------BEGIN_X3_X53_X1->TRANSMISSION_GATE
*.PININFO IN:B OUT:B EN:I EN_B:I
*--------BEGIN_X3_X53_X1_XM1->W'
XM1_X3_X53_X1 X3_X53_NET1 X3_NET29 X3_NET9 X3_VSS X3_X53_X1_SKY130_FD_PR__NFET_01V8 X3_X53_X1_* X3_X53_X1_W/NF X3_X53_X1_* X3_X53_X1_0.29'
+ X3_X53_X1_* X3_X53_X1_W/NF X3_X53_X1_* X3_X53_X1_0.29' X3_X53_X1_* X3_X53_X1_(W/NF X3_X53_X1_+ X3_X53_X1_0.29)'
+ X3_X53_X1_* X3_X53_X1_(W/NF X3_X53_X1_+ X3_X53_X1_0.29)' X3_X53_X1_/ X3_X53_X1_W' X3_X53_X1_/  W' L='L_N' W='W_N' NF=1 AD='INT((NF+1)/2)
+ AS='INT((NF+2)/2) PD='2*INT((NF+1)/2) PS='2*INT((NF+2)/2) NRD='0.29 NRS='0.29 SA=0 SB=0 SD=0 MULT='N' M='N' 
*--------END___X3_X53_X1_XM1->W'
*--------BEGIN_X3_X53_X1_XM2->W'
XM2_X3_X53_X1 X3_X53_NET1 VDD X3_NET9 VDD X3_X53_X1_SKY130_FD_PR__PFET_01V8 X3_X53_X1_* X3_X53_X1_W/NF X3_X53_X1_* X3_X53_X1_0.29'
+ X3_X53_X1_* X3_X53_X1_W/NF X3_X53_X1_* X3_X53_X1_0.29' X3_X53_X1_* X3_X53_X1_(W/NF X3_X53_X1_+ X3_X53_X1_0.29)'
+ X3_X53_X1_* X3_X53_X1_(W/NF X3_X53_X1_+ X3_X53_X1_0.29)' X3_X53_X1_/ X3_X53_X1_W' X3_X53_X1_/  W' L='L_P' W='W_P' NF=1 AD='INT((NF+1)/2)
+ AS='INT((NF+2)/2) PD='2*INT((NF+1)/2) PS='2*INT((NF+2)/2) NRD='0.29 NRS='0.29 SA=0 SB=0 SD=0 MULT='N' M='N' 
*--------END___X3_X53_X1_XM2->W'
*--------END___X3_X53_X1->TRANSMISSION_GATE
*--------BEGIN_X3_X53_X2->TRANSMISSION_GATE
*.PININFO IN:B OUT:B EN:I EN_B:I
*--------BEGIN_X3_X53_X2_XM1->W'
XM1_X3_X53_X2 OUT32 X3_NET29 X3_X53_NET1 X3_VSS X3_X53_X2_SKY130_FD_PR__NFET_01V8 X3_X53_X2_* X3_X53_X2_W/NF X3_X53_X2_* X3_X53_X2_0.29'
+ X3_X53_X2_* X3_X53_X2_W/NF X3_X53_X2_* X3_X53_X2_0.29' X3_X53_X2_* X3_X53_X2_(W/NF X3_X53_X2_+ X3_X53_X2_0.29)'
+ X3_X53_X2_* X3_X53_X2_(W/NF X3_X53_X2_+ X3_X53_X2_0.29)' X3_X53_X2_/ X3_X53_X2_W' X3_X53_X2_/  W' L='L_N' W='W_N' NF=1 AD='INT((NF+1)/2)
+ AS='INT((NF+2)/2) PD='2*INT((NF+1)/2) PS='2*INT((NF+2)/2) NRD='0.29 NRS='0.29 SA=0 SB=0 SD=0 MULT='N' M='N' 
*--------END___X3_X53_X2_XM1->W'
*--------BEGIN_X3_X53_X2_XM2->W'
XM2_X3_X53_X2 OUT32 VDD X3_X53_NET1 VDD X3_X53_X2_SKY130_FD_PR__PFET_01V8 X3_X53_X2_* X3_X53_X2_W/NF X3_X53_X2_* X3_X53_X2_0.29'
+ X3_X53_X2_* X3_X53_X2_W/NF X3_X53_X2_* X3_X53_X2_0.29' X3_X53_X2_* X3_X53_X2_(W/NF X3_X53_X2_+ X3_X53_X2_0.29)'
+ X3_X53_X2_* X3_X53_X2_(W/NF X3_X53_X2_+ X3_X53_X2_0.29)' X3_X53_X2_/ X3_X53_X2_W' X3_X53_X2_/  W' L='L_P' W='W_P' NF=1 AD='INT((NF+1)/2)
+ AS='INT((NF+2)/2) PD='2*INT((NF+1)/2) PS='2*INT((NF+2)/2) NRD='0.29 NRS='0.29 SA=0 SB=0 SD=0 MULT='N' M='N' 
*--------END___X3_X53_X2_XM2->W'
*--------END___X3_X53_X2->TRANSMISSION_GATE
*--------BEGIN_X3_X53_XM1->W'
XM1_X3_X53 X3_X53_NET1 VDD X3_VSS X3_VSS X3_X53_SKY130_FD_PR__NFET_01V8 X3_X53_* X3_X53_W/NF X3_X53_* X3_X53_0.29'
+ X3_X53_* X3_X53_W/NF X3_X53_* X3_X53_0.29' X3_X53_* X3_X53_(W/NF X3_X53_+ X3_X53_0.29)' X3_X53_* X3_X53_(W/NF
+ X3_X53_+ X3_X53_0.29)' X3_X53_/ X3_X53_W' X3_X53_/  W' L=0.15 W=0.5 NF=1 AD='INT((NF+1)/2) AS='INT((NF+2)/2) PD='2*INT((NF+1)/2)
+ PS='2*INT((NF+2)/2) NRD='0.29 NRS='0.29 SA=0 SB=0 SD=0 MULT=1 M=1 
*--------END___X3_X53_XM1->W'
*--------END___X3_X53->SWITCH_5T
*--------BEGIN_X3_X54->SKY130_FD_SC_HD__INV_1
X54_X3 VDD X3_VGND X3_VNB X3_VPB X3_VPWR X3_NET29  SKY130_FD_SC_HD__INV_1
*--------END___X3_X54->SKY130_FD_SC_HD__INV_1
*--------BEGIN_X3_X55->TRANSMISSION_GATE
*.PININFO IN:B OUT:B EN:I EN_B:I
*--------BEGIN_X3_X55_XM1->W'
XM1_X3_X55 X3_NET10 VDD IN19 X3_VSS X3_X55_SKY130_FD_PR__NFET_01V8 X3_X55_* X3_X55_W/NF X3_X55_* X3_X55_0.29'
+ X3_X55_* X3_X55_W/NF X3_X55_* X3_X55_0.29' X3_X55_* X3_X55_(W/NF X3_X55_+ X3_X55_0.29)' X3_X55_* X3_X55_(W/NF
+ X3_X55_+ X3_X55_0.29)' X3_X55_/ X3_X55_W' X3_X55_/  W' L='L_N' W='W_N' NF=1 AD='INT((NF+1)/2) AS='INT((NF+2)/2) PD='2*INT((NF+1)/2)
+ PS='2*INT((NF+2)/2) NRD='0.29 NRS='0.29 SA=0 SB=0 SD=0 MULT='N' M='N' 
*--------END___X3_X55_XM1->W'
*--------BEGIN_X3_X55_XM2->W'
XM2_X3_X55 X3_NET10 GND IN19 VDD X3_X55_SKY130_FD_PR__PFET_01V8 X3_X55_* X3_X55_W/NF X3_X55_* X3_X55_0.29'
+ X3_X55_* X3_X55_W/NF X3_X55_* X3_X55_0.29' X3_X55_* X3_X55_(W/NF X3_X55_+ X3_X55_0.29)' X3_X55_* X3_X55_(W/NF
+ X3_X55_+ X3_X55_0.29)' X3_X55_/ X3_X55_W' X3_X55_/  W' L='L_P' W='W_P' NF=1 AD='INT((NF+1)/2) AS='INT((NF+2)/2) PD='2*INT((NF+1)/2)
+ PS='2*INT((NF+2)/2) NRD='0.29 NRS='0.29 SA=0 SB=0 SD=0 MULT='N' M='N' 
*--------END___X3_X55_XM2->W'
*--------END___X3_X55->TRANSMISSION_GATE
*--------BEGIN_X3_X56->SWITCH_5T
*.PININFO IN:B OUT:B EN:I EN_B:I
*--------BEGIN_X3_X56_X1->TRANSMISSION_GATE
*.PININFO IN:B OUT:B EN:I EN_B:I
*--------BEGIN_X3_X56_X1_XM1->W'
XM1_X3_X56_X1 X3_X56_NET1 X3_NET30 X3_NET10 X3_VSS X3_X56_X1_SKY130_FD_PR__NFET_01V8 X3_X56_X1_* X3_X56_X1_W/NF X3_X56_X1_* X3_X56_X1_0.29'
+ X3_X56_X1_* X3_X56_X1_W/NF X3_X56_X1_* X3_X56_X1_0.29' X3_X56_X1_* X3_X56_X1_(W/NF X3_X56_X1_+ X3_X56_X1_0.29)'
+ X3_X56_X1_* X3_X56_X1_(W/NF X3_X56_X1_+ X3_X56_X1_0.29)' X3_X56_X1_/ X3_X56_X1_W' X3_X56_X1_/  W' L='L_N' W='W_N' NF=1 AD='INT((NF+1)/2)
+ AS='INT((NF+2)/2) PD='2*INT((NF+1)/2) PS='2*INT((NF+2)/2) NRD='0.29 NRS='0.29 SA=0 SB=0 SD=0 MULT='N' M='N' 
*--------END___X3_X56_X1_XM1->W'
*--------BEGIN_X3_X56_X1_XM2->W'
XM2_X3_X56_X1 X3_X56_NET1 VDD X3_NET10 VDD X3_X56_X1_SKY130_FD_PR__PFET_01V8 X3_X56_X1_* X3_X56_X1_W/NF X3_X56_X1_* X3_X56_X1_0.29'
+ X3_X56_X1_* X3_X56_X1_W/NF X3_X56_X1_* X3_X56_X1_0.29' X3_X56_X1_* X3_X56_X1_(W/NF X3_X56_X1_+ X3_X56_X1_0.29)'
+ X3_X56_X1_* X3_X56_X1_(W/NF X3_X56_X1_+ X3_X56_X1_0.29)' X3_X56_X1_/ X3_X56_X1_W' X3_X56_X1_/  W' L='L_P' W='W_P' NF=1 AD='INT((NF+1)/2)
+ AS='INT((NF+2)/2) PD='2*INT((NF+1)/2) PS='2*INT((NF+2)/2) NRD='0.29 NRS='0.29 SA=0 SB=0 SD=0 MULT='N' M='N' 
*--------END___X3_X56_X1_XM2->W'
*--------END___X3_X56_X1->TRANSMISSION_GATE
*--------BEGIN_X3_X56_X2->TRANSMISSION_GATE
*.PININFO IN:B OUT:B EN:I EN_B:I
*--------BEGIN_X3_X56_X2_XM1->W'
XM1_X3_X56_X2 OUT32 X3_NET30 X3_X56_NET1 X3_VSS X3_X56_X2_SKY130_FD_PR__NFET_01V8 X3_X56_X2_* X3_X56_X2_W/NF X3_X56_X2_* X3_X56_X2_0.29'
+ X3_X56_X2_* X3_X56_X2_W/NF X3_X56_X2_* X3_X56_X2_0.29' X3_X56_X2_* X3_X56_X2_(W/NF X3_X56_X2_+ X3_X56_X2_0.29)'
+ X3_X56_X2_* X3_X56_X2_(W/NF X3_X56_X2_+ X3_X56_X2_0.29)' X3_X56_X2_/ X3_X56_X2_W' X3_X56_X2_/  W' L='L_N' W='W_N' NF=1 AD='INT((NF+1)/2)
+ AS='INT((NF+2)/2) PD='2*INT((NF+1)/2) PS='2*INT((NF+2)/2) NRD='0.29 NRS='0.29 SA=0 SB=0 SD=0 MULT='N' M='N' 
*--------END___X3_X56_X2_XM1->W'
*--------BEGIN_X3_X56_X2_XM2->W'
XM2_X3_X56_X2 OUT32 VDD X3_X56_NET1 VDD X3_X56_X2_SKY130_FD_PR__PFET_01V8 X3_X56_X2_* X3_X56_X2_W/NF X3_X56_X2_* X3_X56_X2_0.29'
+ X3_X56_X2_* X3_X56_X2_W/NF X3_X56_X2_* X3_X56_X2_0.29' X3_X56_X2_* X3_X56_X2_(W/NF X3_X56_X2_+ X3_X56_X2_0.29)'
+ X3_X56_X2_* X3_X56_X2_(W/NF X3_X56_X2_+ X3_X56_X2_0.29)' X3_X56_X2_/ X3_X56_X2_W' X3_X56_X2_/  W' L='L_P' W='W_P' NF=1 AD='INT((NF+1)/2)
+ AS='INT((NF+2)/2) PD='2*INT((NF+1)/2) PS='2*INT((NF+2)/2) NRD='0.29 NRS='0.29 SA=0 SB=0 SD=0 MULT='N' M='N' 
*--------END___X3_X56_X2_XM2->W'
*--------END___X3_X56_X2->TRANSMISSION_GATE
*--------BEGIN_X3_X56_XM1->W'
XM1_X3_X56 X3_X56_NET1 VDD X3_VSS X3_VSS X3_X56_SKY130_FD_PR__NFET_01V8 X3_X56_* X3_X56_W/NF X3_X56_* X3_X56_0.29'
+ X3_X56_* X3_X56_W/NF X3_X56_* X3_X56_0.29' X3_X56_* X3_X56_(W/NF X3_X56_+ X3_X56_0.29)' X3_X56_* X3_X56_(W/NF
+ X3_X56_+ X3_X56_0.29)' X3_X56_/ X3_X56_W' X3_X56_/  W' L=0.15 W=0.5 NF=1 AD='INT((NF+1)/2) AS='INT((NF+2)/2) PD='2*INT((NF+1)/2)
+ PS='2*INT((NF+2)/2) NRD='0.29 NRS='0.29 SA=0 SB=0 SD=0 MULT=1 M=1 
*--------END___X3_X56_XM1->W'
*--------END___X3_X56->SWITCH_5T
*--------BEGIN_X3_X57->SKY130_FD_SC_HD__INV_1
X57_X3 VDD X3_VGND X3_VNB X3_VPB X3_VPWR X3_NET30  SKY130_FD_SC_HD__INV_1
*--------END___X3_X57->SKY130_FD_SC_HD__INV_1
*--------BEGIN_X3_X2->TRANSMISSION_GATE
*.PININFO IN:B OUT:B EN:I EN_B:I
*--------BEGIN_X3_X2_XM1->W'
XM1_X3_X2 X3_NET11 VDD IN4 X3_VSS X3_X2_SKY130_FD_PR__NFET_01V8 X3_X2_* X3_X2_W/NF X3_X2_* X3_X2_0.29'
+ X3_X2_* X3_X2_W/NF X3_X2_* X3_X2_0.29' X3_X2_* X3_X2_(W/NF X3_X2_+ X3_X2_0.29)' X3_X2_* X3_X2_(W/NF X3_X2_+
+ X3_X2_0.29)' X3_X2_/ X3_X2_W' X3_X2_/  W' L='L_N' W='W_N' NF=1 AD='INT((NF+1)/2) AS='INT((NF+2)/2) PD='2*INT((NF+1)/2)
+ PS='2*INT((NF+2)/2) NRD='0.29 NRS='0.29 SA=0 SB=0 SD=0 MULT='N' M='N' 
*--------END___X3_X2_XM1->W'
*--------BEGIN_X3_X2_XM2->W'
XM2_X3_X2 X3_NET11 GND IN4 VDD X3_X2_SKY130_FD_PR__PFET_01V8 X3_X2_* X3_X2_W/NF X3_X2_* X3_X2_0.29' X3_X2_*
+ X3_X2_W/NF X3_X2_* X3_X2_0.29' X3_X2_* X3_X2_(W/NF X3_X2_+ X3_X2_0.29)' X3_X2_* X3_X2_(W/NF X3_X2_+ X3_X2_0.29)' X3_X2_/ X3_X2_W'
+ X3_X2_/  W' L='L_P' W='W_P' NF=1 AD='INT((NF+1)/2) AS='INT((NF+2)/2) PD='2*INT((NF+1)/2) PS='2*INT((NF+2)/2) NRD='0.29
+ NRS='0.29 SA=0 SB=0 SD=0 MULT='N' M='N' 
*--------END___X3_X2_XM2->W'
*--------END___X3_X2->TRANSMISSION_GATE
*--------BEGIN_X3_X3->SWITCH_5T
*.PININFO IN:B OUT:B EN:I EN_B:I
*--------BEGIN_X3_X3_X1->TRANSMISSION_GATE
*.PININFO IN:B OUT:B EN:I EN_B:I
*--------BEGIN_X3_X3_X1_XM1->W'
XM1_X3_X3_X1 X3_X3_NET1 X3_NET31 X3_NET11 X3_VSS X3_X3_X1_SKY130_FD_PR__NFET_01V8 X3_X3_X1_* X3_X3_X1_W/NF X3_X3_X1_* X3_X3_X1_0.29'
+ X3_X3_X1_* X3_X3_X1_W/NF X3_X3_X1_* X3_X3_X1_0.29' X3_X3_X1_* X3_X3_X1_(W/NF X3_X3_X1_+ X3_X3_X1_0.29)'
+ X3_X3_X1_* X3_X3_X1_(W/NF X3_X3_X1_+ X3_X3_X1_0.29)' X3_X3_X1_/ X3_X3_X1_W' X3_X3_X1_/  W' L='L_N' W='W_N' NF=1 AD='INT((NF+1)/2)
+ AS='INT((NF+2)/2) PD='2*INT((NF+1)/2) PS='2*INT((NF+2)/2) NRD='0.29 NRS='0.29 SA=0 SB=0 SD=0 MULT='N' M='N' 
*--------END___X3_X3_X1_XM1->W'
*--------BEGIN_X3_X3_X1_XM2->W'
XM2_X3_X3_X1 X3_X3_NET1 VDD X3_NET11 VDD X3_X3_X1_SKY130_FD_PR__PFET_01V8 X3_X3_X1_* X3_X3_X1_W/NF X3_X3_X1_* X3_X3_X1_0.29'
+ X3_X3_X1_* X3_X3_X1_W/NF X3_X3_X1_* X3_X3_X1_0.29' X3_X3_X1_* X3_X3_X1_(W/NF X3_X3_X1_+ X3_X3_X1_0.29)'
+ X3_X3_X1_* X3_X3_X1_(W/NF X3_X3_X1_+ X3_X3_X1_0.29)' X3_X3_X1_/ X3_X3_X1_W' X3_X3_X1_/  W' L='L_P' W='W_P' NF=1 AD='INT((NF+1)/2)
+ AS='INT((NF+2)/2) PD='2*INT((NF+1)/2) PS='2*INT((NF+2)/2) NRD='0.29 NRS='0.29 SA=0 SB=0 SD=0 MULT='N' M='N' 
*--------END___X3_X3_X1_XM2->W'
*--------END___X3_X3_X1->TRANSMISSION_GATE
*--------BEGIN_X3_X3_X2->TRANSMISSION_GATE
*.PININFO IN:B OUT:B EN:I EN_B:I
*--------BEGIN_X3_X3_X2_XM1->W'
XM1_X3_X3_X2 OUT32 X3_NET31 X3_X3_NET1 X3_VSS X3_X3_X2_SKY130_FD_PR__NFET_01V8 X3_X3_X2_* X3_X3_X2_W/NF X3_X3_X2_* X3_X3_X2_0.29'
+ X3_X3_X2_* X3_X3_X2_W/NF X3_X3_X2_* X3_X3_X2_0.29' X3_X3_X2_* X3_X3_X2_(W/NF X3_X3_X2_+ X3_X3_X2_0.29)'
+ X3_X3_X2_* X3_X3_X2_(W/NF X3_X3_X2_+ X3_X3_X2_0.29)' X3_X3_X2_/ X3_X3_X2_W' X3_X3_X2_/  W' L='L_N' W='W_N' NF=1 AD='INT((NF+1)/2)
+ AS='INT((NF+2)/2) PD='2*INT((NF+1)/2) PS='2*INT((NF+2)/2) NRD='0.29 NRS='0.29 SA=0 SB=0 SD=0 MULT='N' M='N' 
*--------END___X3_X3_X2_XM1->W'
*--------BEGIN_X3_X3_X2_XM2->W'
XM2_X3_X3_X2 OUT32 VDD X3_X3_NET1 VDD X3_X3_X2_SKY130_FD_PR__PFET_01V8 X3_X3_X2_* X3_X3_X2_W/NF X3_X3_X2_* X3_X3_X2_0.29'
+ X3_X3_X2_* X3_X3_X2_W/NF X3_X3_X2_* X3_X3_X2_0.29' X3_X3_X2_* X3_X3_X2_(W/NF X3_X3_X2_+ X3_X3_X2_0.29)'
+ X3_X3_X2_* X3_X3_X2_(W/NF X3_X3_X2_+ X3_X3_X2_0.29)' X3_X3_X2_/ X3_X3_X2_W' X3_X3_X2_/  W' L='L_P' W='W_P' NF=1 AD='INT((NF+1)/2)
+ AS='INT((NF+2)/2) PD='2*INT((NF+1)/2) PS='2*INT((NF+2)/2) NRD='0.29 NRS='0.29 SA=0 SB=0 SD=0 MULT='N' M='N' 
*--------END___X3_X3_X2_XM2->W'
*--------END___X3_X3_X2->TRANSMISSION_GATE
*--------BEGIN_X3_X3_XM1->W'
XM1_X3_X3 X3_X3_NET1 VDD X3_VSS X3_VSS X3_X3_SKY130_FD_PR__NFET_01V8 X3_X3_* X3_X3_W/NF X3_X3_* X3_X3_0.29'
+ X3_X3_* X3_X3_W/NF X3_X3_* X3_X3_0.29' X3_X3_* X3_X3_(W/NF X3_X3_+ X3_X3_0.29)' X3_X3_* X3_X3_(W/NF X3_X3_+
+ X3_X3_0.29)' X3_X3_/ X3_X3_W' X3_X3_/  W' L=0.15 W=0.5 NF=1 AD='INT((NF+1)/2) AS='INT((NF+2)/2) PD='2*INT((NF+1)/2)
+ PS='2*INT((NF+2)/2) NRD='0.29 NRS='0.29 SA=0 SB=0 SD=0 MULT=1 M=1 
*--------END___X3_X3_XM1->W'
*--------END___X3_X3->SWITCH_5T
*--------BEGIN_X3_X4->SKY130_FD_SC_HD__INV_1
X4_X3 VDD X3_VGND X3_VNB X3_VPB X3_VPWR X3_NET31  SKY130_FD_SC_HD__INV_1
*--------END___X3_X4->SKY130_FD_SC_HD__INV_1
*--------BEGIN_X3_X5->TRANSMISSION_GATE
*.PININFO IN:B OUT:B EN:I EN_B:I
*--------BEGIN_X3_X5_XM1->W'
XM1_X3_X5 X3_NET12 VDD IN5 X3_VSS X3_X5_SKY130_FD_PR__NFET_01V8 X3_X5_* X3_X5_W/NF X3_X5_* X3_X5_0.29'
+ X3_X5_* X3_X5_W/NF X3_X5_* X3_X5_0.29' X3_X5_* X3_X5_(W/NF X3_X5_+ X3_X5_0.29)' X3_X5_* X3_X5_(W/NF X3_X5_+
+ X3_X5_0.29)' X3_X5_/ X3_X5_W' X3_X5_/  W' L='L_N' W='W_N' NF=1 AD='INT((NF+1)/2) AS='INT((NF+2)/2) PD='2*INT((NF+1)/2)
+ PS='2*INT((NF+2)/2) NRD='0.29 NRS='0.29 SA=0 SB=0 SD=0 MULT='N' M='N' 
*--------END___X3_X5_XM1->W'
*--------BEGIN_X3_X5_XM2->W'
XM2_X3_X5 X3_NET12 GND IN5 VDD X3_X5_SKY130_FD_PR__PFET_01V8 X3_X5_* X3_X5_W/NF X3_X5_* X3_X5_0.29' X3_X5_*
+ X3_X5_W/NF X3_X5_* X3_X5_0.29' X3_X5_* X3_X5_(W/NF X3_X5_+ X3_X5_0.29)' X3_X5_* X3_X5_(W/NF X3_X5_+ X3_X5_0.29)' X3_X5_/ X3_X5_W'
+ X3_X5_/  W' L='L_P' W='W_P' NF=1 AD='INT((NF+1)/2) AS='INT((NF+2)/2) PD='2*INT((NF+1)/2) PS='2*INT((NF+2)/2) NRD='0.29
+ NRS='0.29 SA=0 SB=0 SD=0 MULT='N' M='N' 
*--------END___X3_X5_XM2->W'
*--------END___X3_X5->TRANSMISSION_GATE
*--------BEGIN_X3_X6->SWITCH_5T
*.PININFO IN:B OUT:B EN:I EN_B:I
*--------BEGIN_X3_X6_X1->TRANSMISSION_GATE
*.PININFO IN:B OUT:B EN:I EN_B:I
*--------BEGIN_X3_X6_X1_XM1->W'
XM1_X3_X6_X1 X3_X6_NET1 X3_NET32 X3_NET12 X3_VSS X3_X6_X1_SKY130_FD_PR__NFET_01V8 X3_X6_X1_* X3_X6_X1_W/NF X3_X6_X1_* X3_X6_X1_0.29'
+ X3_X6_X1_* X3_X6_X1_W/NF X3_X6_X1_* X3_X6_X1_0.29' X3_X6_X1_* X3_X6_X1_(W/NF X3_X6_X1_+ X3_X6_X1_0.29)'
+ X3_X6_X1_* X3_X6_X1_(W/NF X3_X6_X1_+ X3_X6_X1_0.29)' X3_X6_X1_/ X3_X6_X1_W' X3_X6_X1_/  W' L='L_N' W='W_N' NF=1 AD='INT((NF+1)/2)
+ AS='INT((NF+2)/2) PD='2*INT((NF+1)/2) PS='2*INT((NF+2)/2) NRD='0.29 NRS='0.29 SA=0 SB=0 SD=0 MULT='N' M='N' 
*--------END___X3_X6_X1_XM1->W'
*--------BEGIN_X3_X6_X1_XM2->W'
XM2_X3_X6_X1 X3_X6_NET1 VDD X3_NET12 VDD X3_X6_X1_SKY130_FD_PR__PFET_01V8 X3_X6_X1_* X3_X6_X1_W/NF X3_X6_X1_* X3_X6_X1_0.29'
+ X3_X6_X1_* X3_X6_X1_W/NF X3_X6_X1_* X3_X6_X1_0.29' X3_X6_X1_* X3_X6_X1_(W/NF X3_X6_X1_+ X3_X6_X1_0.29)'
+ X3_X6_X1_* X3_X6_X1_(W/NF X3_X6_X1_+ X3_X6_X1_0.29)' X3_X6_X1_/ X3_X6_X1_W' X3_X6_X1_/  W' L='L_P' W='W_P' NF=1 AD='INT((NF+1)/2)
+ AS='INT((NF+2)/2) PD='2*INT((NF+1)/2) PS='2*INT((NF+2)/2) NRD='0.29 NRS='0.29 SA=0 SB=0 SD=0 MULT='N' M='N' 
*--------END___X3_X6_X1_XM2->W'
*--------END___X3_X6_X1->TRANSMISSION_GATE
*--------BEGIN_X3_X6_X2->TRANSMISSION_GATE
*.PININFO IN:B OUT:B EN:I EN_B:I
*--------BEGIN_X3_X6_X2_XM1->W'
XM1_X3_X6_X2 OUT32 X3_NET32 X3_X6_NET1 X3_VSS X3_X6_X2_SKY130_FD_PR__NFET_01V8 X3_X6_X2_* X3_X6_X2_W/NF X3_X6_X2_* X3_X6_X2_0.29'
+ X3_X6_X2_* X3_X6_X2_W/NF X3_X6_X2_* X3_X6_X2_0.29' X3_X6_X2_* X3_X6_X2_(W/NF X3_X6_X2_+ X3_X6_X2_0.29)'
+ X3_X6_X2_* X3_X6_X2_(W/NF X3_X6_X2_+ X3_X6_X2_0.29)' X3_X6_X2_/ X3_X6_X2_W' X3_X6_X2_/  W' L='L_N' W='W_N' NF=1 AD='INT((NF+1)/2)
+ AS='INT((NF+2)/2) PD='2*INT((NF+1)/2) PS='2*INT((NF+2)/2) NRD='0.29 NRS='0.29 SA=0 SB=0 SD=0 MULT='N' M='N' 
*--------END___X3_X6_X2_XM1->W'
*--------BEGIN_X3_X6_X2_XM2->W'
XM2_X3_X6_X2 OUT32 VDD X3_X6_NET1 VDD X3_X6_X2_SKY130_FD_PR__PFET_01V8 X3_X6_X2_* X3_X6_X2_W/NF X3_X6_X2_* X3_X6_X2_0.29'
+ X3_X6_X2_* X3_X6_X2_W/NF X3_X6_X2_* X3_X6_X2_0.29' X3_X6_X2_* X3_X6_X2_(W/NF X3_X6_X2_+ X3_X6_X2_0.29)'
+ X3_X6_X2_* X3_X6_X2_(W/NF X3_X6_X2_+ X3_X6_X2_0.29)' X3_X6_X2_/ X3_X6_X2_W' X3_X6_X2_/  W' L='L_P' W='W_P' NF=1 AD='INT((NF+1)/2)
+ AS='INT((NF+2)/2) PD='2*INT((NF+1)/2) PS='2*INT((NF+2)/2) NRD='0.29 NRS='0.29 SA=0 SB=0 SD=0 MULT='N' M='N' 
*--------END___X3_X6_X2_XM2->W'
*--------END___X3_X6_X2->TRANSMISSION_GATE
*--------BEGIN_X3_X6_XM1->W'
XM1_X3_X6 X3_X6_NET1 VDD X3_VSS X3_VSS X3_X6_SKY130_FD_PR__NFET_01V8 X3_X6_* X3_X6_W/NF X3_X6_* X3_X6_0.29'
+ X3_X6_* X3_X6_W/NF X3_X6_* X3_X6_0.29' X3_X6_* X3_X6_(W/NF X3_X6_+ X3_X6_0.29)' X3_X6_* X3_X6_(W/NF X3_X6_+
+ X3_X6_0.29)' X3_X6_/ X3_X6_W' X3_X6_/  W' L=0.15 W=0.5 NF=1 AD='INT((NF+1)/2) AS='INT((NF+2)/2) PD='2*INT((NF+1)/2)
+ PS='2*INT((NF+2)/2) NRD='0.29 NRS='0.29 SA=0 SB=0 SD=0 MULT=1 M=1 
*--------END___X3_X6_XM1->W'
*--------END___X3_X6->SWITCH_5T
*--------BEGIN_X3_X7->SKY130_FD_SC_HD__INV_1
X7_X3 VDD X3_VGND X3_VNB X3_VPB X3_VPWR X3_NET32  SKY130_FD_SC_HD__INV_1
*--------END___X3_X7->SKY130_FD_SC_HD__INV_1
*--------BEGIN_X3_X8->TRANSMISSION_GATE
*.PININFO IN:B OUT:B EN:I EN_B:I
*--------BEGIN_X3_X8_XM1->W'
XM1_X3_X8 X3_NET13 VDD IN6 X3_VSS X3_X8_SKY130_FD_PR__NFET_01V8 X3_X8_* X3_X8_W/NF X3_X8_* X3_X8_0.29'
+ X3_X8_* X3_X8_W/NF X3_X8_* X3_X8_0.29' X3_X8_* X3_X8_(W/NF X3_X8_+ X3_X8_0.29)' X3_X8_* X3_X8_(W/NF X3_X8_+
+ X3_X8_0.29)' X3_X8_/ X3_X8_W' X3_X8_/  W' L='L_N' W='W_N' NF=1 AD='INT((NF+1)/2) AS='INT((NF+2)/2) PD='2*INT((NF+1)/2)
+ PS='2*INT((NF+2)/2) NRD='0.29 NRS='0.29 SA=0 SB=0 SD=0 MULT='N' M='N' 
*--------END___X3_X8_XM1->W'
*--------BEGIN_X3_X8_XM2->W'
XM2_X3_X8 X3_NET13 GND IN6 VDD X3_X8_SKY130_FD_PR__PFET_01V8 X3_X8_* X3_X8_W/NF X3_X8_* X3_X8_0.29' X3_X8_*
+ X3_X8_W/NF X3_X8_* X3_X8_0.29' X3_X8_* X3_X8_(W/NF X3_X8_+ X3_X8_0.29)' X3_X8_* X3_X8_(W/NF X3_X8_+ X3_X8_0.29)' X3_X8_/ X3_X8_W'
+ X3_X8_/  W' L='L_P' W='W_P' NF=1 AD='INT((NF+1)/2) AS='INT((NF+2)/2) PD='2*INT((NF+1)/2) PS='2*INT((NF+2)/2) NRD='0.29
+ NRS='0.29 SA=0 SB=0 SD=0 MULT='N' M='N' 
*--------END___X3_X8_XM2->W'
*--------END___X3_X8->TRANSMISSION_GATE
*--------BEGIN_X3_X9->SWITCH_5T
*.PININFO IN:B OUT:B EN:I EN_B:I
*--------BEGIN_X3_X9_X1->TRANSMISSION_GATE
*.PININFO IN:B OUT:B EN:I EN_B:I
*--------BEGIN_X3_X9_X1_XM1->W'
XM1_X3_X9_X1 X3_X9_NET1 X3_NET33 X3_NET13 X3_VSS X3_X9_X1_SKY130_FD_PR__NFET_01V8 X3_X9_X1_* X3_X9_X1_W/NF X3_X9_X1_* X3_X9_X1_0.29'
+ X3_X9_X1_* X3_X9_X1_W/NF X3_X9_X1_* X3_X9_X1_0.29' X3_X9_X1_* X3_X9_X1_(W/NF X3_X9_X1_+ X3_X9_X1_0.29)'
+ X3_X9_X1_* X3_X9_X1_(W/NF X3_X9_X1_+ X3_X9_X1_0.29)' X3_X9_X1_/ X3_X9_X1_W' X3_X9_X1_/  W' L='L_N' W='W_N' NF=1 AD='INT((NF+1)/2)
+ AS='INT((NF+2)/2) PD='2*INT((NF+1)/2) PS='2*INT((NF+2)/2) NRD='0.29 NRS='0.29 SA=0 SB=0 SD=0 MULT='N' M='N' 
*--------END___X3_X9_X1_XM1->W'
*--------BEGIN_X3_X9_X1_XM2->W'
XM2_X3_X9_X1 X3_X9_NET1 VDD X3_NET13 VDD X3_X9_X1_SKY130_FD_PR__PFET_01V8 X3_X9_X1_* X3_X9_X1_W/NF X3_X9_X1_* X3_X9_X1_0.29'
+ X3_X9_X1_* X3_X9_X1_W/NF X3_X9_X1_* X3_X9_X1_0.29' X3_X9_X1_* X3_X9_X1_(W/NF X3_X9_X1_+ X3_X9_X1_0.29)'
+ X3_X9_X1_* X3_X9_X1_(W/NF X3_X9_X1_+ X3_X9_X1_0.29)' X3_X9_X1_/ X3_X9_X1_W' X3_X9_X1_/  W' L='L_P' W='W_P' NF=1 AD='INT((NF+1)/2)
+ AS='INT((NF+2)/2) PD='2*INT((NF+1)/2) PS='2*INT((NF+2)/2) NRD='0.29 NRS='0.29 SA=0 SB=0 SD=0 MULT='N' M='N' 
*--------END___X3_X9_X1_XM2->W'
*--------END___X3_X9_X1->TRANSMISSION_GATE
*--------BEGIN_X3_X9_X2->TRANSMISSION_GATE
*.PININFO IN:B OUT:B EN:I EN_B:I
*--------BEGIN_X3_X9_X2_XM1->W'
XM1_X3_X9_X2 OUT32 X3_NET33 X3_X9_NET1 X3_VSS X3_X9_X2_SKY130_FD_PR__NFET_01V8 X3_X9_X2_* X3_X9_X2_W/NF X3_X9_X2_* X3_X9_X2_0.29'
+ X3_X9_X2_* X3_X9_X2_W/NF X3_X9_X2_* X3_X9_X2_0.29' X3_X9_X2_* X3_X9_X2_(W/NF X3_X9_X2_+ X3_X9_X2_0.29)'
+ X3_X9_X2_* X3_X9_X2_(W/NF X3_X9_X2_+ X3_X9_X2_0.29)' X3_X9_X2_/ X3_X9_X2_W' X3_X9_X2_/  W' L='L_N' W='W_N' NF=1 AD='INT((NF+1)/2)
+ AS='INT((NF+2)/2) PD='2*INT((NF+1)/2) PS='2*INT((NF+2)/2) NRD='0.29 NRS='0.29 SA=0 SB=0 SD=0 MULT='N' M='N' 
*--------END___X3_X9_X2_XM1->W'
*--------BEGIN_X3_X9_X2_XM2->W'
XM2_X3_X9_X2 OUT32 VDD X3_X9_NET1 VDD X3_X9_X2_SKY130_FD_PR__PFET_01V8 X3_X9_X2_* X3_X9_X2_W/NF X3_X9_X2_* X3_X9_X2_0.29'
+ X3_X9_X2_* X3_X9_X2_W/NF X3_X9_X2_* X3_X9_X2_0.29' X3_X9_X2_* X3_X9_X2_(W/NF X3_X9_X2_+ X3_X9_X2_0.29)'
+ X3_X9_X2_* X3_X9_X2_(W/NF X3_X9_X2_+ X3_X9_X2_0.29)' X3_X9_X2_/ X3_X9_X2_W' X3_X9_X2_/  W' L='L_P' W='W_P' NF=1 AD='INT((NF+1)/2)
+ AS='INT((NF+2)/2) PD='2*INT((NF+1)/2) PS='2*INT((NF+2)/2) NRD='0.29 NRS='0.29 SA=0 SB=0 SD=0 MULT='N' M='N' 
*--------END___X3_X9_X2_XM2->W'
*--------END___X3_X9_X2->TRANSMISSION_GATE
*--------BEGIN_X3_X9_XM1->W'
XM1_X3_X9 X3_X9_NET1 VDD X3_VSS X3_VSS X3_X9_SKY130_FD_PR__NFET_01V8 X3_X9_* X3_X9_W/NF X3_X9_* X3_X9_0.29'
+ X3_X9_* X3_X9_W/NF X3_X9_* X3_X9_0.29' X3_X9_* X3_X9_(W/NF X3_X9_+ X3_X9_0.29)' X3_X9_* X3_X9_(W/NF X3_X9_+
+ X3_X9_0.29)' X3_X9_/ X3_X9_W' X3_X9_/  W' L=0.15 W=0.5 NF=1 AD='INT((NF+1)/2) AS='INT((NF+2)/2) PD='2*INT((NF+1)/2)
+ PS='2*INT((NF+2)/2) NRD='0.29 NRS='0.29 SA=0 SB=0 SD=0 MULT=1 M=1 
*--------END___X3_X9_XM1->W'
*--------END___X3_X9->SWITCH_5T
*--------BEGIN_X3_X10->SKY130_FD_SC_HD__INV_1
X10_X3 VDD X3_VGND X3_VNB X3_VPB X3_VPWR X3_NET33  SKY130_FD_SC_HD__INV_1
*--------END___X3_X10->SKY130_FD_SC_HD__INV_1
*--------BEGIN_X3_X11->TRANSMISSION_GATE
*.PININFO IN:B OUT:B EN:I EN_B:I
*--------BEGIN_X3_X11_XM1->W'
XM1_X3_X11 X3_NET14 VDD IN7 X3_VSS X3_X11_SKY130_FD_PR__NFET_01V8 X3_X11_* X3_X11_W/NF X3_X11_* X3_X11_0.29'
+ X3_X11_* X3_X11_W/NF X3_X11_* X3_X11_0.29' X3_X11_* X3_X11_(W/NF X3_X11_+ X3_X11_0.29)' X3_X11_* X3_X11_(W/NF
+ X3_X11_+ X3_X11_0.29)' X3_X11_/ X3_X11_W' X3_X11_/  W' L='L_N' W='W_N' NF=1 AD='INT((NF+1)/2) AS='INT((NF+2)/2) PD='2*INT((NF+1)/2)
+ PS='2*INT((NF+2)/2) NRD='0.29 NRS='0.29 SA=0 SB=0 SD=0 MULT='N' M='N' 
*--------END___X3_X11_XM1->W'
*--------BEGIN_X3_X11_XM2->W'
XM2_X3_X11 X3_NET14 GND IN7 VDD X3_X11_SKY130_FD_PR__PFET_01V8 X3_X11_* X3_X11_W/NF X3_X11_* X3_X11_0.29'
+ X3_X11_* X3_X11_W/NF X3_X11_* X3_X11_0.29' X3_X11_* X3_X11_(W/NF X3_X11_+ X3_X11_0.29)' X3_X11_* X3_X11_(W/NF
+ X3_X11_+ X3_X11_0.29)' X3_X11_/ X3_X11_W' X3_X11_/  W' L='L_P' W='W_P' NF=1 AD='INT((NF+1)/2) AS='INT((NF+2)/2) PD='2*INT((NF+1)/2)
+ PS='2*INT((NF+2)/2) NRD='0.29 NRS='0.29 SA=0 SB=0 SD=0 MULT='N' M='N' 
*--------END___X3_X11_XM2->W'
*--------END___X3_X11->TRANSMISSION_GATE
*--------BEGIN_X3_X12->SWITCH_5T
*.PININFO IN:B OUT:B EN:I EN_B:I
*--------BEGIN_X3_X12_X1->TRANSMISSION_GATE
*.PININFO IN:B OUT:B EN:I EN_B:I
*--------BEGIN_X3_X12_X1_XM1->W'
XM1_X3_X12_X1 X3_X12_NET1 X3_NET34 X3_NET14 X3_VSS X3_X12_X1_SKY130_FD_PR__NFET_01V8 X3_X12_X1_* X3_X12_X1_W/NF X3_X12_X1_* X3_X12_X1_0.29'
+ X3_X12_X1_* X3_X12_X1_W/NF X3_X12_X1_* X3_X12_X1_0.29' X3_X12_X1_* X3_X12_X1_(W/NF X3_X12_X1_+ X3_X12_X1_0.29)'
+ X3_X12_X1_* X3_X12_X1_(W/NF X3_X12_X1_+ X3_X12_X1_0.29)' X3_X12_X1_/ X3_X12_X1_W' X3_X12_X1_/  W' L='L_N' W='W_N' NF=1 AD='INT((NF+1)/2)
+ AS='INT((NF+2)/2) PD='2*INT((NF+1)/2) PS='2*INT((NF+2)/2) NRD='0.29 NRS='0.29 SA=0 SB=0 SD=0 MULT='N' M='N' 
*--------END___X3_X12_X1_XM1->W'
*--------BEGIN_X3_X12_X1_XM2->W'
XM2_X3_X12_X1 X3_X12_NET1 VDD X3_NET14 VDD X3_X12_X1_SKY130_FD_PR__PFET_01V8 X3_X12_X1_* X3_X12_X1_W/NF X3_X12_X1_* X3_X12_X1_0.29'
+ X3_X12_X1_* X3_X12_X1_W/NF X3_X12_X1_* X3_X12_X1_0.29' X3_X12_X1_* X3_X12_X1_(W/NF X3_X12_X1_+ X3_X12_X1_0.29)'
+ X3_X12_X1_* X3_X12_X1_(W/NF X3_X12_X1_+ X3_X12_X1_0.29)' X3_X12_X1_/ X3_X12_X1_W' X3_X12_X1_/  W' L='L_P' W='W_P' NF=1 AD='INT((NF+1)/2)
+ AS='INT((NF+2)/2) PD='2*INT((NF+1)/2) PS='2*INT((NF+2)/2) NRD='0.29 NRS='0.29 SA=0 SB=0 SD=0 MULT='N' M='N' 
*--------END___X3_X12_X1_XM2->W'
*--------END___X3_X12_X1->TRANSMISSION_GATE
*--------BEGIN_X3_X12_X2->TRANSMISSION_GATE
*.PININFO IN:B OUT:B EN:I EN_B:I
*--------BEGIN_X3_X12_X2_XM1->W'
XM1_X3_X12_X2 OUT32 X3_NET34 X3_X12_NET1 X3_VSS X3_X12_X2_SKY130_FD_PR__NFET_01V8 X3_X12_X2_* X3_X12_X2_W/NF X3_X12_X2_* X3_X12_X2_0.29'
+ X3_X12_X2_* X3_X12_X2_W/NF X3_X12_X2_* X3_X12_X2_0.29' X3_X12_X2_* X3_X12_X2_(W/NF X3_X12_X2_+ X3_X12_X2_0.29)'
+ X3_X12_X2_* X3_X12_X2_(W/NF X3_X12_X2_+ X3_X12_X2_0.29)' X3_X12_X2_/ X3_X12_X2_W' X3_X12_X2_/  W' L='L_N' W='W_N' NF=1 AD='INT((NF+1)/2)
+ AS='INT((NF+2)/2) PD='2*INT((NF+1)/2) PS='2*INT((NF+2)/2) NRD='0.29 NRS='0.29 SA=0 SB=0 SD=0 MULT='N' M='N' 
*--------END___X3_X12_X2_XM1->W'
*--------BEGIN_X3_X12_X2_XM2->W'
XM2_X3_X12_X2 OUT32 VDD X3_X12_NET1 VDD X3_X12_X2_SKY130_FD_PR__PFET_01V8 X3_X12_X2_* X3_X12_X2_W/NF X3_X12_X2_* X3_X12_X2_0.29'
+ X3_X12_X2_* X3_X12_X2_W/NF X3_X12_X2_* X3_X12_X2_0.29' X3_X12_X2_* X3_X12_X2_(W/NF X3_X12_X2_+ X3_X12_X2_0.29)'
+ X3_X12_X2_* X3_X12_X2_(W/NF X3_X12_X2_+ X3_X12_X2_0.29)' X3_X12_X2_/ X3_X12_X2_W' X3_X12_X2_/  W' L='L_P' W='W_P' NF=1 AD='INT((NF+1)/2)
+ AS='INT((NF+2)/2) PD='2*INT((NF+1)/2) PS='2*INT((NF+2)/2) NRD='0.29 NRS='0.29 SA=0 SB=0 SD=0 MULT='N' M='N' 
*--------END___X3_X12_X2_XM2->W'
*--------END___X3_X12_X2->TRANSMISSION_GATE
*--------BEGIN_X3_X12_XM1->W'
XM1_X3_X12 X3_X12_NET1 VDD X3_VSS X3_VSS X3_X12_SKY130_FD_PR__NFET_01V8 X3_X12_* X3_X12_W/NF X3_X12_* X3_X12_0.29'
+ X3_X12_* X3_X12_W/NF X3_X12_* X3_X12_0.29' X3_X12_* X3_X12_(W/NF X3_X12_+ X3_X12_0.29)' X3_X12_* X3_X12_(W/NF
+ X3_X12_+ X3_X12_0.29)' X3_X12_/ X3_X12_W' X3_X12_/  W' L=0.15 W=0.5 NF=1 AD='INT((NF+1)/2) AS='INT((NF+2)/2) PD='2*INT((NF+1)/2)
+ PS='2*INT((NF+2)/2) NRD='0.29 NRS='0.29 SA=0 SB=0 SD=0 MULT=1 M=1 
*--------END___X3_X12_XM1->W'
*--------END___X3_X12->SWITCH_5T
*--------BEGIN_X3_X13->SKY130_FD_SC_HD__INV_1
X13_X3 VDD X3_VGND X3_VNB X3_VPB X3_VPWR X3_NET34  SKY130_FD_SC_HD__INV_1
*--------END___X3_X13->SKY130_FD_SC_HD__INV_1
*--------BEGIN_X3_X14->TRANSMISSION_GATE
*.PININFO IN:B OUT:B EN:I EN_B:I
*--------BEGIN_X3_X14_XM1->W'
XM1_X3_X14 X3_NET15 VDD IN8 X3_VSS X3_X14_SKY130_FD_PR__NFET_01V8 X3_X14_* X3_X14_W/NF X3_X14_* X3_X14_0.29'
+ X3_X14_* X3_X14_W/NF X3_X14_* X3_X14_0.29' X3_X14_* X3_X14_(W/NF X3_X14_+ X3_X14_0.29)' X3_X14_* X3_X14_(W/NF
+ X3_X14_+ X3_X14_0.29)' X3_X14_/ X3_X14_W' X3_X14_/  W' L='L_N' W='W_N' NF=1 AD='INT((NF+1)/2) AS='INT((NF+2)/2) PD='2*INT((NF+1)/2)
+ PS='2*INT((NF+2)/2) NRD='0.29 NRS='0.29 SA=0 SB=0 SD=0 MULT='N' M='N' 
*--------END___X3_X14_XM1->W'
*--------BEGIN_X3_X14_XM2->W'
XM2_X3_X14 X3_NET15 GND IN8 VDD X3_X14_SKY130_FD_PR__PFET_01V8 X3_X14_* X3_X14_W/NF X3_X14_* X3_X14_0.29'
+ X3_X14_* X3_X14_W/NF X3_X14_* X3_X14_0.29' X3_X14_* X3_X14_(W/NF X3_X14_+ X3_X14_0.29)' X3_X14_* X3_X14_(W/NF
+ X3_X14_+ X3_X14_0.29)' X3_X14_/ X3_X14_W' X3_X14_/  W' L='L_P' W='W_P' NF=1 AD='INT((NF+1)/2) AS='INT((NF+2)/2) PD='2*INT((NF+1)/2)
+ PS='2*INT((NF+2)/2) NRD='0.29 NRS='0.29 SA=0 SB=0 SD=0 MULT='N' M='N' 
*--------END___X3_X14_XM2->W'
*--------END___X3_X14->TRANSMISSION_GATE
*--------BEGIN_X3_X15->SWITCH_5T
*.PININFO IN:B OUT:B EN:I EN_B:I
*--------BEGIN_X3_X15_X1->TRANSMISSION_GATE
*.PININFO IN:B OUT:B EN:I EN_B:I
*--------BEGIN_X3_X15_X1_XM1->W'
XM1_X3_X15_X1 X3_X15_NET1 X3_NET35 X3_NET15 X3_VSS X3_X15_X1_SKY130_FD_PR__NFET_01V8 X3_X15_X1_* X3_X15_X1_W/NF X3_X15_X1_* X3_X15_X1_0.29'
+ X3_X15_X1_* X3_X15_X1_W/NF X3_X15_X1_* X3_X15_X1_0.29' X3_X15_X1_* X3_X15_X1_(W/NF X3_X15_X1_+ X3_X15_X1_0.29)'
+ X3_X15_X1_* X3_X15_X1_(W/NF X3_X15_X1_+ X3_X15_X1_0.29)' X3_X15_X1_/ X3_X15_X1_W' X3_X15_X1_/  W' L='L_N' W='W_N' NF=1 AD='INT((NF+1)/2)
+ AS='INT((NF+2)/2) PD='2*INT((NF+1)/2) PS='2*INT((NF+2)/2) NRD='0.29 NRS='0.29 SA=0 SB=0 SD=0 MULT='N' M='N' 
*--------END___X3_X15_X1_XM1->W'
*--------BEGIN_X3_X15_X1_XM2->W'
XM2_X3_X15_X1 X3_X15_NET1 GND X3_NET15 VDD X3_X15_X1_SKY130_FD_PR__PFET_01V8 X3_X15_X1_* X3_X15_X1_W/NF X3_X15_X1_* X3_X15_X1_0.29'
+ X3_X15_X1_* X3_X15_X1_W/NF X3_X15_X1_* X3_X15_X1_0.29' X3_X15_X1_* X3_X15_X1_(W/NF X3_X15_X1_+ X3_X15_X1_0.29)'
+ X3_X15_X1_* X3_X15_X1_(W/NF X3_X15_X1_+ X3_X15_X1_0.29)' X3_X15_X1_/ X3_X15_X1_W' X3_X15_X1_/  W' L='L_P' W='W_P' NF=1 AD='INT((NF+1)/2)
+ AS='INT((NF+2)/2) PD='2*INT((NF+1)/2) PS='2*INT((NF+2)/2) NRD='0.29 NRS='0.29 SA=0 SB=0 SD=0 MULT='N' M='N' 
*--------END___X3_X15_X1_XM2->W'
*--------END___X3_X15_X1->TRANSMISSION_GATE
*--------BEGIN_X3_X15_X2->TRANSMISSION_GATE
*.PININFO IN:B OUT:B EN:I EN_B:I
*--------BEGIN_X3_X15_X2_XM1->W'
XM1_X3_X15_X2 OUT32 X3_NET35 X3_X15_NET1 X3_VSS X3_X15_X2_SKY130_FD_PR__NFET_01V8 X3_X15_X2_* X3_X15_X2_W/NF X3_X15_X2_* X3_X15_X2_0.29'
+ X3_X15_X2_* X3_X15_X2_W/NF X3_X15_X2_* X3_X15_X2_0.29' X3_X15_X2_* X3_X15_X2_(W/NF X3_X15_X2_+ X3_X15_X2_0.29)'
+ X3_X15_X2_* X3_X15_X2_(W/NF X3_X15_X2_+ X3_X15_X2_0.29)' X3_X15_X2_/ X3_X15_X2_W' X3_X15_X2_/  W' L='L_N' W='W_N' NF=1 AD='INT((NF+1)/2)
+ AS='INT((NF+2)/2) PD='2*INT((NF+1)/2) PS='2*INT((NF+2)/2) NRD='0.29 NRS='0.29 SA=0 SB=0 SD=0 MULT='N' M='N' 
*--------END___X3_X15_X2_XM1->W'
*--------BEGIN_X3_X15_X2_XM2->W'
XM2_X3_X15_X2 OUT32 GND X3_X15_NET1 VDD X3_X15_X2_SKY130_FD_PR__PFET_01V8 X3_X15_X2_* X3_X15_X2_W/NF X3_X15_X2_* X3_X15_X2_0.29'
+ X3_X15_X2_* X3_X15_X2_W/NF X3_X15_X2_* X3_X15_X2_0.29' X3_X15_X2_* X3_X15_X2_(W/NF X3_X15_X2_+ X3_X15_X2_0.29)'
+ X3_X15_X2_* X3_X15_X2_(W/NF X3_X15_X2_+ X3_X15_X2_0.29)' X3_X15_X2_/ X3_X15_X2_W' X3_X15_X2_/  W' L='L_P' W='W_P' NF=1 AD='INT((NF+1)/2)
+ AS='INT((NF+2)/2) PD='2*INT((NF+1)/2) PS='2*INT((NF+2)/2) NRD='0.29 NRS='0.29 SA=0 SB=0 SD=0 MULT='N' M='N' 
*--------END___X3_X15_X2_XM2->W'
*--------END___X3_X15_X2->TRANSMISSION_GATE
*--------BEGIN_X3_X15_XM1->W'
XM1_X3_X15 X3_X15_NET1 GND X3_VSS X3_VSS X3_X15_SKY130_FD_PR__NFET_01V8 X3_X15_* X3_X15_W/NF X3_X15_* X3_X15_0.29'
+ X3_X15_* X3_X15_W/NF X3_X15_* X3_X15_0.29' X3_X15_* X3_X15_(W/NF X3_X15_+ X3_X15_0.29)' X3_X15_* X3_X15_(W/NF
+ X3_X15_+ X3_X15_0.29)' X3_X15_/ X3_X15_W' X3_X15_/  W' L=0.15 W=0.5 NF=1 AD='INT((NF+1)/2) AS='INT((NF+2)/2) PD='2*INT((NF+1)/2)
+ PS='2*INT((NF+2)/2) NRD='0.29 NRS='0.29 SA=0 SB=0 SD=0 MULT=1 M=1 
*--------END___X3_X15_XM1->W'
*--------END___X3_X15->SWITCH_5T
*--------BEGIN_X3_X16->SKY130_FD_SC_HD__INV_1
X16_X3 GND X3_VGND X3_VNB X3_VPB X3_VPWR X3_NET35  SKY130_FD_SC_HD__INV_1
*--------END___X3_X16->SKY130_FD_SC_HD__INV_1
*--------BEGIN_X3_X17->TRANSMISSION_GATE
*.PININFO IN:B OUT:B EN:I EN_B:I
*--------BEGIN_X3_X17_XM1->W'
XM1_X3_X17 X3_NET16 VDD IN9 X3_VSS X3_X17_SKY130_FD_PR__NFET_01V8 X3_X17_* X3_X17_W/NF X3_X17_* X3_X17_0.29'
+ X3_X17_* X3_X17_W/NF X3_X17_* X3_X17_0.29' X3_X17_* X3_X17_(W/NF X3_X17_+ X3_X17_0.29)' X3_X17_* X3_X17_(W/NF
+ X3_X17_+ X3_X17_0.29)' X3_X17_/ X3_X17_W' X3_X17_/  W' L='L_N' W='W_N' NF=1 AD='INT((NF+1)/2) AS='INT((NF+2)/2) PD='2*INT((NF+1)/2)
+ PS='2*INT((NF+2)/2) NRD='0.29 NRS='0.29 SA=0 SB=0 SD=0 MULT='N' M='N' 
*--------END___X3_X17_XM1->W'
*--------BEGIN_X3_X17_XM2->W'
XM2_X3_X17 X3_NET16 GND IN9 VDD X3_X17_SKY130_FD_PR__PFET_01V8 X3_X17_* X3_X17_W/NF X3_X17_* X3_X17_0.29'
+ X3_X17_* X3_X17_W/NF X3_X17_* X3_X17_0.29' X3_X17_* X3_X17_(W/NF X3_X17_+ X3_X17_0.29)' X3_X17_* X3_X17_(W/NF
+ X3_X17_+ X3_X17_0.29)' X3_X17_/ X3_X17_W' X3_X17_/  W' L='L_P' W='W_P' NF=1 AD='INT((NF+1)/2) AS='INT((NF+2)/2) PD='2*INT((NF+1)/2)
+ PS='2*INT((NF+2)/2) NRD='0.29 NRS='0.29 SA=0 SB=0 SD=0 MULT='N' M='N' 
*--------END___X3_X17_XM2->W'
*--------END___X3_X17->TRANSMISSION_GATE
*--------BEGIN_X3_X18->SWITCH_5T
*.PININFO IN:B OUT:B EN:I EN_B:I
*--------BEGIN_X3_X18_X1->TRANSMISSION_GATE
*.PININFO IN:B OUT:B EN:I EN_B:I
*--------BEGIN_X3_X18_X1_XM1->W'
XM1_X3_X18_X1 X3_X18_NET1 X3_NET36 X3_NET16 X3_VSS X3_X18_X1_SKY130_FD_PR__NFET_01V8 X3_X18_X1_* X3_X18_X1_W/NF X3_X18_X1_* X3_X18_X1_0.29'
+ X3_X18_X1_* X3_X18_X1_W/NF X3_X18_X1_* X3_X18_X1_0.29' X3_X18_X1_* X3_X18_X1_(W/NF X3_X18_X1_+ X3_X18_X1_0.29)'
+ X3_X18_X1_* X3_X18_X1_(W/NF X3_X18_X1_+ X3_X18_X1_0.29)' X3_X18_X1_/ X3_X18_X1_W' X3_X18_X1_/  W' L='L_N' W='W_N' NF=1 AD='INT((NF+1)/2)
+ AS='INT((NF+2)/2) PD='2*INT((NF+1)/2) PS='2*INT((NF+2)/2) NRD='0.29 NRS='0.29 SA=0 SB=0 SD=0 MULT='N' M='N' 
*--------END___X3_X18_X1_XM1->W'
*--------BEGIN_X3_X18_X1_XM2->W'
XM2_X3_X18_X1 X3_X18_NET1 VDD X3_NET16 VDD X3_X18_X1_SKY130_FD_PR__PFET_01V8 X3_X18_X1_* X3_X18_X1_W/NF X3_X18_X1_* X3_X18_X1_0.29'
+ X3_X18_X1_* X3_X18_X1_W/NF X3_X18_X1_* X3_X18_X1_0.29' X3_X18_X1_* X3_X18_X1_(W/NF X3_X18_X1_+ X3_X18_X1_0.29)'
+ X3_X18_X1_* X3_X18_X1_(W/NF X3_X18_X1_+ X3_X18_X1_0.29)' X3_X18_X1_/ X3_X18_X1_W' X3_X18_X1_/  W' L='L_P' W='W_P' NF=1 AD='INT((NF+1)/2)
+ AS='INT((NF+2)/2) PD='2*INT((NF+1)/2) PS='2*INT((NF+2)/2) NRD='0.29 NRS='0.29 SA=0 SB=0 SD=0 MULT='N' M='N' 
*--------END___X3_X18_X1_XM2->W'
*--------END___X3_X18_X1->TRANSMISSION_GATE
*--------BEGIN_X3_X18_X2->TRANSMISSION_GATE
*.PININFO IN:B OUT:B EN:I EN_B:I
*--------BEGIN_X3_X18_X2_XM1->W'
XM1_X3_X18_X2 OUT32 X3_NET36 X3_X18_NET1 X3_VSS X3_X18_X2_SKY130_FD_PR__NFET_01V8 X3_X18_X2_* X3_X18_X2_W/NF X3_X18_X2_* X3_X18_X2_0.29'
+ X3_X18_X2_* X3_X18_X2_W/NF X3_X18_X2_* X3_X18_X2_0.29' X3_X18_X2_* X3_X18_X2_(W/NF X3_X18_X2_+ X3_X18_X2_0.29)'
+ X3_X18_X2_* X3_X18_X2_(W/NF X3_X18_X2_+ X3_X18_X2_0.29)' X3_X18_X2_/ X3_X18_X2_W' X3_X18_X2_/  W' L='L_N' W='W_N' NF=1 AD='INT((NF+1)/2)
+ AS='INT((NF+2)/2) PD='2*INT((NF+1)/2) PS='2*INT((NF+2)/2) NRD='0.29 NRS='0.29 SA=0 SB=0 SD=0 MULT='N' M='N' 
*--------END___X3_X18_X2_XM1->W'
*--------BEGIN_X3_X18_X2_XM2->W'
XM2_X3_X18_X2 OUT32 VDD X3_X18_NET1 VDD X3_X18_X2_SKY130_FD_PR__PFET_01V8 X3_X18_X2_* X3_X18_X2_W/NF X3_X18_X2_* X3_X18_X2_0.29'
+ X3_X18_X2_* X3_X18_X2_W/NF X3_X18_X2_* X3_X18_X2_0.29' X3_X18_X2_* X3_X18_X2_(W/NF X3_X18_X2_+ X3_X18_X2_0.29)'
+ X3_X18_X2_* X3_X18_X2_(W/NF X3_X18_X2_+ X3_X18_X2_0.29)' X3_X18_X2_/ X3_X18_X2_W' X3_X18_X2_/  W' L='L_P' W='W_P' NF=1 AD='INT((NF+1)/2)
+ AS='INT((NF+2)/2) PD='2*INT((NF+1)/2) PS='2*INT((NF+2)/2) NRD='0.29 NRS='0.29 SA=0 SB=0 SD=0 MULT='N' M='N' 
*--------END___X3_X18_X2_XM2->W'
*--------END___X3_X18_X2->TRANSMISSION_GATE
*--------BEGIN_X3_X18_XM1->W'
XM1_X3_X18 X3_X18_NET1 VDD X3_VSS X3_VSS X3_X18_SKY130_FD_PR__NFET_01V8 X3_X18_* X3_X18_W/NF X3_X18_* X3_X18_0.29'
+ X3_X18_* X3_X18_W/NF X3_X18_* X3_X18_0.29' X3_X18_* X3_X18_(W/NF X3_X18_+ X3_X18_0.29)' X3_X18_* X3_X18_(W/NF
+ X3_X18_+ X3_X18_0.29)' X3_X18_/ X3_X18_W' X3_X18_/  W' L=0.15 W=0.5 NF=1 AD='INT((NF+1)/2) AS='INT((NF+2)/2) PD='2*INT((NF+1)/2)
+ PS='2*INT((NF+2)/2) NRD='0.29 NRS='0.29 SA=0 SB=0 SD=0 MULT=1 M=1 
*--------END___X3_X18_XM1->W'
*--------END___X3_X18->SWITCH_5T
*--------BEGIN_X3_X19->SKY130_FD_SC_HD__INV_1
X19_X3 VDD X3_VGND X3_VNB X3_VPB X3_VPWR X3_NET36  SKY130_FD_SC_HD__INV_1
*--------END___X3_X19->SKY130_FD_SC_HD__INV_1
*--------BEGIN_X3_X20->TRANSMISSION_GATE
*.PININFO IN:B OUT:B EN:I EN_B:I
*--------BEGIN_X3_X20_XM1->W'
XM1_X3_X20 X3_NET17 VDD IN1 X3_VSS X3_X20_SKY130_FD_PR__NFET_01V8 X3_X20_* X3_X20_W/NF X3_X20_* X3_X20_0.29'
+ X3_X20_* X3_X20_W/NF X3_X20_* X3_X20_0.29' X3_X20_* X3_X20_(W/NF X3_X20_+ X3_X20_0.29)' X3_X20_* X3_X20_(W/NF
+ X3_X20_+ X3_X20_0.29)' X3_X20_/ X3_X20_W' X3_X20_/  W' L='L_N' W='W_N' NF=1 AD='INT((NF+1)/2) AS='INT((NF+2)/2) PD='2*INT((NF+1)/2)
+ PS='2*INT((NF+2)/2) NRD='0.29 NRS='0.29 SA=0 SB=0 SD=0 MULT='N' M='N' 
*--------END___X3_X20_XM1->W'
*--------BEGIN_X3_X20_XM2->W'
XM2_X3_X20 X3_NET17 GND IN1 VDD X3_X20_SKY130_FD_PR__PFET_01V8 X3_X20_* X3_X20_W/NF X3_X20_* X3_X20_0.29'
+ X3_X20_* X3_X20_W/NF X3_X20_* X3_X20_0.29' X3_X20_* X3_X20_(W/NF X3_X20_+ X3_X20_0.29)' X3_X20_* X3_X20_(W/NF
+ X3_X20_+ X3_X20_0.29)' X3_X20_/ X3_X20_W' X3_X20_/  W' L='L_P' W='W_P' NF=1 AD='INT((NF+1)/2) AS='INT((NF+2)/2) PD='2*INT((NF+1)/2)
+ PS='2*INT((NF+2)/2) NRD='0.29 NRS='0.29 SA=0 SB=0 SD=0 MULT='N' M='N' 
*--------END___X3_X20_XM2->W'
*--------END___X3_X20->TRANSMISSION_GATE
*--------BEGIN_X3_X21->SWITCH_5T
*.PININFO IN:B OUT:B EN:I EN_B:I
*--------BEGIN_X3_X21_X1->TRANSMISSION_GATE
*.PININFO IN:B OUT:B EN:I EN_B:I
*--------BEGIN_X3_X21_X1_XM1->W'
XM1_X3_X21_X1 X3_X21_NET1 X3_NET37 X3_NET17 X3_VSS X3_X21_X1_SKY130_FD_PR__NFET_01V8 X3_X21_X1_* X3_X21_X1_W/NF X3_X21_X1_* X3_X21_X1_0.29'
+ X3_X21_X1_* X3_X21_X1_W/NF X3_X21_X1_* X3_X21_X1_0.29' X3_X21_X1_* X3_X21_X1_(W/NF X3_X21_X1_+ X3_X21_X1_0.29)'
+ X3_X21_X1_* X3_X21_X1_(W/NF X3_X21_X1_+ X3_X21_X1_0.29)' X3_X21_X1_/ X3_X21_X1_W' X3_X21_X1_/  W' L='L_N' W='W_N' NF=1 AD='INT((NF+1)/2)
+ AS='INT((NF+2)/2) PD='2*INT((NF+1)/2) PS='2*INT((NF+2)/2) NRD='0.29 NRS='0.29 SA=0 SB=0 SD=0 MULT='N' M='N' 
*--------END___X3_X21_X1_XM1->W'
*--------BEGIN_X3_X21_X1_XM2->W'
XM2_X3_X21_X1 X3_X21_NET1 VDD X3_NET17 VDD X3_X21_X1_SKY130_FD_PR__PFET_01V8 X3_X21_X1_* X3_X21_X1_W/NF X3_X21_X1_* X3_X21_X1_0.29'
+ X3_X21_X1_* X3_X21_X1_W/NF X3_X21_X1_* X3_X21_X1_0.29' X3_X21_X1_* X3_X21_X1_(W/NF X3_X21_X1_+ X3_X21_X1_0.29)'
+ X3_X21_X1_* X3_X21_X1_(W/NF X3_X21_X1_+ X3_X21_X1_0.29)' X3_X21_X1_/ X3_X21_X1_W' X3_X21_X1_/  W' L='L_P' W='W_P' NF=1 AD='INT((NF+1)/2)
+ AS='INT((NF+2)/2) PD='2*INT((NF+1)/2) PS='2*INT((NF+2)/2) NRD='0.29 NRS='0.29 SA=0 SB=0 SD=0 MULT='N' M='N' 
*--------END___X3_X21_X1_XM2->W'
*--------END___X3_X21_X1->TRANSMISSION_GATE
*--------BEGIN_X3_X21_X2->TRANSMISSION_GATE
*.PININFO IN:B OUT:B EN:I EN_B:I
*--------BEGIN_X3_X21_X2_XM1->W'
XM1_X3_X21_X2 OUT32 X3_NET37 X3_X21_NET1 X3_VSS X3_X21_X2_SKY130_FD_PR__NFET_01V8 X3_X21_X2_* X3_X21_X2_W/NF X3_X21_X2_* X3_X21_X2_0.29'
+ X3_X21_X2_* X3_X21_X2_W/NF X3_X21_X2_* X3_X21_X2_0.29' X3_X21_X2_* X3_X21_X2_(W/NF X3_X21_X2_+ X3_X21_X2_0.29)'
+ X3_X21_X2_* X3_X21_X2_(W/NF X3_X21_X2_+ X3_X21_X2_0.29)' X3_X21_X2_/ X3_X21_X2_W' X3_X21_X2_/  W' L='L_N' W='W_N' NF=1 AD='INT((NF+1)/2)
+ AS='INT((NF+2)/2) PD='2*INT((NF+1)/2) PS='2*INT((NF+2)/2) NRD='0.29 NRS='0.29 SA=0 SB=0 SD=0 MULT='N' M='N' 
*--------END___X3_X21_X2_XM1->W'
*--------BEGIN_X3_X21_X2_XM2->W'
XM2_X3_X21_X2 OUT32 VDD X3_X21_NET1 VDD X3_X21_X2_SKY130_FD_PR__PFET_01V8 X3_X21_X2_* X3_X21_X2_W/NF X3_X21_X2_* X3_X21_X2_0.29'
+ X3_X21_X2_* X3_X21_X2_W/NF X3_X21_X2_* X3_X21_X2_0.29' X3_X21_X2_* X3_X21_X2_(W/NF X3_X21_X2_+ X3_X21_X2_0.29)'
+ X3_X21_X2_* X3_X21_X2_(W/NF X3_X21_X2_+ X3_X21_X2_0.29)' X3_X21_X2_/ X3_X21_X2_W' X3_X21_X2_/  W' L='L_P' W='W_P' NF=1 AD='INT((NF+1)/2)
+ AS='INT((NF+2)/2) PD='2*INT((NF+1)/2) PS='2*INT((NF+2)/2) NRD='0.29 NRS='0.29 SA=0 SB=0 SD=0 MULT='N' M='N' 
*--------END___X3_X21_X2_XM2->W'
*--------END___X3_X21_X2->TRANSMISSION_GATE
*--------BEGIN_X3_X21_XM1->W'
XM1_X3_X21 X3_X21_NET1 VDD X3_VSS X3_VSS X3_X21_SKY130_FD_PR__NFET_01V8 X3_X21_* X3_X21_W/NF X3_X21_* X3_X21_0.29'
+ X3_X21_* X3_X21_W/NF X3_X21_* X3_X21_0.29' X3_X21_* X3_X21_(W/NF X3_X21_+ X3_X21_0.29)' X3_X21_* X3_X21_(W/NF
+ X3_X21_+ X3_X21_0.29)' X3_X21_/ X3_X21_W' X3_X21_/  W' L=0.15 W=0.5 NF=1 AD='INT((NF+1)/2) AS='INT((NF+2)/2) PD='2*INT((NF+1)/2)
+ PS='2*INT((NF+2)/2) NRD='0.29 NRS='0.29 SA=0 SB=0 SD=0 MULT=1 M=1 
*--------END___X3_X21_XM1->W'
*--------END___X3_X21->SWITCH_5T
*--------BEGIN_X3_X22->SKY130_FD_SC_HD__INV_1
X22_X3 VDD X3_VGND X3_VNB X3_VPB X3_VPWR X3_NET37  SKY130_FD_SC_HD__INV_1
*--------END___X3_X22->SKY130_FD_SC_HD__INV_1
*--------BEGIN_X3_X23->TRANSMISSION_GATE
*.PININFO IN:B OUT:B EN:I EN_B:I
*--------BEGIN_X3_X23_XM1->W'
XM1_X3_X23 X3_NET18 VDD IN2 X3_VSS X3_X23_SKY130_FD_PR__NFET_01V8 X3_X23_* X3_X23_W/NF X3_X23_* X3_X23_0.29'
+ X3_X23_* X3_X23_W/NF X3_X23_* X3_X23_0.29' X3_X23_* X3_X23_(W/NF X3_X23_+ X3_X23_0.29)' X3_X23_* X3_X23_(W/NF
+ X3_X23_+ X3_X23_0.29)' X3_X23_/ X3_X23_W' X3_X23_/  W' L='L_N' W='W_N' NF=1 AD='INT((NF+1)/2) AS='INT((NF+2)/2) PD='2*INT((NF+1)/2)
+ PS='2*INT((NF+2)/2) NRD='0.29 NRS='0.29 SA=0 SB=0 SD=0 MULT='N' M='N' 
*--------END___X3_X23_XM1->W'
*--------BEGIN_X3_X23_XM2->W'
XM2_X3_X23 X3_NET18 GND IN2 VDD X3_X23_SKY130_FD_PR__PFET_01V8 X3_X23_* X3_X23_W/NF X3_X23_* X3_X23_0.29'
+ X3_X23_* X3_X23_W/NF X3_X23_* X3_X23_0.29' X3_X23_* X3_X23_(W/NF X3_X23_+ X3_X23_0.29)' X3_X23_* X3_X23_(W/NF
+ X3_X23_+ X3_X23_0.29)' X3_X23_/ X3_X23_W' X3_X23_/  W' L='L_P' W='W_P' NF=1 AD='INT((NF+1)/2) AS='INT((NF+2)/2) PD='2*INT((NF+1)/2)
+ PS='2*INT((NF+2)/2) NRD='0.29 NRS='0.29 SA=0 SB=0 SD=0 MULT='N' M='N' 
*--------END___X3_X23_XM2->W'
*--------END___X3_X23->TRANSMISSION_GATE
*--------BEGIN_X3_X24->SWITCH_5T
*.PININFO IN:B OUT:B EN:I EN_B:I
*--------BEGIN_X3_X24_X1->TRANSMISSION_GATE
*.PININFO IN:B OUT:B EN:I EN_B:I
*--------BEGIN_X3_X24_X1_XM1->W'
XM1_X3_X24_X1 X3_X24_NET1 X3_NET38 X3_NET18 X3_VSS X3_X24_X1_SKY130_FD_PR__NFET_01V8 X3_X24_X1_* X3_X24_X1_W/NF X3_X24_X1_* X3_X24_X1_0.29'
+ X3_X24_X1_* X3_X24_X1_W/NF X3_X24_X1_* X3_X24_X1_0.29' X3_X24_X1_* X3_X24_X1_(W/NF X3_X24_X1_+ X3_X24_X1_0.29)'
+ X3_X24_X1_* X3_X24_X1_(W/NF X3_X24_X1_+ X3_X24_X1_0.29)' X3_X24_X1_/ X3_X24_X1_W' X3_X24_X1_/  W' L='L_N' W='W_N' NF=1 AD='INT((NF+1)/2)
+ AS='INT((NF+2)/2) PD='2*INT((NF+1)/2) PS='2*INT((NF+2)/2) NRD='0.29 NRS='0.29 SA=0 SB=0 SD=0 MULT='N' M='N' 
*--------END___X3_X24_X1_XM1->W'
*--------BEGIN_X3_X24_X1_XM2->W'
XM2_X3_X24_X1 X3_X24_NET1 VDD X3_NET18 VDD X3_X24_X1_SKY130_FD_PR__PFET_01V8 X3_X24_X1_* X3_X24_X1_W/NF X3_X24_X1_* X3_X24_X1_0.29'
+ X3_X24_X1_* X3_X24_X1_W/NF X3_X24_X1_* X3_X24_X1_0.29' X3_X24_X1_* X3_X24_X1_(W/NF X3_X24_X1_+ X3_X24_X1_0.29)'
+ X3_X24_X1_* X3_X24_X1_(W/NF X3_X24_X1_+ X3_X24_X1_0.29)' X3_X24_X1_/ X3_X24_X1_W' X3_X24_X1_/  W' L='L_P' W='W_P' NF=1 AD='INT((NF+1)/2)
+ AS='INT((NF+2)/2) PD='2*INT((NF+1)/2) PS='2*INT((NF+2)/2) NRD='0.29 NRS='0.29 SA=0 SB=0 SD=0 MULT='N' M='N' 
*--------END___X3_X24_X1_XM2->W'
*--------END___X3_X24_X1->TRANSMISSION_GATE
*--------BEGIN_X3_X24_X2->TRANSMISSION_GATE
*.PININFO IN:B OUT:B EN:I EN_B:I
*--------BEGIN_X3_X24_X2_XM1->W'
XM1_X3_X24_X2 OUT32 X3_NET38 X3_X24_NET1 X3_VSS X3_X24_X2_SKY130_FD_PR__NFET_01V8 X3_X24_X2_* X3_X24_X2_W/NF X3_X24_X2_* X3_X24_X2_0.29'
+ X3_X24_X2_* X3_X24_X2_W/NF X3_X24_X2_* X3_X24_X2_0.29' X3_X24_X2_* X3_X24_X2_(W/NF X3_X24_X2_+ X3_X24_X2_0.29)'
+ X3_X24_X2_* X3_X24_X2_(W/NF X3_X24_X2_+ X3_X24_X2_0.29)' X3_X24_X2_/ X3_X24_X2_W' X3_X24_X2_/  W' L='L_N' W='W_N' NF=1 AD='INT((NF+1)/2)
+ AS='INT((NF+2)/2) PD='2*INT((NF+1)/2) PS='2*INT((NF+2)/2) NRD='0.29 NRS='0.29 SA=0 SB=0 SD=0 MULT='N' M='N' 
*--------END___X3_X24_X2_XM1->W'
*--------BEGIN_X3_X24_X2_XM2->W'
XM2_X3_X24_X2 OUT32 VDD X3_X24_NET1 VDD X3_X24_X2_SKY130_FD_PR__PFET_01V8 X3_X24_X2_* X3_X24_X2_W/NF X3_X24_X2_* X3_X24_X2_0.29'
+ X3_X24_X2_* X3_X24_X2_W/NF X3_X24_X2_* X3_X24_X2_0.29' X3_X24_X2_* X3_X24_X2_(W/NF X3_X24_X2_+ X3_X24_X2_0.29)'
+ X3_X24_X2_* X3_X24_X2_(W/NF X3_X24_X2_+ X3_X24_X2_0.29)' X3_X24_X2_/ X3_X24_X2_W' X3_X24_X2_/  W' L='L_P' W='W_P' NF=1 AD='INT((NF+1)/2)
+ AS='INT((NF+2)/2) PD='2*INT((NF+1)/2) PS='2*INT((NF+2)/2) NRD='0.29 NRS='0.29 SA=0 SB=0 SD=0 MULT='N' M='N' 
*--------END___X3_X24_X2_XM2->W'
*--------END___X3_X24_X2->TRANSMISSION_GATE
*--------BEGIN_X3_X24_XM1->W'
XM1_X3_X24 X3_X24_NET1 VDD X3_VSS X3_VSS X3_X24_SKY130_FD_PR__NFET_01V8 X3_X24_* X3_X24_W/NF X3_X24_* X3_X24_0.29'
+ X3_X24_* X3_X24_W/NF X3_X24_* X3_X24_0.29' X3_X24_* X3_X24_(W/NF X3_X24_+ X3_X24_0.29)' X3_X24_* X3_X24_(W/NF
+ X3_X24_+ X3_X24_0.29)' X3_X24_/ X3_X24_W' X3_X24_/  W' L=0.15 W=0.5 NF=1 AD='INT((NF+1)/2) AS='INT((NF+2)/2) PD='2*INT((NF+1)/2)
+ PS='2*INT((NF+2)/2) NRD='0.29 NRS='0.29 SA=0 SB=0 SD=0 MULT=1 M=1 
*--------END___X3_X24_XM1->W'
*--------END___X3_X24->SWITCH_5T
*--------BEGIN_X3_X25->SKY130_FD_SC_HD__INV_1
X25_X3 VDD X3_VGND X3_VNB X3_VPB X3_VPWR X3_NET38  SKY130_FD_SC_HD__INV_1
*--------END___X3_X25->SKY130_FD_SC_HD__INV_1
*--------BEGIN_X3_X26->TRANSMISSION_GATE
*.PININFO IN:B OUT:B EN:I EN_B:I
*--------BEGIN_X3_X26_XM1->W'
XM1_X3_X26 X3_NET19 VDD IN3 X3_VSS X3_X26_SKY130_FD_PR__NFET_01V8 X3_X26_* X3_X26_W/NF X3_X26_* X3_X26_0.29'
+ X3_X26_* X3_X26_W/NF X3_X26_* X3_X26_0.29' X3_X26_* X3_X26_(W/NF X3_X26_+ X3_X26_0.29)' X3_X26_* X3_X26_(W/NF
+ X3_X26_+ X3_X26_0.29)' X3_X26_/ X3_X26_W' X3_X26_/  W' L='L_N' W='W_N' NF=1 AD='INT((NF+1)/2) AS='INT((NF+2)/2) PD='2*INT((NF+1)/2)
+ PS='2*INT((NF+2)/2) NRD='0.29 NRS='0.29 SA=0 SB=0 SD=0 MULT='N' M='N' 
*--------END___X3_X26_XM1->W'
*--------BEGIN_X3_X26_XM2->W'
XM2_X3_X26 X3_NET19 GND IN3 VDD X3_X26_SKY130_FD_PR__PFET_01V8 X3_X26_* X3_X26_W/NF X3_X26_* X3_X26_0.29'
+ X3_X26_* X3_X26_W/NF X3_X26_* X3_X26_0.29' X3_X26_* X3_X26_(W/NF X3_X26_+ X3_X26_0.29)' X3_X26_* X3_X26_(W/NF
+ X3_X26_+ X3_X26_0.29)' X3_X26_/ X3_X26_W' X3_X26_/  W' L='L_P' W='W_P' NF=1 AD='INT((NF+1)/2) AS='INT((NF+2)/2) PD='2*INT((NF+1)/2)
+ PS='2*INT((NF+2)/2) NRD='0.29 NRS='0.29 SA=0 SB=0 SD=0 MULT='N' M='N' 
*--------END___X3_X26_XM2->W'
*--------END___X3_X26->TRANSMISSION_GATE
*--------BEGIN_X3_X27->SWITCH_5T
*.PININFO IN:B OUT:B EN:I EN_B:I
*--------BEGIN_X3_X27_X1->TRANSMISSION_GATE
*.PININFO IN:B OUT:B EN:I EN_B:I
*--------BEGIN_X3_X27_X1_XM1->W'
XM1_X3_X27_X1 X3_X27_NET1 X3_NET39 X3_NET19 X3_VSS X3_X27_X1_SKY130_FD_PR__NFET_01V8 X3_X27_X1_* X3_X27_X1_W/NF X3_X27_X1_* X3_X27_X1_0.29'
+ X3_X27_X1_* X3_X27_X1_W/NF X3_X27_X1_* X3_X27_X1_0.29' X3_X27_X1_* X3_X27_X1_(W/NF X3_X27_X1_+ X3_X27_X1_0.29)'
+ X3_X27_X1_* X3_X27_X1_(W/NF X3_X27_X1_+ X3_X27_X1_0.29)' X3_X27_X1_/ X3_X27_X1_W' X3_X27_X1_/  W' L='L_N' W='W_N' NF=1 AD='INT((NF+1)/2)
+ AS='INT((NF+2)/2) PD='2*INT((NF+1)/2) PS='2*INT((NF+2)/2) NRD='0.29 NRS='0.29 SA=0 SB=0 SD=0 MULT='N' M='N' 
*--------END___X3_X27_X1_XM1->W'
*--------BEGIN_X3_X27_X1_XM2->W'
XM2_X3_X27_X1 X3_X27_NET1 VDD X3_NET19 VDD X3_X27_X1_SKY130_FD_PR__PFET_01V8 X3_X27_X1_* X3_X27_X1_W/NF X3_X27_X1_* X3_X27_X1_0.29'
+ X3_X27_X1_* X3_X27_X1_W/NF X3_X27_X1_* X3_X27_X1_0.29' X3_X27_X1_* X3_X27_X1_(W/NF X3_X27_X1_+ X3_X27_X1_0.29)'
+ X3_X27_X1_* X3_X27_X1_(W/NF X3_X27_X1_+ X3_X27_X1_0.29)' X3_X27_X1_/ X3_X27_X1_W' X3_X27_X1_/  W' L='L_P' W='W_P' NF=1 AD='INT((NF+1)/2)
+ AS='INT((NF+2)/2) PD='2*INT((NF+1)/2) PS='2*INT((NF+2)/2) NRD='0.29 NRS='0.29 SA=0 SB=0 SD=0 MULT='N' M='N' 
*--------END___X3_X27_X1_XM2->W'
*--------END___X3_X27_X1->TRANSMISSION_GATE
*--------BEGIN_X3_X27_X2->TRANSMISSION_GATE
*.PININFO IN:B OUT:B EN:I EN_B:I
*--------BEGIN_X3_X27_X2_XM1->W'
XM1_X3_X27_X2 OUT32 X3_NET39 X3_X27_NET1 X3_VSS X3_X27_X2_SKY130_FD_PR__NFET_01V8 X3_X27_X2_* X3_X27_X2_W/NF X3_X27_X2_* X3_X27_X2_0.29'
+ X3_X27_X2_* X3_X27_X2_W/NF X3_X27_X2_* X3_X27_X2_0.29' X3_X27_X2_* X3_X27_X2_(W/NF X3_X27_X2_+ X3_X27_X2_0.29)'
+ X3_X27_X2_* X3_X27_X2_(W/NF X3_X27_X2_+ X3_X27_X2_0.29)' X3_X27_X2_/ X3_X27_X2_W' X3_X27_X2_/  W' L='L_N' W='W_N' NF=1 AD='INT((NF+1)/2)
+ AS='INT((NF+2)/2) PD='2*INT((NF+1)/2) PS='2*INT((NF+2)/2) NRD='0.29 NRS='0.29 SA=0 SB=0 SD=0 MULT='N' M='N' 
*--------END___X3_X27_X2_XM1->W'
*--------BEGIN_X3_X27_X2_XM2->W'
XM2_X3_X27_X2 OUT32 VDD X3_X27_NET1 VDD X3_X27_X2_SKY130_FD_PR__PFET_01V8 X3_X27_X2_* X3_X27_X2_W/NF X3_X27_X2_* X3_X27_X2_0.29'
+ X3_X27_X2_* X3_X27_X2_W/NF X3_X27_X2_* X3_X27_X2_0.29' X3_X27_X2_* X3_X27_X2_(W/NF X3_X27_X2_+ X3_X27_X2_0.29)'
+ X3_X27_X2_* X3_X27_X2_(W/NF X3_X27_X2_+ X3_X27_X2_0.29)' X3_X27_X2_/ X3_X27_X2_W' X3_X27_X2_/  W' L='L_P' W='W_P' NF=1 AD='INT((NF+1)/2)
+ AS='INT((NF+2)/2) PD='2*INT((NF+1)/2) PS='2*INT((NF+2)/2) NRD='0.29 NRS='0.29 SA=0 SB=0 SD=0 MULT='N' M='N' 
*--------END___X3_X27_X2_XM2->W'
*--------END___X3_X27_X2->TRANSMISSION_GATE
*--------BEGIN_X3_X27_XM1->W'
XM1_X3_X27 X3_X27_NET1 VDD X3_VSS X3_VSS X3_X27_SKY130_FD_PR__NFET_01V8 X3_X27_* X3_X27_W/NF X3_X27_* X3_X27_0.29'
+ X3_X27_* X3_X27_W/NF X3_X27_* X3_X27_0.29' X3_X27_* X3_X27_(W/NF X3_X27_+ X3_X27_0.29)' X3_X27_* X3_X27_(W/NF
+ X3_X27_+ X3_X27_0.29)' X3_X27_/ X3_X27_W' X3_X27_/  W' L=0.15 W=0.5 NF=1 AD='INT((NF+1)/2) AS='INT((NF+2)/2) PD='2*INT((NF+1)/2)
+ PS='2*INT((NF+2)/2) NRD='0.29 NRS='0.29 SA=0 SB=0 SD=0 MULT=1 M=1 
*--------END___X3_X27_XM1->W'
*--------END___X3_X27->SWITCH_5T
*--------BEGIN_X3_X58->SKY130_FD_SC_HD__INV_1
X58_X3 VDD X3_VGND X3_VNB X3_VPB X3_VPWR X3_NET39  SKY130_FD_SC_HD__INV_1
*--------END___X3_X58->SKY130_FD_SC_HD__INV_1
*--------BEGIN_X3_X59->TRANSMISSION_GATE
*.PININFO IN:B OUT:B EN:I EN_B:I
*--------BEGIN_X3_X59_XM1->W'
XM1_X3_X59 X3_NET20 VDD IN0 X3_VSS X3_X59_SKY130_FD_PR__NFET_01V8 X3_X59_* X3_X59_W/NF X3_X59_* X3_X59_0.29'
+ X3_X59_* X3_X59_W/NF X3_X59_* X3_X59_0.29' X3_X59_* X3_X59_(W/NF X3_X59_+ X3_X59_0.29)' X3_X59_* X3_X59_(W/NF
+ X3_X59_+ X3_X59_0.29)' X3_X59_/ X3_X59_W' X3_X59_/  W' L='L_N' W='W_N' NF=1 AD='INT((NF+1)/2) AS='INT((NF+2)/2) PD='2*INT((NF+1)/2)
+ PS='2*INT((NF+2)/2) NRD='0.29 NRS='0.29 SA=0 SB=0 SD=0 MULT='N' M='N' 
*--------END___X3_X59_XM1->W'
*--------BEGIN_X3_X59_XM2->W'
XM2_X3_X59 X3_NET20 GND IN0 VDD X3_X59_SKY130_FD_PR__PFET_01V8 X3_X59_* X3_X59_W/NF X3_X59_* X3_X59_0.29'
+ X3_X59_* X3_X59_W/NF X3_X59_* X3_X59_0.29' X3_X59_* X3_X59_(W/NF X3_X59_+ X3_X59_0.29)' X3_X59_* X3_X59_(W/NF
+ X3_X59_+ X3_X59_0.29)' X3_X59_/ X3_X59_W' X3_X59_/  W' L='L_P' W='W_P' NF=1 AD='INT((NF+1)/2) AS='INT((NF+2)/2) PD='2*INT((NF+1)/2)
+ PS='2*INT((NF+2)/2) NRD='0.29 NRS='0.29 SA=0 SB=0 SD=0 MULT='N' M='N' 
*--------END___X3_X59_XM2->W'
*--------END___X3_X59->TRANSMISSION_GATE
*--------BEGIN_X3_X60->SWITCH_5T
*.PININFO IN:B OUT:B EN:I EN_B:I
*--------BEGIN_X3_X60_X1->TRANSMISSION_GATE
*.PININFO IN:B OUT:B EN:I EN_B:I
*--------BEGIN_X3_X60_X1_XM1->W'
XM1_X3_X60_X1 X3_X60_NET1 X3_NET40 X3_NET20 X3_VSS X3_X60_X1_SKY130_FD_PR__NFET_01V8 X3_X60_X1_* X3_X60_X1_W/NF X3_X60_X1_* X3_X60_X1_0.29'
+ X3_X60_X1_* X3_X60_X1_W/NF X3_X60_X1_* X3_X60_X1_0.29' X3_X60_X1_* X3_X60_X1_(W/NF X3_X60_X1_+ X3_X60_X1_0.29)'
+ X3_X60_X1_* X3_X60_X1_(W/NF X3_X60_X1_+ X3_X60_X1_0.29)' X3_X60_X1_/ X3_X60_X1_W' X3_X60_X1_/  W' L='L_N' W='W_N' NF=1 AD='INT((NF+1)/2)
+ AS='INT((NF+2)/2) PD='2*INT((NF+1)/2) PS='2*INT((NF+2)/2) NRD='0.29 NRS='0.29 SA=0 SB=0 SD=0 MULT='N' M='N' 
*--------END___X3_X60_X1_XM1->W'
*--------BEGIN_X3_X60_X1_XM2->W'
XM2_X3_X60_X1 X3_X60_NET1 VDD X3_NET20 VDD X3_X60_X1_SKY130_FD_PR__PFET_01V8 X3_X60_X1_* X3_X60_X1_W/NF X3_X60_X1_* X3_X60_X1_0.29'
+ X3_X60_X1_* X3_X60_X1_W/NF X3_X60_X1_* X3_X60_X1_0.29' X3_X60_X1_* X3_X60_X1_(W/NF X3_X60_X1_+ X3_X60_X1_0.29)'
+ X3_X60_X1_* X3_X60_X1_(W/NF X3_X60_X1_+ X3_X60_X1_0.29)' X3_X60_X1_/ X3_X60_X1_W' X3_X60_X1_/  W' L='L_P' W='W_P' NF=1 AD='INT((NF+1)/2)
+ AS='INT((NF+2)/2) PD='2*INT((NF+1)/2) PS='2*INT((NF+2)/2) NRD='0.29 NRS='0.29 SA=0 SB=0 SD=0 MULT='N' M='N' 
*--------END___X3_X60_X1_XM2->W'
*--------END___X3_X60_X1->TRANSMISSION_GATE
*--------BEGIN_X3_X60_X2->TRANSMISSION_GATE
*.PININFO IN:B OUT:B EN:I EN_B:I
*--------BEGIN_X3_X60_X2_XM1->W'
XM1_X3_X60_X2 OUT32 X3_NET40 X3_X60_NET1 X3_VSS X3_X60_X2_SKY130_FD_PR__NFET_01V8 X3_X60_X2_* X3_X60_X2_W/NF X3_X60_X2_* X3_X60_X2_0.29'
+ X3_X60_X2_* X3_X60_X2_W/NF X3_X60_X2_* X3_X60_X2_0.29' X3_X60_X2_* X3_X60_X2_(W/NF X3_X60_X2_+ X3_X60_X2_0.29)'
+ X3_X60_X2_* X3_X60_X2_(W/NF X3_X60_X2_+ X3_X60_X2_0.29)' X3_X60_X2_/ X3_X60_X2_W' X3_X60_X2_/  W' L='L_N' W='W_N' NF=1 AD='INT((NF+1)/2)
+ AS='INT((NF+2)/2) PD='2*INT((NF+1)/2) PS='2*INT((NF+2)/2) NRD='0.29 NRS='0.29 SA=0 SB=0 SD=0 MULT='N' M='N' 
*--------END___X3_X60_X2_XM1->W'
*--------BEGIN_X3_X60_X2_XM2->W'
XM2_X3_X60_X2 OUT32 VDD X3_X60_NET1 VDD X3_X60_X2_SKY130_FD_PR__PFET_01V8 X3_X60_X2_* X3_X60_X2_W/NF X3_X60_X2_* X3_X60_X2_0.29'
+ X3_X60_X2_* X3_X60_X2_W/NF X3_X60_X2_* X3_X60_X2_0.29' X3_X60_X2_* X3_X60_X2_(W/NF X3_X60_X2_+ X3_X60_X2_0.29)'
+ X3_X60_X2_* X3_X60_X2_(W/NF X3_X60_X2_+ X3_X60_X2_0.29)' X3_X60_X2_/ X3_X60_X2_W' X3_X60_X2_/  W' L='L_P' W='W_P' NF=1 AD='INT((NF+1)/2)
+ AS='INT((NF+2)/2) PD='2*INT((NF+1)/2) PS='2*INT((NF+2)/2) NRD='0.29 NRS='0.29 SA=0 SB=0 SD=0 MULT='N' M='N' 
*--------END___X3_X60_X2_XM2->W'
*--------END___X3_X60_X2->TRANSMISSION_GATE
*--------BEGIN_X3_X60_XM1->W'
XM1_X3_X60 X3_X60_NET1 VDD X3_VSS X3_VSS X3_X60_SKY130_FD_PR__NFET_01V8 X3_X60_* X3_X60_W/NF X3_X60_* X3_X60_0.29'
+ X3_X60_* X3_X60_W/NF X3_X60_* X3_X60_0.29' X3_X60_* X3_X60_(W/NF X3_X60_+ X3_X60_0.29)' X3_X60_* X3_X60_(W/NF
+ X3_X60_+ X3_X60_0.29)' X3_X60_/ X3_X60_W' X3_X60_/  W' L=0.15 W=0.5 NF=1 AD='INT((NF+1)/2) AS='INT((NF+2)/2) PD='2*INT((NF+1)/2)
+ PS='2*INT((NF+2)/2) NRD='0.29 NRS='0.29 SA=0 SB=0 SD=0 MULT=1 M=1 
*--------END___X3_X60_XM1->W'
*--------END___X3_X60->SWITCH_5T
*--------BEGIN_X3_X61->SKY130_FD_SC_HD__INV_1
X61_X3 VDD X3_VGND X3_VNB X3_VPB X3_VPWR X3_NET40  SKY130_FD_SC_HD__INV_1
*--------END___X3_X61->SKY130_FD_SC_HD__INV_1
*--------END___X3->LINE_SWITCHES
V8 IN4 GND 0.5
V9 IN5 GND 0.6
V10 IN6 GND 0.7
V11 IN7 GND 0.8
V12 IN8 GND 0.9
V13 IN9 GND 1.0
V14 IN10 GND 1.1
V15 IN11 GND 1.2
V16 IN12 GND 1.3
V17 IN13 GND 1.4
V18 IN14 GND 1.5
V19 IN15 GND 1.6
V20 IN16 GND 1.7
V21 IN17 GND 1.8
V22 IN18 GND 1.9
V23 IN19 GND 2.0
**** BEGIN USER ARCHITECTURE CODE


.OPTIONS SAVECURRENTS
.CONTROL
TRAN 0.1N 30N
WRITE A_MUX_TB.RAW
.ENDC



** OPENCIRCUITDESIGN PDKS INSTALL
.LIB /FARMSHARE/HOME/CLASSES/EE/372/PDKS/OPEN_PDKS_1.0.310/SKY130/SKY130A/LIBS.TECH/NGSPICE/SKY130.LIB.SPICE TT
.INC /FARMSHARE/HOME/CLASSES/EE/372/PDKS/OPEN_PDKS_1.0.310/SKY130/SKY130A/LIBS.REF/SKY130_FD_SC_HD/SPICE/SKY130_FD_SC_HD.SPICE

**** END USER ARCHITECTURE CODE
.end
