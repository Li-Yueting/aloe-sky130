VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO sky130_asc_pfet_01v8_lvt_9
  CLASS CORE ;
  FOREIGN sky130_asc_pfet_01v8_lvt_9 ;
  ORIGIN 0.000 0.000 ;
  SIZE 2.940 BY 9.400 ;
  SITE unitasc ;
  PIN GATE
    DIRECTION INOUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 116.099998 ;
    PORT
      LAYER li1 ;
        RECT 0.000 0.520 21.260 0.820 ;
    END
  END GATE
  PIN SOURCE
    DIRECTION INOUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 9.352500 ;
    PORT
      LAYER li1 ;
        RECT 0.000 8.650 21.260 8.950 ;
        RECT 2.525 8.245 2.695 8.650 ;
        RECT 7.105 8.245 7.275 8.650 ;
        RECT 11.685 8.245 11.855 8.650 ;
        RECT 16.265 8.245 16.435 8.650 ;
        RECT 20.845 8.245 21.015 8.650 ;
        RECT 2.525 8.130 2.700 8.245 ;
        RECT 7.105 8.130 7.280 8.245 ;
        RECT 11.685 8.130 11.860 8.245 ;
        RECT 16.265 8.130 16.440 8.245 ;
        RECT 20.845 8.130 21.020 8.245 ;
        RECT 2.530 1.755 2.700 8.130 ;
        RECT 7.110 1.755 7.280 8.130 ;
        RECT 11.690 1.755 11.860 8.130 ;
        RECT 16.270 1.755 16.440 8.130 ;
        RECT 20.850 1.755 21.020 8.130 ;
      LAYER mcon ;
        RECT 2.530 1.835 2.700 8.165 ;
        RECT 7.110 1.835 7.280 8.165 ;
        RECT 11.690 1.835 11.860 8.165 ;
        RECT 16.270 1.835 16.440 8.165 ;
        RECT 20.850 1.835 21.020 8.165 ;
      LAYER met1 ;
        RECT 2.500 1.775 2.730 8.225 ;
        RECT 7.080 1.775 7.310 8.225 ;
        RECT 11.660 1.775 11.890 8.225 ;
        RECT 16.240 1.775 16.470 8.225 ;
        RECT 20.820 1.775 21.050 8.225 ;
    END
  END SOURCE
  PIN DRAIN
    DIRECTION INOUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 9.352500 ;
    PORT
      LAYER li1 ;
        RECT 0.240 1.870 0.410 8.245 ;
        RECT 4.820 1.870 4.990 8.245 ;
        RECT 9.400 1.870 9.570 8.245 ;
        RECT 13.980 1.870 14.150 8.245 ;
        RECT 18.560 1.870 18.730 8.245 ;
        RECT 0.235 1.755 0.410 1.870 ;
        RECT 4.815 1.755 4.990 1.870 ;
        RECT 9.395 1.755 9.570 1.870 ;
        RECT 13.975 1.755 14.150 1.870 ;
        RECT 18.555 1.755 18.730 1.870 ;
        RECT 0.235 1.350 0.405 1.755 ;
        RECT 4.815 1.350 4.985 1.755 ;
        RECT 9.395 1.350 9.565 1.755 ;
        RECT 13.975 1.350 14.145 1.755 ;
        RECT 18.555 1.350 18.725 1.755 ;
        RECT 0.000 1.050 21.260 1.350 ;
      LAYER mcon ;
        RECT 0.240 1.835 0.410 8.165 ;
        RECT 4.820 1.835 4.990 8.165 ;
        RECT 9.400 1.835 9.570 8.165 ;
        RECT 13.980 1.835 14.150 8.165 ;
        RECT 18.560 1.835 18.730 8.165 ;
      LAYER met1 ;
        RECT 0.210 1.775 0.440 8.225 ;
        RECT 4.790 1.775 5.020 8.225 ;
        RECT 9.370 1.775 9.600 8.225 ;
        RECT 13.950 1.775 14.180 8.225 ;
        RECT 18.530 1.775 18.760 8.225 ;
    END
  END DRAIN
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT 0.000 1.465 21.260 9.700 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER li1 ;
        RECT 0.000 9.250 21.260 9.550 ;
      LAYER mcon ;
        RECT 0.850 9.250 1.150 9.550 ;
        RECT 2.850 9.250 3.150 9.550 ;
        RECT 4.850 9.250 5.150 9.550 ;
        RECT 6.850 9.250 7.150 9.550 ;
        RECT 8.850 9.250 9.150 9.550 ;
        RECT 10.850 9.250 11.150 9.550 ;
        RECT 12.850 9.250 13.150 9.550 ;
        RECT 14.850 9.250 15.150 9.550 ;
        RECT 16.850 9.250 17.150 9.550 ;
        RECT 18.850 9.250 19.150 9.550 ;
      LAYER met1 ;
        RECT 0.000 9.100 21.260 9.700 ;
    END
  END VPWR
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER li1 ;
        RECT 0.000 -0.150 21.260 0.150 ;
      LAYER mcon ;
        RECT 0.850 -0.150 1.150 0.150 ;
        RECT 2.850 -0.150 3.150 0.150 ;
        RECT 4.850 -0.150 5.150 0.150 ;
        RECT 6.850 -0.150 7.150 0.150 ;
        RECT 8.850 -0.150 9.150 0.150 ;
        RECT 10.850 -0.150 11.150 0.150 ;
        RECT 12.850 -0.150 13.150 0.150 ;
        RECT 14.850 -0.150 15.150 0.150 ;
        RECT 16.850 -0.150 17.150 0.150 ;
        RECT 18.850 -0.150 19.150 0.150 ;
      LAYER met1 ;
        RECT 0.000 -0.300 21.260 0.300 ;
    END
  END VGND
END sky130_asc_pfet_01v8_lvt_9
END LIBRARY

