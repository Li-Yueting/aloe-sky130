magic
tech sky130A
magscale 1 2
timestamp 1652937205
<< nwell >>
rect 90 1707 27796 1940
rect 90 294 27797 1707
rect 187 293 27797 294
<< pmoslvt >>
rect 281 355 681 1645
rect 739 355 1139 1645
rect 1197 355 1597 1645
rect 1655 355 2055 1645
rect 2113 355 2513 1645
rect 2571 355 2971 1645
rect 3029 355 3429 1645
rect 3487 355 3887 1645
rect 3945 355 4345 1645
rect 4403 355 4803 1645
rect 4861 355 5261 1645
rect 5319 355 5719 1645
rect 5777 355 6177 1645
rect 6235 355 6635 1645
rect 6693 355 7093 1645
rect 7151 355 7551 1645
rect 7609 355 8009 1645
rect 8067 355 8467 1645
rect 8525 355 8925 1645
rect 8983 355 9383 1645
rect 9441 355 9841 1645
rect 9899 355 10299 1645
rect 10357 355 10757 1645
rect 10815 355 11215 1645
rect 11273 355 11673 1645
rect 11731 355 12131 1645
rect 12189 355 12589 1645
rect 12647 355 13047 1645
rect 13105 355 13505 1645
rect 13563 355 13963 1645
rect 14021 355 14421 1645
rect 14479 355 14879 1645
rect 14937 355 15337 1645
rect 15395 355 15795 1645
rect 15853 355 16253 1645
rect 16311 355 16711 1645
rect 16769 355 17169 1645
rect 17227 355 17627 1645
rect 17685 355 18085 1645
rect 18143 355 18543 1645
rect 18601 355 19001 1645
rect 19059 355 19459 1645
rect 19517 355 19917 1645
rect 19975 355 20375 1645
rect 20433 355 20833 1645
rect 20891 355 21291 1645
rect 21349 355 21749 1645
rect 21807 355 22207 1645
rect 22265 355 22665 1645
rect 22723 355 23123 1645
rect 23181 355 23581 1645
rect 23639 355 24039 1645
rect 24097 355 24497 1645
rect 24555 355 24955 1645
rect 25013 355 25413 1645
rect 25471 355 25871 1645
rect 25929 355 26329 1645
rect 26387 355 26787 1645
rect 26845 355 27245 1645
rect 27303 355 27703 1645
<< pdiff >>
rect 223 1633 281 1645
rect 223 367 235 1633
rect 269 367 281 1633
rect 223 355 281 367
rect 681 1633 739 1645
rect 681 367 693 1633
rect 727 367 739 1633
rect 681 355 739 367
rect 1139 1633 1197 1645
rect 1139 367 1151 1633
rect 1185 367 1197 1633
rect 1139 355 1197 367
rect 1597 1633 1655 1645
rect 1597 367 1609 1633
rect 1643 367 1655 1633
rect 1597 355 1655 367
rect 2055 1633 2113 1645
rect 2055 367 2067 1633
rect 2101 367 2113 1633
rect 2055 355 2113 367
rect 2513 1633 2571 1645
rect 2513 367 2525 1633
rect 2559 367 2571 1633
rect 2513 355 2571 367
rect 2971 1633 3029 1645
rect 2971 367 2983 1633
rect 3017 367 3029 1633
rect 2971 355 3029 367
rect 3429 1633 3487 1645
rect 3429 367 3441 1633
rect 3475 367 3487 1633
rect 3429 355 3487 367
rect 3887 1633 3945 1645
rect 3887 367 3899 1633
rect 3933 367 3945 1633
rect 3887 355 3945 367
rect 4345 1633 4403 1645
rect 4345 367 4357 1633
rect 4391 367 4403 1633
rect 4345 355 4403 367
rect 4803 1633 4861 1645
rect 4803 367 4815 1633
rect 4849 367 4861 1633
rect 4803 355 4861 367
rect 5261 1633 5319 1645
rect 5261 367 5273 1633
rect 5307 367 5319 1633
rect 5261 355 5319 367
rect 5719 1633 5777 1645
rect 5719 367 5731 1633
rect 5765 367 5777 1633
rect 5719 355 5777 367
rect 6177 1633 6235 1645
rect 6177 367 6189 1633
rect 6223 367 6235 1633
rect 6177 355 6235 367
rect 6635 1633 6693 1645
rect 6635 367 6647 1633
rect 6681 367 6693 1633
rect 6635 355 6693 367
rect 7093 1633 7151 1645
rect 7093 367 7105 1633
rect 7139 367 7151 1633
rect 7093 355 7151 367
rect 7551 1633 7609 1645
rect 7551 367 7563 1633
rect 7597 367 7609 1633
rect 7551 355 7609 367
rect 8009 1633 8067 1645
rect 8009 367 8021 1633
rect 8055 367 8067 1633
rect 8009 355 8067 367
rect 8467 1633 8525 1645
rect 8467 367 8479 1633
rect 8513 367 8525 1633
rect 8467 355 8525 367
rect 8925 1633 8983 1645
rect 8925 367 8937 1633
rect 8971 367 8983 1633
rect 8925 355 8983 367
rect 9383 1633 9441 1645
rect 9383 367 9395 1633
rect 9429 367 9441 1633
rect 9383 355 9441 367
rect 9841 1633 9899 1645
rect 9841 367 9853 1633
rect 9887 367 9899 1633
rect 9841 355 9899 367
rect 10299 1633 10357 1645
rect 10299 367 10311 1633
rect 10345 367 10357 1633
rect 10299 355 10357 367
rect 10757 1633 10815 1645
rect 10757 367 10769 1633
rect 10803 367 10815 1633
rect 10757 355 10815 367
rect 11215 1633 11273 1645
rect 11215 367 11227 1633
rect 11261 367 11273 1633
rect 11215 355 11273 367
rect 11673 1633 11731 1645
rect 11673 367 11685 1633
rect 11719 367 11731 1633
rect 11673 355 11731 367
rect 12131 1633 12189 1645
rect 12131 367 12143 1633
rect 12177 367 12189 1633
rect 12131 355 12189 367
rect 12589 1633 12647 1645
rect 12589 367 12601 1633
rect 12635 367 12647 1633
rect 12589 355 12647 367
rect 13047 1633 13105 1645
rect 13047 367 13059 1633
rect 13093 367 13105 1633
rect 13047 355 13105 367
rect 13505 1633 13563 1645
rect 13505 367 13517 1633
rect 13551 367 13563 1633
rect 13505 355 13563 367
rect 13963 1633 14021 1645
rect 13963 367 13975 1633
rect 14009 367 14021 1633
rect 13963 355 14021 367
rect 14421 1633 14479 1645
rect 14421 367 14433 1633
rect 14467 367 14479 1633
rect 14421 355 14479 367
rect 14879 1633 14937 1645
rect 14879 367 14891 1633
rect 14925 367 14937 1633
rect 14879 355 14937 367
rect 15337 1633 15395 1645
rect 15337 367 15349 1633
rect 15383 367 15395 1633
rect 15337 355 15395 367
rect 15795 1633 15853 1645
rect 15795 367 15807 1633
rect 15841 367 15853 1633
rect 15795 355 15853 367
rect 16253 1633 16311 1645
rect 16253 367 16265 1633
rect 16299 367 16311 1633
rect 16253 355 16311 367
rect 16711 1633 16769 1645
rect 16711 367 16723 1633
rect 16757 367 16769 1633
rect 16711 355 16769 367
rect 17169 1633 17227 1645
rect 17169 367 17181 1633
rect 17215 367 17227 1633
rect 17169 355 17227 367
rect 17627 1633 17685 1645
rect 17627 367 17639 1633
rect 17673 367 17685 1633
rect 17627 355 17685 367
rect 18085 1633 18143 1645
rect 18085 367 18097 1633
rect 18131 367 18143 1633
rect 18085 355 18143 367
rect 18543 1633 18601 1645
rect 18543 367 18555 1633
rect 18589 367 18601 1633
rect 18543 355 18601 367
rect 19001 1633 19059 1645
rect 19001 367 19013 1633
rect 19047 367 19059 1633
rect 19001 355 19059 367
rect 19459 1633 19517 1645
rect 19459 367 19471 1633
rect 19505 367 19517 1633
rect 19459 355 19517 367
rect 19917 1633 19975 1645
rect 19917 367 19929 1633
rect 19963 367 19975 1633
rect 19917 355 19975 367
rect 20375 1633 20433 1645
rect 20375 367 20387 1633
rect 20421 367 20433 1633
rect 20375 355 20433 367
rect 20833 1633 20891 1645
rect 20833 367 20845 1633
rect 20879 367 20891 1633
rect 20833 355 20891 367
rect 21291 1633 21349 1645
rect 21291 367 21303 1633
rect 21337 367 21349 1633
rect 21291 355 21349 367
rect 21749 1633 21807 1645
rect 21749 367 21761 1633
rect 21795 367 21807 1633
rect 21749 355 21807 367
rect 22207 1633 22265 1645
rect 22207 367 22219 1633
rect 22253 367 22265 1633
rect 22207 355 22265 367
rect 22665 1633 22723 1645
rect 22665 367 22677 1633
rect 22711 367 22723 1633
rect 22665 355 22723 367
rect 23123 1633 23181 1645
rect 23123 367 23135 1633
rect 23169 367 23181 1633
rect 23123 355 23181 367
rect 23581 1633 23639 1645
rect 23581 367 23593 1633
rect 23627 367 23639 1633
rect 23581 355 23639 367
rect 24039 1633 24097 1645
rect 24039 367 24051 1633
rect 24085 367 24097 1633
rect 24039 355 24097 367
rect 24497 1633 24555 1645
rect 24497 367 24509 1633
rect 24543 367 24555 1633
rect 24497 355 24555 367
rect 24955 1633 25013 1645
rect 24955 367 24967 1633
rect 25001 367 25013 1633
rect 24955 355 25013 367
rect 25413 1633 25471 1645
rect 25413 367 25425 1633
rect 25459 367 25471 1633
rect 25413 355 25471 367
rect 25871 1633 25929 1645
rect 25871 367 25883 1633
rect 25917 367 25929 1633
rect 25871 355 25929 367
rect 26329 1633 26387 1645
rect 26329 367 26341 1633
rect 26375 367 26387 1633
rect 26329 355 26387 367
rect 26787 1633 26845 1645
rect 26787 367 26799 1633
rect 26833 367 26845 1633
rect 26787 355 26845 367
rect 27245 1633 27303 1645
rect 27245 367 27257 1633
rect 27291 367 27303 1633
rect 27245 355 27303 367
rect 27703 1633 27761 1645
rect 27703 367 27715 1633
rect 27749 367 27761 1633
rect 27703 355 27761 367
<< pdiffc >>
rect 235 367 269 1633
rect 693 367 727 1633
rect 1151 367 1185 1633
rect 1609 367 1643 1633
rect 2067 367 2101 1633
rect 2525 367 2559 1633
rect 2983 367 3017 1633
rect 3441 367 3475 1633
rect 3899 367 3933 1633
rect 4357 367 4391 1633
rect 4815 367 4849 1633
rect 5273 367 5307 1633
rect 5731 367 5765 1633
rect 6189 367 6223 1633
rect 6647 367 6681 1633
rect 7105 367 7139 1633
rect 7563 367 7597 1633
rect 8021 367 8055 1633
rect 8479 367 8513 1633
rect 8937 367 8971 1633
rect 9395 367 9429 1633
rect 9853 367 9887 1633
rect 10311 367 10345 1633
rect 10769 367 10803 1633
rect 11227 367 11261 1633
rect 11685 367 11719 1633
rect 12143 367 12177 1633
rect 12601 367 12635 1633
rect 13059 367 13093 1633
rect 13517 367 13551 1633
rect 13975 367 14009 1633
rect 14433 367 14467 1633
rect 14891 367 14925 1633
rect 15349 367 15383 1633
rect 15807 367 15841 1633
rect 16265 367 16299 1633
rect 16723 367 16757 1633
rect 17181 367 17215 1633
rect 17639 367 17673 1633
rect 18097 367 18131 1633
rect 18555 367 18589 1633
rect 19013 367 19047 1633
rect 19471 367 19505 1633
rect 19929 367 19963 1633
rect 20387 367 20421 1633
rect 20845 367 20879 1633
rect 21303 367 21337 1633
rect 21761 367 21795 1633
rect 22219 367 22253 1633
rect 22677 367 22711 1633
rect 23135 367 23169 1633
rect 23593 367 23627 1633
rect 24051 367 24085 1633
rect 24509 367 24543 1633
rect 24967 367 25001 1633
rect 25425 367 25459 1633
rect 25883 367 25917 1633
rect 26341 367 26375 1633
rect 26799 367 26833 1633
rect 27257 367 27291 1633
rect 27715 367 27749 1633
<< nsubdiff >>
rect 1186 1808 1306 1810
rect 128 1760 168 1800
rect 1186 1772 1226 1808
rect 1270 1772 1306 1808
rect 1186 1770 1306 1772
rect 2486 1808 2606 1810
rect 2486 1772 2526 1808
rect 2570 1772 2606 1808
rect 2486 1770 2606 1772
rect 3786 1808 3906 1810
rect 3786 1772 3826 1808
rect 3870 1772 3906 1808
rect 3786 1770 3906 1772
rect 5086 1808 5206 1810
rect 5086 1772 5126 1808
rect 5170 1772 5206 1808
rect 5086 1770 5206 1772
rect 6386 1808 6506 1810
rect 6386 1772 6426 1808
rect 6470 1772 6506 1808
rect 6386 1770 6506 1772
rect 7686 1808 7806 1810
rect 7686 1772 7726 1808
rect 7770 1772 7806 1808
rect 7686 1770 7806 1772
rect 8986 1808 9106 1810
rect 8986 1772 9026 1808
rect 9070 1772 9106 1808
rect 8986 1770 9106 1772
rect 10286 1808 10406 1810
rect 10286 1772 10326 1808
rect 10370 1772 10406 1808
rect 10286 1770 10406 1772
rect 11586 1808 11706 1810
rect 11586 1772 11626 1808
rect 11670 1772 11706 1808
rect 11586 1770 11706 1772
rect 12886 1808 13006 1810
rect 12886 1772 12926 1808
rect 12970 1772 13006 1808
rect 12886 1770 13006 1772
rect 14186 1808 14306 1810
rect 14186 1772 14226 1808
rect 14270 1772 14306 1808
rect 14186 1770 14306 1772
rect 15486 1808 15606 1810
rect 15486 1772 15526 1808
rect 15570 1772 15606 1808
rect 15486 1770 15606 1772
rect 16786 1808 16906 1810
rect 16786 1772 16826 1808
rect 16870 1772 16906 1808
rect 16786 1770 16906 1772
rect 18086 1808 18206 1810
rect 18086 1772 18126 1808
rect 18170 1772 18206 1808
rect 18086 1770 18206 1772
rect 19386 1808 19506 1810
rect 19386 1772 19426 1808
rect 19470 1772 19506 1808
rect 19386 1770 19506 1772
rect 20686 1808 20806 1810
rect 20686 1772 20726 1808
rect 20770 1772 20806 1808
rect 20686 1770 20806 1772
rect 21986 1808 22106 1810
rect 21986 1772 22026 1808
rect 22070 1772 22106 1808
rect 21986 1770 22106 1772
rect 23286 1808 23406 1810
rect 23286 1772 23326 1808
rect 23370 1772 23406 1808
rect 23286 1770 23406 1772
rect 24586 1808 24706 1810
rect 24586 1772 24626 1808
rect 24670 1772 24706 1808
rect 24586 1770 24706 1772
rect 25886 1808 26006 1810
rect 25886 1772 25926 1808
rect 25970 1772 26006 1808
rect 25886 1770 26006 1772
rect 128 1680 168 1720
<< nsubdiffcont >>
rect 1226 1772 1270 1808
rect 2526 1772 2570 1808
rect 3826 1772 3870 1808
rect 5126 1772 5170 1808
rect 6426 1772 6470 1808
rect 7726 1772 7770 1808
rect 9026 1772 9070 1808
rect 10326 1772 10370 1808
rect 11626 1772 11670 1808
rect 12926 1772 12970 1808
rect 14226 1772 14270 1808
rect 15526 1772 15570 1808
rect 16826 1772 16870 1808
rect 18126 1772 18170 1808
rect 19426 1772 19470 1808
rect 20726 1772 20770 1808
rect 22026 1772 22070 1808
rect 23326 1772 23370 1808
rect 24626 1772 24670 1808
rect 25926 1772 25970 1808
rect 128 1720 168 1760
<< poly >>
rect 281 1645 681 1671
rect 739 1645 1139 1671
rect 1197 1645 1597 1671
rect 1655 1645 2055 1671
rect 2113 1645 2513 1671
rect 2571 1645 2971 1671
rect 3029 1645 3429 1671
rect 3487 1645 3887 1671
rect 3945 1645 4345 1671
rect 4403 1645 4803 1671
rect 4861 1645 5261 1671
rect 5319 1645 5719 1671
rect 5777 1645 6177 1671
rect 6235 1645 6635 1671
rect 6693 1645 7093 1671
rect 7151 1645 7551 1671
rect 7609 1645 8009 1671
rect 8067 1645 8467 1671
rect 8525 1645 8925 1671
rect 8983 1645 9383 1671
rect 9441 1645 9841 1671
rect 9899 1645 10299 1671
rect 10357 1645 10757 1671
rect 10815 1645 11215 1671
rect 11273 1645 11673 1671
rect 11731 1645 12131 1671
rect 12189 1645 12589 1671
rect 12647 1645 13047 1671
rect 13105 1645 13505 1671
rect 13563 1645 13963 1671
rect 14021 1645 14421 1671
rect 14479 1645 14879 1671
rect 14937 1645 15337 1671
rect 15395 1645 15795 1671
rect 15853 1645 16253 1671
rect 16311 1645 16711 1671
rect 16769 1645 17169 1671
rect 17227 1645 17627 1671
rect 17685 1645 18085 1671
rect 18143 1645 18543 1671
rect 18601 1645 19001 1671
rect 19059 1645 19459 1671
rect 19517 1645 19917 1671
rect 19975 1645 20375 1671
rect 20433 1645 20833 1671
rect 20891 1645 21291 1671
rect 21349 1645 21749 1671
rect 21807 1645 22207 1671
rect 22265 1645 22665 1671
rect 22723 1645 23123 1671
rect 23181 1645 23581 1671
rect 23639 1645 24039 1671
rect 24097 1645 24497 1671
rect 24555 1645 24955 1671
rect 25013 1645 25413 1671
rect 25471 1645 25871 1671
rect 25929 1645 26329 1671
rect 26387 1645 26787 1671
rect 26845 1645 27245 1671
rect 27303 1645 27703 1671
rect 281 329 681 355
rect 739 329 1139 355
rect 1197 329 1597 355
rect 1655 329 2055 355
rect 2113 329 2513 355
rect 2571 329 2971 355
rect 3029 329 3429 355
rect 3487 329 3887 355
rect 3945 329 4345 355
rect 4403 329 4803 355
rect 4861 329 5261 355
rect 5319 329 5719 355
rect 5777 329 6177 355
rect 6235 329 6635 355
rect 6693 329 7093 355
rect 7151 329 7551 355
rect 7609 329 8009 355
rect 8067 329 8467 355
rect 8525 329 8925 355
rect 8983 329 9383 355
rect 9441 329 9841 355
rect 9899 329 10299 355
rect 10357 329 10757 355
rect 10815 329 11215 355
rect 11273 329 11673 355
rect 11731 329 12131 355
rect 12189 329 12589 355
rect 12647 329 13047 355
rect 13105 329 13505 355
rect 13563 329 13963 355
rect 14021 329 14421 355
rect 14479 329 14879 355
rect 14937 329 15337 355
rect 15395 329 15795 355
rect 15853 329 16253 355
rect 16311 329 16711 355
rect 16769 329 17169 355
rect 17227 329 17627 355
rect 17685 329 18085 355
rect 18143 329 18543 355
rect 18601 329 19001 355
rect 19059 329 19459 355
rect 19517 329 19917 355
rect 19975 329 20375 355
rect 20433 329 20833 355
rect 20891 329 21291 355
rect 21349 329 21749 355
rect 21807 329 22207 355
rect 22265 329 22665 355
rect 22723 329 23123 355
rect 23181 329 23581 355
rect 23639 329 24039 355
rect 24097 329 24497 355
rect 24555 329 24955 355
rect 25013 329 25413 355
rect 25471 329 25871 355
rect 25929 329 26329 355
rect 26387 329 26787 355
rect 26845 329 27245 355
rect 27303 329 27703 355
rect 428 184 548 329
rect 884 184 1004 329
rect 1340 184 1460 329
rect 1796 184 1916 329
rect 2252 184 2372 329
rect 2708 184 2828 329
rect 3164 184 3284 329
rect 3620 184 3740 329
rect 4076 184 4196 329
rect 4532 184 4652 329
rect 4988 184 5108 329
rect 5444 184 5564 329
rect 5900 184 6020 329
rect 6356 184 6476 329
rect 6812 184 6932 329
rect 7268 184 7388 329
rect 7724 184 7844 329
rect 8180 184 8300 329
rect 8636 184 8756 329
rect 9092 184 9212 329
rect 9548 184 9668 329
rect 10004 184 10124 329
rect 10460 184 10580 329
rect 10916 184 11036 329
rect 11372 184 11492 329
rect 11828 184 11948 329
rect 12284 184 12404 329
rect 12740 184 12860 329
rect 13196 184 13316 329
rect 13652 184 13772 329
rect 14108 184 14228 329
rect 14564 184 14684 329
rect 15020 184 15140 329
rect 15476 184 15596 329
rect 15932 184 16052 329
rect 16388 184 16508 329
rect 16844 184 16964 329
rect 17300 184 17420 329
rect 17756 184 17876 329
rect 18212 184 18332 329
rect 18668 184 18788 329
rect 19124 184 19244 329
rect 19580 184 19700 329
rect 20036 184 20156 329
rect 20492 184 20612 329
rect 20948 184 21068 329
rect 21404 184 21524 329
rect 21860 184 21980 329
rect 22316 184 22436 329
rect 22772 184 22892 329
rect 23228 184 23348 329
rect 23684 184 23804 329
rect 24140 184 24260 329
rect 24596 184 24716 329
rect 25052 184 25172 329
rect 25508 184 25628 329
rect 25964 184 26084 329
rect 26420 184 26540 329
rect 26876 184 26996 329
rect 27332 184 27452 329
rect 188 164 27796 184
rect 188 104 358 164
rect 418 104 758 164
rect 818 104 1158 164
rect 1218 104 1558 164
rect 1618 104 1958 164
rect 2018 104 2358 164
rect 2418 104 2758 164
rect 2818 104 3158 164
rect 3218 104 3558 164
rect 3618 104 3958 164
rect 4018 104 4358 164
rect 4418 104 4758 164
rect 4818 104 5158 164
rect 5218 104 5558 164
rect 5618 104 5958 164
rect 6018 104 6358 164
rect 6418 104 6758 164
rect 6818 104 7158 164
rect 7218 104 7558 164
rect 7618 104 7958 164
rect 8018 104 8358 164
rect 8418 104 8758 164
rect 8818 104 9158 164
rect 9218 104 9558 164
rect 9618 104 9958 164
rect 10018 104 10358 164
rect 10418 104 10758 164
rect 10818 104 11158 164
rect 11218 104 11558 164
rect 11618 104 11958 164
rect 12018 104 12358 164
rect 12418 104 12758 164
rect 12818 104 13158 164
rect 13218 104 13558 164
rect 13618 104 13958 164
rect 14018 104 14358 164
rect 14418 104 14758 164
rect 14818 104 15158 164
rect 15218 104 15558 164
rect 15618 104 15958 164
rect 16018 104 16358 164
rect 16418 104 16758 164
rect 16818 104 17158 164
rect 17218 104 17558 164
rect 17618 104 17958 164
rect 18018 104 18358 164
rect 18418 104 18758 164
rect 18818 104 19158 164
rect 19218 104 19558 164
rect 19618 104 19958 164
rect 20018 104 20358 164
rect 20418 104 20758 164
rect 20818 104 21158 164
rect 21218 104 21558 164
rect 21618 104 21958 164
rect 22018 104 22358 164
rect 22418 104 22758 164
rect 22818 104 23158 164
rect 23218 104 23558 164
rect 23618 104 23958 164
rect 24018 104 24358 164
rect 24418 104 24758 164
rect 24818 104 25158 164
rect 25218 104 25558 164
rect 25618 104 25958 164
rect 26018 104 26358 164
rect 26418 104 26758 164
rect 26818 104 27158 164
rect 27218 104 27558 164
rect 27618 104 27796 164
rect 188 84 27796 104
<< polycont >>
rect 358 104 418 164
rect 758 104 818 164
rect 1158 104 1218 164
rect 1558 104 1618 164
rect 1958 104 2018 164
rect 2358 104 2418 164
rect 2758 104 2818 164
rect 3158 104 3218 164
rect 3558 104 3618 164
rect 3958 104 4018 164
rect 4358 104 4418 164
rect 4758 104 4818 164
rect 5158 104 5218 164
rect 5558 104 5618 164
rect 5958 104 6018 164
rect 6358 104 6418 164
rect 6758 104 6818 164
rect 7158 104 7218 164
rect 7558 104 7618 164
rect 7958 104 8018 164
rect 8358 104 8418 164
rect 8758 104 8818 164
rect 9158 104 9218 164
rect 9558 104 9618 164
rect 9958 104 10018 164
rect 10358 104 10418 164
rect 10758 104 10818 164
rect 11158 104 11218 164
rect 11558 104 11618 164
rect 11958 104 12018 164
rect 12358 104 12418 164
rect 12758 104 12818 164
rect 13158 104 13218 164
rect 13558 104 13618 164
rect 13958 104 14018 164
rect 14358 104 14418 164
rect 14758 104 14818 164
rect 15158 104 15218 164
rect 15558 104 15618 164
rect 15958 104 16018 164
rect 16358 104 16418 164
rect 16758 104 16818 164
rect 17158 104 17218 164
rect 17558 104 17618 164
rect 17958 104 18018 164
rect 18358 104 18418 164
rect 18758 104 18818 164
rect 19158 104 19218 164
rect 19558 104 19618 164
rect 19958 104 20018 164
rect 20358 104 20418 164
rect 20758 104 20818 164
rect 21158 104 21218 164
rect 21558 104 21618 164
rect 21958 104 22018 164
rect 22358 104 22418 164
rect 22758 104 22818 164
rect 23158 104 23218 164
rect 23558 104 23618 164
rect 23958 104 24018 164
rect 24358 104 24418 164
rect 24758 104 24818 164
rect 25158 104 25218 164
rect 25558 104 25618 164
rect 25958 104 26018 164
rect 26358 104 26418 164
rect 26758 104 26818 164
rect 27158 104 27218 164
rect 27558 104 27618 164
<< locali >>
rect 90 1850 358 1910
rect 418 1850 758 1910
rect 818 1850 1158 1910
rect 1218 1850 1558 1910
rect 1618 1850 1958 1910
rect 2018 1850 2358 1910
rect 2418 1850 2758 1910
rect 2818 1850 3158 1910
rect 3218 1850 3558 1910
rect 3618 1850 3958 1910
rect 4018 1850 4358 1910
rect 4418 1850 4758 1910
rect 4818 1850 5158 1910
rect 5218 1850 5558 1910
rect 5618 1850 5958 1910
rect 6018 1850 6358 1910
rect 6418 1850 6758 1910
rect 6818 1850 7158 1910
rect 7218 1850 7558 1910
rect 7618 1850 7958 1910
rect 8018 1850 8358 1910
rect 8418 1850 8758 1910
rect 8818 1850 9158 1910
rect 9218 1850 9558 1910
rect 9618 1850 9958 1910
rect 10018 1850 10358 1910
rect 10418 1850 10758 1910
rect 10818 1850 11158 1910
rect 11218 1850 11558 1910
rect 11618 1850 11958 1910
rect 12018 1850 12358 1910
rect 12418 1850 12758 1910
rect 12818 1850 13158 1910
rect 13218 1850 13558 1910
rect 13618 1850 13958 1910
rect 14018 1850 14358 1910
rect 14418 1850 14758 1910
rect 14818 1850 15158 1910
rect 15218 1850 15558 1910
rect 15618 1850 15958 1910
rect 16018 1850 16358 1910
rect 16418 1850 16758 1910
rect 16818 1850 17158 1910
rect 17218 1850 17558 1910
rect 17618 1850 17958 1910
rect 18018 1850 18358 1910
rect 18418 1850 18758 1910
rect 18818 1850 19158 1910
rect 19218 1850 19558 1910
rect 19618 1850 19958 1910
rect 20018 1850 20358 1910
rect 20418 1850 20758 1910
rect 20818 1850 21158 1910
rect 21218 1850 21558 1910
rect 21618 1850 21958 1910
rect 22018 1850 22358 1910
rect 22418 1850 22758 1910
rect 22818 1850 23158 1910
rect 23218 1850 23558 1910
rect 23618 1850 23958 1910
rect 24018 1850 24358 1910
rect 24418 1850 24758 1910
rect 24818 1850 25158 1910
rect 25218 1850 25558 1910
rect 25618 1850 25958 1910
rect 26018 1850 26358 1910
rect 26418 1850 26758 1910
rect 26818 1850 27158 1910
rect 27218 1850 27558 1910
rect 27618 1850 27796 1910
rect 118 1760 178 1850
rect 1166 1808 1326 1850
rect 1166 1772 1226 1808
rect 1270 1772 1326 1808
rect 1166 1770 1326 1772
rect 2466 1808 2626 1850
rect 2466 1772 2526 1808
rect 2570 1772 2626 1808
rect 2466 1770 2626 1772
rect 3766 1808 3926 1850
rect 3766 1772 3826 1808
rect 3870 1772 3926 1808
rect 3766 1770 3926 1772
rect 5066 1808 5226 1850
rect 5066 1772 5126 1808
rect 5170 1772 5226 1808
rect 5066 1770 5226 1772
rect 6366 1808 6526 1850
rect 6366 1772 6426 1808
rect 6470 1772 6526 1808
rect 6366 1770 6526 1772
rect 7666 1808 7826 1850
rect 7666 1772 7726 1808
rect 7770 1772 7826 1808
rect 7666 1770 7826 1772
rect 8966 1808 9126 1850
rect 8966 1772 9026 1808
rect 9070 1772 9126 1808
rect 8966 1770 9126 1772
rect 10266 1808 10426 1850
rect 10266 1772 10326 1808
rect 10370 1772 10426 1808
rect 10266 1770 10426 1772
rect 11566 1808 11726 1850
rect 11566 1772 11626 1808
rect 11670 1772 11726 1808
rect 11566 1770 11726 1772
rect 12866 1808 13026 1850
rect 12866 1772 12926 1808
rect 12970 1772 13026 1808
rect 12866 1770 13026 1772
rect 14166 1808 14326 1850
rect 14166 1772 14226 1808
rect 14270 1772 14326 1808
rect 14166 1770 14326 1772
rect 15466 1808 15626 1850
rect 15466 1772 15526 1808
rect 15570 1772 15626 1808
rect 15466 1770 15626 1772
rect 16766 1808 16926 1850
rect 16766 1772 16826 1808
rect 16870 1772 16926 1808
rect 16766 1770 16926 1772
rect 18066 1808 18226 1850
rect 18066 1772 18126 1808
rect 18170 1772 18226 1808
rect 18066 1770 18226 1772
rect 19366 1808 19526 1850
rect 19366 1772 19426 1808
rect 19470 1772 19526 1808
rect 19366 1770 19526 1772
rect 20666 1808 20826 1850
rect 20666 1772 20726 1808
rect 20770 1772 20826 1808
rect 20666 1770 20826 1772
rect 21966 1808 22126 1850
rect 21966 1772 22026 1808
rect 22070 1772 22126 1808
rect 21966 1770 22126 1772
rect 23266 1808 23426 1850
rect 23266 1772 23326 1808
rect 23370 1772 23426 1808
rect 23266 1770 23426 1772
rect 24566 1808 24726 1850
rect 24566 1772 24626 1808
rect 24670 1772 24726 1808
rect 24566 1770 24726 1772
rect 25866 1808 26026 1850
rect 25866 1772 25926 1808
rect 25970 1772 26026 1808
rect 25866 1770 26026 1772
rect 118 1720 128 1760
rect 168 1720 178 1760
rect 118 1640 178 1720
rect 248 1690 27796 1730
rect 235 1633 269 1649
rect 235 270 269 367
rect 693 1633 727 1690
rect 693 351 727 367
rect 1151 1633 1185 1649
rect 1151 270 1185 367
rect 1609 1633 1643 1690
rect 1609 351 1643 367
rect 2067 1633 2101 1649
rect 2067 270 2101 367
rect 2525 1633 2559 1690
rect 2525 351 2559 367
rect 2983 1633 3017 1649
rect 2983 270 3017 367
rect 3441 1633 3475 1690
rect 3441 351 3475 367
rect 3899 1633 3933 1649
rect 3899 270 3933 367
rect 4357 1633 4391 1690
rect 4357 351 4391 367
rect 4815 1633 4849 1649
rect 4815 270 4849 367
rect 5273 1633 5307 1690
rect 5273 351 5307 367
rect 5731 1633 5765 1649
rect 5731 270 5765 367
rect 6189 1633 6223 1690
rect 6189 351 6223 367
rect 6647 1633 6681 1649
rect 6647 270 6681 367
rect 7105 1633 7139 1690
rect 7105 351 7139 367
rect 7563 1633 7597 1649
rect 7563 270 7597 367
rect 8021 1633 8055 1690
rect 8021 351 8055 367
rect 8479 1633 8513 1649
rect 8479 270 8513 367
rect 8937 1633 8971 1690
rect 8937 351 8971 367
rect 9395 1633 9429 1649
rect 9395 270 9429 367
rect 9853 1633 9887 1690
rect 9853 351 9887 367
rect 10311 1633 10345 1649
rect 10311 270 10345 367
rect 10769 1633 10803 1690
rect 10769 351 10803 367
rect 11227 1633 11261 1649
rect 11227 270 11261 367
rect 11685 1633 11719 1690
rect 11685 351 11719 367
rect 12143 1633 12177 1649
rect 12143 270 12177 367
rect 12601 1633 12635 1690
rect 12601 351 12635 367
rect 13059 1633 13093 1649
rect 13059 270 13093 367
rect 13517 1633 13551 1690
rect 13517 351 13551 367
rect 13975 1633 14009 1649
rect 13975 270 14009 367
rect 14433 1633 14467 1690
rect 14433 351 14467 367
rect 14891 1633 14925 1649
rect 14891 270 14925 367
rect 15349 1633 15383 1690
rect 15349 351 15383 367
rect 15807 1633 15841 1649
rect 15807 270 15841 367
rect 16265 1633 16299 1690
rect 16265 351 16299 367
rect 16723 1633 16757 1649
rect 16723 270 16757 367
rect 17181 1633 17215 1690
rect 17181 351 17215 367
rect 17639 1633 17673 1649
rect 17639 270 17673 367
rect 18097 1633 18131 1690
rect 18097 351 18131 367
rect 18555 1633 18589 1649
rect 18555 270 18589 367
rect 19013 1633 19047 1690
rect 19013 351 19047 367
rect 19471 1633 19505 1649
rect 19471 270 19505 367
rect 19929 1633 19963 1690
rect 19929 351 19963 367
rect 20387 1633 20421 1649
rect 20387 270 20421 367
rect 20845 1633 20879 1690
rect 20845 351 20879 367
rect 21303 1633 21337 1649
rect 21303 270 21337 367
rect 21761 1633 21795 1690
rect 21761 351 21795 367
rect 22219 1633 22253 1649
rect 22219 270 22253 367
rect 22677 1633 22711 1690
rect 22677 351 22711 367
rect 23135 1633 23169 1649
rect 23135 270 23169 367
rect 23593 1633 23627 1690
rect 23593 351 23627 367
rect 24051 1633 24085 1649
rect 24051 270 24085 367
rect 24509 1633 24543 1690
rect 24509 351 24543 367
rect 24967 1633 25001 1649
rect 24967 270 25001 367
rect 25425 1633 25459 1690
rect 25425 351 25459 367
rect 25883 1633 25917 1649
rect 25883 270 25917 367
rect 26341 1633 26375 1690
rect 26341 351 26375 367
rect 26799 1633 26833 1649
rect 26799 270 26833 367
rect 27257 1633 27291 1690
rect 27257 351 27291 367
rect 27715 1633 27749 1649
rect 27715 270 27749 367
rect 188 210 27796 270
rect 188 104 358 164
rect 418 104 758 164
rect 818 104 1158 164
rect 1218 104 1558 164
rect 1618 104 1958 164
rect 2018 104 2358 164
rect 2418 104 2758 164
rect 2818 104 3158 164
rect 3218 104 3558 164
rect 3618 104 3958 164
rect 4018 104 4358 164
rect 4418 104 4758 164
rect 4818 104 5158 164
rect 5218 104 5558 164
rect 5618 104 5958 164
rect 6018 104 6358 164
rect 6418 104 6758 164
rect 6818 104 7158 164
rect 7218 104 7558 164
rect 7618 104 7958 164
rect 8018 104 8358 164
rect 8418 104 8758 164
rect 8818 104 9158 164
rect 9218 104 9558 164
rect 9618 104 9958 164
rect 10018 104 10358 164
rect 10418 104 10758 164
rect 10818 104 11158 164
rect 11218 104 11558 164
rect 11618 104 11958 164
rect 12018 104 12358 164
rect 12418 104 12758 164
rect 12818 104 13158 164
rect 13218 104 13558 164
rect 13618 104 13958 164
rect 14018 104 14358 164
rect 14418 104 14758 164
rect 14818 104 15158 164
rect 15218 104 15558 164
rect 15618 104 15958 164
rect 16018 104 16358 164
rect 16418 104 16758 164
rect 16818 104 17158 164
rect 17218 104 17558 164
rect 17618 104 17958 164
rect 18018 104 18358 164
rect 18418 104 18758 164
rect 18818 104 19158 164
rect 19218 104 19558 164
rect 19618 104 19958 164
rect 20018 104 20358 164
rect 20418 104 20758 164
rect 20818 104 21158 164
rect 21218 104 21558 164
rect 21618 104 21958 164
rect 22018 104 22358 164
rect 22418 104 22758 164
rect 22818 104 23158 164
rect 23218 104 23558 164
rect 23618 104 23958 164
rect 24018 104 24358 164
rect 24418 104 24758 164
rect 24818 104 25158 164
rect 25218 104 25558 164
rect 25618 104 25958 164
rect 26018 104 26358 164
rect 26418 104 26758 164
rect 26818 104 27158 164
rect 27218 104 27558 164
rect 27618 104 27796 164
rect 90 -30 358 30
rect 418 -30 758 30
rect 818 -30 1158 30
rect 1218 -30 1558 30
rect 1618 -30 1958 30
rect 2018 -30 2358 30
rect 2418 -30 2758 30
rect 2818 -30 3158 30
rect 3218 -30 3558 30
rect 3618 -30 3958 30
rect 4018 -30 4358 30
rect 4418 -30 4758 30
rect 4818 -30 5158 30
rect 5218 -30 5558 30
rect 5618 -30 5958 30
rect 6018 -30 6358 30
rect 6418 -30 6758 30
rect 6818 -30 7158 30
rect 7218 -30 7558 30
rect 7618 -30 7958 30
rect 8018 -30 8358 30
rect 8418 -30 8758 30
rect 8818 -30 9158 30
rect 9218 -30 9558 30
rect 9618 -30 9958 30
rect 10018 -30 10358 30
rect 10418 -30 10758 30
rect 10818 -30 11158 30
rect 11218 -30 11558 30
rect 11618 -30 11958 30
rect 12018 -30 12358 30
rect 12418 -30 12758 30
rect 12818 -30 13158 30
rect 13218 -30 13558 30
rect 13618 -30 13958 30
rect 14018 -30 14358 30
rect 14418 -30 14758 30
rect 14818 -30 15158 30
rect 15218 -30 15558 30
rect 15618 -30 15958 30
rect 16018 -30 16358 30
rect 16418 -30 16758 30
rect 16818 -30 17158 30
rect 17218 -30 17558 30
rect 17618 -30 17958 30
rect 18018 -30 18358 30
rect 18418 -30 18758 30
rect 18818 -30 19158 30
rect 19218 -30 19558 30
rect 19618 -30 19958 30
rect 20018 -30 20358 30
rect 20418 -30 20758 30
rect 20818 -30 21158 30
rect 21218 -30 21558 30
rect 21618 -30 21958 30
rect 22018 -30 22358 30
rect 22418 -30 22758 30
rect 22818 -30 23158 30
rect 23218 -30 23558 30
rect 23618 -30 23958 30
rect 24018 -30 24358 30
rect 24418 -30 24758 30
rect 24818 -30 25158 30
rect 25218 -30 25558 30
rect 25618 -30 25958 30
rect 26018 -30 26358 30
rect 26418 -30 26758 30
rect 26818 -30 27158 30
rect 27218 -30 27558 30
rect 27618 -30 27796 30
<< viali >>
rect 358 1850 418 1910
rect 758 1850 818 1910
rect 1158 1850 1218 1910
rect 1558 1850 1618 1910
rect 1958 1850 2018 1910
rect 2358 1850 2418 1910
rect 2758 1850 2818 1910
rect 3158 1850 3218 1910
rect 3558 1850 3618 1910
rect 3958 1850 4018 1910
rect 4358 1850 4418 1910
rect 4758 1850 4818 1910
rect 5158 1850 5218 1910
rect 5558 1850 5618 1910
rect 5958 1850 6018 1910
rect 6358 1850 6418 1910
rect 6758 1850 6818 1910
rect 7158 1850 7218 1910
rect 7558 1850 7618 1910
rect 7958 1850 8018 1910
rect 8358 1850 8418 1910
rect 8758 1850 8818 1910
rect 9158 1850 9218 1910
rect 9558 1850 9618 1910
rect 9958 1850 10018 1910
rect 10358 1850 10418 1910
rect 10758 1850 10818 1910
rect 11158 1850 11218 1910
rect 11558 1850 11618 1910
rect 11958 1850 12018 1910
rect 12358 1850 12418 1910
rect 12758 1850 12818 1910
rect 13158 1850 13218 1910
rect 13558 1850 13618 1910
rect 13958 1850 14018 1910
rect 14358 1850 14418 1910
rect 14758 1850 14818 1910
rect 15158 1850 15218 1910
rect 15558 1850 15618 1910
rect 15958 1850 16018 1910
rect 16358 1850 16418 1910
rect 16758 1850 16818 1910
rect 17158 1850 17218 1910
rect 17558 1850 17618 1910
rect 17958 1850 18018 1910
rect 18358 1850 18418 1910
rect 18758 1850 18818 1910
rect 19158 1850 19218 1910
rect 19558 1850 19618 1910
rect 19958 1850 20018 1910
rect 20358 1850 20418 1910
rect 20758 1850 20818 1910
rect 21158 1850 21218 1910
rect 21558 1850 21618 1910
rect 21958 1850 22018 1910
rect 22358 1850 22418 1910
rect 22758 1850 22818 1910
rect 23158 1850 23218 1910
rect 23558 1850 23618 1910
rect 23958 1850 24018 1910
rect 24358 1850 24418 1910
rect 24758 1850 24818 1910
rect 25158 1850 25218 1910
rect 25558 1850 25618 1910
rect 25958 1850 26018 1910
rect 26358 1850 26418 1910
rect 26758 1850 26818 1910
rect 27158 1850 27218 1910
rect 27558 1850 27618 1910
rect 235 367 269 1633
rect 693 367 727 1633
rect 1151 367 1185 1633
rect 1609 367 1643 1633
rect 2067 367 2101 1633
rect 2525 367 2559 1633
rect 2983 367 3017 1633
rect 3441 367 3475 1633
rect 3899 367 3933 1633
rect 4357 367 4391 1633
rect 4815 367 4849 1633
rect 5273 367 5307 1633
rect 5731 367 5765 1633
rect 6189 367 6223 1633
rect 6647 367 6681 1633
rect 7105 367 7139 1633
rect 7563 367 7597 1633
rect 8021 367 8055 1633
rect 8479 367 8513 1633
rect 8937 367 8971 1633
rect 9395 367 9429 1633
rect 9853 367 9887 1633
rect 10311 367 10345 1633
rect 10769 367 10803 1633
rect 11227 367 11261 1633
rect 11685 367 11719 1633
rect 12143 367 12177 1633
rect 12601 367 12635 1633
rect 13059 367 13093 1633
rect 13517 367 13551 1633
rect 13975 367 14009 1633
rect 14433 367 14467 1633
rect 14891 367 14925 1633
rect 15349 367 15383 1633
rect 15807 367 15841 1633
rect 16265 367 16299 1633
rect 16723 367 16757 1633
rect 17181 367 17215 1633
rect 17639 367 17673 1633
rect 18097 367 18131 1633
rect 18555 367 18589 1633
rect 19013 367 19047 1633
rect 19471 367 19505 1633
rect 19929 367 19963 1633
rect 20387 367 20421 1633
rect 20845 367 20879 1633
rect 21303 367 21337 1633
rect 21761 367 21795 1633
rect 22219 367 22253 1633
rect 22677 367 22711 1633
rect 23135 367 23169 1633
rect 23593 367 23627 1633
rect 24051 367 24085 1633
rect 24509 367 24543 1633
rect 24967 367 25001 1633
rect 25425 367 25459 1633
rect 25883 367 25917 1633
rect 26341 367 26375 1633
rect 26799 367 26833 1633
rect 27257 367 27291 1633
rect 27715 367 27749 1633
rect 358 -30 418 30
rect 758 -30 818 30
rect 1158 -30 1218 30
rect 1558 -30 1618 30
rect 1958 -30 2018 30
rect 2358 -30 2418 30
rect 2758 -30 2818 30
rect 3158 -30 3218 30
rect 3558 -30 3618 30
rect 3958 -30 4018 30
rect 4358 -30 4418 30
rect 4758 -30 4818 30
rect 5158 -30 5218 30
rect 5558 -30 5618 30
rect 5958 -30 6018 30
rect 6358 -30 6418 30
rect 6758 -30 6818 30
rect 7158 -30 7218 30
rect 7558 -30 7618 30
rect 7958 -30 8018 30
rect 8358 -30 8418 30
rect 8758 -30 8818 30
rect 9158 -30 9218 30
rect 9558 -30 9618 30
rect 9958 -30 10018 30
rect 10358 -30 10418 30
rect 10758 -30 10818 30
rect 11158 -30 11218 30
rect 11558 -30 11618 30
rect 11958 -30 12018 30
rect 12358 -30 12418 30
rect 12758 -30 12818 30
rect 13158 -30 13218 30
rect 13558 -30 13618 30
rect 13958 -30 14018 30
rect 14358 -30 14418 30
rect 14758 -30 14818 30
rect 15158 -30 15218 30
rect 15558 -30 15618 30
rect 15958 -30 16018 30
rect 16358 -30 16418 30
rect 16758 -30 16818 30
rect 17158 -30 17218 30
rect 17558 -30 17618 30
rect 17958 -30 18018 30
rect 18358 -30 18418 30
rect 18758 -30 18818 30
rect 19158 -30 19218 30
rect 19558 -30 19618 30
rect 19958 -30 20018 30
rect 20358 -30 20418 30
rect 20758 -30 20818 30
rect 21158 -30 21218 30
rect 21558 -30 21618 30
rect 21958 -30 22018 30
rect 22358 -30 22418 30
rect 22758 -30 22818 30
rect 23158 -30 23218 30
rect 23558 -30 23618 30
rect 23958 -30 24018 30
rect 24358 -30 24418 30
rect 24758 -30 24818 30
rect 25158 -30 25218 30
rect 25558 -30 25618 30
rect 25958 -30 26018 30
rect 26358 -30 26418 30
rect 26758 -30 26818 30
rect 27158 -30 27218 30
rect 27558 -30 27618 30
<< metal1 >>
rect 90 1910 27796 1940
rect 90 1850 358 1910
rect 418 1850 758 1910
rect 818 1850 1158 1910
rect 1218 1850 1558 1910
rect 1618 1850 1958 1910
rect 2018 1850 2358 1910
rect 2418 1850 2758 1910
rect 2818 1850 3158 1910
rect 3218 1850 3558 1910
rect 3618 1850 3958 1910
rect 4018 1850 4358 1910
rect 4418 1850 4758 1910
rect 4818 1850 5158 1910
rect 5218 1850 5558 1910
rect 5618 1850 5958 1910
rect 6018 1850 6358 1910
rect 6418 1850 6758 1910
rect 6818 1850 7158 1910
rect 7218 1850 7558 1910
rect 7618 1850 7958 1910
rect 8018 1850 8358 1910
rect 8418 1850 8758 1910
rect 8818 1850 9158 1910
rect 9218 1850 9558 1910
rect 9618 1850 9958 1910
rect 10018 1850 10358 1910
rect 10418 1850 10758 1910
rect 10818 1850 11158 1910
rect 11218 1850 11558 1910
rect 11618 1850 11958 1910
rect 12018 1850 12358 1910
rect 12418 1850 12758 1910
rect 12818 1850 13158 1910
rect 13218 1850 13558 1910
rect 13618 1850 13958 1910
rect 14018 1850 14358 1910
rect 14418 1850 14758 1910
rect 14818 1850 15158 1910
rect 15218 1850 15558 1910
rect 15618 1850 15958 1910
rect 16018 1850 16358 1910
rect 16418 1850 16758 1910
rect 16818 1850 17158 1910
rect 17218 1850 17558 1910
rect 17618 1850 17958 1910
rect 18018 1850 18358 1910
rect 18418 1850 18758 1910
rect 18818 1850 19158 1910
rect 19218 1850 19558 1910
rect 19618 1850 19958 1910
rect 20018 1850 20358 1910
rect 20418 1850 20758 1910
rect 20818 1850 21158 1910
rect 21218 1850 21558 1910
rect 21618 1850 21958 1910
rect 22018 1850 22358 1910
rect 22418 1850 22758 1910
rect 22818 1850 23158 1910
rect 23218 1850 23558 1910
rect 23618 1850 23958 1910
rect 24018 1850 24358 1910
rect 24418 1850 24758 1910
rect 24818 1850 25158 1910
rect 25218 1850 25558 1910
rect 25618 1850 25958 1910
rect 26018 1850 26358 1910
rect 26418 1850 26758 1910
rect 26818 1850 27158 1910
rect 27218 1850 27558 1910
rect 27618 1850 27796 1910
rect 90 1820 27796 1850
rect 229 1633 275 1645
rect 229 367 235 1633
rect 269 367 275 1633
rect 229 355 275 367
rect 687 1633 733 1645
rect 687 367 693 1633
rect 727 367 733 1633
rect 687 355 733 367
rect 1145 1633 1191 1645
rect 1145 367 1151 1633
rect 1185 367 1191 1633
rect 1145 355 1191 367
rect 1603 1633 1649 1645
rect 1603 367 1609 1633
rect 1643 367 1649 1633
rect 1603 355 1649 367
rect 2061 1633 2107 1645
rect 2061 367 2067 1633
rect 2101 367 2107 1633
rect 2061 355 2107 367
rect 2519 1633 2565 1645
rect 2519 367 2525 1633
rect 2559 367 2565 1633
rect 2519 355 2565 367
rect 2977 1633 3023 1645
rect 2977 367 2983 1633
rect 3017 367 3023 1633
rect 2977 355 3023 367
rect 3435 1633 3481 1645
rect 3435 367 3441 1633
rect 3475 367 3481 1633
rect 3435 355 3481 367
rect 3893 1633 3939 1645
rect 3893 367 3899 1633
rect 3933 367 3939 1633
rect 3893 355 3939 367
rect 4351 1633 4397 1645
rect 4351 367 4357 1633
rect 4391 367 4397 1633
rect 4351 355 4397 367
rect 4809 1633 4855 1645
rect 4809 367 4815 1633
rect 4849 367 4855 1633
rect 4809 355 4855 367
rect 5267 1633 5313 1645
rect 5267 367 5273 1633
rect 5307 367 5313 1633
rect 5267 355 5313 367
rect 5725 1633 5771 1645
rect 5725 367 5731 1633
rect 5765 367 5771 1633
rect 5725 355 5771 367
rect 6183 1633 6229 1645
rect 6183 367 6189 1633
rect 6223 367 6229 1633
rect 6183 355 6229 367
rect 6641 1633 6687 1645
rect 6641 367 6647 1633
rect 6681 367 6687 1633
rect 6641 355 6687 367
rect 7099 1633 7145 1645
rect 7099 367 7105 1633
rect 7139 367 7145 1633
rect 7099 355 7145 367
rect 7557 1633 7603 1645
rect 7557 367 7563 1633
rect 7597 367 7603 1633
rect 7557 355 7603 367
rect 8015 1633 8061 1645
rect 8015 367 8021 1633
rect 8055 367 8061 1633
rect 8015 355 8061 367
rect 8473 1633 8519 1645
rect 8473 367 8479 1633
rect 8513 367 8519 1633
rect 8473 355 8519 367
rect 8931 1633 8977 1645
rect 8931 367 8937 1633
rect 8971 367 8977 1633
rect 8931 355 8977 367
rect 9389 1633 9435 1645
rect 9389 367 9395 1633
rect 9429 367 9435 1633
rect 9389 355 9435 367
rect 9847 1633 9893 1645
rect 9847 367 9853 1633
rect 9887 367 9893 1633
rect 9847 355 9893 367
rect 10305 1633 10351 1645
rect 10305 367 10311 1633
rect 10345 367 10351 1633
rect 10305 355 10351 367
rect 10763 1633 10809 1645
rect 10763 367 10769 1633
rect 10803 367 10809 1633
rect 10763 355 10809 367
rect 11221 1633 11267 1645
rect 11221 367 11227 1633
rect 11261 367 11267 1633
rect 11221 355 11267 367
rect 11679 1633 11725 1645
rect 11679 367 11685 1633
rect 11719 367 11725 1633
rect 11679 355 11725 367
rect 12137 1633 12183 1645
rect 12137 367 12143 1633
rect 12177 367 12183 1633
rect 12137 355 12183 367
rect 12595 1633 12641 1645
rect 12595 367 12601 1633
rect 12635 367 12641 1633
rect 12595 355 12641 367
rect 13053 1633 13099 1645
rect 13053 367 13059 1633
rect 13093 367 13099 1633
rect 13053 355 13099 367
rect 13511 1633 13557 1645
rect 13511 367 13517 1633
rect 13551 367 13557 1633
rect 13511 355 13557 367
rect 13969 1633 14015 1645
rect 13969 367 13975 1633
rect 14009 367 14015 1633
rect 13969 355 14015 367
rect 14427 1633 14473 1645
rect 14427 367 14433 1633
rect 14467 367 14473 1633
rect 14427 355 14473 367
rect 14885 1633 14931 1645
rect 14885 367 14891 1633
rect 14925 367 14931 1633
rect 14885 355 14931 367
rect 15343 1633 15389 1645
rect 15343 367 15349 1633
rect 15383 367 15389 1633
rect 15343 355 15389 367
rect 15801 1633 15847 1645
rect 15801 367 15807 1633
rect 15841 367 15847 1633
rect 15801 355 15847 367
rect 16259 1633 16305 1645
rect 16259 367 16265 1633
rect 16299 367 16305 1633
rect 16259 355 16305 367
rect 16717 1633 16763 1645
rect 16717 367 16723 1633
rect 16757 367 16763 1633
rect 16717 355 16763 367
rect 17175 1633 17221 1645
rect 17175 367 17181 1633
rect 17215 367 17221 1633
rect 17175 355 17221 367
rect 17633 1633 17679 1645
rect 17633 367 17639 1633
rect 17673 367 17679 1633
rect 17633 355 17679 367
rect 18091 1633 18137 1645
rect 18091 367 18097 1633
rect 18131 367 18137 1633
rect 18091 355 18137 367
rect 18549 1633 18595 1645
rect 18549 367 18555 1633
rect 18589 367 18595 1633
rect 18549 355 18595 367
rect 19007 1633 19053 1645
rect 19007 367 19013 1633
rect 19047 367 19053 1633
rect 19007 355 19053 367
rect 19465 1633 19511 1645
rect 19465 367 19471 1633
rect 19505 367 19511 1633
rect 19465 355 19511 367
rect 19923 1633 19969 1645
rect 19923 367 19929 1633
rect 19963 367 19969 1633
rect 19923 355 19969 367
rect 20381 1633 20427 1645
rect 20381 367 20387 1633
rect 20421 367 20427 1633
rect 20381 355 20427 367
rect 20839 1633 20885 1645
rect 20839 367 20845 1633
rect 20879 367 20885 1633
rect 20839 355 20885 367
rect 21297 1633 21343 1645
rect 21297 367 21303 1633
rect 21337 367 21343 1633
rect 21297 355 21343 367
rect 21755 1633 21801 1645
rect 21755 367 21761 1633
rect 21795 367 21801 1633
rect 21755 355 21801 367
rect 22213 1633 22259 1645
rect 22213 367 22219 1633
rect 22253 367 22259 1633
rect 22213 355 22259 367
rect 22671 1633 22717 1645
rect 22671 367 22677 1633
rect 22711 367 22717 1633
rect 22671 355 22717 367
rect 23129 1633 23175 1645
rect 23129 367 23135 1633
rect 23169 367 23175 1633
rect 23129 355 23175 367
rect 23587 1633 23633 1645
rect 23587 367 23593 1633
rect 23627 367 23633 1633
rect 23587 355 23633 367
rect 24045 1633 24091 1645
rect 24045 367 24051 1633
rect 24085 367 24091 1633
rect 24045 355 24091 367
rect 24503 1633 24549 1645
rect 24503 367 24509 1633
rect 24543 367 24549 1633
rect 24503 355 24549 367
rect 24961 1633 25007 1645
rect 24961 367 24967 1633
rect 25001 367 25007 1633
rect 24961 355 25007 367
rect 25419 1633 25465 1645
rect 25419 367 25425 1633
rect 25459 367 25465 1633
rect 25419 355 25465 367
rect 25877 1633 25923 1645
rect 25877 367 25883 1633
rect 25917 367 25923 1633
rect 25877 355 25923 367
rect 26335 1633 26381 1645
rect 26335 367 26341 1633
rect 26375 367 26381 1633
rect 26335 355 26381 367
rect 26793 1633 26839 1645
rect 26793 367 26799 1633
rect 26833 367 26839 1633
rect 26793 355 26839 367
rect 27251 1633 27297 1645
rect 27251 367 27257 1633
rect 27291 367 27297 1633
rect 27251 355 27297 367
rect 27709 1633 27755 1645
rect 27709 367 27715 1633
rect 27749 367 27755 1633
rect 27709 355 27755 367
rect 90 30 27796 60
rect 90 -30 358 30
rect 418 -30 758 30
rect 818 -30 1158 30
rect 1218 -30 1558 30
rect 1618 -30 1958 30
rect 2018 -30 2358 30
rect 2418 -30 2758 30
rect 2818 -30 3158 30
rect 3218 -30 3558 30
rect 3618 -30 3958 30
rect 4018 -30 4358 30
rect 4418 -30 4758 30
rect 4818 -30 5158 30
rect 5218 -30 5558 30
rect 5618 -30 5958 30
rect 6018 -30 6358 30
rect 6418 -30 6758 30
rect 6818 -30 7158 30
rect 7218 -30 7558 30
rect 7618 -30 7958 30
rect 8018 -30 8358 30
rect 8418 -30 8758 30
rect 8818 -30 9158 30
rect 9218 -30 9558 30
rect 9618 -30 9958 30
rect 10018 -30 10358 30
rect 10418 -30 10758 30
rect 10818 -30 11158 30
rect 11218 -30 11558 30
rect 11618 -30 11958 30
rect 12018 -30 12358 30
rect 12418 -30 12758 30
rect 12818 -30 13158 30
rect 13218 -30 13558 30
rect 13618 -30 13958 30
rect 14018 -30 14358 30
rect 14418 -30 14758 30
rect 14818 -30 15158 30
rect 15218 -30 15558 30
rect 15618 -30 15958 30
rect 16018 -30 16358 30
rect 16418 -30 16758 30
rect 16818 -30 17158 30
rect 17218 -30 17558 30
rect 17618 -30 17958 30
rect 18018 -30 18358 30
rect 18418 -30 18758 30
rect 18818 -30 19158 30
rect 19218 -30 19558 30
rect 19618 -30 19958 30
rect 20018 -30 20358 30
rect 20418 -30 20758 30
rect 20818 -30 21158 30
rect 21218 -30 21558 30
rect 21618 -30 21958 30
rect 22018 -30 22358 30
rect 22418 -30 22758 30
rect 22818 -30 23158 30
rect 23218 -30 23558 30
rect 23618 -30 23958 30
rect 24018 -30 24358 30
rect 24418 -30 24758 30
rect 24818 -30 25158 30
rect 25218 -30 25558 30
rect 25618 -30 25958 30
rect 26018 -30 26358 30
rect 26418 -30 26758 30
rect 26818 -30 27158 30
rect 27218 -30 27558 30
rect 27618 -30 27796 30
rect 90 -60 27796 -30
<< labels >>
flabel nwell 90 1850 150 1910 1 FreeSans 800 0 0 0 VPWR
port 4 n power bidirectional
flabel metal1 90 -30 248 30 1 FreeSans 800 0 0 0 VGND
port 5 n ground bidirectional
flabel locali 27736 1690 27796 1730 1 FreeSans 800 0 0 0 SOURCE
port 2 n signal bidirectional
flabel locali 27736 210 27796 270 1 FreeSans 800 0 0 0 DRAIN
port 3 n signal bidirectional
flabel locali 27736 104 27796 164 1 FreeSans 800 0 0 0 GATE
port 1 n signal bidirectional
<< properties >>
string FIXED_BBOX 0 0 27887 1880
string LEFclass CORE
string LEFsite unitasc
<< end >>
