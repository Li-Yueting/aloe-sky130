magic
tech sky130A
magscale 1 2
timestamp 1653532055
<< pwell >>
rect 428 -60 2868 1650
<< psubdiff >>
rect 1340 940 1956 970
rect 1340 820 1400 940
rect 1896 820 1956 940
rect 1340 790 1956 820
<< psubdiffcont >>
rect 1400 820 1896 940
<< xpolycontact >>
rect 141 1075 573 1645
rect 2723 1075 3155 1645
rect 141 115 573 685
rect 2723 115 3155 685
<< xpolyres >>
rect 573 1075 2723 1645
rect 573 115 2723 685
<< locali >>
rect 142 1850 312 1910
rect 372 1850 512 1910
rect 572 1850 712 1910
rect 772 1850 912 1910
rect 972 1850 1112 1910
rect 1172 1850 1312 1910
rect 1372 1850 1512 1910
rect 1572 1850 1712 1910
rect 1772 1850 1912 1910
rect 1972 1850 2112 1910
rect 2172 1850 2312 1910
rect 2372 1850 2512 1910
rect 2572 1850 2712 1910
rect 2772 1850 2912 1910
rect 2972 1850 3154 1910
rect 1340 940 1956 970
rect 1340 820 1400 940
rect 1896 820 1956 940
rect 1340 30 1956 820
rect 2723 685 3155 1075
rect 142 -30 312 30
rect 372 -30 512 30
rect 572 -30 712 30
rect 772 -30 912 30
rect 972 -30 1112 30
rect 1172 -30 1312 30
rect 1372 -30 1512 30
rect 1572 -30 1712 30
rect 1772 -30 1912 30
rect 1972 -30 2112 30
rect 2172 -30 2312 30
rect 2372 -30 2512 30
rect 2572 -30 2712 30
rect 2772 -30 2912 30
rect 2972 -30 3154 30
<< viali >>
rect 312 1850 372 1910
rect 512 1850 572 1910
rect 712 1850 772 1910
rect 912 1850 972 1910
rect 1112 1850 1172 1910
rect 1312 1850 1372 1910
rect 1512 1850 1572 1910
rect 1712 1850 1772 1910
rect 1912 1850 1972 1910
rect 2112 1850 2172 1910
rect 2312 1850 2372 1910
rect 2512 1850 2572 1910
rect 2712 1850 2772 1910
rect 2912 1850 2972 1910
rect 159 1091 556 1629
rect 2740 1091 3137 1629
rect 159 131 556 669
rect 2740 131 3137 669
rect 312 -30 372 30
rect 512 -30 572 30
rect 712 -30 772 30
rect 912 -30 972 30
rect 1112 -30 1172 30
rect 1312 -30 1372 30
rect 1512 -30 1572 30
rect 1712 -30 1772 30
rect 1912 -30 1972 30
rect 2112 -30 2172 30
rect 2312 -30 2372 30
rect 2512 -30 2572 30
rect 2712 -30 2772 30
rect 2912 -30 2972 30
<< metal1 >>
rect 142 1910 3154 1940
rect 142 1850 312 1910
rect 372 1850 512 1910
rect 572 1850 712 1910
rect 772 1850 912 1910
rect 972 1850 1112 1910
rect 1172 1850 1312 1910
rect 1372 1850 1512 1910
rect 1572 1850 1712 1910
rect 1772 1850 1912 1910
rect 1972 1850 2112 1910
rect 2172 1850 2312 1910
rect 2372 1850 2512 1910
rect 2572 1850 2712 1910
rect 2772 1850 2912 1910
rect 2972 1850 3154 1910
rect 142 1820 3154 1850
rect 152 1629 562 1641
rect 152 1091 159 1629
rect 556 1091 562 1629
rect 152 1079 562 1091
rect 2734 1629 3144 1641
rect 2734 1091 2740 1629
rect 3137 1091 3144 1629
rect 2734 1079 3144 1091
rect 152 669 562 681
rect 152 131 159 669
rect 556 131 562 669
rect 152 119 562 131
rect 2723 669 3155 1079
rect 2723 131 2740 669
rect 3137 131 3155 669
rect 2723 115 3155 131
rect 142 30 3154 60
rect 142 -30 312 30
rect 372 -30 512 30
rect 572 -30 712 30
rect 772 -30 912 30
rect 972 -30 1112 30
rect 1172 -30 1312 30
rect 1372 -30 1512 30
rect 1572 -30 1712 30
rect 1772 -30 1912 30
rect 1972 -30 2112 30
rect 2172 -30 2312 30
rect 2372 -30 2512 30
rect 2572 -30 2712 30
rect 2772 -30 2912 30
rect 2972 -30 3154 30
rect 142 -60 3154 -30
<< labels >>
flabel metal1 261 1300 381 1420 1 FreeSans 480 0 0 0 Rin
port 1 n default bidirectional
flabel metal1 261 340 381 460 1 FreeSans 480 0 0 0 Rout
port 2 n default bidirectional
flabel metal1 142 1850 202 1910 1 FreeSans 800 0 0 0 VPWR
port 3 n power bidirectional
flabel metal1 142 -30 202 30 1 FreeSans 800 0 0 0 VGND
port 4 n ground bidirectional
<< properties >>
string FIXED_BBOX 0 0 3294 1880
string LEFclass CORE
string LEFsite unitasc
<< end >>
