magic
tech sky130A
magscale 1 2
timestamp 1651893041
<< nwell >>
rect 0 293 4252 1940
<< pmoslvt >>
rect 94 355 494 1645
rect 552 355 952 1645
rect 1010 355 1410 1645
rect 1468 355 1868 1645
rect 1926 355 2326 1645
rect 2384 355 2784 1645
rect 2842 355 3242 1645
rect 3300 355 3700 1645
rect 3758 355 4158 1645
<< pdiff >>
rect 36 1633 94 1645
rect 36 367 48 1633
rect 82 367 94 1633
rect 36 355 94 367
rect 494 1633 552 1645
rect 494 367 506 1633
rect 540 367 552 1633
rect 494 355 552 367
rect 952 1633 1010 1645
rect 952 367 964 1633
rect 998 367 1010 1633
rect 952 355 1010 367
rect 1410 1633 1468 1645
rect 1410 367 1422 1633
rect 1456 367 1468 1633
rect 1410 355 1468 367
rect 1868 1633 1926 1645
rect 1868 367 1880 1633
rect 1914 367 1926 1633
rect 1868 355 1926 367
rect 2326 1633 2384 1645
rect 2326 367 2338 1633
rect 2372 367 2384 1633
rect 2326 355 2384 367
rect 2784 1633 2842 1645
rect 2784 367 2796 1633
rect 2830 367 2842 1633
rect 2784 355 2842 367
rect 3242 1633 3300 1645
rect 3242 367 3254 1633
rect 3288 367 3300 1633
rect 3242 355 3300 367
rect 3700 1633 3758 1645
rect 3700 367 3712 1633
rect 3746 367 3758 1633
rect 3700 355 3758 367
rect 4158 1633 4216 1645
rect 4158 367 4170 1633
rect 4204 367 4216 1633
rect 4158 355 4216 367
<< pdiffc >>
rect 48 367 82 1633
rect 506 367 540 1633
rect 964 367 998 1633
rect 1422 367 1456 1633
rect 1880 367 1914 1633
rect 2338 367 2372 1633
rect 2796 367 2830 1633
rect 3254 367 3288 1633
rect 3712 367 3746 1633
rect 4170 367 4204 1633
<< poly >>
rect 94 1645 494 1671
rect 552 1645 952 1671
rect 1010 1645 1410 1671
rect 1468 1645 1868 1671
rect 1926 1645 2326 1671
rect 2384 1645 2784 1671
rect 2842 1645 3242 1671
rect 3300 1645 3700 1671
rect 3758 1645 4158 1671
rect 94 329 494 355
rect 552 329 952 355
rect 1010 329 1410 355
rect 1468 329 1868 355
rect 1926 329 2326 355
rect 2384 329 2784 355
rect 2842 329 3242 355
rect 3300 329 3700 355
rect 3758 329 4158 355
rect 240 184 360 329
rect 696 184 816 329
rect 1152 184 1272 329
rect 1608 184 1728 329
rect 2064 184 2184 329
rect 2520 184 2640 329
rect 2976 184 3096 329
rect 3432 184 3552 329
rect 3888 184 4008 329
rect 0 164 4252 184
rect 0 104 170 164
rect 230 104 570 164
rect 630 104 970 164
rect 1030 104 1370 164
rect 1430 104 1770 164
rect 1830 104 2170 164
rect 2230 104 2570 164
rect 2630 104 2970 164
rect 3030 104 3370 164
rect 3430 104 3770 164
rect 3830 104 4252 164
rect 0 84 4252 104
<< polycont >>
rect 170 104 230 164
rect 570 104 630 164
rect 970 104 1030 164
rect 1370 104 1430 164
rect 1770 104 1830 164
rect 2170 104 2230 164
rect 2570 104 2630 164
rect 2970 104 3030 164
rect 3370 104 3430 164
rect 3770 104 3830 164
<< locali >>
rect 0 1850 170 1910
rect 230 1850 570 1910
rect 630 1850 970 1910
rect 1030 1850 1370 1910
rect 1430 1850 1770 1910
rect 1830 1850 2170 1910
rect 2230 1850 2570 1910
rect 2630 1850 2970 1910
rect 3030 1850 3370 1910
rect 3430 1850 3770 1910
rect 3830 1850 4252 1910
rect 0 1730 4252 1790
rect 505 1649 539 1730
rect 1421 1649 1455 1730
rect 2337 1649 2371 1730
rect 3253 1649 3287 1730
rect 4169 1649 4203 1730
rect 48 1633 82 1649
rect 47 367 48 374
rect 505 1633 540 1649
rect 505 1626 506 1633
rect 47 351 82 367
rect 964 1633 998 1649
rect 506 351 540 367
rect 963 367 964 374
rect 1421 1633 1456 1649
rect 1421 1626 1422 1633
rect 963 351 998 367
rect 1880 1633 1914 1649
rect 1422 351 1456 367
rect 1879 367 1880 374
rect 2337 1633 2372 1649
rect 2337 1626 2338 1633
rect 1879 351 1914 367
rect 2796 1633 2830 1649
rect 2338 351 2372 367
rect 2795 367 2796 374
rect 3253 1633 3288 1649
rect 3253 1626 3254 1633
rect 2795 351 2830 367
rect 3712 1633 3746 1649
rect 3254 351 3288 367
rect 3711 367 3712 374
rect 4169 1633 4204 1649
rect 4169 1626 4170 1633
rect 3711 351 3746 367
rect 4170 351 4204 367
rect 47 270 81 351
rect 963 270 997 351
rect 1879 270 1913 351
rect 2795 270 2829 351
rect 3711 270 3745 351
rect 0 210 4252 270
rect 0 104 170 164
rect 230 104 570 164
rect 630 104 970 164
rect 1030 104 1370 164
rect 1430 104 1770 164
rect 1830 104 2170 164
rect 2230 104 2570 164
rect 2630 104 2970 164
rect 3030 104 3370 164
rect 3430 104 3770 164
rect 3830 104 4252 164
rect 0 -30 170 30
rect 230 -30 570 30
rect 630 -30 970 30
rect 1030 -30 1370 30
rect 1430 -30 1770 30
rect 1830 -30 2170 30
rect 2230 -30 2570 30
rect 2630 -30 2970 30
rect 3030 -30 3370 30
rect 3430 -30 3770 30
rect 3830 -30 4252 30
<< viali >>
rect 170 1850 230 1910
rect 570 1850 630 1910
rect 970 1850 1030 1910
rect 1370 1850 1430 1910
rect 1770 1850 1830 1910
rect 2170 1850 2230 1910
rect 2570 1850 2630 1910
rect 2970 1850 3030 1910
rect 3370 1850 3430 1910
rect 3770 1850 3830 1910
rect 48 367 82 1633
rect 506 367 540 1633
rect 964 367 998 1633
rect 1422 367 1456 1633
rect 1880 367 1914 1633
rect 2338 367 2372 1633
rect 2796 367 2830 1633
rect 3254 367 3288 1633
rect 3712 367 3746 1633
rect 4170 367 4204 1633
rect 170 -30 230 30
rect 570 -30 630 30
rect 970 -30 1030 30
rect 1370 -30 1430 30
rect 1770 -30 1830 30
rect 2170 -30 2230 30
rect 2570 -30 2630 30
rect 2970 -30 3030 30
rect 3370 -30 3430 30
rect 3770 -30 3830 30
<< metal1 >>
rect 0 1910 4252 1940
rect 0 1850 170 1910
rect 230 1850 570 1910
rect 630 1850 970 1910
rect 1030 1850 1370 1910
rect 1430 1850 1770 1910
rect 1830 1850 2170 1910
rect 2230 1850 2570 1910
rect 2630 1850 2970 1910
rect 3030 1850 3370 1910
rect 3430 1850 3770 1910
rect 3830 1850 4252 1910
rect 0 1820 4252 1850
rect 42 1633 88 1645
rect 42 367 48 1633
rect 82 367 88 1633
rect 42 355 88 367
rect 500 1633 546 1645
rect 500 367 506 1633
rect 540 367 546 1633
rect 500 355 546 367
rect 958 1633 1004 1645
rect 958 367 964 1633
rect 998 367 1004 1633
rect 958 355 1004 367
rect 1416 1633 1462 1645
rect 1416 367 1422 1633
rect 1456 367 1462 1633
rect 1416 355 1462 367
rect 1874 1633 1920 1645
rect 1874 367 1880 1633
rect 1914 367 1920 1633
rect 1874 355 1920 367
rect 2332 1633 2378 1645
rect 2332 367 2338 1633
rect 2372 367 2378 1633
rect 2332 355 2378 367
rect 2790 1633 2836 1645
rect 2790 367 2796 1633
rect 2830 367 2836 1633
rect 2790 355 2836 367
rect 3248 1633 3294 1645
rect 3248 367 3254 1633
rect 3288 367 3294 1633
rect 3248 355 3294 367
rect 3706 1633 3752 1645
rect 3706 367 3712 1633
rect 3746 367 3752 1633
rect 3706 355 3752 367
rect 4164 1633 4210 1645
rect 4164 367 4170 1633
rect 4204 367 4210 1633
rect 4164 355 4210 367
rect 0 30 4252 60
rect 0 -30 170 30
rect 230 -30 570 30
rect 630 -30 970 30
rect 1030 -30 1370 30
rect 1430 -30 1770 30
rect 1830 -30 2170 30
rect 2230 -30 2570 30
rect 2630 -30 2970 30
rect 3030 -30 3370 30
rect 3430 -30 3770 30
rect 3830 -30 4252 30
rect 0 -60 4252 -30
<< labels >>
flabel nwell 170 1850 230 1910 1 FreeSans 800 0 0 0 VPB
port 4 n power bidirectional
flabel metal1 0 1850 60 1910 1 FreeSans 800 0 0 0 VPWR
port 5 n power bidirectional
flabel metal1 0 -30 60 30 1 FreeSans 800 0 0 0 VGND
port 6 n ground bidirectional
flabel locali 4192 1730 4252 1790 1 FreeSans 800 0 0 0 SOURCE
port 2 n signal bidirectional
flabel locali 4192 210 4252 270 1 FreeSans 800 0 0 0 DRAIN
port 3 n signal bidirectional
flabel locali 4192 104 4252 164 1 FreeSans 800 0 0 0 GATE
port 1 n signal bidirectional
<< properties >>
string FIXED_BBOX 0 0 588 1880
string LEFclass CORE
string LEFsite unitasc
<< end >>
