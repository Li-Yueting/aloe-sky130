../../11-open-magic-def2spice/outputs/design_extracted.spice