../results/ringosc.lef