VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO sky130_asc_pfet_01v8_lvt_6
  CLASS CORE ;
  FOREIGN sky130_asc_pfet_01v8_lvt_6 ;
  ORIGIN 0.000 0.000 ;
  SIZE 14.875 BY 9.400 ;
  SITE unitasc ;
  PIN GATE
    DIRECTION INOUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 77.400002 ;
    PORT
      LAYER li1 ;
        RECT 0.490 0.520 14.870 0.820 ;
    END
  END GATE
  PIN SOURCE
    DIRECTION INOUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 5.611500 ;
    PORT
      LAYER li1 ;
        RECT 0.790 8.650 14.870 8.950 ;
        RECT 3.015 1.755 3.185 8.650 ;
        RECT 7.595 1.755 7.765 8.650 ;
        RECT 12.175 1.755 12.345 8.650 ;
      LAYER mcon ;
        RECT 3.015 1.835 3.185 8.165 ;
        RECT 7.595 1.835 7.765 8.165 ;
        RECT 12.175 1.835 12.345 8.165 ;
      LAYER met1 ;
        RECT 2.985 1.775 3.215 8.225 ;
        RECT 7.565 1.775 7.795 8.225 ;
        RECT 12.145 1.775 12.375 8.225 ;
    END
  END SOURCE
  PIN DRAIN
    DIRECTION INOUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 7.482000 ;
    PORT
      LAYER li1 ;
        RECT 0.725 1.350 0.895 8.245 ;
        RECT 5.305 1.350 5.475 8.245 ;
        RECT 9.885 1.350 10.055 8.245 ;
        RECT 14.465 1.350 14.635 8.245 ;
        RECT 0.490 1.050 14.870 1.350 ;
      LAYER mcon ;
        RECT 0.725 1.835 0.895 8.165 ;
        RECT 5.305 1.835 5.475 8.165 ;
        RECT 9.885 1.835 10.055 8.165 ;
        RECT 14.465 1.835 14.635 8.165 ;
      LAYER met1 ;
        RECT 0.695 1.775 0.925 8.225 ;
        RECT 5.275 1.775 5.505 8.225 ;
        RECT 9.855 1.775 10.085 8.225 ;
        RECT 14.435 1.775 14.665 8.225 ;
    END
  END DRAIN
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT 0.000 8.535 14.870 9.700 ;
        RECT 0.000 1.470 14.875 8.535 ;
        RECT 0.485 1.465 14.875 1.470 ;
      LAYER li1 ;
        RECT 0.000 9.250 14.870 9.550 ;
        RECT 0.140 8.200 0.440 9.250 ;
      LAYER mcon ;
        RECT 1.340 9.250 1.640 9.550 ;
        RECT 3.340 9.250 3.640 9.550 ;
        RECT 5.340 9.250 5.640 9.550 ;
        RECT 7.340 9.250 7.640 9.550 ;
        RECT 9.340 9.250 9.640 9.550 ;
        RECT 11.340 9.250 11.640 9.550 ;
        RECT 13.340 9.250 13.640 9.550 ;
      LAYER met1 ;
        RECT 0.000 9.100 14.870 9.700 ;
    END
  END VPWR
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER li1 ;
        RECT 0.000 -0.150 14.870 0.150 ;
      LAYER mcon ;
        RECT 1.340 -0.150 1.640 0.150 ;
        RECT 3.340 -0.150 3.640 0.150 ;
        RECT 5.340 -0.150 5.640 0.150 ;
        RECT 7.340 -0.150 7.640 0.150 ;
        RECT 9.340 -0.150 9.640 0.150 ;
        RECT 11.340 -0.150 11.640 0.150 ;
        RECT 13.340 -0.150 13.640 0.150 ;
      LAYER met1 ;
        RECT 0.000 -0.300 14.870 0.300 ;
    END
  END VGND
END sky130_asc_pfet_01v8_lvt_6
END LIBRARY

