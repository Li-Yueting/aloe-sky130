VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO sky130_asc_pfet_01v8_lvt_1
  CLASS CORE ;
  FOREIGN sky130_asc_pfet_01v8_lvt_1 ;
  ORIGIN 0.000 0.000 ;
  SIZE 2.940 BY 9.400 ;
  SITE unitasc ;
  PIN GATE
    DIRECTION INOUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 12.900000 ;
    PORT
      LAYER li1 ;
        RECT 0.000 0.520 2.940 0.820 ;
    END
  END GATE
  PIN SOURCE
    DIRECTION INOUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.870500 ;
    PORT
      LAYER li1 ;
        RECT 0.000 8.650 2.940 8.950 ;
        RECT 2.525 8.245 2.695 8.650 ;
        RECT 2.525 8.130 2.700 8.245 ;
        RECT 2.530 1.755 2.700 8.130 ;
      LAYER mcon ;
        RECT 2.530 1.835 2.700 8.165 ;
      LAYER met1 ;
        RECT 2.500 1.775 2.730 8.225 ;
    END
  END SOURCE
  PIN DRAIN
    DIRECTION INOUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.870500 ;
    PORT
      LAYER li1 ;
        RECT 0.240 1.870 0.410 8.245 ;
        RECT 0.235 1.755 0.410 1.870 ;
        RECT 0.235 1.350 0.405 1.755 ;
        RECT 0.000 1.050 2.940 1.350 ;
      LAYER mcon ;
        RECT 0.240 1.835 0.410 8.165 ;
      LAYER met1 ;
        RECT 0.210 1.775 0.440 8.225 ;
    END
  END DRAIN
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT 0.000 1.465 2.940 9.700 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER li1 ;
        RECT 0.000 9.250 2.940 9.550 ;
      LAYER mcon ;
        RECT 0.850 9.250 1.150 9.550 ;
      LAYER met1 ;
        RECT 0.000 9.100 2.940 9.700 ;
    END
  END VPWR
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER li1 ;
        RECT 0.000 -0.150 2.940 0.150 ;
      LAYER mcon ;
        RECT 0.850 -0.150 1.150 0.150 ;
      LAYER met1 ;
        RECT 0.000 -0.300 2.940 0.300 ;
    END
  END VGND
END sky130_asc_pfet_01v8_lvt_1

#--------EOF---------

MACRO sky130_asc_nfet_01v8_lvt_1
  CLASS CORE ;
  FOREIGN sky130_asc_nfet_01v8_lvt_1 ;
  ORIGIN 0.000 0.000 ;
  SIZE 2.580 BY 9.400 ;
  SITE unitasc ;
  PIN VNB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER pwell ;
        RECT 0.000 0.150 2.580 5.000 ;
        RECT 0.150 -0.150 0.450 0.150 ;
    END
  END VNB
  PIN GATE
    DIRECTION INOUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 8.000000 ;
    PORT
      LAYER li1 ;
        RECT 0.000 0.720 2.580 1.020 ;
    END
  END GATE
  PIN SOURCE
    DIRECTION INOUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.160000 ;
    PORT
      LAYER li1 ;
        RECT 0.000 8.250 2.580 8.550 ;
        RECT 2.345 7.020 2.515 8.250 ;
        RECT 2.345 6.730 2.520 7.020 ;
        RECT 2.350 2.980 2.520 6.730 ;
      LAYER mcon ;
        RECT 2.350 3.060 2.520 6.940 ;
      LAYER met1 ;
        RECT 2.320 3.000 2.550 7.000 ;
    END
  END SOURCE
  PIN DRAIN
    DIRECTION INOUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.160000 ;
    PORT
      LAYER li1 ;
        RECT 0.060 3.270 0.230 7.020 ;
        RECT 0.055 2.980 0.230 3.270 ;
        RECT 0.055 2.520 0.225 2.980 ;
        RECT 0.000 2.220 2.580 2.520 ;
      LAYER mcon ;
        RECT 0.060 3.060 0.230 6.940 ;
      LAYER met1 ;
        RECT 0.030 3.000 0.260 7.000 ;
    END
  END DRAIN
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER li1 ;
        RECT 0.000 9.250 2.580 9.550 ;
      LAYER mcon ;
        RECT 0.850 9.250 1.150 9.550 ;
      LAYER met1 ;
        RECT 0.000 9.100 2.580 9.700 ;
    END
  END VPWR
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER li1 ;
        RECT 0.000 -0.150 2.580 0.150 ;
      LAYER mcon ;
        RECT 0.850 -0.150 1.150 0.150 ;
      LAYER met1 ;
        RECT 0.000 -0.300 2.580 0.300 ;
    END
  END VGND
END sky130_asc_nfet_01v8_lvt_1

# -------------EOF--------------------

MACRO sky130_asc_pfet_01v8_lvt_6
  CLASS CORE ;
  FOREIGN sky130_asc_pfet_01v8_lvt_6 ;
  ORIGIN 0.000 0.000 ;
  SIZE 14.395 BY 9.400 ;
  SITE unitasc ;
  PIN GATE
    DIRECTION INOUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 77.400002 ;
    PORT
      LAYER li1 ;
        RECT 0.010 0.520 14.390 0.820 ;
    END
  END GATE
  PIN SOURCE
    DIRECTION INOUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 5.611500 ;
    PORT
      LAYER li1 ;
        RECT 0.010 8.650 14.390 8.950 ;
        RECT 2.535 1.755 2.705 8.650 ;
        RECT 7.115 1.755 7.285 8.650 ;
        RECT 11.695 1.755 11.865 8.650 ;
      LAYER mcon ;
        RECT 2.535 1.835 2.705 8.165 ;
        RECT 7.115 1.835 7.285 8.165 ;
        RECT 11.695 1.835 11.865 8.165 ;
      LAYER met1 ;
        RECT 2.505 1.775 2.735 8.225 ;
        RECT 7.085 1.775 7.315 8.225 ;
        RECT 11.665 1.775 11.895 8.225 ;
    END
  END SOURCE
  PIN DRAIN
    DIRECTION INOUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 7.482000 ;
    PORT
      LAYER li1 ;
        RECT 0.245 1.350 0.415 8.245 ;
        RECT 4.825 1.350 4.995 8.245 ;
        RECT 9.405 1.350 9.575 8.245 ;
        RECT 13.985 1.350 14.155 8.245 ;
        RECT 0.010 1.050 14.390 1.350 ;
      LAYER mcon ;
        RECT 0.245 1.835 0.415 8.165 ;
        RECT 4.825 1.835 4.995 8.165 ;
        RECT 9.405 1.835 9.575 8.165 ;
        RECT 13.985 1.835 14.155 8.165 ;
      LAYER met1 ;
        RECT 0.215 1.775 0.445 8.225 ;
        RECT 4.795 1.775 5.025 8.225 ;
        RECT 9.375 1.775 9.605 8.225 ;
        RECT 13.955 1.775 14.185 8.225 ;
    END
  END DRAIN
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT 0.010 8.535 14.390 9.700 ;
        RECT 0.005 1.465 14.395 8.535 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER li1 ;
        RECT 0.010 9.250 14.390 9.550 ;
      LAYER mcon ;
        RECT 0.860 9.250 1.160 9.550 ;
        RECT 2.860 9.250 3.160 9.550 ;
        RECT 4.860 9.250 5.160 9.550 ;
        RECT 6.860 9.250 7.160 9.550 ;
        RECT 8.860 9.250 9.160 9.550 ;
        RECT 10.860 9.250 11.160 9.550 ;
        RECT 12.860 9.250 13.160 9.550 ;
      LAYER met1 ;
        RECT 0.010 9.100 14.390 9.700 ;
    END
  END VPWR
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER li1 ;
        RECT 0.010 -0.150 14.390 0.150 ;
      LAYER mcon ;
        RECT 0.860 -0.150 1.160 0.150 ;
        RECT 2.860 -0.150 3.160 0.150 ;
        RECT 4.860 -0.150 5.160 0.150 ;
        RECT 6.860 -0.150 7.160 0.150 ;
        RECT 8.860 -0.150 9.160 0.150 ;
        RECT 10.860 -0.150 11.160 0.150 ;
        RECT 12.860 -0.150 13.160 0.150 ;
      LAYER met1 ;
        RECT 0.010 -0.300 14.390 0.300 ;
    END
  END VGND
END sky130_asc_pfet_01v8_lvt_6

# -------------EOF--------------------

MACRO sky130_asc_pfet_01v8_lvt_9
  CLASS CORE ;
  FOREIGN sky130_asc_pfet_01v8_lvt_9 ;
  ORIGIN 0.000 0.000 ;
  SIZE 21.260 BY 9.400 ;
  SITE unitasc ;
  PIN GATE
    DIRECTION INOUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 116.099998 ;
    PORT
      LAYER li1 ;
        RECT 0.000 0.520 21.260 0.820 ;
    END
  END GATE
  PIN SOURCE
    DIRECTION INOUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 9.352500 ;
    PORT
      LAYER li1 ;
        RECT 0.000 8.650 21.260 8.950 ;
        RECT 2.525 8.245 2.695 8.650 ;
        RECT 7.105 8.245 7.275 8.650 ;
        RECT 11.685 8.245 11.855 8.650 ;
        RECT 16.265 8.245 16.435 8.650 ;
        RECT 20.845 8.245 21.015 8.650 ;
        RECT 2.525 8.130 2.700 8.245 ;
        RECT 7.105 8.130 7.280 8.245 ;
        RECT 11.685 8.130 11.860 8.245 ;
        RECT 16.265 8.130 16.440 8.245 ;
        RECT 20.845 8.130 21.020 8.245 ;
        RECT 2.530 1.755 2.700 8.130 ;
        RECT 7.110 1.755 7.280 8.130 ;
        RECT 11.690 1.755 11.860 8.130 ;
        RECT 16.270 1.755 16.440 8.130 ;
        RECT 20.850 1.755 21.020 8.130 ;
      LAYER mcon ;
        RECT 2.530 1.835 2.700 8.165 ;
        RECT 7.110 1.835 7.280 8.165 ;
        RECT 11.690 1.835 11.860 8.165 ;
        RECT 16.270 1.835 16.440 8.165 ;
        RECT 20.850 1.835 21.020 8.165 ;
      LAYER met1 ;
        RECT 2.500 1.775 2.730 8.225 ;
        RECT 7.080 1.775 7.310 8.225 ;
        RECT 11.660 1.775 11.890 8.225 ;
        RECT 16.240 1.775 16.470 8.225 ;
        RECT 20.820 1.775 21.050 8.225 ;
    END
  END SOURCE
  PIN DRAIN
    DIRECTION INOUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 9.352500 ;
    PORT
      LAYER li1 ;
        RECT 0.240 1.870 0.410 8.245 ;
        RECT 4.820 1.870 4.990 8.245 ;
        RECT 9.400 1.870 9.570 8.245 ;
        RECT 13.980 1.870 14.150 8.245 ;
        RECT 18.560 1.870 18.730 8.245 ;
        RECT 0.235 1.755 0.410 1.870 ;
        RECT 4.815 1.755 4.990 1.870 ;
        RECT 9.395 1.755 9.570 1.870 ;
        RECT 13.975 1.755 14.150 1.870 ;
        RECT 18.555 1.755 18.730 1.870 ;
        RECT 0.235 1.350 0.405 1.755 ;
        RECT 4.815 1.350 4.985 1.755 ;
        RECT 9.395 1.350 9.565 1.755 ;
        RECT 13.975 1.350 14.145 1.755 ;
        RECT 18.555 1.350 18.725 1.755 ;
        RECT 0.000 1.050 21.260 1.350 ;
      LAYER mcon ;
        RECT 0.240 1.835 0.410 8.165 ;
        RECT 4.820 1.835 4.990 8.165 ;
        RECT 9.400 1.835 9.570 8.165 ;
        RECT 13.980 1.835 14.150 8.165 ;
        RECT 18.560 1.835 18.730 8.165 ;
      LAYER met1 ;
        RECT 0.210 1.775 0.440 8.225 ;
        RECT 4.790 1.775 5.020 8.225 ;
        RECT 9.370 1.775 9.600 8.225 ;
        RECT 13.950 1.775 14.180 8.225 ;
        RECT 18.530 1.775 18.760 8.225 ;
    END
  END DRAIN
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT 0.000 1.465 21.260 9.700 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER li1 ;
        RECT 0.000 9.250 21.260 9.550 ;
      LAYER mcon ;
        RECT 0.850 9.250 1.150 9.550 ;
        RECT 2.850 9.250 3.150 9.550 ;
        RECT 4.850 9.250 5.150 9.550 ;
        RECT 6.850 9.250 7.150 9.550 ;
        RECT 8.850 9.250 9.150 9.550 ;
        RECT 10.850 9.250 11.150 9.550 ;
        RECT 12.850 9.250 13.150 9.550 ;
        RECT 14.850 9.250 15.150 9.550 ;
        RECT 16.850 9.250 17.150 9.550 ;
        RECT 18.850 9.250 19.150 9.550 ;
      LAYER met1 ;
        RECT 0.000 9.100 21.260 9.700 ;
    END
  END VPWR
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER li1 ;
        RECT 0.000 -0.150 21.260 0.150 ;
      LAYER mcon ;
        RECT 0.850 -0.150 1.150 0.150 ;
        RECT 2.850 -0.150 3.150 0.150 ;
        RECT 4.850 -0.150 5.150 0.150 ;
        RECT 6.850 -0.150 7.150 0.150 ;
        RECT 8.850 -0.150 9.150 0.150 ;
        RECT 10.850 -0.150 11.150 0.150 ;
        RECT 12.850 -0.150 13.150 0.150 ;
        RECT 14.850 -0.150 15.150 0.150 ;
        RECT 16.850 -0.150 17.150 0.150 ;
        RECT 18.850 -0.150 19.150 0.150 ;
      LAYER met1 ;
        RECT 0.000 -0.300 21.260 0.300 ;
    END
  END VGND
END sky130_asc_pfet_01v8_lvt_9

# -------------EOF--------------------

MACRO sky130_asc_pfet_01v8_lvt_12
  CLASS CORE ;
  FOREIGN sky130_asc_pfet_01v8_lvt_12 ;
  ORIGIN 0.000 0.000 ;
  SIZE 28.135 BY 9.400 ;
  SITE unitasc ;
  PIN GATE
    DIRECTION INOUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 154.800003 ;
    PORT
      LAYER li1 ;
        RECT 0.010 0.520 28.130 0.820 ;
    END
  END GATE
  PIN SOURCE
    DIRECTION INOUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 11.223000 ;
    PORT
      LAYER li1 ;
        RECT 0.010 8.650 28.130 8.950 ;
        RECT 2.535 1.755 2.705 8.650 ;
        RECT 7.115 1.755 7.285 8.650 ;
        RECT 11.695 1.755 11.865 8.650 ;
        RECT 16.275 1.755 16.445 8.650 ;
        RECT 20.855 1.755 21.025 8.650 ;
        RECT 25.435 1.755 25.605 8.650 ;
      LAYER mcon ;
        RECT 2.535 1.835 2.705 8.165 ;
        RECT 7.115 1.835 7.285 8.165 ;
        RECT 11.695 1.835 11.865 8.165 ;
        RECT 16.275 1.835 16.445 8.165 ;
        RECT 20.855 1.835 21.025 8.165 ;
        RECT 25.435 1.835 25.605 8.165 ;
      LAYER met1 ;
        RECT 2.505 1.775 2.735 8.225 ;
        RECT 7.085 1.775 7.315 8.225 ;
        RECT 11.665 1.775 11.895 8.225 ;
        RECT 16.245 1.775 16.475 8.225 ;
        RECT 20.825 1.775 21.055 8.225 ;
        RECT 25.405 1.775 25.635 8.225 ;
    END
  END SOURCE
  PIN DRAIN
    DIRECTION INOUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 13.093500 ;
    PORT
      LAYER li1 ;
        RECT 0.245 1.350 0.415 8.245 ;
        RECT 4.825 1.350 4.995 8.245 ;
        RECT 9.405 1.350 9.575 8.245 ;
        RECT 13.985 1.350 14.155 8.245 ;
        RECT 18.565 1.350 18.735 8.245 ;
        RECT 23.145 1.350 23.315 8.245 ;
        RECT 27.725 1.350 27.895 8.245 ;
        RECT 0.010 1.050 28.130 1.350 ;
      LAYER mcon ;
        RECT 0.245 1.835 0.415 8.165 ;
        RECT 4.825 1.835 4.995 8.165 ;
        RECT 9.405 1.835 9.575 8.165 ;
        RECT 13.985 1.835 14.155 8.165 ;
        RECT 18.565 1.835 18.735 8.165 ;
        RECT 23.145 1.835 23.315 8.165 ;
        RECT 27.725 1.835 27.895 8.165 ;
      LAYER met1 ;
        RECT 0.215 1.775 0.445 8.225 ;
        RECT 4.795 1.775 5.025 8.225 ;
        RECT 9.375 1.775 9.605 8.225 ;
        RECT 13.955 1.775 14.185 8.225 ;
        RECT 18.535 1.775 18.765 8.225 ;
        RECT 23.115 1.775 23.345 8.225 ;
        RECT 27.695 1.775 27.925 8.225 ;
    END
  END DRAIN
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT 0.010 8.535 28.130 9.700 ;
        RECT 0.005 1.465 28.135 8.535 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER li1 ;
        RECT 0.010 9.250 28.130 9.550 ;
      LAYER mcon ;
        RECT 0.860 9.250 1.160 9.550 ;
        RECT 2.860 9.250 3.160 9.550 ;
        RECT 4.860 9.250 5.160 9.550 ;
        RECT 6.860 9.250 7.160 9.550 ;
        RECT 8.860 9.250 9.160 9.550 ;
        RECT 10.860 9.250 11.160 9.550 ;
        RECT 12.860 9.250 13.160 9.550 ;
        RECT 14.860 9.250 15.160 9.550 ;
        RECT 16.860 9.250 17.160 9.550 ;
        RECT 18.860 9.250 19.160 9.550 ;
        RECT 20.860 9.250 21.160 9.550 ;
        RECT 22.860 9.250 23.160 9.550 ;
        RECT 24.860 9.250 25.160 9.550 ;
        RECT 26.860 9.250 27.160 9.550 ;
      LAYER met1 ;
        RECT 0.010 9.100 28.130 9.700 ;
    END
  END VPWR
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER li1 ;
        RECT 0.010 -0.150 28.130 0.150 ;
      LAYER mcon ;
        RECT 0.860 -0.150 1.160 0.150 ;
        RECT 2.860 -0.150 3.160 0.150 ;
        RECT 4.860 -0.150 5.160 0.150 ;
        RECT 6.860 -0.150 7.160 0.150 ;
        RECT 8.860 -0.150 9.160 0.150 ;
        RECT 10.860 -0.150 11.160 0.150 ;
        RECT 12.860 -0.150 13.160 0.150 ;
        RECT 14.860 -0.150 15.160 0.150 ;
        RECT 16.860 -0.150 17.160 0.150 ;
        RECT 18.860 -0.150 19.160 0.150 ;
        RECT 20.860 -0.150 21.160 0.150 ;
        RECT 22.860 -0.150 23.160 0.150 ;
        RECT 24.860 -0.150 25.160 0.150 ;
        RECT 26.860 -0.150 27.160 0.150 ;
      LAYER met1 ;
        RECT 0.010 -0.300 28.130 0.300 ;
    END
  END VGND
END sky130_asc_pfet_01v8_lvt_12

# -------------EOF--------------------

MACRO sky130_asc_pfet_01v8_lvt_60
  CLASS CORE ;
  FOREIGN sky130_asc_pfet_01v8_lvt_60 ;
  ORIGIN 0.000 0.000 ;
  SIZE 138.055 BY 9.400 ;
  SITE unitasc ;
  PIN GATE
    DIRECTION INOUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 774.000000 ;
    PORT
      LAYER li1 ;
        RECT 0.010 0.520 138.050 0.820 ;
    END
  END GATE
  PIN SOURCE
    DIRECTION INOUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 56.114998 ;
    PORT
      LAYER li1 ;
        RECT 0.010 8.650 138.050 8.950 ;
        RECT 2.535 1.755 2.705 8.650 ;
        RECT 7.115 1.755 7.285 8.650 ;
        RECT 11.695 1.755 11.865 8.650 ;
        RECT 16.275 1.755 16.445 8.650 ;
        RECT 20.855 1.755 21.025 8.650 ;
        RECT 25.435 1.755 25.605 8.650 ;
        RECT 30.015 1.755 30.185 8.650 ;
        RECT 34.595 1.755 34.765 8.650 ;
        RECT 39.175 1.755 39.345 8.650 ;
        RECT 43.755 1.755 43.925 8.650 ;
        RECT 48.335 1.755 48.505 8.650 ;
        RECT 52.915 1.755 53.085 8.650 ;
        RECT 57.495 1.755 57.665 8.650 ;
        RECT 62.075 1.755 62.245 8.650 ;
        RECT 66.655 1.755 66.825 8.650 ;
        RECT 71.235 1.755 71.405 8.650 ;
        RECT 75.815 1.755 75.985 8.650 ;
        RECT 80.395 1.755 80.565 8.650 ;
        RECT 84.975 1.755 85.145 8.650 ;
        RECT 89.555 1.755 89.725 8.650 ;
        RECT 94.135 1.755 94.305 8.650 ;
        RECT 98.715 1.755 98.885 8.650 ;
        RECT 103.295 1.755 103.465 8.650 ;
        RECT 107.875 1.755 108.045 8.650 ;
        RECT 112.455 1.755 112.625 8.650 ;
        RECT 117.035 1.755 117.205 8.650 ;
        RECT 121.615 1.755 121.785 8.650 ;
        RECT 126.195 1.755 126.365 8.650 ;
        RECT 130.775 1.755 130.945 8.650 ;
        RECT 135.355 1.755 135.525 8.650 ;
      LAYER mcon ;
        RECT 2.535 1.835 2.705 8.165 ;
        RECT 7.115 1.835 7.285 8.165 ;
        RECT 11.695 1.835 11.865 8.165 ;
        RECT 16.275 1.835 16.445 8.165 ;
        RECT 20.855 1.835 21.025 8.165 ;
        RECT 25.435 1.835 25.605 8.165 ;
        RECT 30.015 1.835 30.185 8.165 ;
        RECT 34.595 1.835 34.765 8.165 ;
        RECT 39.175 1.835 39.345 8.165 ;
        RECT 43.755 1.835 43.925 8.165 ;
        RECT 48.335 1.835 48.505 8.165 ;
        RECT 52.915 1.835 53.085 8.165 ;
        RECT 57.495 1.835 57.665 8.165 ;
        RECT 62.075 1.835 62.245 8.165 ;
        RECT 66.655 1.835 66.825 8.165 ;
        RECT 71.235 1.835 71.405 8.165 ;
        RECT 75.815 1.835 75.985 8.165 ;
        RECT 80.395 1.835 80.565 8.165 ;
        RECT 84.975 1.835 85.145 8.165 ;
        RECT 89.555 1.835 89.725 8.165 ;
        RECT 94.135 1.835 94.305 8.165 ;
        RECT 98.715 1.835 98.885 8.165 ;
        RECT 103.295 1.835 103.465 8.165 ;
        RECT 107.875 1.835 108.045 8.165 ;
        RECT 112.455 1.835 112.625 8.165 ;
        RECT 117.035 1.835 117.205 8.165 ;
        RECT 121.615 1.835 121.785 8.165 ;
        RECT 126.195 1.835 126.365 8.165 ;
        RECT 130.775 1.835 130.945 8.165 ;
        RECT 135.355 1.835 135.525 8.165 ;
      LAYER met1 ;
        RECT 2.505 1.775 2.735 8.225 ;
        RECT 7.085 1.775 7.315 8.225 ;
        RECT 11.665 1.775 11.895 8.225 ;
        RECT 16.245 1.775 16.475 8.225 ;
        RECT 20.825 1.775 21.055 8.225 ;
        RECT 25.405 1.775 25.635 8.225 ;
        RECT 29.985 1.775 30.215 8.225 ;
        RECT 34.565 1.775 34.795 8.225 ;
        RECT 39.145 1.775 39.375 8.225 ;
        RECT 43.725 1.775 43.955 8.225 ;
        RECT 48.305 1.775 48.535 8.225 ;
        RECT 52.885 1.775 53.115 8.225 ;
        RECT 57.465 1.775 57.695 8.225 ;
        RECT 62.045 1.775 62.275 8.225 ;
        RECT 66.625 1.775 66.855 8.225 ;
        RECT 71.205 1.775 71.435 8.225 ;
        RECT 75.785 1.775 76.015 8.225 ;
        RECT 80.365 1.775 80.595 8.225 ;
        RECT 84.945 1.775 85.175 8.225 ;
        RECT 89.525 1.775 89.755 8.225 ;
        RECT 94.105 1.775 94.335 8.225 ;
        RECT 98.685 1.775 98.915 8.225 ;
        RECT 103.265 1.775 103.495 8.225 ;
        RECT 107.845 1.775 108.075 8.225 ;
        RECT 112.425 1.775 112.655 8.225 ;
        RECT 117.005 1.775 117.235 8.225 ;
        RECT 121.585 1.775 121.815 8.225 ;
        RECT 126.165 1.775 126.395 8.225 ;
        RECT 130.745 1.775 130.975 8.225 ;
        RECT 135.325 1.775 135.555 8.225 ;
    END
  END SOURCE
  PIN DRAIN
    DIRECTION INOUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 57.985500 ;
    PORT
      LAYER li1 ;
        RECT 0.245 1.350 0.415 8.245 ;
        RECT 4.825 1.350 4.995 8.245 ;
        RECT 9.405 1.350 9.575 8.245 ;
        RECT 13.985 1.350 14.155 8.245 ;
        RECT 18.565 1.350 18.735 8.245 ;
        RECT 23.145 1.350 23.315 8.245 ;
        RECT 27.725 1.350 27.895 8.245 ;
        RECT 32.305 1.350 32.475 8.245 ;
        RECT 36.885 1.350 37.055 8.245 ;
        RECT 41.465 1.350 41.635 8.245 ;
        RECT 46.045 1.350 46.215 8.245 ;
        RECT 50.625 1.350 50.795 8.245 ;
        RECT 55.205 1.350 55.375 8.245 ;
        RECT 59.785 1.350 59.955 8.245 ;
        RECT 64.365 1.350 64.535 8.245 ;
        RECT 68.945 1.350 69.115 8.245 ;
        RECT 73.525 1.350 73.695 8.245 ;
        RECT 78.105 1.350 78.275 8.245 ;
        RECT 82.685 1.350 82.855 8.245 ;
        RECT 87.265 1.350 87.435 8.245 ;
        RECT 91.845 1.350 92.015 8.245 ;
        RECT 96.425 1.350 96.595 8.245 ;
        RECT 101.005 1.350 101.175 8.245 ;
        RECT 105.585 1.350 105.755 8.245 ;
        RECT 110.165 1.350 110.335 8.245 ;
        RECT 114.745 1.350 114.915 8.245 ;
        RECT 119.325 1.350 119.495 8.245 ;
        RECT 123.905 1.350 124.075 8.245 ;
        RECT 128.485 1.350 128.655 8.245 ;
        RECT 133.065 1.350 133.235 8.245 ;
        RECT 137.645 1.350 137.815 8.245 ;
        RECT 0.010 1.050 138.050 1.350 ;
      LAYER mcon ;
        RECT 0.245 1.835 0.415 8.165 ;
        RECT 4.825 1.835 4.995 8.165 ;
        RECT 9.405 1.835 9.575 8.165 ;
        RECT 13.985 1.835 14.155 8.165 ;
        RECT 18.565 1.835 18.735 8.165 ;
        RECT 23.145 1.835 23.315 8.165 ;
        RECT 27.725 1.835 27.895 8.165 ;
        RECT 32.305 1.835 32.475 8.165 ;
        RECT 36.885 1.835 37.055 8.165 ;
        RECT 41.465 1.835 41.635 8.165 ;
        RECT 46.045 1.835 46.215 8.165 ;
        RECT 50.625 1.835 50.795 8.165 ;
        RECT 55.205 1.835 55.375 8.165 ;
        RECT 59.785 1.835 59.955 8.165 ;
        RECT 64.365 1.835 64.535 8.165 ;
        RECT 68.945 1.835 69.115 8.165 ;
        RECT 73.525 1.835 73.695 8.165 ;
        RECT 78.105 1.835 78.275 8.165 ;
        RECT 82.685 1.835 82.855 8.165 ;
        RECT 87.265 1.835 87.435 8.165 ;
        RECT 91.845 1.835 92.015 8.165 ;
        RECT 96.425 1.835 96.595 8.165 ;
        RECT 101.005 1.835 101.175 8.165 ;
        RECT 105.585 1.835 105.755 8.165 ;
        RECT 110.165 1.835 110.335 8.165 ;
        RECT 114.745 1.835 114.915 8.165 ;
        RECT 119.325 1.835 119.495 8.165 ;
        RECT 123.905 1.835 124.075 8.165 ;
        RECT 128.485 1.835 128.655 8.165 ;
        RECT 133.065 1.835 133.235 8.165 ;
        RECT 137.645 1.835 137.815 8.165 ;
      LAYER met1 ;
        RECT 0.215 1.775 0.445 8.225 ;
        RECT 4.795 1.775 5.025 8.225 ;
        RECT 9.375 1.775 9.605 8.225 ;
        RECT 13.955 1.775 14.185 8.225 ;
        RECT 18.535 1.775 18.765 8.225 ;
        RECT 23.115 1.775 23.345 8.225 ;
        RECT 27.695 1.775 27.925 8.225 ;
        RECT 32.275 1.775 32.505 8.225 ;
        RECT 36.855 1.775 37.085 8.225 ;
        RECT 41.435 1.775 41.665 8.225 ;
        RECT 46.015 1.775 46.245 8.225 ;
        RECT 50.595 1.775 50.825 8.225 ;
        RECT 55.175 1.775 55.405 8.225 ;
        RECT 59.755 1.775 59.985 8.225 ;
        RECT 64.335 1.775 64.565 8.225 ;
        RECT 68.915 1.775 69.145 8.225 ;
        RECT 73.495 1.775 73.725 8.225 ;
        RECT 78.075 1.775 78.305 8.225 ;
        RECT 82.655 1.775 82.885 8.225 ;
        RECT 87.235 1.775 87.465 8.225 ;
        RECT 91.815 1.775 92.045 8.225 ;
        RECT 96.395 1.775 96.625 8.225 ;
        RECT 100.975 1.775 101.205 8.225 ;
        RECT 105.555 1.775 105.785 8.225 ;
        RECT 110.135 1.775 110.365 8.225 ;
        RECT 114.715 1.775 114.945 8.225 ;
        RECT 119.295 1.775 119.525 8.225 ;
        RECT 123.875 1.775 124.105 8.225 ;
        RECT 128.455 1.775 128.685 8.225 ;
        RECT 133.035 1.775 133.265 8.225 ;
        RECT 137.615 1.775 137.845 8.225 ;
    END
  END DRAIN
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT 0.010 8.535 138.050 9.700 ;
        RECT 0.005 1.465 138.055 8.535 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER li1 ;
        RECT 0.010 9.250 138.050 9.550 ;
      LAYER mcon ;
        RECT 0.860 9.250 1.160 9.550 ;
        RECT 2.860 9.250 3.160 9.550 ;
        RECT 4.860 9.250 5.160 9.550 ;
        RECT 6.860 9.250 7.160 9.550 ;
        RECT 8.860 9.250 9.160 9.550 ;
        RECT 10.860 9.250 11.160 9.550 ;
        RECT 12.860 9.250 13.160 9.550 ;
        RECT 14.860 9.250 15.160 9.550 ;
        RECT 16.860 9.250 17.160 9.550 ;
        RECT 18.860 9.250 19.160 9.550 ;
        RECT 20.860 9.250 21.160 9.550 ;
        RECT 22.860 9.250 23.160 9.550 ;
        RECT 24.860 9.250 25.160 9.550 ;
        RECT 26.860 9.250 27.160 9.550 ;
        RECT 28.860 9.250 29.160 9.550 ;
        RECT 30.860 9.250 31.160 9.550 ;
        RECT 32.860 9.250 33.160 9.550 ;
        RECT 34.860 9.250 35.160 9.550 ;
        RECT 36.860 9.250 37.160 9.550 ;
        RECT 38.860 9.250 39.160 9.550 ;
        RECT 40.860 9.250 41.160 9.550 ;
        RECT 42.860 9.250 43.160 9.550 ;
        RECT 44.860 9.250 45.160 9.550 ;
        RECT 46.860 9.250 47.160 9.550 ;
        RECT 48.860 9.250 49.160 9.550 ;
        RECT 50.860 9.250 51.160 9.550 ;
        RECT 52.860 9.250 53.160 9.550 ;
        RECT 54.860 9.250 55.160 9.550 ;
        RECT 56.860 9.250 57.160 9.550 ;
        RECT 58.860 9.250 59.160 9.550 ;
        RECT 60.860 9.250 61.160 9.550 ;
        RECT 62.860 9.250 63.160 9.550 ;
        RECT 64.860 9.250 65.160 9.550 ;
        RECT 66.860 9.250 67.160 9.550 ;
        RECT 68.860 9.250 69.160 9.550 ;
        RECT 70.860 9.250 71.160 9.550 ;
        RECT 72.860 9.250 73.160 9.550 ;
        RECT 74.860 9.250 75.160 9.550 ;
        RECT 76.860 9.250 77.160 9.550 ;
        RECT 78.860 9.250 79.160 9.550 ;
        RECT 80.860 9.250 81.160 9.550 ;
        RECT 82.860 9.250 83.160 9.550 ;
        RECT 84.860 9.250 85.160 9.550 ;
        RECT 86.860 9.250 87.160 9.550 ;
        RECT 88.860 9.250 89.160 9.550 ;
        RECT 90.860 9.250 91.160 9.550 ;
        RECT 92.860 9.250 93.160 9.550 ;
        RECT 94.860 9.250 95.160 9.550 ;
        RECT 96.860 9.250 97.160 9.550 ;
        RECT 98.860 9.250 99.160 9.550 ;
        RECT 100.860 9.250 101.160 9.550 ;
        RECT 102.860 9.250 103.160 9.550 ;
        RECT 104.860 9.250 105.160 9.550 ;
        RECT 106.860 9.250 107.160 9.550 ;
        RECT 108.860 9.250 109.160 9.550 ;
        RECT 110.860 9.250 111.160 9.550 ;
        RECT 112.860 9.250 113.160 9.550 ;
        RECT 114.860 9.250 115.160 9.550 ;
        RECT 116.860 9.250 117.160 9.550 ;
        RECT 118.860 9.250 119.160 9.550 ;
        RECT 120.860 9.250 121.160 9.550 ;
        RECT 122.860 9.250 123.160 9.550 ;
        RECT 124.860 9.250 125.160 9.550 ;
        RECT 126.860 9.250 127.160 9.550 ;
        RECT 128.860 9.250 129.160 9.550 ;
        RECT 130.860 9.250 131.160 9.550 ;
        RECT 132.860 9.250 133.160 9.550 ;
        RECT 134.860 9.250 135.160 9.550 ;
        RECT 136.860 9.250 137.160 9.550 ;
      LAYER met1 ;
        RECT 0.010 9.100 138.050 9.700 ;
    END
  END VPWR
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER li1 ;
        RECT 0.010 -0.150 138.050 0.150 ;
      LAYER mcon ;
        RECT 0.860 -0.150 1.160 0.150 ;
        RECT 2.860 -0.150 3.160 0.150 ;
        RECT 4.860 -0.150 5.160 0.150 ;
        RECT 6.860 -0.150 7.160 0.150 ;
        RECT 8.860 -0.150 9.160 0.150 ;
        RECT 10.860 -0.150 11.160 0.150 ;
        RECT 12.860 -0.150 13.160 0.150 ;
        RECT 14.860 -0.150 15.160 0.150 ;
        RECT 16.860 -0.150 17.160 0.150 ;
        RECT 18.860 -0.150 19.160 0.150 ;
        RECT 20.860 -0.150 21.160 0.150 ;
        RECT 22.860 -0.150 23.160 0.150 ;
        RECT 24.860 -0.150 25.160 0.150 ;
        RECT 26.860 -0.150 27.160 0.150 ;
        RECT 28.860 -0.150 29.160 0.150 ;
        RECT 30.860 -0.150 31.160 0.150 ;
        RECT 32.860 -0.150 33.160 0.150 ;
        RECT 34.860 -0.150 35.160 0.150 ;
        RECT 36.860 -0.150 37.160 0.150 ;
        RECT 38.860 -0.150 39.160 0.150 ;
        RECT 40.860 -0.150 41.160 0.150 ;
        RECT 42.860 -0.150 43.160 0.150 ;
        RECT 44.860 -0.150 45.160 0.150 ;
        RECT 46.860 -0.150 47.160 0.150 ;
        RECT 48.860 -0.150 49.160 0.150 ;
        RECT 50.860 -0.150 51.160 0.150 ;
        RECT 52.860 -0.150 53.160 0.150 ;
        RECT 54.860 -0.150 55.160 0.150 ;
        RECT 56.860 -0.150 57.160 0.150 ;
        RECT 58.860 -0.150 59.160 0.150 ;
        RECT 60.860 -0.150 61.160 0.150 ;
        RECT 62.860 -0.150 63.160 0.150 ;
        RECT 64.860 -0.150 65.160 0.150 ;
        RECT 66.860 -0.150 67.160 0.150 ;
        RECT 68.860 -0.150 69.160 0.150 ;
        RECT 70.860 -0.150 71.160 0.150 ;
        RECT 72.860 -0.150 73.160 0.150 ;
        RECT 74.860 -0.150 75.160 0.150 ;
        RECT 76.860 -0.150 77.160 0.150 ;
        RECT 78.860 -0.150 79.160 0.150 ;
        RECT 80.860 -0.150 81.160 0.150 ;
        RECT 82.860 -0.150 83.160 0.150 ;
        RECT 84.860 -0.150 85.160 0.150 ;
        RECT 86.860 -0.150 87.160 0.150 ;
        RECT 88.860 -0.150 89.160 0.150 ;
        RECT 90.860 -0.150 91.160 0.150 ;
        RECT 92.860 -0.150 93.160 0.150 ;
        RECT 94.860 -0.150 95.160 0.150 ;
        RECT 96.860 -0.150 97.160 0.150 ;
        RECT 98.860 -0.150 99.160 0.150 ;
        RECT 100.860 -0.150 101.160 0.150 ;
        RECT 102.860 -0.150 103.160 0.150 ;
        RECT 104.860 -0.150 105.160 0.150 ;
        RECT 106.860 -0.150 107.160 0.150 ;
        RECT 108.860 -0.150 109.160 0.150 ;
        RECT 110.860 -0.150 111.160 0.150 ;
        RECT 112.860 -0.150 113.160 0.150 ;
        RECT 114.860 -0.150 115.160 0.150 ;
        RECT 116.860 -0.150 117.160 0.150 ;
        RECT 118.860 -0.150 119.160 0.150 ;
        RECT 120.860 -0.150 121.160 0.150 ;
        RECT 122.860 -0.150 123.160 0.150 ;
        RECT 124.860 -0.150 125.160 0.150 ;
        RECT 126.860 -0.150 127.160 0.150 ;
        RECT 128.860 -0.150 129.160 0.150 ;
        RECT 130.860 -0.150 131.160 0.150 ;
        RECT 132.860 -0.150 133.160 0.150 ;
        RECT 134.860 -0.150 135.160 0.150 ;
        RECT 136.860 -0.150 137.160 0.150 ;
      LAYER met1 ;
        RECT 0.010 -0.300 138.050 0.300 ;
    END
  END VGND
END sky130_asc_pfet_01v8_lvt_60

# -------------EOF--------------------

MACRO sky130_asc_nfet_01v8_lvt_9
  CLASS CORE ;
  FOREIGN sky130_asc_nfet_01v8_lvt_9 ;
  ORIGIN 0.000 0.000 ;
  SIZE 20.900 BY 9.400 ;
  SITE unitasc ;
  PIN GATE
    DIRECTION INOUT ;
    ANTENNAGATEAREA 54.000000 ;
    PORT
      LAYER li1 ;
        RECT 0.000 1.220 20.900 1.520 ;
    END
  END GATE
  PIN SOURCE
    DIRECTION INOUT ;
    ANTENNADIFFAREA 4.350000 ;
    PORT
      LAYER li1 ;
        RECT 0.000 8.450 20.900 8.750 ;
        RECT 2.345 6.520 2.515 8.450 ;
        RECT 6.925 6.520 7.095 8.450 ;
        RECT 11.505 6.520 11.675 8.450 ;
        RECT 16.085 6.520 16.255 8.450 ;
        RECT 20.665 6.520 20.835 8.450 ;
        RECT 2.345 6.430 2.520 6.520 ;
        RECT 6.925 6.430 7.100 6.520 ;
        RECT 11.505 6.430 11.680 6.520 ;
        RECT 16.085 6.430 16.260 6.520 ;
        RECT 20.665 6.430 20.840 6.520 ;
        RECT 2.350 3.480 2.520 6.430 ;
        RECT 6.930 3.480 7.100 6.430 ;
        RECT 11.510 3.480 11.680 6.430 ;
        RECT 16.090 3.480 16.260 6.430 ;
        RECT 20.670 3.480 20.840 6.430 ;
      LAYER mcon ;
        RECT 2.350 3.560 2.520 6.440 ;
        RECT 6.930 3.560 7.100 6.440 ;
        RECT 11.510 3.560 11.680 6.440 ;
        RECT 16.090 3.560 16.260 6.440 ;
        RECT 20.670 3.560 20.840 6.440 ;
      LAYER met1 ;
        RECT 2.320 3.500 2.550 6.500 ;
        RECT 6.900 3.500 7.130 6.500 ;
        RECT 11.480 3.500 11.710 6.500 ;
        RECT 16.060 3.500 16.290 6.500 ;
        RECT 20.640 3.500 20.870 6.500 ;
    END
  END SOURCE
  PIN DRAIN
    DIRECTION INOUT ;
    ANTENNADIFFAREA 4.350000 ;
    PORT
      LAYER li1 ;
        RECT 0.060 3.770 0.230 6.520 ;
        RECT 4.640 3.770 4.810 6.520 ;
        RECT 9.220 3.770 9.390 6.520 ;
        RECT 13.800 3.770 13.970 6.520 ;
        RECT 18.380 3.770 18.550 6.520 ;
        RECT 0.055 3.480 0.230 3.770 ;
        RECT 4.635 3.480 4.810 3.770 ;
        RECT 9.215 3.480 9.390 3.770 ;
        RECT 13.795 3.480 13.970 3.770 ;
        RECT 18.375 3.480 18.550 3.770 ;
        RECT 0.055 2.150 0.225 3.480 ;
        RECT 4.635 2.150 4.805 3.480 ;
        RECT 9.215 2.150 9.385 3.480 ;
        RECT 13.795 2.150 13.965 3.480 ;
        RECT 18.375 2.150 18.545 3.480 ;
        RECT 0.000 1.850 20.900 2.150 ;
      LAYER mcon ;
        RECT 0.060 3.560 0.230 6.440 ;
        RECT 4.640 3.560 4.810 6.440 ;
        RECT 9.220 3.560 9.390 6.440 ;
        RECT 13.800 3.560 13.970 6.440 ;
        RECT 18.380 3.560 18.550 6.440 ;
      LAYER met1 ;
        RECT 0.030 3.500 0.260 6.500 ;
        RECT 4.610 3.500 4.840 6.500 ;
        RECT 9.190 3.500 9.420 6.500 ;
        RECT 13.770 3.500 14.000 6.500 ;
        RECT 18.350 3.500 18.580 6.500 ;
    END
  END DRAIN
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.000 0.150 20.900 5.000 ;
        RECT 20.600 -0.150 20.900 0.150 ;
    END
  END VNB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER li1 ;
        RECT 0.000 9.250 20.900 9.550 ;
      LAYER mcon ;
        RECT 0.850 9.250 1.150 9.550 ;
        RECT 2.850 9.250 3.150 9.550 ;
        RECT 4.850 9.250 5.150 9.550 ;
        RECT 6.850 9.250 7.150 9.550 ;
        RECT 8.850 9.250 9.150 9.550 ;
        RECT 10.850 9.250 11.150 9.550 ;
        RECT 12.850 9.250 13.150 9.550 ;
        RECT 14.850 9.250 15.150 9.550 ;
        RECT 16.850 9.250 17.150 9.550 ;
        RECT 18.850 9.250 19.150 9.550 ;
      LAYER met1 ;
        RECT 0.000 9.100 20.900 9.700 ;
    END
  END VPWR
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER li1 ;
        RECT 0.000 -0.150 20.900 0.150 ;
      LAYER mcon ;
        RECT 0.850 -0.150 1.150 0.150 ;
        RECT 2.850 -0.150 3.150 0.150 ;
        RECT 4.850 -0.150 5.150 0.150 ;
        RECT 6.850 -0.150 7.150 0.150 ;
        RECT 8.850 -0.150 9.150 0.150 ;
        RECT 10.850 -0.150 11.150 0.150 ;
        RECT 12.850 -0.150 13.150 0.150 ;
        RECT 14.850 -0.150 15.150 0.150 ;
        RECT 16.850 -0.150 17.150 0.150 ;
        RECT 18.850 -0.150 19.150 0.150 ;
      LAYER met1 ;
        RECT 0.000 -0.300 20.900 0.300 ;
    END
  END VGND
END sky130_asc_nfet_01v8_lvt_9

# -------------EOF--------------------

MACRO sky130_asc_res
  CLASS CORE ;
  FOREIGN sky130_asc_res ;
  ORIGIN 0.000 0.000 ;
  SIZE 12.200 BY 9.400 ;
  SITE unitasc ;
  PIN Rin
    DIRECTION INOUT ;
    PORT
      LAYER li1 ;
        RECT 0.000 5.375 2.160 8.225 ;
      LAYER mcon ;
        RECT 0.090 5.455 2.075 8.145 ;
      LAYER met1 ;
        RECT 0.055 5.395 2.105 8.205 ;
    END
  END Rin
  PIN Rout
    DIRECTION INOUT ;
    PORT
      LAYER li1 ;
        RECT 0.000 0.575 2.160 3.425 ;
      LAYER mcon ;
        RECT 0.090 0.655 2.075 3.345 ;
      LAYER met1 ;
        RECT 0.055 0.595 2.105 3.405 ;
    END
  END Rout
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER li1 ;
        RECT 0.000 8.650 12.200 8.950 ;
      LAYER mcon ;
        RECT 0.850 8.650 1.150 8.950 ;
        RECT 1.850 8.650 2.150 8.950 ;
        RECT 2.850 8.650 3.150 8.950 ;
        RECT 3.850 8.650 4.150 8.950 ;
        RECT 4.850 8.650 5.150 8.950 ;
        RECT 5.850 8.650 6.150 8.950 ;
        RECT 6.850 8.650 7.150 8.950 ;
        RECT 7.850 8.650 8.150 8.950 ;
        RECT 8.850 8.650 9.150 8.950 ;
        RECT 9.850 8.650 10.150 8.950 ;
        RECT 10.850 8.650 11.150 8.950 ;
      LAYER met1 ;
        RECT 0.000 8.500 12.200 9.100 ;
    END
  END VPWR
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.000 -0.300 12.200 8.250 ;
      LAYER li1 ;
        RECT 4.560 0.150 7.640 4.850 ;
        RECT 0.000 -0.150 12.200 0.150 ;
      LAYER mcon ;
        RECT 0.850 -0.150 1.150 0.150 ;
        RECT 1.850 -0.150 2.150 0.150 ;
        RECT 2.850 -0.150 3.150 0.150 ;
        RECT 3.850 -0.150 4.150 0.150 ;
        RECT 4.850 -0.150 5.150 0.150 ;
        RECT 5.850 -0.150 6.150 0.150 ;
        RECT 6.850 -0.150 7.150 0.150 ;
        RECT 7.850 -0.150 8.150 0.150 ;
        RECT 8.850 -0.150 9.150 0.150 ;
        RECT 9.850 -0.150 10.150 0.150 ;
        RECT 10.850 -0.150 11.150 0.150 ;
      LAYER met1 ;
        RECT 0.000 -0.300 12.200 0.300 ;
    END
  END VGND
  OBS
      LAYER li1 ;
        RECT 10.040 0.575 12.200 8.225 ;
      LAYER mcon ;
        RECT 10.125 5.455 12.110 8.145 ;
        RECT 10.125 0.655 12.110 3.345 ;
      LAYER met1 ;
        RECT 10.095 5.395 12.145 8.205 ;
        RECT 10.040 0.575 12.200 5.395 ;
  END
END sky130_asc_res

# -------------EOF--------------------

MACRO sky130_asc_res_2
  CLASS CORE ;
  FOREIGN sky130_asc_res_2 ;
  ORIGIN 0.000 0.000 ;
  SIZE 15.070 BY 9.400 ;
  SITE unitasc ;
  PIN Rin
    DIRECTION INOUT ;
    PORT
      LAYER li1 ;
        RECT 0.005 5.375 2.165 8.225 ;
      LAYER mcon ;
        RECT 0.095 5.455 2.080 8.145 ;
      LAYER met1 ;
        RECT 0.060 5.395 2.110 8.205 ;
    END
  END Rin
  PIN Rout
    DIRECTION INOUT ;
    PORT
      LAYER li1 ;
        RECT 0.005 0.575 2.165 3.425 ;
      LAYER mcon ;
        RECT 0.095 0.655 2.080 3.345 ;
      LAYER met1 ;
        RECT 0.060 0.595 2.110 3.405 ;
    END
  END Rout
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER li1 ;
        RECT 0.010 8.650 15.070 8.950 ;
      LAYER mcon ;
        RECT 0.860 8.650 1.160 8.950 ;
        RECT 1.860 8.650 2.160 8.950 ;
        RECT 2.860 8.650 3.160 8.950 ;
        RECT 3.860 8.650 4.160 8.950 ;
        RECT 4.860 8.650 5.160 8.950 ;
        RECT 5.860 8.650 6.160 8.950 ;
        RECT 6.860 8.650 7.160 8.950 ;
        RECT 7.860 8.650 8.160 8.950 ;
        RECT 8.860 8.650 9.160 8.950 ;
        RECT 9.860 8.650 10.160 8.950 ;
        RECT 10.860 8.650 11.160 8.950 ;
        RECT 11.860 8.650 12.160 8.950 ;
        RECT 12.860 8.650 13.160 8.950 ;
        RECT 13.860 8.650 14.160 8.950 ;
      LAYER met1 ;
        RECT 0.010 8.500 15.070 9.100 ;
    END
  END VPWR
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 1.440 -0.300 13.640 8.250 ;
      LAYER li1 ;
        RECT 6.000 0.150 9.080 4.850 ;
        RECT 0.010 -0.150 15.070 0.150 ;
      LAYER mcon ;
        RECT 0.860 -0.150 1.160 0.150 ;
        RECT 1.860 -0.150 2.160 0.150 ;
        RECT 2.860 -0.150 3.160 0.150 ;
        RECT 3.860 -0.150 4.160 0.150 ;
        RECT 4.860 -0.150 5.160 0.150 ;
        RECT 5.860 -0.150 6.160 0.150 ;
        RECT 6.860 -0.150 7.160 0.150 ;
        RECT 7.860 -0.150 8.160 0.150 ;
        RECT 8.860 -0.150 9.160 0.150 ;
        RECT 9.860 -0.150 10.160 0.150 ;
        RECT 10.860 -0.150 11.160 0.150 ;
        RECT 11.860 -0.150 12.160 0.150 ;
        RECT 12.860 -0.150 13.160 0.150 ;
        RECT 13.860 -0.150 14.160 0.150 ;
      LAYER met1 ;
        RECT 0.010 -0.300 15.070 0.300 ;
    END
  END VGND
  OBS
      LAYER li1 ;
        RECT 12.915 0.575 15.075 8.225 ;
      LAYER mcon ;
        RECT 13.000 5.455 14.985 8.145 ;
        RECT 13.000 0.655 14.985 3.345 ;
      LAYER met1 ;
        RECT 12.970 5.395 15.020 8.205 ;
        RECT 12.915 0.575 15.075 5.395 ;
  END
END sky130_asc_res_2

# -------------EOF--------------------

MACRO sky130_asc_pnp_0
  CLASS CORE ;
  FOREIGN sky130_asc_pnp_0 ;
  ORIGIN 0.000 0.000 ;
  SIZE 6.700 BY 9.400 ;
  SITE unitasc ;
  PIN Emitter
    DIRECTION INOUT ;
    ANTENNADIFFAREA 11.559999 ;
    PORT
      LAYER li1 ;
        RECT 1.615 2.665 5.085 6.135 ;
      LAYER mcon ;
        RECT 1.980 5.530 2.150 5.700 ;
        RECT 2.480 5.530 2.650 5.700 ;
        RECT 2.980 5.530 3.150 5.700 ;
        RECT 3.480 5.530 3.650 5.700 ;
        RECT 3.980 5.530 4.150 5.700 ;
        RECT 4.480 5.530 4.650 5.700 ;
        RECT 1.980 5.030 2.150 5.200 ;
        RECT 2.480 5.030 2.650 5.200 ;
        RECT 2.980 5.030 3.150 5.200 ;
        RECT 3.480 5.030 3.650 5.200 ;
        RECT 3.980 5.030 4.150 5.200 ;
        RECT 4.480 5.030 4.650 5.200 ;
        RECT 1.980 4.530 2.150 4.700 ;
        RECT 2.480 4.530 2.650 4.700 ;
        RECT 2.980 4.530 3.150 4.700 ;
        RECT 3.480 4.530 3.650 4.700 ;
        RECT 3.980 4.530 4.150 4.700 ;
        RECT 4.480 4.530 4.650 4.700 ;
        RECT 1.980 4.030 2.150 4.200 ;
        RECT 2.480 4.030 2.650 4.200 ;
        RECT 2.980 4.030 3.150 4.200 ;
        RECT 3.480 4.030 3.650 4.200 ;
        RECT 3.980 4.030 4.150 4.200 ;
        RECT 4.480 4.030 4.650 4.200 ;
        RECT 1.980 3.530 2.150 3.700 ;
        RECT 2.480 3.530 2.650 3.700 ;
        RECT 2.980 3.530 3.150 3.700 ;
        RECT 3.480 3.530 3.650 3.700 ;
        RECT 3.980 3.530 4.150 3.700 ;
        RECT 4.480 3.530 4.650 3.700 ;
        RECT 1.980 3.030 2.150 3.200 ;
        RECT 2.480 3.030 2.650 3.200 ;
        RECT 2.980 3.030 3.150 3.200 ;
        RECT 3.480 3.030 3.650 3.200 ;
        RECT 3.980 3.030 4.150 3.200 ;
        RECT 4.480 3.030 4.650 3.200 ;
      LAYER met1 ;
        RECT 1.825 2.875 4.875 5.925 ;
    END
  END Emitter
  PIN Base
    DIRECTION INOUT ;
    ANTENNAGATEAREA 26.728899 ;
    ANTENNADIFFAREA 6.408000 ;
    PORT
      LAYER li1 ;
        RECT 0.945 6.445 5.755 6.805 ;
        RECT 0.945 2.355 1.305 6.445 ;
        RECT 5.395 2.355 5.755 6.445 ;
        RECT 0.945 1.995 5.755 2.355 ;
    END
  END Base
  PIN Collector
    DIRECTION INOUT ;
    ANTENNADIFFAREA 11.988700 ;
    PORT
      LAYER pwell ;
        RECT 0.000 6.985 6.700 7.750 ;
        RECT 0.000 1.815 0.765 6.985 ;
        RECT 5.935 1.815 6.700 6.985 ;
        RECT 0.000 1.050 6.700 1.815 ;
      LAYER li1 ;
        RECT 0.130 7.125 6.570 7.620 ;
        RECT 0.130 1.675 0.625 7.125 ;
        RECT 6.075 1.675 6.570 7.125 ;
        RECT 0.130 1.180 6.570 1.675 ;
    END
  END Collector
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER li1 ;
        RECT 0.000 8.650 6.700 8.950 ;
      LAYER mcon ;
        RECT 0.850 8.650 1.150 8.950 ;
        RECT 1.850 8.650 2.150 8.950 ;
        RECT 2.850 8.650 3.150 8.950 ;
        RECT 3.850 8.650 4.150 8.950 ;
        RECT 4.850 8.650 5.150 8.950 ;
        RECT 5.850 8.650 6.150 8.950 ;
      LAYER met1 ;
        RECT 0.000 8.500 6.700 9.100 ;
    END
  END VPWR
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER li1 ;
        RECT 0.000 -0.150 6.700 0.150 ;
      LAYER mcon ;
        RECT 0.850 -0.150 1.150 0.150 ;
        RECT 1.850 -0.150 2.150 0.150 ;
        RECT 2.850 -0.150 3.150 0.150 ;
        RECT 3.850 -0.150 4.150 0.150 ;
        RECT 4.850 -0.150 5.150 0.150 ;
        RECT 5.850 -0.150 6.150 0.150 ;
      LAYER met1 ;
        RECT 0.000 -0.300 6.700 0.300 ;
    END
  END VGND
END sky130_asc_pnp_0

# -------------EOF--------------------

MACRO sky130_asc_pnp_8
  CLASS CORE ;
  FOREIGN sky130_asc_pnp_8 ;
  ORIGIN 0.000 0.000 ;
  SIZE 53.600 BY 9.400 ;
  SITE unitasc ;
  PIN Emitter
    DIRECTION INOUT ;
    ANTENNADIFFAREA 92.479996 ;
    PORT
      LAYER li1 ;
        RECT 1.615 2.665 5.085 6.135 ;
        RECT 8.315 2.665 11.785 6.135 ;
        RECT 15.015 2.665 18.485 6.135 ;
        RECT 21.715 2.665 25.185 6.135 ;
        RECT 28.415 2.665 31.885 6.135 ;
        RECT 35.115 2.665 38.585 6.135 ;
        RECT 41.815 2.665 45.285 6.135 ;
        RECT 48.515 2.665 51.985 6.135 ;
      LAYER mcon ;
        RECT 1.980 5.530 2.150 5.700 ;
        RECT 2.480 5.530 2.650 5.700 ;
        RECT 2.980 5.530 3.150 5.700 ;
        RECT 3.480 5.530 3.650 5.700 ;
        RECT 3.980 5.530 4.150 5.700 ;
        RECT 4.480 5.530 4.650 5.700 ;
        RECT 1.980 5.030 2.150 5.200 ;
        RECT 2.480 5.030 2.650 5.200 ;
        RECT 2.980 5.030 3.150 5.200 ;
        RECT 3.480 5.030 3.650 5.200 ;
        RECT 3.980 5.030 4.150 5.200 ;
        RECT 4.480 5.030 4.650 5.200 ;
        RECT 1.980 4.530 2.150 4.700 ;
        RECT 2.480 4.530 2.650 4.700 ;
        RECT 2.980 4.530 3.150 4.700 ;
        RECT 3.480 4.530 3.650 4.700 ;
        RECT 3.980 4.530 4.150 4.700 ;
        RECT 4.480 4.530 4.650 4.700 ;
        RECT 1.980 4.030 2.150 4.200 ;
        RECT 2.480 4.030 2.650 4.200 ;
        RECT 2.980 4.030 3.150 4.200 ;
        RECT 3.480 4.030 3.650 4.200 ;
        RECT 3.980 4.030 4.150 4.200 ;
        RECT 4.480 4.030 4.650 4.200 ;
        RECT 1.980 3.530 2.150 3.700 ;
        RECT 2.480 3.530 2.650 3.700 ;
        RECT 2.980 3.530 3.150 3.700 ;
        RECT 3.480 3.530 3.650 3.700 ;
        RECT 3.980 3.530 4.150 3.700 ;
        RECT 4.480 3.530 4.650 3.700 ;
        RECT 1.980 3.030 2.150 3.200 ;
        RECT 2.480 3.030 2.650 3.200 ;
        RECT 2.980 3.030 3.150 3.200 ;
        RECT 3.480 3.030 3.650 3.200 ;
        RECT 3.980 3.030 4.150 3.200 ;
        RECT 4.480 3.030 4.650 3.200 ;
        RECT 8.680 5.530 8.850 5.700 ;
        RECT 9.180 5.530 9.350 5.700 ;
        RECT 9.680 5.530 9.850 5.700 ;
        RECT 10.180 5.530 10.350 5.700 ;
        RECT 10.680 5.530 10.850 5.700 ;
        RECT 11.180 5.530 11.350 5.700 ;
        RECT 8.680 5.030 8.850 5.200 ;
        RECT 9.180 5.030 9.350 5.200 ;
        RECT 9.680 5.030 9.850 5.200 ;
        RECT 10.180 5.030 10.350 5.200 ;
        RECT 10.680 5.030 10.850 5.200 ;
        RECT 11.180 5.030 11.350 5.200 ;
        RECT 8.680 4.530 8.850 4.700 ;
        RECT 9.180 4.530 9.350 4.700 ;
        RECT 9.680 4.530 9.850 4.700 ;
        RECT 10.180 4.530 10.350 4.700 ;
        RECT 10.680 4.530 10.850 4.700 ;
        RECT 11.180 4.530 11.350 4.700 ;
        RECT 8.680 4.030 8.850 4.200 ;
        RECT 9.180 4.030 9.350 4.200 ;
        RECT 9.680 4.030 9.850 4.200 ;
        RECT 10.180 4.030 10.350 4.200 ;
        RECT 10.680 4.030 10.850 4.200 ;
        RECT 11.180 4.030 11.350 4.200 ;
        RECT 8.680 3.530 8.850 3.700 ;
        RECT 9.180 3.530 9.350 3.700 ;
        RECT 9.680 3.530 9.850 3.700 ;
        RECT 10.180 3.530 10.350 3.700 ;
        RECT 10.680 3.530 10.850 3.700 ;
        RECT 11.180 3.530 11.350 3.700 ;
        RECT 8.680 3.030 8.850 3.200 ;
        RECT 9.180 3.030 9.350 3.200 ;
        RECT 9.680 3.030 9.850 3.200 ;
        RECT 10.180 3.030 10.350 3.200 ;
        RECT 10.680 3.030 10.850 3.200 ;
        RECT 11.180 3.030 11.350 3.200 ;
        RECT 15.380 5.530 15.550 5.700 ;
        RECT 15.880 5.530 16.050 5.700 ;
        RECT 16.380 5.530 16.550 5.700 ;
        RECT 16.880 5.530 17.050 5.700 ;
        RECT 17.380 5.530 17.550 5.700 ;
        RECT 17.880 5.530 18.050 5.700 ;
        RECT 15.380 5.030 15.550 5.200 ;
        RECT 15.880 5.030 16.050 5.200 ;
        RECT 16.380 5.030 16.550 5.200 ;
        RECT 16.880 5.030 17.050 5.200 ;
        RECT 17.380 5.030 17.550 5.200 ;
        RECT 17.880 5.030 18.050 5.200 ;
        RECT 15.380 4.530 15.550 4.700 ;
        RECT 15.880 4.530 16.050 4.700 ;
        RECT 16.380 4.530 16.550 4.700 ;
        RECT 16.880 4.530 17.050 4.700 ;
        RECT 17.380 4.530 17.550 4.700 ;
        RECT 17.880 4.530 18.050 4.700 ;
        RECT 15.380 4.030 15.550 4.200 ;
        RECT 15.880 4.030 16.050 4.200 ;
        RECT 16.380 4.030 16.550 4.200 ;
        RECT 16.880 4.030 17.050 4.200 ;
        RECT 17.380 4.030 17.550 4.200 ;
        RECT 17.880 4.030 18.050 4.200 ;
        RECT 15.380 3.530 15.550 3.700 ;
        RECT 15.880 3.530 16.050 3.700 ;
        RECT 16.380 3.530 16.550 3.700 ;
        RECT 16.880 3.530 17.050 3.700 ;
        RECT 17.380 3.530 17.550 3.700 ;
        RECT 17.880 3.530 18.050 3.700 ;
        RECT 15.380 3.030 15.550 3.200 ;
        RECT 15.880 3.030 16.050 3.200 ;
        RECT 16.380 3.030 16.550 3.200 ;
        RECT 16.880 3.030 17.050 3.200 ;
        RECT 17.380 3.030 17.550 3.200 ;
        RECT 17.880 3.030 18.050 3.200 ;
        RECT 22.080 5.530 22.250 5.700 ;
        RECT 22.580 5.530 22.750 5.700 ;
        RECT 23.080 5.530 23.250 5.700 ;
        RECT 23.580 5.530 23.750 5.700 ;
        RECT 24.080 5.530 24.250 5.700 ;
        RECT 24.580 5.530 24.750 5.700 ;
        RECT 22.080 5.030 22.250 5.200 ;
        RECT 22.580 5.030 22.750 5.200 ;
        RECT 23.080 5.030 23.250 5.200 ;
        RECT 23.580 5.030 23.750 5.200 ;
        RECT 24.080 5.030 24.250 5.200 ;
        RECT 24.580 5.030 24.750 5.200 ;
        RECT 22.080 4.530 22.250 4.700 ;
        RECT 22.580 4.530 22.750 4.700 ;
        RECT 23.080 4.530 23.250 4.700 ;
        RECT 23.580 4.530 23.750 4.700 ;
        RECT 24.080 4.530 24.250 4.700 ;
        RECT 24.580 4.530 24.750 4.700 ;
        RECT 22.080 4.030 22.250 4.200 ;
        RECT 22.580 4.030 22.750 4.200 ;
        RECT 23.080 4.030 23.250 4.200 ;
        RECT 23.580 4.030 23.750 4.200 ;
        RECT 24.080 4.030 24.250 4.200 ;
        RECT 24.580 4.030 24.750 4.200 ;
        RECT 22.080 3.530 22.250 3.700 ;
        RECT 22.580 3.530 22.750 3.700 ;
        RECT 23.080 3.530 23.250 3.700 ;
        RECT 23.580 3.530 23.750 3.700 ;
        RECT 24.080 3.530 24.250 3.700 ;
        RECT 24.580 3.530 24.750 3.700 ;
        RECT 22.080 3.030 22.250 3.200 ;
        RECT 22.580 3.030 22.750 3.200 ;
        RECT 23.080 3.030 23.250 3.200 ;
        RECT 23.580 3.030 23.750 3.200 ;
        RECT 24.080 3.030 24.250 3.200 ;
        RECT 24.580 3.030 24.750 3.200 ;
        RECT 28.780 5.530 28.950 5.700 ;
        RECT 29.280 5.530 29.450 5.700 ;
        RECT 29.780 5.530 29.950 5.700 ;
        RECT 30.280 5.530 30.450 5.700 ;
        RECT 30.780 5.530 30.950 5.700 ;
        RECT 31.280 5.530 31.450 5.700 ;
        RECT 28.780 5.030 28.950 5.200 ;
        RECT 29.280 5.030 29.450 5.200 ;
        RECT 29.780 5.030 29.950 5.200 ;
        RECT 30.280 5.030 30.450 5.200 ;
        RECT 30.780 5.030 30.950 5.200 ;
        RECT 31.280 5.030 31.450 5.200 ;
        RECT 28.780 4.530 28.950 4.700 ;
        RECT 29.280 4.530 29.450 4.700 ;
        RECT 29.780 4.530 29.950 4.700 ;
        RECT 30.280 4.530 30.450 4.700 ;
        RECT 30.780 4.530 30.950 4.700 ;
        RECT 31.280 4.530 31.450 4.700 ;
        RECT 28.780 4.030 28.950 4.200 ;
        RECT 29.280 4.030 29.450 4.200 ;
        RECT 29.780 4.030 29.950 4.200 ;
        RECT 30.280 4.030 30.450 4.200 ;
        RECT 30.780 4.030 30.950 4.200 ;
        RECT 31.280 4.030 31.450 4.200 ;
        RECT 28.780 3.530 28.950 3.700 ;
        RECT 29.280 3.530 29.450 3.700 ;
        RECT 29.780 3.530 29.950 3.700 ;
        RECT 30.280 3.530 30.450 3.700 ;
        RECT 30.780 3.530 30.950 3.700 ;
        RECT 31.280 3.530 31.450 3.700 ;
        RECT 28.780 3.030 28.950 3.200 ;
        RECT 29.280 3.030 29.450 3.200 ;
        RECT 29.780 3.030 29.950 3.200 ;
        RECT 30.280 3.030 30.450 3.200 ;
        RECT 30.780 3.030 30.950 3.200 ;
        RECT 31.280 3.030 31.450 3.200 ;
        RECT 35.480 5.530 35.650 5.700 ;
        RECT 35.980 5.530 36.150 5.700 ;
        RECT 36.480 5.530 36.650 5.700 ;
        RECT 36.980 5.530 37.150 5.700 ;
        RECT 37.480 5.530 37.650 5.700 ;
        RECT 37.980 5.530 38.150 5.700 ;
        RECT 35.480 5.030 35.650 5.200 ;
        RECT 35.980 5.030 36.150 5.200 ;
        RECT 36.480 5.030 36.650 5.200 ;
        RECT 36.980 5.030 37.150 5.200 ;
        RECT 37.480 5.030 37.650 5.200 ;
        RECT 37.980 5.030 38.150 5.200 ;
        RECT 35.480 4.530 35.650 4.700 ;
        RECT 35.980 4.530 36.150 4.700 ;
        RECT 36.480 4.530 36.650 4.700 ;
        RECT 36.980 4.530 37.150 4.700 ;
        RECT 37.480 4.530 37.650 4.700 ;
        RECT 37.980 4.530 38.150 4.700 ;
        RECT 35.480 4.030 35.650 4.200 ;
        RECT 35.980 4.030 36.150 4.200 ;
        RECT 36.480 4.030 36.650 4.200 ;
        RECT 36.980 4.030 37.150 4.200 ;
        RECT 37.480 4.030 37.650 4.200 ;
        RECT 37.980 4.030 38.150 4.200 ;
        RECT 35.480 3.530 35.650 3.700 ;
        RECT 35.980 3.530 36.150 3.700 ;
        RECT 36.480 3.530 36.650 3.700 ;
        RECT 36.980 3.530 37.150 3.700 ;
        RECT 37.480 3.530 37.650 3.700 ;
        RECT 37.980 3.530 38.150 3.700 ;
        RECT 35.480 3.030 35.650 3.200 ;
        RECT 35.980 3.030 36.150 3.200 ;
        RECT 36.480 3.030 36.650 3.200 ;
        RECT 36.980 3.030 37.150 3.200 ;
        RECT 37.480 3.030 37.650 3.200 ;
        RECT 37.980 3.030 38.150 3.200 ;
        RECT 42.180 5.530 42.350 5.700 ;
        RECT 42.680 5.530 42.850 5.700 ;
        RECT 43.180 5.530 43.350 5.700 ;
        RECT 43.680 5.530 43.850 5.700 ;
        RECT 44.180 5.530 44.350 5.700 ;
        RECT 44.680 5.530 44.850 5.700 ;
        RECT 42.180 5.030 42.350 5.200 ;
        RECT 42.680 5.030 42.850 5.200 ;
        RECT 43.180 5.030 43.350 5.200 ;
        RECT 43.680 5.030 43.850 5.200 ;
        RECT 44.180 5.030 44.350 5.200 ;
        RECT 44.680 5.030 44.850 5.200 ;
        RECT 42.180 4.530 42.350 4.700 ;
        RECT 42.680 4.530 42.850 4.700 ;
        RECT 43.180 4.530 43.350 4.700 ;
        RECT 43.680 4.530 43.850 4.700 ;
        RECT 44.180 4.530 44.350 4.700 ;
        RECT 44.680 4.530 44.850 4.700 ;
        RECT 42.180 4.030 42.350 4.200 ;
        RECT 42.680 4.030 42.850 4.200 ;
        RECT 43.180 4.030 43.350 4.200 ;
        RECT 43.680 4.030 43.850 4.200 ;
        RECT 44.180 4.030 44.350 4.200 ;
        RECT 44.680 4.030 44.850 4.200 ;
        RECT 42.180 3.530 42.350 3.700 ;
        RECT 42.680 3.530 42.850 3.700 ;
        RECT 43.180 3.530 43.350 3.700 ;
        RECT 43.680 3.530 43.850 3.700 ;
        RECT 44.180 3.530 44.350 3.700 ;
        RECT 44.680 3.530 44.850 3.700 ;
        RECT 42.180 3.030 42.350 3.200 ;
        RECT 42.680 3.030 42.850 3.200 ;
        RECT 43.180 3.030 43.350 3.200 ;
        RECT 43.680 3.030 43.850 3.200 ;
        RECT 44.180 3.030 44.350 3.200 ;
        RECT 44.680 3.030 44.850 3.200 ;
        RECT 48.880 5.530 49.050 5.700 ;
        RECT 49.380 5.530 49.550 5.700 ;
        RECT 49.880 5.530 50.050 5.700 ;
        RECT 50.380 5.530 50.550 5.700 ;
        RECT 50.880 5.530 51.050 5.700 ;
        RECT 51.380 5.530 51.550 5.700 ;
        RECT 48.880 5.030 49.050 5.200 ;
        RECT 49.380 5.030 49.550 5.200 ;
        RECT 49.880 5.030 50.050 5.200 ;
        RECT 50.380 5.030 50.550 5.200 ;
        RECT 50.880 5.030 51.050 5.200 ;
        RECT 51.380 5.030 51.550 5.200 ;
        RECT 48.880 4.530 49.050 4.700 ;
        RECT 49.380 4.530 49.550 4.700 ;
        RECT 49.880 4.530 50.050 4.700 ;
        RECT 50.380 4.530 50.550 4.700 ;
        RECT 50.880 4.530 51.050 4.700 ;
        RECT 51.380 4.530 51.550 4.700 ;
        RECT 48.880 4.030 49.050 4.200 ;
        RECT 49.380 4.030 49.550 4.200 ;
        RECT 49.880 4.030 50.050 4.200 ;
        RECT 50.380 4.030 50.550 4.200 ;
        RECT 50.880 4.030 51.050 4.200 ;
        RECT 51.380 4.030 51.550 4.200 ;
        RECT 48.880 3.530 49.050 3.700 ;
        RECT 49.380 3.530 49.550 3.700 ;
        RECT 49.880 3.530 50.050 3.700 ;
        RECT 50.380 3.530 50.550 3.700 ;
        RECT 50.880 3.530 51.050 3.700 ;
        RECT 51.380 3.530 51.550 3.700 ;
        RECT 48.880 3.030 49.050 3.200 ;
        RECT 49.380 3.030 49.550 3.200 ;
        RECT 49.880 3.030 50.050 3.200 ;
        RECT 50.380 3.030 50.550 3.200 ;
        RECT 50.880 3.030 51.050 3.200 ;
        RECT 51.380 3.030 51.550 3.200 ;
      LAYER met1 ;
        RECT 1.820 2.870 51.780 5.930 ;
    END
  END Emitter
  PIN Base
    DIRECTION INOUT ;
    ANTENNAGATEAREA 213.831192 ;
    ANTENNADIFFAREA 158.894394 ;
    PORT
      LAYER pwell ;
        RECT 0.000 6.985 53.600 7.750 ;
        RECT 0.000 1.815 0.765 6.985 ;
        RECT 5.935 1.815 7.465 6.985 ;
        RECT 12.635 1.815 14.165 6.985 ;
        RECT 19.335 1.815 20.865 6.985 ;
        RECT 26.035 1.815 27.565 6.985 ;
        RECT 32.735 1.815 34.265 6.985 ;
        RECT 39.435 1.815 40.965 6.985 ;
        RECT 46.135 1.815 47.665 6.985 ;
        RECT 52.835 1.815 53.600 6.985 ;
        RECT 0.000 1.050 53.600 1.815 ;
      LAYER li1 ;
        RECT 0.130 6.750 53.470 7.620 ;
        RECT 0.130 2.050 0.625 6.750 ;
        RECT 0.945 6.445 5.755 6.750 ;
        RECT 0.945 2.355 1.305 6.445 ;
        RECT 5.395 2.355 5.755 6.445 ;
        RECT 0.945 2.050 5.755 2.355 ;
        RECT 6.075 2.050 7.325 6.750 ;
        RECT 7.645 6.445 12.455 6.750 ;
        RECT 7.645 2.355 8.005 6.445 ;
        RECT 12.095 2.355 12.455 6.445 ;
        RECT 7.645 2.050 12.455 2.355 ;
        RECT 12.775 2.050 14.025 6.750 ;
        RECT 14.345 6.445 19.155 6.750 ;
        RECT 14.345 2.355 14.705 6.445 ;
        RECT 18.795 2.355 19.155 6.445 ;
        RECT 14.345 2.050 19.155 2.355 ;
        RECT 19.475 2.050 20.725 6.750 ;
        RECT 21.045 6.445 25.855 6.750 ;
        RECT 21.045 2.355 21.405 6.445 ;
        RECT 25.495 2.355 25.855 6.445 ;
        RECT 21.045 2.050 25.855 2.355 ;
        RECT 26.175 2.050 27.425 6.750 ;
        RECT 27.745 6.445 32.555 6.750 ;
        RECT 27.745 2.355 28.105 6.445 ;
        RECT 32.195 2.355 32.555 6.445 ;
        RECT 27.745 2.050 32.555 2.355 ;
        RECT 32.875 2.050 34.125 6.750 ;
        RECT 34.445 6.445 39.255 6.750 ;
        RECT 34.445 2.355 34.805 6.445 ;
        RECT 38.895 2.355 39.255 6.445 ;
        RECT 34.445 2.050 39.255 2.355 ;
        RECT 39.575 2.050 40.825 6.750 ;
        RECT 41.145 6.445 45.955 6.750 ;
        RECT 41.145 2.355 41.505 6.445 ;
        RECT 45.595 2.355 45.955 6.445 ;
        RECT 41.145 2.050 45.955 2.355 ;
        RECT 46.275 2.050 47.525 6.750 ;
        RECT 47.845 6.445 52.655 6.750 ;
        RECT 47.845 2.355 48.205 6.445 ;
        RECT 52.295 2.355 52.655 6.445 ;
        RECT 47.845 2.050 52.655 2.355 ;
        RECT 52.975 2.050 53.470 6.750 ;
        RECT 0.130 1.180 53.470 2.050 ;
    END
  END Base
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER li1 ;
        RECT 0.000 8.650 53.600 8.950 ;
      LAYER mcon ;
        RECT 0.850 8.650 1.150 8.950 ;
        RECT 1.850 8.650 2.150 8.950 ;
        RECT 2.850 8.650 3.150 8.950 ;
        RECT 3.850 8.650 4.150 8.950 ;
        RECT 4.850 8.650 5.150 8.950 ;
        RECT 5.850 8.650 6.150 8.950 ;
        RECT 6.850 8.650 7.150 8.950 ;
        RECT 7.850 8.650 8.150 8.950 ;
        RECT 8.850 8.650 9.150 8.950 ;
        RECT 9.850 8.650 10.150 8.950 ;
        RECT 10.850 8.650 11.150 8.950 ;
        RECT 11.850 8.650 12.150 8.950 ;
        RECT 12.850 8.650 13.150 8.950 ;
        RECT 13.850 8.650 14.150 8.950 ;
        RECT 14.850 8.650 15.150 8.950 ;
        RECT 15.850 8.650 16.150 8.950 ;
        RECT 16.850 8.650 17.150 8.950 ;
        RECT 17.850 8.650 18.150 8.950 ;
        RECT 18.850 8.650 19.150 8.950 ;
        RECT 19.850 8.650 20.150 8.950 ;
        RECT 20.850 8.650 21.150 8.950 ;
        RECT 21.850 8.650 22.150 8.950 ;
        RECT 22.850 8.650 23.150 8.950 ;
        RECT 23.850 8.650 24.150 8.950 ;
        RECT 24.850 8.650 25.150 8.950 ;
        RECT 25.850 8.650 26.150 8.950 ;
        RECT 26.850 8.650 27.150 8.950 ;
        RECT 27.850 8.650 28.150 8.950 ;
        RECT 28.850 8.650 29.150 8.950 ;
        RECT 29.850 8.650 30.150 8.950 ;
        RECT 30.850 8.650 31.150 8.950 ;
        RECT 31.850 8.650 32.150 8.950 ;
        RECT 32.850 8.650 33.150 8.950 ;
        RECT 33.850 8.650 34.150 8.950 ;
        RECT 34.850 8.650 35.150 8.950 ;
        RECT 35.850 8.650 36.150 8.950 ;
        RECT 36.850 8.650 37.150 8.950 ;
        RECT 37.850 8.650 38.150 8.950 ;
        RECT 38.850 8.650 39.150 8.950 ;
        RECT 39.850 8.650 40.150 8.950 ;
        RECT 40.850 8.650 41.150 8.950 ;
        RECT 41.850 8.650 42.150 8.950 ;
        RECT 42.850 8.650 43.150 8.950 ;
        RECT 43.850 8.650 44.150 8.950 ;
        RECT 44.850 8.650 45.150 8.950 ;
        RECT 45.850 8.650 46.150 8.950 ;
        RECT 46.850 8.650 47.150 8.950 ;
        RECT 47.850 8.650 48.150 8.950 ;
        RECT 48.850 8.650 49.150 8.950 ;
        RECT 49.850 8.650 50.150 8.950 ;
        RECT 50.850 8.650 51.150 8.950 ;
        RECT 51.850 8.650 52.150 8.950 ;
        RECT 52.850 8.650 53.150 8.950 ;
      LAYER met1 ;
        RECT 0.000 8.500 53.600 9.100 ;
    END
  END VPWR
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER li1 ;
        RECT 0.000 -0.150 53.600 0.150 ;
      LAYER mcon ;
        RECT 0.850 -0.150 1.150 0.150 ;
        RECT 1.850 -0.150 2.150 0.150 ;
        RECT 2.850 -0.150 3.150 0.150 ;
        RECT 3.850 -0.150 4.150 0.150 ;
        RECT 4.850 -0.150 5.150 0.150 ;
        RECT 5.850 -0.150 6.150 0.150 ;
        RECT 6.850 -0.150 7.150 0.150 ;
        RECT 7.850 -0.150 8.150 0.150 ;
        RECT 8.850 -0.150 9.150 0.150 ;
        RECT 9.850 -0.150 10.150 0.150 ;
        RECT 10.850 -0.150 11.150 0.150 ;
        RECT 11.850 -0.150 12.150 0.150 ;
        RECT 12.850 -0.150 13.150 0.150 ;
        RECT 13.850 -0.150 14.150 0.150 ;
        RECT 14.850 -0.150 15.150 0.150 ;
        RECT 15.850 -0.150 16.150 0.150 ;
        RECT 16.850 -0.150 17.150 0.150 ;
        RECT 17.850 -0.150 18.150 0.150 ;
        RECT 18.850 -0.150 19.150 0.150 ;
        RECT 19.850 -0.150 20.150 0.150 ;
        RECT 20.850 -0.150 21.150 0.150 ;
        RECT 21.850 -0.150 22.150 0.150 ;
        RECT 22.850 -0.150 23.150 0.150 ;
        RECT 23.850 -0.150 24.150 0.150 ;
        RECT 24.850 -0.150 25.150 0.150 ;
        RECT 25.850 -0.150 26.150 0.150 ;
        RECT 26.850 -0.150 27.150 0.150 ;
        RECT 27.850 -0.150 28.150 0.150 ;
        RECT 28.850 -0.150 29.150 0.150 ;
        RECT 29.850 -0.150 30.150 0.150 ;
        RECT 30.850 -0.150 31.150 0.150 ;
        RECT 31.850 -0.150 32.150 0.150 ;
        RECT 32.850 -0.150 33.150 0.150 ;
        RECT 33.850 -0.150 34.150 0.150 ;
        RECT 34.850 -0.150 35.150 0.150 ;
        RECT 35.850 -0.150 36.150 0.150 ;
        RECT 36.850 -0.150 37.150 0.150 ;
        RECT 37.850 -0.150 38.150 0.150 ;
        RECT 38.850 -0.150 39.150 0.150 ;
        RECT 39.850 -0.150 40.150 0.150 ;
        RECT 40.850 -0.150 41.150 0.150 ;
        RECT 41.850 -0.150 42.150 0.150 ;
        RECT 42.850 -0.150 43.150 0.150 ;
        RECT 43.850 -0.150 44.150 0.150 ;
        RECT 44.850 -0.150 45.150 0.150 ;
        RECT 45.850 -0.150 46.150 0.150 ;
        RECT 46.850 -0.150 47.150 0.150 ;
        RECT 47.850 -0.150 48.150 0.150 ;
        RECT 48.850 -0.150 49.150 0.150 ;
        RECT 49.850 -0.150 50.150 0.150 ;
        RECT 50.850 -0.150 51.150 0.150 ;
        RECT 51.850 -0.150 52.150 0.150 ;
        RECT 52.850 -0.150 53.150 0.150 ;
      LAYER met1 ;
        RECT 0.000 -0.300 53.600 0.300 ;
    END
  END VGND
END sky130_asc_pnp_8

# -------------EOF--------------------

MACRO sky130_asc_pnp_7
  CLASS CORE ;
  FOREIGN sky130_asc_pnp_7 ;
  ORIGIN 0.000 0.000 ;
  SIZE 46.900 BY 9.400 ;
  SITE unitasc ;
  PIN Emitter
    DIRECTION INOUT ;
    ANTENNADIFFAREA 80.919998 ;
    PORT
      LAYER li1 ;
        RECT 1.615 2.665 5.085 6.135 ;
        RECT 8.315 2.665 11.785 6.135 ;
        RECT 15.015 2.665 18.485 6.135 ;
        RECT 21.715 2.665 25.185 6.135 ;
        RECT 28.415 2.665 31.885 6.135 ;
        RECT 35.115 2.665 38.585 6.135 ;
        RECT 41.815 2.665 45.285 6.135 ;
      LAYER mcon ;
        RECT 1.980 5.530 2.150 5.700 ;
        RECT 2.480 5.530 2.650 5.700 ;
        RECT 2.980 5.530 3.150 5.700 ;
        RECT 3.480 5.530 3.650 5.700 ;
        RECT 3.980 5.530 4.150 5.700 ;
        RECT 4.480 5.530 4.650 5.700 ;
        RECT 1.980 5.030 2.150 5.200 ;
        RECT 2.480 5.030 2.650 5.200 ;
        RECT 2.980 5.030 3.150 5.200 ;
        RECT 3.480 5.030 3.650 5.200 ;
        RECT 3.980 5.030 4.150 5.200 ;
        RECT 4.480 5.030 4.650 5.200 ;
        RECT 1.980 4.530 2.150 4.700 ;
        RECT 2.480 4.530 2.650 4.700 ;
        RECT 2.980 4.530 3.150 4.700 ;
        RECT 3.480 4.530 3.650 4.700 ;
        RECT 3.980 4.530 4.150 4.700 ;
        RECT 4.480 4.530 4.650 4.700 ;
        RECT 1.980 4.030 2.150 4.200 ;
        RECT 2.480 4.030 2.650 4.200 ;
        RECT 2.980 4.030 3.150 4.200 ;
        RECT 3.480 4.030 3.650 4.200 ;
        RECT 3.980 4.030 4.150 4.200 ;
        RECT 4.480 4.030 4.650 4.200 ;
        RECT 1.980 3.530 2.150 3.700 ;
        RECT 2.480 3.530 2.650 3.700 ;
        RECT 2.980 3.530 3.150 3.700 ;
        RECT 3.480 3.530 3.650 3.700 ;
        RECT 3.980 3.530 4.150 3.700 ;
        RECT 4.480 3.530 4.650 3.700 ;
        RECT 1.980 3.030 2.150 3.200 ;
        RECT 2.480 3.030 2.650 3.200 ;
        RECT 2.980 3.030 3.150 3.200 ;
        RECT 3.480 3.030 3.650 3.200 ;
        RECT 3.980 3.030 4.150 3.200 ;
        RECT 4.480 3.030 4.650 3.200 ;
        RECT 8.680 5.530 8.850 5.700 ;
        RECT 9.180 5.530 9.350 5.700 ;
        RECT 9.680 5.530 9.850 5.700 ;
        RECT 10.180 5.530 10.350 5.700 ;
        RECT 10.680 5.530 10.850 5.700 ;
        RECT 11.180 5.530 11.350 5.700 ;
        RECT 8.680 5.030 8.850 5.200 ;
        RECT 9.180 5.030 9.350 5.200 ;
        RECT 9.680 5.030 9.850 5.200 ;
        RECT 10.180 5.030 10.350 5.200 ;
        RECT 10.680 5.030 10.850 5.200 ;
        RECT 11.180 5.030 11.350 5.200 ;
        RECT 8.680 4.530 8.850 4.700 ;
        RECT 9.180 4.530 9.350 4.700 ;
        RECT 9.680 4.530 9.850 4.700 ;
        RECT 10.180 4.530 10.350 4.700 ;
        RECT 10.680 4.530 10.850 4.700 ;
        RECT 11.180 4.530 11.350 4.700 ;
        RECT 8.680 4.030 8.850 4.200 ;
        RECT 9.180 4.030 9.350 4.200 ;
        RECT 9.680 4.030 9.850 4.200 ;
        RECT 10.180 4.030 10.350 4.200 ;
        RECT 10.680 4.030 10.850 4.200 ;
        RECT 11.180 4.030 11.350 4.200 ;
        RECT 8.680 3.530 8.850 3.700 ;
        RECT 9.180 3.530 9.350 3.700 ;
        RECT 9.680 3.530 9.850 3.700 ;
        RECT 10.180 3.530 10.350 3.700 ;
        RECT 10.680 3.530 10.850 3.700 ;
        RECT 11.180 3.530 11.350 3.700 ;
        RECT 8.680 3.030 8.850 3.200 ;
        RECT 9.180 3.030 9.350 3.200 ;
        RECT 9.680 3.030 9.850 3.200 ;
        RECT 10.180 3.030 10.350 3.200 ;
        RECT 10.680 3.030 10.850 3.200 ;
        RECT 11.180 3.030 11.350 3.200 ;
        RECT 15.380 5.530 15.550 5.700 ;
        RECT 15.880 5.530 16.050 5.700 ;
        RECT 16.380 5.530 16.550 5.700 ;
        RECT 16.880 5.530 17.050 5.700 ;
        RECT 17.380 5.530 17.550 5.700 ;
        RECT 17.880 5.530 18.050 5.700 ;
        RECT 15.380 5.030 15.550 5.200 ;
        RECT 15.880 5.030 16.050 5.200 ;
        RECT 16.380 5.030 16.550 5.200 ;
        RECT 16.880 5.030 17.050 5.200 ;
        RECT 17.380 5.030 17.550 5.200 ;
        RECT 17.880 5.030 18.050 5.200 ;
        RECT 15.380 4.530 15.550 4.700 ;
        RECT 15.880 4.530 16.050 4.700 ;
        RECT 16.380 4.530 16.550 4.700 ;
        RECT 16.880 4.530 17.050 4.700 ;
        RECT 17.380 4.530 17.550 4.700 ;
        RECT 17.880 4.530 18.050 4.700 ;
        RECT 15.380 4.030 15.550 4.200 ;
        RECT 15.880 4.030 16.050 4.200 ;
        RECT 16.380 4.030 16.550 4.200 ;
        RECT 16.880 4.030 17.050 4.200 ;
        RECT 17.380 4.030 17.550 4.200 ;
        RECT 17.880 4.030 18.050 4.200 ;
        RECT 15.380 3.530 15.550 3.700 ;
        RECT 15.880 3.530 16.050 3.700 ;
        RECT 16.380 3.530 16.550 3.700 ;
        RECT 16.880 3.530 17.050 3.700 ;
        RECT 17.380 3.530 17.550 3.700 ;
        RECT 17.880 3.530 18.050 3.700 ;
        RECT 15.380 3.030 15.550 3.200 ;
        RECT 15.880 3.030 16.050 3.200 ;
        RECT 16.380 3.030 16.550 3.200 ;
        RECT 16.880 3.030 17.050 3.200 ;
        RECT 17.380 3.030 17.550 3.200 ;
        RECT 17.880 3.030 18.050 3.200 ;
        RECT 22.080 5.530 22.250 5.700 ;
        RECT 22.580 5.530 22.750 5.700 ;
        RECT 23.080 5.530 23.250 5.700 ;
        RECT 23.580 5.530 23.750 5.700 ;
        RECT 24.080 5.530 24.250 5.700 ;
        RECT 24.580 5.530 24.750 5.700 ;
        RECT 22.080 5.030 22.250 5.200 ;
        RECT 22.580 5.030 22.750 5.200 ;
        RECT 23.080 5.030 23.250 5.200 ;
        RECT 23.580 5.030 23.750 5.200 ;
        RECT 24.080 5.030 24.250 5.200 ;
        RECT 24.580 5.030 24.750 5.200 ;
        RECT 22.080 4.530 22.250 4.700 ;
        RECT 22.580 4.530 22.750 4.700 ;
        RECT 23.080 4.530 23.250 4.700 ;
        RECT 23.580 4.530 23.750 4.700 ;
        RECT 24.080 4.530 24.250 4.700 ;
        RECT 24.580 4.530 24.750 4.700 ;
        RECT 22.080 4.030 22.250 4.200 ;
        RECT 22.580 4.030 22.750 4.200 ;
        RECT 23.080 4.030 23.250 4.200 ;
        RECT 23.580 4.030 23.750 4.200 ;
        RECT 24.080 4.030 24.250 4.200 ;
        RECT 24.580 4.030 24.750 4.200 ;
        RECT 22.080 3.530 22.250 3.700 ;
        RECT 22.580 3.530 22.750 3.700 ;
        RECT 23.080 3.530 23.250 3.700 ;
        RECT 23.580 3.530 23.750 3.700 ;
        RECT 24.080 3.530 24.250 3.700 ;
        RECT 24.580 3.530 24.750 3.700 ;
        RECT 22.080 3.030 22.250 3.200 ;
        RECT 22.580 3.030 22.750 3.200 ;
        RECT 23.080 3.030 23.250 3.200 ;
        RECT 23.580 3.030 23.750 3.200 ;
        RECT 24.080 3.030 24.250 3.200 ;
        RECT 24.580 3.030 24.750 3.200 ;
        RECT 28.780 5.530 28.950 5.700 ;
        RECT 29.280 5.530 29.450 5.700 ;
        RECT 29.780 5.530 29.950 5.700 ;
        RECT 30.280 5.530 30.450 5.700 ;
        RECT 30.780 5.530 30.950 5.700 ;
        RECT 31.280 5.530 31.450 5.700 ;
        RECT 28.780 5.030 28.950 5.200 ;
        RECT 29.280 5.030 29.450 5.200 ;
        RECT 29.780 5.030 29.950 5.200 ;
        RECT 30.280 5.030 30.450 5.200 ;
        RECT 30.780 5.030 30.950 5.200 ;
        RECT 31.280 5.030 31.450 5.200 ;
        RECT 28.780 4.530 28.950 4.700 ;
        RECT 29.280 4.530 29.450 4.700 ;
        RECT 29.780 4.530 29.950 4.700 ;
        RECT 30.280 4.530 30.450 4.700 ;
        RECT 30.780 4.530 30.950 4.700 ;
        RECT 31.280 4.530 31.450 4.700 ;
        RECT 28.780 4.030 28.950 4.200 ;
        RECT 29.280 4.030 29.450 4.200 ;
        RECT 29.780 4.030 29.950 4.200 ;
        RECT 30.280 4.030 30.450 4.200 ;
        RECT 30.780 4.030 30.950 4.200 ;
        RECT 31.280 4.030 31.450 4.200 ;
        RECT 28.780 3.530 28.950 3.700 ;
        RECT 29.280 3.530 29.450 3.700 ;
        RECT 29.780 3.530 29.950 3.700 ;
        RECT 30.280 3.530 30.450 3.700 ;
        RECT 30.780 3.530 30.950 3.700 ;
        RECT 31.280 3.530 31.450 3.700 ;
        RECT 28.780 3.030 28.950 3.200 ;
        RECT 29.280 3.030 29.450 3.200 ;
        RECT 29.780 3.030 29.950 3.200 ;
        RECT 30.280 3.030 30.450 3.200 ;
        RECT 30.780 3.030 30.950 3.200 ;
        RECT 31.280 3.030 31.450 3.200 ;
        RECT 35.480 5.530 35.650 5.700 ;
        RECT 35.980 5.530 36.150 5.700 ;
        RECT 36.480 5.530 36.650 5.700 ;
        RECT 36.980 5.530 37.150 5.700 ;
        RECT 37.480 5.530 37.650 5.700 ;
        RECT 37.980 5.530 38.150 5.700 ;
        RECT 35.480 5.030 35.650 5.200 ;
        RECT 35.980 5.030 36.150 5.200 ;
        RECT 36.480 5.030 36.650 5.200 ;
        RECT 36.980 5.030 37.150 5.200 ;
        RECT 37.480 5.030 37.650 5.200 ;
        RECT 37.980 5.030 38.150 5.200 ;
        RECT 35.480 4.530 35.650 4.700 ;
        RECT 35.980 4.530 36.150 4.700 ;
        RECT 36.480 4.530 36.650 4.700 ;
        RECT 36.980 4.530 37.150 4.700 ;
        RECT 37.480 4.530 37.650 4.700 ;
        RECT 37.980 4.530 38.150 4.700 ;
        RECT 35.480 4.030 35.650 4.200 ;
        RECT 35.980 4.030 36.150 4.200 ;
        RECT 36.480 4.030 36.650 4.200 ;
        RECT 36.980 4.030 37.150 4.200 ;
        RECT 37.480 4.030 37.650 4.200 ;
        RECT 37.980 4.030 38.150 4.200 ;
        RECT 35.480 3.530 35.650 3.700 ;
        RECT 35.980 3.530 36.150 3.700 ;
        RECT 36.480 3.530 36.650 3.700 ;
        RECT 36.980 3.530 37.150 3.700 ;
        RECT 37.480 3.530 37.650 3.700 ;
        RECT 37.980 3.530 38.150 3.700 ;
        RECT 35.480 3.030 35.650 3.200 ;
        RECT 35.980 3.030 36.150 3.200 ;
        RECT 36.480 3.030 36.650 3.200 ;
        RECT 36.980 3.030 37.150 3.200 ;
        RECT 37.480 3.030 37.650 3.200 ;
        RECT 37.980 3.030 38.150 3.200 ;
        RECT 42.180 5.530 42.350 5.700 ;
        RECT 42.680 5.530 42.850 5.700 ;
        RECT 43.180 5.530 43.350 5.700 ;
        RECT 43.680 5.530 43.850 5.700 ;
        RECT 44.180 5.530 44.350 5.700 ;
        RECT 44.680 5.530 44.850 5.700 ;
        RECT 42.180 5.030 42.350 5.200 ;
        RECT 42.680 5.030 42.850 5.200 ;
        RECT 43.180 5.030 43.350 5.200 ;
        RECT 43.680 5.030 43.850 5.200 ;
        RECT 44.180 5.030 44.350 5.200 ;
        RECT 44.680 5.030 44.850 5.200 ;
        RECT 42.180 4.530 42.350 4.700 ;
        RECT 42.680 4.530 42.850 4.700 ;
        RECT 43.180 4.530 43.350 4.700 ;
        RECT 43.680 4.530 43.850 4.700 ;
        RECT 44.180 4.530 44.350 4.700 ;
        RECT 44.680 4.530 44.850 4.700 ;
        RECT 42.180 4.030 42.350 4.200 ;
        RECT 42.680 4.030 42.850 4.200 ;
        RECT 43.180 4.030 43.350 4.200 ;
        RECT 43.680 4.030 43.850 4.200 ;
        RECT 44.180 4.030 44.350 4.200 ;
        RECT 44.680 4.030 44.850 4.200 ;
        RECT 42.180 3.530 42.350 3.700 ;
        RECT 42.680 3.530 42.850 3.700 ;
        RECT 43.180 3.530 43.350 3.700 ;
        RECT 43.680 3.530 43.850 3.700 ;
        RECT 44.180 3.530 44.350 3.700 ;
        RECT 44.680 3.530 44.850 3.700 ;
        RECT 42.180 3.030 42.350 3.200 ;
        RECT 42.680 3.030 42.850 3.200 ;
        RECT 43.180 3.030 43.350 3.200 ;
        RECT 43.680 3.030 43.850 3.200 ;
        RECT 44.180 3.030 44.350 3.200 ;
        RECT 44.680 3.030 44.850 3.200 ;
      LAYER met1 ;
        RECT 1.820 2.870 45.310 5.930 ;
    END
  END Emitter
  PIN Base
    DIRECTION INOUT ;
    ANTENNAGATEAREA 187.102295 ;
    ANTENNADIFFAREA 138.823303 ;
    PORT
      LAYER pwell ;
        RECT 0.000 6.985 46.900 7.750 ;
        RECT 0.000 1.815 0.765 6.985 ;
        RECT 5.935 1.815 7.465 6.985 ;
        RECT 12.635 1.815 14.165 6.985 ;
        RECT 19.335 1.815 20.865 6.985 ;
        RECT 26.035 1.815 27.565 6.985 ;
        RECT 32.735 1.815 34.265 6.985 ;
        RECT 39.435 1.815 40.965 6.985 ;
        RECT 46.135 1.815 46.900 6.985 ;
        RECT 0.000 1.050 46.900 1.815 ;
      LAYER li1 ;
        RECT 0.130 6.750 46.785 7.620 ;
        RECT 0.130 2.050 0.625 6.750 ;
        RECT 0.945 6.445 5.755 6.750 ;
        RECT 0.945 2.355 1.305 6.445 ;
        RECT 5.395 2.355 5.755 6.445 ;
        RECT 0.945 2.050 5.755 2.355 ;
        RECT 6.075 2.050 7.325 6.750 ;
        RECT 7.645 6.445 12.455 6.750 ;
        RECT 7.645 2.355 8.005 6.445 ;
        RECT 12.095 2.355 12.455 6.445 ;
        RECT 7.645 2.050 12.455 2.355 ;
        RECT 12.775 2.050 14.025 6.750 ;
        RECT 14.345 6.445 19.155 6.750 ;
        RECT 14.345 2.355 14.705 6.445 ;
        RECT 18.795 2.355 19.155 6.445 ;
        RECT 14.345 2.050 19.155 2.355 ;
        RECT 19.475 2.050 20.725 6.750 ;
        RECT 21.045 6.445 25.855 6.750 ;
        RECT 21.045 2.355 21.405 6.445 ;
        RECT 25.495 2.355 25.855 6.445 ;
        RECT 21.045 2.050 25.855 2.355 ;
        RECT 26.175 2.050 27.425 6.750 ;
        RECT 27.745 6.445 32.555 6.750 ;
        RECT 27.745 2.355 28.105 6.445 ;
        RECT 32.195 2.355 32.555 6.445 ;
        RECT 27.745 2.050 32.555 2.355 ;
        RECT 32.875 2.050 34.125 6.750 ;
        RECT 34.445 6.445 39.255 6.750 ;
        RECT 34.445 2.355 34.805 6.445 ;
        RECT 38.895 2.355 39.255 6.445 ;
        RECT 34.445 2.050 39.255 2.355 ;
        RECT 39.575 2.050 40.825 6.750 ;
        RECT 41.145 6.445 45.955 6.750 ;
        RECT 41.145 2.355 41.505 6.445 ;
        RECT 45.595 2.355 45.955 6.445 ;
        RECT 41.145 2.050 45.955 2.355 ;
        RECT 46.275 2.050 46.770 6.750 ;
        RECT 0.130 1.180 46.785 2.050 ;
    END
  END Base
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER li1 ;
        RECT 0.000 8.650 46.900 8.950 ;
      LAYER mcon ;
        RECT 0.850 8.650 1.150 8.950 ;
        RECT 1.850 8.650 2.150 8.950 ;
        RECT 2.850 8.650 3.150 8.950 ;
        RECT 3.850 8.650 4.150 8.950 ;
        RECT 4.850 8.650 5.150 8.950 ;
        RECT 5.850 8.650 6.150 8.950 ;
        RECT 6.850 8.650 7.150 8.950 ;
        RECT 7.850 8.650 8.150 8.950 ;
        RECT 8.850 8.650 9.150 8.950 ;
        RECT 9.850 8.650 10.150 8.950 ;
        RECT 10.850 8.650 11.150 8.950 ;
        RECT 11.850 8.650 12.150 8.950 ;
        RECT 12.850 8.650 13.150 8.950 ;
        RECT 13.850 8.650 14.150 8.950 ;
        RECT 14.850 8.650 15.150 8.950 ;
        RECT 15.850 8.650 16.150 8.950 ;
        RECT 16.850 8.650 17.150 8.950 ;
        RECT 17.850 8.650 18.150 8.950 ;
        RECT 18.850 8.650 19.150 8.950 ;
        RECT 19.850 8.650 20.150 8.950 ;
        RECT 20.850 8.650 21.150 8.950 ;
        RECT 21.850 8.650 22.150 8.950 ;
        RECT 22.850 8.650 23.150 8.950 ;
        RECT 23.850 8.650 24.150 8.950 ;
        RECT 24.850 8.650 25.150 8.950 ;
        RECT 25.850 8.650 26.150 8.950 ;
        RECT 26.850 8.650 27.150 8.950 ;
        RECT 27.850 8.650 28.150 8.950 ;
        RECT 28.850 8.650 29.150 8.950 ;
        RECT 29.850 8.650 30.150 8.950 ;
        RECT 30.850 8.650 31.150 8.950 ;
        RECT 31.850 8.650 32.150 8.950 ;
        RECT 32.850 8.650 33.150 8.950 ;
        RECT 33.850 8.650 34.150 8.950 ;
        RECT 34.850 8.650 35.150 8.950 ;
        RECT 35.850 8.650 36.150 8.950 ;
        RECT 36.850 8.650 37.150 8.950 ;
        RECT 37.850 8.650 38.150 8.950 ;
        RECT 38.850 8.650 39.150 8.950 ;
        RECT 39.850 8.650 40.150 8.950 ;
        RECT 40.850 8.650 41.150 8.950 ;
        RECT 41.850 8.650 42.150 8.950 ;
        RECT 42.850 8.650 43.150 8.950 ;
        RECT 43.850 8.650 44.150 8.950 ;
        RECT 44.850 8.650 45.150 8.950 ;
        RECT 45.850 8.650 46.150 8.950 ;
      LAYER met1 ;
        RECT 0.000 8.500 46.900 9.100 ;
    END
  END VPWR
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER li1 ;
        RECT 0.000 -0.150 46.900 0.150 ;
      LAYER mcon ;
        RECT 0.850 -0.150 1.150 0.150 ;
        RECT 1.850 -0.150 2.150 0.150 ;
        RECT 2.850 -0.150 3.150 0.150 ;
        RECT 3.850 -0.150 4.150 0.150 ;
        RECT 4.850 -0.150 5.150 0.150 ;
        RECT 5.850 -0.150 6.150 0.150 ;
        RECT 6.850 -0.150 7.150 0.150 ;
        RECT 7.850 -0.150 8.150 0.150 ;
        RECT 8.850 -0.150 9.150 0.150 ;
        RECT 9.850 -0.150 10.150 0.150 ;
        RECT 10.850 -0.150 11.150 0.150 ;
        RECT 11.850 -0.150 12.150 0.150 ;
        RECT 12.850 -0.150 13.150 0.150 ;
        RECT 13.850 -0.150 14.150 0.150 ;
        RECT 14.850 -0.150 15.150 0.150 ;
        RECT 15.850 -0.150 16.150 0.150 ;
        RECT 16.850 -0.150 17.150 0.150 ;
        RECT 17.850 -0.150 18.150 0.150 ;
        RECT 18.850 -0.150 19.150 0.150 ;
        RECT 19.850 -0.150 20.150 0.150 ;
        RECT 20.850 -0.150 21.150 0.150 ;
        RECT 21.850 -0.150 22.150 0.150 ;
        RECT 22.850 -0.150 23.150 0.150 ;
        RECT 23.850 -0.150 24.150 0.150 ;
        RECT 24.850 -0.150 25.150 0.150 ;
        RECT 25.850 -0.150 26.150 0.150 ;
        RECT 26.850 -0.150 27.150 0.150 ;
        RECT 27.850 -0.150 28.150 0.150 ;
        RECT 28.850 -0.150 29.150 0.150 ;
        RECT 29.850 -0.150 30.150 0.150 ;
        RECT 30.850 -0.150 31.150 0.150 ;
        RECT 31.850 -0.150 32.150 0.150 ;
        RECT 32.850 -0.150 33.150 0.150 ;
        RECT 33.850 -0.150 34.150 0.150 ;
        RECT 34.850 -0.150 35.150 0.150 ;
        RECT 35.850 -0.150 36.150 0.150 ;
        RECT 36.850 -0.150 37.150 0.150 ;
        RECT 37.850 -0.150 38.150 0.150 ;
        RECT 38.850 -0.150 39.150 0.150 ;
        RECT 39.850 -0.150 40.150 0.150 ;
        RECT 40.850 -0.150 41.150 0.150 ;
        RECT 41.850 -0.150 42.150 0.150 ;
        RECT 42.850 -0.150 43.150 0.150 ;
        RECT 43.850 -0.150 44.150 0.150 ;
        RECT 44.850 -0.150 45.150 0.150 ;
        RECT 45.850 -0.150 46.150 0.150 ;
      LAYER met1 ;
        RECT 0.000 -0.300 46.900 0.300 ;
    END
  END VGND
END sky130_asc_pnp_7

# -------------EOF--------------------

MACRO sky130_fd_sc_hd__inv_2
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__inv_2 ;
  ORIGIN 0.000 0.000 ;
  SIZE 1.380 BY 2.720 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.495000 ;
    PORT
      LAYER li1 ;
        RECT 0.105 1.075 0.435 1.325 ;
    END
  END A
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met1 ;
        RECT 0.000 -0.240 1.380 0.240 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.015 0.105 1.365 1.015 ;
        RECT 0.145 -0.085 0.315 0.105 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190 1.305 1.570 2.910 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met1 ;
        RECT 0.000 2.480 1.380 2.960 ;
    END
  END VPWR
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER li1 ;
        RECT 0.525 1.485 0.855 2.465 ;
        RECT 0.605 0.885 0.855 1.485 ;
        RECT 0.525 0.255 0.855 0.885 ;
    END
  END Y
  OBS
      LAYER li1 ;
        RECT 0.000 2.635 1.380 2.805 ;
        RECT 0.125 1.495 0.355 2.635 ;
        RECT 1.025 1.495 1.235 2.635 ;
        RECT 0.125 0.085 0.355 0.905 ;
        RECT 1.025 0.085 1.235 0.905 ;
        RECT 0.000 -0.085 1.380 0.085 ;
      LAYER mcon ;
        RECT 0.145 2.635 0.315 2.805 ;
        RECT 0.605 2.635 0.775 2.805 ;
        RECT 1.065 2.635 1.235 2.805 ;
        RECT 0.145 -0.085 0.315 0.085 ;
        RECT 0.605 -0.085 0.775 0.085 ;
        RECT 1.065 -0.085 1.235 0.085 ;
  END
END sky130_fd_sc_hd__inv_2

END LIBRARY





