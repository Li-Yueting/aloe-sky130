magic
tech sky130A
magscale 1 2
timestamp 1654322491
<< nwell >>
rect 1774 552 5048 556
rect -379 190 5048 552
rect -379 -94 5046 190
rect -379 -98 1941 -94
rect 4694 -113 5046 -94
<< pwell >>
rect 3042 -106 3298 -94
rect 611 -110 4579 -106
rect -369 -170 4579 -110
rect -369 -171 4852 -170
rect -369 -233 4966 -171
rect -369 -357 4967 -233
rect -369 -391 4979 -357
rect -369 -494 4967 -391
rect -369 -498 3298 -494
rect -369 -552 905 -498
rect 1784 -548 3298 -498
rect 3305 -547 4967 -494
rect 3305 -548 4579 -547
rect 3042 -558 3298 -548
<< nmos >>
rect -179 -352 -149 -248
rect -83 -352 -53 -248
rect 13 -352 43 -248
rect 109 -352 139 -248
rect 205 -352 235 -248
rect 301 -352 331 -248
rect 397 -352 427 -248
rect 493 -352 523 -248
rect 589 -352 619 -248
rect 685 -352 715 -248
rect 1974 -348 2004 -244
rect 2070 -348 2100 -244
rect 2166 -348 2196 -244
rect 2262 -348 2292 -244
rect 2358 -348 2388 -244
rect 2454 -348 2484 -244
rect 2550 -348 2580 -244
rect 2646 -348 2676 -244
rect 2742 -348 2772 -244
rect 2838 -348 2868 -244
rect 3151 -340 3181 -240
rect 3495 -348 3525 -244
rect 3591 -348 3621 -244
rect 3687 -348 3717 -244
rect 3783 -348 3813 -244
rect 3879 -348 3909 -244
rect 3975 -348 4005 -244
rect 4071 -348 4101 -244
rect 4167 -348 4197 -244
rect 4263 -348 4293 -244
rect 4359 -348 4389 -244
<< scnmos >>
rect 4858 -327 4888 -197
<< pmos >>
rect -179 60 -149 332
rect -83 60 -53 332
rect 13 60 43 332
rect 109 60 139 332
rect 205 60 235 332
rect 301 60 331 332
rect 397 60 427 332
rect 493 60 523 332
rect 589 60 619 332
rect 685 60 715 332
rect 1974 64 2004 336
rect 2070 64 2100 336
rect 2166 64 2196 336
rect 2262 64 2292 336
rect 2358 64 2388 336
rect 2454 64 2484 336
rect 2550 64 2580 336
rect 2646 64 2676 336
rect 2742 64 2772 336
rect 2838 64 2868 336
rect 3495 64 3525 336
rect 3591 64 3621 336
rect 3687 64 3717 336
rect 3783 64 3813 336
rect 3879 64 3909 336
rect 3975 64 4005 336
rect 4071 64 4101 336
rect 4167 64 4197 336
rect 4263 64 4293 336
rect 4359 64 4389 336
<< scpmoshvt >>
rect 4858 -77 4888 123
<< ndiff >>
rect -241 -283 -179 -248
rect -241 -317 -229 -283
rect -195 -317 -179 -283
rect -241 -352 -179 -317
rect -149 -283 -83 -248
rect -149 -317 -133 -283
rect -99 -317 -83 -283
rect -149 -352 -83 -317
rect -53 -283 13 -248
rect -53 -317 -37 -283
rect -3 -317 13 -283
rect -53 -352 13 -317
rect 43 -283 109 -248
rect 43 -317 59 -283
rect 93 -317 109 -283
rect 43 -352 109 -317
rect 139 -283 205 -248
rect 139 -317 155 -283
rect 189 -317 205 -283
rect 139 -352 205 -317
rect 235 -283 301 -248
rect 235 -317 251 -283
rect 285 -317 301 -283
rect 235 -352 301 -317
rect 331 -283 397 -248
rect 331 -317 347 -283
rect 381 -317 397 -283
rect 331 -352 397 -317
rect 427 -283 493 -248
rect 427 -317 443 -283
rect 477 -317 493 -283
rect 427 -352 493 -317
rect 523 -283 589 -248
rect 523 -317 539 -283
rect 573 -317 589 -283
rect 523 -352 589 -317
rect 619 -283 685 -248
rect 619 -317 635 -283
rect 669 -317 685 -283
rect 619 -352 685 -317
rect 715 -283 777 -248
rect 715 -317 731 -283
rect 765 -317 777 -283
rect 715 -352 777 -317
rect 1912 -279 1974 -244
rect 1912 -313 1924 -279
rect 1958 -313 1974 -279
rect 1912 -348 1974 -313
rect 2004 -279 2070 -244
rect 2004 -313 2020 -279
rect 2054 -313 2070 -279
rect 2004 -348 2070 -313
rect 2100 -279 2166 -244
rect 2100 -313 2116 -279
rect 2150 -313 2166 -279
rect 2100 -348 2166 -313
rect 2196 -279 2262 -244
rect 2196 -313 2212 -279
rect 2246 -313 2262 -279
rect 2196 -348 2262 -313
rect 2292 -279 2358 -244
rect 2292 -313 2308 -279
rect 2342 -313 2358 -279
rect 2292 -348 2358 -313
rect 2388 -279 2454 -244
rect 2388 -313 2404 -279
rect 2438 -313 2454 -279
rect 2388 -348 2454 -313
rect 2484 -279 2550 -244
rect 2484 -313 2500 -279
rect 2534 -313 2550 -279
rect 2484 -348 2550 -313
rect 2580 -279 2646 -244
rect 2580 -313 2596 -279
rect 2630 -313 2646 -279
rect 2580 -348 2646 -313
rect 2676 -279 2742 -244
rect 2676 -313 2692 -279
rect 2726 -313 2742 -279
rect 2676 -348 2742 -313
rect 2772 -279 2838 -244
rect 2772 -313 2788 -279
rect 2822 -313 2838 -279
rect 2772 -348 2838 -313
rect 2868 -279 2930 -244
rect 2868 -313 2884 -279
rect 2918 -313 2930 -279
rect 2868 -348 2930 -313
rect 3093 -252 3151 -240
rect 3093 -328 3105 -252
rect 3139 -328 3151 -252
rect 3093 -340 3151 -328
rect 3181 -252 3239 -240
rect 3181 -328 3193 -252
rect 3227 -328 3239 -252
rect 3181 -340 3239 -328
rect 3433 -279 3495 -244
rect 3433 -313 3445 -279
rect 3479 -313 3495 -279
rect 3433 -348 3495 -313
rect 3525 -279 3591 -244
rect 3525 -313 3541 -279
rect 3575 -313 3591 -279
rect 3525 -348 3591 -313
rect 3621 -279 3687 -244
rect 3621 -313 3637 -279
rect 3671 -313 3687 -279
rect 3621 -348 3687 -313
rect 3717 -279 3783 -244
rect 3717 -313 3733 -279
rect 3767 -313 3783 -279
rect 3717 -348 3783 -313
rect 3813 -279 3879 -244
rect 3813 -313 3829 -279
rect 3863 -313 3879 -279
rect 3813 -348 3879 -313
rect 3909 -279 3975 -244
rect 3909 -313 3925 -279
rect 3959 -313 3975 -279
rect 3909 -348 3975 -313
rect 4005 -279 4071 -244
rect 4005 -313 4021 -279
rect 4055 -313 4071 -279
rect 4005 -348 4071 -313
rect 4101 -279 4167 -244
rect 4101 -313 4117 -279
rect 4151 -313 4167 -279
rect 4101 -348 4167 -313
rect 4197 -279 4263 -244
rect 4197 -313 4213 -279
rect 4247 -313 4263 -279
rect 4197 -348 4263 -313
rect 4293 -279 4359 -244
rect 4293 -313 4309 -279
rect 4343 -313 4359 -279
rect 4293 -348 4359 -313
rect 4389 -279 4451 -244
rect 4389 -313 4405 -279
rect 4439 -313 4451 -279
rect 4389 -348 4451 -313
rect 4806 -209 4858 -197
rect 4806 -243 4814 -209
rect 4848 -243 4858 -209
rect 4806 -277 4858 -243
rect 4806 -311 4814 -277
rect 4848 -311 4858 -277
rect 4806 -327 4858 -311
rect 4888 -209 4940 -197
rect 4888 -243 4898 -209
rect 4932 -243 4940 -209
rect 4888 -277 4940 -243
rect 4888 -311 4898 -277
rect 4932 -311 4940 -277
rect 4888 -327 4940 -311
<< pdiff >>
rect -241 315 -179 332
rect -241 281 -229 315
rect -195 281 -179 315
rect -241 247 -179 281
rect -241 213 -229 247
rect -195 213 -179 247
rect -241 179 -179 213
rect -241 145 -229 179
rect -195 145 -179 179
rect -241 111 -179 145
rect -241 77 -229 111
rect -195 77 -179 111
rect -241 60 -179 77
rect -149 315 -83 332
rect -149 281 -133 315
rect -99 281 -83 315
rect -149 247 -83 281
rect -149 213 -133 247
rect -99 213 -83 247
rect -149 179 -83 213
rect -149 145 -133 179
rect -99 145 -83 179
rect -149 111 -83 145
rect -149 77 -133 111
rect -99 77 -83 111
rect -149 60 -83 77
rect -53 315 13 332
rect -53 281 -37 315
rect -3 281 13 315
rect -53 247 13 281
rect -53 213 -37 247
rect -3 213 13 247
rect -53 179 13 213
rect -53 145 -37 179
rect -3 145 13 179
rect -53 111 13 145
rect -53 77 -37 111
rect -3 77 13 111
rect -53 60 13 77
rect 43 315 109 332
rect 43 281 59 315
rect 93 281 109 315
rect 43 247 109 281
rect 43 213 59 247
rect 93 213 109 247
rect 43 179 109 213
rect 43 145 59 179
rect 93 145 109 179
rect 43 111 109 145
rect 43 77 59 111
rect 93 77 109 111
rect 43 60 109 77
rect 139 315 205 332
rect 139 281 155 315
rect 189 281 205 315
rect 139 247 205 281
rect 139 213 155 247
rect 189 213 205 247
rect 139 179 205 213
rect 139 145 155 179
rect 189 145 205 179
rect 139 111 205 145
rect 139 77 155 111
rect 189 77 205 111
rect 139 60 205 77
rect 235 315 301 332
rect 235 281 251 315
rect 285 281 301 315
rect 235 247 301 281
rect 235 213 251 247
rect 285 213 301 247
rect 235 179 301 213
rect 235 145 251 179
rect 285 145 301 179
rect 235 111 301 145
rect 235 77 251 111
rect 285 77 301 111
rect 235 60 301 77
rect 331 315 397 332
rect 331 281 347 315
rect 381 281 397 315
rect 331 247 397 281
rect 331 213 347 247
rect 381 213 397 247
rect 331 179 397 213
rect 331 145 347 179
rect 381 145 397 179
rect 331 111 397 145
rect 331 77 347 111
rect 381 77 397 111
rect 331 60 397 77
rect 427 315 493 332
rect 427 281 443 315
rect 477 281 493 315
rect 427 247 493 281
rect 427 213 443 247
rect 477 213 493 247
rect 427 179 493 213
rect 427 145 443 179
rect 477 145 493 179
rect 427 111 493 145
rect 427 77 443 111
rect 477 77 493 111
rect 427 60 493 77
rect 523 315 589 332
rect 523 281 539 315
rect 573 281 589 315
rect 523 247 589 281
rect 523 213 539 247
rect 573 213 589 247
rect 523 179 589 213
rect 523 145 539 179
rect 573 145 589 179
rect 523 111 589 145
rect 523 77 539 111
rect 573 77 589 111
rect 523 60 589 77
rect 619 315 685 332
rect 619 281 635 315
rect 669 281 685 315
rect 619 247 685 281
rect 619 213 635 247
rect 669 213 685 247
rect 619 179 685 213
rect 619 145 635 179
rect 669 145 685 179
rect 619 111 685 145
rect 619 77 635 111
rect 669 77 685 111
rect 619 60 685 77
rect 715 315 777 332
rect 715 281 731 315
rect 765 281 777 315
rect 715 247 777 281
rect 715 213 731 247
rect 765 213 777 247
rect 715 179 777 213
rect 715 145 731 179
rect 765 145 777 179
rect 715 111 777 145
rect 715 77 731 111
rect 765 77 777 111
rect 715 60 777 77
rect 1912 319 1974 336
rect 1912 285 1924 319
rect 1958 285 1974 319
rect 1912 251 1974 285
rect 1912 217 1924 251
rect 1958 217 1974 251
rect 1912 183 1974 217
rect 1912 149 1924 183
rect 1958 149 1974 183
rect 1912 115 1974 149
rect 1912 81 1924 115
rect 1958 81 1974 115
rect 1912 64 1974 81
rect 2004 319 2070 336
rect 2004 285 2020 319
rect 2054 285 2070 319
rect 2004 251 2070 285
rect 2004 217 2020 251
rect 2054 217 2070 251
rect 2004 183 2070 217
rect 2004 149 2020 183
rect 2054 149 2070 183
rect 2004 115 2070 149
rect 2004 81 2020 115
rect 2054 81 2070 115
rect 2004 64 2070 81
rect 2100 319 2166 336
rect 2100 285 2116 319
rect 2150 285 2166 319
rect 2100 251 2166 285
rect 2100 217 2116 251
rect 2150 217 2166 251
rect 2100 183 2166 217
rect 2100 149 2116 183
rect 2150 149 2166 183
rect 2100 115 2166 149
rect 2100 81 2116 115
rect 2150 81 2166 115
rect 2100 64 2166 81
rect 2196 319 2262 336
rect 2196 285 2212 319
rect 2246 285 2262 319
rect 2196 251 2262 285
rect 2196 217 2212 251
rect 2246 217 2262 251
rect 2196 183 2262 217
rect 2196 149 2212 183
rect 2246 149 2262 183
rect 2196 115 2262 149
rect 2196 81 2212 115
rect 2246 81 2262 115
rect 2196 64 2262 81
rect 2292 319 2358 336
rect 2292 285 2308 319
rect 2342 285 2358 319
rect 2292 251 2358 285
rect 2292 217 2308 251
rect 2342 217 2358 251
rect 2292 183 2358 217
rect 2292 149 2308 183
rect 2342 149 2358 183
rect 2292 115 2358 149
rect 2292 81 2308 115
rect 2342 81 2358 115
rect 2292 64 2358 81
rect 2388 319 2454 336
rect 2388 285 2404 319
rect 2438 285 2454 319
rect 2388 251 2454 285
rect 2388 217 2404 251
rect 2438 217 2454 251
rect 2388 183 2454 217
rect 2388 149 2404 183
rect 2438 149 2454 183
rect 2388 115 2454 149
rect 2388 81 2404 115
rect 2438 81 2454 115
rect 2388 64 2454 81
rect 2484 319 2550 336
rect 2484 285 2500 319
rect 2534 285 2550 319
rect 2484 251 2550 285
rect 2484 217 2500 251
rect 2534 217 2550 251
rect 2484 183 2550 217
rect 2484 149 2500 183
rect 2534 149 2550 183
rect 2484 115 2550 149
rect 2484 81 2500 115
rect 2534 81 2550 115
rect 2484 64 2550 81
rect 2580 319 2646 336
rect 2580 285 2596 319
rect 2630 285 2646 319
rect 2580 251 2646 285
rect 2580 217 2596 251
rect 2630 217 2646 251
rect 2580 183 2646 217
rect 2580 149 2596 183
rect 2630 149 2646 183
rect 2580 115 2646 149
rect 2580 81 2596 115
rect 2630 81 2646 115
rect 2580 64 2646 81
rect 2676 319 2742 336
rect 2676 285 2692 319
rect 2726 285 2742 319
rect 2676 251 2742 285
rect 2676 217 2692 251
rect 2726 217 2742 251
rect 2676 183 2742 217
rect 2676 149 2692 183
rect 2726 149 2742 183
rect 2676 115 2742 149
rect 2676 81 2692 115
rect 2726 81 2742 115
rect 2676 64 2742 81
rect 2772 319 2838 336
rect 2772 285 2788 319
rect 2822 285 2838 319
rect 2772 251 2838 285
rect 2772 217 2788 251
rect 2822 217 2838 251
rect 2772 183 2838 217
rect 2772 149 2788 183
rect 2822 149 2838 183
rect 2772 115 2838 149
rect 2772 81 2788 115
rect 2822 81 2838 115
rect 2772 64 2838 81
rect 2868 319 2930 336
rect 2868 285 2884 319
rect 2918 285 2930 319
rect 2868 251 2930 285
rect 2868 217 2884 251
rect 2918 217 2930 251
rect 2868 183 2930 217
rect 2868 149 2884 183
rect 2918 149 2930 183
rect 2868 115 2930 149
rect 2868 81 2884 115
rect 2918 81 2930 115
rect 2868 64 2930 81
rect 3433 319 3495 336
rect 3433 285 3445 319
rect 3479 285 3495 319
rect 3433 251 3495 285
rect 3433 217 3445 251
rect 3479 217 3495 251
rect 3433 183 3495 217
rect 3433 149 3445 183
rect 3479 149 3495 183
rect 3433 115 3495 149
rect 3433 81 3445 115
rect 3479 81 3495 115
rect 3433 64 3495 81
rect 3525 319 3591 336
rect 3525 285 3541 319
rect 3575 285 3591 319
rect 3525 251 3591 285
rect 3525 217 3541 251
rect 3575 217 3591 251
rect 3525 183 3591 217
rect 3525 149 3541 183
rect 3575 149 3591 183
rect 3525 115 3591 149
rect 3525 81 3541 115
rect 3575 81 3591 115
rect 3525 64 3591 81
rect 3621 319 3687 336
rect 3621 285 3637 319
rect 3671 285 3687 319
rect 3621 251 3687 285
rect 3621 217 3637 251
rect 3671 217 3687 251
rect 3621 183 3687 217
rect 3621 149 3637 183
rect 3671 149 3687 183
rect 3621 115 3687 149
rect 3621 81 3637 115
rect 3671 81 3687 115
rect 3621 64 3687 81
rect 3717 319 3783 336
rect 3717 285 3733 319
rect 3767 285 3783 319
rect 3717 251 3783 285
rect 3717 217 3733 251
rect 3767 217 3783 251
rect 3717 183 3783 217
rect 3717 149 3733 183
rect 3767 149 3783 183
rect 3717 115 3783 149
rect 3717 81 3733 115
rect 3767 81 3783 115
rect 3717 64 3783 81
rect 3813 319 3879 336
rect 3813 285 3829 319
rect 3863 285 3879 319
rect 3813 251 3879 285
rect 3813 217 3829 251
rect 3863 217 3879 251
rect 3813 183 3879 217
rect 3813 149 3829 183
rect 3863 149 3879 183
rect 3813 115 3879 149
rect 3813 81 3829 115
rect 3863 81 3879 115
rect 3813 64 3879 81
rect 3909 319 3975 336
rect 3909 285 3925 319
rect 3959 285 3975 319
rect 3909 251 3975 285
rect 3909 217 3925 251
rect 3959 217 3975 251
rect 3909 183 3975 217
rect 3909 149 3925 183
rect 3959 149 3975 183
rect 3909 115 3975 149
rect 3909 81 3925 115
rect 3959 81 3975 115
rect 3909 64 3975 81
rect 4005 319 4071 336
rect 4005 285 4021 319
rect 4055 285 4071 319
rect 4005 251 4071 285
rect 4005 217 4021 251
rect 4055 217 4071 251
rect 4005 183 4071 217
rect 4005 149 4021 183
rect 4055 149 4071 183
rect 4005 115 4071 149
rect 4005 81 4021 115
rect 4055 81 4071 115
rect 4005 64 4071 81
rect 4101 319 4167 336
rect 4101 285 4117 319
rect 4151 285 4167 319
rect 4101 251 4167 285
rect 4101 217 4117 251
rect 4151 217 4167 251
rect 4101 183 4167 217
rect 4101 149 4117 183
rect 4151 149 4167 183
rect 4101 115 4167 149
rect 4101 81 4117 115
rect 4151 81 4167 115
rect 4101 64 4167 81
rect 4197 319 4263 336
rect 4197 285 4213 319
rect 4247 285 4263 319
rect 4197 251 4263 285
rect 4197 217 4213 251
rect 4247 217 4263 251
rect 4197 183 4263 217
rect 4197 149 4213 183
rect 4247 149 4263 183
rect 4197 115 4263 149
rect 4197 81 4213 115
rect 4247 81 4263 115
rect 4197 64 4263 81
rect 4293 319 4359 336
rect 4293 285 4309 319
rect 4343 285 4359 319
rect 4293 251 4359 285
rect 4293 217 4309 251
rect 4343 217 4359 251
rect 4293 183 4359 217
rect 4293 149 4309 183
rect 4343 149 4359 183
rect 4293 115 4359 149
rect 4293 81 4309 115
rect 4343 81 4359 115
rect 4293 64 4359 81
rect 4389 319 4451 336
rect 4389 285 4405 319
rect 4439 285 4451 319
rect 4389 251 4451 285
rect 4389 217 4405 251
rect 4439 217 4451 251
rect 4389 183 4451 217
rect 4389 149 4405 183
rect 4439 149 4451 183
rect 4389 115 4451 149
rect 4389 81 4405 115
rect 4439 81 4451 115
rect 4389 64 4451 81
rect 4806 111 4858 123
rect 4806 77 4814 111
rect 4848 77 4858 111
rect 4806 43 4858 77
rect 4806 9 4814 43
rect 4848 9 4858 43
rect 4806 -25 4858 9
rect 4806 -59 4814 -25
rect 4848 -59 4858 -25
rect 4806 -77 4858 -59
rect 4888 111 4940 123
rect 4888 77 4898 111
rect 4932 77 4940 111
rect 4888 43 4940 77
rect 4888 9 4898 43
rect 4932 9 4940 43
rect 4888 -25 4940 9
rect 4888 -59 4898 -25
rect 4932 -59 4940 -25
rect 4888 -77 4940 -59
<< ndiffc >>
rect -229 -317 -195 -283
rect -133 -317 -99 -283
rect -37 -317 -3 -283
rect 59 -317 93 -283
rect 155 -317 189 -283
rect 251 -317 285 -283
rect 347 -317 381 -283
rect 443 -317 477 -283
rect 539 -317 573 -283
rect 635 -317 669 -283
rect 731 -317 765 -283
rect 1924 -313 1958 -279
rect 2020 -313 2054 -279
rect 2116 -313 2150 -279
rect 2212 -313 2246 -279
rect 2308 -313 2342 -279
rect 2404 -313 2438 -279
rect 2500 -313 2534 -279
rect 2596 -313 2630 -279
rect 2692 -313 2726 -279
rect 2788 -313 2822 -279
rect 2884 -313 2918 -279
rect 3105 -328 3139 -252
rect 3193 -328 3227 -252
rect 3445 -313 3479 -279
rect 3541 -313 3575 -279
rect 3637 -313 3671 -279
rect 3733 -313 3767 -279
rect 3829 -313 3863 -279
rect 3925 -313 3959 -279
rect 4021 -313 4055 -279
rect 4117 -313 4151 -279
rect 4213 -313 4247 -279
rect 4309 -313 4343 -279
rect 4405 -313 4439 -279
rect 4814 -243 4848 -209
rect 4814 -311 4848 -277
rect 4898 -243 4932 -209
rect 4898 -311 4932 -277
<< pdiffc >>
rect -229 281 -195 315
rect -229 213 -195 247
rect -229 145 -195 179
rect -229 77 -195 111
rect -133 281 -99 315
rect -133 213 -99 247
rect -133 145 -99 179
rect -133 77 -99 111
rect -37 281 -3 315
rect -37 213 -3 247
rect -37 145 -3 179
rect -37 77 -3 111
rect 59 281 93 315
rect 59 213 93 247
rect 59 145 93 179
rect 59 77 93 111
rect 155 281 189 315
rect 155 213 189 247
rect 155 145 189 179
rect 155 77 189 111
rect 251 281 285 315
rect 251 213 285 247
rect 251 145 285 179
rect 251 77 285 111
rect 347 281 381 315
rect 347 213 381 247
rect 347 145 381 179
rect 347 77 381 111
rect 443 281 477 315
rect 443 213 477 247
rect 443 145 477 179
rect 443 77 477 111
rect 539 281 573 315
rect 539 213 573 247
rect 539 145 573 179
rect 539 77 573 111
rect 635 281 669 315
rect 635 213 669 247
rect 635 145 669 179
rect 635 77 669 111
rect 731 281 765 315
rect 731 213 765 247
rect 731 145 765 179
rect 731 77 765 111
rect 1924 285 1958 319
rect 1924 217 1958 251
rect 1924 149 1958 183
rect 1924 81 1958 115
rect 2020 285 2054 319
rect 2020 217 2054 251
rect 2020 149 2054 183
rect 2020 81 2054 115
rect 2116 285 2150 319
rect 2116 217 2150 251
rect 2116 149 2150 183
rect 2116 81 2150 115
rect 2212 285 2246 319
rect 2212 217 2246 251
rect 2212 149 2246 183
rect 2212 81 2246 115
rect 2308 285 2342 319
rect 2308 217 2342 251
rect 2308 149 2342 183
rect 2308 81 2342 115
rect 2404 285 2438 319
rect 2404 217 2438 251
rect 2404 149 2438 183
rect 2404 81 2438 115
rect 2500 285 2534 319
rect 2500 217 2534 251
rect 2500 149 2534 183
rect 2500 81 2534 115
rect 2596 285 2630 319
rect 2596 217 2630 251
rect 2596 149 2630 183
rect 2596 81 2630 115
rect 2692 285 2726 319
rect 2692 217 2726 251
rect 2692 149 2726 183
rect 2692 81 2726 115
rect 2788 285 2822 319
rect 2788 217 2822 251
rect 2788 149 2822 183
rect 2788 81 2822 115
rect 2884 285 2918 319
rect 2884 217 2918 251
rect 2884 149 2918 183
rect 2884 81 2918 115
rect 3445 285 3479 319
rect 3445 217 3479 251
rect 3445 149 3479 183
rect 3445 81 3479 115
rect 3541 285 3575 319
rect 3541 217 3575 251
rect 3541 149 3575 183
rect 3541 81 3575 115
rect 3637 285 3671 319
rect 3637 217 3671 251
rect 3637 149 3671 183
rect 3637 81 3671 115
rect 3733 285 3767 319
rect 3733 217 3767 251
rect 3733 149 3767 183
rect 3733 81 3767 115
rect 3829 285 3863 319
rect 3829 217 3863 251
rect 3829 149 3863 183
rect 3829 81 3863 115
rect 3925 285 3959 319
rect 3925 217 3959 251
rect 3925 149 3959 183
rect 3925 81 3959 115
rect 4021 285 4055 319
rect 4021 217 4055 251
rect 4021 149 4055 183
rect 4021 81 4055 115
rect 4117 285 4151 319
rect 4117 217 4151 251
rect 4117 149 4151 183
rect 4117 81 4151 115
rect 4213 285 4247 319
rect 4213 217 4247 251
rect 4213 149 4247 183
rect 4213 81 4247 115
rect 4309 285 4343 319
rect 4309 217 4343 251
rect 4309 149 4343 183
rect 4309 81 4343 115
rect 4405 285 4439 319
rect 4405 217 4439 251
rect 4405 149 4439 183
rect 4405 81 4439 115
rect 4814 77 4848 111
rect 4814 9 4848 43
rect 4814 -59 4848 -25
rect 4898 77 4932 111
rect 4898 9 4932 43
rect 4898 -59 4932 -25
<< psubdiff >>
rect -343 -170 -225 -136
rect -191 -170 -157 -136
rect -123 -170 -89 -136
rect -55 -170 -21 -136
rect 13 -170 47 -136
rect 81 -170 115 -136
rect 149 -170 183 -136
rect 217 -170 251 -136
rect 285 -170 319 -136
rect 353 -170 387 -136
rect 421 -170 455 -136
rect 489 -170 523 -136
rect 557 -170 591 -136
rect 625 -170 659 -136
rect 693 -170 727 -136
rect 761 -170 879 -136
rect -343 -246 -309 -170
rect 845 -246 879 -170
rect -343 -314 -309 -280
rect -343 -382 -309 -348
rect 845 -314 879 -280
rect -343 -492 -309 -416
rect 845 -382 879 -348
rect 845 -492 879 -416
rect -343 -526 -225 -492
rect -191 -526 -157 -492
rect -123 -526 -89 -492
rect -55 -526 -21 -492
rect 13 -526 47 -492
rect 81 -526 115 -492
rect 149 -526 183 -492
rect 217 -526 251 -492
rect 285 -526 319 -492
rect 353 -526 387 -492
rect 421 -526 455 -492
rect 489 -526 523 -492
rect 557 -526 591 -492
rect 625 -526 659 -492
rect 693 -526 727 -492
rect 761 -526 879 -492
rect 1810 -166 1928 -132
rect 1962 -166 1996 -132
rect 2030 -166 2064 -132
rect 2098 -166 2132 -132
rect 2166 -166 2200 -132
rect 2234 -166 2268 -132
rect 2302 -166 2336 -132
rect 2370 -166 2404 -132
rect 2438 -166 2472 -132
rect 2506 -166 2540 -132
rect 2574 -166 2608 -132
rect 2642 -166 2676 -132
rect 2710 -166 2744 -132
rect 2778 -166 2812 -132
rect 2846 -166 2880 -132
rect 2914 -166 3032 -132
rect 1810 -242 1844 -166
rect 2998 -242 3032 -166
rect 3331 -166 3449 -132
rect 3483 -166 3517 -132
rect 3551 -166 3585 -132
rect 3619 -166 3653 -132
rect 3687 -166 3721 -132
rect 3755 -166 3789 -132
rect 3823 -166 3857 -132
rect 3891 -166 3925 -132
rect 3959 -166 3993 -132
rect 4027 -166 4061 -132
rect 4095 -166 4129 -132
rect 4163 -166 4197 -132
rect 4231 -166 4265 -132
rect 4299 -166 4333 -132
rect 4367 -166 4401 -132
rect 4435 -166 4553 -132
rect 1810 -310 1844 -276
rect 1810 -378 1844 -344
rect 2998 -310 3032 -276
rect 3331 -242 3365 -166
rect 4519 -242 4553 -166
rect 3331 -310 3365 -276
rect 1810 -488 1844 -412
rect 2998 -378 3032 -344
rect 2998 -488 3032 -412
rect 1810 -522 1928 -488
rect 1962 -522 1996 -488
rect 2030 -522 2064 -488
rect 2098 -522 2132 -488
rect 2166 -522 2200 -488
rect 2234 -522 2268 -488
rect 2302 -522 2336 -488
rect 2370 -522 2404 -488
rect 2438 -522 2472 -488
rect 2506 -522 2540 -488
rect 2574 -522 2608 -488
rect 2642 -522 2676 -488
rect 2710 -522 2744 -488
rect 2778 -522 2812 -488
rect 2846 -522 2880 -488
rect 2914 -522 3032 -488
rect 3331 -378 3365 -344
rect 4519 -310 4553 -276
rect 3331 -488 3365 -412
rect 4519 -378 4553 -344
rect 4519 -488 4553 -412
rect 3331 -522 3449 -488
rect 3483 -522 3517 -488
rect 3551 -522 3585 -488
rect 3619 -522 3653 -488
rect 3687 -522 3721 -488
rect 3755 -522 3789 -488
rect 3823 -522 3857 -488
rect 3891 -522 3925 -488
rect 3959 -522 3993 -488
rect 4027 -522 4061 -488
rect 4095 -522 4129 -488
rect 4163 -522 4197 -488
rect 4231 -522 4265 -488
rect 4299 -522 4333 -488
rect 4367 -522 4401 -488
rect 4435 -522 4553 -488
<< nsubdiff >>
rect -343 482 -225 516
rect -191 482 -157 516
rect -123 482 -89 516
rect -55 482 -21 516
rect 13 482 47 516
rect 81 482 115 516
rect 149 482 183 516
rect 217 482 251 516
rect 285 482 319 516
rect 353 482 387 516
rect 421 482 455 516
rect 489 482 523 516
rect 557 482 591 516
rect 625 482 659 516
rect 693 482 727 516
rect 761 482 879 516
rect -343 414 -309 482
rect -343 346 -309 380
rect 845 414 879 482
rect 845 346 879 380
rect -343 278 -309 312
rect -343 210 -309 244
rect -343 142 -309 176
rect -343 74 -309 108
rect 845 278 879 312
rect 845 210 879 244
rect 845 142 879 176
rect 845 74 879 108
rect -343 -28 -309 40
rect 845 -28 879 40
rect -343 -62 -225 -28
rect -191 -62 -157 -28
rect -123 -62 -89 -28
rect -55 -62 -21 -28
rect 13 -62 47 -28
rect 81 -62 115 -28
rect 149 -62 183 -28
rect 217 -62 251 -28
rect 285 -62 319 -28
rect 353 -62 387 -28
rect 421 -62 455 -28
rect 489 -62 523 -28
rect 557 -62 591 -28
rect 625 -62 659 -28
rect 693 -62 727 -28
rect 761 -62 879 -28
rect 1810 486 1928 520
rect 1962 486 1996 520
rect 2030 486 2064 520
rect 2098 486 2132 520
rect 2166 486 2200 520
rect 2234 486 2268 520
rect 2302 486 2336 520
rect 2370 486 2404 520
rect 2438 486 2472 520
rect 2506 486 2540 520
rect 2574 486 2608 520
rect 2642 486 2676 520
rect 2710 486 2744 520
rect 2778 486 2812 520
rect 2846 486 2880 520
rect 2914 486 3032 520
rect 1810 418 1844 486
rect 1810 350 1844 384
rect 2998 418 3032 486
rect 2998 350 3032 384
rect 1810 282 1844 316
rect 1810 214 1844 248
rect 1810 146 1844 180
rect 1810 78 1844 112
rect 2998 282 3032 316
rect 2998 214 3032 248
rect 2998 146 3032 180
rect 2998 78 3032 112
rect 1810 -24 1844 44
rect 2998 -24 3032 44
rect 1810 -58 1928 -24
rect 1962 -58 1996 -24
rect 2030 -58 2064 -24
rect 2098 -58 2132 -24
rect 2166 -58 2200 -24
rect 2234 -58 2268 -24
rect 2302 -58 2336 -24
rect 2370 -58 2404 -24
rect 2438 -58 2472 -24
rect 2506 -58 2540 -24
rect 2574 -58 2608 -24
rect 2642 -58 2676 -24
rect 2710 -58 2744 -24
rect 2778 -58 2812 -24
rect 2846 -58 2880 -24
rect 2914 -58 3032 -24
rect 3331 486 3449 520
rect 3483 486 3517 520
rect 3551 486 3585 520
rect 3619 486 3653 520
rect 3687 486 3721 520
rect 3755 486 3789 520
rect 3823 486 3857 520
rect 3891 486 3925 520
rect 3959 486 3993 520
rect 4027 486 4061 520
rect 4095 486 4129 520
rect 4163 486 4197 520
rect 4231 486 4265 520
rect 4299 486 4333 520
rect 4367 486 4401 520
rect 4435 486 4553 520
rect 3331 418 3365 486
rect 3331 350 3365 384
rect 4519 418 4553 486
rect 4519 350 4553 384
rect 3331 282 3365 316
rect 3331 214 3365 248
rect 3331 146 3365 180
rect 3331 78 3365 112
rect 4519 282 4553 316
rect 4519 214 4553 248
rect 4519 146 4553 180
rect 4519 78 4553 112
rect 3331 -24 3365 44
rect 4519 -24 4553 44
rect 3331 -58 3449 -24
rect 3483 -58 3517 -24
rect 3551 -58 3585 -24
rect 3619 -58 3653 -24
rect 3687 -58 3721 -24
rect 3755 -58 3789 -24
rect 3823 -58 3857 -24
rect 3891 -58 3925 -24
rect 3959 -58 3993 -24
rect 4027 -58 4061 -24
rect 4095 -58 4129 -24
rect 4163 -58 4197 -24
rect 4231 -58 4265 -24
rect 4299 -58 4333 -24
rect 4367 -58 4401 -24
rect 4435 -58 4553 -24
<< psubdiffcont >>
rect -225 -170 -191 -136
rect -157 -170 -123 -136
rect -89 -170 -55 -136
rect -21 -170 13 -136
rect 47 -170 81 -136
rect 115 -170 149 -136
rect 183 -170 217 -136
rect 251 -170 285 -136
rect 319 -170 353 -136
rect 387 -170 421 -136
rect 455 -170 489 -136
rect 523 -170 557 -136
rect 591 -170 625 -136
rect 659 -170 693 -136
rect 727 -170 761 -136
rect -343 -280 -309 -246
rect -343 -348 -309 -314
rect 845 -280 879 -246
rect 845 -348 879 -314
rect -343 -416 -309 -382
rect 845 -416 879 -382
rect -225 -526 -191 -492
rect -157 -526 -123 -492
rect -89 -526 -55 -492
rect -21 -526 13 -492
rect 47 -526 81 -492
rect 115 -526 149 -492
rect 183 -526 217 -492
rect 251 -526 285 -492
rect 319 -526 353 -492
rect 387 -526 421 -492
rect 455 -526 489 -492
rect 523 -526 557 -492
rect 591 -526 625 -492
rect 659 -526 693 -492
rect 727 -526 761 -492
rect 1928 -166 1962 -132
rect 1996 -166 2030 -132
rect 2064 -166 2098 -132
rect 2132 -166 2166 -132
rect 2200 -166 2234 -132
rect 2268 -166 2302 -132
rect 2336 -166 2370 -132
rect 2404 -166 2438 -132
rect 2472 -166 2506 -132
rect 2540 -166 2574 -132
rect 2608 -166 2642 -132
rect 2676 -166 2710 -132
rect 2744 -166 2778 -132
rect 2812 -166 2846 -132
rect 2880 -166 2914 -132
rect 1810 -276 1844 -242
rect 3449 -166 3483 -132
rect 3517 -166 3551 -132
rect 3585 -166 3619 -132
rect 3653 -166 3687 -132
rect 3721 -166 3755 -132
rect 3789 -166 3823 -132
rect 3857 -166 3891 -132
rect 3925 -166 3959 -132
rect 3993 -166 4027 -132
rect 4061 -166 4095 -132
rect 4129 -166 4163 -132
rect 4197 -166 4231 -132
rect 4265 -166 4299 -132
rect 4333 -166 4367 -132
rect 4401 -166 4435 -132
rect 1810 -344 1844 -310
rect 2998 -276 3032 -242
rect 2998 -344 3032 -310
rect 3331 -276 3365 -242
rect 1810 -412 1844 -378
rect 3331 -344 3365 -310
rect 2998 -412 3032 -378
rect 1928 -522 1962 -488
rect 1996 -522 2030 -488
rect 2064 -522 2098 -488
rect 2132 -522 2166 -488
rect 2200 -522 2234 -488
rect 2268 -522 2302 -488
rect 2336 -522 2370 -488
rect 2404 -522 2438 -488
rect 2472 -522 2506 -488
rect 2540 -522 2574 -488
rect 2608 -522 2642 -488
rect 2676 -522 2710 -488
rect 2744 -522 2778 -488
rect 2812 -522 2846 -488
rect 2880 -522 2914 -488
rect 4519 -276 4553 -242
rect 4519 -344 4553 -310
rect 3331 -412 3365 -378
rect 4519 -412 4553 -378
rect 3449 -522 3483 -488
rect 3517 -522 3551 -488
rect 3585 -522 3619 -488
rect 3653 -522 3687 -488
rect 3721 -522 3755 -488
rect 3789 -522 3823 -488
rect 3857 -522 3891 -488
rect 3925 -522 3959 -488
rect 3993 -522 4027 -488
rect 4061 -522 4095 -488
rect 4129 -522 4163 -488
rect 4197 -522 4231 -488
rect 4265 -522 4299 -488
rect 4333 -522 4367 -488
rect 4401 -522 4435 -488
<< nsubdiffcont >>
rect -225 482 -191 516
rect -157 482 -123 516
rect -89 482 -55 516
rect -21 482 13 516
rect 47 482 81 516
rect 115 482 149 516
rect 183 482 217 516
rect 251 482 285 516
rect 319 482 353 516
rect 387 482 421 516
rect 455 482 489 516
rect 523 482 557 516
rect 591 482 625 516
rect 659 482 693 516
rect 727 482 761 516
rect -343 380 -309 414
rect 845 380 879 414
rect -343 312 -309 346
rect -343 244 -309 278
rect -343 176 -309 210
rect -343 108 -309 142
rect -343 40 -309 74
rect 845 312 879 346
rect 845 244 879 278
rect 845 176 879 210
rect 845 108 879 142
rect 845 40 879 74
rect -225 -62 -191 -28
rect -157 -62 -123 -28
rect -89 -62 -55 -28
rect -21 -62 13 -28
rect 47 -62 81 -28
rect 115 -62 149 -28
rect 183 -62 217 -28
rect 251 -62 285 -28
rect 319 -62 353 -28
rect 387 -62 421 -28
rect 455 -62 489 -28
rect 523 -62 557 -28
rect 591 -62 625 -28
rect 659 -62 693 -28
rect 727 -62 761 -28
rect 1928 486 1962 520
rect 1996 486 2030 520
rect 2064 486 2098 520
rect 2132 486 2166 520
rect 2200 486 2234 520
rect 2268 486 2302 520
rect 2336 486 2370 520
rect 2404 486 2438 520
rect 2472 486 2506 520
rect 2540 486 2574 520
rect 2608 486 2642 520
rect 2676 486 2710 520
rect 2744 486 2778 520
rect 2812 486 2846 520
rect 2880 486 2914 520
rect 1810 384 1844 418
rect 2998 384 3032 418
rect 1810 316 1844 350
rect 1810 248 1844 282
rect 1810 180 1844 214
rect 1810 112 1844 146
rect 1810 44 1844 78
rect 2998 316 3032 350
rect 2998 248 3032 282
rect 2998 180 3032 214
rect 2998 112 3032 146
rect 2998 44 3032 78
rect 1928 -58 1962 -24
rect 1996 -58 2030 -24
rect 2064 -58 2098 -24
rect 2132 -58 2166 -24
rect 2200 -58 2234 -24
rect 2268 -58 2302 -24
rect 2336 -58 2370 -24
rect 2404 -58 2438 -24
rect 2472 -58 2506 -24
rect 2540 -58 2574 -24
rect 2608 -58 2642 -24
rect 2676 -58 2710 -24
rect 2744 -58 2778 -24
rect 2812 -58 2846 -24
rect 2880 -58 2914 -24
rect 3449 486 3483 520
rect 3517 486 3551 520
rect 3585 486 3619 520
rect 3653 486 3687 520
rect 3721 486 3755 520
rect 3789 486 3823 520
rect 3857 486 3891 520
rect 3925 486 3959 520
rect 3993 486 4027 520
rect 4061 486 4095 520
rect 4129 486 4163 520
rect 4197 486 4231 520
rect 4265 486 4299 520
rect 4333 486 4367 520
rect 4401 486 4435 520
rect 3331 384 3365 418
rect 4519 384 4553 418
rect 3331 316 3365 350
rect 3331 248 3365 282
rect 3331 180 3365 214
rect 3331 112 3365 146
rect 3331 44 3365 78
rect 4519 316 4553 350
rect 4519 248 4553 282
rect 4519 180 4553 214
rect 4519 112 4553 146
rect 4519 44 4553 78
rect 3449 -58 3483 -24
rect 3517 -58 3551 -24
rect 3585 -58 3619 -24
rect 3653 -58 3687 -24
rect 3721 -58 3755 -24
rect 3789 -58 3823 -24
rect 3857 -58 3891 -24
rect 3925 -58 3959 -24
rect 3993 -58 4027 -24
rect 4061 -58 4095 -24
rect 4129 -58 4163 -24
rect 4197 -58 4231 -24
rect 4265 -58 4299 -24
rect 4333 -58 4367 -24
rect 4401 -58 4435 -24
<< poly >>
rect -245 414 781 430
rect -245 380 -229 414
rect -195 380 -37 414
rect -3 380 155 414
rect 189 380 347 414
rect 381 380 539 414
rect 573 380 731 414
rect 765 380 781 414
rect -245 364 781 380
rect -179 332 -149 364
rect -83 332 -53 364
rect 13 332 43 364
rect 109 332 139 364
rect 205 332 235 364
rect 301 332 331 364
rect 397 332 427 364
rect 493 332 523 364
rect 589 332 619 364
rect 685 332 715 364
rect -179 34 -149 60
rect -83 34 -53 60
rect 13 34 43 60
rect 109 34 139 60
rect 205 34 235 60
rect 301 34 331 60
rect 397 34 427 60
rect 493 34 523 60
rect 589 34 619 60
rect 685 34 715 60
rect 1908 418 2934 434
rect 1908 384 1924 418
rect 1958 384 2116 418
rect 2150 384 2308 418
rect 2342 384 2500 418
rect 2534 384 2692 418
rect 2726 384 2884 418
rect 2918 384 2934 418
rect 1908 368 2934 384
rect 1974 336 2004 368
rect 2070 336 2100 368
rect 2166 336 2196 368
rect 2262 336 2292 368
rect 2358 336 2388 368
rect 2454 336 2484 368
rect 2550 336 2580 368
rect 2646 336 2676 368
rect 2742 336 2772 368
rect 2838 336 2868 368
rect 1974 38 2004 64
rect 2070 38 2100 64
rect 2166 38 2196 64
rect 2262 38 2292 64
rect 2358 38 2388 64
rect 2454 38 2484 64
rect 2550 38 2580 64
rect 2646 38 2676 64
rect 2742 38 2772 64
rect 2838 38 2868 64
rect 3429 418 4455 434
rect 3429 384 3445 418
rect 3479 384 3637 418
rect 3671 384 3829 418
rect 3863 384 4021 418
rect 4055 384 4213 418
rect 4247 384 4405 418
rect 4439 384 4455 418
rect 3429 368 4455 384
rect 3495 336 3525 368
rect 3591 336 3621 368
rect 3687 336 3717 368
rect 3783 336 3813 368
rect 3879 336 3909 368
rect 3975 336 4005 368
rect 4071 336 4101 368
rect 4167 336 4197 368
rect 4263 336 4293 368
rect 4359 336 4389 368
rect 4858 123 4888 149
rect 3495 38 3525 64
rect 3591 38 3621 64
rect 3687 38 3717 64
rect 3783 38 3813 64
rect 3879 38 3909 64
rect 3975 38 4005 64
rect 4071 38 4101 64
rect 4167 38 4197 64
rect 4263 38 4293 64
rect 4359 38 4389 64
rect 4858 -109 4888 -77
rect 4858 -125 4944 -109
rect -179 -248 -149 -222
rect -83 -248 -53 -222
rect 13 -248 43 -222
rect 109 -248 139 -222
rect 205 -248 235 -222
rect 301 -248 331 -222
rect 397 -248 427 -222
rect 493 -248 523 -222
rect 589 -248 619 -222
rect 685 -248 715 -222
rect -179 -374 -149 -352
rect -83 -374 -53 -352
rect 13 -374 43 -352
rect 109 -374 139 -352
rect 205 -374 235 -352
rect 301 -374 331 -352
rect 397 -374 427 -352
rect 493 -374 523 -352
rect 589 -374 619 -352
rect 685 -374 715 -352
rect -245 -394 781 -374
rect -245 -428 -229 -394
rect -195 -428 -37 -394
rect -3 -428 155 -394
rect 189 -428 347 -394
rect 381 -428 539 -394
rect 573 -428 731 -394
rect 765 -428 781 -394
rect -245 -440 781 -428
rect 1974 -244 2004 -218
rect 2070 -244 2100 -218
rect 2166 -244 2196 -218
rect 2262 -244 2292 -218
rect 2358 -244 2388 -218
rect 2454 -244 2484 -218
rect 2550 -244 2580 -218
rect 2646 -244 2676 -218
rect 2742 -244 2772 -218
rect 2838 -244 2868 -218
rect 3133 -168 3199 -152
rect 3133 -202 3149 -168
rect 3183 -202 3199 -168
rect 3133 -218 3199 -202
rect 3151 -240 3181 -218
rect 3495 -244 3525 -218
rect 3591 -244 3621 -218
rect 3687 -244 3717 -218
rect 3783 -244 3813 -218
rect 3879 -244 3909 -218
rect 3975 -244 4005 -218
rect 4071 -244 4101 -218
rect 4167 -244 4197 -218
rect 4263 -244 4293 -218
rect 4359 -244 4389 -218
rect 4858 -159 4894 -125
rect 4928 -159 4944 -125
rect 4858 -175 4944 -159
rect 4858 -197 4888 -175
rect 1974 -370 2004 -348
rect 2070 -370 2100 -348
rect 2166 -370 2196 -348
rect 2262 -370 2292 -348
rect 2358 -370 2388 -348
rect 2454 -370 2484 -348
rect 2550 -370 2580 -348
rect 2646 -370 2676 -348
rect 2742 -370 2772 -348
rect 2838 -370 2868 -348
rect 1908 -390 2934 -370
rect 1908 -424 1924 -390
rect 1958 -424 2116 -390
rect 2150 -424 2308 -390
rect 2342 -424 2500 -390
rect 2534 -424 2692 -390
rect 2726 -424 2884 -390
rect 2918 -424 2934 -390
rect 1908 -436 2934 -424
rect 3151 -366 3181 -340
rect 3495 -370 3525 -348
rect 3591 -370 3621 -348
rect 3687 -370 3717 -348
rect 3783 -370 3813 -348
rect 3879 -370 3909 -348
rect 3975 -370 4005 -348
rect 4071 -370 4101 -348
rect 4167 -370 4197 -348
rect 4263 -370 4293 -348
rect 4359 -370 4389 -348
rect 3429 -390 4455 -370
rect 3429 -424 3445 -390
rect 3479 -424 3637 -390
rect 3671 -424 3829 -390
rect 3863 -424 4021 -390
rect 4055 -424 4213 -390
rect 4247 -424 4405 -390
rect 4439 -424 4455 -390
rect 3429 -436 4455 -424
rect 4858 -353 4888 -327
<< polycont >>
rect -229 380 -195 414
rect -37 380 -3 414
rect 155 380 189 414
rect 347 380 381 414
rect 539 380 573 414
rect 731 380 765 414
rect 1924 384 1958 418
rect 2116 384 2150 418
rect 2308 384 2342 418
rect 2500 384 2534 418
rect 2692 384 2726 418
rect 2884 384 2918 418
rect 3445 384 3479 418
rect 3637 384 3671 418
rect 3829 384 3863 418
rect 4021 384 4055 418
rect 4213 384 4247 418
rect 4405 384 4439 418
rect -229 -428 -195 -394
rect -37 -428 -3 -394
rect 155 -428 189 -394
rect 347 -428 381 -394
rect 539 -428 573 -394
rect 731 -428 765 -394
rect 3149 -202 3183 -168
rect 4894 -159 4928 -125
rect 1924 -424 1958 -390
rect 2116 -424 2150 -390
rect 2308 -424 2342 -390
rect 2500 -424 2534 -390
rect 2692 -424 2726 -390
rect 2884 -424 2918 -390
rect 3445 -424 3479 -390
rect 3637 -424 3671 -390
rect 3829 -424 3863 -390
rect 4021 -424 4055 -390
rect 4213 -424 4247 -390
rect 4405 -424 4439 -390
<< locali >>
rect -343 482 -225 516
rect -191 482 -157 516
rect -123 482 -89 516
rect -55 482 -21 516
rect 13 482 47 516
rect 81 482 115 516
rect 149 482 183 516
rect 217 482 251 516
rect 285 482 319 516
rect 353 482 387 516
rect 421 482 455 516
rect 489 482 523 516
rect 557 482 591 516
rect 625 482 659 516
rect 693 482 727 516
rect 761 482 879 516
rect -343 414 -309 482
rect 845 414 879 482
rect -245 380 -229 414
rect -195 380 -179 414
rect -53 380 -37 414
rect -3 380 13 414
rect 139 380 155 414
rect 189 380 205 414
rect 331 380 347 414
rect 381 380 397 414
rect 523 380 539 414
rect 573 380 589 414
rect 715 380 731 414
rect 765 380 781 414
rect -343 346 -309 380
rect 845 346 879 354
rect -343 278 -309 312
rect -343 210 -309 244
rect -343 142 -309 176
rect -343 74 -309 108
rect -229 315 -195 336
rect -229 247 -195 251
rect -229 141 -195 145
rect -229 56 -195 77
rect -133 315 -99 336
rect -133 247 -99 251
rect -133 141 -99 145
rect -133 56 -99 77
rect -37 315 -3 336
rect -37 247 -3 251
rect -37 141 -3 145
rect -37 56 -3 77
rect 59 315 93 336
rect 59 247 93 251
rect 59 141 93 145
rect 59 56 93 77
rect 155 315 189 336
rect 155 247 189 251
rect 155 141 189 145
rect 155 56 189 77
rect 251 315 285 336
rect 251 247 285 251
rect 251 141 285 145
rect 251 56 285 77
rect 347 315 381 336
rect 347 247 381 251
rect 347 141 381 145
rect 347 56 381 77
rect 443 315 477 336
rect 443 247 477 251
rect 443 141 477 145
rect 443 56 477 77
rect 539 315 573 336
rect 539 247 573 251
rect 539 141 573 145
rect 539 56 573 77
rect 635 315 669 336
rect 635 247 669 251
rect 635 141 669 145
rect 635 56 669 77
rect 731 315 765 336
rect 731 247 765 251
rect 731 141 765 145
rect 731 56 765 77
rect 845 278 879 282
rect 845 172 879 176
rect 845 100 879 108
rect -343 -28 -309 40
rect 845 -28 879 40
rect -343 -62 -225 -28
rect -191 -62 -157 -28
rect -123 -62 -89 -28
rect -55 -62 -21 -28
rect 13 -62 47 -28
rect 81 -62 115 -28
rect 149 -62 183 -28
rect 217 -62 251 -28
rect 285 -62 319 -28
rect 353 -62 387 -28
rect 421 -62 455 -28
rect 489 -62 523 -28
rect 557 -62 591 -28
rect 625 -62 659 -28
rect 693 -62 727 -28
rect 761 -62 879 -28
rect 1810 486 1928 520
rect 1962 486 1996 520
rect 2030 486 2064 520
rect 2098 486 2132 520
rect 2166 486 2200 520
rect 2234 486 2268 520
rect 2302 486 2336 520
rect 2370 486 2404 520
rect 2438 486 2472 520
rect 2506 486 2540 520
rect 2574 486 2608 520
rect 2642 486 2676 520
rect 2710 486 2744 520
rect 2778 486 2812 520
rect 2846 486 2880 520
rect 2914 486 3032 520
rect 1810 418 1844 486
rect 2998 418 3032 486
rect 1908 384 1924 418
rect 1958 384 1974 418
rect 2100 384 2116 418
rect 2150 384 2166 418
rect 2292 384 2308 418
rect 2342 384 2358 418
rect 2484 384 2500 418
rect 2534 384 2550 418
rect 2676 384 2692 418
rect 2726 384 2742 418
rect 2868 384 2884 418
rect 2918 384 2934 418
rect 1810 350 1844 384
rect 2998 350 3032 358
rect 1810 282 1844 316
rect 1810 214 1844 248
rect 1810 146 1844 180
rect 1810 78 1844 112
rect 1924 319 1958 340
rect 1924 251 1958 255
rect 1924 145 1958 149
rect 1924 60 1958 81
rect 2020 319 2054 340
rect 2020 251 2054 255
rect 2020 145 2054 149
rect 2020 60 2054 81
rect 2116 319 2150 340
rect 2116 251 2150 255
rect 2116 145 2150 149
rect 2116 60 2150 81
rect 2212 319 2246 340
rect 2212 251 2246 255
rect 2212 145 2246 149
rect 2212 60 2246 81
rect 2308 319 2342 340
rect 2308 251 2342 255
rect 2308 145 2342 149
rect 2308 60 2342 81
rect 2404 319 2438 340
rect 2404 251 2438 255
rect 2404 145 2438 149
rect 2404 60 2438 81
rect 2500 319 2534 340
rect 2500 251 2534 255
rect 2500 145 2534 149
rect 2500 60 2534 81
rect 2596 319 2630 340
rect 2596 251 2630 255
rect 2596 145 2630 149
rect 2596 60 2630 81
rect 2692 319 2726 340
rect 2692 251 2726 255
rect 2692 145 2726 149
rect 2692 60 2726 81
rect 2788 319 2822 340
rect 2788 251 2822 255
rect 2788 145 2822 149
rect 2788 60 2822 81
rect 2884 319 2918 340
rect 2884 251 2918 255
rect 2884 145 2918 149
rect 2884 60 2918 81
rect 2998 282 3032 286
rect 2998 176 3032 180
rect 2998 104 3032 112
rect 1810 -24 1844 44
rect 2998 -24 3032 44
rect 1810 -58 1928 -24
rect 1962 -58 1996 -24
rect 2030 -58 2064 -24
rect 2098 -58 2132 -24
rect 2166 -58 2200 -24
rect 2234 -58 2268 -24
rect 2302 -58 2336 -24
rect 2370 -58 2404 -24
rect 2438 -58 2472 -24
rect 2506 -58 2540 -24
rect 2574 -58 2608 -24
rect 2642 -58 2676 -24
rect 2710 -58 2744 -24
rect 2778 -58 2812 -24
rect 2846 -58 2880 -24
rect 2914 -58 3032 -24
rect 3331 486 3449 520
rect 3483 486 3517 520
rect 3551 486 3585 520
rect 3619 486 3653 520
rect 3687 486 3721 520
rect 3755 486 3789 520
rect 3823 486 3857 520
rect 3891 486 3925 520
rect 3959 486 3993 520
rect 4027 486 4061 520
rect 4095 486 4129 520
rect 4163 486 4197 520
rect 4231 486 4265 520
rect 4299 486 4333 520
rect 4367 486 4401 520
rect 4435 486 4553 520
rect 3331 418 3365 486
rect 4519 418 4553 486
rect 3429 384 3445 418
rect 3479 384 3495 418
rect 3621 384 3637 418
rect 3671 384 3687 418
rect 3813 384 3829 418
rect 3863 384 3879 418
rect 4005 384 4021 418
rect 4055 384 4071 418
rect 4197 384 4213 418
rect 4247 384 4263 418
rect 4389 384 4405 418
rect 4439 384 4455 418
rect 3331 350 3365 384
rect 4519 350 4553 358
rect 3331 282 3365 316
rect 3331 214 3365 248
rect 3331 146 3365 180
rect 3331 78 3365 112
rect 3445 319 3479 340
rect 3445 251 3479 255
rect 3445 145 3479 149
rect 3445 60 3479 81
rect 3541 319 3575 340
rect 3541 251 3575 255
rect 3541 145 3575 149
rect 3541 60 3575 81
rect 3637 319 3671 340
rect 3637 251 3671 255
rect 3637 145 3671 149
rect 3637 60 3671 81
rect 3733 319 3767 340
rect 3733 251 3767 255
rect 3733 145 3767 149
rect 3733 60 3767 81
rect 3829 319 3863 340
rect 3829 251 3863 255
rect 3829 145 3863 149
rect 3829 60 3863 81
rect 3925 319 3959 340
rect 3925 251 3959 255
rect 3925 145 3959 149
rect 3925 60 3959 81
rect 4021 319 4055 340
rect 4021 251 4055 255
rect 4021 145 4055 149
rect 4021 60 4055 81
rect 4117 319 4151 340
rect 4117 251 4151 255
rect 4117 145 4151 149
rect 4117 60 4151 81
rect 4213 319 4247 340
rect 4213 251 4247 255
rect 4213 145 4247 149
rect 4213 60 4247 81
rect 4309 319 4343 340
rect 4309 251 4343 255
rect 4309 145 4343 149
rect 4309 60 4343 81
rect 4405 319 4439 340
rect 4405 251 4439 255
rect 4405 145 4439 149
rect 4405 60 4439 81
rect 4519 282 4553 286
rect 4519 176 4553 180
rect 4732 153 4761 187
rect 4795 153 4853 187
rect 4887 153 4945 187
rect 4979 153 5008 187
rect 4519 104 4553 112
rect 3331 -24 3365 44
rect 4519 -24 4553 44
rect 3331 -58 3449 -24
rect 3483 -58 3517 -24
rect 3551 -58 3585 -24
rect 3619 -58 3653 -24
rect 3687 -58 3721 -24
rect 3755 -58 3789 -24
rect 3823 -58 3857 -24
rect 3891 -58 3925 -24
rect 3959 -58 3993 -24
rect 4027 -58 4061 -24
rect 4095 -58 4129 -24
rect 4163 -58 4197 -24
rect 4231 -58 4265 -24
rect 4299 -58 4333 -24
rect 4367 -58 4401 -24
rect 4435 -58 4553 -24
rect 4798 111 4864 119
rect 4798 77 4814 111
rect 4848 77 4864 111
rect 4798 43 4864 77
rect 4798 9 4814 43
rect 4848 9 4864 43
rect 4798 -25 4864 9
rect 4798 -59 4814 -25
rect 4848 -59 4864 -25
rect 4798 -77 4864 -59
rect 4898 111 4940 153
rect 4932 77 4940 111
rect 4898 43 4940 77
rect 4932 9 4940 43
rect 4898 -25 4940 9
rect 4932 -59 4940 -25
rect 4898 -75 4940 -59
rect 4798 -127 4844 -77
rect -343 -170 -225 -136
rect -191 -170 -157 -136
rect -123 -170 -89 -136
rect -55 -170 -21 -136
rect 13 -170 47 -136
rect 81 -170 115 -136
rect 149 -170 183 -136
rect 217 -170 251 -136
rect 285 -170 319 -136
rect 353 -170 387 -136
rect 421 -170 455 -136
rect 489 -170 523 -136
rect 557 -170 591 -136
rect 625 -170 659 -136
rect 693 -170 727 -136
rect 761 -170 879 -136
rect -343 -246 -309 -170
rect 845 -241 879 -170
rect -343 -314 -309 -280
rect -343 -382 -309 -348
rect -229 -283 -195 -244
rect -229 -356 -195 -317
rect -133 -283 -99 -244
rect -133 -356 -99 -317
rect -37 -283 -3 -244
rect -37 -356 -3 -317
rect 59 -283 93 -244
rect 59 -356 93 -317
rect 155 -283 189 -244
rect 155 -356 189 -317
rect 251 -283 285 -244
rect 251 -356 285 -317
rect 347 -283 381 -244
rect 347 -356 381 -317
rect 443 -283 477 -244
rect 443 -356 477 -317
rect 539 -283 573 -244
rect 539 -356 573 -317
rect 635 -283 669 -244
rect 635 -356 669 -317
rect 731 -283 765 -244
rect 731 -356 765 -317
rect 845 -313 879 -280
rect 845 -382 879 -348
rect -343 -492 -309 -416
rect -245 -428 -229 -394
rect -195 -428 -179 -394
rect -53 -428 -37 -394
rect -3 -428 13 -394
rect 139 -428 155 -394
rect 189 -428 205 -394
rect 331 -428 347 -394
rect 381 -428 397 -394
rect 523 -428 539 -394
rect 573 -428 589 -394
rect 715 -428 731 -394
rect 765 -428 781 -394
rect 845 -492 879 -419
rect -343 -526 -225 -492
rect -191 -526 -157 -492
rect -123 -526 -89 -492
rect -55 -526 -21 -492
rect 13 -526 47 -492
rect 81 -526 115 -492
rect 149 -526 183 -492
rect 217 -526 251 -492
rect 285 -526 319 -492
rect 353 -526 387 -492
rect 421 -526 455 -492
rect 489 -526 523 -492
rect 557 -526 591 -492
rect 625 -526 659 -492
rect 693 -526 727 -492
rect 761 -526 879 -492
rect 1810 -166 1928 -132
rect 1962 -166 1996 -132
rect 2030 -166 2064 -132
rect 2098 -166 2132 -132
rect 2166 -166 2200 -132
rect 2234 -166 2268 -132
rect 2302 -166 2336 -132
rect 2370 -166 2404 -132
rect 2438 -166 2472 -132
rect 2506 -166 2540 -132
rect 2574 -166 2608 -132
rect 2642 -166 2676 -132
rect 2710 -166 2744 -132
rect 2778 -166 2812 -132
rect 2846 -166 2880 -132
rect 2914 -166 3032 -132
rect 1810 -242 1844 -166
rect 2998 -237 3032 -166
rect 3331 -166 3449 -132
rect 3483 -166 3517 -132
rect 3551 -166 3585 -132
rect 3619 -166 3653 -132
rect 3687 -166 3721 -132
rect 3755 -166 3789 -132
rect 3823 -166 3857 -132
rect 3891 -166 3925 -132
rect 3959 -166 3993 -132
rect 4027 -166 4061 -132
rect 4095 -166 4129 -132
rect 4163 -166 4197 -132
rect 4231 -166 4265 -132
rect 4299 -166 4333 -132
rect 4367 -166 4401 -132
rect 4435 -166 4553 -132
rect 3133 -202 3149 -168
rect 3183 -202 3199 -168
rect 1810 -310 1844 -276
rect 1810 -378 1844 -344
rect 1924 -279 1958 -240
rect 1924 -352 1958 -313
rect 2020 -279 2054 -240
rect 2020 -352 2054 -313
rect 2116 -279 2150 -240
rect 2116 -352 2150 -313
rect 2212 -279 2246 -240
rect 2212 -352 2246 -313
rect 2308 -279 2342 -240
rect 2308 -352 2342 -313
rect 2404 -279 2438 -240
rect 2404 -352 2438 -313
rect 2500 -279 2534 -240
rect 2500 -352 2534 -313
rect 2596 -279 2630 -240
rect 2596 -352 2630 -313
rect 2692 -279 2726 -240
rect 2692 -352 2726 -313
rect 2788 -279 2822 -240
rect 2788 -352 2822 -313
rect 2884 -279 2918 -240
rect 2884 -352 2918 -313
rect 2998 -309 3032 -276
rect 3105 -252 3139 -236
rect 3105 -344 3139 -328
rect 3193 -252 3227 -236
rect 3193 -344 3227 -328
rect 3331 -242 3365 -166
rect 4519 -237 4553 -166
rect 3331 -310 3365 -276
rect 2998 -378 3032 -344
rect 1810 -488 1844 -412
rect 1908 -424 1924 -390
rect 1958 -424 1974 -390
rect 2100 -424 2116 -390
rect 2150 -424 2166 -390
rect 2292 -424 2308 -390
rect 2342 -424 2358 -390
rect 2484 -424 2500 -390
rect 2534 -424 2550 -390
rect 2676 -424 2692 -390
rect 2726 -424 2742 -390
rect 2868 -424 2884 -390
rect 2918 -424 2934 -390
rect 2998 -488 3032 -415
rect 1810 -522 1928 -488
rect 1962 -522 1996 -488
rect 2030 -522 2064 -488
rect 2098 -522 2132 -488
rect 2166 -522 2200 -488
rect 2234 -522 2268 -488
rect 2302 -522 2336 -488
rect 2370 -522 2404 -488
rect 2438 -522 2472 -488
rect 2506 -522 2540 -488
rect 2574 -522 2608 -488
rect 2642 -522 2676 -488
rect 2710 -522 2744 -488
rect 2778 -522 2812 -488
rect 2846 -522 2880 -488
rect 2914 -522 3032 -488
rect 3331 -378 3365 -344
rect 3445 -279 3479 -240
rect 3445 -352 3479 -313
rect 3541 -279 3575 -240
rect 3541 -352 3575 -313
rect 3637 -279 3671 -240
rect 3637 -352 3671 -313
rect 3733 -279 3767 -240
rect 3733 -352 3767 -313
rect 3829 -279 3863 -240
rect 3829 -352 3863 -313
rect 3925 -279 3959 -240
rect 3925 -352 3959 -313
rect 4021 -279 4055 -240
rect 4021 -352 4055 -313
rect 4117 -279 4151 -240
rect 4117 -352 4151 -313
rect 4213 -279 4247 -240
rect 4213 -352 4247 -313
rect 4309 -279 4343 -240
rect 4309 -352 4343 -313
rect 4405 -279 4439 -240
rect 4405 -352 4439 -313
rect 4519 -309 4553 -276
rect 4798 -161 4806 -127
rect 4840 -161 4844 -127
rect 4878 -122 4944 -111
rect 4878 -125 4908 -122
rect 4878 -159 4894 -125
rect 4942 -156 4944 -122
rect 4928 -159 4944 -156
rect 4798 -197 4844 -161
rect 4798 -209 4864 -197
rect 4798 -243 4814 -209
rect 4848 -243 4864 -209
rect 4798 -277 4864 -243
rect 4798 -311 4814 -277
rect 4848 -311 4864 -277
rect 4798 -323 4864 -311
rect 4898 -209 4944 -193
rect 4932 -243 4944 -209
rect 4898 -277 4944 -243
rect 4932 -311 4944 -277
rect 4519 -378 4553 -344
rect 4898 -357 4944 -311
rect 3331 -488 3365 -412
rect 3429 -424 3445 -390
rect 3479 -424 3495 -390
rect 3621 -424 3637 -390
rect 3671 -424 3687 -390
rect 3813 -424 3829 -390
rect 3863 -424 3879 -390
rect 4005 -424 4021 -390
rect 4055 -424 4071 -390
rect 4197 -424 4213 -390
rect 4247 -424 4263 -390
rect 4389 -424 4405 -390
rect 4439 -424 4455 -390
rect 4732 -391 4761 -357
rect 4795 -391 4853 -357
rect 4887 -391 4945 -357
rect 4979 -391 5008 -357
rect 4519 -488 4553 -415
rect 3331 -522 3449 -488
rect 3483 -522 3517 -488
rect 3551 -522 3585 -488
rect 3619 -522 3653 -488
rect 3687 -522 3721 -488
rect 3755 -522 3789 -488
rect 3823 -522 3857 -488
rect 3891 -522 3925 -488
rect 3959 -522 3993 -488
rect 4027 -522 4061 -488
rect 4095 -522 4129 -488
rect 4163 -522 4197 -488
rect 4231 -522 4265 -488
rect 4299 -522 4333 -488
rect 4367 -522 4401 -488
rect 4435 -522 4553 -488
<< viali >>
rect -229 380 -195 414
rect -37 380 -3 414
rect 155 380 189 414
rect 347 380 381 414
rect 539 380 573 414
rect 731 380 765 414
rect 845 380 879 388
rect 845 354 879 380
rect -229 281 -195 285
rect -229 251 -195 281
rect -229 179 -195 213
rect -229 111 -195 141
rect -229 107 -195 111
rect -133 281 -99 285
rect -133 251 -99 281
rect -133 179 -99 213
rect -133 111 -99 141
rect -133 107 -99 111
rect -37 281 -3 285
rect -37 251 -3 281
rect -37 179 -3 213
rect -37 111 -3 141
rect -37 107 -3 111
rect 59 281 93 285
rect 59 251 93 281
rect 59 179 93 213
rect 59 111 93 141
rect 59 107 93 111
rect 155 281 189 285
rect 155 251 189 281
rect 155 179 189 213
rect 155 111 189 141
rect 155 107 189 111
rect 251 281 285 285
rect 251 251 285 281
rect 251 179 285 213
rect 251 111 285 141
rect 251 107 285 111
rect 347 281 381 285
rect 347 251 381 281
rect 347 179 381 213
rect 347 111 381 141
rect 347 107 381 111
rect 443 281 477 285
rect 443 251 477 281
rect 443 179 477 213
rect 443 111 477 141
rect 443 107 477 111
rect 539 281 573 285
rect 539 251 573 281
rect 539 179 573 213
rect 539 111 573 141
rect 539 107 573 111
rect 635 281 669 285
rect 635 251 669 281
rect 635 179 669 213
rect 635 111 669 141
rect 635 107 669 111
rect 731 281 765 285
rect 731 251 765 281
rect 731 179 765 213
rect 731 111 765 141
rect 731 107 765 111
rect 845 312 879 316
rect 845 282 879 312
rect 845 210 879 244
rect 845 142 879 172
rect 845 138 879 142
rect 845 74 879 100
rect 845 66 879 74
rect 1924 384 1958 418
rect 2116 384 2150 418
rect 2308 384 2342 418
rect 2500 384 2534 418
rect 2692 384 2726 418
rect 2884 384 2918 418
rect 2998 384 3032 392
rect 2998 358 3032 384
rect 1924 285 1958 289
rect 1924 255 1958 285
rect 1924 183 1958 217
rect 1924 115 1958 145
rect 1924 111 1958 115
rect 2020 285 2054 289
rect 2020 255 2054 285
rect 2020 183 2054 217
rect 2020 115 2054 145
rect 2020 111 2054 115
rect 2116 285 2150 289
rect 2116 255 2150 285
rect 2116 183 2150 217
rect 2116 115 2150 145
rect 2116 111 2150 115
rect 2212 285 2246 289
rect 2212 255 2246 285
rect 2212 183 2246 217
rect 2212 115 2246 145
rect 2212 111 2246 115
rect 2308 285 2342 289
rect 2308 255 2342 285
rect 2308 183 2342 217
rect 2308 115 2342 145
rect 2308 111 2342 115
rect 2404 285 2438 289
rect 2404 255 2438 285
rect 2404 183 2438 217
rect 2404 115 2438 145
rect 2404 111 2438 115
rect 2500 285 2534 289
rect 2500 255 2534 285
rect 2500 183 2534 217
rect 2500 115 2534 145
rect 2500 111 2534 115
rect 2596 285 2630 289
rect 2596 255 2630 285
rect 2596 183 2630 217
rect 2596 115 2630 145
rect 2596 111 2630 115
rect 2692 285 2726 289
rect 2692 255 2726 285
rect 2692 183 2726 217
rect 2692 115 2726 145
rect 2692 111 2726 115
rect 2788 285 2822 289
rect 2788 255 2822 285
rect 2788 183 2822 217
rect 2788 115 2822 145
rect 2788 111 2822 115
rect 2884 285 2918 289
rect 2884 255 2918 285
rect 2884 183 2918 217
rect 2884 115 2918 145
rect 2884 111 2918 115
rect 2998 316 3032 320
rect 2998 286 3032 316
rect 2998 214 3032 248
rect 2998 146 3032 176
rect 2998 142 3032 146
rect 2998 78 3032 104
rect 2998 70 3032 78
rect 3445 384 3479 418
rect 3637 384 3671 418
rect 3829 384 3863 418
rect 4021 384 4055 418
rect 4213 384 4247 418
rect 4405 384 4439 418
rect 4519 384 4553 392
rect 4519 358 4553 384
rect 3445 285 3479 289
rect 3445 255 3479 285
rect 3445 183 3479 217
rect 3445 115 3479 145
rect 3445 111 3479 115
rect 3541 285 3575 289
rect 3541 255 3575 285
rect 3541 183 3575 217
rect 3541 115 3575 145
rect 3541 111 3575 115
rect 3637 285 3671 289
rect 3637 255 3671 285
rect 3637 183 3671 217
rect 3637 115 3671 145
rect 3637 111 3671 115
rect 3733 285 3767 289
rect 3733 255 3767 285
rect 3733 183 3767 217
rect 3733 115 3767 145
rect 3733 111 3767 115
rect 3829 285 3863 289
rect 3829 255 3863 285
rect 3829 183 3863 217
rect 3829 115 3863 145
rect 3829 111 3863 115
rect 3925 285 3959 289
rect 3925 255 3959 285
rect 3925 183 3959 217
rect 3925 115 3959 145
rect 3925 111 3959 115
rect 4021 285 4055 289
rect 4021 255 4055 285
rect 4021 183 4055 217
rect 4021 115 4055 145
rect 4021 111 4055 115
rect 4117 285 4151 289
rect 4117 255 4151 285
rect 4117 183 4151 217
rect 4117 115 4151 145
rect 4117 111 4151 115
rect 4213 285 4247 289
rect 4213 255 4247 285
rect 4213 183 4247 217
rect 4213 115 4247 145
rect 4213 111 4247 115
rect 4309 285 4343 289
rect 4309 255 4343 285
rect 4309 183 4343 217
rect 4309 115 4343 145
rect 4309 111 4343 115
rect 4405 285 4439 289
rect 4405 255 4439 285
rect 4405 183 4439 217
rect 4405 115 4439 145
rect 4405 111 4439 115
rect 4519 316 4553 320
rect 4519 286 4553 316
rect 4519 214 4553 248
rect 4519 146 4553 176
rect 4761 153 4795 187
rect 4853 153 4887 187
rect 4945 153 4979 187
rect 4519 142 4553 146
rect 4519 78 4553 104
rect 4519 70 4553 78
rect -229 -317 -195 -283
rect -133 -317 -99 -283
rect -37 -317 -3 -283
rect 59 -317 93 -283
rect 155 -317 189 -283
rect 251 -317 285 -283
rect 347 -317 381 -283
rect 443 -317 477 -283
rect 539 -317 573 -283
rect 635 -317 669 -283
rect 731 -317 765 -283
rect 845 -246 879 -241
rect 845 -275 879 -246
rect 845 -314 879 -313
rect 845 -347 879 -314
rect -229 -428 -195 -394
rect -37 -428 -3 -394
rect 155 -428 189 -394
rect 347 -428 381 -394
rect 539 -428 573 -394
rect 731 -428 765 -394
rect 845 -416 879 -385
rect 845 -419 879 -416
rect 3149 -202 3183 -168
rect 1924 -313 1958 -279
rect 2020 -313 2054 -279
rect 2116 -313 2150 -279
rect 2212 -313 2246 -279
rect 2308 -313 2342 -279
rect 2404 -313 2438 -279
rect 2500 -313 2534 -279
rect 2596 -313 2630 -279
rect 2692 -313 2726 -279
rect 2788 -313 2822 -279
rect 2884 -313 2918 -279
rect 2998 -242 3032 -237
rect 2998 -271 3032 -242
rect 2998 -310 3032 -309
rect 2998 -343 3032 -310
rect 3105 -328 3139 -252
rect 3193 -328 3227 -252
rect 1924 -424 1958 -390
rect 2116 -424 2150 -390
rect 2308 -424 2342 -390
rect 2500 -424 2534 -390
rect 2692 -424 2726 -390
rect 2884 -424 2918 -390
rect 2998 -412 3032 -381
rect 2998 -415 3032 -412
rect 3445 -313 3479 -279
rect 3541 -313 3575 -279
rect 3637 -313 3671 -279
rect 3733 -313 3767 -279
rect 3829 -313 3863 -279
rect 3925 -313 3959 -279
rect 4021 -313 4055 -279
rect 4117 -313 4151 -279
rect 4213 -313 4247 -279
rect 4309 -313 4343 -279
rect 4405 -313 4439 -279
rect 4519 -242 4553 -237
rect 4519 -271 4553 -242
rect 4519 -310 4553 -309
rect 4519 -343 4553 -310
rect 4806 -161 4840 -127
rect 4908 -125 4942 -122
rect 4908 -156 4928 -125
rect 4928 -156 4942 -125
rect 3445 -424 3479 -390
rect 3637 -424 3671 -390
rect 3829 -424 3863 -390
rect 4021 -424 4055 -390
rect 4213 -424 4247 -390
rect 4405 -424 4439 -390
rect 4519 -412 4553 -381
rect 4761 -391 4795 -357
rect 4853 -391 4887 -357
rect 4945 -391 4979 -357
rect 4519 -415 4553 -412
<< metal1 >>
rect -413 482 669 516
rect -413 -81 -379 482
rect -248 372 -238 424
rect -186 372 -176 424
rect -133 332 -99 482
rect -55 372 -45 424
rect 7 372 17 424
rect 59 332 93 482
rect 136 372 146 424
rect 198 372 208 424
rect 251 332 285 482
rect 328 372 338 424
rect 390 372 400 424
rect 443 332 477 482
rect 520 372 530 424
rect 582 372 592 424
rect 635 332 669 482
rect 712 372 722 424
rect 774 372 784 424
rect 839 388 885 552
rect 1740 486 2822 520
rect 839 354 845 388
rect 879 354 885 388
rect 970 365 980 425
rect 1036 365 1250 425
rect 1310 365 1320 425
rect -235 285 -189 332
rect -235 251 -229 285
rect -195 251 -189 285
rect -235 213 -189 251
rect -235 179 -229 213
rect -195 179 -189 213
rect -235 141 -189 179
rect -235 107 -229 141
rect -195 107 -189 141
rect -235 60 -189 107
rect -139 285 -93 332
rect -139 251 -133 285
rect -99 251 -93 285
rect -139 213 -93 251
rect -139 179 -133 213
rect -99 179 -93 213
rect -139 141 -93 179
rect -139 107 -133 141
rect -99 107 -93 141
rect -139 60 -93 107
rect -43 285 3 332
rect -43 251 -37 285
rect -3 251 3 285
rect -43 213 3 251
rect -43 179 -37 213
rect -3 179 3 213
rect -43 141 3 179
rect -43 107 -37 141
rect -3 107 3 141
rect -43 60 3 107
rect 53 285 99 332
rect 53 251 59 285
rect 93 251 99 285
rect 53 213 99 251
rect 53 179 59 213
rect 93 179 99 213
rect 53 141 99 179
rect 53 107 59 141
rect 93 107 99 141
rect 53 60 99 107
rect 149 285 195 332
rect 149 251 155 285
rect 189 251 195 285
rect 149 213 195 251
rect 149 179 155 213
rect 189 179 195 213
rect 149 141 195 179
rect 149 107 155 141
rect 189 107 195 141
rect 149 60 195 107
rect 245 285 291 332
rect 245 251 251 285
rect 285 251 291 285
rect 245 213 291 251
rect 245 179 251 213
rect 285 179 291 213
rect 245 141 291 179
rect 245 107 251 141
rect 285 107 291 141
rect 245 60 291 107
rect 341 285 387 332
rect 341 251 347 285
rect 381 251 387 285
rect 341 213 387 251
rect 341 179 347 213
rect 381 179 387 213
rect 341 141 387 179
rect 341 107 347 141
rect 381 107 387 141
rect 341 60 387 107
rect 437 285 483 332
rect 437 251 443 285
rect 477 251 483 285
rect 437 213 483 251
rect 437 179 443 213
rect 477 179 483 213
rect 437 141 483 179
rect 437 107 443 141
rect 477 107 483 141
rect 437 60 483 107
rect 533 285 579 332
rect 533 251 539 285
rect 573 251 579 285
rect 533 213 579 251
rect 533 179 539 213
rect 573 179 579 213
rect 533 141 579 179
rect 533 107 539 141
rect 573 107 579 141
rect 533 60 579 107
rect 629 285 675 332
rect 629 251 635 285
rect 669 251 675 285
rect 629 213 675 251
rect 629 179 635 213
rect 669 179 675 213
rect 629 141 675 179
rect 629 107 635 141
rect 669 107 675 141
rect 629 60 675 107
rect 725 285 771 332
rect 725 251 731 285
rect 765 251 771 285
rect 725 213 771 251
rect 725 179 731 213
rect 765 179 771 213
rect 725 141 771 179
rect 725 107 731 141
rect 765 107 771 141
rect 725 60 771 107
rect 839 316 885 354
rect 839 282 845 316
rect 879 282 885 316
rect 839 244 885 282
rect 839 210 845 244
rect 879 210 885 244
rect 839 172 885 210
rect 839 138 845 172
rect 879 138 885 172
rect 839 100 885 138
rect 839 75 845 100
rect 838 66 845 75
rect 879 76 885 100
rect 879 66 1508 76
rect -542 -115 -379 -81
rect -413 -492 -379 -115
rect -229 -81 -195 60
rect -37 -81 -3 60
rect 155 -81 189 60
rect 347 -81 381 60
rect 539 -81 573 60
rect 731 -81 765 60
rect 838 16 1508 66
rect 1562 16 1572 76
rect 1740 -77 1774 486
rect 1905 376 1915 428
rect 1967 376 1977 428
rect 2020 336 2054 486
rect 2098 376 2108 428
rect 2160 376 2170 428
rect 2212 336 2246 486
rect 2289 376 2299 428
rect 2351 376 2361 428
rect 2404 336 2438 486
rect 2481 376 2491 428
rect 2543 376 2553 428
rect 2596 336 2630 486
rect 2673 376 2683 428
rect 2735 376 2745 428
rect 2788 336 2822 486
rect 2865 376 2875 428
rect 2927 376 2937 428
rect 2992 392 3038 600
rect 2992 358 2998 392
rect 3032 358 3038 392
rect 1918 289 1964 336
rect 1918 255 1924 289
rect 1958 255 1964 289
rect 1918 217 1964 255
rect 1918 183 1924 217
rect 1958 183 1964 217
rect 1918 145 1964 183
rect 1918 111 1924 145
rect 1958 111 1964 145
rect 1918 64 1964 111
rect 2014 289 2060 336
rect 2014 255 2020 289
rect 2054 255 2060 289
rect 2014 217 2060 255
rect 2014 183 2020 217
rect 2054 183 2060 217
rect 2014 145 2060 183
rect 2014 111 2020 145
rect 2054 111 2060 145
rect 2014 64 2060 111
rect 2110 289 2156 336
rect 2110 255 2116 289
rect 2150 255 2156 289
rect 2110 217 2156 255
rect 2110 183 2116 217
rect 2150 183 2156 217
rect 2110 145 2156 183
rect 2110 111 2116 145
rect 2150 111 2156 145
rect 2110 64 2156 111
rect 2206 289 2252 336
rect 2206 255 2212 289
rect 2246 255 2252 289
rect 2206 217 2252 255
rect 2206 183 2212 217
rect 2246 183 2252 217
rect 2206 145 2252 183
rect 2206 111 2212 145
rect 2246 111 2252 145
rect 2206 64 2252 111
rect 2302 289 2348 336
rect 2302 255 2308 289
rect 2342 255 2348 289
rect 2302 217 2348 255
rect 2302 183 2308 217
rect 2342 183 2348 217
rect 2302 145 2348 183
rect 2302 111 2308 145
rect 2342 111 2348 145
rect 2302 64 2348 111
rect 2398 289 2444 336
rect 2398 255 2404 289
rect 2438 255 2444 289
rect 2398 217 2444 255
rect 2398 183 2404 217
rect 2438 183 2444 217
rect 2398 145 2444 183
rect 2398 111 2404 145
rect 2438 111 2444 145
rect 2398 64 2444 111
rect 2494 289 2540 336
rect 2494 255 2500 289
rect 2534 255 2540 289
rect 2494 217 2540 255
rect 2494 183 2500 217
rect 2534 183 2540 217
rect 2494 145 2540 183
rect 2494 111 2500 145
rect 2534 111 2540 145
rect 2494 64 2540 111
rect 2590 289 2636 336
rect 2590 255 2596 289
rect 2630 255 2636 289
rect 2590 217 2636 255
rect 2590 183 2596 217
rect 2630 183 2636 217
rect 2590 145 2636 183
rect 2590 111 2596 145
rect 2630 111 2636 145
rect 2590 64 2636 111
rect 2686 289 2732 336
rect 2686 255 2692 289
rect 2726 255 2732 289
rect 2686 217 2732 255
rect 2686 183 2692 217
rect 2726 183 2732 217
rect 2686 145 2732 183
rect 2686 111 2692 145
rect 2726 111 2732 145
rect 2686 64 2732 111
rect 2782 289 2828 336
rect 2782 255 2788 289
rect 2822 255 2828 289
rect 2782 217 2828 255
rect 2782 183 2788 217
rect 2822 183 2828 217
rect 2782 145 2828 183
rect 2782 111 2788 145
rect 2822 111 2828 145
rect 2782 64 2828 111
rect 2878 289 2924 336
rect 2878 255 2884 289
rect 2918 255 2924 289
rect 2878 217 2924 255
rect 2878 183 2884 217
rect 2918 183 2924 217
rect 2878 145 2924 183
rect 2878 111 2884 145
rect 2918 111 2924 145
rect 2878 64 2924 111
rect 2992 320 3038 358
rect 2992 286 2998 320
rect 3032 286 3038 320
rect 2992 248 3038 286
rect 2992 214 2998 248
rect 3032 214 3038 248
rect 2992 176 3038 214
rect 2992 142 2998 176
rect 3032 142 3038 176
rect 2992 104 3038 142
rect 2992 70 2998 104
rect 3032 70 3038 104
rect 1559 -81 1774 -77
rect -229 -111 1774 -81
rect -229 -115 1599 -111
rect -229 -248 -195 -115
rect -37 -248 -3 -115
rect 155 -248 189 -115
rect 347 -248 381 -115
rect 539 -248 573 -115
rect 731 -248 765 -115
rect 839 -241 885 -218
rect -235 -283 -189 -248
rect -235 -317 -229 -283
rect -195 -317 -189 -283
rect -235 -352 -189 -317
rect -139 -283 -93 -248
rect -139 -317 -133 -283
rect -99 -317 -93 -283
rect -139 -352 -93 -317
rect -43 -283 3 -248
rect -43 -317 -37 -283
rect -3 -317 3 -283
rect -43 -352 3 -317
rect 53 -283 99 -248
rect 53 -317 59 -283
rect 93 -317 99 -283
rect 53 -352 99 -317
rect 149 -283 195 -248
rect 149 -317 155 -283
rect 189 -317 195 -283
rect 149 -352 195 -317
rect 245 -283 291 -248
rect 245 -317 251 -283
rect 285 -317 291 -283
rect 245 -352 291 -317
rect 341 -283 387 -248
rect 341 -317 347 -283
rect 381 -317 387 -283
rect 341 -352 387 -317
rect 437 -283 483 -248
rect 437 -317 443 -283
rect 477 -317 483 -283
rect 437 -352 483 -317
rect 533 -283 579 -248
rect 533 -317 539 -283
rect 573 -317 579 -283
rect 533 -352 579 -317
rect 629 -283 675 -248
rect 629 -317 635 -283
rect 669 -317 675 -283
rect 629 -352 675 -317
rect 725 -283 771 -248
rect 725 -317 731 -283
rect 765 -317 771 -283
rect 725 -352 771 -317
rect 839 -275 845 -241
rect 879 -275 885 -241
rect 839 -313 885 -275
rect 839 -347 845 -313
rect 879 -347 885 -313
rect -245 -383 -179 -380
rect -248 -435 -238 -383
rect -186 -435 -176 -383
rect -245 -440 -179 -435
rect -133 -492 -99 -352
rect -53 -383 13 -380
rect -57 -435 -47 -383
rect 5 -435 15 -383
rect -53 -440 13 -435
rect 59 -492 93 -352
rect 139 -383 205 -380
rect 135 -435 145 -383
rect 197 -435 207 -383
rect 139 -440 205 -435
rect 251 -492 285 -352
rect 331 -383 397 -380
rect 327 -435 337 -383
rect 389 -435 399 -383
rect 331 -440 397 -435
rect 443 -492 477 -352
rect 523 -384 589 -380
rect 520 -436 530 -384
rect 582 -436 592 -384
rect 523 -440 589 -436
rect 635 -492 669 -352
rect 715 -384 781 -380
rect 712 -436 722 -384
rect 774 -436 784 -384
rect 839 -385 885 -347
rect 839 -419 845 -385
rect 879 -419 885 -385
rect 715 -440 781 -436
rect -413 -526 669 -492
rect 839 -562 885 -419
rect 1740 -488 1774 -111
rect 1924 -77 1958 64
rect 2116 -77 2150 64
rect 2308 -77 2342 64
rect 2500 -77 2534 64
rect 2692 -77 2726 64
rect 2884 -77 2918 64
rect 2992 26 3038 70
rect 3261 486 4343 520
rect 3261 -77 3295 486
rect 3426 376 3436 428
rect 3488 376 3498 428
rect 3541 336 3575 486
rect 3619 376 3629 428
rect 3681 376 3691 428
rect 3733 336 3767 486
rect 3810 376 3820 428
rect 3872 376 3882 428
rect 3925 336 3959 486
rect 4002 376 4012 428
rect 4064 376 4074 428
rect 4117 336 4151 486
rect 4194 376 4204 428
rect 4256 376 4266 428
rect 4309 336 4343 486
rect 4386 376 4396 428
rect 4448 376 4458 428
rect 4513 392 4559 597
rect 4513 358 4519 392
rect 4553 358 4559 392
rect 3439 289 3485 336
rect 3439 255 3445 289
rect 3479 255 3485 289
rect 3439 217 3485 255
rect 3439 183 3445 217
rect 3479 183 3485 217
rect 3439 145 3485 183
rect 3439 111 3445 145
rect 3479 111 3485 145
rect 3439 64 3485 111
rect 3535 289 3581 336
rect 3535 255 3541 289
rect 3575 255 3581 289
rect 3535 217 3581 255
rect 3535 183 3541 217
rect 3575 183 3581 217
rect 3535 145 3581 183
rect 3535 111 3541 145
rect 3575 111 3581 145
rect 3535 64 3581 111
rect 3631 289 3677 336
rect 3631 255 3637 289
rect 3671 255 3677 289
rect 3631 217 3677 255
rect 3631 183 3637 217
rect 3671 183 3677 217
rect 3631 145 3677 183
rect 3631 111 3637 145
rect 3671 111 3677 145
rect 3631 64 3677 111
rect 3727 289 3773 336
rect 3727 255 3733 289
rect 3767 255 3773 289
rect 3727 217 3773 255
rect 3727 183 3733 217
rect 3767 183 3773 217
rect 3727 145 3773 183
rect 3727 111 3733 145
rect 3767 111 3773 145
rect 3727 64 3773 111
rect 3823 289 3869 336
rect 3823 255 3829 289
rect 3863 255 3869 289
rect 3823 217 3869 255
rect 3823 183 3829 217
rect 3863 183 3869 217
rect 3823 145 3869 183
rect 3823 111 3829 145
rect 3863 111 3869 145
rect 3823 64 3869 111
rect 3919 289 3965 336
rect 3919 255 3925 289
rect 3959 255 3965 289
rect 3919 217 3965 255
rect 3919 183 3925 217
rect 3959 183 3965 217
rect 3919 145 3965 183
rect 3919 111 3925 145
rect 3959 111 3965 145
rect 3919 64 3965 111
rect 4015 289 4061 336
rect 4015 255 4021 289
rect 4055 255 4061 289
rect 4015 217 4061 255
rect 4015 183 4021 217
rect 4055 183 4061 217
rect 4015 145 4061 183
rect 4015 111 4021 145
rect 4055 111 4061 145
rect 4015 64 4061 111
rect 4111 289 4157 336
rect 4111 255 4117 289
rect 4151 255 4157 289
rect 4111 217 4157 255
rect 4111 183 4117 217
rect 4151 183 4157 217
rect 4111 145 4157 183
rect 4111 111 4117 145
rect 4151 111 4157 145
rect 4111 64 4157 111
rect 4207 289 4253 336
rect 4207 255 4213 289
rect 4247 255 4253 289
rect 4207 217 4253 255
rect 4207 183 4213 217
rect 4247 183 4253 217
rect 4207 145 4253 183
rect 4207 111 4213 145
rect 4247 111 4253 145
rect 4207 64 4253 111
rect 4303 289 4349 336
rect 4303 255 4309 289
rect 4343 255 4349 289
rect 4303 217 4349 255
rect 4303 183 4309 217
rect 4343 183 4349 217
rect 4303 145 4349 183
rect 4303 111 4309 145
rect 4343 111 4349 145
rect 4303 64 4349 111
rect 4399 289 4445 336
rect 4399 255 4405 289
rect 4439 255 4445 289
rect 4399 217 4445 255
rect 4399 183 4405 217
rect 4439 183 4445 217
rect 4399 145 4445 183
rect 4399 111 4405 145
rect 4439 111 4445 145
rect 4399 64 4445 111
rect 4513 320 4559 358
rect 4513 286 4519 320
rect 4553 286 4559 320
rect 4513 248 4559 286
rect 4513 214 4519 248
rect 4553 217 4559 248
rect 4732 217 5008 218
rect 4553 214 5008 217
rect 4513 187 5008 214
rect 4513 176 4761 187
rect 4513 142 4519 176
rect 4553 153 4761 176
rect 4795 153 4853 187
rect 4887 153 4945 187
rect 4979 153 5008 187
rect 4553 142 5008 153
rect 4513 122 5008 142
rect 4513 104 4559 122
rect 4513 70 4519 104
rect 4553 70 4559 104
rect 1924 -111 3295 -77
rect 1924 -244 1958 -111
rect 2116 -244 2150 -111
rect 2308 -244 2342 -111
rect 2500 -244 2534 -111
rect 2692 -244 2726 -111
rect 2884 -244 2918 -111
rect 3129 -201 3139 -149
rect 3191 -201 3201 -149
rect 3137 -202 3149 -201
rect 3183 -202 3195 -201
rect 3137 -208 3195 -202
rect 2992 -237 3038 -214
rect 1918 -279 1964 -244
rect 1918 -313 1924 -279
rect 1958 -313 1964 -279
rect 1918 -348 1964 -313
rect 2014 -279 2060 -244
rect 2014 -313 2020 -279
rect 2054 -313 2060 -279
rect 2014 -348 2060 -313
rect 2110 -279 2156 -244
rect 2110 -313 2116 -279
rect 2150 -313 2156 -279
rect 2110 -348 2156 -313
rect 2206 -279 2252 -244
rect 2206 -313 2212 -279
rect 2246 -313 2252 -279
rect 2206 -348 2252 -313
rect 2302 -279 2348 -244
rect 2302 -313 2308 -279
rect 2342 -313 2348 -279
rect 2302 -348 2348 -313
rect 2398 -279 2444 -244
rect 2398 -313 2404 -279
rect 2438 -313 2444 -279
rect 2398 -348 2444 -313
rect 2494 -279 2540 -244
rect 2494 -313 2500 -279
rect 2534 -313 2540 -279
rect 2494 -348 2540 -313
rect 2590 -279 2636 -244
rect 2590 -313 2596 -279
rect 2630 -313 2636 -279
rect 2590 -348 2636 -313
rect 2686 -279 2732 -244
rect 2686 -313 2692 -279
rect 2726 -313 2732 -279
rect 2686 -348 2732 -313
rect 2782 -279 2828 -244
rect 2782 -313 2788 -279
rect 2822 -313 2828 -279
rect 2782 -348 2828 -313
rect 2878 -279 2924 -244
rect 2878 -313 2884 -279
rect 2918 -313 2924 -279
rect 2878 -348 2924 -313
rect 2992 -271 2998 -237
rect 3032 -239 3038 -237
rect 3261 -239 3295 -111
rect 3032 -240 3138 -239
rect 3192 -240 3295 -239
rect 3032 -252 3145 -240
rect 3032 -271 3105 -252
rect 2992 -309 3105 -271
rect 2992 -343 2998 -309
rect 3032 -328 3105 -309
rect 3139 -328 3145 -252
rect 3032 -339 3145 -328
rect 3032 -343 3038 -339
rect 3099 -340 3145 -339
rect 3187 -252 3295 -240
rect 3445 -77 3479 64
rect 3637 -77 3671 64
rect 3829 -77 3863 64
rect 4021 -77 4055 64
rect 4213 -77 4247 64
rect 4405 -77 4439 64
rect 4513 26 4559 70
rect 4635 -57 5242 -23
rect 4635 -77 4669 -57
rect 3445 -111 4669 -77
rect 3445 -244 3479 -111
rect 3637 -244 3671 -111
rect 3829 -244 3863 -111
rect 4021 -244 4055 -111
rect 4213 -244 4247 -111
rect 4405 -244 4439 -111
rect 4896 -115 4970 -114
rect 4784 -117 4858 -116
rect 4784 -169 4795 -117
rect 4847 -169 4858 -117
rect 4896 -167 4907 -115
rect 4959 -167 4970 -115
rect 4896 -168 4970 -167
rect 4784 -170 4858 -169
rect 4513 -237 4559 -214
rect 3187 -328 3193 -252
rect 3227 -328 3295 -252
rect 3187 -339 3295 -328
rect 3187 -340 3233 -339
rect 1908 -379 1974 -376
rect 1905 -431 1915 -379
rect 1967 -431 1977 -379
rect 1908 -436 1974 -431
rect 2020 -488 2054 -348
rect 2100 -379 2166 -376
rect 2096 -431 2106 -379
rect 2158 -431 2168 -379
rect 2100 -436 2166 -431
rect 2212 -488 2246 -348
rect 2292 -379 2358 -376
rect 2288 -431 2298 -379
rect 2350 -431 2360 -379
rect 2292 -436 2358 -431
rect 2404 -488 2438 -348
rect 2484 -379 2550 -376
rect 2480 -431 2490 -379
rect 2542 -431 2552 -379
rect 2484 -436 2550 -431
rect 2596 -488 2630 -348
rect 2676 -380 2742 -376
rect 2673 -432 2683 -380
rect 2735 -432 2745 -380
rect 2676 -436 2742 -432
rect 2788 -488 2822 -348
rect 2868 -380 2934 -376
rect 2865 -432 2875 -380
rect 2927 -432 2937 -380
rect 2992 -381 3038 -343
rect 2992 -415 2998 -381
rect 3032 -415 3038 -381
rect 2868 -436 2934 -432
rect 1740 -522 2822 -488
rect 2992 -598 3038 -415
rect 3261 -488 3295 -339
rect 3439 -279 3485 -244
rect 3439 -313 3445 -279
rect 3479 -313 3485 -279
rect 3439 -348 3485 -313
rect 3535 -279 3581 -244
rect 3535 -313 3541 -279
rect 3575 -313 3581 -279
rect 3535 -348 3581 -313
rect 3631 -279 3677 -244
rect 3631 -313 3637 -279
rect 3671 -313 3677 -279
rect 3631 -348 3677 -313
rect 3727 -279 3773 -244
rect 3727 -313 3733 -279
rect 3767 -313 3773 -279
rect 3727 -348 3773 -313
rect 3823 -279 3869 -244
rect 3823 -313 3829 -279
rect 3863 -313 3869 -279
rect 3823 -348 3869 -313
rect 3919 -279 3965 -244
rect 3919 -313 3925 -279
rect 3959 -313 3965 -279
rect 3919 -348 3965 -313
rect 4015 -279 4061 -244
rect 4015 -313 4021 -279
rect 4055 -313 4061 -279
rect 4015 -348 4061 -313
rect 4111 -279 4157 -244
rect 4111 -313 4117 -279
rect 4151 -313 4157 -279
rect 4111 -348 4157 -313
rect 4207 -279 4253 -244
rect 4207 -313 4213 -279
rect 4247 -313 4253 -279
rect 4207 -348 4253 -313
rect 4303 -279 4349 -244
rect 4303 -313 4309 -279
rect 4343 -313 4349 -279
rect 4303 -348 4349 -313
rect 4399 -279 4445 -244
rect 4399 -313 4405 -279
rect 4439 -313 4445 -279
rect 4399 -348 4445 -313
rect 4513 -271 4519 -237
rect 4553 -271 4559 -237
rect 4513 -309 4559 -271
rect 4513 -343 4519 -309
rect 4553 -326 4559 -309
rect 4553 -343 5008 -326
rect 3429 -379 3495 -376
rect 3426 -431 3436 -379
rect 3488 -431 3498 -379
rect 3429 -436 3495 -431
rect 3541 -488 3575 -348
rect 3621 -379 3687 -376
rect 3617 -431 3627 -379
rect 3679 -431 3689 -379
rect 3621 -436 3687 -431
rect 3733 -488 3767 -348
rect 3813 -379 3879 -376
rect 3809 -431 3819 -379
rect 3871 -431 3881 -379
rect 3813 -436 3879 -431
rect 3925 -488 3959 -348
rect 4005 -379 4071 -376
rect 4001 -431 4011 -379
rect 4063 -431 4073 -379
rect 4005 -436 4071 -431
rect 4117 -488 4151 -348
rect 4197 -380 4263 -376
rect 4194 -432 4204 -380
rect 4256 -432 4266 -380
rect 4197 -436 4263 -432
rect 4309 -488 4343 -348
rect 4513 -357 5008 -343
rect 4389 -380 4455 -376
rect 4386 -432 4396 -380
rect 4448 -432 4458 -380
rect 4513 -381 4761 -357
rect 4513 -415 4519 -381
rect 4553 -391 4761 -381
rect 4795 -391 4853 -357
rect 4887 -391 4945 -357
rect 4979 -391 5008 -357
rect 4553 -415 5008 -391
rect 4513 -422 5008 -415
rect 4389 -436 4455 -432
rect 3261 -522 4343 -488
rect 4513 -597 4559 -422
<< via1 >>
rect -238 414 -186 424
rect -238 380 -229 414
rect -229 380 -195 414
rect -195 380 -186 414
rect -238 372 -186 380
rect -45 414 7 424
rect -45 380 -37 414
rect -37 380 -3 414
rect -3 380 7 414
rect -45 372 7 380
rect 146 414 198 424
rect 146 380 155 414
rect 155 380 189 414
rect 189 380 198 414
rect 146 372 198 380
rect 338 414 390 424
rect 338 380 347 414
rect 347 380 381 414
rect 381 380 390 414
rect 338 372 390 380
rect 530 414 582 424
rect 530 380 539 414
rect 539 380 573 414
rect 573 380 582 414
rect 530 372 582 380
rect 722 414 774 424
rect 722 380 731 414
rect 731 380 765 414
rect 765 380 774 414
rect 722 372 774 380
rect 980 365 1036 425
rect 1250 365 1310 425
rect 1508 16 1562 76
rect 1915 418 1967 428
rect 1915 384 1924 418
rect 1924 384 1958 418
rect 1958 384 1967 418
rect 1915 376 1967 384
rect 2108 418 2160 428
rect 2108 384 2116 418
rect 2116 384 2150 418
rect 2150 384 2160 418
rect 2108 376 2160 384
rect 2299 418 2351 428
rect 2299 384 2308 418
rect 2308 384 2342 418
rect 2342 384 2351 418
rect 2299 376 2351 384
rect 2491 418 2543 428
rect 2491 384 2500 418
rect 2500 384 2534 418
rect 2534 384 2543 418
rect 2491 376 2543 384
rect 2683 418 2735 428
rect 2683 384 2692 418
rect 2692 384 2726 418
rect 2726 384 2735 418
rect 2683 376 2735 384
rect 2875 418 2927 428
rect 2875 384 2884 418
rect 2884 384 2918 418
rect 2918 384 2927 418
rect 2875 376 2927 384
rect -238 -394 -186 -383
rect -238 -428 -229 -394
rect -229 -428 -195 -394
rect -195 -428 -186 -394
rect -238 -435 -186 -428
rect -47 -394 5 -383
rect -47 -428 -37 -394
rect -37 -428 -3 -394
rect -3 -428 5 -394
rect -47 -435 5 -428
rect 145 -394 197 -383
rect 145 -428 155 -394
rect 155 -428 189 -394
rect 189 -428 197 -394
rect 145 -435 197 -428
rect 337 -394 389 -383
rect 337 -428 347 -394
rect 347 -428 381 -394
rect 381 -428 389 -394
rect 337 -435 389 -428
rect 530 -394 582 -384
rect 530 -428 539 -394
rect 539 -428 573 -394
rect 573 -428 582 -394
rect 530 -436 582 -428
rect 722 -394 774 -384
rect 722 -428 731 -394
rect 731 -428 765 -394
rect 765 -428 774 -394
rect 722 -436 774 -428
rect 3436 418 3488 428
rect 3436 384 3445 418
rect 3445 384 3479 418
rect 3479 384 3488 418
rect 3436 376 3488 384
rect 3629 418 3681 428
rect 3629 384 3637 418
rect 3637 384 3671 418
rect 3671 384 3681 418
rect 3629 376 3681 384
rect 3820 418 3872 428
rect 3820 384 3829 418
rect 3829 384 3863 418
rect 3863 384 3872 418
rect 3820 376 3872 384
rect 4012 418 4064 428
rect 4012 384 4021 418
rect 4021 384 4055 418
rect 4055 384 4064 418
rect 4012 376 4064 384
rect 4204 418 4256 428
rect 4204 384 4213 418
rect 4213 384 4247 418
rect 4247 384 4256 418
rect 4204 376 4256 384
rect 4396 418 4448 428
rect 4396 384 4405 418
rect 4405 384 4439 418
rect 4439 384 4448 418
rect 4396 376 4448 384
rect 3139 -168 3191 -149
rect 3139 -201 3149 -168
rect 3149 -201 3183 -168
rect 3183 -201 3191 -168
rect 4795 -127 4847 -117
rect 4795 -161 4806 -127
rect 4806 -161 4840 -127
rect 4840 -161 4847 -127
rect 4795 -169 4847 -161
rect 4907 -122 4959 -115
rect 4907 -156 4908 -122
rect 4908 -156 4942 -122
rect 4942 -156 4959 -122
rect 4907 -167 4959 -156
rect 1915 -390 1967 -379
rect 1915 -424 1924 -390
rect 1924 -424 1958 -390
rect 1958 -424 1967 -390
rect 1915 -431 1967 -424
rect 2106 -390 2158 -379
rect 2106 -424 2116 -390
rect 2116 -424 2150 -390
rect 2150 -424 2158 -390
rect 2106 -431 2158 -424
rect 2298 -390 2350 -379
rect 2298 -424 2308 -390
rect 2308 -424 2342 -390
rect 2342 -424 2350 -390
rect 2298 -431 2350 -424
rect 2490 -390 2542 -379
rect 2490 -424 2500 -390
rect 2500 -424 2534 -390
rect 2534 -424 2542 -390
rect 2490 -431 2542 -424
rect 2683 -390 2735 -380
rect 2683 -424 2692 -390
rect 2692 -424 2726 -390
rect 2726 -424 2735 -390
rect 2683 -432 2735 -424
rect 2875 -390 2927 -380
rect 2875 -424 2884 -390
rect 2884 -424 2918 -390
rect 2918 -424 2927 -390
rect 2875 -432 2927 -424
rect 3436 -390 3488 -379
rect 3436 -424 3445 -390
rect 3445 -424 3479 -390
rect 3479 -424 3488 -390
rect 3436 -431 3488 -424
rect 3627 -390 3679 -379
rect 3627 -424 3637 -390
rect 3637 -424 3671 -390
rect 3671 -424 3679 -390
rect 3627 -431 3679 -424
rect 3819 -390 3871 -379
rect 3819 -424 3829 -390
rect 3829 -424 3863 -390
rect 3863 -424 3871 -390
rect 3819 -431 3871 -424
rect 4011 -390 4063 -379
rect 4011 -424 4021 -390
rect 4021 -424 4055 -390
rect 4055 -424 4063 -390
rect 4011 -431 4063 -424
rect 4204 -390 4256 -380
rect 4204 -424 4213 -390
rect 4213 -424 4247 -390
rect 4247 -424 4256 -390
rect 4204 -432 4256 -424
rect 4396 -390 4448 -380
rect 4396 -424 4405 -390
rect 4405 -424 4439 -390
rect 4439 -424 4448 -390
rect 4396 -432 4448 -424
<< metal2 >>
rect -238 424 -186 434
rect -45 424 7 434
rect 146 424 198 434
rect 338 424 390 434
rect 530 424 582 434
rect 722 424 774 434
rect 980 425 1036 435
rect -516 372 -238 424
rect -186 372 -45 424
rect 7 372 146 424
rect 198 372 338 424
rect 390 372 530 424
rect 582 372 722 424
rect 774 372 980 424
rect -238 362 -186 372
rect -45 362 7 372
rect 146 362 198 372
rect 338 362 390 372
rect 530 362 582 372
rect 722 362 774 372
rect 980 355 1036 365
rect 1250 425 1310 435
rect 1915 428 1967 438
rect 2108 428 2160 438
rect 2299 428 2351 438
rect 2491 428 2543 438
rect 2683 428 2735 438
rect 2875 428 2927 438
rect 3436 428 3488 438
rect 3629 428 3681 438
rect 3820 428 3872 438
rect 4012 428 4064 438
rect 4204 428 4256 438
rect 4396 428 4448 438
rect 1637 376 1915 428
rect 1967 376 2108 428
rect 2160 376 2299 428
rect 2351 376 2491 428
rect 2543 376 2683 428
rect 2735 376 2875 428
rect 2927 376 3436 428
rect 3488 376 3629 428
rect 3681 376 3820 428
rect 3872 376 4012 428
rect 4064 376 4204 428
rect 4256 376 4396 428
rect 4448 376 5274 428
rect 1915 366 1967 376
rect 2108 366 2160 376
rect 2299 366 2351 376
rect 2491 366 2543 376
rect 2683 366 2735 376
rect 2875 366 2927 376
rect 1250 229 1310 365
rect 1508 76 1562 86
rect 1562 16 1564 76
rect 1508 -44 1564 16
rect -238 -383 -186 -373
rect -47 -383 5 -373
rect 145 -383 197 -373
rect 337 -383 389 -373
rect 530 -383 582 -374
rect 722 -383 774 -374
rect -515 -435 -238 -383
rect -186 -435 -47 -383
rect 5 -435 145 -383
rect 197 -435 337 -383
rect 389 -384 1182 -383
rect 389 -435 530 -384
rect -238 -445 -186 -435
rect -47 -445 5 -435
rect 145 -445 197 -435
rect 337 -445 389 -435
rect 582 -435 722 -384
rect 530 -446 582 -436
rect 774 -435 1182 -384
rect 722 -446 774 -436
rect 1509 -521 1564 -44
rect 3139 -149 3191 376
rect 3436 366 3488 376
rect 3629 366 3681 376
rect 3820 366 3872 376
rect 4012 366 4064 376
rect 4204 366 4256 376
rect 4396 366 4448 376
rect 4794 -117 4848 -106
rect 4794 -124 4795 -117
rect 3139 -211 3191 -201
rect 4636 -169 4795 -124
rect 4847 -169 4848 -117
rect 4636 -176 4848 -169
rect 1915 -379 1967 -369
rect 2106 -379 2158 -369
rect 2298 -379 2350 -369
rect 2490 -379 2542 -369
rect 2683 -379 2735 -370
rect 2875 -379 2927 -370
rect 3436 -379 3488 -369
rect 3627 -379 3679 -369
rect 3819 -379 3871 -369
rect 4011 -379 4063 -369
rect 4204 -379 4256 -370
rect 4396 -379 4448 -370
rect 4636 -379 4688 -176
rect 4794 -180 4848 -176
rect 4906 -108 4960 -104
rect 5066 -108 5118 376
rect 4906 -115 5118 -108
rect 4906 -167 4907 -115
rect 4959 -160 5118 -115
rect 4959 -167 4960 -160
rect 4906 -178 4960 -167
rect 1638 -431 1915 -379
rect 1967 -431 2106 -379
rect 2158 -431 2298 -379
rect 2350 -431 2490 -379
rect 2542 -380 3436 -379
rect 2542 -431 2683 -380
rect 1915 -441 1967 -431
rect 2106 -441 2158 -431
rect 2298 -441 2350 -431
rect 2490 -441 2542 -431
rect 2735 -431 2875 -380
rect 2683 -442 2735 -432
rect 2927 -431 3436 -380
rect 3488 -431 3627 -379
rect 3679 -431 3819 -379
rect 3871 -431 4011 -379
rect 4063 -380 4688 -379
rect 4063 -431 4204 -380
rect 2875 -442 2927 -432
rect 3436 -441 3488 -431
rect 3627 -441 3679 -431
rect 3819 -441 3871 -431
rect 4011 -441 4063 -431
rect 4256 -431 4396 -380
rect 4204 -442 4256 -432
rect 4448 -431 4688 -380
rect 4396 -442 4448 -432
<< labels >>
flabel metal2 5222 376 5274 428 1 FreeSans 480 0 0 0 con_en_b
flabel space 5142 -58 5182 -22 1 FreeSans 480 0 0 0 out
flabel metal2 -516 372 -464 424 1 FreeSans 480 0 0 0 tgate_flat_0/en_b
flabel metal2 -514 -435 -454 -383 1 FreeSans 480 0 0 0 tgate_flat_0/en
flabel metal1 862 -559 862 -559 1 FreeSans 500 0 0 0 tgate_flat_0/VSS
flabel metal1 862 547 862 547 5 FreeSans 500 0 0 0 tgate_flat_0/VDD
flabel metal1 953 -99 953 -99 7 FreeSans 500 0 0 0 tgate_flat_0/out
flabel metal1 -538 -98 -538 -98 3 FreeSans 500 0 0 0 tgate_flat_0/in
flabel metal1 3015 591 3015 591 1 FreeSans 400 0 0 0 switch_5t_0/VDD
flabel metal1 3015 -591 3015 -591 1 FreeSans 400 0 0 0 switch_5t_0/VSS
flabel metal1 1568 -94 1568 -94 1 FreeSans 400 0 0 0 switch_5t_0/in
flabel metal1 4663 -95 4663 -95 7 FreeSans 400 0 0 0 switch_5t_0/out
flabel metal1 4536 592 4536 592 1 FreeSans 400 0 0 0 switch_5t_0/VDD
flabel metal1 4536 -590 4536 -590 1 FreeSans 400 0 0 0 switch_5t_0/VSS
flabel metal1 1615 -94 1615 -94 3 FreeSans 500 0 0 0 switch_5t_0/transmission_gate_0/in
flabel metal1 3106 -95 3106 -95 7 FreeSans 500 0 0 0 switch_5t_0/transmission_gate_0/out
flabel metal1 3015 551 3015 551 5 FreeSans 500 0 0 0 switch_5t_0/transmission_gate_0/VDD
flabel metal1 3015 -555 3015 -555 1 FreeSans 500 0 0 0 switch_5t_0/transmission_gate_0/VSS
flabel metal2 1639 -431 1699 -379 1 FreeSans 480 0 0 0 switch_5t_0/transmission_gate_0/en
flabel metal2 1637 376 1689 428 1 FreeSans 480 0 0 0 switch_5t_0/transmission_gate_0/en_b
flabel metal1 3136 -94 3136 -94 3 FreeSans 500 0 0 0 switch_5t_0/transmission_gate_1/in
flabel metal1 4627 -95 4627 -95 7 FreeSans 500 0 0 0 switch_5t_0/transmission_gate_1/out
flabel metal1 4536 551 4536 551 5 FreeSans 500 0 0 0 switch_5t_0/transmission_gate_1/VDD
flabel metal1 4536 -555 4536 -555 1 FreeSans 500 0 0 0 switch_5t_0/transmission_gate_1/VSS
flabel metal2 3160 -431 3220 -379 1 FreeSans 480 0 0 0 switch_5t_0/transmission_gate_1/en
flabel metal2 3158 376 3210 428 1 FreeSans 480 0 0 0 switch_5t_0/transmission_gate_1/en_b
flabel locali 4810 -85 4844 -51 0 FreeSans 340 0 0 0 sky130_fd_sc_hd__inv_1_0/Y
flabel locali 4810 -153 4844 -119 0 FreeSans 340 0 0 0 sky130_fd_sc_hd__inv_1_0/Y
flabel locali 4902 -153 4936 -119 0 FreeSans 340 0 0 0 sky130_fd_sc_hd__inv_1_0/A
flabel nwell 4945 153 4979 187 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__inv_1_0/VPB
flabel pwell 4945 -391 4979 -357 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__inv_1_0/VNB
flabel metal1 4945 -391 4979 -357 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__inv_1_0/VGND
flabel metal1 4945 153 4979 187 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__inv_1_0/VPWR
rlabel comment 5008 -374 5008 -374 6 sky130_fd_sc_hd__inv_1_0/inv_1
<< end >>
