//-----------------------------------------------------------------------------
// GcdUnit
//-----------------------------------------------------------------------------
// dump-vcd: False
// verilator-xinit: zeros
module macro (
    inout porst,
    inout va, 
    inout vb,
    inout vbg
 );
endmodule


