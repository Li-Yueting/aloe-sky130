VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO sky130_asc_nfet_01v8_lvt_9
  CLASS CORE ;
  FOREIGN sky130_asc_nfet_01v8_lvt_9 ;
  ORIGIN 0.000 0.000 ;
  SIZE 22.590 BY 9.400 ;
  SITE unitasc ;
  PIN GATE
    DIRECTION INOUT ;
    ANTENNAGATEAREA 72.000000 ;
    PORT
      LAYER li1 ;
        RECT 1.490 1.520 21.990 1.820 ;
    END
  END GATE
  PIN SOURCE
    DIRECTION INOUT ;
    ANTENNADIFFAREA 5.800000 ;
    PORT
      LAYER li1 ;
        RECT 1.090 8.450 21.990 8.750 ;
        RECT 3.435 7.020 3.605 8.450 ;
        RECT 8.015 7.020 8.185 8.450 ;
        RECT 12.595 7.020 12.765 8.450 ;
        RECT 17.175 7.020 17.345 8.450 ;
        RECT 21.755 7.020 21.925 8.450 ;
        RECT 3.435 6.930 3.610 7.020 ;
        RECT 8.015 6.930 8.190 7.020 ;
        RECT 12.595 6.930 12.770 7.020 ;
        RECT 17.175 6.930 17.350 7.020 ;
        RECT 21.755 6.930 21.930 7.020 ;
        RECT 3.440 2.980 3.610 6.930 ;
        RECT 8.020 2.980 8.190 6.930 ;
        RECT 12.600 2.980 12.770 6.930 ;
        RECT 17.180 2.980 17.350 6.930 ;
        RECT 21.760 2.980 21.930 6.930 ;
      LAYER mcon ;
        RECT 3.440 3.060 3.610 6.940 ;
        RECT 8.020 3.060 8.190 6.940 ;
        RECT 12.600 3.060 12.770 6.940 ;
        RECT 17.180 3.060 17.350 6.940 ;
        RECT 21.760 3.060 21.930 6.940 ;
      LAYER met1 ;
        RECT 3.410 3.000 3.640 7.000 ;
        RECT 7.990 3.000 8.220 7.000 ;
        RECT 12.570 3.000 12.800 7.000 ;
        RECT 17.150 3.000 17.380 7.000 ;
        RECT 21.730 3.000 21.960 7.000 ;
    END
  END SOURCE
  PIN DRAIN
    DIRECTION INOUT ;
    ANTENNADIFFAREA 5.800000 ;
    PORT
      LAYER li1 ;
        RECT 1.150 3.270 1.320 7.020 ;
        RECT 5.730 3.270 5.900 7.020 ;
        RECT 10.310 3.270 10.480 7.020 ;
        RECT 14.890 3.270 15.060 7.020 ;
        RECT 19.470 3.270 19.640 7.020 ;
        RECT 1.145 2.980 1.320 3.270 ;
        RECT 5.725 2.980 5.900 3.270 ;
        RECT 10.305 2.980 10.480 3.270 ;
        RECT 14.885 2.980 15.060 3.270 ;
        RECT 19.465 2.980 19.640 3.270 ;
        RECT 1.145 2.650 1.315 2.980 ;
        RECT 5.725 2.650 5.895 2.980 ;
        RECT 10.305 2.650 10.475 2.980 ;
        RECT 14.885 2.650 15.055 2.980 ;
        RECT 19.465 2.650 19.635 2.980 ;
        RECT 1.090 2.350 21.990 2.650 ;
      LAYER mcon ;
        RECT 1.150 3.060 1.320 6.940 ;
        RECT 5.730 3.060 5.900 6.940 ;
        RECT 10.310 3.060 10.480 6.940 ;
        RECT 14.890 3.060 15.060 6.940 ;
        RECT 19.470 3.060 19.640 6.940 ;
      LAYER met1 ;
        RECT 1.120 3.000 1.350 7.000 ;
        RECT 5.700 3.000 5.930 7.000 ;
        RECT 10.280 3.000 10.510 7.000 ;
        RECT 14.860 3.000 15.090 7.000 ;
        RECT 19.440 3.000 19.670 7.000 ;
    END
  END DRAIN
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER li1 ;
        RECT 0.600 9.250 21.990 9.550 ;
      LAYER mcon ;
        RECT 1.940 9.250 2.240 9.550 ;
        RECT 3.940 9.250 4.240 9.550 ;
        RECT 5.940 9.250 6.240 9.550 ;
        RECT 7.940 9.250 8.240 9.550 ;
        RECT 9.940 9.250 10.240 9.550 ;
        RECT 11.940 9.250 12.240 9.550 ;
        RECT 13.940 9.250 14.240 9.550 ;
        RECT 15.940 9.250 16.240 9.550 ;
        RECT 17.940 9.250 18.240 9.550 ;
        RECT 19.940 9.250 20.240 9.550 ;
      LAYER met1 ;
        RECT 0.600 9.100 21.990 9.700 ;
    END
  END VPWR
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.600 0.150 21.990 7.130 ;
      LAYER li1 ;
        RECT 0.740 0.150 1.040 1.200 ;
        RECT 5.990 0.150 6.790 0.750 ;
        RECT 12.490 0.150 13.290 0.750 ;
        RECT 0.600 -0.150 21.990 0.150 ;
      LAYER mcon ;
        RECT 1.940 -0.150 2.240 0.150 ;
        RECT 3.940 -0.150 4.240 0.150 ;
        RECT 5.940 -0.150 6.240 0.150 ;
        RECT 7.940 -0.150 8.240 0.150 ;
        RECT 9.940 -0.150 10.240 0.150 ;
        RECT 11.940 -0.150 12.240 0.150 ;
        RECT 13.940 -0.150 14.240 0.150 ;
        RECT 15.940 -0.150 16.240 0.150 ;
        RECT 17.940 -0.150 18.240 0.150 ;
        RECT 19.940 -0.150 20.240 0.150 ;
      LAYER met1 ;
        RECT 0.600 -0.300 21.990 0.300 ;
    END
  END VGND
END sky130_asc_nfet_01v8_lvt_9
END LIBRARY

