* NGSPICE file created from bgr_top.ext - technology: sky130A

.subckt sky130_asc_res_xhigh_po_2p85_1 Rin Rout VPWR VGND a_2148_115#
X0 Rin a_2148_115# VGND sky130_fd_pr__res_xhigh_po_2p85 l=7.88e+06u
X1 Rout a_2148_115# VGND sky130_fd_pr__res_xhigh_po_2p85 l=7.88e+06u
C0 Rin Rout 0.12fF
C1 Rin VPWR 0.17fF
C2 VPWR a_2148_115# 0.17fF
C3 VPWR VGND 2.31fF
C4 Rout VGND 1.26fF
C5 Rin VGND 0.78fF
C6 a_2148_115# VGND 2.70fF
.ends

.subckt sky130_asc_pfet_01v8_lvt_60 GATE SOURCE DRAIN VGND VPWR VSUBS
X0 DRAIN GATE SOURCE VPWR sky130_fd_pr__pfet_01v8_lvt ad=5.79855e+13p pd=4.1788e+08u as=5.6115e+13p ps=4.044e+08u w=6.45e+06u l=2e+06u
X1 SOURCE GATE DRAIN VPWR sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=6.45e+06u l=2e+06u
X2 DRAIN GATE SOURCE VPWR sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=6.45e+06u l=2e+06u
X3 SOURCE GATE DRAIN VPWR sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=6.45e+06u l=2e+06u
X4 DRAIN GATE SOURCE VPWR sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=6.45e+06u l=2e+06u
X5 DRAIN GATE SOURCE VPWR sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=6.45e+06u l=2e+06u
X6 DRAIN GATE SOURCE VPWR sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=6.45e+06u l=2e+06u
X7 DRAIN GATE SOURCE VPWR sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=6.45e+06u l=2e+06u
X8 DRAIN GATE SOURCE VPWR sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=6.45e+06u l=2e+06u
X9 SOURCE GATE DRAIN VPWR sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=6.45e+06u l=2e+06u
X10 DRAIN GATE SOURCE VPWR sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=6.45e+06u l=2e+06u
X11 SOURCE GATE DRAIN VPWR sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=6.45e+06u l=2e+06u
X12 SOURCE GATE DRAIN VPWR sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=6.45e+06u l=2e+06u
X13 DRAIN GATE SOURCE VPWR sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=6.45e+06u l=2e+06u
X14 DRAIN GATE SOURCE VPWR sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=6.45e+06u l=2e+06u
X15 SOURCE GATE DRAIN VPWR sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=6.45e+06u l=2e+06u
X16 SOURCE GATE DRAIN VPWR sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=6.45e+06u l=2e+06u
X17 DRAIN GATE SOURCE VPWR sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=6.45e+06u l=2e+06u
X18 SOURCE GATE DRAIN VPWR sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=6.45e+06u l=2e+06u
X19 DRAIN GATE SOURCE VPWR sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=6.45e+06u l=2e+06u
X20 SOURCE GATE DRAIN VPWR sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=6.45e+06u l=2e+06u
X21 DRAIN GATE SOURCE VPWR sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=6.45e+06u l=2e+06u
X22 SOURCE GATE DRAIN VPWR sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=6.45e+06u l=2e+06u
X23 DRAIN GATE SOURCE VPWR sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=6.45e+06u l=2e+06u
X24 SOURCE GATE DRAIN VPWR sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=6.45e+06u l=2e+06u
X25 DRAIN GATE SOURCE VPWR sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=6.45e+06u l=2e+06u
X26 SOURCE GATE DRAIN VPWR sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=6.45e+06u l=2e+06u
X27 SOURCE GATE DRAIN VPWR sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=6.45e+06u l=2e+06u
X28 DRAIN GATE SOURCE VPWR sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=6.45e+06u l=2e+06u
X29 SOURCE GATE DRAIN VPWR sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=6.45e+06u l=2e+06u
X30 DRAIN GATE SOURCE VPWR sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=6.45e+06u l=2e+06u
X31 SOURCE GATE DRAIN VPWR sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=6.45e+06u l=2e+06u
X32 DRAIN GATE SOURCE VPWR sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=6.45e+06u l=2e+06u
X33 SOURCE GATE DRAIN VPWR sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=6.45e+06u l=2e+06u
X34 DRAIN GATE SOURCE VPWR sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=6.45e+06u l=2e+06u
X35 SOURCE GATE DRAIN VPWR sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=6.45e+06u l=2e+06u
X36 DRAIN GATE SOURCE VPWR sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=6.45e+06u l=2e+06u
X37 SOURCE GATE DRAIN VPWR sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=6.45e+06u l=2e+06u
X38 DRAIN GATE SOURCE VPWR sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=6.45e+06u l=2e+06u
X39 SOURCE GATE DRAIN VPWR sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=6.45e+06u l=2e+06u
X40 SOURCE GATE DRAIN VPWR sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=6.45e+06u l=2e+06u
X41 DRAIN GATE SOURCE VPWR sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=6.45e+06u l=2e+06u
X42 DRAIN GATE SOURCE VPWR sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=6.45e+06u l=2e+06u
X43 DRAIN GATE SOURCE VPWR sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=6.45e+06u l=2e+06u
X44 SOURCE GATE DRAIN VPWR sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=6.45e+06u l=2e+06u
X45 SOURCE GATE DRAIN VPWR sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=6.45e+06u l=2e+06u
X46 DRAIN GATE SOURCE VPWR sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=6.45e+06u l=2e+06u
X47 SOURCE GATE DRAIN VPWR sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=6.45e+06u l=2e+06u
X48 SOURCE GATE DRAIN VPWR sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=6.45e+06u l=2e+06u
X49 SOURCE GATE DRAIN VPWR sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=6.45e+06u l=2e+06u
X50 DRAIN GATE SOURCE VPWR sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=6.45e+06u l=2e+06u
X51 SOURCE GATE DRAIN VPWR sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=6.45e+06u l=2e+06u
X52 SOURCE GATE DRAIN VPWR sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=6.45e+06u l=2e+06u
X53 SOURCE GATE DRAIN VPWR sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=6.45e+06u l=2e+06u
X54 DRAIN GATE SOURCE VPWR sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=6.45e+06u l=2e+06u
X55 SOURCE GATE DRAIN VPWR sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=6.45e+06u l=2e+06u
X56 DRAIN GATE SOURCE VPWR sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=6.45e+06u l=2e+06u
X57 DRAIN GATE SOURCE VPWR sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=6.45e+06u l=2e+06u
X58 SOURCE GATE DRAIN VPWR sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=6.45e+06u l=2e+06u
X59 DRAIN GATE SOURCE VPWR sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=6.45e+06u l=2e+06u
C0 DRAIN VPWR 1.83fF
C1 DRAIN VGND 5.28fF
C2 VPWR SOURCE 22.83fF
C3 VGND SOURCE 0.32fF
C4 DRAIN SOURCE 1.25fF
C5 GATE VPWR 27.32fF
C6 VGND GATE 12.31fF
C7 DRAIN GATE 25.46fF
C8 GATE SOURCE 0.18fF
C9 VGND VSUBS 25.41fF
C10 SOURCE VSUBS 0.00fF
C11 DRAIN VSUBS 9.62fF
C12 GATE VSUBS 30.27fF
C13 VPWR VSUBS 142.65fF
.ends

.subckt sky130_asc_pnp_05v5_W3p40L3p40_7 Emitter Base Collector VPWR VGND
X0 Collector Base Emitter sky130_fd_pr__pnp_05v5_W3p40L3p40
X1 Collector Base Emitter sky130_fd_pr__pnp_05v5_W3p40L3p40
X2 Collector Base Emitter sky130_fd_pr__pnp_05v5_W3p40L3p40
X3 Collector Base Emitter sky130_fd_pr__pnp_05v5_W3p40L3p40
X4 Collector Base Emitter sky130_fd_pr__pnp_05v5_W3p40L3p40
X5 Collector Base Emitter sky130_fd_pr__pnp_05v5_W3p40L3p40
X6 Collector Base Emitter sky130_fd_pr__pnp_05v5_W3p40L3p40
C0 Base Emitter 18.67fF
C1 VGND Collector 9.81fF
C2 VPWR Collector 11.49fF
C3 Emitter Collector 9.06fF
C4 Base Collector 28.86fF
.ends

.subckt sky130_asc_res_xhigh_po_2p85_2 Rin Rout VPWR a_2723_115# VGND
X0 Rout a_2723_115# VGND sky130_fd_pr__res_xhigh_po w=2.85e+06u l=1.075e+07u
X1 Rin a_2723_115# VGND sky130_fd_pr__res_xhigh_po w=2.85e+06u l=1.075e+07u
C0 VPWR Rin 0.17fF
C1 Rout Rin 0.12fF
C2 VPWR a_2723_115# 0.17fF
C3 VPWR VGND 2.83fF
C4 Rout VGND 1.26fF
C5 Rin VGND 0.78fF
C6 a_2723_115# VGND 2.70fF
.ends

.subckt sky130_asc_pfet_01v8_lvt_12 GATE SOURCE DRAIN VGND VPWR VSUBS
X0 SOURCE GATE DRAIN VPWR sky130_fd_pr__pfet_01v8_lvt ad=1.1223e+13p pd=8.088e+07u as=1.30935e+13p ps=9.436e+07u w=6.45e+06u l=2e+06u
X1 DRAIN GATE SOURCE VPWR sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=6.45e+06u l=2e+06u
X2 DRAIN GATE SOURCE VPWR sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=6.45e+06u l=2e+06u
X3 SOURCE GATE DRAIN VPWR sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=6.45e+06u l=2e+06u
X4 SOURCE GATE DRAIN VPWR sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=6.45e+06u l=2e+06u
X5 DRAIN GATE SOURCE VPWR sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=6.45e+06u l=2e+06u
X6 SOURCE GATE DRAIN VPWR sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=6.45e+06u l=2e+06u
X7 DRAIN GATE SOURCE VPWR sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=6.45e+06u l=2e+06u
X8 DRAIN GATE SOURCE VPWR sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=6.45e+06u l=2e+06u
X9 SOURCE GATE DRAIN VPWR sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=6.45e+06u l=2e+06u
X10 SOURCE GATE DRAIN VPWR sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=6.45e+06u l=2e+06u
X11 DRAIN GATE SOURCE VPWR sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=6.45e+06u l=2e+06u
C0 SOURCE VGND 0.06fF
C1 GATE SOURCE 0.04fF
C2 GATE VGND 2.51fF
C3 SOURCE VPWR 4.54fF
C4 GATE VPWR 5.46fF
C5 DRAIN SOURCE 0.26fF
C6 DRAIN VGND 1.08fF
C7 GATE DRAIN 5.17fF
C8 DRAIN VPWR 0.42fF
C9 VGND VSUBS 5.31fF
C10 SOURCE VSUBS 0.00fF
C11 DRAIN VSUBS 1.99fF
C12 GATE VSUBS 6.20fF
C13 VPWR VSUBS 29.52fF
.ends

.subckt sky130_asc_nfet_01v8_lvt_9 GATE SOURCE DRAIN VPWR VGND
X0 SOURCE GATE DRAIN VGND sky130_fd_pr__nfet_01v8_lvt ad=5.8e+12p pd=4.29e+07u as=5.8e+12p ps=4.29e+07u w=4e+06u l=2e+06u
X1 SOURCE GATE DRAIN VGND sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=2e+06u
X2 DRAIN GATE SOURCE VGND sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=2e+06u
X3 SOURCE GATE DRAIN VGND sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=2e+06u
X4 DRAIN GATE SOURCE VGND sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=2e+06u
X5 SOURCE GATE DRAIN VGND sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=2e+06u
X6 DRAIN GATE SOURCE VGND sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=2e+06u
X7 SOURCE GATE DRAIN VGND sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=2e+06u
X8 DRAIN GATE SOURCE VGND sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=2e+06u
C0 VPWR SOURCE 1.38fF
C1 GATE SOURCE 0.01fF
C2 SOURCE DRAIN 0.05fF
C3 GATE DRAIN 1.66fF
C4 VPWR VGND 3.99fF
C5 SOURCE VGND 2.64fF
C6 DRAIN VGND 2.28fF
C7 GATE VGND 11.48fF
.ends

.subckt sky130_asc_pfet_01v8_lvt_6 GATE SOURCE DRAIN VGND VPWR VSUBS
X0 SOURCE GATE DRAIN VPWR sky130_fd_pr__pfet_01v8_lvt ad=5.6115e+12p pd=4.044e+07u as=7.482e+12p ps=5.392e+07u w=6.45e+06u l=2e+06u
X1 SOURCE GATE DRAIN VPWR sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=6.45e+06u l=2e+06u
X2 DRAIN GATE SOURCE VPWR sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=6.45e+06u l=2e+06u
X3 DRAIN GATE SOURCE VPWR sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=6.45e+06u l=2e+06u
X4 SOURCE GATE DRAIN VPWR sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=6.45e+06u l=2e+06u
X5 DRAIN GATE SOURCE VPWR sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=6.45e+06u l=2e+06u
C0 GATE VGND 1.28fF
C1 GATE VPWR 2.73fF
C2 GATE DRAIN 2.63fF
C3 DRAIN VGND 0.56fF
C4 VPWR DRAIN 0.24fF
C5 GATE SOURCE 0.02fF
C6 SOURCE VGND 0.03fF
C7 VPWR SOURCE 2.27fF
C8 SOURCE DRAIN 0.14fF
C9 VGND VSUBS 2.79fF
C10 SOURCE VSUBS 0.00fF
C11 DRAIN VSUBS 1.04fF
C12 GATE VSUBS 3.19fF
C13 VPWR VSUBS 15.38fF
.ends

.subckt sky130_asc_pnp_05v5_W3p40L3p40_1 Emitter Base Collector VPWR VGND
X0 Collector Base Emitter sky130_fd_pr__pnp_05v5_W3p40L3p40
C0 Emitter Base 1.55fF
C1 VGND Collector 1.50fF
C2 VPWR Collector 1.46fF
C3 Emitter Collector 0.40fF
C4 Base Collector 3.33fF
.ends

.subckt sky130_asc_cap_mim_m3_1 Cin Cout VPWR VGND VSUBS
X0 Cout Cin sky130_fd_pr__cap_mim_m3_1 l=2e+06u w=2e+06u
X1 Cout Cin sky130_fd_pr__cap_mim_m3_1 l=2e+06u w=2e+06u
X2 Cout Cin sky130_fd_pr__cap_mim_m3_1 l=2e+06u w=2e+06u
X3 Cout Cin sky130_fd_pr__cap_mim_m3_1 l=2e+06u w=2e+06u
X4 Cout Cin sky130_fd_pr__cap_mim_m3_1 l=2e+06u w=2e+06u
X5 Cout Cin sky130_fd_pr__cap_mim_m3_1 l=2e+06u w=2e+06u
X6 Cout Cin sky130_fd_pr__cap_mim_m3_1 l=2e+06u w=2e+06u
X7 Cout Cin sky130_fd_pr__cap_mim_m3_1 l=2e+06u w=2e+06u
X8 Cout Cin sky130_fd_pr__cap_mim_m3_1 l=2e+06u w=2e+06u
X9 Cout Cin sky130_fd_pr__cap_mim_m3_1 l=2e+06u w=2e+06u
X10 Cout Cin sky130_fd_pr__cap_mim_m3_1 l=2e+06u w=2e+06u
X11 Cout Cin sky130_fd_pr__cap_mim_m3_1 l=2e+06u w=2e+06u
X12 Cout Cin sky130_fd_pr__cap_mim_m3_1 l=2e+06u w=2e+06u
X13 Cout Cin sky130_fd_pr__cap_mim_m3_1 l=2e+06u w=2e+06u
X14 Cout Cin sky130_fd_pr__cap_mim_m3_1 l=2e+06u w=2e+06u
X15 Cout Cin sky130_fd_pr__cap_mim_m3_1 l=2e+06u w=2e+06u
X16 Cout Cin sky130_fd_pr__cap_mim_m3_1 l=2e+06u w=2e+06u
X17 Cout Cin sky130_fd_pr__cap_mim_m3_1 l=2e+06u w=2e+06u
X18 Cout Cin sky130_fd_pr__cap_mim_m3_1 l=2e+06u w=2e+06u
X19 Cout Cin sky130_fd_pr__cap_mim_m3_1 l=2e+06u w=2e+06u
C0 Cin Cout 28.31fF
C1 Cout VSUBS 2.81fF
C2 Cin VSUBS 6.38fF
C3 VGND VSUBS 6.63fF
C4 VPWR VSUBS 6.63fF
.ends

.subckt sky130_asc_pnp_05v5_W3p40L3p40_8 Emitter Base Collector VPWR VGND
X0 Collector Base Emitter sky130_fd_pr__pnp_05v5_W3p40L3p40
X1 Collector Base Emitter sky130_fd_pr__pnp_05v5_W3p40L3p40
X2 Collector Base Emitter sky130_fd_pr__pnp_05v5_W3p40L3p40
X3 Collector Base Emitter sky130_fd_pr__pnp_05v5_W3p40L3p40
X4 Collector Base Emitter sky130_fd_pr__pnp_05v5_W3p40L3p40
X5 Collector Base Emitter sky130_fd_pr__pnp_05v5_W3p40L3p40
X6 Collector Base Emitter sky130_fd_pr__pnp_05v5_W3p40L3p40
X7 Collector Base Emitter sky130_fd_pr__pnp_05v5_W3p40L3p40
C0 Base Emitter 21.50fF
C1 VGND Collector 11.20fF
C2 VPWR Collector 13.12fF
C3 Emitter Collector 10.49fF
C4 Base Collector 33.06fF
.ends

.subckt sky130_asc_nfet_01v8_lvt_1 GATE SOURCE DRAIN VPWR VGND
X0 SOURCE GATE DRAIN VGND sky130_fd_pr__nfet_01v8_lvt ad=1.16e+12p pd=8.58e+06u as=1.16e+12p ps=8.58e+06u w=4e+06u l=2e+06u
C0 SOURCE GATE 0.00fF
C1 SOURCE VPWR 0.17fF
C2 SOURCE DRAIN 0.01fF
C3 GATE DRAIN 0.18fF
C4 VPWR VGND 0.64fF
C5 SOURCE VGND 0.40fF
C6 DRAIN VGND 0.34fF
C7 GATE VGND 1.34fF
.ends

.subckt bgr_top porst va vb vbg VSS VDD
Xsky130_asc_res_xhigh_po_2p85_1_7 sky130_asc_res_xhigh_po_2p85_1_7/Rin sky130_asc_res_xhigh_po_2p85_1_6/Rin
+ VDD VSS sky130_asc_res_xhigh_po_2p85_1_7/a_2148_115# sky130_asc_res_xhigh_po_2p85_1
Xsky130_asc_res_xhigh_po_2p85_1_8 vbg sky130_asc_res_xhigh_po_2p85_1_7/Rin VDD VSS
+ sky130_asc_res_xhigh_po_2p85_1_8/a_2148_115# sky130_asc_res_xhigh_po_2p85_1
Xsky130_asc_res_xhigh_po_2p85_1_9 sky130_asc_res_xhigh_po_2p85_1_9/Rin sky130_asc_res_xhigh_po_2p85_2_0/Rin
+ VDD VSS sky130_asc_res_xhigh_po_2p85_1_9/a_2148_115# sky130_asc_res_xhigh_po_2p85_1
Xsky130_asc_pfet_01v8_lvt_60_0 sky130_asc_cap_mim_m3_1_4/Cout VDD vbg VSS VDD VSS
+ sky130_asc_pfet_01v8_lvt_60
Xsky130_asc_pfet_01v8_lvt_60_1 sky130_asc_cap_mim_m3_1_4/Cout VDD vb VSS VDD VSS sky130_asc_pfet_01v8_lvt_60
Xsky130_asc_pfet_01v8_lvt_60_2 sky130_asc_cap_mim_m3_1_4/Cout VDD va VSS VDD VSS sky130_asc_pfet_01v8_lvt_60
Xsky130_asc_res_xhigh_po_2p85_1_30 va sky130_asc_res_xhigh_po_2p85_1_29/Rin VDD VSS
+ sky130_asc_res_xhigh_po_2p85_1_30/a_2148_115# sky130_asc_res_xhigh_po_2p85_1
Xsky130_asc_res_xhigh_po_2p85_1_20 vb sky130_asc_res_xhigh_po_2p85_1_19/Rin VDD VSS
+ sky130_asc_res_xhigh_po_2p85_1_20/a_2148_115# sky130_asc_res_xhigh_po_2p85_1
Xsky130_asc_pnp_05v5_W3p40L3p40_7_0 sky130_asc_res_xhigh_po_2p85_1_19/Rout VSS VSS
+ VDD VSS sky130_asc_pnp_05v5_W3p40L3p40_7
Xsky130_asc_res_xhigh_po_2p85_1_21 sky130_asc_res_xhigh_po_2p85_1_21/Rin sky130_asc_res_xhigh_po_2p85_2_1/Rin
+ VDD VSS sky130_asc_res_xhigh_po_2p85_1_21/a_2148_115# sky130_asc_res_xhigh_po_2p85_1
Xsky130_asc_res_xhigh_po_2p85_1_10 sky130_asc_res_xhigh_po_2p85_1_10/Rin sky130_asc_res_xhigh_po_2p85_1_9/Rin
+ VDD VSS sky130_asc_res_xhigh_po_2p85_1_10/a_2148_115# sky130_asc_res_xhigh_po_2p85_1
Xsky130_asc_res_xhigh_po_2p85_2_0 sky130_asc_res_xhigh_po_2p85_2_0/Rin VSS VDD sky130_asc_res_xhigh_po_2p85_2_0/a_2723_115#
+ VSS sky130_asc_res_xhigh_po_2p85_2
Xsky130_asc_res_xhigh_po_2p85_1_22 sky130_asc_res_xhigh_po_2p85_1_22/Rin sky130_asc_res_xhigh_po_2p85_1_21/Rin
+ VDD VSS sky130_asc_res_xhigh_po_2p85_1_22/a_2148_115# sky130_asc_res_xhigh_po_2p85_1
Xsky130_asc_res_xhigh_po_2p85_1_11 sky130_asc_res_xhigh_po_2p85_1_11/Rin sky130_asc_res_xhigh_po_2p85_1_10/Rin
+ VDD VSS sky130_asc_res_xhigh_po_2p85_1_11/a_2148_115# sky130_asc_res_xhigh_po_2p85_1
Xsky130_asc_res_xhigh_po_2p85_2_1 sky130_asc_res_xhigh_po_2p85_2_1/Rin VSS VDD sky130_asc_res_xhigh_po_2p85_2_1/a_2723_115#
+ VSS sky130_asc_res_xhigh_po_2p85_2
Xsky130_asc_res_xhigh_po_2p85_1_12 sky130_asc_res_xhigh_po_2p85_1_12/Rin sky130_asc_res_xhigh_po_2p85_1_11/Rin
+ VDD VSS sky130_asc_res_xhigh_po_2p85_1_12/a_2148_115# sky130_asc_res_xhigh_po_2p85_1
Xsky130_asc_res_xhigh_po_2p85_1_23 sky130_asc_res_xhigh_po_2p85_1_23/Rin sky130_asc_res_xhigh_po_2p85_1_22/Rin
+ VDD VSS sky130_asc_res_xhigh_po_2p85_1_23/a_2148_115# sky130_asc_res_xhigh_po_2p85_1
Xsky130_asc_res_xhigh_po_2p85_1_24 sky130_asc_res_xhigh_po_2p85_1_24/Rin sky130_asc_res_xhigh_po_2p85_1_23/Rin
+ VDD VSS sky130_asc_res_xhigh_po_2p85_1_24/a_2148_115# sky130_asc_res_xhigh_po_2p85_1
Xsky130_asc_res_xhigh_po_2p85_1_13 sky130_asc_res_xhigh_po_2p85_1_13/Rin sky130_asc_res_xhigh_po_2p85_1_12/Rin
+ VDD VSS sky130_asc_res_xhigh_po_2p85_1_13/a_2148_115# sky130_asc_res_xhigh_po_2p85_1
Xsky130_asc_pfet_01v8_lvt_12_0 VDD VDD va VSS VDD VSS sky130_asc_pfet_01v8_lvt_12
Xsky130_asc_res_xhigh_po_2p85_1_25 sky130_asc_res_xhigh_po_2p85_1_25/Rin sky130_asc_res_xhigh_po_2p85_1_24/Rin
+ VDD VSS sky130_asc_res_xhigh_po_2p85_1_25/a_2148_115# sky130_asc_res_xhigh_po_2p85_1
Xsky130_asc_res_xhigh_po_2p85_1_14 sky130_asc_res_xhigh_po_2p85_1_14/Rin sky130_asc_res_xhigh_po_2p85_1_13/Rin
+ VDD VSS sky130_asc_res_xhigh_po_2p85_1_14/a_2148_115# sky130_asc_res_xhigh_po_2p85_1
Xsky130_asc_pfet_01v8_lvt_12_1 sky130_asc_cap_mim_m3_1_4/Cout VDD sky130_asc_nfet_01v8_lvt_1_1/GATE
+ VSS VDD VSS sky130_asc_pfet_01v8_lvt_12
Xsky130_asc_res_xhigh_po_2p85_1_15 sky130_asc_res_xhigh_po_2p85_1_15/Rin sky130_asc_res_xhigh_po_2p85_1_14/Rin
+ VDD VSS sky130_asc_res_xhigh_po_2p85_1_15/a_2148_115# sky130_asc_res_xhigh_po_2p85_1
Xsky130_asc_res_xhigh_po_2p85_1_26 sky130_asc_res_xhigh_po_2p85_1_26/Rin sky130_asc_res_xhigh_po_2p85_1_25/Rin
+ VDD VSS sky130_asc_res_xhigh_po_2p85_1_26/a_2148_115# sky130_asc_res_xhigh_po_2p85_1
Xsky130_asc_res_xhigh_po_2p85_1_16 sky130_asc_res_xhigh_po_2p85_1_18/Rin sky130_asc_res_xhigh_po_2p85_1_15/Rin
+ VDD VSS sky130_asc_res_xhigh_po_2p85_1_16/a_2148_115# sky130_asc_res_xhigh_po_2p85_1
Xsky130_asc_res_xhigh_po_2p85_1_27 sky130_asc_res_xhigh_po_2p85_1_27/Rin sky130_asc_res_xhigh_po_2p85_1_26/Rin
+ VDD VSS sky130_asc_res_xhigh_po_2p85_1_27/a_2148_115# sky130_asc_res_xhigh_po_2p85_1
Xsky130_asc_res_xhigh_po_2p85_1_17 sky130_asc_res_xhigh_po_2p85_1_17/Rin vb VDD VSS
+ sky130_asc_res_xhigh_po_2p85_1_17/a_2148_115# sky130_asc_res_xhigh_po_2p85_1
Xsky130_asc_res_xhigh_po_2p85_1_28 sky130_asc_res_xhigh_po_2p85_1_28/Rin sky130_asc_res_xhigh_po_2p85_1_27/Rin
+ VDD VSS sky130_asc_res_xhigh_po_2p85_1_28/a_2148_115# sky130_asc_res_xhigh_po_2p85_1
Xsky130_asc_nfet_01v8_lvt_9_0 porst VSS sky130_asc_cap_mim_m3_1_4/Cout VDD VSS sky130_asc_nfet_01v8_lvt_9
Xsky130_asc_res_xhigh_po_2p85_1_18 sky130_asc_res_xhigh_po_2p85_1_18/Rin sky130_asc_res_xhigh_po_2p85_1_17/Rin
+ VDD VSS sky130_asc_res_xhigh_po_2p85_1_18/a_2148_115# sky130_asc_res_xhigh_po_2p85_1
Xsky130_asc_res_xhigh_po_2p85_1_29 sky130_asc_res_xhigh_po_2p85_1_29/Rin sky130_asc_res_xhigh_po_2p85_1_28/Rin
+ VDD VSS sky130_asc_res_xhigh_po_2p85_1_29/a_2148_115# sky130_asc_res_xhigh_po_2p85_1
Xsky130_asc_pfet_01v8_lvt_6_0 sky130_asc_pfet_01v8_lvt_6_1/GATE VDD sky130_asc_cap_mim_m3_1_4/Cout
+ VSS VDD VSS sky130_asc_pfet_01v8_lvt_6
Xsky130_asc_nfet_01v8_lvt_9_1 va sky130_asc_nfet_01v8_lvt_1_1/DRAIN sky130_asc_cap_mim_m3_1_4/Cout
+ VDD VSS sky130_asc_nfet_01v8_lvt_9
Xsky130_asc_res_xhigh_po_2p85_1_19 sky130_asc_res_xhigh_po_2p85_1_19/Rin sky130_asc_res_xhigh_po_2p85_1_19/Rout
+ VDD VSS sky130_asc_res_xhigh_po_2p85_1_19/a_2148_115# sky130_asc_res_xhigh_po_2p85_1
Xsky130_asc_pfet_01v8_lvt_6_1 sky130_asc_pfet_01v8_lvt_6_1/GATE VDD sky130_asc_pfet_01v8_lvt_6_1/GATE
+ VSS VDD VSS sky130_asc_pfet_01v8_lvt_6
Xsky130_asc_pnp_05v5_W3p40L3p40_1_0 va VSS VSS VDD VSS sky130_asc_pnp_05v5_W3p40L3p40_1
Xsky130_asc_nfet_01v8_lvt_9_2 vb sky130_asc_nfet_01v8_lvt_1_1/DRAIN sky130_asc_pfet_01v8_lvt_6_1/GATE
+ VDD VSS sky130_asc_nfet_01v8_lvt_9
Xsky130_asc_cap_mim_m3_1_0 VDD sky130_asc_cap_mim_m3_1_4/Cout VDD VSS VSS sky130_asc_cap_mim_m3_1
Xsky130_asc_cap_mim_m3_1_1 VDD sky130_asc_cap_mim_m3_1_4/Cout VDD VSS VSS sky130_asc_cap_mim_m3_1
Xsky130_asc_pnp_05v5_W3p40L3p40_8_0 sky130_asc_res_xhigh_po_2p85_1_19/Rout VSS VSS
+ VDD VSS sky130_asc_pnp_05v5_W3p40L3p40_8
Xsky130_asc_cap_mim_m3_1_2 VDD sky130_asc_cap_mim_m3_1_4/Cout VDD VSS VSS sky130_asc_cap_mim_m3_1
Xsky130_asc_pnp_05v5_W3p40L3p40_8_1 sky130_asc_res_xhigh_po_2p85_1_19/Rout VSS VSS
+ VDD VSS sky130_asc_pnp_05v5_W3p40L3p40_8
Xsky130_asc_cap_mim_m3_1_3 VDD sky130_asc_cap_mim_m3_1_4/Cout VDD VSS VSS sky130_asc_cap_mim_m3_1
Xsky130_asc_pnp_05v5_W3p40L3p40_8_2 sky130_asc_res_xhigh_po_2p85_1_19/Rout VSS VSS
+ VDD VSS sky130_asc_pnp_05v5_W3p40L3p40_8
Xsky130_asc_cap_mim_m3_1_4 VDD sky130_asc_cap_mim_m3_1_4/Cout VDD VSS VSS sky130_asc_cap_mim_m3_1
Xsky130_asc_pnp_05v5_W3p40L3p40_8_3 sky130_asc_res_xhigh_po_2p85_1_19/Rout VSS VSS
+ VDD VSS sky130_asc_pnp_05v5_W3p40L3p40_8
Xsky130_asc_cap_mim_m3_1_5 va VSS VDD VSS VSS sky130_asc_cap_mim_m3_1
Xsky130_asc_res_xhigh_po_2p85_1_0 sky130_asc_res_xhigh_po_2p85_1_0/Rin VSS VDD VSS
+ sky130_asc_res_xhigh_po_2p85_1_0/a_2148_115# sky130_asc_res_xhigh_po_2p85_1
Xsky130_asc_cap_mim_m3_1_6 va VSS VDD VSS VSS sky130_asc_cap_mim_m3_1
Xsky130_asc_nfet_01v8_lvt_1_0 sky130_asc_nfet_01v8_lvt_1_1/GATE VSS sky130_asc_nfet_01v8_lvt_1_1/GATE
+ VDD VSS sky130_asc_nfet_01v8_lvt_1
Xsky130_asc_res_xhigh_po_2p85_1_1 sky130_asc_res_xhigh_po_2p85_1_1/Rin sky130_asc_res_xhigh_po_2p85_1_0/Rin
+ VDD VSS sky130_asc_res_xhigh_po_2p85_1_1/a_2148_115# sky130_asc_res_xhigh_po_2p85_1
Xsky130_asc_cap_mim_m3_1_7 va VSS VDD VSS VSS sky130_asc_cap_mim_m3_1
Xsky130_asc_nfet_01v8_lvt_1_1 sky130_asc_nfet_01v8_lvt_1_1/GATE VSS sky130_asc_nfet_01v8_lvt_1_1/DRAIN
+ VDD VSS sky130_asc_nfet_01v8_lvt_1
Xsky130_asc_res_xhigh_po_2p85_1_2 sky130_asc_res_xhigh_po_2p85_1_2/Rin sky130_asc_res_xhigh_po_2p85_1_1/Rin
+ VDD VSS sky130_asc_res_xhigh_po_2p85_1_2/a_2148_115# sky130_asc_res_xhigh_po_2p85_1
Xsky130_asc_cap_mim_m3_1_8 va VSS VDD VSS VSS sky130_asc_cap_mim_m3_1
Xsky130_asc_res_xhigh_po_2p85_1_3 sky130_asc_res_xhigh_po_2p85_1_3/Rin sky130_asc_res_xhigh_po_2p85_1_2/Rin
+ VDD VSS sky130_asc_res_xhigh_po_2p85_1_3/a_2148_115# sky130_asc_res_xhigh_po_2p85_1
Xsky130_asc_cap_mim_m3_1_9 va VSS VDD VSS VSS sky130_asc_cap_mim_m3_1
Xsky130_asc_res_xhigh_po_2p85_1_4 sky130_asc_res_xhigh_po_2p85_1_4/Rin sky130_asc_res_xhigh_po_2p85_1_3/Rin
+ VDD VSS sky130_asc_res_xhigh_po_2p85_1_4/a_2148_115# sky130_asc_res_xhigh_po_2p85_1
Xsky130_asc_res_xhigh_po_2p85_1_5 sky130_asc_res_xhigh_po_2p85_1_5/Rin sky130_asc_res_xhigh_po_2p85_1_4/Rin
+ VDD VSS sky130_asc_res_xhigh_po_2p85_1_5/a_2148_115# sky130_asc_res_xhigh_po_2p85_1
Xsky130_asc_res_xhigh_po_2p85_1_6 sky130_asc_res_xhigh_po_2p85_1_6/Rin sky130_asc_res_xhigh_po_2p85_1_5/Rin
+ VDD VSS sky130_asc_res_xhigh_po_2p85_1_6/a_2148_115# sky130_asc_res_xhigh_po_2p85_1
C0 sky130_asc_res_xhigh_po_2p85_1_8/a_2148_115# sky130_asc_res_xhigh_po_2p85_1_7/Rin 0.45fF
C1 sky130_asc_res_xhigh_po_2p85_1_22/Rin VDD 0.93fF
C2 sky130_asc_nfet_01v8_lvt_1_1/DRAIN VDD 2.65fF
C3 VDD sky130_asc_res_xhigh_po_2p85_1_5/Rin -0.12fF
C4 sky130_asc_res_xhigh_po_2p85_1_22/a_2148_115# sky130_asc_res_xhigh_po_2p85_1_23/Rin 0.20fF
C5 sky130_asc_res_xhigh_po_2p85_1_24/a_2148_115# sky130_asc_res_xhigh_po_2p85_1_10/Rin 0.20fF
C6 sky130_asc_cap_mim_m3_1_4/Cout VDD 3.00fF
C7 sky130_asc_res_xhigh_po_2p85_1_5/Rin sky130_asc_res_xhigh_po_2p85_1_7/Rin 0.11fF
C8 sky130_asc_res_xhigh_po_2p85_1_24/Rin sky130_asc_res_xhigh_po_2p85_1_18/Rin 0.25fF
C9 sky130_asc_res_xhigh_po_2p85_1_11/Rin sky130_asc_res_xhigh_po_2p85_1_10/Rin 0.53fF
C10 sky130_asc_res_xhigh_po_2p85_1_14/Rin sky130_asc_res_xhigh_po_2p85_1_9/Rin 0.03fF
C11 sky130_asc_res_xhigh_po_2p85_1_3/Rin sky130_asc_res_xhigh_po_2p85_1_0/a_2148_115# 0.29fF
C12 vbg VDD 1.93fF
C13 sky130_asc_res_xhigh_po_2p85_1_3/Rin sky130_asc_res_xhigh_po_2p85_1_2/Rin 0.46fF
C14 sky130_asc_res_xhigh_po_2p85_1_27/Rin VDD 0.13fF
C15 sky130_asc_cap_mim_m3_1_4/Cout porst 0.00fF
C16 vbg sky130_asc_res_xhigh_po_2p85_1_7/Rin 0.03fF
C17 sky130_asc_res_xhigh_po_2p85_1_26/a_2148_115# sky130_asc_res_xhigh_po_2p85_1_27/Rin 0.20fF
C18 sky130_asc_res_xhigh_po_2p85_1_22/Rin sky130_asc_res_xhigh_po_2p85_1_21/Rin 0.06fF
C19 sky130_asc_res_xhigh_po_2p85_1_13/Rin sky130_asc_res_xhigh_po_2p85_2_0/a_2723_115# 0.47fF
C20 sky130_asc_res_xhigh_po_2p85_2_1/Rin sky130_asc_cap_mim_m3_1_4/Cout -0.10fF
C21 VDD sky130_asc_res_xhigh_po_2p85_1_29/Rin 0.11fF
C22 sky130_asc_res_xhigh_po_2p85_1_24/Rin VDD 5.52fF
C23 VDD sky130_asc_res_xhigh_po_2p85_1_10/Rin 0.11fF
C24 sky130_asc_res_xhigh_po_2p85_1_24/Rin sky130_asc_res_xhigh_po_2p85_1_15/Rin 0.01fF
C25 sky130_asc_res_xhigh_po_2p85_1_14/Rin sky130_asc_res_xhigh_po_2p85_2_0/Rin 0.03fF
C26 sky130_asc_cap_mim_m3_1_4/Cout sky130_asc_res_xhigh_po_2p85_1_21/Rin 0.14fF
C27 sky130_asc_res_xhigh_po_2p85_1_17/Rin VDD 2.87fF
C28 sky130_asc_res_xhigh_po_2p85_1_19/a_2148_115# sky130_asc_res_xhigh_po_2p85_1_19/Rin 0.54fF
C29 sky130_asc_res_xhigh_po_2p85_1_14/a_2148_115# sky130_asc_res_xhigh_po_2p85_1_23/Rin 0.20fF
C30 sky130_asc_res_xhigh_po_2p85_1_0/a_2148_115# vbg 0.20fF
C31 sky130_asc_pfet_01v8_lvt_6_1/GATE sky130_asc_nfet_01v8_lvt_1_1/DRAIN 0.23fF
C32 sky130_asc_pfet_01v8_lvt_6_1/GATE sky130_asc_cap_mim_m3_1_4/Cout 0.08fF
C33 sky130_asc_res_xhigh_po_2p85_1_26/Rin VDD 0.97fF
C34 sky130_asc_res_xhigh_po_2p85_1_28/Rin sky130_asc_res_xhigh_po_2p85_1_23/a_2148_115# 0.20fF
C35 sky130_asc_res_xhigh_po_2p85_1_17/a_2148_115# sky130_asc_res_xhigh_po_2p85_1_17/Rin 0.23fF
C36 sky130_asc_res_xhigh_po_2p85_1_26/Rin sky130_asc_res_xhigh_po_2p85_1_26/a_2148_115# 0.62fF
C37 sky130_asc_res_xhigh_po_2p85_1_23/a_2148_115# sky130_asc_res_xhigh_po_2p85_1_21/Rin 0.06fF
C38 sky130_asc_nfet_01v8_lvt_1_1/DRAIN vb 0.98fF
C39 sky130_asc_res_xhigh_po_2p85_1_14/Rin sky130_asc_res_xhigh_po_2p85_1_24/Rin 0.03fF
C40 sky130_asc_res_xhigh_po_2p85_1_14/Rin sky130_asc_res_xhigh_po_2p85_1_10/Rin 0.03fF
C41 sky130_asc_res_xhigh_po_2p85_1_8/a_2148_115# sky130_asc_res_xhigh_po_2p85_1_6/Rin 0.20fF
C42 sky130_asc_res_xhigh_po_2p85_1_4/Rin sky130_asc_res_xhigh_po_2p85_1_3/Rin 1.17fF
C43 sky130_asc_cap_mim_m3_1_4/Cout vb 0.23fF
C44 sky130_asc_res_xhigh_po_2p85_1_12/Rin sky130_asc_res_xhigh_po_2p85_1_18/Rin 0.38fF
C45 sky130_asc_res_xhigh_po_2p85_1_4/Rin sky130_asc_res_xhigh_po_2p85_1_0/Rin 0.35fF
C46 sky130_asc_res_xhigh_po_2p85_1_9/a_2148_115# sky130_asc_res_xhigh_po_2p85_1_11/Rin 0.20fF
C47 sky130_asc_res_xhigh_po_2p85_1_11/Rin sky130_asc_res_xhigh_po_2p85_1_12/Rin 1.56fF
C48 sky130_asc_res_xhigh_po_2p85_1_22/a_2148_115# sky130_asc_res_xhigh_po_2p85_1_21/Rin 0.14fF
C49 sky130_asc_res_xhigh_po_2p85_1_4/Rin sky130_asc_res_xhigh_po_2p85_1_5/Rin 0.55fF
C50 VDD sky130_asc_res_xhigh_po_2p85_1_23/Rin 3.93fF
C51 sky130_asc_res_xhigh_po_2p85_1_29/a_2148_115# sky130_asc_res_xhigh_po_2p85_1_21/Rin 1.25fF
C52 sky130_asc_res_xhigh_po_2p85_1_19/a_2148_115# vb 0.20fF
C53 sky130_asc_res_xhigh_po_2p85_1_9/Rin sky130_asc_res_xhigh_po_2p85_2_0/Rin 0.72fF
C54 sky130_asc_nfet_01v8_lvt_1_1/GATE sky130_asc_nfet_01v8_lvt_1_1/DRAIN 0.15fF
C55 sky130_asc_res_xhigh_po_2p85_1_12/Rin VDD 0.32fF
C56 sky130_asc_res_xhigh_po_2p85_1_11/Rin sky130_asc_res_xhigh_po_2p85_1_18/Rin 0.03fF
C57 sky130_asc_res_xhigh_po_2p85_1_24/Rin vb 0.03fF
C58 sky130_asc_res_xhigh_po_2p85_1_12/Rin sky130_asc_res_xhigh_po_2p85_1_15/Rin 0.09fF
C59 sky130_asc_res_xhigh_po_2p85_1_4/Rin vbg 0.05fF
C60 sky130_asc_nfet_01v8_lvt_1_1/GATE sky130_asc_cap_mim_m3_1_4/Cout -0.10fF
C61 sky130_asc_res_xhigh_po_2p85_1_17/Rin vb 0.49fF
C62 sky130_asc_res_xhigh_po_2p85_1_1/Rin VDD 0.24fF
C63 sky130_asc_res_xhigh_po_2p85_1_3/Rin sky130_asc_res_xhigh_po_2p85_1_5/Rin 1.98fF
C64 sky130_asc_res_xhigh_po_2p85_1_8/a_2148_115# sky130_asc_res_xhigh_po_2p85_1_5/Rin 0.36fF
C65 sky130_asc_res_xhigh_po_2p85_1_4/Rin sky130_asc_res_xhigh_po_2p85_1_1/a_2148_115# 0.21fF
C66 sky130_asc_res_xhigh_po_2p85_1_1/Rin sky130_asc_res_xhigh_po_2p85_1_3/a_2148_115# 0.32fF
C67 sky130_asc_res_xhigh_po_2p85_2_0/Rin sky130_asc_nfet_01v8_lvt_1_1/DRAIN 0.12fF
C68 sky130_asc_res_xhigh_po_2p85_1_18/Rin VDD 4.14fF
C69 va VDD 3.41fF
C70 sky130_asc_res_xhigh_po_2p85_1_15/a_2148_115# sky130_asc_res_xhigh_po_2p85_1_17/Rin 0.26fF
C71 sky130_asc_res_xhigh_po_2p85_1_23/Rin sky130_asc_res_xhigh_po_2p85_1_21/Rin 0.03fF
C72 sky130_asc_res_xhigh_po_2p85_1_18/Rin sky130_asc_res_xhigh_po_2p85_1_15/Rin 1.10fF
C73 sky130_asc_res_xhigh_po_2p85_1_11/Rin VDD 0.11fF
C74 sky130_asc_res_xhigh_po_2p85_1_11/Rin sky130_asc_res_xhigh_po_2p85_1_15/Rin 0.03fF
C75 sky130_asc_res_xhigh_po_2p85_1_3/Rin vbg 0.45fF
C76 sky130_asc_nfet_01v8_lvt_1_1/DRAIN sky130_asc_cap_mim_m3_1_4/Cout 0.12fF
C77 sky130_asc_res_xhigh_po_2p85_1_14/Rin sky130_asc_res_xhigh_po_2p85_1_23/Rin 0.42fF
C78 sky130_asc_res_xhigh_po_2p85_1_9/Rin sky130_asc_res_xhigh_po_2p85_1_24/Rin 0.03fF
C79 sky130_asc_res_xhigh_po_2p85_1_27/a_2148_115# sky130_asc_res_xhigh_po_2p85_1_9/Rin 0.20fF
C80 sky130_asc_res_xhigh_po_2p85_1_9/Rin sky130_asc_res_xhigh_po_2p85_1_10/Rin 0.59fF
C81 sky130_asc_res_xhigh_po_2p85_1_5/a_2148_115# sky130_asc_res_xhigh_po_2p85_1_7/Rin 0.25fF
C82 sky130_asc_res_xhigh_po_2p85_1_13/Rin VDD 1.98fF
C83 sky130_asc_res_xhigh_po_2p85_1_27/Rin sky130_asc_res_xhigh_po_2p85_1_25/Rin 0.03fF
C84 sky130_asc_res_xhigh_po_2p85_1_14/Rin sky130_asc_res_xhigh_po_2p85_1_12/Rin 0.03fF
C85 sky130_asc_res_xhigh_po_2p85_1_12/a_2148_115# sky130_asc_res_xhigh_po_2p85_1_18/Rin 0.28fF
C86 vbg sky130_asc_res_xhigh_po_2p85_1_5/Rin 0.33fF
C87 sky130_asc_res_xhigh_po_2p85_1_15/Rin VDD 4.23fF
C88 vbg sky130_asc_cap_mim_m3_1_4/Cout 1.01fF
C89 sky130_asc_res_xhigh_po_2p85_1_27/Rin sky130_asc_cap_mim_m3_1_4/Cout 0.02fF
C90 VDD sky130_asc_res_xhigh_po_2p85_1_7/Rin 0.11fF
C91 sky130_asc_res_xhigh_po_2p85_1_27/a_2148_115# sky130_asc_res_xhigh_po_2p85_2_0/Rin 0.20fF
C92 sky130_asc_res_xhigh_po_2p85_1_1/a_2148_115# sky130_asc_res_xhigh_po_2p85_1_5/Rin 0.20fF
C93 sky130_asc_res_xhigh_po_2p85_1_4/Rin sky130_asc_res_xhigh_po_2p85_1_4/a_2148_115# 0.36fF
C94 sky130_asc_res_xhigh_po_2p85_1_19/Rin VDD 0.68fF
C95 sky130_asc_res_xhigh_po_2p85_1_14/Rin sky130_asc_res_xhigh_po_2p85_1_18/Rin 0.03fF
C96 porst VDD 1.76fF
C97 sky130_asc_res_xhigh_po_2p85_1_23/Rin vb 0.03fF
C98 sky130_asc_res_xhigh_po_2p85_1_12/a_2148_115# sky130_asc_res_xhigh_po_2p85_1_15/Rin 0.28fF
C99 sky130_asc_res_xhigh_po_2p85_2_1/Rin VDD 1.13fF
C100 sky130_asc_res_xhigh_po_2p85_1_28/Rin VDD 0.11fF
C101 sky130_asc_res_xhigh_po_2p85_1_13/Rin sky130_asc_res_xhigh_po_2p85_1_14/Rin 0.21fF
C102 VDD sky130_asc_res_xhigh_po_2p85_1_21/Rin 0.99fF
C103 sky130_asc_res_xhigh_po_2p85_1_22/a_2148_115# sky130_asc_res_xhigh_po_2p85_1_22/Rin 0.68fF
C104 sky130_asc_res_xhigh_po_2p85_1_3/Rin sky130_asc_res_xhigh_po_2p85_1_4/a_2148_115# 0.33fF
C105 sky130_asc_res_xhigh_po_2p85_1_0/a_2148_115# sky130_asc_res_xhigh_po_2p85_1_7/Rin 0.20fF
C106 sky130_asc_res_xhigh_po_2p85_1_14/Rin VDD 0.21fF
C107 sky130_asc_res_xhigh_po_2p85_1_14/Rin sky130_asc_res_xhigh_po_2p85_1_15/Rin 0.45fF
C108 sky130_asc_res_xhigh_po_2p85_1_4/a_2148_115# sky130_asc_res_xhigh_po_2p85_1_0/Rin 0.20fF
C109 sky130_asc_res_xhigh_po_2p85_1_2/Rin sky130_asc_res_xhigh_po_2p85_1_3/a_2148_115# 0.70fF
C110 sky130_asc_res_xhigh_po_2p85_1_23/a_2148_115# sky130_asc_res_xhigh_po_2p85_1_29/Rin 0.20fF
C111 va vb 0.04fF
C112 sky130_asc_res_xhigh_po_2p85_1_9/Rin sky130_asc_res_xhigh_po_2p85_1_23/Rin 0.14fF
C113 sky130_asc_pfet_01v8_lvt_6_1/GATE VDD 0.46fF
C114 sky130_asc_res_xhigh_po_2p85_1_16/a_2148_115# sky130_asc_res_xhigh_po_2p85_1_12/Rin 0.20fF
C115 sky130_asc_res_xhigh_po_2p85_2_1/Rin sky130_asc_res_xhigh_po_2p85_1_21/Rin 0.03fF
C116 sky130_asc_res_xhigh_po_2p85_1_14/a_2148_115# sky130_asc_res_xhigh_po_2p85_1_9/Rin 0.02fF
C117 sky130_asc_res_xhigh_po_2p85_1_28/Rin sky130_asc_res_xhigh_po_2p85_1_21/Rin 0.10fF
C118 sky130_asc_res_xhigh_po_2p85_1_25/a_2148_115# sky130_asc_res_xhigh_po_2p85_1_24/Rin 0.09fF
C119 sky130_asc_res_xhigh_po_2p85_1_9/Rin sky130_asc_res_xhigh_po_2p85_1_12/Rin 0.03fF
C120 sky130_asc_res_xhigh_po_2p85_1_14/Rin sky130_asc_res_xhigh_po_2p85_1_12/a_2148_115# 0.20fF
C121 sky130_asc_res_xhigh_po_2p85_1_26/Rin sky130_asc_res_xhigh_po_2p85_1_27/Rin 0.56fF
C122 sky130_asc_res_xhigh_po_2p85_1_13/Rin vb 3.88fF
C123 sky130_asc_res_xhigh_po_2p85_1_5/a_2148_115# sky130_asc_res_xhigh_po_2p85_1_6/Rin 0.20fF
C124 sky130_asc_res_xhigh_po_2p85_1_15/a_2148_115# sky130_asc_res_xhigh_po_2p85_1_18/Rin 0.53fF
C125 sky130_asc_res_xhigh_po_2p85_2_0/Rin sky130_asc_res_xhigh_po_2p85_1_23/Rin 0.03fF
C126 VDD vb 3.15fF
C127 sky130_asc_res_xhigh_po_2p85_1_3/Rin sky130_asc_res_xhigh_po_2p85_1_1/Rin 0.03fF
C128 sky130_asc_res_xhigh_po_2p85_1_16/a_2148_115# sky130_asc_res_xhigh_po_2p85_1_18/Rin 0.28fF
C129 sky130_asc_res_xhigh_po_2p85_1_9/Rin sky130_asc_res_xhigh_po_2p85_1_24/a_2148_115# 0.29fF
C130 va sky130_asc_nfet_01v8_lvt_1_1/GATE 0.04fF
C131 sky130_asc_res_xhigh_po_2p85_1_16/a_2148_115# sky130_asc_res_xhigh_po_2p85_1_11/Rin 0.20fF
C132 sky130_asc_res_xhigh_po_2p85_2_1/Rin sky130_asc_res_xhigh_po_2p85_1_30/a_2148_115# 0.09fF
C133 sky130_asc_cap_mim_m3_1_4/Cout sky130_asc_res_xhigh_po_2p85_1_23/Rin 0.02fF
C134 VDD sky130_asc_res_xhigh_po_2p85_1_6/Rin 0.11fF
C135 sky130_asc_res_xhigh_po_2p85_1_19/Rin vb 0.60fF
C136 sky130_asc_res_xhigh_po_2p85_1_4/Rin VDD 2.19fF
C137 sky130_asc_res_xhigh_po_2p85_1_7/Rin sky130_asc_res_xhigh_po_2p85_1_6/Rin 0.48fF
C138 sky130_asc_nfet_01v8_lvt_1_1/GATE VDD 0.01fF
C139 sky130_asc_res_xhigh_po_2p85_1_16/a_2148_115# sky130_asc_res_xhigh_po_2p85_1_15/Rin 0.08fF
C140 sky130_asc_res_xhigh_po_2p85_1_19/Rout VDD 0.53fF
C141 sky130_asc_res_xhigh_po_2p85_1_9/Rin VDD 0.11fF
C142 va sky130_asc_nfet_01v8_lvt_1_1/DRAIN 0.06fF
C143 sky130_asc_res_xhigh_po_2p85_1_23/Rin sky130_asc_res_xhigh_po_2p85_1_29/Rin 0.03fF
C144 sky130_asc_res_xhigh_po_2p85_1_24/Rin sky130_asc_res_xhigh_po_2p85_1_23/Rin 1.91fF
C145 sky130_asc_res_xhigh_po_2p85_1_14/Rin vb 2.02fF
C146 sky130_asc_res_xhigh_po_2p85_1_14/a_2148_115# sky130_asc_res_xhigh_po_2p85_1_24/Rin 0.20fF
C147 va sky130_asc_cap_mim_m3_1_4/Cout 4.38fF
C148 sky130_asc_res_xhigh_po_2p85_1_13/Rin sky130_asc_res_xhigh_po_2p85_2_0/Rin 0.69fF
C149 sky130_asc_res_xhigh_po_2p85_1_3/Rin VDD 0.21fF
C150 sky130_asc_res_xhigh_po_2p85_1_9/a_2148_115# sky130_asc_res_xhigh_po_2p85_1_10/Rin 0.20fF
C151 sky130_asc_res_xhigh_po_2p85_2_1/Rin sky130_asc_res_xhigh_po_2p85_2_1/a_2723_115# 0.06fF
C152 sky130_asc_res_xhigh_po_2p85_1_19/Rout sky130_asc_res_xhigh_po_2p85_1_19/Rin 0.45fF
C153 sky130_asc_res_xhigh_po_2p85_1_13/Rin sky130_asc_nfet_01v8_lvt_1_1/DRAIN 0.06fF
C154 VDD sky130_asc_res_xhigh_po_2p85_1_25/Rin 0.11fF
C155 sky130_asc_res_xhigh_po_2p85_1_0/Rin VDD 0.11fF
C156 sky130_asc_res_xhigh_po_2p85_1_4/Rin sky130_asc_res_xhigh_po_2p85_1_0/a_2148_115# 0.31fF
C157 sky130_asc_res_xhigh_po_2p85_1_3/Rin sky130_asc_res_xhigh_po_2p85_1_7/Rin 0.60fF
C158 sky130_asc_res_xhigh_po_2p85_2_0/a_2723_115# sky130_asc_res_xhigh_po_2p85_1_12/Rin 0.20fF
C159 sky130_asc_res_xhigh_po_2p85_2_0/Rin VDD 0.21fF
C160 sky130_asc_pfet_01v8_lvt_6_1/GATE vb -0.07fF
C161 VDD VSS 1039.96fF
C162 porst VSS 17.65fF
C163 sky130_asc_res_xhigh_po_2p85_1_6/Rin VSS 2.91fF
C164 sky130_asc_res_xhigh_po_2p85_1_5/Rin VSS 5.78fF
C165 sky130_asc_res_xhigh_po_2p85_1_0/Rin VSS 2.75fF
C166 sky130_asc_res_xhigh_po_2p85_1_19/Rout VSS 58.63fF
C167 sky130_asc_res_xhigh_po_2p85_1_11/Rin VSS 2.70fF
C168 sky130_asc_res_xhigh_po_2p85_1_9/Rin VSS 5.79fF
C169 vb VSS 39.34fF
C170 sky130_asc_res_xhigh_po_2p85_1_25/Rin VSS 2.91fF
C171 sky130_asc_res_xhigh_po_2p85_1_26/Rin VSS 4.12fF
C172 sky130_asc_res_xhigh_po_2p85_1_14/Rin VSS 7.17fF
C173 sky130_asc_res_xhigh_po_2p85_1_28/Rin VSS 2.95fF
C174 sky130_asc_res_xhigh_po_2p85_1_21/Rin VSS 9.19fF
C175 sky130_asc_res_xhigh_po_2p85_1_29/Rin VSS 3.55fF
C176 sky130_asc_res_xhigh_po_2p85_1_23/Rin VSS 4.76fF
C177 sky130_asc_res_xhigh_po_2p85_2_1/Rin VSS 4.37fF
C178 sky130_asc_nfet_01v8_lvt_1_1/DRAIN VSS 8.91fF
C179 sky130_asc_res_xhigh_po_2p85_1_6/a_2148_115# VSS 2.70fF
C180 sky130_asc_res_xhigh_po_2p85_1_5/a_2148_115# VSS 2.70fF
C181 sky130_asc_res_xhigh_po_2p85_1_3/Rin VSS 5.58fF
C182 sky130_asc_res_xhigh_po_2p85_1_4/Rin VSS 3.34fF
C183 sky130_asc_res_xhigh_po_2p85_1_4/a_2148_115# VSS 2.90fF
C184 sky130_asc_res_xhigh_po_2p85_1_2/Rin VSS 3.25fF
C185 sky130_asc_res_xhigh_po_2p85_1_3/a_2148_115# VSS 2.70fF
C186 sky130_asc_res_xhigh_po_2p85_1_2/a_2148_115# VSS 2.70fF
C187 sky130_asc_res_xhigh_po_2p85_1_1/Rin VSS 5.40fF
C188 sky130_asc_res_xhigh_po_2p85_1_1/a_2148_115# VSS 2.70fF
C189 sky130_asc_nfet_01v8_lvt_1_1/GATE VSS 6.59fF
C190 sky130_asc_res_xhigh_po_2p85_1_0/a_2148_115# VSS 2.70fF
C191 sky130_asc_pfet_01v8_lvt_6_1/GATE VSS 11.29fF
C192 sky130_asc_res_xhigh_po_2p85_1_19/a_2148_115# VSS 2.70fF
C193 sky130_asc_res_xhigh_po_2p85_1_29/a_2148_115# VSS 2.70fF
C194 sky130_asc_res_xhigh_po_2p85_1_18/a_2148_115# VSS 2.70fF
C195 sky130_asc_res_xhigh_po_2p85_1_27/Rin VSS 5.23fF
C196 sky130_asc_res_xhigh_po_2p85_1_28/a_2148_115# VSS 2.70fF
C197 sky130_asc_res_xhigh_po_2p85_1_17/Rin VSS 4.79fF
C198 sky130_asc_res_xhigh_po_2p85_1_17/a_2148_115# VSS 2.70fF
C199 sky130_asc_res_xhigh_po_2p85_1_27/a_2148_115# VSS 2.70fF
C200 sky130_asc_res_xhigh_po_2p85_1_15/Rin VSS 4.73fF
C201 sky130_asc_res_xhigh_po_2p85_1_18/Rin VSS 2.83fF
C202 sky130_asc_res_xhigh_po_2p85_1_16/a_2148_115# VSS 2.70fF
C203 sky130_asc_res_xhigh_po_2p85_1_26/a_2148_115# VSS 2.70fF
C204 sky130_asc_res_xhigh_po_2p85_1_15/a_2148_115# VSS 2.70fF
C205 sky130_asc_res_xhigh_po_2p85_1_13/Rin VSS 5.15fF
C206 sky130_asc_res_xhigh_po_2p85_1_14/a_2148_115# VSS 2.70fF
C207 sky130_asc_res_xhigh_po_2p85_1_24/Rin VSS 6.72fF
C208 sky130_asc_res_xhigh_po_2p85_1_25/a_2148_115# VSS 2.70fF
C209 va VSS 73.00fF
C210 sky130_asc_res_xhigh_po_2p85_1_13/a_2148_115# VSS 2.70fF
C211 sky130_asc_res_xhigh_po_2p85_1_24/a_2148_115# VSS 2.70fF
C212 sky130_asc_res_xhigh_po_2p85_1_22/Rin VSS 4.15fF
C213 sky130_asc_res_xhigh_po_2p85_1_23/a_2148_115# VSS 2.70fF
C214 sky130_asc_res_xhigh_po_2p85_1_12/Rin VSS 4.35fF
C215 sky130_asc_res_xhigh_po_2p85_1_12/a_2148_115# VSS 2.70fF
C216 sky130_asc_res_xhigh_po_2p85_2_1/a_2723_115# VSS 2.70fF
C217 sky130_asc_res_xhigh_po_2p85_1_10/Rin VSS 3.17fF
C218 sky130_asc_res_xhigh_po_2p85_1_11/a_2148_115# VSS 2.70fF
C219 sky130_asc_res_xhigh_po_2p85_1_22/a_2148_115# VSS 2.70fF
C220 sky130_asc_res_xhigh_po_2p85_2_0/a_2723_115# VSS 2.70fF
C221 sky130_asc_res_xhigh_po_2p85_1_10/a_2148_115# VSS 2.70fF
C222 sky130_asc_res_xhigh_po_2p85_1_21/a_2148_115# VSS 2.70fF
C223 sky130_asc_res_xhigh_po_2p85_1_19/Rin VSS 3.69fF
C224 sky130_asc_res_xhigh_po_2p85_1_20/a_2148_115# VSS 2.70fF
C225 sky130_asc_res_xhigh_po_2p85_1_30/a_2148_115# VSS 2.70fF
C226 vbg VSS 16.97fF
C227 sky130_asc_cap_mim_m3_1_4/Cout VSS 132.21fF
C228 sky130_asc_res_xhigh_po_2p85_2_0/Rin VSS 3.38fF
C229 sky130_asc_res_xhigh_po_2p85_1_9/a_2148_115# VSS 2.70fF
C230 sky130_asc_res_xhigh_po_2p85_1_7/Rin VSS 4.29fF
C231 sky130_asc_res_xhigh_po_2p85_1_8/a_2148_115# VSS 2.70fF
C232 sky130_asc_res_xhigh_po_2p85_1_7/a_2148_115# VSS 2.70fF
.ends

