magic
tech sky130A
magscale 1 2
timestamp 1658609783
<< nwell >>
rect 130 1707 27740 1940
rect 130 1000 27741 1707
rect 131 293 27741 1000
<< pmoslvt >>
rect 225 355 625 1645
rect 683 355 1083 1645
rect 1141 355 1541 1645
rect 1599 355 1999 1645
rect 2057 355 2457 1645
rect 2515 355 2915 1645
rect 2973 355 3373 1645
rect 3431 355 3831 1645
rect 3889 355 4289 1645
rect 4347 355 4747 1645
rect 4805 355 5205 1645
rect 5263 355 5663 1645
rect 5721 355 6121 1645
rect 6179 355 6579 1645
rect 6637 355 7037 1645
rect 7095 355 7495 1645
rect 7553 355 7953 1645
rect 8011 355 8411 1645
rect 8469 355 8869 1645
rect 8927 355 9327 1645
rect 9385 355 9785 1645
rect 9843 355 10243 1645
rect 10301 355 10701 1645
rect 10759 355 11159 1645
rect 11217 355 11617 1645
rect 11675 355 12075 1645
rect 12133 355 12533 1645
rect 12591 355 12991 1645
rect 13049 355 13449 1645
rect 13507 355 13907 1645
rect 13965 355 14365 1645
rect 14423 355 14823 1645
rect 14881 355 15281 1645
rect 15339 355 15739 1645
rect 15797 355 16197 1645
rect 16255 355 16655 1645
rect 16713 355 17113 1645
rect 17171 355 17571 1645
rect 17629 355 18029 1645
rect 18087 355 18487 1645
rect 18545 355 18945 1645
rect 19003 355 19403 1645
rect 19461 355 19861 1645
rect 19919 355 20319 1645
rect 20377 355 20777 1645
rect 20835 355 21235 1645
rect 21293 355 21693 1645
rect 21751 355 22151 1645
rect 22209 355 22609 1645
rect 22667 355 23067 1645
rect 23125 355 23525 1645
rect 23583 355 23983 1645
rect 24041 355 24441 1645
rect 24499 355 24899 1645
rect 24957 355 25357 1645
rect 25415 355 25815 1645
rect 25873 355 26273 1645
rect 26331 355 26731 1645
rect 26789 355 27189 1645
rect 27247 355 27647 1645
<< pdiff >>
rect 167 1633 225 1645
rect 167 367 179 1633
rect 213 367 225 1633
rect 167 355 225 367
rect 625 1633 683 1645
rect 625 367 637 1633
rect 671 367 683 1633
rect 625 355 683 367
rect 1083 1633 1141 1645
rect 1083 367 1095 1633
rect 1129 367 1141 1633
rect 1083 355 1141 367
rect 1541 1633 1599 1645
rect 1541 367 1553 1633
rect 1587 367 1599 1633
rect 1541 355 1599 367
rect 1999 1633 2057 1645
rect 1999 367 2011 1633
rect 2045 367 2057 1633
rect 1999 355 2057 367
rect 2457 1633 2515 1645
rect 2457 367 2469 1633
rect 2503 367 2515 1633
rect 2457 355 2515 367
rect 2915 1633 2973 1645
rect 2915 367 2927 1633
rect 2961 367 2973 1633
rect 2915 355 2973 367
rect 3373 1633 3431 1645
rect 3373 367 3385 1633
rect 3419 367 3431 1633
rect 3373 355 3431 367
rect 3831 1633 3889 1645
rect 3831 367 3843 1633
rect 3877 367 3889 1633
rect 3831 355 3889 367
rect 4289 1633 4347 1645
rect 4289 367 4301 1633
rect 4335 367 4347 1633
rect 4289 355 4347 367
rect 4747 1633 4805 1645
rect 4747 367 4759 1633
rect 4793 367 4805 1633
rect 4747 355 4805 367
rect 5205 1633 5263 1645
rect 5205 367 5217 1633
rect 5251 367 5263 1633
rect 5205 355 5263 367
rect 5663 1633 5721 1645
rect 5663 367 5675 1633
rect 5709 367 5721 1633
rect 5663 355 5721 367
rect 6121 1633 6179 1645
rect 6121 367 6133 1633
rect 6167 367 6179 1633
rect 6121 355 6179 367
rect 6579 1633 6637 1645
rect 6579 367 6591 1633
rect 6625 367 6637 1633
rect 6579 355 6637 367
rect 7037 1633 7095 1645
rect 7037 367 7049 1633
rect 7083 367 7095 1633
rect 7037 355 7095 367
rect 7495 1633 7553 1645
rect 7495 367 7507 1633
rect 7541 367 7553 1633
rect 7495 355 7553 367
rect 7953 1633 8011 1645
rect 7953 367 7965 1633
rect 7999 367 8011 1633
rect 7953 355 8011 367
rect 8411 1633 8469 1645
rect 8411 367 8423 1633
rect 8457 367 8469 1633
rect 8411 355 8469 367
rect 8869 1633 8927 1645
rect 8869 367 8881 1633
rect 8915 367 8927 1633
rect 8869 355 8927 367
rect 9327 1633 9385 1645
rect 9327 367 9339 1633
rect 9373 367 9385 1633
rect 9327 355 9385 367
rect 9785 1633 9843 1645
rect 9785 367 9797 1633
rect 9831 367 9843 1633
rect 9785 355 9843 367
rect 10243 1633 10301 1645
rect 10243 367 10255 1633
rect 10289 367 10301 1633
rect 10243 355 10301 367
rect 10701 1633 10759 1645
rect 10701 367 10713 1633
rect 10747 367 10759 1633
rect 10701 355 10759 367
rect 11159 1633 11217 1645
rect 11159 367 11171 1633
rect 11205 367 11217 1633
rect 11159 355 11217 367
rect 11617 1633 11675 1645
rect 11617 367 11629 1633
rect 11663 367 11675 1633
rect 11617 355 11675 367
rect 12075 1633 12133 1645
rect 12075 367 12087 1633
rect 12121 367 12133 1633
rect 12075 355 12133 367
rect 12533 1633 12591 1645
rect 12533 367 12545 1633
rect 12579 367 12591 1633
rect 12533 355 12591 367
rect 12991 1633 13049 1645
rect 12991 367 13003 1633
rect 13037 367 13049 1633
rect 12991 355 13049 367
rect 13449 1633 13507 1645
rect 13449 367 13461 1633
rect 13495 367 13507 1633
rect 13449 355 13507 367
rect 13907 1633 13965 1645
rect 13907 367 13919 1633
rect 13953 367 13965 1633
rect 13907 355 13965 367
rect 14365 1633 14423 1645
rect 14365 367 14377 1633
rect 14411 367 14423 1633
rect 14365 355 14423 367
rect 14823 1633 14881 1645
rect 14823 367 14835 1633
rect 14869 367 14881 1633
rect 14823 355 14881 367
rect 15281 1633 15339 1645
rect 15281 367 15293 1633
rect 15327 367 15339 1633
rect 15281 355 15339 367
rect 15739 1633 15797 1645
rect 15739 367 15751 1633
rect 15785 367 15797 1633
rect 15739 355 15797 367
rect 16197 1633 16255 1645
rect 16197 367 16209 1633
rect 16243 367 16255 1633
rect 16197 355 16255 367
rect 16655 1633 16713 1645
rect 16655 367 16667 1633
rect 16701 367 16713 1633
rect 16655 355 16713 367
rect 17113 1633 17171 1645
rect 17113 367 17125 1633
rect 17159 367 17171 1633
rect 17113 355 17171 367
rect 17571 1633 17629 1645
rect 17571 367 17583 1633
rect 17617 367 17629 1633
rect 17571 355 17629 367
rect 18029 1633 18087 1645
rect 18029 367 18041 1633
rect 18075 367 18087 1633
rect 18029 355 18087 367
rect 18487 1633 18545 1645
rect 18487 367 18499 1633
rect 18533 367 18545 1633
rect 18487 355 18545 367
rect 18945 1633 19003 1645
rect 18945 367 18957 1633
rect 18991 367 19003 1633
rect 18945 355 19003 367
rect 19403 1633 19461 1645
rect 19403 367 19415 1633
rect 19449 367 19461 1633
rect 19403 355 19461 367
rect 19861 1633 19919 1645
rect 19861 367 19873 1633
rect 19907 367 19919 1633
rect 19861 355 19919 367
rect 20319 1633 20377 1645
rect 20319 367 20331 1633
rect 20365 367 20377 1633
rect 20319 355 20377 367
rect 20777 1633 20835 1645
rect 20777 367 20789 1633
rect 20823 367 20835 1633
rect 20777 355 20835 367
rect 21235 1633 21293 1645
rect 21235 367 21247 1633
rect 21281 367 21293 1633
rect 21235 355 21293 367
rect 21693 1633 21751 1645
rect 21693 367 21705 1633
rect 21739 367 21751 1633
rect 21693 355 21751 367
rect 22151 1633 22209 1645
rect 22151 367 22163 1633
rect 22197 367 22209 1633
rect 22151 355 22209 367
rect 22609 1633 22667 1645
rect 22609 367 22621 1633
rect 22655 367 22667 1633
rect 22609 355 22667 367
rect 23067 1633 23125 1645
rect 23067 367 23079 1633
rect 23113 367 23125 1633
rect 23067 355 23125 367
rect 23525 1633 23583 1645
rect 23525 367 23537 1633
rect 23571 367 23583 1633
rect 23525 355 23583 367
rect 23983 1633 24041 1645
rect 23983 367 23995 1633
rect 24029 367 24041 1633
rect 23983 355 24041 367
rect 24441 1633 24499 1645
rect 24441 367 24453 1633
rect 24487 367 24499 1633
rect 24441 355 24499 367
rect 24899 1633 24957 1645
rect 24899 367 24911 1633
rect 24945 367 24957 1633
rect 24899 355 24957 367
rect 25357 1633 25415 1645
rect 25357 367 25369 1633
rect 25403 367 25415 1633
rect 25357 355 25415 367
rect 25815 1633 25873 1645
rect 25815 367 25827 1633
rect 25861 367 25873 1633
rect 25815 355 25873 367
rect 26273 1633 26331 1645
rect 26273 367 26285 1633
rect 26319 367 26331 1633
rect 26273 355 26331 367
rect 26731 1633 26789 1645
rect 26731 367 26743 1633
rect 26777 367 26789 1633
rect 26731 355 26789 367
rect 27189 1633 27247 1645
rect 27189 367 27201 1633
rect 27235 367 27247 1633
rect 27189 355 27247 367
rect 27647 1633 27705 1645
rect 27647 367 27659 1633
rect 27693 367 27705 1633
rect 27647 355 27705 367
<< pdiffc >>
rect 179 367 213 1633
rect 637 367 671 1633
rect 1095 367 1129 1633
rect 1553 367 1587 1633
rect 2011 367 2045 1633
rect 2469 367 2503 1633
rect 2927 367 2961 1633
rect 3385 367 3419 1633
rect 3843 367 3877 1633
rect 4301 367 4335 1633
rect 4759 367 4793 1633
rect 5217 367 5251 1633
rect 5675 367 5709 1633
rect 6133 367 6167 1633
rect 6591 367 6625 1633
rect 7049 367 7083 1633
rect 7507 367 7541 1633
rect 7965 367 7999 1633
rect 8423 367 8457 1633
rect 8881 367 8915 1633
rect 9339 367 9373 1633
rect 9797 367 9831 1633
rect 10255 367 10289 1633
rect 10713 367 10747 1633
rect 11171 367 11205 1633
rect 11629 367 11663 1633
rect 12087 367 12121 1633
rect 12545 367 12579 1633
rect 13003 367 13037 1633
rect 13461 367 13495 1633
rect 13919 367 13953 1633
rect 14377 367 14411 1633
rect 14835 367 14869 1633
rect 15293 367 15327 1633
rect 15751 367 15785 1633
rect 16209 367 16243 1633
rect 16667 367 16701 1633
rect 17125 367 17159 1633
rect 17583 367 17617 1633
rect 18041 367 18075 1633
rect 18499 367 18533 1633
rect 18957 367 18991 1633
rect 19415 367 19449 1633
rect 19873 367 19907 1633
rect 20331 367 20365 1633
rect 20789 367 20823 1633
rect 21247 367 21281 1633
rect 21705 367 21739 1633
rect 22163 367 22197 1633
rect 22621 367 22655 1633
rect 23079 367 23113 1633
rect 23537 367 23571 1633
rect 23995 367 24029 1633
rect 24453 367 24487 1633
rect 24911 367 24945 1633
rect 25369 367 25403 1633
rect 25827 367 25861 1633
rect 26285 367 26319 1633
rect 26743 367 26777 1633
rect 27201 367 27235 1633
rect 27659 367 27693 1633
<< poly >>
rect 225 1645 625 1671
rect 683 1645 1083 1671
rect 1141 1645 1541 1671
rect 1599 1645 1999 1671
rect 2057 1645 2457 1671
rect 2515 1645 2915 1671
rect 2973 1645 3373 1671
rect 3431 1645 3831 1671
rect 3889 1645 4289 1671
rect 4347 1645 4747 1671
rect 4805 1645 5205 1671
rect 5263 1645 5663 1671
rect 5721 1645 6121 1671
rect 6179 1645 6579 1671
rect 6637 1645 7037 1671
rect 7095 1645 7495 1671
rect 7553 1645 7953 1671
rect 8011 1645 8411 1671
rect 8469 1645 8869 1671
rect 8927 1645 9327 1671
rect 9385 1645 9785 1671
rect 9843 1645 10243 1671
rect 10301 1645 10701 1671
rect 10759 1645 11159 1671
rect 11217 1645 11617 1671
rect 11675 1645 12075 1671
rect 12133 1645 12533 1671
rect 12591 1645 12991 1671
rect 13049 1645 13449 1671
rect 13507 1645 13907 1671
rect 13965 1645 14365 1671
rect 14423 1645 14823 1671
rect 14881 1645 15281 1671
rect 15339 1645 15739 1671
rect 15797 1645 16197 1671
rect 16255 1645 16655 1671
rect 16713 1645 17113 1671
rect 17171 1645 17571 1671
rect 17629 1645 18029 1671
rect 18087 1645 18487 1671
rect 18545 1645 18945 1671
rect 19003 1645 19403 1671
rect 19461 1645 19861 1671
rect 19919 1645 20319 1671
rect 20377 1645 20777 1671
rect 20835 1645 21235 1671
rect 21293 1645 21693 1671
rect 21751 1645 22151 1671
rect 22209 1645 22609 1671
rect 22667 1645 23067 1671
rect 23125 1645 23525 1671
rect 23583 1645 23983 1671
rect 24041 1645 24441 1671
rect 24499 1645 24899 1671
rect 24957 1645 25357 1671
rect 25415 1645 25815 1671
rect 25873 1645 26273 1671
rect 26331 1645 26731 1671
rect 26789 1645 27189 1671
rect 27247 1645 27647 1671
rect 225 329 625 355
rect 683 329 1083 355
rect 1141 329 1541 355
rect 1599 329 1999 355
rect 2057 329 2457 355
rect 2515 329 2915 355
rect 2973 329 3373 355
rect 3431 329 3831 355
rect 3889 329 4289 355
rect 4347 329 4747 355
rect 4805 329 5205 355
rect 5263 329 5663 355
rect 5721 329 6121 355
rect 6179 329 6579 355
rect 6637 329 7037 355
rect 7095 329 7495 355
rect 7553 329 7953 355
rect 8011 329 8411 355
rect 8469 329 8869 355
rect 8927 329 9327 355
rect 9385 329 9785 355
rect 9843 329 10243 355
rect 10301 329 10701 355
rect 10759 329 11159 355
rect 11217 329 11617 355
rect 11675 329 12075 355
rect 12133 329 12533 355
rect 12591 329 12991 355
rect 13049 329 13449 355
rect 13507 329 13907 355
rect 13965 329 14365 355
rect 14423 329 14823 355
rect 14881 329 15281 355
rect 15339 329 15739 355
rect 15797 329 16197 355
rect 16255 329 16655 355
rect 16713 329 17113 355
rect 17171 329 17571 355
rect 17629 329 18029 355
rect 18087 329 18487 355
rect 18545 329 18945 355
rect 19003 329 19403 355
rect 19461 329 19861 355
rect 19919 329 20319 355
rect 20377 329 20777 355
rect 20835 329 21235 355
rect 21293 329 21693 355
rect 21751 329 22151 355
rect 22209 329 22609 355
rect 22667 329 23067 355
rect 23125 329 23525 355
rect 23583 329 23983 355
rect 24041 329 24441 355
rect 24499 329 24899 355
rect 24957 329 25357 355
rect 25415 329 25815 355
rect 25873 329 26273 355
rect 26331 329 26731 355
rect 26789 329 27189 355
rect 27247 329 27647 355
rect 370 182 490 329
rect 826 182 946 329
rect 1282 182 1402 329
rect 1738 182 1858 329
rect 2194 182 2314 329
rect 2650 182 2770 329
rect 3106 182 3226 329
rect 3562 182 3682 329
rect 4018 182 4138 329
rect 4474 182 4594 329
rect 4930 182 5050 329
rect 5386 182 5506 329
rect 5842 182 5962 329
rect 6298 182 6418 329
rect 6754 182 6874 329
rect 7210 182 7330 329
rect 7666 182 7786 329
rect 8122 182 8242 329
rect 8578 182 8698 329
rect 9034 182 9154 329
rect 9490 182 9610 329
rect 9946 182 10066 329
rect 10402 182 10522 329
rect 10858 182 10978 329
rect 11314 182 11434 329
rect 11770 182 11890 329
rect 12226 182 12346 329
rect 12682 182 12802 329
rect 13138 182 13258 329
rect 13594 182 13714 329
rect 14050 182 14170 329
rect 14506 182 14626 329
rect 14962 182 15082 329
rect 15418 182 15538 329
rect 15874 182 15994 329
rect 16330 182 16450 329
rect 16786 182 16906 329
rect 17242 182 17362 329
rect 17698 182 17818 329
rect 18154 182 18274 329
rect 18610 182 18730 329
rect 19066 182 19186 329
rect 19522 182 19642 329
rect 19978 182 20098 329
rect 20434 182 20554 329
rect 20890 182 21010 329
rect 21346 182 21466 329
rect 21802 182 21922 329
rect 22258 182 22378 329
rect 22714 182 22834 329
rect 23170 182 23290 329
rect 23626 182 23746 329
rect 24082 182 24202 329
rect 24538 182 24658 329
rect 24994 182 25114 329
rect 25450 182 25570 329
rect 25906 182 26026 329
rect 26362 182 26482 329
rect 26818 182 26938 329
rect 27274 182 27394 329
rect 130 162 27740 182
rect 130 102 300 162
rect 360 102 700 162
rect 760 102 1100 162
rect 1160 102 1500 162
rect 1560 102 1900 162
rect 1960 102 2300 162
rect 2360 102 2700 162
rect 2760 102 3100 162
rect 3160 102 3500 162
rect 3560 102 3900 162
rect 3960 102 4300 162
rect 4360 102 4700 162
rect 4760 102 5100 162
rect 5160 102 5500 162
rect 5560 102 5900 162
rect 5960 102 6300 162
rect 6360 102 6700 162
rect 6760 102 7100 162
rect 7160 102 7500 162
rect 7560 102 7900 162
rect 7960 102 8300 162
rect 8360 102 8700 162
rect 8760 102 9100 162
rect 9160 102 9500 162
rect 9560 102 9900 162
rect 9960 102 10300 162
rect 10360 102 10700 162
rect 10760 102 11100 162
rect 11160 102 11500 162
rect 11560 102 11900 162
rect 11960 102 12300 162
rect 12360 102 12700 162
rect 12760 102 13100 162
rect 13160 102 13500 162
rect 13560 102 13900 162
rect 13960 102 14300 162
rect 14360 102 14700 162
rect 14760 102 15100 162
rect 15160 102 15500 162
rect 15560 102 15900 162
rect 15960 102 16300 162
rect 16360 102 16700 162
rect 16760 102 17100 162
rect 17160 102 17500 162
rect 17560 102 17900 162
rect 17960 102 18300 162
rect 18360 102 18700 162
rect 18760 102 19100 162
rect 19160 102 19500 162
rect 19560 102 19900 162
rect 19960 102 20300 162
rect 20360 102 20700 162
rect 20760 102 21100 162
rect 21160 102 21500 162
rect 21560 102 21900 162
rect 21960 102 22300 162
rect 22360 102 22700 162
rect 22760 102 23100 162
rect 23160 102 23500 162
rect 23560 102 23900 162
rect 23960 102 24300 162
rect 24360 102 24700 162
rect 24760 102 25100 162
rect 25160 102 25500 162
rect 25560 102 25900 162
rect 25960 102 26300 162
rect 26360 102 26700 162
rect 26760 102 27100 162
rect 27160 102 27500 162
rect 27560 102 27740 162
rect 130 82 27740 102
<< polycont >>
rect 300 102 360 162
rect 700 102 760 162
rect 1100 102 1160 162
rect 1500 102 1560 162
rect 1900 102 1960 162
rect 2300 102 2360 162
rect 2700 102 2760 162
rect 3100 102 3160 162
rect 3500 102 3560 162
rect 3900 102 3960 162
rect 4300 102 4360 162
rect 4700 102 4760 162
rect 5100 102 5160 162
rect 5500 102 5560 162
rect 5900 102 5960 162
rect 6300 102 6360 162
rect 6700 102 6760 162
rect 7100 102 7160 162
rect 7500 102 7560 162
rect 7900 102 7960 162
rect 8300 102 8360 162
rect 8700 102 8760 162
rect 9100 102 9160 162
rect 9500 102 9560 162
rect 9900 102 9960 162
rect 10300 102 10360 162
rect 10700 102 10760 162
rect 11100 102 11160 162
rect 11500 102 11560 162
rect 11900 102 11960 162
rect 12300 102 12360 162
rect 12700 102 12760 162
rect 13100 102 13160 162
rect 13500 102 13560 162
rect 13900 102 13960 162
rect 14300 102 14360 162
rect 14700 102 14760 162
rect 15100 102 15160 162
rect 15500 102 15560 162
rect 15900 102 15960 162
rect 16300 102 16360 162
rect 16700 102 16760 162
rect 17100 102 17160 162
rect 17500 102 17560 162
rect 17900 102 17960 162
rect 18300 102 18360 162
rect 18700 102 18760 162
rect 19100 102 19160 162
rect 19500 102 19560 162
rect 19900 102 19960 162
rect 20300 102 20360 162
rect 20700 102 20760 162
rect 21100 102 21160 162
rect 21500 102 21560 162
rect 21900 102 21960 162
rect 22300 102 22360 162
rect 22700 102 22760 162
rect 23100 102 23160 162
rect 23500 102 23560 162
rect 23900 102 23960 162
rect 24300 102 24360 162
rect 24700 102 24760 162
rect 25100 102 25160 162
rect 25500 102 25560 162
rect 25900 102 25960 162
rect 26300 102 26360 162
rect 26700 102 26760 162
rect 27100 102 27160 162
rect 27500 102 27560 162
<< locali >>
rect 130 1850 300 1910
rect 360 1850 700 1910
rect 760 1850 1100 1910
rect 1160 1850 1500 1910
rect 1560 1850 1900 1910
rect 1960 1850 2300 1910
rect 2360 1850 2700 1910
rect 2760 1850 3100 1910
rect 3160 1850 3500 1910
rect 3560 1850 3900 1910
rect 3960 1850 4300 1910
rect 4360 1850 4700 1910
rect 4760 1850 5100 1910
rect 5160 1850 5500 1910
rect 5560 1850 5900 1910
rect 5960 1850 6300 1910
rect 6360 1850 6700 1910
rect 6760 1850 7100 1910
rect 7160 1850 7500 1910
rect 7560 1850 7900 1910
rect 7960 1850 8300 1910
rect 8360 1850 8700 1910
rect 8760 1850 9100 1910
rect 9160 1850 9500 1910
rect 9560 1850 9900 1910
rect 9960 1850 10300 1910
rect 10360 1850 10700 1910
rect 10760 1850 11100 1910
rect 11160 1850 11500 1910
rect 11560 1850 11900 1910
rect 11960 1850 12300 1910
rect 12360 1850 12700 1910
rect 12760 1850 13100 1910
rect 13160 1850 13500 1910
rect 13560 1850 13900 1910
rect 13960 1850 14300 1910
rect 14360 1850 14700 1910
rect 14760 1850 15100 1910
rect 15160 1850 15500 1910
rect 15560 1850 15900 1910
rect 15960 1850 16300 1910
rect 16360 1850 16700 1910
rect 16760 1850 17100 1910
rect 17160 1850 17500 1910
rect 17560 1850 17900 1910
rect 17960 1850 18300 1910
rect 18360 1850 18700 1910
rect 18760 1850 19100 1910
rect 19160 1850 19500 1910
rect 19560 1850 19900 1910
rect 19960 1850 20300 1910
rect 20360 1850 20700 1910
rect 20760 1850 21100 1910
rect 21160 1850 21500 1910
rect 21560 1850 21900 1910
rect 21960 1850 22300 1910
rect 22360 1850 22700 1910
rect 22760 1850 23100 1910
rect 23160 1850 23500 1910
rect 23560 1850 23900 1910
rect 23960 1850 24300 1910
rect 24360 1850 24700 1910
rect 24760 1850 25100 1910
rect 25160 1850 25500 1910
rect 25560 1850 25900 1910
rect 25960 1850 26300 1910
rect 26360 1850 26700 1910
rect 26760 1850 27100 1910
rect 27160 1850 27500 1910
rect 27560 1850 27740 1910
rect 130 1730 27740 1790
rect 635 1649 669 1730
rect 1551 1649 1585 1730
rect 2467 1649 2501 1730
rect 3383 1649 3417 1730
rect 4299 1649 4333 1730
rect 5215 1649 5249 1730
rect 6131 1649 6165 1730
rect 7047 1649 7081 1730
rect 7963 1649 7997 1730
rect 8879 1649 8913 1730
rect 9795 1649 9829 1730
rect 10711 1649 10745 1730
rect 11627 1649 11661 1730
rect 12543 1649 12577 1730
rect 13459 1649 13493 1730
rect 14375 1649 14409 1730
rect 15291 1649 15325 1730
rect 16207 1649 16241 1730
rect 17123 1649 17157 1730
rect 18039 1649 18073 1730
rect 18955 1649 18989 1730
rect 19871 1649 19905 1730
rect 20787 1649 20821 1730
rect 21703 1649 21737 1730
rect 22619 1649 22653 1730
rect 23535 1649 23569 1730
rect 24451 1649 24485 1730
rect 25367 1649 25401 1730
rect 26283 1649 26317 1730
rect 27199 1649 27233 1730
rect 179 1633 213 1649
rect 177 367 179 372
rect 635 1633 671 1649
rect 635 1626 637 1633
rect 177 351 213 367
rect 1095 1633 1129 1649
rect 637 351 671 367
rect 1093 367 1095 372
rect 1551 1633 1587 1649
rect 1551 1626 1553 1633
rect 1093 351 1129 367
rect 2011 1633 2045 1649
rect 1553 351 1587 367
rect 2009 367 2011 372
rect 2467 1633 2503 1649
rect 2467 1626 2469 1633
rect 2009 351 2045 367
rect 2927 1633 2961 1649
rect 2469 351 2503 367
rect 2925 367 2927 372
rect 3383 1633 3419 1649
rect 3383 1626 3385 1633
rect 2925 351 2961 367
rect 3843 1633 3877 1649
rect 3385 351 3419 367
rect 3841 367 3843 372
rect 4299 1633 4335 1649
rect 4299 1626 4301 1633
rect 3841 351 3877 367
rect 4759 1633 4793 1649
rect 4301 351 4335 367
rect 4757 367 4759 372
rect 5215 1633 5251 1649
rect 5215 1626 5217 1633
rect 4757 351 4793 367
rect 5675 1633 5709 1649
rect 5217 351 5251 367
rect 5673 367 5675 372
rect 6131 1633 6167 1649
rect 6131 1626 6133 1633
rect 5673 351 5709 367
rect 6591 1633 6625 1649
rect 6133 351 6167 367
rect 6589 367 6591 372
rect 7047 1633 7083 1649
rect 7047 1626 7049 1633
rect 6589 351 6625 367
rect 7507 1633 7541 1649
rect 7049 351 7083 367
rect 7505 367 7507 372
rect 7963 1633 7999 1649
rect 7963 1626 7965 1633
rect 7505 351 7541 367
rect 8423 1633 8457 1649
rect 7965 351 7999 367
rect 8421 367 8423 372
rect 8879 1633 8915 1649
rect 8879 1626 8881 1633
rect 8421 351 8457 367
rect 9339 1633 9373 1649
rect 8881 351 8915 367
rect 9337 367 9339 372
rect 9795 1633 9831 1649
rect 9795 1626 9797 1633
rect 9337 351 9373 367
rect 10255 1633 10289 1649
rect 9797 351 9831 367
rect 10253 367 10255 372
rect 10711 1633 10747 1649
rect 10711 1626 10713 1633
rect 10253 351 10289 367
rect 11171 1633 11205 1649
rect 10713 351 10747 367
rect 11169 367 11171 372
rect 11627 1633 11663 1649
rect 11627 1626 11629 1633
rect 11169 351 11205 367
rect 12087 1633 12121 1649
rect 11629 351 11663 367
rect 12085 367 12087 372
rect 12543 1633 12579 1649
rect 12543 1626 12545 1633
rect 12085 351 12121 367
rect 13003 1633 13037 1649
rect 12545 351 12579 367
rect 13001 367 13003 372
rect 13459 1633 13495 1649
rect 13459 1626 13461 1633
rect 13001 351 13037 367
rect 13919 1633 13953 1649
rect 13461 351 13495 367
rect 13917 367 13919 372
rect 14375 1633 14411 1649
rect 14375 1626 14377 1633
rect 13917 351 13953 367
rect 14835 1633 14869 1649
rect 14377 351 14411 367
rect 14833 367 14835 372
rect 15291 1633 15327 1649
rect 15291 1626 15293 1633
rect 14833 351 14869 367
rect 15751 1633 15785 1649
rect 15293 351 15327 367
rect 15749 367 15751 372
rect 16207 1633 16243 1649
rect 16207 1626 16209 1633
rect 15749 351 15785 367
rect 16667 1633 16701 1649
rect 16209 351 16243 367
rect 16665 367 16667 372
rect 17123 1633 17159 1649
rect 17123 1626 17125 1633
rect 16665 351 16701 367
rect 17583 1633 17617 1649
rect 17125 351 17159 367
rect 17581 367 17583 372
rect 18039 1633 18075 1649
rect 18039 1626 18041 1633
rect 17581 351 17617 367
rect 18499 1633 18533 1649
rect 18041 351 18075 367
rect 18497 367 18499 372
rect 18955 1633 18991 1649
rect 18955 1626 18957 1633
rect 18497 351 18533 367
rect 19415 1633 19449 1649
rect 18957 351 18991 367
rect 19413 367 19415 372
rect 19871 1633 19907 1649
rect 19871 1626 19873 1633
rect 19413 351 19449 367
rect 20331 1633 20365 1649
rect 19873 351 19907 367
rect 20329 367 20331 372
rect 20787 1633 20823 1649
rect 20787 1626 20789 1633
rect 20329 351 20365 367
rect 21247 1633 21281 1649
rect 20789 351 20823 367
rect 21245 367 21247 372
rect 21703 1633 21739 1649
rect 21703 1626 21705 1633
rect 21245 351 21281 367
rect 22163 1633 22197 1649
rect 21705 351 21739 367
rect 22161 367 22163 372
rect 22619 1633 22655 1649
rect 22619 1626 22621 1633
rect 22161 351 22197 367
rect 23079 1633 23113 1649
rect 22621 351 22655 367
rect 23077 367 23079 372
rect 23535 1633 23571 1649
rect 23535 1626 23537 1633
rect 23077 351 23113 367
rect 23995 1633 24029 1649
rect 23537 351 23571 367
rect 23993 367 23995 372
rect 24451 1633 24487 1649
rect 24451 1626 24453 1633
rect 23993 351 24029 367
rect 24911 1633 24945 1649
rect 24453 351 24487 367
rect 24909 367 24911 372
rect 25367 1633 25403 1649
rect 25367 1626 25369 1633
rect 24909 351 24945 367
rect 25827 1633 25861 1649
rect 25369 351 25403 367
rect 25825 367 25827 372
rect 26283 1633 26319 1649
rect 26283 1626 26285 1633
rect 25825 351 25861 367
rect 26743 1633 26777 1649
rect 26285 351 26319 367
rect 26741 367 26743 372
rect 27199 1633 27235 1649
rect 27199 1626 27201 1633
rect 26741 351 26777 367
rect 27659 1633 27693 1649
rect 27201 351 27235 367
rect 27657 367 27659 372
rect 27657 351 27693 367
rect 177 270 211 351
rect 1093 270 1127 351
rect 2009 270 2043 351
rect 2925 270 2959 351
rect 3841 270 3875 351
rect 4757 270 4791 351
rect 5673 270 5707 351
rect 6589 270 6623 351
rect 7505 270 7539 351
rect 8421 270 8455 351
rect 9337 270 9371 351
rect 10253 270 10287 351
rect 11169 270 11203 351
rect 12085 270 12119 351
rect 13001 270 13035 351
rect 13917 270 13951 351
rect 14833 270 14867 351
rect 15749 270 15783 351
rect 16665 270 16699 351
rect 17581 270 17615 351
rect 18497 270 18531 351
rect 19413 270 19447 351
rect 20329 270 20363 351
rect 21245 270 21279 351
rect 22161 270 22195 351
rect 23077 270 23111 351
rect 23993 270 24027 351
rect 24909 270 24943 351
rect 25825 270 25859 351
rect 26741 270 26775 351
rect 27657 270 27691 351
rect 130 210 27740 270
rect 130 102 300 162
rect 360 102 700 162
rect 760 102 1100 162
rect 1160 102 1500 162
rect 1560 102 1900 162
rect 1960 102 2300 162
rect 2360 102 2700 162
rect 2760 102 3100 162
rect 3160 102 3500 162
rect 3560 102 3900 162
rect 3960 102 4300 162
rect 4360 102 4700 162
rect 4760 102 5100 162
rect 5160 102 5500 162
rect 5560 102 5900 162
rect 5960 102 6300 162
rect 6360 102 6700 162
rect 6760 102 7100 162
rect 7160 102 7500 162
rect 7560 102 7900 162
rect 7960 102 8300 162
rect 8360 102 8700 162
rect 8760 102 9100 162
rect 9160 102 9500 162
rect 9560 102 9900 162
rect 9960 102 10300 162
rect 10360 102 10700 162
rect 10760 102 11100 162
rect 11160 102 11500 162
rect 11560 102 11900 162
rect 11960 102 12300 162
rect 12360 102 12700 162
rect 12760 102 13100 162
rect 13160 102 13500 162
rect 13560 102 13900 162
rect 13960 102 14300 162
rect 14360 102 14700 162
rect 14760 102 15100 162
rect 15160 102 15500 162
rect 15560 102 15900 162
rect 15960 102 16300 162
rect 16360 102 16700 162
rect 16760 102 17100 162
rect 17160 102 17500 162
rect 17560 102 17900 162
rect 17960 102 18300 162
rect 18360 102 18700 162
rect 18760 102 19100 162
rect 19160 102 19500 162
rect 19560 102 19900 162
rect 19960 102 20300 162
rect 20360 102 20700 162
rect 20760 102 21100 162
rect 21160 102 21500 162
rect 21560 102 21900 162
rect 21960 102 22300 162
rect 22360 102 22700 162
rect 22760 102 23100 162
rect 23160 102 23500 162
rect 23560 102 23900 162
rect 23960 102 24300 162
rect 24360 102 24700 162
rect 24760 102 25100 162
rect 25160 102 25500 162
rect 25560 102 25900 162
rect 25960 102 26300 162
rect 26360 102 26700 162
rect 26760 102 27100 162
rect 27160 102 27500 162
rect 27560 102 27740 162
rect 130 -30 300 30
rect 360 -30 700 30
rect 760 -30 1100 30
rect 1160 -30 1500 30
rect 1560 -30 1900 30
rect 1960 -30 2300 30
rect 2360 -30 2700 30
rect 2760 -30 3100 30
rect 3160 -30 3500 30
rect 3560 -30 3900 30
rect 3960 -30 4300 30
rect 4360 -30 4700 30
rect 4760 -30 5100 30
rect 5160 -30 5500 30
rect 5560 -30 5900 30
rect 5960 -30 6300 30
rect 6360 -30 6700 30
rect 6760 -30 7100 30
rect 7160 -30 7500 30
rect 7560 -30 7900 30
rect 7960 -30 8300 30
rect 8360 -30 8700 30
rect 8760 -30 9100 30
rect 9160 -30 9500 30
rect 9560 -30 9900 30
rect 9960 -30 10300 30
rect 10360 -30 10700 30
rect 10760 -30 11100 30
rect 11160 -30 11500 30
rect 11560 -30 11900 30
rect 11960 -30 12300 30
rect 12360 -30 12700 30
rect 12760 -30 13100 30
rect 13160 -30 13500 30
rect 13560 -30 13900 30
rect 13960 -30 14300 30
rect 14360 -30 14700 30
rect 14760 -30 15100 30
rect 15160 -30 15500 30
rect 15560 -30 15900 30
rect 15960 -30 16300 30
rect 16360 -30 16700 30
rect 16760 -30 17100 30
rect 17160 -30 17500 30
rect 17560 -30 17900 30
rect 17960 -30 18300 30
rect 18360 -30 18700 30
rect 18760 -30 19100 30
rect 19160 -30 19500 30
rect 19560 -30 19900 30
rect 19960 -30 20300 30
rect 20360 -30 20700 30
rect 20760 -30 21100 30
rect 21160 -30 21500 30
rect 21560 -30 21900 30
rect 21960 -30 22300 30
rect 22360 -30 22700 30
rect 22760 -30 23100 30
rect 23160 -30 23500 30
rect 23560 -30 23900 30
rect 23960 -30 24300 30
rect 24360 -30 24700 30
rect 24760 -30 25100 30
rect 25160 -30 25500 30
rect 25560 -30 25900 30
rect 25960 -30 26300 30
rect 26360 -30 26700 30
rect 26760 -30 27100 30
rect 27160 -30 27500 30
rect 27560 -30 27740 30
<< viali >>
rect 300 1850 360 1910
rect 700 1850 760 1910
rect 1100 1850 1160 1910
rect 1500 1850 1560 1910
rect 1900 1850 1960 1910
rect 2300 1850 2360 1910
rect 2700 1850 2760 1910
rect 3100 1850 3160 1910
rect 3500 1850 3560 1910
rect 3900 1850 3960 1910
rect 4300 1850 4360 1910
rect 4700 1850 4760 1910
rect 5100 1850 5160 1910
rect 5500 1850 5560 1910
rect 5900 1850 5960 1910
rect 6300 1850 6360 1910
rect 6700 1850 6760 1910
rect 7100 1850 7160 1910
rect 7500 1850 7560 1910
rect 7900 1850 7960 1910
rect 8300 1850 8360 1910
rect 8700 1850 8760 1910
rect 9100 1850 9160 1910
rect 9500 1850 9560 1910
rect 9900 1850 9960 1910
rect 10300 1850 10360 1910
rect 10700 1850 10760 1910
rect 11100 1850 11160 1910
rect 11500 1850 11560 1910
rect 11900 1850 11960 1910
rect 12300 1850 12360 1910
rect 12700 1850 12760 1910
rect 13100 1850 13160 1910
rect 13500 1850 13560 1910
rect 13900 1850 13960 1910
rect 14300 1850 14360 1910
rect 14700 1850 14760 1910
rect 15100 1850 15160 1910
rect 15500 1850 15560 1910
rect 15900 1850 15960 1910
rect 16300 1850 16360 1910
rect 16700 1850 16760 1910
rect 17100 1850 17160 1910
rect 17500 1850 17560 1910
rect 17900 1850 17960 1910
rect 18300 1850 18360 1910
rect 18700 1850 18760 1910
rect 19100 1850 19160 1910
rect 19500 1850 19560 1910
rect 19900 1850 19960 1910
rect 20300 1850 20360 1910
rect 20700 1850 20760 1910
rect 21100 1850 21160 1910
rect 21500 1850 21560 1910
rect 21900 1850 21960 1910
rect 22300 1850 22360 1910
rect 22700 1850 22760 1910
rect 23100 1850 23160 1910
rect 23500 1850 23560 1910
rect 23900 1850 23960 1910
rect 24300 1850 24360 1910
rect 24700 1850 24760 1910
rect 25100 1850 25160 1910
rect 25500 1850 25560 1910
rect 25900 1850 25960 1910
rect 26300 1850 26360 1910
rect 26700 1850 26760 1910
rect 27100 1850 27160 1910
rect 27500 1850 27560 1910
rect 179 367 213 1633
rect 637 367 671 1633
rect 1095 367 1129 1633
rect 1553 367 1587 1633
rect 2011 367 2045 1633
rect 2469 367 2503 1633
rect 2927 367 2961 1633
rect 3385 367 3419 1633
rect 3843 367 3877 1633
rect 4301 367 4335 1633
rect 4759 367 4793 1633
rect 5217 367 5251 1633
rect 5675 367 5709 1633
rect 6133 367 6167 1633
rect 6591 367 6625 1633
rect 7049 367 7083 1633
rect 7507 367 7541 1633
rect 7965 367 7999 1633
rect 8423 367 8457 1633
rect 8881 367 8915 1633
rect 9339 367 9373 1633
rect 9797 367 9831 1633
rect 10255 367 10289 1633
rect 10713 367 10747 1633
rect 11171 367 11205 1633
rect 11629 367 11663 1633
rect 12087 367 12121 1633
rect 12545 367 12579 1633
rect 13003 367 13037 1633
rect 13461 367 13495 1633
rect 13919 367 13953 1633
rect 14377 367 14411 1633
rect 14835 367 14869 1633
rect 15293 367 15327 1633
rect 15751 367 15785 1633
rect 16209 367 16243 1633
rect 16667 367 16701 1633
rect 17125 367 17159 1633
rect 17583 367 17617 1633
rect 18041 367 18075 1633
rect 18499 367 18533 1633
rect 18957 367 18991 1633
rect 19415 367 19449 1633
rect 19873 367 19907 1633
rect 20331 367 20365 1633
rect 20789 367 20823 1633
rect 21247 367 21281 1633
rect 21705 367 21739 1633
rect 22163 367 22197 1633
rect 22621 367 22655 1633
rect 23079 367 23113 1633
rect 23537 367 23571 1633
rect 23995 367 24029 1633
rect 24453 367 24487 1633
rect 24911 367 24945 1633
rect 25369 367 25403 1633
rect 25827 367 25861 1633
rect 26285 367 26319 1633
rect 26743 367 26777 1633
rect 27201 367 27235 1633
rect 27659 367 27693 1633
rect 300 -30 360 30
rect 700 -30 760 30
rect 1100 -30 1160 30
rect 1500 -30 1560 30
rect 1900 -30 1960 30
rect 2300 -30 2360 30
rect 2700 -30 2760 30
rect 3100 -30 3160 30
rect 3500 -30 3560 30
rect 3900 -30 3960 30
rect 4300 -30 4360 30
rect 4700 -30 4760 30
rect 5100 -30 5160 30
rect 5500 -30 5560 30
rect 5900 -30 5960 30
rect 6300 -30 6360 30
rect 6700 -30 6760 30
rect 7100 -30 7160 30
rect 7500 -30 7560 30
rect 7900 -30 7960 30
rect 8300 -30 8360 30
rect 8700 -30 8760 30
rect 9100 -30 9160 30
rect 9500 -30 9560 30
rect 9900 -30 9960 30
rect 10300 -30 10360 30
rect 10700 -30 10760 30
rect 11100 -30 11160 30
rect 11500 -30 11560 30
rect 11900 -30 11960 30
rect 12300 -30 12360 30
rect 12700 -30 12760 30
rect 13100 -30 13160 30
rect 13500 -30 13560 30
rect 13900 -30 13960 30
rect 14300 -30 14360 30
rect 14700 -30 14760 30
rect 15100 -30 15160 30
rect 15500 -30 15560 30
rect 15900 -30 15960 30
rect 16300 -30 16360 30
rect 16700 -30 16760 30
rect 17100 -30 17160 30
rect 17500 -30 17560 30
rect 17900 -30 17960 30
rect 18300 -30 18360 30
rect 18700 -30 18760 30
rect 19100 -30 19160 30
rect 19500 -30 19560 30
rect 19900 -30 19960 30
rect 20300 -30 20360 30
rect 20700 -30 20760 30
rect 21100 -30 21160 30
rect 21500 -30 21560 30
rect 21900 -30 21960 30
rect 22300 -30 22360 30
rect 22700 -30 22760 30
rect 23100 -30 23160 30
rect 23500 -30 23560 30
rect 23900 -30 23960 30
rect 24300 -30 24360 30
rect 24700 -30 24760 30
rect 25100 -30 25160 30
rect 25500 -30 25560 30
rect 25900 -30 25960 30
rect 26300 -30 26360 30
rect 26700 -30 26760 30
rect 27100 -30 27160 30
rect 27500 -30 27560 30
<< metal1 >>
rect 130 1910 27740 1940
rect 130 1850 300 1910
rect 360 1850 700 1910
rect 760 1850 1100 1910
rect 1160 1850 1500 1910
rect 1560 1850 1900 1910
rect 1960 1850 2300 1910
rect 2360 1850 2700 1910
rect 2760 1850 3100 1910
rect 3160 1850 3500 1910
rect 3560 1850 3900 1910
rect 3960 1850 4300 1910
rect 4360 1850 4700 1910
rect 4760 1850 5100 1910
rect 5160 1850 5500 1910
rect 5560 1850 5900 1910
rect 5960 1850 6300 1910
rect 6360 1850 6700 1910
rect 6760 1850 7100 1910
rect 7160 1850 7500 1910
rect 7560 1850 7900 1910
rect 7960 1850 8300 1910
rect 8360 1850 8700 1910
rect 8760 1850 9100 1910
rect 9160 1850 9500 1910
rect 9560 1850 9900 1910
rect 9960 1850 10300 1910
rect 10360 1850 10700 1910
rect 10760 1850 11100 1910
rect 11160 1850 11500 1910
rect 11560 1850 11900 1910
rect 11960 1850 12300 1910
rect 12360 1850 12700 1910
rect 12760 1850 13100 1910
rect 13160 1850 13500 1910
rect 13560 1850 13900 1910
rect 13960 1850 14300 1910
rect 14360 1850 14700 1910
rect 14760 1850 15100 1910
rect 15160 1850 15500 1910
rect 15560 1850 15900 1910
rect 15960 1850 16300 1910
rect 16360 1850 16700 1910
rect 16760 1850 17100 1910
rect 17160 1850 17500 1910
rect 17560 1850 17900 1910
rect 17960 1850 18300 1910
rect 18360 1850 18700 1910
rect 18760 1850 19100 1910
rect 19160 1850 19500 1910
rect 19560 1850 19900 1910
rect 19960 1850 20300 1910
rect 20360 1850 20700 1910
rect 20760 1850 21100 1910
rect 21160 1850 21500 1910
rect 21560 1850 21900 1910
rect 21960 1850 22300 1910
rect 22360 1850 22700 1910
rect 22760 1850 23100 1910
rect 23160 1850 23500 1910
rect 23560 1850 23900 1910
rect 23960 1850 24300 1910
rect 24360 1850 24700 1910
rect 24760 1850 25100 1910
rect 25160 1850 25500 1910
rect 25560 1850 25900 1910
rect 25960 1850 26300 1910
rect 26360 1850 26700 1910
rect 26760 1850 27100 1910
rect 27160 1850 27500 1910
rect 27560 1850 27740 1910
rect 130 1820 27740 1850
rect 173 1633 219 1645
rect 173 367 179 1633
rect 213 367 219 1633
rect 173 355 219 367
rect 631 1633 677 1645
rect 631 367 637 1633
rect 671 367 677 1633
rect 631 355 677 367
rect 1089 1633 1135 1645
rect 1089 367 1095 1633
rect 1129 367 1135 1633
rect 1089 355 1135 367
rect 1547 1633 1593 1645
rect 1547 367 1553 1633
rect 1587 367 1593 1633
rect 1547 355 1593 367
rect 2005 1633 2051 1645
rect 2005 367 2011 1633
rect 2045 367 2051 1633
rect 2005 355 2051 367
rect 2463 1633 2509 1645
rect 2463 367 2469 1633
rect 2503 367 2509 1633
rect 2463 355 2509 367
rect 2921 1633 2967 1645
rect 2921 367 2927 1633
rect 2961 367 2967 1633
rect 2921 355 2967 367
rect 3379 1633 3425 1645
rect 3379 367 3385 1633
rect 3419 367 3425 1633
rect 3379 355 3425 367
rect 3837 1633 3883 1645
rect 3837 367 3843 1633
rect 3877 367 3883 1633
rect 3837 355 3883 367
rect 4295 1633 4341 1645
rect 4295 367 4301 1633
rect 4335 367 4341 1633
rect 4295 355 4341 367
rect 4753 1633 4799 1645
rect 4753 367 4759 1633
rect 4793 367 4799 1633
rect 4753 355 4799 367
rect 5211 1633 5257 1645
rect 5211 367 5217 1633
rect 5251 367 5257 1633
rect 5211 355 5257 367
rect 5669 1633 5715 1645
rect 5669 367 5675 1633
rect 5709 367 5715 1633
rect 5669 355 5715 367
rect 6127 1633 6173 1645
rect 6127 367 6133 1633
rect 6167 367 6173 1633
rect 6127 355 6173 367
rect 6585 1633 6631 1645
rect 6585 367 6591 1633
rect 6625 367 6631 1633
rect 6585 355 6631 367
rect 7043 1633 7089 1645
rect 7043 367 7049 1633
rect 7083 367 7089 1633
rect 7043 355 7089 367
rect 7501 1633 7547 1645
rect 7501 367 7507 1633
rect 7541 367 7547 1633
rect 7501 355 7547 367
rect 7959 1633 8005 1645
rect 7959 367 7965 1633
rect 7999 367 8005 1633
rect 7959 355 8005 367
rect 8417 1633 8463 1645
rect 8417 367 8423 1633
rect 8457 367 8463 1633
rect 8417 355 8463 367
rect 8875 1633 8921 1645
rect 8875 367 8881 1633
rect 8915 367 8921 1633
rect 8875 355 8921 367
rect 9333 1633 9379 1645
rect 9333 367 9339 1633
rect 9373 367 9379 1633
rect 9333 355 9379 367
rect 9791 1633 9837 1645
rect 9791 367 9797 1633
rect 9831 367 9837 1633
rect 9791 355 9837 367
rect 10249 1633 10295 1645
rect 10249 367 10255 1633
rect 10289 367 10295 1633
rect 10249 355 10295 367
rect 10707 1633 10753 1645
rect 10707 367 10713 1633
rect 10747 367 10753 1633
rect 10707 355 10753 367
rect 11165 1633 11211 1645
rect 11165 367 11171 1633
rect 11205 367 11211 1633
rect 11165 355 11211 367
rect 11623 1633 11669 1645
rect 11623 367 11629 1633
rect 11663 367 11669 1633
rect 11623 355 11669 367
rect 12081 1633 12127 1645
rect 12081 367 12087 1633
rect 12121 367 12127 1633
rect 12081 355 12127 367
rect 12539 1633 12585 1645
rect 12539 367 12545 1633
rect 12579 367 12585 1633
rect 12539 355 12585 367
rect 12997 1633 13043 1645
rect 12997 367 13003 1633
rect 13037 367 13043 1633
rect 12997 355 13043 367
rect 13455 1633 13501 1645
rect 13455 367 13461 1633
rect 13495 367 13501 1633
rect 13455 355 13501 367
rect 13913 1633 13959 1645
rect 13913 367 13919 1633
rect 13953 367 13959 1633
rect 13913 355 13959 367
rect 14371 1633 14417 1645
rect 14371 367 14377 1633
rect 14411 367 14417 1633
rect 14371 355 14417 367
rect 14829 1633 14875 1645
rect 14829 367 14835 1633
rect 14869 367 14875 1633
rect 14829 355 14875 367
rect 15287 1633 15333 1645
rect 15287 367 15293 1633
rect 15327 367 15333 1633
rect 15287 355 15333 367
rect 15745 1633 15791 1645
rect 15745 367 15751 1633
rect 15785 367 15791 1633
rect 15745 355 15791 367
rect 16203 1633 16249 1645
rect 16203 367 16209 1633
rect 16243 367 16249 1633
rect 16203 355 16249 367
rect 16661 1633 16707 1645
rect 16661 367 16667 1633
rect 16701 367 16707 1633
rect 16661 355 16707 367
rect 17119 1633 17165 1645
rect 17119 367 17125 1633
rect 17159 367 17165 1633
rect 17119 355 17165 367
rect 17577 1633 17623 1645
rect 17577 367 17583 1633
rect 17617 367 17623 1633
rect 17577 355 17623 367
rect 18035 1633 18081 1645
rect 18035 367 18041 1633
rect 18075 367 18081 1633
rect 18035 355 18081 367
rect 18493 1633 18539 1645
rect 18493 367 18499 1633
rect 18533 367 18539 1633
rect 18493 355 18539 367
rect 18951 1633 18997 1645
rect 18951 367 18957 1633
rect 18991 367 18997 1633
rect 18951 355 18997 367
rect 19409 1633 19455 1645
rect 19409 367 19415 1633
rect 19449 367 19455 1633
rect 19409 355 19455 367
rect 19867 1633 19913 1645
rect 19867 367 19873 1633
rect 19907 367 19913 1633
rect 19867 355 19913 367
rect 20325 1633 20371 1645
rect 20325 367 20331 1633
rect 20365 367 20371 1633
rect 20325 355 20371 367
rect 20783 1633 20829 1645
rect 20783 367 20789 1633
rect 20823 367 20829 1633
rect 20783 355 20829 367
rect 21241 1633 21287 1645
rect 21241 367 21247 1633
rect 21281 367 21287 1633
rect 21241 355 21287 367
rect 21699 1633 21745 1645
rect 21699 367 21705 1633
rect 21739 367 21745 1633
rect 21699 355 21745 367
rect 22157 1633 22203 1645
rect 22157 367 22163 1633
rect 22197 367 22203 1633
rect 22157 355 22203 367
rect 22615 1633 22661 1645
rect 22615 367 22621 1633
rect 22655 367 22661 1633
rect 22615 355 22661 367
rect 23073 1633 23119 1645
rect 23073 367 23079 1633
rect 23113 367 23119 1633
rect 23073 355 23119 367
rect 23531 1633 23577 1645
rect 23531 367 23537 1633
rect 23571 367 23577 1633
rect 23531 355 23577 367
rect 23989 1633 24035 1645
rect 23989 367 23995 1633
rect 24029 367 24035 1633
rect 23989 355 24035 367
rect 24447 1633 24493 1645
rect 24447 367 24453 1633
rect 24487 367 24493 1633
rect 24447 355 24493 367
rect 24905 1633 24951 1645
rect 24905 367 24911 1633
rect 24945 367 24951 1633
rect 24905 355 24951 367
rect 25363 1633 25409 1645
rect 25363 367 25369 1633
rect 25403 367 25409 1633
rect 25363 355 25409 367
rect 25821 1633 25867 1645
rect 25821 367 25827 1633
rect 25861 367 25867 1633
rect 25821 355 25867 367
rect 26279 1633 26325 1645
rect 26279 367 26285 1633
rect 26319 367 26325 1633
rect 26279 355 26325 367
rect 26737 1633 26783 1645
rect 26737 367 26743 1633
rect 26777 367 26783 1633
rect 26737 355 26783 367
rect 27195 1633 27241 1645
rect 27195 367 27201 1633
rect 27235 367 27241 1633
rect 27195 355 27241 367
rect 27653 1633 27699 1645
rect 27653 367 27659 1633
rect 27693 367 27699 1633
rect 27653 355 27699 367
rect 130 30 27740 60
rect 130 -30 300 30
rect 360 -30 700 30
rect 760 -30 1100 30
rect 1160 -30 1500 30
rect 1560 -30 1900 30
rect 1960 -30 2300 30
rect 2360 -30 2700 30
rect 2760 -30 3100 30
rect 3160 -30 3500 30
rect 3560 -30 3900 30
rect 3960 -30 4300 30
rect 4360 -30 4700 30
rect 4760 -30 5100 30
rect 5160 -30 5500 30
rect 5560 -30 5900 30
rect 5960 -30 6300 30
rect 6360 -30 6700 30
rect 6760 -30 7100 30
rect 7160 -30 7500 30
rect 7560 -30 7900 30
rect 7960 -30 8300 30
rect 8360 -30 8700 30
rect 8760 -30 9100 30
rect 9160 -30 9500 30
rect 9560 -30 9900 30
rect 9960 -30 10300 30
rect 10360 -30 10700 30
rect 10760 -30 11100 30
rect 11160 -30 11500 30
rect 11560 -30 11900 30
rect 11960 -30 12300 30
rect 12360 -30 12700 30
rect 12760 -30 13100 30
rect 13160 -30 13500 30
rect 13560 -30 13900 30
rect 13960 -30 14300 30
rect 14360 -30 14700 30
rect 14760 -30 15100 30
rect 15160 -30 15500 30
rect 15560 -30 15900 30
rect 15960 -30 16300 30
rect 16360 -30 16700 30
rect 16760 -30 17100 30
rect 17160 -30 17500 30
rect 17560 -30 17900 30
rect 17960 -30 18300 30
rect 18360 -30 18700 30
rect 18760 -30 19100 30
rect 19160 -30 19500 30
rect 19560 -30 19900 30
rect 19960 -30 20300 30
rect 20360 -30 20700 30
rect 20760 -30 21100 30
rect 21160 -30 21500 30
rect 21560 -30 21900 30
rect 21960 -30 22300 30
rect 22360 -30 22700 30
rect 22760 -30 23100 30
rect 23160 -30 23500 30
rect 23560 -30 23900 30
rect 23960 -30 24300 30
rect 24360 -30 24700 30
rect 24760 -30 25100 30
rect 25160 -30 25500 30
rect 25560 -30 25900 30
rect 25960 -30 26300 30
rect 26360 -30 26700 30
rect 26760 -30 27100 30
rect 27160 -30 27500 30
rect 27560 -30 27740 30
rect 130 -60 27740 -30
<< labels >>
flabel metal1 130 1850 190 1910 1 FreeSans 480 0 0 0 VPWR
port 4 n power bidirectional
flabel space 120 1850 180 1910 1 FreeSans 480 0 0 0 VPB
flabel metal1 130 -30 190 30 1 FreeSans 480 0 0 0 VGND
port 5 n ground bidirectional
flabel locali 27680 1730 27740 1790 1 FreeSans 480 0 0 0 SOURCE
port 2 n signal bidirectional
flabel locali 27680 210 27740 270 1 FreeSans 480 0 0 0 DRAIN
port 3 n signal bidirectional
flabel locali 27680 102 27740 162 1 FreeSans 480 0 0 0 GATE
port 1 n signal bidirectional
<< properties >>
string FIXED_BBOX 0 0 27947 1880
string LEFclass CORE
string LEFsite unitasc
<< end >>
