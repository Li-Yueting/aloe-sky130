magic
tech sky130A
magscale 1 2
timestamp 1653531887
<< pwell >>
rect 140 -60 2580 1650
<< psubdiff >>
rect 1052 940 1668 970
rect 1052 820 1112 940
rect 1608 820 1668 940
rect 1052 790 1668 820
<< psubdiffcont >>
rect 1112 820 1608 940
<< xpolycontact >>
rect 140 1075 572 1645
rect 2148 1075 2580 1645
rect 140 115 572 685
rect 2148 115 2580 685
<< xpolyres >>
rect 572 1075 2148 1645
rect 572 115 2148 685
<< locali >>
rect 140 1850 310 1910
rect 370 1850 510 1910
rect 570 1850 710 1910
rect 770 1850 910 1910
rect 970 1850 1110 1910
rect 1170 1850 1310 1910
rect 1370 1850 1510 1910
rect 1570 1850 1710 1910
rect 1770 1850 1910 1910
rect 1970 1850 2110 1910
rect 2170 1850 2310 1910
rect 2370 1850 2580 1910
rect 1052 940 1668 970
rect 1052 820 1112 940
rect 1608 820 1668 940
rect 1052 30 1668 820
rect 2148 685 2580 1075
rect 140 -30 310 30
rect 370 -30 510 30
rect 570 -30 710 30
rect 770 -30 910 30
rect 970 -30 1110 30
rect 1170 -30 1310 30
rect 1370 -30 1510 30
rect 1570 -30 1710 30
rect 1770 -30 1910 30
rect 1970 -30 2110 30
rect 2170 -30 2310 30
rect 2370 -30 2580 30
<< viali >>
rect 310 1850 370 1910
rect 510 1850 570 1910
rect 710 1850 770 1910
rect 910 1850 970 1910
rect 1110 1850 1170 1910
rect 1310 1850 1370 1910
rect 1510 1850 1570 1910
rect 1710 1850 1770 1910
rect 1910 1850 1970 1910
rect 2110 1850 2170 1910
rect 2310 1850 2370 1910
rect 158 1091 555 1629
rect 2165 1091 2562 1629
rect 158 131 555 669
rect 2165 131 2562 669
rect 310 -30 370 30
rect 510 -30 570 30
rect 710 -30 770 30
rect 910 -30 970 30
rect 1110 -30 1170 30
rect 1310 -30 1370 30
rect 1510 -30 1570 30
rect 1710 -30 1770 30
rect 1910 -30 1970 30
rect 2110 -30 2170 30
rect 2310 -30 2370 30
<< metal1 >>
rect 140 1910 2580 1940
rect 140 1850 310 1910
rect 370 1850 510 1910
rect 570 1850 710 1910
rect 770 1850 910 1910
rect 970 1850 1110 1910
rect 1170 1850 1310 1910
rect 1370 1850 1510 1910
rect 1570 1850 1710 1910
rect 1770 1850 1910 1910
rect 1970 1850 2110 1910
rect 2170 1850 2310 1910
rect 2370 1850 2580 1910
rect 140 1820 2580 1850
rect 151 1629 561 1641
rect 151 1091 158 1629
rect 555 1091 561 1629
rect 151 1079 561 1091
rect 2159 1629 2569 1641
rect 2159 1091 2165 1629
rect 2562 1091 2569 1629
rect 2159 1079 2569 1091
rect 151 669 561 681
rect 151 131 158 669
rect 555 131 561 669
rect 151 119 561 131
rect 2148 669 2580 1079
rect 2148 131 2165 669
rect 2562 131 2580 669
rect 2148 115 2580 131
rect 140 30 2580 60
rect 140 -30 310 30
rect 370 -30 510 30
rect 570 -30 710 30
rect 770 -30 910 30
rect 970 -30 1110 30
rect 1170 -30 1310 30
rect 1370 -30 1510 30
rect 1570 -30 1710 30
rect 1770 -30 1910 30
rect 1970 -30 2110 30
rect 2170 -30 2310 30
rect 2370 -30 2580 30
rect 140 -60 2580 -30
<< labels >>
flabel metal1 260 1300 380 1420 1 FreeSans 480 0 0 0 Rin
port 1 n default bidirectional
flabel metal1 260 340 380 460 1 FreeSans 480 0 0 0 Rout
port 2 n default bidirectional
flabel metal1 140 1850 200 1910 1 FreeSans 800 0 0 0 VPWR
port 3 n power bidirectional
flabel metal1 140 -30 200 30 1 FreeSans 800 0 0 0 VGND
port 4 n ground bidirectional
<< properties >>
string FIXED_BBOX 0 0 2720 1880
string LEFclass CORE
string LEFsite unitasc
<< end >>
