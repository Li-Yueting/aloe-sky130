magic
tech sky130A
magscale 1 2
timestamp 1653339094
<< pwell >>
rect 90 1457 1430 1610
rect 90 423 243 1457
rect 1277 423 1430 1457
rect 90 270 1430 423
<< nbase >>
rect 243 423 1277 1457
<< pdiff >>
rect 420 1228 1100 1280
rect 420 1194 474 1228
rect 508 1194 564 1228
rect 598 1194 654 1228
rect 688 1194 744 1228
rect 778 1194 834 1228
rect 868 1194 924 1228
rect 958 1194 1014 1228
rect 1048 1194 1100 1228
rect 420 1138 1100 1194
rect 420 1104 474 1138
rect 508 1104 564 1138
rect 598 1104 654 1138
rect 688 1104 744 1138
rect 778 1104 834 1138
rect 868 1104 924 1138
rect 958 1104 1014 1138
rect 1048 1104 1100 1138
rect 420 1048 1100 1104
rect 420 1014 474 1048
rect 508 1014 564 1048
rect 598 1014 654 1048
rect 688 1014 744 1048
rect 778 1014 834 1048
rect 868 1014 924 1048
rect 958 1014 1014 1048
rect 1048 1014 1100 1048
rect 420 958 1100 1014
rect 420 924 474 958
rect 508 924 564 958
rect 598 924 654 958
rect 688 924 744 958
rect 778 924 834 958
rect 868 924 924 958
rect 958 924 1014 958
rect 1048 924 1100 958
rect 420 868 1100 924
rect 420 834 474 868
rect 508 834 564 868
rect 598 834 654 868
rect 688 834 744 868
rect 778 834 834 868
rect 868 834 924 868
rect 958 834 1014 868
rect 1048 834 1100 868
rect 420 778 1100 834
rect 420 744 474 778
rect 508 744 564 778
rect 598 744 654 778
rect 688 744 744 778
rect 778 744 834 778
rect 868 744 924 778
rect 958 744 1014 778
rect 1048 744 1100 778
rect 420 688 1100 744
rect 420 654 474 688
rect 508 654 564 688
rect 598 654 654 688
rect 688 654 744 688
rect 778 654 834 688
rect 868 654 924 688
rect 958 654 1014 688
rect 1048 654 1100 688
rect 420 600 1100 654
<< pdiffc >>
rect 474 1194 508 1228
rect 564 1194 598 1228
rect 654 1194 688 1228
rect 744 1194 778 1228
rect 834 1194 868 1228
rect 924 1194 958 1228
rect 1014 1194 1048 1228
rect 474 1104 508 1138
rect 564 1104 598 1138
rect 654 1104 688 1138
rect 744 1104 778 1138
rect 834 1104 868 1138
rect 924 1104 958 1138
rect 1014 1104 1048 1138
rect 474 1014 508 1048
rect 564 1014 598 1048
rect 654 1014 688 1048
rect 744 1014 778 1048
rect 834 1014 868 1048
rect 924 1014 958 1048
rect 1014 1014 1048 1048
rect 474 924 508 958
rect 564 924 598 958
rect 654 924 688 958
rect 744 924 778 958
rect 834 924 868 958
rect 924 924 958 958
rect 1014 924 1048 958
rect 474 834 508 868
rect 564 834 598 868
rect 654 834 688 868
rect 744 834 778 868
rect 834 834 868 868
rect 924 834 958 868
rect 1014 834 1048 868
rect 474 744 508 778
rect 564 744 598 778
rect 654 744 688 778
rect 744 744 778 778
rect 834 744 868 778
rect 924 744 958 778
rect 1014 744 1048 778
rect 474 654 508 688
rect 564 654 598 688
rect 654 654 688 688
rect 744 654 778 688
rect 834 654 868 688
rect 924 654 958 688
rect 1014 654 1048 688
<< psubdiff >>
rect 116 1549 1404 1584
rect 116 1526 246 1549
rect 116 1492 150 1526
rect 184 1515 246 1526
rect 280 1515 336 1549
rect 370 1515 426 1549
rect 460 1515 516 1549
rect 550 1515 606 1549
rect 640 1515 696 1549
rect 730 1515 786 1549
rect 820 1515 876 1549
rect 910 1515 966 1549
rect 1000 1515 1056 1549
rect 1090 1515 1146 1549
rect 1180 1515 1236 1549
rect 1270 1526 1404 1549
rect 1270 1515 1337 1526
rect 184 1492 1337 1515
rect 1371 1492 1404 1526
rect 116 1483 1404 1492
rect 116 1436 217 1483
rect 116 1402 150 1436
rect 184 1402 217 1436
rect 1303 1436 1404 1483
rect 116 1346 217 1402
rect 116 1312 150 1346
rect 184 1312 217 1346
rect 116 1256 217 1312
rect 116 1222 150 1256
rect 184 1222 217 1256
rect 116 1166 217 1222
rect 116 1132 150 1166
rect 184 1132 217 1166
rect 116 1076 217 1132
rect 116 1042 150 1076
rect 184 1042 217 1076
rect 116 986 217 1042
rect 116 952 150 986
rect 184 952 217 986
rect 116 896 217 952
rect 116 862 150 896
rect 184 862 217 896
rect 116 806 217 862
rect 116 772 150 806
rect 184 772 217 806
rect 116 716 217 772
rect 116 682 150 716
rect 184 682 217 716
rect 116 626 217 682
rect 116 592 150 626
rect 184 592 217 626
rect 116 536 217 592
rect 116 502 150 536
rect 184 502 217 536
rect 116 446 217 502
rect 1303 1402 1337 1436
rect 1371 1402 1404 1436
rect 1303 1346 1404 1402
rect 1303 1312 1337 1346
rect 1371 1312 1404 1346
rect 1303 1256 1404 1312
rect 1303 1222 1337 1256
rect 1371 1222 1404 1256
rect 1303 1166 1404 1222
rect 1303 1132 1337 1166
rect 1371 1132 1404 1166
rect 1303 1076 1404 1132
rect 1303 1042 1337 1076
rect 1371 1042 1404 1076
rect 1303 986 1404 1042
rect 1303 952 1337 986
rect 1371 952 1404 986
rect 1303 896 1404 952
rect 1303 862 1337 896
rect 1371 862 1404 896
rect 1303 806 1404 862
rect 1303 772 1337 806
rect 1371 772 1404 806
rect 1303 716 1404 772
rect 1303 682 1337 716
rect 1371 682 1404 716
rect 1303 626 1404 682
rect 1303 592 1337 626
rect 1371 592 1404 626
rect 1303 536 1404 592
rect 1303 502 1337 536
rect 1371 502 1404 536
rect 116 412 150 446
rect 184 412 217 446
rect 116 397 217 412
rect 1303 446 1404 502
rect 1303 412 1337 446
rect 1371 412 1404 446
rect 1303 397 1404 412
rect 116 362 1404 397
rect 116 328 246 362
rect 280 328 336 362
rect 370 328 426 362
rect 460 328 516 362
rect 550 328 606 362
rect 640 328 696 362
rect 730 328 786 362
rect 820 328 876 362
rect 910 328 966 362
rect 1000 328 1056 362
rect 1090 328 1146 362
rect 1180 328 1236 362
rect 1270 328 1404 362
rect 116 296 1404 328
<< nsubdiff >>
rect 279 1402 1241 1421
rect 279 1368 410 1402
rect 444 1368 500 1402
rect 534 1368 590 1402
rect 624 1368 680 1402
rect 714 1368 770 1402
rect 804 1368 860 1402
rect 894 1368 950 1402
rect 984 1368 1040 1402
rect 1074 1368 1130 1402
rect 1164 1368 1241 1402
rect 279 1349 1241 1368
rect 279 1345 351 1349
rect 279 1311 298 1345
rect 332 1311 351 1345
rect 279 1255 351 1311
rect 1169 1326 1241 1349
rect 1169 1292 1188 1326
rect 1222 1292 1241 1326
rect 279 1221 298 1255
rect 332 1221 351 1255
rect 279 1165 351 1221
rect 279 1131 298 1165
rect 332 1131 351 1165
rect 279 1075 351 1131
rect 279 1041 298 1075
rect 332 1041 351 1075
rect 279 985 351 1041
rect 279 951 298 985
rect 332 951 351 985
rect 279 895 351 951
rect 279 861 298 895
rect 332 861 351 895
rect 279 805 351 861
rect 279 771 298 805
rect 332 771 351 805
rect 279 715 351 771
rect 279 681 298 715
rect 332 681 351 715
rect 279 625 351 681
rect 279 591 298 625
rect 332 591 351 625
rect 1169 1236 1241 1292
rect 1169 1202 1188 1236
rect 1222 1202 1241 1236
rect 1169 1146 1241 1202
rect 1169 1112 1188 1146
rect 1222 1112 1241 1146
rect 1169 1056 1241 1112
rect 1169 1022 1188 1056
rect 1222 1022 1241 1056
rect 1169 966 1241 1022
rect 1169 932 1188 966
rect 1222 932 1241 966
rect 1169 876 1241 932
rect 1169 842 1188 876
rect 1222 842 1241 876
rect 1169 786 1241 842
rect 1169 752 1188 786
rect 1222 752 1241 786
rect 1169 696 1241 752
rect 1169 662 1188 696
rect 1222 662 1241 696
rect 1169 606 1241 662
rect 279 531 351 591
rect 1169 572 1188 606
rect 1222 572 1241 606
rect 1169 531 1241 572
rect 279 512 1241 531
rect 279 478 376 512
rect 410 478 466 512
rect 500 478 556 512
rect 590 478 646 512
rect 680 478 736 512
rect 770 478 826 512
rect 860 478 916 512
rect 950 478 1006 512
rect 1040 478 1096 512
rect 1130 478 1241 512
rect 279 459 1241 478
<< psubdiffcont >>
rect 150 1492 184 1526
rect 246 1515 280 1549
rect 336 1515 370 1549
rect 426 1515 460 1549
rect 516 1515 550 1549
rect 606 1515 640 1549
rect 696 1515 730 1549
rect 786 1515 820 1549
rect 876 1515 910 1549
rect 966 1515 1000 1549
rect 1056 1515 1090 1549
rect 1146 1515 1180 1549
rect 1236 1515 1270 1549
rect 1337 1492 1371 1526
rect 150 1402 184 1436
rect 150 1312 184 1346
rect 150 1222 184 1256
rect 150 1132 184 1166
rect 150 1042 184 1076
rect 150 952 184 986
rect 150 862 184 896
rect 150 772 184 806
rect 150 682 184 716
rect 150 592 184 626
rect 150 502 184 536
rect 1337 1402 1371 1436
rect 1337 1312 1371 1346
rect 1337 1222 1371 1256
rect 1337 1132 1371 1166
rect 1337 1042 1371 1076
rect 1337 952 1371 986
rect 1337 862 1371 896
rect 1337 772 1371 806
rect 1337 682 1371 716
rect 1337 592 1371 626
rect 1337 502 1371 536
rect 150 412 184 446
rect 1337 412 1371 446
rect 246 328 280 362
rect 336 328 370 362
rect 426 328 460 362
rect 516 328 550 362
rect 606 328 640 362
rect 696 328 730 362
rect 786 328 820 362
rect 876 328 910 362
rect 966 328 1000 362
rect 1056 328 1090 362
rect 1146 328 1180 362
rect 1236 328 1270 362
<< nsubdiffcont >>
rect 410 1368 444 1402
rect 500 1368 534 1402
rect 590 1368 624 1402
rect 680 1368 714 1402
rect 770 1368 804 1402
rect 860 1368 894 1402
rect 950 1368 984 1402
rect 1040 1368 1074 1402
rect 1130 1368 1164 1402
rect 298 1311 332 1345
rect 1188 1292 1222 1326
rect 298 1221 332 1255
rect 298 1131 332 1165
rect 298 1041 332 1075
rect 298 951 332 985
rect 298 861 332 895
rect 298 771 332 805
rect 298 681 332 715
rect 298 591 332 625
rect 1188 1202 1222 1236
rect 1188 1112 1222 1146
rect 1188 1022 1222 1056
rect 1188 932 1222 966
rect 1188 842 1222 876
rect 1188 752 1222 786
rect 1188 662 1222 696
rect 1188 572 1222 606
rect 376 478 410 512
rect 466 478 500 512
rect 556 478 590 512
rect 646 478 680 512
rect 736 478 770 512
rect 826 478 860 512
rect 916 478 950 512
rect 1006 478 1040 512
rect 1096 478 1130 512
<< locali >>
rect 90 1850 260 1910
rect 320 1850 460 1910
rect 520 1850 660 1910
rect 720 1850 860 1910
rect 920 1850 1060 1910
rect 1120 1850 1260 1910
rect 1320 1850 1430 1910
rect 116 1549 1404 1584
rect 116 1526 246 1549
rect 116 1492 150 1526
rect 184 1515 246 1526
rect 280 1515 336 1549
rect 370 1515 426 1549
rect 460 1515 516 1549
rect 550 1515 606 1549
rect 640 1515 696 1549
rect 730 1515 786 1549
rect 820 1515 876 1549
rect 910 1515 966 1549
rect 1000 1515 1056 1549
rect 1090 1515 1146 1549
rect 1180 1515 1236 1549
rect 1270 1526 1404 1549
rect 1270 1515 1337 1526
rect 184 1492 1337 1515
rect 1371 1492 1404 1526
rect 116 1485 1404 1492
rect 116 1436 215 1485
rect 116 1402 150 1436
rect 184 1402 215 1436
rect 1305 1436 1404 1485
rect 116 1346 215 1402
rect 116 1312 150 1346
rect 184 1312 215 1346
rect 116 1256 215 1312
rect 116 1222 150 1256
rect 184 1222 215 1256
rect 116 1166 215 1222
rect 116 1132 150 1166
rect 184 1132 215 1166
rect 116 1076 215 1132
rect 116 1042 150 1076
rect 184 1042 215 1076
rect 116 986 215 1042
rect 116 952 150 986
rect 184 952 215 986
rect 116 896 215 952
rect 116 862 150 896
rect 184 862 215 896
rect 116 806 215 862
rect 116 772 150 806
rect 184 772 215 806
rect 116 716 215 772
rect 116 682 150 716
rect 184 682 215 716
rect 116 626 215 682
rect 116 592 150 626
rect 184 592 215 626
rect 116 536 215 592
rect 116 502 150 536
rect 184 502 215 536
rect 116 446 215 502
rect 279 1402 1241 1421
rect 279 1368 410 1402
rect 444 1368 500 1402
rect 534 1368 590 1402
rect 624 1368 680 1402
rect 714 1368 770 1402
rect 804 1368 860 1402
rect 894 1368 950 1402
rect 984 1368 1040 1402
rect 1074 1368 1130 1402
rect 1164 1368 1241 1402
rect 279 1349 1241 1368
rect 279 1345 351 1349
rect 279 1311 298 1345
rect 332 1311 351 1345
rect 279 1255 351 1311
rect 1169 1326 1241 1349
rect 1169 1292 1188 1326
rect 1222 1292 1241 1326
rect 279 1221 298 1255
rect 332 1221 351 1255
rect 279 1165 351 1221
rect 279 1131 298 1165
rect 332 1131 351 1165
rect 279 1075 351 1131
rect 279 1041 298 1075
rect 332 1041 351 1075
rect 279 985 351 1041
rect 279 951 298 985
rect 332 951 351 985
rect 279 895 351 951
rect 279 861 298 895
rect 332 861 351 895
rect 279 805 351 861
rect 279 771 298 805
rect 332 771 351 805
rect 279 715 351 771
rect 279 681 298 715
rect 332 681 351 715
rect 279 625 351 681
rect 279 591 298 625
rect 332 591 351 625
rect 413 1228 1107 1287
rect 413 1194 474 1228
rect 508 1200 564 1228
rect 598 1200 654 1228
rect 688 1200 744 1228
rect 520 1194 564 1200
rect 620 1194 654 1200
rect 720 1194 744 1200
rect 778 1200 834 1228
rect 778 1194 786 1200
rect 413 1166 486 1194
rect 520 1166 586 1194
rect 620 1166 686 1194
rect 720 1166 786 1194
rect 820 1194 834 1200
rect 868 1200 924 1228
rect 868 1194 886 1200
rect 820 1166 886 1194
rect 920 1194 924 1200
rect 958 1200 1014 1228
rect 958 1194 986 1200
rect 1048 1194 1107 1228
rect 920 1166 986 1194
rect 1020 1166 1107 1194
rect 413 1138 1107 1166
rect 413 1104 474 1138
rect 508 1104 564 1138
rect 598 1104 654 1138
rect 688 1104 744 1138
rect 778 1104 834 1138
rect 868 1104 924 1138
rect 958 1104 1014 1138
rect 1048 1104 1107 1138
rect 413 1100 1107 1104
rect 413 1066 486 1100
rect 520 1066 586 1100
rect 620 1066 686 1100
rect 720 1066 786 1100
rect 820 1066 886 1100
rect 920 1066 986 1100
rect 1020 1066 1107 1100
rect 413 1048 1107 1066
rect 413 1014 474 1048
rect 508 1014 564 1048
rect 598 1014 654 1048
rect 688 1014 744 1048
rect 778 1014 834 1048
rect 868 1014 924 1048
rect 958 1014 1014 1048
rect 1048 1014 1107 1048
rect 413 1000 1107 1014
rect 413 966 486 1000
rect 520 966 586 1000
rect 620 966 686 1000
rect 720 966 786 1000
rect 820 966 886 1000
rect 920 966 986 1000
rect 1020 966 1107 1000
rect 413 958 1107 966
rect 413 924 474 958
rect 508 924 564 958
rect 598 924 654 958
rect 688 924 744 958
rect 778 924 834 958
rect 868 924 924 958
rect 958 924 1014 958
rect 1048 924 1107 958
rect 413 900 1107 924
rect 413 868 486 900
rect 520 868 586 900
rect 620 868 686 900
rect 720 868 786 900
rect 413 834 474 868
rect 520 866 564 868
rect 620 866 654 868
rect 720 866 744 868
rect 508 834 564 866
rect 598 834 654 866
rect 688 834 744 866
rect 778 866 786 868
rect 820 868 886 900
rect 820 866 834 868
rect 778 834 834 866
rect 868 866 886 868
rect 920 868 986 900
rect 1020 868 1107 900
rect 920 866 924 868
rect 868 834 924 866
rect 958 866 986 868
rect 958 834 1014 866
rect 1048 834 1107 868
rect 413 800 1107 834
rect 413 778 486 800
rect 520 778 586 800
rect 620 778 686 800
rect 720 778 786 800
rect 413 744 474 778
rect 520 766 564 778
rect 620 766 654 778
rect 720 766 744 778
rect 508 744 564 766
rect 598 744 654 766
rect 688 744 744 766
rect 778 766 786 778
rect 820 778 886 800
rect 820 766 834 778
rect 778 744 834 766
rect 868 766 886 778
rect 920 778 986 800
rect 1020 778 1107 800
rect 920 766 924 778
rect 868 744 924 766
rect 958 766 986 778
rect 958 744 1014 766
rect 1048 744 1107 778
rect 413 700 1107 744
rect 413 688 486 700
rect 520 688 586 700
rect 620 688 686 700
rect 720 688 786 700
rect 413 654 474 688
rect 520 666 564 688
rect 620 666 654 688
rect 720 666 744 688
rect 508 654 564 666
rect 598 654 654 666
rect 688 654 744 666
rect 778 666 786 688
rect 820 688 886 700
rect 820 666 834 688
rect 778 654 834 666
rect 868 666 886 688
rect 920 688 986 700
rect 1020 688 1107 700
rect 920 666 924 688
rect 868 654 924 666
rect 958 666 986 688
rect 958 654 1014 666
rect 1048 654 1107 688
rect 413 593 1107 654
rect 1169 1236 1241 1292
rect 1169 1202 1188 1236
rect 1222 1202 1241 1236
rect 1169 1146 1241 1202
rect 1169 1112 1188 1146
rect 1222 1112 1241 1146
rect 1169 1056 1241 1112
rect 1169 1022 1188 1056
rect 1222 1022 1241 1056
rect 1169 966 1241 1022
rect 1169 932 1188 966
rect 1222 932 1241 966
rect 1169 876 1241 932
rect 1169 842 1188 876
rect 1222 842 1241 876
rect 1169 786 1241 842
rect 1169 752 1188 786
rect 1222 752 1241 786
rect 1169 696 1241 752
rect 1169 662 1188 696
rect 1222 662 1241 696
rect 1169 606 1241 662
rect 279 531 351 591
rect 1169 572 1188 606
rect 1222 572 1241 606
rect 1169 531 1241 572
rect 279 512 1241 531
rect 279 478 376 512
rect 410 478 466 512
rect 500 478 556 512
rect 590 478 646 512
rect 680 478 736 512
rect 770 478 826 512
rect 860 478 916 512
rect 958 478 1006 512
rect 1040 478 1096 512
rect 1130 478 1241 512
rect 279 459 1241 478
rect 1305 1402 1337 1436
rect 1371 1402 1404 1436
rect 1305 1346 1404 1402
rect 1305 1312 1337 1346
rect 1371 1312 1404 1346
rect 1305 1256 1404 1312
rect 1305 1222 1337 1256
rect 1371 1222 1404 1256
rect 1305 1166 1404 1222
rect 1305 1132 1337 1166
rect 1371 1132 1404 1166
rect 1305 1076 1404 1132
rect 1305 1042 1337 1076
rect 1371 1042 1404 1076
rect 1305 986 1404 1042
rect 1305 952 1337 986
rect 1371 952 1404 986
rect 1305 896 1404 952
rect 1305 862 1337 896
rect 1371 862 1404 896
rect 1305 806 1404 862
rect 1305 772 1337 806
rect 1371 772 1404 806
rect 1305 716 1404 772
rect 1305 682 1337 716
rect 1371 682 1404 716
rect 1305 626 1404 682
rect 1305 592 1337 626
rect 1371 592 1404 626
rect 1305 536 1404 592
rect 1305 502 1337 536
rect 1371 502 1404 536
rect 116 412 150 446
rect 184 412 215 446
rect 116 395 215 412
rect 1305 446 1404 502
rect 1305 412 1337 446
rect 1371 412 1404 446
rect 1305 395 1404 412
rect 116 362 1404 395
rect 116 328 246 362
rect 280 328 336 362
rect 370 328 426 362
rect 460 328 516 362
rect 550 328 606 362
rect 640 328 696 362
rect 730 328 786 362
rect 820 328 876 362
rect 910 352 966 362
rect 910 328 922 352
rect 116 318 922 328
rect 958 328 966 352
rect 1000 328 1056 362
rect 1090 328 1146 362
rect 1180 328 1236 362
rect 1270 328 1404 362
rect 958 318 1404 328
rect 116 296 1404 318
rect 90 -30 260 30
rect 320 -30 460 30
rect 520 -30 660 30
rect 720 -30 860 30
rect 920 -30 1060 30
rect 1120 -30 1260 30
rect 1320 -30 1430 30
<< viali >>
rect 260 1850 320 1910
rect 460 1850 520 1910
rect 660 1850 720 1910
rect 860 1850 920 1910
rect 1060 1850 1120 1910
rect 1260 1850 1320 1910
rect 486 1194 508 1200
rect 508 1194 520 1200
rect 586 1194 598 1200
rect 598 1194 620 1200
rect 686 1194 688 1200
rect 688 1194 720 1200
rect 486 1166 520 1194
rect 586 1166 620 1194
rect 686 1166 720 1194
rect 786 1166 820 1200
rect 886 1166 920 1200
rect 986 1194 1014 1200
rect 1014 1194 1020 1200
rect 986 1166 1020 1194
rect 486 1066 520 1100
rect 586 1066 620 1100
rect 686 1066 720 1100
rect 786 1066 820 1100
rect 886 1066 920 1100
rect 986 1066 1020 1100
rect 486 966 520 1000
rect 586 966 620 1000
rect 686 966 720 1000
rect 786 966 820 1000
rect 886 966 920 1000
rect 986 966 1020 1000
rect 486 868 520 900
rect 586 868 620 900
rect 686 868 720 900
rect 486 866 508 868
rect 508 866 520 868
rect 586 866 598 868
rect 598 866 620 868
rect 686 866 688 868
rect 688 866 720 868
rect 786 866 820 900
rect 886 866 920 900
rect 986 868 1020 900
rect 986 866 1014 868
rect 1014 866 1020 868
rect 486 778 520 800
rect 586 778 620 800
rect 686 778 720 800
rect 486 766 508 778
rect 508 766 520 778
rect 586 766 598 778
rect 598 766 620 778
rect 686 766 688 778
rect 688 766 720 778
rect 786 766 820 800
rect 886 766 920 800
rect 986 778 1020 800
rect 986 766 1014 778
rect 1014 766 1020 778
rect 486 688 520 700
rect 586 688 620 700
rect 686 688 720 700
rect 486 666 508 688
rect 508 666 520 688
rect 586 666 598 688
rect 598 666 620 688
rect 686 666 688 688
rect 688 666 720 688
rect 786 666 820 700
rect 886 666 920 700
rect 986 688 1020 700
rect 986 666 1014 688
rect 1014 666 1020 688
rect 922 478 950 512
rect 950 478 958 512
rect 922 318 958 352
rect 260 -30 320 30
rect 460 -30 520 30
rect 660 -30 720 30
rect 860 -30 920 30
rect 1060 -30 1120 30
rect 1260 -30 1320 30
<< metal1 >>
rect 90 1910 1430 1940
rect 90 1850 260 1910
rect 320 1850 460 1910
rect 520 1850 660 1910
rect 720 1850 860 1910
rect 920 1850 1060 1910
rect 1120 1850 1260 1910
rect 1320 1850 1430 1910
rect 90 1820 1430 1850
rect 455 1200 1065 1245
rect 455 1166 486 1200
rect 520 1166 586 1200
rect 620 1166 686 1200
rect 720 1166 786 1200
rect 820 1166 886 1200
rect 920 1166 986 1200
rect 1020 1166 1065 1200
rect 455 1100 1065 1166
rect 455 1066 486 1100
rect 520 1066 586 1100
rect 620 1066 686 1100
rect 720 1066 786 1100
rect 820 1066 886 1100
rect 920 1066 986 1100
rect 1020 1066 1065 1100
rect 455 1000 1065 1066
rect 455 966 486 1000
rect 520 966 586 1000
rect 620 966 686 1000
rect 720 966 786 1000
rect 820 966 886 1000
rect 920 966 986 1000
rect 1020 966 1065 1000
rect 455 900 1065 966
rect 455 866 486 900
rect 520 866 586 900
rect 620 866 686 900
rect 720 866 786 900
rect 820 866 886 900
rect 920 866 986 900
rect 1020 866 1065 900
rect 455 800 1065 866
rect 455 766 486 800
rect 520 766 586 800
rect 620 766 686 800
rect 720 766 786 800
rect 820 766 886 800
rect 920 766 986 800
rect 1020 766 1065 800
rect 455 700 1065 766
rect 455 666 486 700
rect 520 666 586 700
rect 620 666 686 700
rect 720 666 786 700
rect 820 666 886 700
rect 920 666 986 700
rect 1020 666 1065 700
rect 455 635 1065 666
rect 878 512 1108 522
rect 878 478 922 512
rect 958 478 1108 512
rect 878 462 1108 478
rect 878 352 1108 384
rect 878 318 922 352
rect 958 318 1108 352
rect 878 302 1108 318
rect 90 30 1430 60
rect 90 -30 260 30
rect 320 -30 460 30
rect 520 -30 660 30
rect 720 -30 860 30
rect 920 -30 1060 30
rect 1120 -30 1260 30
rect 1320 -30 1430 30
rect 90 -60 1430 -30
<< pnp3p40 >>
rect 243 423 1277 1457
<< labels >>
flabel metal1 878 302 1108 384 1 FreeSans 480 0 0 0 Collector
port 3 n default bidirectional
flabel metal1 878 462 1108 522 1 FreeSans 480 0 0 0 Base
port 2 n default bidirectional
flabel locali 652 1010 880 1140 1 FreeSans 480 0 0 0 Emitter
port 1 n default bidirectional
flabel metal1 90 1850 150 1910 1 FreeSans 800 0 0 0 VPWR
port 4 n power bidirectional
flabel metal1 90 -30 150 30 1 FreeSans 800 0 0 0 VGND
port 5 n ground bidirectional
flabel locali 644 896 892 1000 0 FreeSans 400 0 0 0 xm2/Emitter
flabel locali 703 1522 804 1571 0 FreeSans 400 0 0 0 xm2/Collector
flabel locali 680 1372 798 1412 0 FreeSans 400 0 0 0 xm2/Base
<< properties >>
string FIXED_BBOX 0 0 1520 1880
string LEFclass CORE
string LEFsite unitasc
<< end >>
