VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO sky130_asc_cap_mim_m3_1
  CLASS CORE ;
  FOREIGN sky130_asc_cap_mim_m3_1 ;
  ORIGIN 0.000 0.000 ;
  SIZE 37.055 BY 9.400 ;
  SITE unitasc ;
  PIN Cin
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 0.600 7.850 1.600 8.250 ;
    END
  END Cin
  PIN Cout
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 0.710 0.700 1.510 1.200 ;
    END
  END Cout
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER li1 ;
        RECT 0.610 9.250 36.450 9.550 ;
      LAYER mcon ;
        RECT 1.460 9.250 1.760 9.550 ;
        RECT 3.460 9.250 3.760 9.550 ;
        RECT 5.460 9.250 5.760 9.550 ;
        RECT 7.460 9.250 7.760 9.550 ;
        RECT 9.460 9.250 9.760 9.550 ;
        RECT 11.460 9.250 11.760 9.550 ;
        RECT 13.460 9.250 13.760 9.550 ;
        RECT 15.460 9.250 15.760 9.550 ;
        RECT 17.460 9.250 17.760 9.550 ;
        RECT 19.460 9.250 19.760 9.550 ;
        RECT 21.460 9.250 21.760 9.550 ;
        RECT 23.460 9.250 23.760 9.550 ;
        RECT 25.460 9.250 25.760 9.550 ;
        RECT 27.460 9.250 27.760 9.550 ;
        RECT 29.460 9.250 29.760 9.550 ;
        RECT 31.460 9.250 31.760 9.550 ;
        RECT 33.460 9.250 33.760 9.550 ;
        RECT 35.460 9.250 35.760 9.550 ;
      LAYER met1 ;
        RECT 0.610 9.100 36.450 9.700 ;
    END
  END VPWR
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER li1 ;
        RECT 0.610 -0.150 36.450 0.150 ;
      LAYER mcon ;
        RECT 1.460 -0.150 1.760 0.150 ;
        RECT 3.460 -0.150 3.760 0.150 ;
        RECT 5.460 -0.150 5.760 0.150 ;
        RECT 7.460 -0.150 7.760 0.150 ;
        RECT 9.460 -0.150 9.760 0.150 ;
        RECT 11.460 -0.150 11.760 0.150 ;
        RECT 13.460 -0.150 13.760 0.150 ;
        RECT 15.460 -0.150 15.760 0.150 ;
        RECT 17.460 -0.150 17.760 0.150 ;
        RECT 19.460 -0.150 19.760 0.150 ;
        RECT 21.460 -0.150 21.760 0.150 ;
        RECT 23.460 -0.150 23.760 0.150 ;
        RECT 25.460 -0.150 25.760 0.150 ;
        RECT 27.460 -0.150 27.760 0.150 ;
        RECT 29.460 -0.150 29.760 0.150 ;
        RECT 31.460 -0.150 31.760 0.150 ;
        RECT 33.460 -0.150 33.760 0.150 ;
        RECT 35.460 -0.150 35.760 0.150 ;
      LAYER met1 ;
        RECT 0.610 -0.300 36.450 0.300 ;
    END
  END VGND
  OBS
      LAYER met3 ;
        RECT 0.600 1.750 37 8.250 ;
      LAYER met4 ;
        RECT 0.4 0.500 36.830 8.870 ;
      LAYER met5 ;
        RECT 0.4 0.500 36.830 8.870 ;
  END
END sky130_asc_cap_mim_m3_1
END LIBRARY

