VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO sky130_asc_nfet_01v8_lvt_1
  CLASS CORE ;
  FOREIGN sky130_asc_nfet_01v8_lvt_1 ;
  ORIGIN 0.000 0.000 ;
  SIZE 4.270 BY 9.400 ;
  SITE unitasc ;
  PIN GATE
    DIRECTION INOUT ;
    ANTENNAGATEAREA 8.000000 ;
    PORT
      LAYER li1 ;
        RECT 0.600 0.570 3.180 0.870 ;
    END
  END GATE
  PIN SOURCE
    DIRECTION INOUT ;
    ANTENNADIFFAREA 1.160000 ;
    PORT
      LAYER li1 ;
        RECT 0.600 5.950 3.180 6.250 ;
        RECT 2.945 5.670 3.115 5.950 ;
        RECT 2.945 5.380 3.120 5.670 ;
        RECT 2.950 1.630 3.120 5.380 ;
      LAYER mcon ;
        RECT 2.950 1.710 3.120 5.590 ;
      LAYER met1 ;
        RECT 2.920 1.650 3.150 5.650 ;
    END
  END SOURCE
  PIN DRAIN
    DIRECTION INOUT ;
    ANTENNADIFFAREA 1.160000 ;
    PORT
      LAYER li1 ;
        RECT 0.660 1.920 0.830 5.670 ;
        RECT 0.655 1.630 0.830 1.920 ;
        RECT 0.655 1.350 0.825 1.630 ;
        RECT 0.600 1.050 3.180 1.350 ;
      LAYER mcon ;
        RECT 0.660 1.710 0.830 5.590 ;
      LAYER met1 ;
        RECT 0.630 1.650 0.860 5.650 ;
    END
  END DRAIN
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER li1 ;
        RECT 0.600 6.550 3.180 6.850 ;
      LAYER mcon ;
        RECT 1.450 6.550 1.750 6.850 ;
      LAYER met1 ;
        RECT 0.600 6.400 3.180 7.000 ;
    END
  END VPWR
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER li1 ;
        RECT 0.600 -0.150 3.180 0.150 ;
      LAYER mcon ;
        RECT 1.450 -0.150 1.750 0.150 ;
      LAYER met1 ;
        RECT 0.600 -0.300 3.180 0.300 ;
    END
  END VGND
  OBS
      LAYER pwell ;
        RECT 0.600 0.150 3.180 3.650 ;
  END
END sky130_asc_nfet_01v8_lvt_1
END LIBRARY

