VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO sky130_asc_cap_mim_m3_1
  CLASS CORE ;
  FOREIGN sky130_asc_cap_mim_m3_1 ;
  ORIGIN 0.000 0.000 ;
  SIZE 35.855 BY 9.400 ;
  SITE unitasc ;
  PIN Cin
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 8.250 35.850 8.450 ;
        RECT 0.000 5.250 35.855 8.250 ;
        RECT 0.000 4.750 35.850 5.250 ;
        RECT 0.000 1.750 35.855 4.750 ;
      LAYER via3 ;
        RECT 3.080 5.390 3.400 8.110 ;
        RECT 6.675 5.390 6.995 8.110 ;
        RECT 10.270 5.390 10.590 8.110 ;
        RECT 13.865 5.390 14.185 8.110 ;
        RECT 17.460 5.390 17.780 8.110 ;
        RECT 21.055 5.390 21.375 8.110 ;
        RECT 24.650 5.390 24.970 8.110 ;
        RECT 28.245 5.390 28.565 8.110 ;
        RECT 31.840 5.390 32.160 8.110 ;
        RECT 35.435 5.390 35.755 8.110 ;
        RECT 3.080 1.890 3.400 4.610 ;
        RECT 6.675 1.890 6.995 4.610 ;
        RECT 10.270 1.890 10.590 4.610 ;
        RECT 13.865 1.890 14.185 4.610 ;
        RECT 17.460 1.890 17.780 4.610 ;
        RECT 21.055 1.890 21.375 4.610 ;
        RECT 24.650 1.890 24.970 4.610 ;
        RECT 28.245 1.890 28.565 4.610 ;
        RECT 31.840 1.890 32.160 4.610 ;
        RECT 35.435 1.890 35.755 4.610 ;
      LAYER met4 ;
        RECT 3.000 5.310 3.480 8.190 ;
        RECT 6.595 5.310 7.075 8.190 ;
        RECT 10.190 5.310 10.670 8.190 ;
        RECT 13.785 5.310 14.265 8.190 ;
        RECT 17.380 5.310 17.860 8.190 ;
        RECT 20.975 5.310 21.455 8.190 ;
        RECT 24.570 5.310 25.050 8.190 ;
        RECT 28.165 5.310 28.645 8.190 ;
        RECT 31.760 5.310 32.240 8.190 ;
        RECT 35.355 5.310 35.835 8.190 ;
        RECT 3.000 1.810 3.480 4.690 ;
        RECT 6.595 1.810 7.075 4.690 ;
        RECT 10.190 1.810 10.670 4.690 ;
        RECT 13.785 1.810 14.265 4.690 ;
        RECT 17.380 1.810 17.860 4.690 ;
        RECT 20.975 1.810 21.455 4.690 ;
        RECT 24.570 1.810 25.050 4.690 ;
        RECT 28.165 1.810 28.645 4.690 ;
        RECT 31.760 1.810 32.240 4.690 ;
        RECT 35.355 1.810 35.835 4.690 ;
    END
  END Cin
  PIN Cout
    DIRECTION INOUT ;
    PORT
      LAYER met4 ;
        RECT 0.700 7.555 2.300 7.650 ;
        RECT 4.300 7.555 5.900 7.650 ;
        RECT 7.900 7.555 9.500 7.650 ;
        RECT 11.500 7.555 13.100 7.650 ;
        RECT 15.100 7.555 16.700 7.650 ;
        RECT 18.700 7.555 20.300 7.650 ;
        RECT 22.300 7.555 23.900 7.650 ;
        RECT 25.900 7.555 27.500 7.650 ;
        RECT 29.500 7.555 31.100 7.650 ;
        RECT 33.100 7.555 34.700 7.650 ;
        RECT 0.700 5.945 2.310 7.555 ;
        RECT 4.295 5.945 5.905 7.555 ;
        RECT 7.890 5.945 9.500 7.555 ;
        RECT 11.485 5.945 13.100 7.555 ;
        RECT 15.080 5.945 16.700 7.555 ;
        RECT 18.675 5.945 20.300 7.555 ;
        RECT 22.270 5.945 23.900 7.555 ;
        RECT 25.865 5.945 27.500 7.555 ;
        RECT 29.460 5.945 31.100 7.555 ;
        RECT 33.055 5.945 34.700 7.555 ;
        RECT 0.700 4.055 2.300 5.945 ;
        RECT 4.300 4.055 5.900 5.945 ;
        RECT 7.900 4.055 9.500 5.945 ;
        RECT 11.500 4.055 13.100 5.945 ;
        RECT 15.100 4.055 16.700 5.945 ;
        RECT 18.700 4.055 20.300 5.945 ;
        RECT 22.300 4.055 23.900 5.945 ;
        RECT 25.900 4.055 27.500 5.945 ;
        RECT 29.500 4.055 31.100 5.945 ;
        RECT 33.100 4.055 34.700 5.945 ;
        RECT 0.700 2.445 2.310 4.055 ;
        RECT 4.295 2.445 5.905 4.055 ;
        RECT 7.890 2.445 9.500 4.055 ;
        RECT 11.485 2.445 13.100 4.055 ;
        RECT 15.080 2.445 16.700 4.055 ;
        RECT 18.675 2.445 20.300 4.055 ;
        RECT 22.270 2.445 23.900 4.055 ;
        RECT 25.865 2.445 27.500 4.055 ;
        RECT 29.460 2.445 31.100 4.055 ;
        RECT 33.055 2.445 34.700 4.055 ;
        RECT 0.700 1.450 2.300 2.445 ;
        RECT 4.300 1.450 5.900 2.445 ;
        RECT 7.900 1.450 9.500 2.445 ;
        RECT 11.500 1.450 13.100 2.445 ;
        RECT 15.100 1.450 16.700 2.445 ;
        RECT 18.700 1.450 20.300 2.445 ;
        RECT 22.300 1.450 23.900 2.445 ;
        RECT 25.900 1.450 27.500 2.445 ;
        RECT 29.500 1.450 31.100 2.445 ;
        RECT 33.100 1.450 34.700 2.445 ;
        RECT 0.010 0.950 35.850 1.450 ;
    END
  END Cout
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER li1 ;
        RECT 0.010 9.250 35.850 9.550 ;
      LAYER mcon ;
        RECT 0.860 9.250 1.160 9.550 ;
        RECT 2.860 9.250 3.160 9.550 ;
        RECT 4.860 9.250 5.160 9.550 ;
        RECT 6.860 9.250 7.160 9.550 ;
        RECT 8.860 9.250 9.160 9.550 ;
        RECT 10.860 9.250 11.160 9.550 ;
        RECT 12.860 9.250 13.160 9.550 ;
        RECT 14.860 9.250 15.160 9.550 ;
        RECT 16.860 9.250 17.160 9.550 ;
        RECT 18.860 9.250 19.160 9.550 ;
        RECT 20.860 9.250 21.160 9.550 ;
        RECT 22.860 9.250 23.160 9.550 ;
        RECT 24.860 9.250 25.160 9.550 ;
        RECT 26.860 9.250 27.160 9.550 ;
        RECT 28.860 9.250 29.160 9.550 ;
        RECT 30.860 9.250 31.160 9.550 ;
        RECT 32.860 9.250 33.160 9.550 ;
        RECT 34.860 9.250 35.160 9.550 ;
      LAYER met1 ;
        RECT 0.010 9.100 35.850 9.700 ;
    END
  END VPWR
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER li1 ;
        RECT 0.010 -0.150 35.850 0.150 ;
      LAYER mcon ;
        RECT 0.860 -0.150 1.160 0.150 ;
        RECT 2.860 -0.150 3.160 0.150 ;
        RECT 4.860 -0.150 5.160 0.150 ;
        RECT 6.860 -0.150 7.160 0.150 ;
        RECT 8.860 -0.150 9.160 0.150 ;
        RECT 10.860 -0.150 11.160 0.150 ;
        RECT 12.860 -0.150 13.160 0.150 ;
        RECT 14.860 -0.150 15.160 0.150 ;
        RECT 16.860 -0.150 17.160 0.150 ;
        RECT 18.860 -0.150 19.160 0.150 ;
        RECT 20.860 -0.150 21.160 0.150 ;
        RECT 22.860 -0.150 23.160 0.150 ;
        RECT 24.860 -0.150 25.160 0.150 ;
        RECT 26.860 -0.150 27.160 0.150 ;
        RECT 28.860 -0.150 29.160 0.150 ;
        RECT 30.860 -0.150 31.160 0.150 ;
        RECT 32.860 -0.150 33.160 0.150 ;
        RECT 34.860 -0.150 35.160 0.150 ;
      LAYER met1 ;
        RECT 0.010 -0.300 35.850 0.300 ;
    END
  END VGND
END sky130_asc_cap_mim_m3_1
END LIBRARY

