//-----------------------------------------------------------------------------
// BGR  
//-----------------------------------------------------------------------------
module bgr_0 (
  `ifdef USE_POWER_PINS
    inout VDD,
    inout VSS,
	`endif
    inout porst,
    inout va, 
    inout vb,
    inout vbg
 );
  // supply1 VDD;
  // supply0 VSS;
endmodule

